magic
tech sky130l
timestamp 1731220575
<< m1 >>
rect 152 3435 156 3483
rect 1272 3435 1276 3483
rect 1520 3447 1524 3483
rect 2816 3435 2820 3491
rect 3192 3455 3196 3491
rect 936 3335 940 3431
rect 3336 3399 3340 3431
rect 552 3295 556 3331
rect 1384 3279 1388 3331
rect 1528 3295 1532 3331
rect 656 3243 660 3275
rect 1480 3243 1484 3275
rect 2824 3267 2828 3327
rect 3080 3291 3084 3327
rect 3000 2947 3004 2983
rect 672 2827 676 2863
rect 2352 2787 2356 2823
rect 2464 2787 2468 2823
rect 704 2671 708 2707
rect 2216 2667 2220 2763
rect 2312 2627 2316 2663
rect 1128 2463 1132 2495
rect 2104 2247 2108 2279
rect 2248 2247 2252 2279
rect 3088 2275 3092 2287
rect 3496 2283 3500 2331
rect 144 2139 148 2187
rect 2848 2099 2852 2159
rect 496 2019 500 2067
rect 1096 2019 1100 2059
rect 680 1823 684 1855
rect 1128 1823 1132 1855
rect 2112 1803 2116 1819
rect 1520 1663 1524 1695
rect 128 1431 132 1531
rect 3480 1459 3484 1511
rect 3488 1475 3492 1671
rect 128 1259 132 1359
rect 1384 1327 1388 1359
rect 1600 1259 1604 1359
rect 2416 1319 2420 1391
rect 2520 1259 2524 1291
rect 208 1227 212 1255
rect 128 1099 132 1195
rect 3488 1191 3492 1291
rect 360 1035 364 1087
rect 768 1035 772 1087
rect 1888 1031 1892 1127
rect 2264 1095 2268 1127
rect 3496 1031 3500 1127
rect 128 923 132 1031
rect 2480 975 2484 1027
rect 2632 975 2636 1027
rect 3344 975 3348 1027
rect 256 883 260 967
rect 960 867 964 919
rect 1216 883 1220 967
rect 752 831 756 863
rect 1888 831 1892 971
rect 3496 863 3500 971
rect 1904 811 1908 859
rect 2168 823 2172 859
rect 2552 811 2556 859
rect 2560 823 2564 859
rect 3496 711 3500 807
rect 2592 671 2596 707
rect 2736 659 2740 699
rect 952 547 956 627
rect 3184 559 3188 655
rect 2352 463 2356 495
rect 536 351 540 411
rect 648 375 652 411
rect 752 375 756 455
rect 128 243 132 347
rect 2232 339 2236 383
rect 2328 355 2332 391
rect 3488 355 3492 431
rect 648 203 652 239
rect 2624 171 2628 231
rect 1248 119 1252 151
rect 1488 119 1492 151
<< m2c >>
rect 136 3595 140 3599
rect 216 3595 220 3599
rect 2056 3591 2060 3595
rect 2144 3591 2148 3595
rect 2248 3591 2252 3595
rect 2360 3591 2364 3595
rect 2472 3591 2476 3595
rect 2584 3591 2588 3595
rect 2696 3591 2700 3595
rect 2808 3591 2812 3595
rect 2912 3591 2916 3595
rect 3008 3591 3012 3595
rect 3104 3591 3108 3595
rect 3200 3591 3204 3595
rect 3296 3591 3300 3595
rect 3392 3591 3396 3595
rect 136 3583 140 3587
rect 216 3583 220 3587
rect 336 3583 340 3587
rect 464 3583 468 3587
rect 600 3583 604 3587
rect 736 3583 740 3587
rect 872 3583 876 3587
rect 992 3583 996 3587
rect 1104 3583 1108 3587
rect 1216 3583 1220 3587
rect 1320 3583 1324 3587
rect 1416 3583 1420 3587
rect 1520 3583 1524 3587
rect 1624 3583 1628 3587
rect 2600 3527 2604 3531
rect 3408 3527 3412 3531
rect 1640 3519 1644 3523
rect 2816 3491 2820 3495
rect 152 3483 156 3487
rect 1272 3483 1276 3487
rect 192 3443 196 3447
rect 328 3443 332 3447
rect 472 3443 476 3447
rect 624 3443 628 3447
rect 776 3443 780 3447
rect 920 3443 924 3447
rect 1056 3443 1060 3447
rect 1184 3443 1188 3447
rect 1520 3483 1524 3487
rect 2088 3451 2092 3455
rect 2168 3451 2172 3455
rect 2264 3451 2268 3455
rect 2368 3451 2372 3455
rect 2488 3451 2492 3455
rect 2616 3451 2620 3455
rect 2744 3451 2748 3455
rect 1312 3443 1316 3447
rect 1440 3443 1444 3447
rect 1520 3443 1524 3447
rect 1568 3443 1572 3447
rect 3192 3491 3196 3495
rect 2872 3451 2876 3455
rect 2992 3451 2996 3455
rect 3120 3451 3124 3455
rect 3192 3451 3196 3455
rect 3248 3451 3252 3455
rect 3376 3451 3380 3455
rect 144 3431 148 3435
rect 152 3431 156 3435
rect 288 3431 292 3435
rect 448 3431 452 3435
rect 616 3431 620 3435
rect 784 3431 788 3435
rect 936 3431 940 3435
rect 952 3431 956 3435
rect 1112 3431 1116 3435
rect 1264 3431 1268 3435
rect 1272 3431 1276 3435
rect 1408 3431 1412 3435
rect 1552 3431 1556 3435
rect 1704 3431 1708 3435
rect 2104 3431 2108 3435
rect 2192 3431 2196 3435
rect 2296 3431 2300 3435
rect 2408 3431 2412 3435
rect 2536 3431 2540 3435
rect 2672 3431 2676 3435
rect 2808 3431 2812 3435
rect 2816 3431 2820 3435
rect 2952 3431 2956 3435
rect 3104 3431 3108 3435
rect 3256 3431 3260 3435
rect 3336 3431 3340 3435
rect 3416 3431 3420 3435
rect 800 3367 804 3371
rect 3336 3395 3340 3399
rect 2312 3367 2316 3371
rect 552 3331 556 3335
rect 936 3331 940 3335
rect 1384 3331 1388 3335
rect 208 3291 212 3295
rect 336 3291 340 3295
rect 472 3291 476 3295
rect 552 3291 556 3295
rect 624 3291 628 3295
rect 784 3291 788 3295
rect 944 3291 948 3295
rect 1104 3291 1108 3295
rect 1264 3291 1268 3295
rect 1528 3331 1532 3335
rect 2824 3327 2828 3331
rect 1424 3291 1428 3295
rect 1528 3291 1532 3295
rect 1584 3291 1588 3295
rect 1744 3291 1748 3295
rect 2128 3287 2132 3291
rect 2224 3287 2228 3291
rect 2336 3287 2340 3291
rect 2456 3287 2460 3291
rect 2584 3287 2588 3291
rect 2720 3287 2724 3291
rect 344 3275 348 3279
rect 448 3275 452 3279
rect 568 3275 572 3279
rect 656 3275 660 3279
rect 696 3275 700 3279
rect 832 3275 836 3279
rect 976 3275 980 3279
rect 1112 3275 1116 3279
rect 1248 3275 1252 3279
rect 1376 3275 1380 3279
rect 1384 3275 1388 3279
rect 1480 3275 1484 3279
rect 1504 3275 1508 3279
rect 1632 3275 1636 3279
rect 1744 3275 1748 3279
rect 656 3239 660 3243
rect 3080 3327 3084 3331
rect 2864 3287 2868 3291
rect 3008 3287 3012 3291
rect 3080 3287 3084 3291
rect 3160 3287 3164 3291
rect 3312 3287 3316 3291
rect 3472 3287 3476 3291
rect 2128 3263 2132 3267
rect 2272 3263 2276 3267
rect 2408 3263 2412 3267
rect 2544 3263 2548 3267
rect 2680 3263 2684 3267
rect 2816 3263 2820 3267
rect 2824 3263 2828 3267
rect 2952 3263 2956 3267
rect 3088 3263 3092 3267
rect 3224 3263 3228 3267
rect 3368 3263 3372 3267
rect 3504 3263 3508 3267
rect 1480 3239 1484 3243
rect 848 3211 852 3215
rect 1760 3211 1764 3215
rect 2560 3199 2564 3203
rect 488 3135 492 3139
rect 576 3135 580 3139
rect 664 3135 668 3139
rect 768 3135 772 3139
rect 888 3135 892 3139
rect 1024 3135 1028 3139
rect 1192 3135 1196 3139
rect 1376 3135 1380 3139
rect 1568 3135 1572 3139
rect 1744 3135 1748 3139
rect 584 3119 588 3123
rect 664 3119 668 3123
rect 752 3119 756 3123
rect 840 3119 844 3123
rect 928 3119 932 3123
rect 1016 3119 1020 3123
rect 1104 3119 1108 3123
rect 1192 3119 1196 3123
rect 1280 3119 1284 3123
rect 1368 3119 1372 3123
rect 1896 3119 1900 3123
rect 1992 3119 1996 3123
rect 2120 3119 2124 3123
rect 2248 3119 2252 3123
rect 2384 3119 2388 3123
rect 2512 3119 2516 3123
rect 2640 3119 2644 3123
rect 2768 3119 2772 3123
rect 2896 3119 2900 3123
rect 3032 3119 3036 3123
rect 3176 3119 3180 3123
rect 3328 3119 3332 3123
rect 3488 3119 3492 3123
rect 1896 3091 1900 3095
rect 2008 3091 2012 3095
rect 2184 3091 2188 3095
rect 2400 3091 2404 3095
rect 2648 3091 2652 3095
rect 2928 3091 2932 3095
rect 3224 3091 3228 3095
rect 3504 3091 3508 3095
rect 3520 3027 3524 3031
rect 3000 2983 3004 2987
rect 544 2975 548 2979
rect 624 2975 628 2979
rect 712 2975 716 2979
rect 808 2975 812 2979
rect 904 2975 908 2979
rect 1000 2975 1004 2979
rect 1088 2975 1092 2979
rect 1184 2975 1188 2979
rect 1280 2975 1284 2979
rect 1376 2975 1380 2979
rect 1472 2975 1476 2979
rect 464 2963 468 2967
rect 568 2963 572 2967
rect 680 2963 684 2967
rect 800 2963 804 2967
rect 936 2963 940 2967
rect 1080 2963 1084 2967
rect 1240 2963 1244 2967
rect 1408 2963 1412 2967
rect 1584 2963 1588 2967
rect 1744 2963 1748 2967
rect 1896 2943 1900 2947
rect 2048 2943 2052 2947
rect 2224 2943 2228 2947
rect 2392 2943 2396 2947
rect 2544 2943 2548 2947
rect 2688 2943 2692 2947
rect 2816 2943 2820 2947
rect 2928 2943 2932 2947
rect 3000 2943 3004 2947
rect 3040 2943 3044 2947
rect 3144 2943 3148 2947
rect 3240 2943 3244 2947
rect 3336 2943 3340 2947
rect 3424 2943 3428 2947
rect 3504 2943 3508 2947
rect 1896 2931 1900 2935
rect 2080 2931 2084 2935
rect 2288 2931 2292 2935
rect 2480 2931 2484 2935
rect 2664 2931 2668 2935
rect 2832 2931 2836 2935
rect 2992 2931 2996 2935
rect 3144 2931 3148 2935
rect 3296 2931 3300 2935
rect 3448 2931 3452 2935
rect 1760 2899 1764 2903
rect 672 2863 676 2867
rect 312 2823 316 2827
rect 432 2823 436 2827
rect 552 2823 556 2827
rect 672 2823 676 2827
rect 680 2823 684 2827
rect 816 2823 820 2827
rect 952 2823 956 2827
rect 1088 2823 1092 2827
rect 1224 2823 1228 2827
rect 1360 2823 1364 2827
rect 1496 2823 1500 2827
rect 1632 2823 1636 2827
rect 1744 2823 1748 2827
rect 2352 2823 2356 2827
rect 160 2811 164 2815
rect 296 2811 300 2815
rect 440 2811 444 2815
rect 600 2811 604 2815
rect 776 2811 780 2815
rect 952 2811 956 2815
rect 1136 2811 1140 2815
rect 1328 2811 1332 2815
rect 1528 2811 1532 2815
rect 1728 2811 1732 2815
rect 2464 2823 2468 2827
rect 2136 2783 2140 2787
rect 2264 2783 2268 2787
rect 2352 2783 2356 2787
rect 2392 2783 2396 2787
rect 2464 2783 2468 2787
rect 2520 2783 2524 2787
rect 2648 2783 2652 2787
rect 2768 2783 2772 2787
rect 2888 2783 2892 2787
rect 3008 2783 3012 2787
rect 3136 2783 3140 2787
rect 2216 2763 2220 2767
rect 2224 2763 2228 2767
rect 2304 2763 2308 2767
rect 2384 2763 2388 2767
rect 2464 2763 2468 2767
rect 2544 2763 2548 2767
rect 2632 2763 2636 2767
rect 2720 2763 2724 2767
rect 2808 2763 2812 2767
rect 2896 2763 2900 2767
rect 2984 2763 2988 2767
rect 792 2747 796 2751
rect 1744 2747 1748 2751
rect 704 2707 708 2711
rect 136 2667 140 2671
rect 248 2667 252 2671
rect 392 2667 396 2671
rect 552 2667 556 2671
rect 704 2667 708 2671
rect 712 2667 716 2671
rect 880 2667 884 2671
rect 1040 2667 1044 2671
rect 1200 2667 1204 2671
rect 1360 2667 1364 2671
rect 1520 2667 1524 2671
rect 1688 2667 1692 2671
rect 2216 2663 2220 2667
rect 2312 2663 2316 2667
rect 136 2655 140 2659
rect 248 2655 252 2659
rect 392 2655 396 2659
rect 544 2655 548 2659
rect 704 2655 708 2659
rect 872 2655 876 2659
rect 1040 2655 1044 2659
rect 1208 2655 1212 2659
rect 1384 2655 1388 2659
rect 1560 2655 1564 2659
rect 2240 2623 2244 2627
rect 2312 2623 2316 2627
rect 2320 2623 2324 2627
rect 2400 2623 2404 2627
rect 2480 2623 2484 2627
rect 2560 2623 2564 2627
rect 2640 2623 2644 2627
rect 2720 2623 2724 2627
rect 2800 2623 2804 2627
rect 2880 2623 2884 2627
rect 2960 2623 2964 2627
rect 2184 2603 2188 2607
rect 2264 2603 2268 2607
rect 2344 2603 2348 2607
rect 2424 2603 2428 2607
rect 2504 2603 2508 2607
rect 2584 2603 2588 2607
rect 2664 2603 2668 2607
rect 2744 2603 2748 2607
rect 2824 2603 2828 2607
rect 2904 2603 2908 2607
rect 2984 2603 2988 2607
rect 720 2591 724 2595
rect 1576 2591 1580 2595
rect 3000 2539 3004 2543
rect 160 2511 164 2515
rect 280 2511 284 2515
rect 416 2511 420 2515
rect 560 2511 564 2515
rect 704 2511 708 2515
rect 848 2511 852 2515
rect 984 2511 988 2515
rect 1120 2511 1124 2515
rect 1256 2511 1260 2515
rect 1392 2511 1396 2515
rect 1528 2511 1532 2515
rect 328 2495 332 2499
rect 408 2495 412 2499
rect 496 2495 500 2499
rect 592 2495 596 2499
rect 696 2495 700 2499
rect 808 2495 812 2499
rect 928 2495 932 2499
rect 1056 2495 1060 2499
rect 1128 2495 1132 2499
rect 1184 2495 1188 2499
rect 1320 2495 1324 2499
rect 1464 2495 1468 2499
rect 1128 2459 1132 2463
rect 2120 2455 2124 2459
rect 2208 2455 2212 2459
rect 2304 2455 2308 2459
rect 2400 2455 2404 2459
rect 2496 2455 2500 2459
rect 2592 2455 2596 2459
rect 2688 2455 2692 2459
rect 2784 2455 2788 2459
rect 2880 2455 2884 2459
rect 2976 2455 2980 2459
rect 3080 2455 3084 2459
rect 1896 2439 1900 2443
rect 1984 2439 1988 2443
rect 2104 2439 2108 2443
rect 2240 2439 2244 2443
rect 2384 2439 2388 2443
rect 2528 2439 2532 2443
rect 2664 2439 2668 2443
rect 2800 2439 2804 2443
rect 2936 2439 2940 2443
rect 3072 2439 3076 2443
rect 3208 2439 3212 2443
rect 824 2431 828 2435
rect 3224 2375 3228 2379
rect 384 2347 388 2351
rect 464 2347 468 2351
rect 544 2347 548 2351
rect 624 2347 628 2351
rect 704 2347 708 2351
rect 784 2347 788 2351
rect 864 2347 868 2351
rect 944 2347 948 2351
rect 1024 2347 1028 2351
rect 1104 2347 1108 2351
rect 1184 2347 1188 2351
rect 1264 2347 1268 2351
rect 1352 2347 1356 2351
rect 1440 2347 1444 2351
rect 1528 2347 1532 2351
rect 1400 2335 1404 2339
rect 1480 2335 1484 2339
rect 1560 2335 1564 2339
rect 1640 2335 1644 2339
rect 3496 2331 3500 2335
rect 1896 2291 1900 2295
rect 2016 2291 2020 2295
rect 2176 2291 2180 2295
rect 2344 2291 2348 2295
rect 2512 2291 2516 2295
rect 2672 2291 2676 2295
rect 2824 2291 2828 2295
rect 2960 2291 2964 2295
rect 3080 2291 3084 2295
rect 3192 2291 3196 2295
rect 3304 2291 3308 2295
rect 3416 2291 3420 2295
rect 3088 2287 3092 2291
rect 1896 2279 1900 2283
rect 2024 2279 2028 2283
rect 2104 2279 2108 2283
rect 2176 2279 2180 2283
rect 2248 2279 2252 2283
rect 2360 2279 2364 2283
rect 2568 2279 2572 2283
rect 2784 2279 2788 2283
rect 3016 2279 3020 2283
rect 1656 2271 1660 2275
rect 2104 2243 2108 2247
rect 3504 2291 3508 2295
rect 3248 2279 3252 2283
rect 3488 2279 3492 2283
rect 3496 2279 3500 2283
rect 3088 2271 3092 2275
rect 2248 2243 2252 2247
rect 2800 2215 2804 2219
rect 136 2187 140 2191
rect 144 2187 148 2191
rect 216 2187 220 2191
rect 296 2187 300 2191
rect 384 2187 388 2191
rect 520 2187 524 2191
rect 672 2187 676 2191
rect 832 2187 836 2191
rect 1000 2187 1004 2191
rect 1160 2187 1164 2191
rect 1312 2187 1316 2191
rect 1456 2187 1460 2191
rect 1608 2187 1612 2191
rect 1744 2187 1748 2191
rect 184 2171 188 2175
rect 304 2171 308 2175
rect 456 2171 460 2175
rect 632 2171 636 2175
rect 816 2171 820 2175
rect 1008 2171 1012 2175
rect 1192 2171 1196 2175
rect 1384 2171 1388 2175
rect 1576 2171 1580 2175
rect 1744 2171 1748 2175
rect 144 2135 148 2139
rect 2848 2159 2852 2163
rect 2200 2119 2204 2123
rect 2296 2119 2300 2123
rect 2400 2119 2404 2123
rect 2520 2119 2524 2123
rect 2640 2119 2644 2123
rect 2760 2119 2764 2123
rect 1760 2107 1764 2111
rect 2880 2119 2884 2123
rect 2992 2119 2996 2123
rect 3096 2119 3100 2123
rect 3200 2119 3204 2123
rect 3304 2119 3308 2123
rect 3408 2119 3412 2123
rect 3504 2119 3508 2123
rect 2168 2095 2172 2099
rect 2264 2095 2268 2099
rect 2368 2095 2372 2099
rect 2480 2095 2484 2099
rect 2600 2095 2604 2099
rect 2720 2095 2724 2099
rect 2840 2095 2844 2099
rect 2848 2095 2852 2099
rect 2960 2095 2964 2099
rect 3072 2095 3076 2099
rect 3184 2095 3188 2099
rect 3296 2095 3300 2099
rect 3408 2095 3412 2099
rect 3504 2095 3508 2099
rect 496 2067 500 2071
rect 216 2027 220 2031
rect 360 2027 364 2031
rect 1096 2059 1100 2063
rect 520 2027 524 2031
rect 704 2027 708 2031
rect 896 2027 900 2031
rect 3088 2031 3092 2035
rect 3520 2031 3524 2035
rect 1104 2027 1108 2031
rect 1312 2027 1316 2031
rect 1528 2027 1532 2031
rect 1744 2027 1748 2031
rect 136 2015 140 2019
rect 256 2015 260 2019
rect 376 2015 380 2019
rect 488 2015 492 2019
rect 496 2015 500 2019
rect 600 2015 604 2019
rect 712 2015 716 2019
rect 816 2015 820 2019
rect 920 2015 924 2019
rect 1016 2015 1020 2019
rect 1096 2015 1100 2019
rect 1104 2015 1108 2019
rect 1200 2015 1204 2019
rect 1288 2015 1292 2019
rect 1384 2015 1388 2019
rect 1480 2015 1484 2019
rect 1576 2015 1580 2019
rect 1664 2015 1668 2019
rect 1744 2015 1748 2019
rect 1496 1951 1500 1955
rect 1760 1951 1764 1955
rect 2072 1951 2076 1955
rect 2208 1951 2212 1955
rect 2360 1951 2364 1955
rect 2520 1951 2524 1955
rect 2680 1951 2684 1955
rect 2848 1951 2852 1955
rect 3016 1951 3020 1955
rect 3184 1951 3188 1955
rect 3352 1951 3356 1955
rect 3504 1951 3508 1955
rect 1896 1939 1900 1943
rect 2000 1939 2004 1943
rect 2128 1939 2132 1943
rect 2248 1939 2252 1943
rect 2368 1939 2372 1943
rect 2480 1939 2484 1943
rect 2592 1939 2596 1943
rect 2712 1939 2716 1943
rect 2832 1939 2836 1943
rect 1912 1875 1916 1879
rect 2848 1875 2852 1879
rect 168 1867 172 1871
rect 328 1867 332 1871
rect 488 1867 492 1871
rect 648 1867 652 1871
rect 800 1867 804 1871
rect 944 1867 948 1871
rect 1080 1867 1084 1871
rect 1216 1867 1220 1871
rect 1352 1867 1356 1871
rect 1488 1867 1492 1871
rect 1624 1867 1628 1871
rect 1744 1867 1748 1871
rect 152 1855 156 1859
rect 296 1855 300 1859
rect 440 1855 444 1859
rect 592 1855 596 1859
rect 680 1855 684 1859
rect 744 1855 748 1859
rect 896 1855 900 1859
rect 1048 1855 1052 1859
rect 1128 1855 1132 1859
rect 1200 1855 1204 1859
rect 1344 1855 1348 1859
rect 1480 1855 1484 1859
rect 1624 1855 1628 1859
rect 1744 1855 1748 1859
rect 680 1819 684 1823
rect 1128 1819 1132 1823
rect 2112 1819 2116 1823
rect 1896 1799 1900 1803
rect 1992 1799 1996 1803
rect 2112 1799 2116 1803
rect 2120 1799 2124 1803
rect 2248 1799 2252 1803
rect 2384 1799 2388 1803
rect 2520 1799 2524 1803
rect 2656 1799 2660 1803
rect 2808 1799 2812 1803
rect 2976 1799 2980 1803
rect 3152 1799 3156 1803
rect 3336 1799 3340 1803
rect 3504 1799 3508 1803
rect 912 1791 916 1795
rect 1896 1775 1900 1779
rect 2024 1775 2028 1779
rect 2184 1775 2188 1779
rect 2352 1775 2356 1779
rect 2520 1775 2524 1779
rect 2680 1775 2684 1779
rect 2832 1775 2836 1779
rect 2976 1775 2980 1779
rect 3112 1775 3116 1779
rect 3248 1775 3252 1779
rect 3384 1775 3388 1779
rect 3504 1775 3508 1779
rect 248 1711 252 1715
rect 424 1711 428 1715
rect 592 1711 596 1715
rect 752 1711 756 1715
rect 896 1711 900 1715
rect 1024 1711 1028 1715
rect 1144 1711 1148 1715
rect 1264 1711 1268 1715
rect 1392 1711 1396 1715
rect 2536 1711 2540 1715
rect 3400 1711 3404 1715
rect 3520 1711 3524 1715
rect 184 1695 188 1699
rect 304 1695 308 1699
rect 440 1695 444 1699
rect 584 1695 588 1699
rect 736 1695 740 1699
rect 888 1695 892 1699
rect 1032 1695 1036 1699
rect 1176 1695 1180 1699
rect 1312 1695 1316 1699
rect 1440 1695 1444 1699
rect 1520 1695 1524 1699
rect 1568 1695 1572 1699
rect 1704 1695 1708 1699
rect 1520 1659 1524 1663
rect 3488 1671 3492 1675
rect 1048 1631 1052 1635
rect 1896 1631 1900 1635
rect 1992 1631 1996 1635
rect 2136 1631 2140 1635
rect 2296 1631 2300 1635
rect 2472 1631 2476 1635
rect 2648 1631 2652 1635
rect 2816 1631 2820 1635
rect 2968 1631 2972 1635
rect 3112 1631 3116 1635
rect 3248 1631 3252 1635
rect 3384 1631 3388 1635
rect 1968 1615 1972 1619
rect 2088 1615 2092 1619
rect 2224 1615 2228 1619
rect 2360 1615 2364 1619
rect 2496 1615 2500 1619
rect 2632 1615 2636 1619
rect 2768 1615 2772 1619
rect 2904 1615 2908 1619
rect 3048 1615 3052 1619
rect 3200 1615 3204 1619
rect 3360 1615 3364 1619
rect 2512 1551 2516 1555
rect 168 1547 172 1551
rect 352 1547 356 1551
rect 544 1547 548 1551
rect 728 1547 732 1551
rect 904 1547 908 1551
rect 1072 1547 1076 1551
rect 1224 1547 1228 1551
rect 1360 1547 1364 1551
rect 1496 1547 1500 1551
rect 1624 1547 1628 1551
rect 1744 1547 1748 1551
rect 128 1531 132 1535
rect 136 1531 140 1535
rect 240 1531 244 1535
rect 376 1531 380 1535
rect 520 1531 524 1535
rect 664 1531 668 1535
rect 808 1531 812 1535
rect 944 1531 948 1535
rect 1072 1531 1076 1535
rect 1200 1531 1204 1535
rect 1328 1531 1332 1535
rect 1464 1531 1468 1535
rect 3480 1511 3484 1515
rect 2088 1471 2092 1475
rect 2168 1471 2172 1475
rect 2256 1471 2260 1475
rect 2344 1471 2348 1475
rect 2440 1471 2444 1475
rect 2536 1471 2540 1475
rect 2648 1471 2652 1475
rect 2784 1471 2788 1475
rect 2944 1471 2948 1475
rect 3120 1471 3124 1475
rect 3304 1471 3308 1475
rect 824 1467 828 1471
rect 3504 1631 3508 1635
rect 3504 1615 3508 1619
rect 3488 1471 3492 1475
rect 3496 1471 3500 1475
rect 2256 1455 2260 1459
rect 2336 1455 2340 1459
rect 2416 1455 2420 1459
rect 2496 1455 2500 1459
rect 2600 1455 2604 1459
rect 2728 1455 2732 1459
rect 2888 1455 2892 1459
rect 3072 1455 3076 1459
rect 3272 1455 3276 1459
rect 3472 1455 3476 1459
rect 3480 1455 3484 1459
rect 128 1427 132 1431
rect 2416 1391 2420 1395
rect 2512 1391 2516 1395
rect 2616 1391 2620 1395
rect 3488 1391 3492 1395
rect 136 1387 140 1391
rect 232 1387 236 1391
rect 360 1387 364 1391
rect 480 1387 484 1391
rect 600 1387 604 1391
rect 720 1387 724 1391
rect 832 1387 836 1391
rect 936 1387 940 1391
rect 1040 1387 1044 1391
rect 1144 1387 1148 1391
rect 1256 1387 1260 1391
rect 128 1359 132 1363
rect 136 1359 140 1363
rect 280 1359 284 1363
rect 424 1359 428 1363
rect 576 1359 580 1363
rect 728 1359 732 1363
rect 872 1359 876 1363
rect 1016 1359 1020 1363
rect 1160 1359 1164 1363
rect 1312 1359 1316 1363
rect 1384 1359 1388 1363
rect 1464 1359 1468 1363
rect 1600 1359 1604 1363
rect 1616 1359 1620 1363
rect 1384 1323 1388 1327
rect 440 1295 444 1299
rect 2264 1315 2268 1319
rect 2344 1315 2348 1319
rect 2416 1315 2420 1319
rect 2424 1315 2428 1319
rect 2504 1315 2508 1319
rect 2592 1315 2596 1319
rect 2696 1315 2700 1319
rect 2808 1315 2812 1319
rect 2920 1315 2924 1319
rect 3040 1315 3044 1319
rect 3160 1315 3164 1319
rect 3280 1315 3284 1319
rect 3400 1315 3404 1319
rect 3504 1315 3508 1319
rect 2208 1291 2212 1295
rect 2288 1291 2292 1295
rect 2368 1291 2372 1295
rect 2448 1291 2452 1295
rect 2520 1291 2524 1295
rect 2544 1291 2548 1295
rect 2656 1291 2660 1295
rect 2784 1291 2788 1295
rect 2920 1291 2924 1295
rect 3064 1291 3068 1295
rect 3208 1291 3212 1295
rect 3360 1291 3364 1295
rect 3488 1291 3492 1295
rect 3504 1291 3508 1295
rect 128 1255 132 1259
rect 208 1255 212 1259
rect 1600 1255 1604 1259
rect 2520 1255 2524 1259
rect 2224 1227 2228 1231
rect 2800 1227 2804 1231
rect 3376 1227 3380 1231
rect 208 1223 212 1227
rect 136 1215 140 1219
rect 264 1215 268 1219
rect 424 1215 428 1219
rect 592 1215 596 1219
rect 760 1215 764 1219
rect 928 1215 932 1219
rect 1080 1215 1084 1219
rect 1224 1215 1228 1219
rect 1352 1215 1356 1219
rect 1480 1215 1484 1219
rect 1608 1215 1612 1219
rect 1736 1215 1740 1219
rect 128 1195 132 1199
rect 136 1195 140 1199
rect 304 1195 308 1199
rect 480 1195 484 1199
rect 664 1195 668 1199
rect 840 1195 844 1199
rect 1000 1195 1004 1199
rect 1152 1195 1156 1199
rect 1288 1195 1292 1199
rect 1408 1195 1412 1199
rect 1528 1195 1532 1199
rect 1648 1195 1652 1199
rect 1744 1195 1748 1199
rect 3488 1187 3492 1191
rect 2112 1147 2116 1151
rect 2208 1147 2212 1151
rect 2304 1147 2308 1151
rect 2408 1147 2412 1151
rect 2528 1147 2532 1151
rect 2648 1147 2652 1151
rect 2776 1147 2780 1151
rect 2912 1147 2916 1151
rect 3056 1147 3060 1151
rect 3200 1147 3204 1151
rect 3344 1147 3348 1151
rect 3496 1147 3500 1151
rect 320 1131 324 1135
rect 128 1095 132 1099
rect 1888 1127 1892 1131
rect 1896 1127 1900 1131
rect 2120 1127 2124 1131
rect 2264 1127 2268 1131
rect 2352 1127 2356 1131
rect 2568 1127 2572 1131
rect 2768 1127 2772 1131
rect 2960 1127 2964 1131
rect 3152 1127 3156 1131
rect 3336 1127 3340 1131
rect 3496 1127 3500 1131
rect 3504 1127 3508 1131
rect 360 1087 364 1091
rect 136 1055 140 1059
rect 248 1055 252 1059
rect 768 1087 772 1091
rect 384 1055 388 1059
rect 520 1055 524 1059
rect 648 1055 652 1059
rect 776 1055 780 1059
rect 896 1055 900 1059
rect 1016 1055 1020 1059
rect 1136 1055 1140 1059
rect 1256 1055 1260 1059
rect 1376 1055 1380 1059
rect 1504 1055 1508 1059
rect 1632 1055 1636 1059
rect 1744 1055 1748 1059
rect 128 1031 132 1035
rect 136 1031 140 1035
rect 232 1031 236 1035
rect 352 1031 356 1035
rect 360 1031 364 1035
rect 464 1031 468 1035
rect 568 1031 572 1035
rect 664 1031 668 1035
rect 760 1031 764 1035
rect 768 1031 772 1035
rect 848 1031 852 1035
rect 936 1031 940 1035
rect 1024 1031 1028 1035
rect 1120 1031 1124 1035
rect 1216 1031 1220 1035
rect 2264 1091 2268 1095
rect 1912 1063 1916 1067
rect 1888 1027 1892 1031
rect 2480 1027 2484 1031
rect 1896 987 1900 991
rect 2016 987 2020 991
rect 2168 987 2172 991
rect 2328 987 2332 991
rect 2632 1027 2636 1031
rect 2488 987 2492 991
rect 3344 1027 3348 1031
rect 3496 1027 3500 1031
rect 2640 987 2644 991
rect 2792 987 2796 991
rect 2936 987 2940 991
rect 3080 987 3084 991
rect 3224 987 3228 991
rect 3376 987 3380 991
rect 3504 987 3508 991
rect 1888 971 1892 975
rect 1896 971 1900 975
rect 1976 971 1980 975
rect 2072 971 2076 975
rect 2192 971 2196 975
rect 2328 971 2332 975
rect 2472 971 2476 975
rect 2480 971 2484 975
rect 2624 971 2628 975
rect 2632 971 2636 975
rect 2784 971 2788 975
rect 2960 971 2964 975
rect 3144 971 3148 975
rect 3336 971 3340 975
rect 3344 971 3348 975
rect 3496 971 3500 975
rect 3504 971 3508 975
rect 248 967 252 971
rect 256 967 260 971
rect 128 919 132 923
rect 1216 967 1220 971
rect 1232 967 1236 971
rect 960 919 964 923
rect 136 879 140 883
rect 256 879 260 883
rect 264 879 268 883
rect 416 879 420 883
rect 560 879 564 883
rect 704 879 708 883
rect 840 879 844 883
rect 976 879 980 883
rect 1104 879 1108 883
rect 1216 879 1220 883
rect 1224 879 1228 883
rect 1336 879 1340 883
rect 1440 879 1444 883
rect 1544 879 1548 883
rect 1656 879 1660 883
rect 1744 879 1748 883
rect 136 863 140 867
rect 240 863 244 867
rect 376 863 380 867
rect 512 863 516 867
rect 656 863 660 867
rect 752 863 756 867
rect 808 863 812 867
rect 952 863 956 867
rect 960 863 964 867
rect 1096 863 1100 867
rect 1240 863 1244 867
rect 1376 863 1380 867
rect 1504 863 1508 867
rect 1632 863 1636 867
rect 1744 863 1748 867
rect 752 827 756 831
rect 2344 907 2348 911
rect 2976 907 2980 911
rect 1888 827 1892 831
rect 1904 859 1908 863
rect 2168 859 2172 863
rect 2552 859 2556 863
rect 1920 819 1924 823
rect 2096 819 2100 823
rect 2168 819 2172 823
rect 2272 819 2276 823
rect 2456 819 2460 823
rect 2560 859 2564 863
rect 3496 859 3500 863
rect 2560 819 2564 823
rect 2656 819 2660 823
rect 2864 819 2868 823
rect 3080 819 3084 823
rect 3304 819 3308 823
rect 3504 819 3508 823
rect 1896 807 1900 811
rect 1904 807 1908 811
rect 2008 807 2012 811
rect 2160 807 2164 811
rect 2320 807 2324 811
rect 2480 807 2484 811
rect 2552 807 2556 811
rect 2640 807 2644 811
rect 2800 807 2804 811
rect 2952 807 2956 811
rect 3096 807 3100 811
rect 3240 807 3244 811
rect 3384 807 3388 811
rect 3496 807 3500 811
rect 3504 807 3508 811
rect 1256 799 1260 803
rect 2496 743 2500 747
rect 3400 743 3404 747
rect 136 711 140 715
rect 216 711 220 715
rect 304 711 308 715
rect 416 711 420 715
rect 544 711 548 715
rect 688 711 692 715
rect 840 711 844 715
rect 992 711 996 715
rect 1144 711 1148 715
rect 1296 711 1300 715
rect 1448 711 1452 715
rect 1608 711 1612 715
rect 2592 707 2596 711
rect 3496 707 3500 711
rect 224 691 228 695
rect 312 691 316 695
rect 416 691 420 695
rect 536 691 540 695
rect 672 691 676 695
rect 808 691 812 695
rect 944 691 948 695
rect 1080 691 1084 695
rect 1208 691 1212 695
rect 1328 691 1332 695
rect 1448 691 1452 695
rect 1576 691 1580 695
rect 2736 699 2740 703
rect 1968 667 1972 671
rect 2064 667 2068 671
rect 2176 667 2180 671
rect 2304 667 2308 671
rect 2448 667 2452 671
rect 2592 667 2596 671
rect 2600 667 2604 671
rect 2752 667 2756 671
rect 2904 667 2908 671
rect 3056 667 3060 671
rect 3208 667 3212 671
rect 3360 667 3364 671
rect 3504 667 3508 671
rect 2168 655 2172 659
rect 2264 655 2268 659
rect 2368 655 2372 659
rect 2480 655 2484 659
rect 2600 655 2604 659
rect 2728 655 2732 659
rect 2736 655 2740 659
rect 2856 655 2860 659
rect 2984 655 2988 659
rect 3112 655 3116 659
rect 3184 655 3188 659
rect 3240 655 3244 659
rect 3368 655 3372 659
rect 3504 655 3508 659
rect 952 627 956 631
rect 960 627 964 631
rect 2616 591 2620 595
rect 3184 555 3188 559
rect 448 543 452 547
rect 528 543 532 547
rect 608 543 612 547
rect 688 543 692 547
rect 776 543 780 547
rect 872 543 876 547
rect 952 543 956 547
rect 960 543 964 547
rect 1048 543 1052 547
rect 1144 543 1148 547
rect 1240 543 1244 547
rect 1336 543 1340 547
rect 1432 543 1436 547
rect 328 519 332 523
rect 416 519 420 523
rect 504 519 508 523
rect 584 519 588 523
rect 664 519 668 523
rect 744 519 748 523
rect 832 519 836 523
rect 920 519 924 523
rect 1008 519 1012 523
rect 1096 519 1100 523
rect 1184 519 1188 523
rect 1272 519 1276 523
rect 2264 515 2268 519
rect 2344 515 2348 519
rect 2424 515 2428 519
rect 2504 515 2508 519
rect 2592 515 2596 519
rect 2696 515 2700 519
rect 2816 515 2820 519
rect 2960 515 2964 519
rect 3112 515 3116 519
rect 3280 515 3284 519
rect 3448 515 3452 519
rect 2184 495 2188 499
rect 2280 495 2284 499
rect 2352 495 2356 499
rect 2376 495 2380 499
rect 2480 495 2484 499
rect 2576 495 2580 499
rect 2680 495 2684 499
rect 2784 495 2788 499
rect 2904 495 2908 499
rect 3032 495 3036 499
rect 3168 495 3172 499
rect 3312 495 3316 499
rect 3464 495 3468 499
rect 2352 459 2356 463
rect 752 455 756 459
rect 760 455 764 459
rect 536 411 540 415
rect 224 371 228 375
rect 336 371 340 375
rect 448 371 452 375
rect 648 411 652 415
rect 2200 431 2204 435
rect 2592 431 2596 435
rect 3480 431 3484 435
rect 3488 431 3492 435
rect 2328 391 2332 395
rect 2232 383 2236 387
rect 560 371 564 375
rect 648 371 652 375
rect 664 371 668 375
rect 752 371 756 375
rect 760 371 764 375
rect 848 371 852 375
rect 936 371 940 375
rect 1024 371 1028 375
rect 1112 371 1116 375
rect 1200 371 1204 375
rect 1296 371 1300 375
rect 1976 351 1980 355
rect 2064 351 2068 355
rect 2160 351 2164 355
rect 128 347 132 351
rect 136 347 140 351
rect 256 347 260 351
rect 392 347 396 351
rect 528 347 532 351
rect 536 347 540 351
rect 664 347 668 351
rect 784 347 788 351
rect 904 347 908 351
rect 1016 347 1020 351
rect 1120 347 1124 351
rect 1224 347 1228 351
rect 1328 347 1332 351
rect 1432 347 1436 351
rect 2256 351 2260 355
rect 2328 351 2332 355
rect 2360 351 2364 355
rect 2472 351 2476 355
rect 2608 351 2612 355
rect 2760 351 2764 355
rect 2928 351 2932 355
rect 3112 351 3116 355
rect 3304 351 3308 355
rect 3488 351 3492 355
rect 3496 351 3500 355
rect 2208 335 2212 339
rect 2232 335 2236 339
rect 2288 335 2292 339
rect 2376 335 2380 339
rect 2472 335 2476 339
rect 2584 335 2588 339
rect 2712 335 2716 339
rect 2840 335 2844 339
rect 2976 335 2980 339
rect 3112 335 3116 339
rect 3248 335 3252 339
rect 3384 335 3388 339
rect 3504 335 3508 339
rect 2728 271 2732 275
rect 3520 271 3524 275
rect 128 239 132 243
rect 648 239 652 243
rect 2624 231 2628 235
rect 136 199 140 203
rect 248 199 252 203
rect 392 199 396 203
rect 544 199 548 203
rect 648 199 652 203
rect 696 199 700 203
rect 848 199 852 203
rect 992 199 996 203
rect 1120 199 1124 203
rect 1240 199 1244 203
rect 1360 199 1364 203
rect 1480 199 1484 203
rect 1600 199 1604 203
rect 1992 191 1996 195
rect 2120 191 2124 195
rect 2256 191 2260 195
rect 2392 191 2396 195
rect 2536 191 2540 195
rect 2680 191 2684 195
rect 2816 191 2820 195
rect 2952 191 2956 195
rect 3096 191 3100 195
rect 3240 191 3244 195
rect 3384 191 3388 195
rect 3504 191 3508 195
rect 1896 167 1900 171
rect 1976 167 1980 171
rect 2080 167 2084 171
rect 2208 167 2212 171
rect 2344 167 2348 171
rect 2480 167 2484 171
rect 2616 167 2620 171
rect 2624 167 2628 171
rect 2736 167 2740 171
rect 2848 167 2852 171
rect 2952 167 2956 171
rect 3056 167 3060 171
rect 3152 167 3156 171
rect 3240 167 3244 171
rect 3336 167 3340 171
rect 3424 167 3428 171
rect 3504 167 3508 171
rect 136 151 140 155
rect 216 151 220 155
rect 296 151 300 155
rect 376 151 380 155
rect 456 151 460 155
rect 536 151 540 155
rect 616 151 620 155
rect 696 151 700 155
rect 776 151 780 155
rect 856 151 860 155
rect 936 151 940 155
rect 1016 151 1020 155
rect 1096 151 1100 155
rect 1176 151 1180 155
rect 1248 151 1252 155
rect 1256 151 1260 155
rect 1336 151 1340 155
rect 1416 151 1420 155
rect 1488 151 1492 155
rect 1504 151 1508 155
rect 1584 151 1588 155
rect 1664 151 1668 155
rect 1744 151 1748 155
rect 1248 115 1252 119
rect 1488 115 1492 119
<< m2 >>
rect 134 3648 140 3649
rect 110 3645 116 3646
rect 110 3641 111 3645
rect 115 3641 116 3645
rect 134 3644 135 3648
rect 139 3644 140 3648
rect 134 3643 140 3644
rect 214 3648 220 3649
rect 214 3644 215 3648
rect 219 3644 220 3648
rect 214 3643 220 3644
rect 294 3648 300 3649
rect 294 3644 295 3648
rect 299 3644 300 3648
rect 294 3643 300 3644
rect 1830 3645 1836 3646
rect 110 3640 116 3641
rect 1830 3641 1831 3645
rect 1835 3641 1836 3645
rect 1830 3640 1836 3641
rect 202 3639 208 3640
rect 136 3636 153 3638
rect 134 3635 140 3636
rect 134 3631 135 3635
rect 139 3631 140 3635
rect 202 3635 203 3639
rect 207 3638 208 3639
rect 282 3639 288 3640
rect 207 3636 233 3638
rect 207 3635 208 3636
rect 202 3634 208 3635
rect 282 3635 283 3639
rect 287 3638 288 3639
rect 287 3636 313 3638
rect 287 3635 288 3636
rect 282 3634 288 3635
rect 134 3630 140 3631
rect 110 3628 116 3629
rect 110 3624 111 3628
rect 115 3624 116 3628
rect 110 3623 116 3624
rect 1830 3628 1836 3629
rect 1830 3624 1831 3628
rect 1835 3624 1836 3628
rect 1830 3623 1836 3624
rect 142 3610 148 3611
rect 142 3606 143 3610
rect 147 3606 148 3610
rect 142 3605 148 3606
rect 222 3610 228 3611
rect 222 3606 223 3610
rect 227 3606 228 3610
rect 222 3605 228 3606
rect 302 3610 308 3611
rect 302 3606 303 3610
rect 307 3606 308 3610
rect 302 3605 308 3606
rect 2826 3603 2832 3604
rect 2826 3602 2827 3603
rect 2748 3600 2827 3602
rect 135 3599 141 3600
rect 135 3595 136 3599
rect 140 3598 141 3599
rect 202 3599 208 3600
rect 202 3598 203 3599
rect 140 3596 203 3598
rect 140 3595 141 3596
rect 135 3594 141 3595
rect 202 3595 203 3596
rect 207 3595 208 3599
rect 202 3594 208 3595
rect 215 3599 221 3600
rect 215 3595 216 3599
rect 220 3598 221 3599
rect 282 3599 288 3600
rect 282 3598 283 3599
rect 220 3596 283 3598
rect 220 3595 221 3596
rect 215 3594 221 3595
rect 282 3595 283 3596
rect 287 3595 288 3599
rect 282 3594 288 3595
rect 2055 3595 2061 3596
rect 2055 3591 2056 3595
rect 2060 3594 2061 3595
rect 2070 3595 2076 3596
rect 2070 3594 2071 3595
rect 2060 3592 2071 3594
rect 2060 3591 2061 3592
rect 2055 3590 2061 3591
rect 2070 3591 2071 3592
rect 2075 3591 2076 3595
rect 2070 3590 2076 3591
rect 2114 3595 2120 3596
rect 2114 3591 2115 3595
rect 2119 3594 2120 3595
rect 2143 3595 2149 3596
rect 2143 3594 2144 3595
rect 2119 3592 2144 3594
rect 2119 3591 2120 3592
rect 2114 3590 2120 3591
rect 2143 3591 2144 3592
rect 2148 3591 2149 3595
rect 2143 3590 2149 3591
rect 2202 3595 2208 3596
rect 2202 3591 2203 3595
rect 2207 3594 2208 3595
rect 2247 3595 2253 3596
rect 2247 3594 2248 3595
rect 2207 3592 2248 3594
rect 2207 3591 2208 3592
rect 2202 3590 2208 3591
rect 2247 3591 2248 3592
rect 2252 3591 2253 3595
rect 2247 3590 2253 3591
rect 2306 3595 2312 3596
rect 2306 3591 2307 3595
rect 2311 3594 2312 3595
rect 2359 3595 2365 3596
rect 2359 3594 2360 3595
rect 2311 3592 2360 3594
rect 2311 3591 2312 3592
rect 2306 3590 2312 3591
rect 2359 3591 2360 3592
rect 2364 3591 2365 3595
rect 2359 3590 2365 3591
rect 2418 3595 2424 3596
rect 2418 3591 2419 3595
rect 2423 3594 2424 3595
rect 2471 3595 2477 3596
rect 2471 3594 2472 3595
rect 2423 3592 2472 3594
rect 2423 3591 2424 3592
rect 2418 3590 2424 3591
rect 2471 3591 2472 3592
rect 2476 3591 2477 3595
rect 2471 3590 2477 3591
rect 2530 3595 2536 3596
rect 2530 3591 2531 3595
rect 2535 3594 2536 3595
rect 2583 3595 2589 3596
rect 2583 3594 2584 3595
rect 2535 3592 2584 3594
rect 2535 3591 2536 3592
rect 2530 3590 2536 3591
rect 2583 3591 2584 3592
rect 2588 3591 2589 3595
rect 2583 3590 2589 3591
rect 2695 3595 2701 3596
rect 2695 3591 2696 3595
rect 2700 3594 2701 3595
rect 2748 3594 2750 3600
rect 2826 3599 2827 3600
rect 2831 3599 2832 3603
rect 2826 3598 2832 3599
rect 2700 3592 2750 3594
rect 2754 3595 2760 3596
rect 2700 3591 2701 3592
rect 2695 3590 2701 3591
rect 2754 3591 2755 3595
rect 2759 3594 2760 3595
rect 2807 3595 2813 3596
rect 2807 3594 2808 3595
rect 2759 3592 2808 3594
rect 2759 3591 2760 3592
rect 2754 3590 2760 3591
rect 2807 3591 2808 3592
rect 2812 3591 2813 3595
rect 2807 3590 2813 3591
rect 2866 3595 2872 3596
rect 2866 3591 2867 3595
rect 2871 3594 2872 3595
rect 2911 3595 2917 3596
rect 2911 3594 2912 3595
rect 2871 3592 2912 3594
rect 2871 3591 2872 3592
rect 2866 3590 2872 3591
rect 2911 3591 2912 3592
rect 2916 3591 2917 3595
rect 2911 3590 2917 3591
rect 2970 3595 2976 3596
rect 2970 3591 2971 3595
rect 2975 3594 2976 3595
rect 3007 3595 3013 3596
rect 3007 3594 3008 3595
rect 2975 3592 3008 3594
rect 2975 3591 2976 3592
rect 2970 3590 2976 3591
rect 3007 3591 3008 3592
rect 3012 3591 3013 3595
rect 3007 3590 3013 3591
rect 3066 3595 3072 3596
rect 3066 3591 3067 3595
rect 3071 3594 3072 3595
rect 3103 3595 3109 3596
rect 3103 3594 3104 3595
rect 3071 3592 3104 3594
rect 3071 3591 3072 3592
rect 3066 3590 3072 3591
rect 3103 3591 3104 3592
rect 3108 3591 3109 3595
rect 3103 3590 3109 3591
rect 3162 3595 3168 3596
rect 3162 3591 3163 3595
rect 3167 3594 3168 3595
rect 3199 3595 3205 3596
rect 3199 3594 3200 3595
rect 3167 3592 3200 3594
rect 3167 3591 3168 3592
rect 3162 3590 3168 3591
rect 3199 3591 3200 3592
rect 3204 3591 3205 3595
rect 3199 3590 3205 3591
rect 3258 3595 3264 3596
rect 3258 3591 3259 3595
rect 3263 3594 3264 3595
rect 3295 3595 3301 3596
rect 3295 3594 3296 3595
rect 3263 3592 3296 3594
rect 3263 3591 3264 3592
rect 3258 3590 3264 3591
rect 3295 3591 3296 3592
rect 3300 3591 3301 3595
rect 3295 3590 3301 3591
rect 3354 3595 3360 3596
rect 3354 3591 3355 3595
rect 3359 3594 3360 3595
rect 3391 3595 3397 3596
rect 3391 3594 3392 3595
rect 3359 3592 3392 3594
rect 3359 3591 3360 3592
rect 3354 3590 3360 3591
rect 3391 3591 3392 3592
rect 3396 3591 3397 3595
rect 3391 3590 3397 3591
rect 134 3587 141 3588
rect 134 3583 135 3587
rect 140 3583 141 3587
rect 134 3582 141 3583
rect 194 3587 200 3588
rect 194 3583 195 3587
rect 199 3586 200 3587
rect 215 3587 221 3588
rect 215 3586 216 3587
rect 199 3584 216 3586
rect 199 3583 200 3584
rect 194 3582 200 3583
rect 215 3583 216 3584
rect 220 3583 221 3587
rect 215 3582 221 3583
rect 274 3587 280 3588
rect 274 3583 275 3587
rect 279 3586 280 3587
rect 335 3587 341 3588
rect 335 3586 336 3587
rect 279 3584 336 3586
rect 279 3583 280 3584
rect 274 3582 280 3583
rect 335 3583 336 3584
rect 340 3583 341 3587
rect 335 3582 341 3583
rect 394 3587 400 3588
rect 394 3583 395 3587
rect 399 3586 400 3587
rect 463 3587 469 3588
rect 463 3586 464 3587
rect 399 3584 464 3586
rect 399 3583 400 3584
rect 394 3582 400 3583
rect 463 3583 464 3584
rect 468 3583 469 3587
rect 463 3582 469 3583
rect 522 3587 528 3588
rect 522 3583 523 3587
rect 527 3586 528 3587
rect 599 3587 605 3588
rect 599 3586 600 3587
rect 527 3584 600 3586
rect 527 3583 528 3584
rect 522 3582 528 3583
rect 599 3583 600 3584
rect 604 3583 605 3587
rect 599 3582 605 3583
rect 658 3587 664 3588
rect 658 3583 659 3587
rect 663 3586 664 3587
rect 735 3587 741 3588
rect 735 3586 736 3587
rect 663 3584 736 3586
rect 663 3583 664 3584
rect 658 3582 664 3583
rect 735 3583 736 3584
rect 740 3583 741 3587
rect 735 3582 741 3583
rect 871 3587 877 3588
rect 871 3583 872 3587
rect 876 3586 877 3587
rect 886 3587 892 3588
rect 886 3586 887 3587
rect 876 3584 887 3586
rect 876 3583 877 3584
rect 871 3582 877 3583
rect 886 3583 887 3584
rect 891 3583 892 3587
rect 886 3582 892 3583
rect 930 3587 936 3588
rect 930 3583 931 3587
rect 935 3586 936 3587
rect 991 3587 997 3588
rect 991 3586 992 3587
rect 935 3584 992 3586
rect 935 3583 936 3584
rect 930 3582 936 3583
rect 991 3583 992 3584
rect 996 3583 997 3587
rect 991 3582 997 3583
rect 1050 3587 1056 3588
rect 1050 3583 1051 3587
rect 1055 3586 1056 3587
rect 1103 3587 1109 3588
rect 1103 3586 1104 3587
rect 1055 3584 1104 3586
rect 1055 3583 1056 3584
rect 1050 3582 1056 3583
rect 1103 3583 1104 3584
rect 1108 3583 1109 3587
rect 1103 3582 1109 3583
rect 1162 3587 1168 3588
rect 1162 3583 1163 3587
rect 1167 3586 1168 3587
rect 1215 3587 1221 3588
rect 1215 3586 1216 3587
rect 1167 3584 1216 3586
rect 1167 3583 1168 3584
rect 1162 3582 1168 3583
rect 1215 3583 1216 3584
rect 1220 3583 1221 3587
rect 1215 3582 1221 3583
rect 1274 3587 1280 3588
rect 1274 3583 1275 3587
rect 1279 3586 1280 3587
rect 1319 3587 1325 3588
rect 1319 3586 1320 3587
rect 1279 3584 1320 3586
rect 1279 3583 1280 3584
rect 1274 3582 1280 3583
rect 1319 3583 1320 3584
rect 1324 3583 1325 3587
rect 1319 3582 1325 3583
rect 1378 3587 1384 3588
rect 1378 3583 1379 3587
rect 1383 3586 1384 3587
rect 1415 3587 1421 3588
rect 1415 3586 1416 3587
rect 1383 3584 1416 3586
rect 1383 3583 1384 3584
rect 1378 3582 1384 3583
rect 1415 3583 1416 3584
rect 1420 3583 1421 3587
rect 1415 3582 1421 3583
rect 1474 3587 1480 3588
rect 1474 3583 1475 3587
rect 1479 3586 1480 3587
rect 1519 3587 1525 3588
rect 1519 3586 1520 3587
rect 1479 3584 1520 3586
rect 1479 3583 1480 3584
rect 1474 3582 1480 3583
rect 1519 3583 1520 3584
rect 1524 3583 1525 3587
rect 1519 3582 1525 3583
rect 1578 3587 1584 3588
rect 1578 3583 1579 3587
rect 1583 3586 1584 3587
rect 1623 3587 1629 3588
rect 1623 3586 1624 3587
rect 1583 3584 1624 3586
rect 1583 3583 1584 3584
rect 1578 3582 1584 3583
rect 1623 3583 1624 3584
rect 1628 3583 1629 3587
rect 1623 3582 1629 3583
rect 2062 3586 2068 3587
rect 2062 3582 2063 3586
rect 2067 3582 2068 3586
rect 2062 3581 2068 3582
rect 2150 3586 2156 3587
rect 2150 3582 2151 3586
rect 2155 3582 2156 3586
rect 2150 3581 2156 3582
rect 2254 3586 2260 3587
rect 2254 3582 2255 3586
rect 2259 3582 2260 3586
rect 2254 3581 2260 3582
rect 2366 3586 2372 3587
rect 2366 3582 2367 3586
rect 2371 3582 2372 3586
rect 2366 3581 2372 3582
rect 2478 3586 2484 3587
rect 2478 3582 2479 3586
rect 2483 3582 2484 3586
rect 2478 3581 2484 3582
rect 2590 3586 2596 3587
rect 2590 3582 2591 3586
rect 2595 3582 2596 3586
rect 2590 3581 2596 3582
rect 2702 3586 2708 3587
rect 2702 3582 2703 3586
rect 2707 3582 2708 3586
rect 2702 3581 2708 3582
rect 2814 3586 2820 3587
rect 2814 3582 2815 3586
rect 2819 3582 2820 3586
rect 2814 3581 2820 3582
rect 2918 3586 2924 3587
rect 2918 3582 2919 3586
rect 2923 3582 2924 3586
rect 2918 3581 2924 3582
rect 3014 3586 3020 3587
rect 3014 3582 3015 3586
rect 3019 3582 3020 3586
rect 3014 3581 3020 3582
rect 3110 3586 3116 3587
rect 3110 3582 3111 3586
rect 3115 3582 3116 3586
rect 3110 3581 3116 3582
rect 3206 3586 3212 3587
rect 3206 3582 3207 3586
rect 3211 3582 3212 3586
rect 3206 3581 3212 3582
rect 3302 3586 3308 3587
rect 3302 3582 3303 3586
rect 3307 3582 3308 3586
rect 3302 3581 3308 3582
rect 3398 3586 3404 3587
rect 3398 3582 3399 3586
rect 3403 3582 3404 3586
rect 3398 3581 3404 3582
rect 142 3578 148 3579
rect 142 3574 143 3578
rect 147 3574 148 3578
rect 142 3573 148 3574
rect 222 3578 228 3579
rect 222 3574 223 3578
rect 227 3574 228 3578
rect 222 3573 228 3574
rect 342 3578 348 3579
rect 342 3574 343 3578
rect 347 3574 348 3578
rect 342 3573 348 3574
rect 470 3578 476 3579
rect 470 3574 471 3578
rect 475 3574 476 3578
rect 470 3573 476 3574
rect 606 3578 612 3579
rect 606 3574 607 3578
rect 611 3574 612 3578
rect 606 3573 612 3574
rect 742 3578 748 3579
rect 742 3574 743 3578
rect 747 3574 748 3578
rect 742 3573 748 3574
rect 878 3578 884 3579
rect 878 3574 879 3578
rect 883 3574 884 3578
rect 878 3573 884 3574
rect 998 3578 1004 3579
rect 998 3574 999 3578
rect 1003 3574 1004 3578
rect 998 3573 1004 3574
rect 1110 3578 1116 3579
rect 1110 3574 1111 3578
rect 1115 3574 1116 3578
rect 1110 3573 1116 3574
rect 1222 3578 1228 3579
rect 1222 3574 1223 3578
rect 1227 3574 1228 3578
rect 1222 3573 1228 3574
rect 1326 3578 1332 3579
rect 1326 3574 1327 3578
rect 1331 3574 1332 3578
rect 1326 3573 1332 3574
rect 1422 3578 1428 3579
rect 1422 3574 1423 3578
rect 1427 3574 1428 3578
rect 1422 3573 1428 3574
rect 1526 3578 1532 3579
rect 1526 3574 1527 3578
rect 1531 3574 1532 3578
rect 1526 3573 1532 3574
rect 1630 3578 1636 3579
rect 1630 3574 1631 3578
rect 1635 3574 1636 3578
rect 1630 3573 1636 3574
rect 1870 3568 1876 3569
rect 1870 3564 1871 3568
rect 1875 3564 1876 3568
rect 1870 3563 1876 3564
rect 3590 3568 3596 3569
rect 3590 3564 3591 3568
rect 3595 3564 3596 3568
rect 3590 3563 3596 3564
rect 110 3560 116 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 1830 3560 1836 3561
rect 1830 3556 1831 3560
rect 1835 3556 1836 3560
rect 1830 3555 1836 3556
rect 2114 3559 2120 3560
rect 2114 3555 2115 3559
rect 2119 3555 2120 3559
rect 2114 3554 2120 3555
rect 2202 3559 2208 3560
rect 2202 3555 2203 3559
rect 2207 3555 2208 3559
rect 2202 3554 2208 3555
rect 2306 3559 2312 3560
rect 2306 3555 2307 3559
rect 2311 3555 2312 3559
rect 2306 3554 2312 3555
rect 2418 3559 2424 3560
rect 2418 3555 2419 3559
rect 2423 3555 2424 3559
rect 2418 3554 2424 3555
rect 2530 3559 2536 3560
rect 2530 3555 2531 3559
rect 2535 3555 2536 3559
rect 2530 3554 2536 3555
rect 2754 3559 2760 3560
rect 2754 3555 2755 3559
rect 2759 3555 2760 3559
rect 2754 3554 2760 3555
rect 2866 3559 2872 3560
rect 2866 3555 2867 3559
rect 2871 3555 2872 3559
rect 2866 3554 2872 3555
rect 2970 3559 2976 3560
rect 2970 3555 2971 3559
rect 2975 3555 2976 3559
rect 2970 3554 2976 3555
rect 3066 3559 3072 3560
rect 3066 3555 3067 3559
rect 3071 3555 3072 3559
rect 3066 3554 3072 3555
rect 3162 3559 3168 3560
rect 3162 3555 3163 3559
rect 3167 3555 3168 3559
rect 3162 3554 3168 3555
rect 3258 3559 3264 3560
rect 3258 3555 3259 3559
rect 3263 3555 3264 3559
rect 3258 3554 3264 3555
rect 3354 3559 3360 3560
rect 3354 3555 3355 3559
rect 3359 3555 3360 3559
rect 3354 3554 3360 3555
rect 194 3551 200 3552
rect 194 3547 195 3551
rect 199 3547 200 3551
rect 194 3546 200 3547
rect 274 3551 280 3552
rect 274 3547 275 3551
rect 279 3547 280 3551
rect 274 3546 280 3547
rect 394 3551 400 3552
rect 394 3547 395 3551
rect 399 3547 400 3551
rect 394 3546 400 3547
rect 522 3551 528 3552
rect 522 3547 523 3551
rect 527 3547 528 3551
rect 522 3546 528 3547
rect 658 3551 664 3552
rect 658 3547 659 3551
rect 663 3547 664 3551
rect 658 3546 664 3547
rect 766 3551 772 3552
rect 766 3547 767 3551
rect 771 3547 772 3551
rect 766 3546 772 3547
rect 930 3551 936 3552
rect 930 3547 931 3551
rect 935 3547 936 3551
rect 930 3546 936 3547
rect 1050 3551 1056 3552
rect 1050 3547 1051 3551
rect 1055 3547 1056 3551
rect 1050 3546 1056 3547
rect 1162 3551 1168 3552
rect 1162 3547 1163 3551
rect 1167 3547 1168 3551
rect 1162 3546 1168 3547
rect 1274 3551 1280 3552
rect 1274 3547 1275 3551
rect 1279 3547 1280 3551
rect 1274 3546 1280 3547
rect 1378 3551 1384 3552
rect 1378 3547 1379 3551
rect 1383 3547 1384 3551
rect 1378 3546 1384 3547
rect 1474 3551 1480 3552
rect 1474 3547 1475 3551
rect 1479 3547 1480 3551
rect 1474 3546 1480 3547
rect 1578 3551 1584 3552
rect 1578 3547 1579 3551
rect 1583 3547 1584 3551
rect 1578 3546 1584 3547
rect 1870 3551 1876 3552
rect 1870 3547 1871 3551
rect 1875 3547 1876 3551
rect 3590 3551 3596 3552
rect 1870 3546 1876 3547
rect 2054 3548 2060 3549
rect 2054 3544 2055 3548
rect 2059 3544 2060 3548
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 1830 3543 1836 3544
rect 2054 3543 2060 3544
rect 2142 3548 2148 3549
rect 2142 3544 2143 3548
rect 2147 3544 2148 3548
rect 2142 3543 2148 3544
rect 2246 3548 2252 3549
rect 2246 3544 2247 3548
rect 2251 3544 2252 3548
rect 2246 3543 2252 3544
rect 2358 3548 2364 3549
rect 2358 3544 2359 3548
rect 2363 3544 2364 3548
rect 2358 3543 2364 3544
rect 2470 3548 2476 3549
rect 2470 3544 2471 3548
rect 2475 3544 2476 3548
rect 2470 3543 2476 3544
rect 2582 3548 2588 3549
rect 2582 3544 2583 3548
rect 2587 3544 2588 3548
rect 2582 3543 2588 3544
rect 2694 3548 2700 3549
rect 2694 3544 2695 3548
rect 2699 3544 2700 3548
rect 2694 3543 2700 3544
rect 2806 3548 2812 3549
rect 2806 3544 2807 3548
rect 2811 3544 2812 3548
rect 2806 3543 2812 3544
rect 2910 3548 2916 3549
rect 2910 3544 2911 3548
rect 2915 3544 2916 3548
rect 2910 3543 2916 3544
rect 3006 3548 3012 3549
rect 3006 3544 3007 3548
rect 3011 3544 3012 3548
rect 3006 3543 3012 3544
rect 3102 3548 3108 3549
rect 3102 3544 3103 3548
rect 3107 3544 3108 3548
rect 3102 3543 3108 3544
rect 3198 3548 3204 3549
rect 3198 3544 3199 3548
rect 3203 3544 3204 3548
rect 3198 3543 3204 3544
rect 3294 3548 3300 3549
rect 3294 3544 3295 3548
rect 3299 3544 3300 3548
rect 3294 3543 3300 3544
rect 3390 3548 3396 3549
rect 3390 3544 3391 3548
rect 3395 3544 3396 3548
rect 3590 3547 3591 3551
rect 3595 3547 3596 3551
rect 3590 3546 3596 3547
rect 3390 3543 3396 3544
rect 110 3538 116 3539
rect 134 3540 140 3541
rect 134 3536 135 3540
rect 139 3536 140 3540
rect 134 3535 140 3536
rect 214 3540 220 3541
rect 214 3536 215 3540
rect 219 3536 220 3540
rect 214 3535 220 3536
rect 334 3540 340 3541
rect 334 3536 335 3540
rect 339 3536 340 3540
rect 334 3535 340 3536
rect 462 3540 468 3541
rect 462 3536 463 3540
rect 467 3536 468 3540
rect 462 3535 468 3536
rect 598 3540 604 3541
rect 598 3536 599 3540
rect 603 3536 604 3540
rect 598 3535 604 3536
rect 734 3540 740 3541
rect 734 3536 735 3540
rect 739 3536 740 3540
rect 734 3535 740 3536
rect 870 3540 876 3541
rect 870 3536 871 3540
rect 875 3536 876 3540
rect 870 3535 876 3536
rect 990 3540 996 3541
rect 990 3536 991 3540
rect 995 3536 996 3540
rect 990 3535 996 3536
rect 1102 3540 1108 3541
rect 1102 3536 1103 3540
rect 1107 3536 1108 3540
rect 1102 3535 1108 3536
rect 1214 3540 1220 3541
rect 1214 3536 1215 3540
rect 1219 3536 1220 3540
rect 1214 3535 1220 3536
rect 1318 3540 1324 3541
rect 1318 3536 1319 3540
rect 1323 3536 1324 3540
rect 1318 3535 1324 3536
rect 1414 3540 1420 3541
rect 1414 3536 1415 3540
rect 1419 3536 1420 3540
rect 1414 3535 1420 3536
rect 1518 3540 1524 3541
rect 1518 3536 1519 3540
rect 1523 3536 1524 3540
rect 1518 3535 1524 3536
rect 1622 3540 1628 3541
rect 1622 3536 1623 3540
rect 1627 3536 1628 3540
rect 1830 3539 1831 3543
rect 1835 3539 1836 3543
rect 1830 3538 1836 3539
rect 1622 3535 1628 3536
rect 2382 3531 2388 3532
rect 2382 3527 2383 3531
rect 2387 3530 2388 3531
rect 2599 3531 2605 3532
rect 2599 3530 2600 3531
rect 2387 3528 2600 3530
rect 2387 3527 2388 3528
rect 2382 3526 2388 3527
rect 2599 3527 2600 3528
rect 2604 3527 2605 3531
rect 2599 3526 2605 3527
rect 3134 3531 3140 3532
rect 3134 3527 3135 3531
rect 3139 3530 3140 3531
rect 3407 3531 3413 3532
rect 3407 3530 3408 3531
rect 3139 3528 3408 3530
rect 3139 3527 3140 3528
rect 3134 3526 3140 3527
rect 3407 3527 3408 3528
rect 3412 3527 3413 3531
rect 3407 3526 3413 3527
rect 1582 3523 1588 3524
rect 1582 3519 1583 3523
rect 1587 3522 1588 3523
rect 1639 3523 1645 3524
rect 1639 3522 1640 3523
rect 1587 3520 1640 3522
rect 1587 3519 1588 3520
rect 1582 3518 1588 3519
rect 1639 3519 1640 3520
rect 1644 3519 1645 3523
rect 1639 3518 1645 3519
rect 2086 3504 2092 3505
rect 1870 3501 1876 3502
rect 1870 3497 1871 3501
rect 1875 3497 1876 3501
rect 2086 3500 2087 3504
rect 2091 3500 2092 3504
rect 2086 3499 2092 3500
rect 2166 3504 2172 3505
rect 2166 3500 2167 3504
rect 2171 3500 2172 3504
rect 2166 3499 2172 3500
rect 2262 3504 2268 3505
rect 2262 3500 2263 3504
rect 2267 3500 2268 3504
rect 2262 3499 2268 3500
rect 2366 3504 2372 3505
rect 2366 3500 2367 3504
rect 2371 3500 2372 3504
rect 2366 3499 2372 3500
rect 2486 3504 2492 3505
rect 2486 3500 2487 3504
rect 2491 3500 2492 3504
rect 2486 3499 2492 3500
rect 2614 3504 2620 3505
rect 2614 3500 2615 3504
rect 2619 3500 2620 3504
rect 2614 3499 2620 3500
rect 2742 3504 2748 3505
rect 2742 3500 2743 3504
rect 2747 3500 2748 3504
rect 2742 3499 2748 3500
rect 2870 3504 2876 3505
rect 2870 3500 2871 3504
rect 2875 3500 2876 3504
rect 2870 3499 2876 3500
rect 2990 3504 2996 3505
rect 2990 3500 2991 3504
rect 2995 3500 2996 3504
rect 2990 3499 2996 3500
rect 3118 3504 3124 3505
rect 3118 3500 3119 3504
rect 3123 3500 3124 3504
rect 3118 3499 3124 3500
rect 3246 3504 3252 3505
rect 3246 3500 3247 3504
rect 3251 3500 3252 3504
rect 3246 3499 3252 3500
rect 3374 3504 3380 3505
rect 3374 3500 3375 3504
rect 3379 3500 3380 3504
rect 3374 3499 3380 3500
rect 3590 3501 3596 3502
rect 190 3496 196 3497
rect 110 3493 116 3494
rect 110 3489 111 3493
rect 115 3489 116 3493
rect 190 3492 191 3496
rect 195 3492 196 3496
rect 190 3491 196 3492
rect 326 3496 332 3497
rect 326 3492 327 3496
rect 331 3492 332 3496
rect 326 3491 332 3492
rect 470 3496 476 3497
rect 470 3492 471 3496
rect 475 3492 476 3496
rect 470 3491 476 3492
rect 622 3496 628 3497
rect 622 3492 623 3496
rect 627 3492 628 3496
rect 622 3491 628 3492
rect 774 3496 780 3497
rect 774 3492 775 3496
rect 779 3492 780 3496
rect 774 3491 780 3492
rect 918 3496 924 3497
rect 918 3492 919 3496
rect 923 3492 924 3496
rect 918 3491 924 3492
rect 1054 3496 1060 3497
rect 1054 3492 1055 3496
rect 1059 3492 1060 3496
rect 1054 3491 1060 3492
rect 1182 3496 1188 3497
rect 1182 3492 1183 3496
rect 1187 3492 1188 3496
rect 1182 3491 1188 3492
rect 1310 3496 1316 3497
rect 1310 3492 1311 3496
rect 1315 3492 1316 3496
rect 1310 3491 1316 3492
rect 1438 3496 1444 3497
rect 1438 3492 1439 3496
rect 1443 3492 1444 3496
rect 1438 3491 1444 3492
rect 1566 3496 1572 3497
rect 1870 3496 1876 3497
rect 3590 3497 3591 3501
rect 3595 3497 3596 3501
rect 3590 3496 3596 3497
rect 1566 3492 1567 3496
rect 1571 3492 1572 3496
rect 2070 3495 2076 3496
rect 1566 3491 1572 3492
rect 1830 3493 1836 3494
rect 110 3488 116 3489
rect 1830 3489 1831 3493
rect 1835 3489 1836 3493
rect 2070 3491 2071 3495
rect 2075 3494 2076 3495
rect 2154 3495 2160 3496
rect 2075 3492 2105 3494
rect 2075 3491 2076 3492
rect 2070 3490 2076 3491
rect 2154 3491 2155 3495
rect 2159 3494 2160 3495
rect 2234 3495 2240 3496
rect 2159 3492 2185 3494
rect 2159 3491 2160 3492
rect 2154 3490 2160 3491
rect 2234 3491 2235 3495
rect 2239 3494 2240 3495
rect 2434 3495 2440 3496
rect 2434 3494 2435 3495
rect 2239 3492 2281 3494
rect 2429 3492 2435 3494
rect 2239 3491 2240 3492
rect 2234 3490 2240 3491
rect 2434 3491 2435 3492
rect 2439 3491 2440 3495
rect 2558 3495 2564 3496
rect 2558 3494 2559 3495
rect 2549 3492 2559 3494
rect 2434 3490 2440 3491
rect 2558 3491 2559 3492
rect 2563 3491 2564 3495
rect 2686 3495 2692 3496
rect 2686 3494 2687 3495
rect 2677 3492 2687 3494
rect 2558 3490 2564 3491
rect 2686 3491 2687 3492
rect 2691 3491 2692 3495
rect 2815 3495 2821 3496
rect 2815 3494 2816 3495
rect 2805 3492 2816 3494
rect 2686 3490 2692 3491
rect 2815 3491 2816 3492
rect 2820 3491 2821 3495
rect 2815 3490 2821 3491
rect 2826 3495 2832 3496
rect 2826 3491 2827 3495
rect 2831 3494 2832 3495
rect 2938 3495 2944 3496
rect 2831 3492 2889 3494
rect 2831 3491 2832 3492
rect 2826 3490 2832 3491
rect 2938 3491 2939 3495
rect 2943 3494 2944 3495
rect 3191 3495 3197 3496
rect 3191 3494 3192 3495
rect 2943 3492 3009 3494
rect 3181 3492 3192 3494
rect 2943 3491 2944 3492
rect 2938 3490 2944 3491
rect 3191 3491 3192 3492
rect 3196 3491 3197 3495
rect 3318 3495 3324 3496
rect 3318 3494 3319 3495
rect 3309 3492 3319 3494
rect 3191 3490 3197 3491
rect 3318 3491 3319 3492
rect 3323 3491 3324 3495
rect 3318 3490 3324 3491
rect 1830 3488 1836 3489
rect 3436 3488 3438 3493
rect 151 3487 157 3488
rect 151 3483 152 3487
rect 156 3486 157 3487
rect 258 3487 264 3488
rect 156 3484 209 3486
rect 156 3483 157 3484
rect 151 3482 157 3483
rect 258 3483 259 3487
rect 263 3486 264 3487
rect 394 3487 400 3488
rect 263 3484 345 3486
rect 263 3483 264 3484
rect 258 3482 264 3483
rect 394 3483 395 3487
rect 399 3486 400 3487
rect 538 3487 544 3488
rect 399 3484 489 3486
rect 399 3483 400 3484
rect 394 3482 400 3483
rect 538 3483 539 3487
rect 543 3486 544 3487
rect 690 3487 696 3488
rect 543 3484 641 3486
rect 543 3483 544 3484
rect 538 3482 544 3483
rect 690 3483 691 3487
rect 695 3486 696 3487
rect 886 3487 892 3488
rect 695 3484 793 3486
rect 695 3483 696 3484
rect 690 3482 696 3483
rect 886 3483 887 3487
rect 891 3486 892 3487
rect 986 3487 992 3488
rect 891 3484 937 3486
rect 891 3483 892 3484
rect 886 3482 892 3483
rect 986 3483 987 3487
rect 991 3486 992 3487
rect 1126 3487 1132 3488
rect 991 3484 1073 3486
rect 991 3483 992 3484
rect 986 3482 992 3483
rect 1126 3483 1127 3487
rect 1131 3486 1132 3487
rect 1271 3487 1277 3488
rect 1131 3484 1201 3486
rect 1131 3483 1132 3484
rect 1126 3482 1132 3483
rect 1271 3483 1272 3487
rect 1276 3486 1277 3487
rect 1378 3487 1384 3488
rect 1276 3484 1329 3486
rect 1276 3483 1277 3484
rect 1271 3482 1277 3483
rect 1378 3483 1379 3487
rect 1383 3486 1384 3487
rect 1519 3487 1525 3488
rect 1383 3484 1457 3486
rect 1383 3483 1384 3484
rect 1378 3482 1384 3483
rect 1519 3483 1520 3487
rect 1524 3486 1525 3487
rect 3434 3487 3440 3488
rect 1524 3484 1585 3486
rect 1870 3484 1876 3485
rect 1524 3483 1525 3484
rect 1519 3482 1525 3483
rect 1870 3480 1871 3484
rect 1875 3480 1876 3484
rect 3434 3483 3435 3487
rect 3439 3483 3440 3487
rect 3434 3482 3440 3483
rect 3590 3484 3596 3485
rect 1870 3479 1876 3480
rect 3590 3480 3591 3484
rect 3595 3480 3596 3484
rect 3590 3479 3596 3480
rect 110 3476 116 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 110 3471 116 3472
rect 1830 3476 1836 3477
rect 1830 3472 1831 3476
rect 1835 3472 1836 3476
rect 1830 3471 1836 3472
rect 2094 3466 2100 3467
rect 2094 3462 2095 3466
rect 2099 3462 2100 3466
rect 2094 3461 2100 3462
rect 2174 3466 2180 3467
rect 2174 3462 2175 3466
rect 2179 3462 2180 3466
rect 2174 3461 2180 3462
rect 2270 3466 2276 3467
rect 2270 3462 2271 3466
rect 2275 3462 2276 3466
rect 2270 3461 2276 3462
rect 2374 3466 2380 3467
rect 2374 3462 2375 3466
rect 2379 3462 2380 3466
rect 2374 3461 2380 3462
rect 2494 3466 2500 3467
rect 2494 3462 2495 3466
rect 2499 3462 2500 3466
rect 2494 3461 2500 3462
rect 2622 3466 2628 3467
rect 2622 3462 2623 3466
rect 2627 3462 2628 3466
rect 2622 3461 2628 3462
rect 2750 3466 2756 3467
rect 2750 3462 2751 3466
rect 2755 3462 2756 3466
rect 2750 3461 2756 3462
rect 2878 3466 2884 3467
rect 2878 3462 2879 3466
rect 2883 3462 2884 3466
rect 2878 3461 2884 3462
rect 2998 3466 3004 3467
rect 2998 3462 2999 3466
rect 3003 3462 3004 3466
rect 2998 3461 3004 3462
rect 3126 3466 3132 3467
rect 3126 3462 3127 3466
rect 3131 3462 3132 3466
rect 3126 3461 3132 3462
rect 3254 3466 3260 3467
rect 3254 3462 3255 3466
rect 3259 3462 3260 3466
rect 3254 3461 3260 3462
rect 3382 3466 3388 3467
rect 3382 3462 3383 3466
rect 3387 3462 3388 3466
rect 3382 3461 3388 3462
rect 198 3458 204 3459
rect 198 3454 199 3458
rect 203 3454 204 3458
rect 198 3453 204 3454
rect 334 3458 340 3459
rect 334 3454 335 3458
rect 339 3454 340 3458
rect 334 3453 340 3454
rect 478 3458 484 3459
rect 478 3454 479 3458
rect 483 3454 484 3458
rect 478 3453 484 3454
rect 630 3458 636 3459
rect 630 3454 631 3458
rect 635 3454 636 3458
rect 630 3453 636 3454
rect 782 3458 788 3459
rect 782 3454 783 3458
rect 787 3454 788 3458
rect 782 3453 788 3454
rect 926 3458 932 3459
rect 926 3454 927 3458
rect 931 3454 932 3458
rect 926 3453 932 3454
rect 1062 3458 1068 3459
rect 1062 3454 1063 3458
rect 1067 3454 1068 3458
rect 1062 3453 1068 3454
rect 1190 3458 1196 3459
rect 1190 3454 1191 3458
rect 1195 3454 1196 3458
rect 1190 3453 1196 3454
rect 1318 3458 1324 3459
rect 1318 3454 1319 3458
rect 1323 3454 1324 3458
rect 1318 3453 1324 3454
rect 1446 3458 1452 3459
rect 1446 3454 1447 3458
rect 1451 3454 1452 3458
rect 1446 3453 1452 3454
rect 1574 3458 1580 3459
rect 1574 3454 1575 3458
rect 1579 3454 1580 3458
rect 1574 3453 1580 3454
rect 2087 3455 2093 3456
rect 2087 3451 2088 3455
rect 2092 3454 2093 3455
rect 2154 3455 2160 3456
rect 2154 3454 2155 3455
rect 2092 3452 2155 3454
rect 2092 3451 2093 3452
rect 2087 3450 2093 3451
rect 2154 3451 2155 3452
rect 2159 3451 2160 3455
rect 2154 3450 2160 3451
rect 2167 3455 2173 3456
rect 2167 3451 2168 3455
rect 2172 3454 2173 3455
rect 2234 3455 2240 3456
rect 2234 3454 2235 3455
rect 2172 3452 2235 3454
rect 2172 3451 2173 3452
rect 2167 3450 2173 3451
rect 2234 3451 2235 3452
rect 2239 3451 2240 3455
rect 2234 3450 2240 3451
rect 2250 3455 2256 3456
rect 2250 3451 2251 3455
rect 2255 3454 2256 3455
rect 2263 3455 2269 3456
rect 2263 3454 2264 3455
rect 2255 3452 2264 3454
rect 2255 3451 2256 3452
rect 2250 3450 2256 3451
rect 2263 3451 2264 3452
rect 2268 3451 2269 3455
rect 2263 3450 2269 3451
rect 2367 3455 2373 3456
rect 2367 3451 2368 3455
rect 2372 3454 2373 3455
rect 2382 3455 2388 3456
rect 2382 3454 2383 3455
rect 2372 3452 2383 3454
rect 2372 3451 2373 3452
rect 2367 3450 2373 3451
rect 2382 3451 2383 3452
rect 2387 3451 2388 3455
rect 2382 3450 2388 3451
rect 2434 3455 2440 3456
rect 2434 3451 2435 3455
rect 2439 3454 2440 3455
rect 2487 3455 2493 3456
rect 2487 3454 2488 3455
rect 2439 3452 2488 3454
rect 2439 3451 2440 3452
rect 2434 3450 2440 3451
rect 2487 3451 2488 3452
rect 2492 3451 2493 3455
rect 2487 3450 2493 3451
rect 2558 3455 2564 3456
rect 2558 3451 2559 3455
rect 2563 3454 2564 3455
rect 2615 3455 2621 3456
rect 2615 3454 2616 3455
rect 2563 3452 2616 3454
rect 2563 3451 2564 3452
rect 2558 3450 2564 3451
rect 2615 3451 2616 3452
rect 2620 3451 2621 3455
rect 2615 3450 2621 3451
rect 2686 3455 2692 3456
rect 2686 3451 2687 3455
rect 2691 3454 2692 3455
rect 2743 3455 2749 3456
rect 2743 3454 2744 3455
rect 2691 3452 2744 3454
rect 2691 3451 2692 3452
rect 2686 3450 2692 3451
rect 2743 3451 2744 3452
rect 2748 3451 2749 3455
rect 2743 3450 2749 3451
rect 2871 3455 2877 3456
rect 2871 3451 2872 3455
rect 2876 3454 2877 3455
rect 2938 3455 2944 3456
rect 2938 3454 2939 3455
rect 2876 3452 2939 3454
rect 2876 3451 2877 3452
rect 2871 3450 2877 3451
rect 2938 3451 2939 3452
rect 2943 3451 2944 3455
rect 2938 3450 2944 3451
rect 2990 3455 2997 3456
rect 2990 3451 2991 3455
rect 2996 3451 2997 3455
rect 2990 3450 2997 3451
rect 3119 3455 3125 3456
rect 3119 3451 3120 3455
rect 3124 3454 3125 3455
rect 3134 3455 3140 3456
rect 3134 3454 3135 3455
rect 3124 3452 3135 3454
rect 3124 3451 3125 3452
rect 3119 3450 3125 3451
rect 3134 3451 3135 3452
rect 3139 3451 3140 3455
rect 3134 3450 3140 3451
rect 3191 3455 3197 3456
rect 3191 3451 3192 3455
rect 3196 3454 3197 3455
rect 3247 3455 3253 3456
rect 3247 3454 3248 3455
rect 3196 3452 3248 3454
rect 3196 3451 3197 3452
rect 3191 3450 3197 3451
rect 3247 3451 3248 3452
rect 3252 3451 3253 3455
rect 3247 3450 3253 3451
rect 3318 3455 3324 3456
rect 3318 3451 3319 3455
rect 3323 3454 3324 3455
rect 3375 3455 3381 3456
rect 3375 3454 3376 3455
rect 3323 3452 3376 3454
rect 3323 3451 3324 3452
rect 3318 3450 3324 3451
rect 3375 3451 3376 3452
rect 3380 3451 3381 3455
rect 3375 3450 3381 3451
rect 191 3447 197 3448
rect 191 3443 192 3447
rect 196 3446 197 3447
rect 258 3447 264 3448
rect 258 3446 259 3447
rect 196 3444 259 3446
rect 196 3443 197 3444
rect 191 3442 197 3443
rect 258 3443 259 3444
rect 263 3443 264 3447
rect 258 3442 264 3443
rect 327 3447 333 3448
rect 327 3443 328 3447
rect 332 3446 333 3447
rect 394 3447 400 3448
rect 394 3446 395 3447
rect 332 3444 395 3446
rect 332 3443 333 3444
rect 327 3442 333 3443
rect 394 3443 395 3444
rect 399 3443 400 3447
rect 394 3442 400 3443
rect 471 3447 477 3448
rect 471 3443 472 3447
rect 476 3446 477 3447
rect 538 3447 544 3448
rect 538 3446 539 3447
rect 476 3444 539 3446
rect 476 3443 477 3444
rect 471 3442 477 3443
rect 538 3443 539 3444
rect 543 3443 544 3447
rect 538 3442 544 3443
rect 623 3447 629 3448
rect 623 3443 624 3447
rect 628 3446 629 3447
rect 690 3447 696 3448
rect 690 3446 691 3447
rect 628 3444 691 3446
rect 628 3443 629 3444
rect 623 3442 629 3443
rect 690 3443 691 3444
rect 695 3443 696 3447
rect 690 3442 696 3443
rect 766 3447 772 3448
rect 766 3443 767 3447
rect 771 3446 772 3447
rect 775 3447 781 3448
rect 775 3446 776 3447
rect 771 3444 776 3446
rect 771 3443 772 3444
rect 766 3442 772 3443
rect 775 3443 776 3444
rect 780 3443 781 3447
rect 775 3442 781 3443
rect 919 3447 925 3448
rect 919 3443 920 3447
rect 924 3446 925 3447
rect 986 3447 992 3448
rect 986 3446 987 3447
rect 924 3444 987 3446
rect 924 3443 925 3444
rect 919 3442 925 3443
rect 986 3443 987 3444
rect 991 3443 992 3447
rect 986 3442 992 3443
rect 1055 3447 1061 3448
rect 1055 3443 1056 3447
rect 1060 3446 1061 3447
rect 1126 3447 1132 3448
rect 1126 3446 1127 3447
rect 1060 3444 1127 3446
rect 1060 3443 1061 3444
rect 1055 3442 1061 3443
rect 1126 3443 1127 3444
rect 1131 3443 1132 3447
rect 1126 3442 1132 3443
rect 1170 3447 1176 3448
rect 1170 3443 1171 3447
rect 1175 3446 1176 3447
rect 1183 3447 1189 3448
rect 1183 3446 1184 3447
rect 1175 3444 1184 3446
rect 1175 3443 1176 3444
rect 1170 3442 1176 3443
rect 1183 3443 1184 3444
rect 1188 3443 1189 3447
rect 1183 3442 1189 3443
rect 1311 3447 1317 3448
rect 1311 3443 1312 3447
rect 1316 3446 1317 3447
rect 1378 3447 1384 3448
rect 1378 3446 1379 3447
rect 1316 3444 1379 3446
rect 1316 3443 1317 3444
rect 1311 3442 1317 3443
rect 1378 3443 1379 3444
rect 1383 3443 1384 3447
rect 1378 3442 1384 3443
rect 1439 3447 1445 3448
rect 1439 3443 1440 3447
rect 1444 3446 1445 3447
rect 1519 3447 1525 3448
rect 1519 3446 1520 3447
rect 1444 3444 1520 3446
rect 1444 3443 1445 3444
rect 1439 3442 1445 3443
rect 1519 3443 1520 3444
rect 1524 3443 1525 3447
rect 1519 3442 1525 3443
rect 1567 3447 1573 3448
rect 1567 3443 1568 3447
rect 1572 3446 1573 3447
rect 1582 3447 1588 3448
rect 1582 3446 1583 3447
rect 1572 3444 1583 3446
rect 1572 3443 1573 3444
rect 1567 3442 1573 3443
rect 1582 3443 1583 3444
rect 1587 3443 1588 3447
rect 1582 3442 1588 3443
rect 143 3435 149 3436
rect 143 3431 144 3435
rect 148 3434 149 3435
rect 151 3435 157 3436
rect 151 3434 152 3435
rect 148 3432 152 3434
rect 148 3431 149 3432
rect 143 3430 149 3431
rect 151 3431 152 3432
rect 156 3431 157 3435
rect 151 3430 157 3431
rect 286 3435 293 3436
rect 286 3431 287 3435
rect 292 3431 293 3435
rect 286 3430 293 3431
rect 346 3435 352 3436
rect 346 3431 347 3435
rect 351 3434 352 3435
rect 447 3435 453 3436
rect 447 3434 448 3435
rect 351 3432 448 3434
rect 351 3431 352 3432
rect 346 3430 352 3431
rect 447 3431 448 3432
rect 452 3431 453 3435
rect 447 3430 453 3431
rect 506 3435 512 3436
rect 506 3431 507 3435
rect 511 3434 512 3435
rect 615 3435 621 3436
rect 615 3434 616 3435
rect 511 3432 616 3434
rect 511 3431 512 3432
rect 506 3430 512 3431
rect 615 3431 616 3432
rect 620 3431 621 3435
rect 615 3430 621 3431
rect 674 3435 680 3436
rect 674 3431 675 3435
rect 679 3434 680 3435
rect 783 3435 789 3436
rect 783 3434 784 3435
rect 679 3432 784 3434
rect 679 3431 680 3432
rect 674 3430 680 3431
rect 783 3431 784 3432
rect 788 3431 789 3435
rect 783 3430 789 3431
rect 935 3435 941 3436
rect 935 3431 936 3435
rect 940 3434 941 3435
rect 951 3435 957 3436
rect 951 3434 952 3435
rect 940 3432 952 3434
rect 940 3431 941 3432
rect 935 3430 941 3431
rect 951 3431 952 3432
rect 956 3431 957 3435
rect 951 3430 957 3431
rect 1010 3435 1016 3436
rect 1010 3431 1011 3435
rect 1015 3434 1016 3435
rect 1111 3435 1117 3436
rect 1111 3434 1112 3435
rect 1015 3432 1112 3434
rect 1015 3431 1016 3432
rect 1010 3430 1016 3431
rect 1111 3431 1112 3432
rect 1116 3431 1117 3435
rect 1111 3430 1117 3431
rect 1263 3435 1269 3436
rect 1263 3431 1264 3435
rect 1268 3434 1269 3435
rect 1271 3435 1277 3436
rect 1271 3434 1272 3435
rect 1268 3432 1272 3434
rect 1268 3431 1269 3432
rect 1263 3430 1269 3431
rect 1271 3431 1272 3432
rect 1276 3431 1277 3435
rect 1271 3430 1277 3431
rect 1350 3435 1356 3436
rect 1350 3431 1351 3435
rect 1355 3434 1356 3435
rect 1407 3435 1413 3436
rect 1407 3434 1408 3435
rect 1355 3432 1408 3434
rect 1355 3431 1356 3432
rect 1350 3430 1356 3431
rect 1407 3431 1408 3432
rect 1412 3431 1413 3435
rect 1407 3430 1413 3431
rect 1466 3435 1472 3436
rect 1466 3431 1467 3435
rect 1471 3434 1472 3435
rect 1551 3435 1557 3436
rect 1551 3434 1552 3435
rect 1471 3432 1552 3434
rect 1471 3431 1472 3432
rect 1466 3430 1472 3431
rect 1551 3431 1552 3432
rect 1556 3431 1557 3435
rect 1551 3430 1557 3431
rect 1610 3435 1616 3436
rect 1610 3431 1611 3435
rect 1615 3434 1616 3435
rect 1703 3435 1709 3436
rect 1703 3434 1704 3435
rect 1615 3432 1704 3434
rect 1615 3431 1616 3432
rect 1610 3430 1616 3431
rect 1703 3431 1704 3432
rect 1708 3431 1709 3435
rect 1703 3430 1709 3431
rect 2103 3435 2109 3436
rect 2103 3431 2104 3435
rect 2108 3434 2109 3435
rect 2154 3435 2160 3436
rect 2154 3434 2155 3435
rect 2108 3432 2155 3434
rect 2108 3431 2109 3432
rect 2103 3430 2109 3431
rect 2154 3431 2155 3432
rect 2159 3431 2160 3435
rect 2154 3430 2160 3431
rect 2162 3435 2168 3436
rect 2162 3431 2163 3435
rect 2167 3434 2168 3435
rect 2191 3435 2197 3436
rect 2191 3434 2192 3435
rect 2167 3432 2192 3434
rect 2167 3431 2168 3432
rect 2162 3430 2168 3431
rect 2191 3431 2192 3432
rect 2196 3431 2197 3435
rect 2191 3430 2197 3431
rect 2294 3435 2301 3436
rect 2294 3431 2295 3435
rect 2300 3431 2301 3435
rect 2294 3430 2301 3431
rect 2407 3435 2413 3436
rect 2407 3431 2408 3435
rect 2412 3434 2413 3435
rect 2422 3435 2428 3436
rect 2422 3434 2423 3435
rect 2412 3432 2423 3434
rect 2412 3431 2413 3432
rect 2407 3430 2413 3431
rect 2422 3431 2423 3432
rect 2427 3431 2428 3435
rect 2422 3430 2428 3431
rect 2535 3435 2541 3436
rect 2535 3431 2536 3435
rect 2540 3434 2541 3435
rect 2602 3435 2608 3436
rect 2602 3434 2603 3435
rect 2540 3432 2603 3434
rect 2540 3431 2541 3432
rect 2535 3430 2541 3431
rect 2602 3431 2603 3432
rect 2607 3431 2608 3435
rect 2602 3430 2608 3431
rect 2671 3435 2677 3436
rect 2671 3431 2672 3435
rect 2676 3434 2677 3435
rect 2738 3435 2744 3436
rect 2738 3434 2739 3435
rect 2676 3432 2739 3434
rect 2676 3431 2677 3432
rect 2671 3430 2677 3431
rect 2738 3431 2739 3432
rect 2743 3431 2744 3435
rect 2738 3430 2744 3431
rect 2807 3435 2813 3436
rect 2807 3431 2808 3435
rect 2812 3434 2813 3435
rect 2815 3435 2821 3436
rect 2815 3434 2816 3435
rect 2812 3432 2816 3434
rect 2812 3431 2813 3432
rect 2807 3430 2813 3431
rect 2815 3431 2816 3432
rect 2820 3431 2821 3435
rect 2815 3430 2821 3431
rect 2951 3435 2957 3436
rect 2951 3431 2952 3435
rect 2956 3434 2957 3435
rect 3030 3435 3036 3436
rect 3030 3434 3031 3435
rect 2956 3432 3031 3434
rect 2956 3431 2957 3432
rect 2951 3430 2957 3431
rect 3030 3431 3031 3432
rect 3035 3431 3036 3435
rect 3030 3430 3036 3431
rect 3103 3435 3109 3436
rect 3103 3431 3104 3435
rect 3108 3434 3109 3435
rect 3134 3435 3140 3436
rect 3134 3434 3135 3435
rect 3108 3432 3135 3434
rect 3108 3431 3109 3432
rect 3103 3430 3109 3431
rect 3134 3431 3135 3432
rect 3139 3431 3140 3435
rect 3134 3430 3140 3431
rect 3255 3435 3261 3436
rect 3255 3431 3256 3435
rect 3260 3434 3261 3435
rect 3335 3435 3341 3436
rect 3335 3434 3336 3435
rect 3260 3432 3336 3434
rect 3260 3431 3261 3432
rect 3255 3430 3261 3431
rect 3335 3431 3336 3432
rect 3340 3431 3341 3435
rect 3335 3430 3341 3431
rect 3415 3435 3421 3436
rect 3415 3431 3416 3435
rect 3420 3434 3421 3435
rect 3434 3435 3440 3436
rect 3434 3434 3435 3435
rect 3420 3432 3435 3434
rect 3420 3431 3421 3432
rect 3415 3430 3421 3431
rect 3434 3431 3435 3432
rect 3439 3431 3440 3435
rect 3434 3430 3440 3431
rect 150 3426 156 3427
rect 150 3422 151 3426
rect 155 3422 156 3426
rect 150 3421 156 3422
rect 294 3426 300 3427
rect 294 3422 295 3426
rect 299 3422 300 3426
rect 294 3421 300 3422
rect 454 3426 460 3427
rect 454 3422 455 3426
rect 459 3422 460 3426
rect 454 3421 460 3422
rect 622 3426 628 3427
rect 622 3422 623 3426
rect 627 3422 628 3426
rect 622 3421 628 3422
rect 790 3426 796 3427
rect 790 3422 791 3426
rect 795 3422 796 3426
rect 790 3421 796 3422
rect 958 3426 964 3427
rect 958 3422 959 3426
rect 963 3422 964 3426
rect 958 3421 964 3422
rect 1118 3426 1124 3427
rect 1118 3422 1119 3426
rect 1123 3422 1124 3426
rect 1118 3421 1124 3422
rect 1270 3426 1276 3427
rect 1270 3422 1271 3426
rect 1275 3422 1276 3426
rect 1270 3421 1276 3422
rect 1414 3426 1420 3427
rect 1414 3422 1415 3426
rect 1419 3422 1420 3426
rect 1414 3421 1420 3422
rect 1558 3426 1564 3427
rect 1558 3422 1559 3426
rect 1563 3422 1564 3426
rect 1558 3421 1564 3422
rect 1710 3426 1716 3427
rect 1710 3422 1711 3426
rect 1715 3422 1716 3426
rect 1710 3421 1716 3422
rect 2110 3426 2116 3427
rect 2110 3422 2111 3426
rect 2115 3422 2116 3426
rect 2110 3421 2116 3422
rect 2198 3426 2204 3427
rect 2198 3422 2199 3426
rect 2203 3422 2204 3426
rect 2198 3421 2204 3422
rect 2302 3426 2308 3427
rect 2302 3422 2303 3426
rect 2307 3422 2308 3426
rect 2302 3421 2308 3422
rect 2414 3426 2420 3427
rect 2414 3422 2415 3426
rect 2419 3422 2420 3426
rect 2414 3421 2420 3422
rect 2542 3426 2548 3427
rect 2542 3422 2543 3426
rect 2547 3422 2548 3426
rect 2542 3421 2548 3422
rect 2678 3426 2684 3427
rect 2678 3422 2679 3426
rect 2683 3422 2684 3426
rect 2678 3421 2684 3422
rect 2814 3426 2820 3427
rect 2814 3422 2815 3426
rect 2819 3422 2820 3426
rect 2814 3421 2820 3422
rect 2958 3426 2964 3427
rect 2958 3422 2959 3426
rect 2963 3422 2964 3426
rect 2958 3421 2964 3422
rect 3110 3426 3116 3427
rect 3110 3422 3111 3426
rect 3115 3422 3116 3426
rect 3110 3421 3116 3422
rect 3262 3426 3268 3427
rect 3262 3422 3263 3426
rect 3267 3422 3268 3426
rect 3262 3421 3268 3422
rect 3422 3426 3428 3427
rect 3422 3422 3423 3426
rect 3427 3422 3428 3426
rect 3422 3421 3428 3422
rect 110 3408 116 3409
rect 110 3404 111 3408
rect 115 3404 116 3408
rect 110 3403 116 3404
rect 1830 3408 1836 3409
rect 1830 3404 1831 3408
rect 1835 3404 1836 3408
rect 1830 3403 1836 3404
rect 1870 3408 1876 3409
rect 1870 3404 1871 3408
rect 1875 3404 1876 3408
rect 3590 3408 3596 3409
rect 3590 3404 3591 3408
rect 3595 3404 3596 3408
rect 1870 3403 1876 3404
rect 2294 3403 2300 3404
rect 3590 3403 3596 3404
rect 286 3399 292 3400
rect 286 3398 287 3399
rect 205 3396 287 3398
rect 286 3395 287 3396
rect 291 3395 292 3399
rect 286 3394 292 3395
rect 346 3399 352 3400
rect 346 3395 347 3399
rect 351 3395 352 3399
rect 346 3394 352 3395
rect 506 3399 512 3400
rect 506 3395 507 3399
rect 511 3395 512 3399
rect 506 3394 512 3395
rect 674 3399 680 3400
rect 674 3395 675 3399
rect 679 3395 680 3399
rect 674 3394 680 3395
rect 1010 3399 1016 3400
rect 1010 3395 1011 3399
rect 1015 3395 1016 3399
rect 1010 3394 1016 3395
rect 1170 3399 1176 3400
rect 1170 3395 1171 3399
rect 1175 3395 1176 3399
rect 1350 3399 1356 3400
rect 1350 3398 1351 3399
rect 1325 3396 1351 3398
rect 1170 3394 1176 3395
rect 1350 3395 1351 3396
rect 1355 3395 1356 3399
rect 1350 3394 1356 3395
rect 1466 3399 1472 3400
rect 1466 3395 1467 3399
rect 1471 3395 1472 3399
rect 1466 3394 1472 3395
rect 1610 3399 1616 3400
rect 1610 3395 1611 3399
rect 1615 3395 1616 3399
rect 1610 3394 1616 3395
rect 1734 3399 1740 3400
rect 1734 3395 1735 3399
rect 1739 3395 1740 3399
rect 1734 3394 1740 3395
rect 2162 3399 2168 3400
rect 2162 3395 2163 3399
rect 2167 3395 2168 3399
rect 2162 3394 2168 3395
rect 2250 3399 2256 3400
rect 2250 3395 2251 3399
rect 2255 3395 2256 3399
rect 2294 3399 2295 3403
rect 2299 3402 2300 3403
rect 2299 3400 2426 3402
rect 2299 3399 2300 3400
rect 2294 3398 2300 3399
rect 2424 3397 2426 3400
rect 2574 3399 2580 3400
rect 2250 3394 2256 3395
rect 2574 3395 2575 3399
rect 2579 3395 2580 3399
rect 2574 3394 2580 3395
rect 2602 3399 2608 3400
rect 2602 3395 2603 3399
rect 2607 3398 2608 3399
rect 2738 3399 2744 3400
rect 2607 3396 2689 3398
rect 2607 3395 2608 3396
rect 2602 3394 2608 3395
rect 2738 3395 2739 3399
rect 2743 3398 2744 3399
rect 2990 3399 2996 3400
rect 2743 3396 2825 3398
rect 2743 3395 2744 3396
rect 2738 3394 2744 3395
rect 2990 3395 2991 3399
rect 2995 3395 2996 3399
rect 2990 3394 2996 3395
rect 3030 3399 3036 3400
rect 3030 3395 3031 3399
rect 3035 3398 3036 3399
rect 3302 3399 3308 3400
rect 3035 3396 3121 3398
rect 3035 3395 3036 3396
rect 3030 3394 3036 3395
rect 3302 3395 3303 3399
rect 3307 3395 3308 3399
rect 3302 3394 3308 3395
rect 3335 3399 3341 3400
rect 3335 3395 3336 3399
rect 3340 3398 3341 3399
rect 3340 3396 3433 3398
rect 3340 3395 3341 3396
rect 3335 3394 3341 3395
rect 110 3391 116 3392
rect 110 3387 111 3391
rect 115 3387 116 3391
rect 1830 3391 1836 3392
rect 110 3386 116 3387
rect 142 3388 148 3389
rect 142 3384 143 3388
rect 147 3384 148 3388
rect 142 3383 148 3384
rect 286 3388 292 3389
rect 286 3384 287 3388
rect 291 3384 292 3388
rect 286 3383 292 3384
rect 446 3388 452 3389
rect 446 3384 447 3388
rect 451 3384 452 3388
rect 446 3383 452 3384
rect 614 3388 620 3389
rect 614 3384 615 3388
rect 619 3384 620 3388
rect 614 3383 620 3384
rect 782 3388 788 3389
rect 782 3384 783 3388
rect 787 3384 788 3388
rect 782 3383 788 3384
rect 950 3388 956 3389
rect 950 3384 951 3388
rect 955 3384 956 3388
rect 950 3383 956 3384
rect 1110 3388 1116 3389
rect 1110 3384 1111 3388
rect 1115 3384 1116 3388
rect 1110 3383 1116 3384
rect 1262 3388 1268 3389
rect 1262 3384 1263 3388
rect 1267 3384 1268 3388
rect 1262 3383 1268 3384
rect 1406 3388 1412 3389
rect 1406 3384 1407 3388
rect 1411 3384 1412 3388
rect 1406 3383 1412 3384
rect 1550 3388 1556 3389
rect 1550 3384 1551 3388
rect 1555 3384 1556 3388
rect 1550 3383 1556 3384
rect 1702 3388 1708 3389
rect 1702 3384 1703 3388
rect 1707 3384 1708 3388
rect 1830 3387 1831 3391
rect 1835 3387 1836 3391
rect 1830 3386 1836 3387
rect 1870 3391 1876 3392
rect 1870 3387 1871 3391
rect 1875 3387 1876 3391
rect 3590 3391 3596 3392
rect 1870 3386 1876 3387
rect 2102 3388 2108 3389
rect 1702 3383 1708 3384
rect 2102 3384 2103 3388
rect 2107 3384 2108 3388
rect 2102 3383 2108 3384
rect 2190 3388 2196 3389
rect 2190 3384 2191 3388
rect 2195 3384 2196 3388
rect 2190 3383 2196 3384
rect 2294 3388 2300 3389
rect 2294 3384 2295 3388
rect 2299 3384 2300 3388
rect 2294 3383 2300 3384
rect 2406 3388 2412 3389
rect 2406 3384 2407 3388
rect 2411 3384 2412 3388
rect 2406 3383 2412 3384
rect 2534 3388 2540 3389
rect 2534 3384 2535 3388
rect 2539 3384 2540 3388
rect 2534 3383 2540 3384
rect 2670 3388 2676 3389
rect 2670 3384 2671 3388
rect 2675 3384 2676 3388
rect 2670 3383 2676 3384
rect 2806 3388 2812 3389
rect 2806 3384 2807 3388
rect 2811 3384 2812 3388
rect 2806 3383 2812 3384
rect 2950 3388 2956 3389
rect 2950 3384 2951 3388
rect 2955 3384 2956 3388
rect 2950 3383 2956 3384
rect 3102 3388 3108 3389
rect 3102 3384 3103 3388
rect 3107 3384 3108 3388
rect 3102 3383 3108 3384
rect 3254 3388 3260 3389
rect 3254 3384 3255 3388
rect 3259 3384 3260 3388
rect 3254 3383 3260 3384
rect 3414 3388 3420 3389
rect 3414 3384 3415 3388
rect 3419 3384 3420 3388
rect 3590 3387 3591 3391
rect 3595 3387 3596 3391
rect 3590 3386 3596 3387
rect 3414 3383 3420 3384
rect 678 3371 684 3372
rect 678 3367 679 3371
rect 683 3370 684 3371
rect 799 3371 805 3372
rect 799 3370 800 3371
rect 683 3368 800 3370
rect 683 3367 684 3368
rect 678 3366 684 3367
rect 799 3367 800 3368
rect 804 3367 805 3371
rect 799 3366 805 3367
rect 2154 3371 2160 3372
rect 2154 3367 2155 3371
rect 2159 3370 2160 3371
rect 2311 3371 2317 3372
rect 2311 3370 2312 3371
rect 2159 3368 2312 3370
rect 2159 3367 2160 3368
rect 2154 3366 2160 3367
rect 2311 3367 2312 3368
rect 2316 3367 2317 3371
rect 2311 3366 2317 3367
rect 206 3344 212 3345
rect 110 3341 116 3342
rect 110 3337 111 3341
rect 115 3337 116 3341
rect 206 3340 207 3344
rect 211 3340 212 3344
rect 206 3339 212 3340
rect 334 3344 340 3345
rect 334 3340 335 3344
rect 339 3340 340 3344
rect 334 3339 340 3340
rect 470 3344 476 3345
rect 470 3340 471 3344
rect 475 3340 476 3344
rect 470 3339 476 3340
rect 622 3344 628 3345
rect 622 3340 623 3344
rect 627 3340 628 3344
rect 622 3339 628 3340
rect 782 3344 788 3345
rect 782 3340 783 3344
rect 787 3340 788 3344
rect 782 3339 788 3340
rect 942 3344 948 3345
rect 942 3340 943 3344
rect 947 3340 948 3344
rect 942 3339 948 3340
rect 1102 3344 1108 3345
rect 1102 3340 1103 3344
rect 1107 3340 1108 3344
rect 1102 3339 1108 3340
rect 1262 3344 1268 3345
rect 1262 3340 1263 3344
rect 1267 3340 1268 3344
rect 1262 3339 1268 3340
rect 1422 3344 1428 3345
rect 1422 3340 1423 3344
rect 1427 3340 1428 3344
rect 1422 3339 1428 3340
rect 1582 3344 1588 3345
rect 1582 3340 1583 3344
rect 1587 3340 1588 3344
rect 1582 3339 1588 3340
rect 1742 3344 1748 3345
rect 1742 3340 1743 3344
rect 1747 3340 1748 3344
rect 1742 3339 1748 3340
rect 1830 3341 1836 3342
rect 110 3336 116 3337
rect 1830 3337 1831 3341
rect 1835 3337 1836 3341
rect 2126 3340 2132 3341
rect 1830 3336 1836 3337
rect 1870 3337 1876 3338
rect 278 3335 284 3336
rect 278 3334 279 3335
rect 269 3332 279 3334
rect 278 3331 279 3332
rect 283 3331 284 3335
rect 410 3335 416 3336
rect 410 3334 411 3335
rect 397 3332 411 3334
rect 278 3330 284 3331
rect 410 3331 411 3332
rect 415 3331 416 3335
rect 551 3335 557 3336
rect 551 3334 552 3335
rect 533 3332 552 3334
rect 410 3330 416 3331
rect 551 3331 552 3332
rect 556 3331 557 3335
rect 706 3335 712 3336
rect 706 3334 707 3335
rect 685 3332 707 3334
rect 551 3330 557 3331
rect 706 3331 707 3332
rect 711 3331 712 3335
rect 935 3335 941 3336
rect 706 3330 712 3331
rect 394 3327 400 3328
rect 110 3324 116 3325
rect 110 3320 111 3324
rect 115 3320 116 3324
rect 394 3323 395 3327
rect 399 3326 400 3327
rect 800 3326 802 3333
rect 935 3331 936 3335
rect 940 3334 941 3335
rect 1010 3335 1016 3336
rect 940 3332 961 3334
rect 940 3331 941 3332
rect 935 3330 941 3331
rect 1010 3331 1011 3335
rect 1015 3334 1016 3335
rect 1170 3335 1176 3336
rect 1015 3332 1121 3334
rect 1015 3331 1016 3332
rect 1010 3330 1016 3331
rect 1170 3331 1171 3335
rect 1175 3334 1176 3335
rect 1383 3335 1389 3336
rect 1175 3332 1281 3334
rect 1175 3331 1176 3332
rect 1170 3330 1176 3331
rect 1383 3331 1384 3335
rect 1388 3334 1389 3335
rect 1527 3335 1533 3336
rect 1388 3332 1441 3334
rect 1388 3331 1389 3332
rect 1383 3330 1389 3331
rect 1527 3331 1528 3335
rect 1532 3334 1533 3335
rect 1650 3335 1656 3336
rect 1532 3332 1601 3334
rect 1532 3331 1533 3332
rect 1527 3330 1533 3331
rect 1650 3331 1651 3335
rect 1655 3334 1656 3335
rect 1655 3332 1761 3334
rect 1870 3333 1871 3337
rect 1875 3333 1876 3337
rect 2126 3336 2127 3340
rect 2131 3336 2132 3340
rect 2126 3335 2132 3336
rect 2222 3340 2228 3341
rect 2222 3336 2223 3340
rect 2227 3336 2228 3340
rect 2222 3335 2228 3336
rect 2334 3340 2340 3341
rect 2334 3336 2335 3340
rect 2339 3336 2340 3340
rect 2334 3335 2340 3336
rect 2454 3340 2460 3341
rect 2454 3336 2455 3340
rect 2459 3336 2460 3340
rect 2454 3335 2460 3336
rect 2582 3340 2588 3341
rect 2582 3336 2583 3340
rect 2587 3336 2588 3340
rect 2582 3335 2588 3336
rect 2718 3340 2724 3341
rect 2718 3336 2719 3340
rect 2723 3336 2724 3340
rect 2718 3335 2724 3336
rect 2862 3340 2868 3341
rect 2862 3336 2863 3340
rect 2867 3336 2868 3340
rect 2862 3335 2868 3336
rect 3006 3340 3012 3341
rect 3006 3336 3007 3340
rect 3011 3336 3012 3340
rect 3006 3335 3012 3336
rect 3158 3340 3164 3341
rect 3158 3336 3159 3340
rect 3163 3336 3164 3340
rect 3158 3335 3164 3336
rect 3310 3340 3316 3341
rect 3310 3336 3311 3340
rect 3315 3336 3316 3340
rect 3310 3335 3316 3336
rect 3470 3340 3476 3341
rect 3470 3336 3471 3340
rect 3475 3336 3476 3340
rect 3470 3335 3476 3336
rect 3590 3337 3596 3338
rect 1870 3332 1876 3333
rect 3590 3333 3591 3337
rect 3595 3333 3596 3337
rect 3590 3332 3596 3333
rect 1655 3331 1656 3332
rect 1650 3330 1656 3331
rect 2194 3331 2200 3332
rect 2194 3330 2195 3331
rect 2189 3328 2195 3330
rect 2194 3327 2195 3328
rect 2199 3327 2200 3331
rect 2290 3331 2296 3332
rect 2290 3330 2291 3331
rect 2285 3328 2291 3330
rect 2194 3326 2200 3327
rect 2290 3327 2291 3328
rect 2295 3327 2296 3331
rect 2402 3331 2408 3332
rect 2402 3330 2403 3331
rect 2397 3328 2403 3330
rect 2290 3326 2296 3327
rect 2402 3327 2403 3328
rect 2407 3327 2408 3331
rect 2402 3326 2408 3327
rect 2422 3331 2428 3332
rect 2422 3327 2423 3331
rect 2427 3330 2428 3331
rect 2650 3331 2656 3332
rect 2650 3330 2651 3331
rect 2427 3328 2473 3330
rect 2645 3328 2651 3330
rect 2427 3327 2428 3328
rect 2422 3326 2428 3327
rect 2650 3327 2651 3328
rect 2655 3327 2656 3331
rect 2798 3331 2804 3332
rect 2798 3330 2799 3331
rect 2781 3328 2799 3330
rect 2650 3326 2656 3327
rect 2798 3327 2799 3328
rect 2803 3327 2804 3331
rect 2798 3326 2804 3327
rect 2823 3331 2829 3332
rect 2823 3327 2824 3331
rect 2828 3330 2829 3331
rect 3079 3331 3085 3332
rect 3079 3330 3080 3331
rect 2828 3328 2881 3330
rect 3069 3328 3080 3330
rect 2828 3327 2829 3328
rect 2823 3326 2829 3327
rect 3079 3327 3080 3328
rect 3084 3327 3085 3331
rect 3079 3326 3085 3327
rect 3134 3331 3140 3332
rect 3134 3327 3135 3331
rect 3139 3330 3140 3331
rect 3394 3331 3400 3332
rect 3394 3330 3395 3331
rect 3139 3328 3177 3330
rect 3373 3328 3395 3330
rect 3139 3327 3140 3328
rect 3134 3326 3140 3327
rect 3394 3327 3395 3328
rect 3399 3327 3400 3331
rect 3394 3326 3400 3327
rect 399 3324 802 3326
rect 1830 3324 1836 3325
rect 3532 3324 3534 3329
rect 399 3323 400 3324
rect 394 3322 400 3323
rect 110 3319 116 3320
rect 1830 3320 1831 3324
rect 1835 3320 1836 3324
rect 3530 3323 3536 3324
rect 1830 3319 1836 3320
rect 1870 3320 1876 3321
rect 1870 3316 1871 3320
rect 1875 3316 1876 3320
rect 3530 3319 3531 3323
rect 3535 3319 3536 3323
rect 3530 3318 3536 3319
rect 3590 3320 3596 3321
rect 1870 3315 1876 3316
rect 3590 3316 3591 3320
rect 3595 3316 3596 3320
rect 3590 3315 3596 3316
rect 214 3306 220 3307
rect 214 3302 215 3306
rect 219 3302 220 3306
rect 214 3301 220 3302
rect 342 3306 348 3307
rect 342 3302 343 3306
rect 347 3302 348 3306
rect 342 3301 348 3302
rect 478 3306 484 3307
rect 478 3302 479 3306
rect 483 3302 484 3306
rect 478 3301 484 3302
rect 630 3306 636 3307
rect 630 3302 631 3306
rect 635 3302 636 3306
rect 630 3301 636 3302
rect 790 3306 796 3307
rect 790 3302 791 3306
rect 795 3302 796 3306
rect 790 3301 796 3302
rect 950 3306 956 3307
rect 950 3302 951 3306
rect 955 3302 956 3306
rect 950 3301 956 3302
rect 1110 3306 1116 3307
rect 1110 3302 1111 3306
rect 1115 3302 1116 3306
rect 1110 3301 1116 3302
rect 1270 3306 1276 3307
rect 1270 3302 1271 3306
rect 1275 3302 1276 3306
rect 1270 3301 1276 3302
rect 1430 3306 1436 3307
rect 1430 3302 1431 3306
rect 1435 3302 1436 3306
rect 1430 3301 1436 3302
rect 1590 3306 1596 3307
rect 1590 3302 1591 3306
rect 1595 3302 1596 3306
rect 1590 3301 1596 3302
rect 1750 3306 1756 3307
rect 1750 3302 1751 3306
rect 1755 3302 1756 3306
rect 1750 3301 1756 3302
rect 2134 3302 2140 3303
rect 2134 3298 2135 3302
rect 2139 3298 2140 3302
rect 2134 3297 2140 3298
rect 2230 3302 2236 3303
rect 2230 3298 2231 3302
rect 2235 3298 2236 3302
rect 2230 3297 2236 3298
rect 2342 3302 2348 3303
rect 2342 3298 2343 3302
rect 2347 3298 2348 3302
rect 2342 3297 2348 3298
rect 2462 3302 2468 3303
rect 2462 3298 2463 3302
rect 2467 3298 2468 3302
rect 2462 3297 2468 3298
rect 2590 3302 2596 3303
rect 2590 3298 2591 3302
rect 2595 3298 2596 3302
rect 2590 3297 2596 3298
rect 2726 3302 2732 3303
rect 2726 3298 2727 3302
rect 2731 3298 2732 3302
rect 2726 3297 2732 3298
rect 2870 3302 2876 3303
rect 2870 3298 2871 3302
rect 2875 3298 2876 3302
rect 2870 3297 2876 3298
rect 3014 3302 3020 3303
rect 3014 3298 3015 3302
rect 3019 3298 3020 3302
rect 3014 3297 3020 3298
rect 3166 3302 3172 3303
rect 3166 3298 3167 3302
rect 3171 3298 3172 3302
rect 3166 3297 3172 3298
rect 3318 3302 3324 3303
rect 3318 3298 3319 3302
rect 3323 3298 3324 3302
rect 3318 3297 3324 3298
rect 3478 3302 3484 3303
rect 3478 3298 3479 3302
rect 3483 3298 3484 3302
rect 3478 3297 3484 3298
rect 207 3295 213 3296
rect 207 3291 208 3295
rect 212 3294 213 3295
rect 222 3295 228 3296
rect 222 3294 223 3295
rect 212 3292 223 3294
rect 212 3291 213 3292
rect 207 3290 213 3291
rect 222 3291 223 3292
rect 227 3291 228 3295
rect 222 3290 228 3291
rect 278 3295 284 3296
rect 278 3291 279 3295
rect 283 3294 284 3295
rect 335 3295 341 3296
rect 335 3294 336 3295
rect 283 3292 336 3294
rect 283 3291 284 3292
rect 278 3290 284 3291
rect 335 3291 336 3292
rect 340 3291 341 3295
rect 335 3290 341 3291
rect 410 3295 416 3296
rect 410 3291 411 3295
rect 415 3294 416 3295
rect 471 3295 477 3296
rect 471 3294 472 3295
rect 415 3292 472 3294
rect 415 3291 416 3292
rect 410 3290 416 3291
rect 471 3291 472 3292
rect 476 3291 477 3295
rect 471 3290 477 3291
rect 551 3295 557 3296
rect 551 3291 552 3295
rect 556 3294 557 3295
rect 623 3295 629 3296
rect 623 3294 624 3295
rect 556 3292 624 3294
rect 556 3291 557 3292
rect 551 3290 557 3291
rect 623 3291 624 3292
rect 628 3291 629 3295
rect 623 3290 629 3291
rect 706 3295 712 3296
rect 706 3291 707 3295
rect 711 3294 712 3295
rect 783 3295 789 3296
rect 783 3294 784 3295
rect 711 3292 784 3294
rect 711 3291 712 3292
rect 706 3290 712 3291
rect 783 3291 784 3292
rect 788 3291 789 3295
rect 783 3290 789 3291
rect 943 3295 949 3296
rect 943 3291 944 3295
rect 948 3294 949 3295
rect 1010 3295 1016 3296
rect 1010 3294 1011 3295
rect 948 3292 1011 3294
rect 948 3291 949 3292
rect 943 3290 949 3291
rect 1010 3291 1011 3292
rect 1015 3291 1016 3295
rect 1010 3290 1016 3291
rect 1103 3295 1109 3296
rect 1103 3291 1104 3295
rect 1108 3294 1109 3295
rect 1170 3295 1176 3296
rect 1170 3294 1171 3295
rect 1108 3292 1171 3294
rect 1108 3291 1109 3292
rect 1103 3290 1109 3291
rect 1170 3291 1171 3292
rect 1175 3291 1176 3295
rect 1170 3290 1176 3291
rect 1262 3295 1269 3296
rect 1262 3291 1263 3295
rect 1268 3291 1269 3295
rect 1262 3290 1269 3291
rect 1423 3295 1429 3296
rect 1423 3291 1424 3295
rect 1428 3294 1429 3295
rect 1527 3295 1533 3296
rect 1527 3294 1528 3295
rect 1428 3292 1528 3294
rect 1428 3291 1429 3292
rect 1423 3290 1429 3291
rect 1527 3291 1528 3292
rect 1532 3291 1533 3295
rect 1527 3290 1533 3291
rect 1583 3295 1589 3296
rect 1583 3291 1584 3295
rect 1588 3294 1589 3295
rect 1650 3295 1656 3296
rect 1650 3294 1651 3295
rect 1588 3292 1651 3294
rect 1588 3291 1589 3292
rect 1583 3290 1589 3291
rect 1650 3291 1651 3292
rect 1655 3291 1656 3295
rect 1650 3290 1656 3291
rect 1734 3295 1740 3296
rect 1734 3291 1735 3295
rect 1739 3294 1740 3295
rect 1743 3295 1749 3296
rect 1743 3294 1744 3295
rect 1739 3292 1744 3294
rect 1739 3291 1740 3292
rect 1734 3290 1740 3291
rect 1743 3291 1744 3292
rect 1748 3291 1749 3295
rect 1743 3290 1749 3291
rect 2127 3291 2133 3292
rect 2127 3287 2128 3291
rect 2132 3290 2133 3291
rect 2142 3291 2148 3292
rect 2142 3290 2143 3291
rect 2132 3288 2143 3290
rect 2132 3287 2133 3288
rect 2127 3286 2133 3287
rect 2142 3287 2143 3288
rect 2147 3287 2148 3291
rect 2142 3286 2148 3287
rect 2194 3291 2200 3292
rect 2194 3287 2195 3291
rect 2199 3290 2200 3291
rect 2223 3291 2229 3292
rect 2223 3290 2224 3291
rect 2199 3288 2224 3290
rect 2199 3287 2200 3288
rect 2194 3286 2200 3287
rect 2223 3287 2224 3288
rect 2228 3287 2229 3291
rect 2223 3286 2229 3287
rect 2290 3291 2296 3292
rect 2290 3287 2291 3291
rect 2295 3290 2296 3291
rect 2335 3291 2341 3292
rect 2335 3290 2336 3291
rect 2295 3288 2336 3290
rect 2295 3287 2296 3288
rect 2290 3286 2296 3287
rect 2335 3287 2336 3288
rect 2340 3287 2341 3291
rect 2335 3286 2341 3287
rect 2402 3291 2408 3292
rect 2402 3287 2403 3291
rect 2407 3290 2408 3291
rect 2455 3291 2461 3292
rect 2455 3290 2456 3291
rect 2407 3288 2456 3290
rect 2407 3287 2408 3288
rect 2402 3286 2408 3287
rect 2455 3287 2456 3288
rect 2460 3287 2461 3291
rect 2455 3286 2461 3287
rect 2574 3291 2580 3292
rect 2574 3287 2575 3291
rect 2579 3290 2580 3291
rect 2583 3291 2589 3292
rect 2583 3290 2584 3291
rect 2579 3288 2584 3290
rect 2579 3287 2580 3288
rect 2574 3286 2580 3287
rect 2583 3287 2584 3288
rect 2588 3287 2589 3291
rect 2583 3286 2589 3287
rect 2650 3291 2656 3292
rect 2650 3287 2651 3291
rect 2655 3290 2656 3291
rect 2719 3291 2725 3292
rect 2719 3290 2720 3291
rect 2655 3288 2720 3290
rect 2655 3287 2656 3288
rect 2650 3286 2656 3287
rect 2719 3287 2720 3288
rect 2724 3287 2725 3291
rect 2719 3286 2725 3287
rect 2798 3291 2804 3292
rect 2798 3287 2799 3291
rect 2803 3290 2804 3291
rect 2863 3291 2869 3292
rect 2863 3290 2864 3291
rect 2803 3288 2864 3290
rect 2803 3287 2804 3288
rect 2798 3286 2804 3287
rect 2863 3287 2864 3288
rect 2868 3287 2869 3291
rect 2863 3286 2869 3287
rect 3006 3291 3013 3292
rect 3006 3287 3007 3291
rect 3012 3287 3013 3291
rect 3006 3286 3013 3287
rect 3079 3291 3085 3292
rect 3079 3287 3080 3291
rect 3084 3290 3085 3291
rect 3159 3291 3165 3292
rect 3159 3290 3160 3291
rect 3084 3288 3160 3290
rect 3084 3287 3085 3288
rect 3079 3286 3085 3287
rect 3159 3287 3160 3288
rect 3164 3287 3165 3291
rect 3159 3286 3165 3287
rect 3302 3291 3308 3292
rect 3302 3287 3303 3291
rect 3307 3290 3308 3291
rect 3311 3291 3317 3292
rect 3311 3290 3312 3291
rect 3307 3288 3312 3290
rect 3307 3287 3308 3288
rect 3302 3286 3308 3287
rect 3311 3287 3312 3288
rect 3316 3287 3317 3291
rect 3311 3286 3317 3287
rect 3394 3291 3400 3292
rect 3394 3287 3395 3291
rect 3399 3290 3400 3291
rect 3471 3291 3477 3292
rect 3471 3290 3472 3291
rect 3399 3288 3472 3290
rect 3399 3287 3400 3288
rect 3394 3286 3400 3287
rect 3471 3287 3472 3288
rect 3476 3287 3477 3291
rect 3471 3286 3477 3287
rect 343 3279 349 3280
rect 343 3275 344 3279
rect 348 3278 349 3279
rect 394 3279 400 3280
rect 394 3278 395 3279
rect 348 3276 395 3278
rect 348 3275 349 3276
rect 343 3274 349 3275
rect 394 3275 395 3276
rect 399 3275 400 3279
rect 394 3274 400 3275
rect 402 3279 408 3280
rect 402 3275 403 3279
rect 407 3278 408 3279
rect 447 3279 453 3280
rect 447 3278 448 3279
rect 407 3276 448 3278
rect 407 3275 408 3276
rect 402 3274 408 3275
rect 447 3275 448 3276
rect 452 3275 453 3279
rect 447 3274 453 3275
rect 506 3279 512 3280
rect 506 3275 507 3279
rect 511 3278 512 3279
rect 567 3279 573 3280
rect 567 3278 568 3279
rect 511 3276 568 3278
rect 511 3275 512 3276
rect 506 3274 512 3275
rect 567 3275 568 3276
rect 572 3275 573 3279
rect 567 3274 573 3275
rect 655 3279 661 3280
rect 655 3275 656 3279
rect 660 3278 661 3279
rect 695 3279 701 3280
rect 695 3278 696 3279
rect 660 3276 696 3278
rect 660 3275 661 3276
rect 655 3274 661 3275
rect 695 3275 696 3276
rect 700 3275 701 3279
rect 695 3274 701 3275
rect 754 3279 760 3280
rect 754 3275 755 3279
rect 759 3278 760 3279
rect 831 3279 837 3280
rect 831 3278 832 3279
rect 759 3276 832 3278
rect 759 3275 760 3276
rect 754 3274 760 3275
rect 831 3275 832 3276
rect 836 3275 837 3279
rect 831 3274 837 3275
rect 975 3279 981 3280
rect 975 3275 976 3279
rect 980 3278 981 3279
rect 990 3279 996 3280
rect 990 3278 991 3279
rect 980 3276 991 3278
rect 980 3275 981 3276
rect 975 3274 981 3275
rect 990 3275 991 3276
rect 995 3275 996 3279
rect 990 3274 996 3275
rect 1034 3279 1040 3280
rect 1034 3275 1035 3279
rect 1039 3278 1040 3279
rect 1111 3279 1117 3280
rect 1111 3278 1112 3279
rect 1039 3276 1112 3278
rect 1039 3275 1040 3276
rect 1034 3274 1040 3275
rect 1111 3275 1112 3276
rect 1116 3275 1117 3279
rect 1111 3274 1117 3275
rect 1170 3279 1176 3280
rect 1170 3275 1171 3279
rect 1175 3278 1176 3279
rect 1247 3279 1253 3280
rect 1247 3278 1248 3279
rect 1175 3276 1248 3278
rect 1175 3275 1176 3276
rect 1170 3274 1176 3275
rect 1247 3275 1248 3276
rect 1252 3275 1253 3279
rect 1247 3274 1253 3275
rect 1375 3279 1381 3280
rect 1375 3275 1376 3279
rect 1380 3278 1381 3279
rect 1383 3279 1389 3280
rect 1383 3278 1384 3279
rect 1380 3276 1384 3278
rect 1380 3275 1381 3276
rect 1375 3274 1381 3275
rect 1383 3275 1384 3276
rect 1388 3275 1389 3279
rect 1383 3274 1389 3275
rect 1479 3279 1485 3280
rect 1479 3275 1480 3279
rect 1484 3278 1485 3279
rect 1503 3279 1509 3280
rect 1503 3278 1504 3279
rect 1484 3276 1504 3278
rect 1484 3275 1485 3276
rect 1479 3274 1485 3275
rect 1503 3275 1504 3276
rect 1508 3275 1509 3279
rect 1503 3274 1509 3275
rect 1562 3279 1568 3280
rect 1562 3275 1563 3279
rect 1567 3278 1568 3279
rect 1631 3279 1637 3280
rect 1631 3278 1632 3279
rect 1567 3276 1632 3278
rect 1567 3275 1568 3276
rect 1562 3274 1568 3275
rect 1631 3275 1632 3276
rect 1636 3275 1637 3279
rect 1631 3274 1637 3275
rect 1690 3279 1696 3280
rect 1690 3275 1691 3279
rect 1695 3278 1696 3279
rect 1743 3279 1749 3280
rect 1743 3278 1744 3279
rect 1695 3276 1744 3278
rect 1695 3275 1696 3276
rect 1690 3274 1696 3275
rect 1743 3275 1744 3276
rect 1748 3275 1749 3279
rect 1743 3274 1749 3275
rect 2422 3275 2428 3276
rect 2422 3274 2423 3275
rect 2212 3272 2423 3274
rect 350 3270 356 3271
rect 350 3266 351 3270
rect 355 3266 356 3270
rect 350 3265 356 3266
rect 454 3270 460 3271
rect 454 3266 455 3270
rect 459 3266 460 3270
rect 454 3265 460 3266
rect 574 3270 580 3271
rect 574 3266 575 3270
rect 579 3266 580 3270
rect 574 3265 580 3266
rect 702 3270 708 3271
rect 702 3266 703 3270
rect 707 3266 708 3270
rect 702 3265 708 3266
rect 838 3270 844 3271
rect 838 3266 839 3270
rect 843 3266 844 3270
rect 838 3265 844 3266
rect 982 3270 988 3271
rect 982 3266 983 3270
rect 987 3266 988 3270
rect 982 3265 988 3266
rect 1118 3270 1124 3271
rect 1118 3266 1119 3270
rect 1123 3266 1124 3270
rect 1118 3265 1124 3266
rect 1254 3270 1260 3271
rect 1254 3266 1255 3270
rect 1259 3266 1260 3270
rect 1254 3265 1260 3266
rect 1382 3270 1388 3271
rect 1382 3266 1383 3270
rect 1387 3266 1388 3270
rect 1382 3265 1388 3266
rect 1510 3270 1516 3271
rect 1510 3266 1511 3270
rect 1515 3266 1516 3270
rect 1510 3265 1516 3266
rect 1638 3270 1644 3271
rect 1638 3266 1639 3270
rect 1643 3266 1644 3270
rect 1638 3265 1644 3266
rect 1750 3270 1756 3271
rect 1750 3266 1751 3270
rect 1755 3266 1756 3270
rect 1750 3265 1756 3266
rect 2127 3267 2133 3268
rect 2127 3263 2128 3267
rect 2132 3266 2133 3267
rect 2212 3266 2214 3272
rect 2422 3271 2423 3272
rect 2427 3271 2428 3275
rect 2422 3270 2428 3271
rect 2132 3264 2214 3266
rect 2254 3267 2260 3268
rect 2132 3263 2133 3264
rect 2127 3262 2133 3263
rect 2254 3263 2255 3267
rect 2259 3266 2260 3267
rect 2271 3267 2277 3268
rect 2271 3266 2272 3267
rect 2259 3264 2272 3266
rect 2259 3263 2260 3264
rect 2254 3262 2260 3263
rect 2271 3263 2272 3264
rect 2276 3263 2277 3267
rect 2271 3262 2277 3263
rect 2330 3267 2336 3268
rect 2330 3263 2331 3267
rect 2335 3266 2336 3267
rect 2407 3267 2413 3268
rect 2407 3266 2408 3267
rect 2335 3264 2408 3266
rect 2335 3263 2336 3264
rect 2330 3262 2336 3263
rect 2407 3263 2408 3264
rect 2412 3263 2413 3267
rect 2407 3262 2413 3263
rect 2543 3267 2549 3268
rect 2543 3263 2544 3267
rect 2548 3266 2549 3267
rect 2610 3267 2616 3268
rect 2610 3266 2611 3267
rect 2548 3264 2611 3266
rect 2548 3263 2549 3264
rect 2543 3262 2549 3263
rect 2610 3263 2611 3264
rect 2615 3263 2616 3267
rect 2610 3262 2616 3263
rect 2679 3267 2685 3268
rect 2679 3263 2680 3267
rect 2684 3266 2685 3267
rect 2746 3267 2752 3268
rect 2746 3266 2747 3267
rect 2684 3264 2747 3266
rect 2684 3263 2685 3264
rect 2679 3262 2685 3263
rect 2746 3263 2747 3264
rect 2751 3263 2752 3267
rect 2746 3262 2752 3263
rect 2815 3267 2821 3268
rect 2815 3263 2816 3267
rect 2820 3266 2821 3267
rect 2823 3267 2829 3268
rect 2823 3266 2824 3267
rect 2820 3264 2824 3266
rect 2820 3263 2821 3264
rect 2815 3262 2821 3263
rect 2823 3263 2824 3264
rect 2828 3263 2829 3267
rect 2823 3262 2829 3263
rect 2951 3267 2957 3268
rect 2951 3263 2952 3267
rect 2956 3266 2957 3267
rect 3022 3267 3028 3268
rect 3022 3266 3023 3267
rect 2956 3264 3023 3266
rect 2956 3263 2957 3264
rect 2951 3262 2957 3263
rect 3022 3263 3023 3264
rect 3027 3263 3028 3267
rect 3022 3262 3028 3263
rect 3087 3267 3093 3268
rect 3087 3263 3088 3267
rect 3092 3266 3093 3267
rect 3186 3267 3192 3268
rect 3186 3266 3187 3267
rect 3092 3264 3187 3266
rect 3092 3263 3093 3264
rect 3087 3262 3093 3263
rect 3186 3263 3187 3264
rect 3191 3263 3192 3267
rect 3186 3262 3192 3263
rect 3223 3267 3229 3268
rect 3223 3263 3224 3267
rect 3228 3266 3229 3267
rect 3266 3267 3272 3268
rect 3266 3266 3267 3267
rect 3228 3264 3267 3266
rect 3228 3263 3229 3264
rect 3223 3262 3229 3263
rect 3266 3263 3267 3264
rect 3271 3263 3272 3267
rect 3266 3262 3272 3263
rect 3367 3267 3373 3268
rect 3367 3263 3368 3267
rect 3372 3266 3373 3267
rect 3434 3267 3440 3268
rect 3434 3266 3435 3267
rect 3372 3264 3435 3266
rect 3372 3263 3373 3264
rect 3367 3262 3373 3263
rect 3434 3263 3435 3264
rect 3439 3263 3440 3267
rect 3434 3262 3440 3263
rect 3503 3267 3509 3268
rect 3503 3263 3504 3267
rect 3508 3266 3509 3267
rect 3530 3267 3536 3268
rect 3530 3266 3531 3267
rect 3508 3264 3531 3266
rect 3508 3263 3509 3264
rect 3503 3262 3509 3263
rect 3530 3263 3531 3264
rect 3535 3263 3536 3267
rect 3530 3262 3536 3263
rect 2134 3258 2140 3259
rect 2134 3254 2135 3258
rect 2139 3254 2140 3258
rect 2134 3253 2140 3254
rect 2278 3258 2284 3259
rect 2278 3254 2279 3258
rect 2283 3254 2284 3258
rect 2278 3253 2284 3254
rect 2414 3258 2420 3259
rect 2414 3254 2415 3258
rect 2419 3254 2420 3258
rect 2414 3253 2420 3254
rect 2550 3258 2556 3259
rect 2550 3254 2551 3258
rect 2555 3254 2556 3258
rect 2550 3253 2556 3254
rect 2686 3258 2692 3259
rect 2686 3254 2687 3258
rect 2691 3254 2692 3258
rect 2686 3253 2692 3254
rect 2822 3258 2828 3259
rect 2822 3254 2823 3258
rect 2827 3254 2828 3258
rect 2822 3253 2828 3254
rect 2958 3258 2964 3259
rect 2958 3254 2959 3258
rect 2963 3254 2964 3258
rect 2958 3253 2964 3254
rect 3094 3258 3100 3259
rect 3094 3254 3095 3258
rect 3099 3254 3100 3258
rect 3094 3253 3100 3254
rect 3230 3258 3236 3259
rect 3230 3254 3231 3258
rect 3235 3254 3236 3258
rect 3230 3253 3236 3254
rect 3374 3258 3380 3259
rect 3374 3254 3375 3258
rect 3379 3254 3380 3258
rect 3374 3253 3380 3254
rect 3510 3258 3516 3259
rect 3510 3254 3511 3258
rect 3515 3254 3516 3258
rect 3510 3253 3516 3254
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 110 3247 116 3248
rect 1830 3252 1836 3253
rect 1830 3248 1831 3252
rect 1835 3248 1836 3252
rect 1830 3247 1836 3248
rect 402 3243 408 3244
rect 402 3239 403 3243
rect 407 3239 408 3243
rect 402 3238 408 3239
rect 506 3243 512 3244
rect 506 3239 507 3243
rect 511 3239 512 3243
rect 655 3243 661 3244
rect 655 3242 656 3243
rect 629 3240 656 3242
rect 506 3238 512 3239
rect 655 3239 656 3240
rect 660 3239 661 3243
rect 655 3238 661 3239
rect 754 3243 760 3244
rect 754 3239 755 3243
rect 759 3239 760 3243
rect 754 3238 760 3239
rect 1034 3243 1040 3244
rect 1034 3239 1035 3243
rect 1039 3239 1040 3243
rect 1034 3238 1040 3239
rect 1170 3243 1176 3244
rect 1170 3239 1171 3243
rect 1175 3239 1176 3243
rect 1170 3238 1176 3239
rect 1262 3243 1268 3244
rect 1262 3239 1263 3243
rect 1267 3239 1268 3243
rect 1479 3243 1485 3244
rect 1479 3242 1480 3243
rect 1437 3240 1480 3242
rect 1262 3238 1268 3239
rect 1479 3239 1480 3240
rect 1484 3239 1485 3243
rect 1479 3238 1485 3239
rect 1562 3243 1568 3244
rect 1562 3239 1563 3243
rect 1567 3239 1568 3243
rect 1562 3238 1568 3239
rect 1690 3243 1696 3244
rect 1690 3239 1691 3243
rect 1695 3239 1696 3243
rect 1690 3238 1696 3239
rect 1870 3240 1876 3241
rect 1870 3236 1871 3240
rect 1875 3236 1876 3240
rect 110 3235 116 3236
rect 110 3231 111 3235
rect 115 3231 116 3235
rect 1830 3235 1836 3236
rect 1870 3235 1876 3236
rect 3590 3240 3596 3241
rect 3590 3236 3591 3240
rect 3595 3236 3596 3240
rect 3590 3235 3596 3236
rect 110 3230 116 3231
rect 342 3232 348 3233
rect 342 3228 343 3232
rect 347 3228 348 3232
rect 342 3227 348 3228
rect 446 3232 452 3233
rect 446 3228 447 3232
rect 451 3228 452 3232
rect 446 3227 452 3228
rect 566 3232 572 3233
rect 566 3228 567 3232
rect 571 3228 572 3232
rect 566 3227 572 3228
rect 694 3232 700 3233
rect 694 3228 695 3232
rect 699 3228 700 3232
rect 694 3227 700 3228
rect 830 3232 836 3233
rect 830 3228 831 3232
rect 835 3228 836 3232
rect 830 3227 836 3228
rect 974 3232 980 3233
rect 974 3228 975 3232
rect 979 3228 980 3232
rect 974 3227 980 3228
rect 1110 3232 1116 3233
rect 1110 3228 1111 3232
rect 1115 3228 1116 3232
rect 1110 3227 1116 3228
rect 1246 3232 1252 3233
rect 1246 3228 1247 3232
rect 1251 3228 1252 3232
rect 1246 3227 1252 3228
rect 1374 3232 1380 3233
rect 1374 3228 1375 3232
rect 1379 3228 1380 3232
rect 1374 3227 1380 3228
rect 1502 3232 1508 3233
rect 1502 3228 1503 3232
rect 1507 3228 1508 3232
rect 1502 3227 1508 3228
rect 1630 3232 1636 3233
rect 1630 3228 1631 3232
rect 1635 3228 1636 3232
rect 1630 3227 1636 3228
rect 1742 3232 1748 3233
rect 1742 3228 1743 3232
rect 1747 3228 1748 3232
rect 1830 3231 1831 3235
rect 1835 3231 1836 3235
rect 1830 3230 1836 3231
rect 2142 3231 2148 3232
rect 1742 3227 1748 3228
rect 2142 3227 2143 3231
rect 2147 3227 2148 3231
rect 2142 3226 2148 3227
rect 2330 3231 2336 3232
rect 2330 3227 2331 3231
rect 2335 3227 2336 3231
rect 2330 3226 2336 3227
rect 2422 3231 2428 3232
rect 2422 3227 2423 3231
rect 2427 3227 2428 3231
rect 2422 3226 2428 3227
rect 2610 3231 2616 3232
rect 2610 3227 2611 3231
rect 2615 3230 2616 3231
rect 2746 3231 2752 3232
rect 2615 3228 2697 3230
rect 2615 3227 2616 3228
rect 2610 3226 2616 3227
rect 2746 3227 2747 3231
rect 2751 3230 2752 3231
rect 3006 3231 3012 3232
rect 2751 3228 2833 3230
rect 2751 3227 2752 3228
rect 2746 3226 2752 3227
rect 3006 3227 3007 3231
rect 3011 3227 3012 3231
rect 3006 3226 3012 3227
rect 3022 3231 3028 3232
rect 3022 3227 3023 3231
rect 3027 3230 3028 3231
rect 3186 3231 3192 3232
rect 3027 3228 3105 3230
rect 3027 3227 3028 3228
rect 3022 3226 3028 3227
rect 3186 3227 3187 3231
rect 3191 3230 3192 3231
rect 3426 3231 3432 3232
rect 3191 3228 3241 3230
rect 3191 3227 3192 3228
rect 3186 3226 3192 3227
rect 3426 3227 3427 3231
rect 3431 3227 3432 3231
rect 3426 3226 3432 3227
rect 3434 3231 3440 3232
rect 3434 3227 3435 3231
rect 3439 3230 3440 3231
rect 3439 3228 3521 3230
rect 3439 3227 3440 3228
rect 3434 3226 3440 3227
rect 1870 3223 1876 3224
rect 1870 3219 1871 3223
rect 1875 3219 1876 3223
rect 3590 3223 3596 3224
rect 1870 3218 1876 3219
rect 2126 3220 2132 3221
rect 2126 3216 2127 3220
rect 2131 3216 2132 3220
rect 502 3215 508 3216
rect 502 3211 503 3215
rect 507 3214 508 3215
rect 847 3215 853 3216
rect 847 3214 848 3215
rect 507 3212 848 3214
rect 507 3211 508 3212
rect 502 3210 508 3211
rect 847 3211 848 3212
rect 852 3211 853 3215
rect 847 3210 853 3211
rect 1758 3215 1765 3216
rect 2126 3215 2132 3216
rect 2270 3220 2276 3221
rect 2270 3216 2271 3220
rect 2275 3216 2276 3220
rect 2270 3215 2276 3216
rect 2406 3220 2412 3221
rect 2406 3216 2407 3220
rect 2411 3216 2412 3220
rect 2406 3215 2412 3216
rect 2542 3220 2548 3221
rect 2542 3216 2543 3220
rect 2547 3216 2548 3220
rect 2542 3215 2548 3216
rect 2678 3220 2684 3221
rect 2678 3216 2679 3220
rect 2683 3216 2684 3220
rect 2678 3215 2684 3216
rect 2814 3220 2820 3221
rect 2814 3216 2815 3220
rect 2819 3216 2820 3220
rect 2814 3215 2820 3216
rect 2950 3220 2956 3221
rect 2950 3216 2951 3220
rect 2955 3216 2956 3220
rect 2950 3215 2956 3216
rect 3086 3220 3092 3221
rect 3086 3216 3087 3220
rect 3091 3216 3092 3220
rect 3086 3215 3092 3216
rect 3222 3220 3228 3221
rect 3222 3216 3223 3220
rect 3227 3216 3228 3220
rect 3222 3215 3228 3216
rect 3366 3220 3372 3221
rect 3366 3216 3367 3220
rect 3371 3216 3372 3220
rect 3366 3215 3372 3216
rect 3502 3220 3508 3221
rect 3502 3216 3503 3220
rect 3507 3216 3508 3220
rect 3590 3219 3591 3223
rect 3595 3219 3596 3223
rect 3590 3218 3596 3219
rect 3502 3215 3508 3216
rect 1758 3211 1759 3215
rect 1764 3211 1765 3215
rect 1758 3210 1765 3211
rect 2550 3203 2556 3204
rect 2550 3199 2551 3203
rect 2555 3202 2556 3203
rect 2559 3203 2565 3204
rect 2559 3202 2560 3203
rect 2555 3200 2560 3202
rect 2555 3199 2556 3200
rect 2550 3198 2556 3199
rect 2559 3199 2560 3200
rect 2564 3199 2565 3203
rect 2559 3198 2565 3199
rect 486 3188 492 3189
rect 110 3185 116 3186
rect 110 3181 111 3185
rect 115 3181 116 3185
rect 486 3184 487 3188
rect 491 3184 492 3188
rect 486 3183 492 3184
rect 574 3188 580 3189
rect 574 3184 575 3188
rect 579 3184 580 3188
rect 574 3183 580 3184
rect 662 3188 668 3189
rect 662 3184 663 3188
rect 667 3184 668 3188
rect 662 3183 668 3184
rect 766 3188 772 3189
rect 766 3184 767 3188
rect 771 3184 772 3188
rect 766 3183 772 3184
rect 886 3188 892 3189
rect 886 3184 887 3188
rect 891 3184 892 3188
rect 886 3183 892 3184
rect 1022 3188 1028 3189
rect 1022 3184 1023 3188
rect 1027 3184 1028 3188
rect 1022 3183 1028 3184
rect 1190 3188 1196 3189
rect 1190 3184 1191 3188
rect 1195 3184 1196 3188
rect 1190 3183 1196 3184
rect 1374 3188 1380 3189
rect 1374 3184 1375 3188
rect 1379 3184 1380 3188
rect 1374 3183 1380 3184
rect 1566 3188 1572 3189
rect 1566 3184 1567 3188
rect 1571 3184 1572 3188
rect 1566 3183 1572 3184
rect 1742 3188 1748 3189
rect 1742 3184 1743 3188
rect 1747 3184 1748 3188
rect 1742 3183 1748 3184
rect 1830 3185 1836 3186
rect 110 3180 116 3181
rect 1830 3181 1831 3185
rect 1835 3181 1836 3185
rect 1830 3180 1836 3181
rect 554 3179 560 3180
rect 554 3178 555 3179
rect 549 3176 555 3178
rect 554 3175 555 3176
rect 559 3175 560 3179
rect 642 3179 648 3180
rect 642 3178 643 3179
rect 637 3176 643 3178
rect 554 3174 560 3175
rect 642 3175 643 3176
rect 647 3175 648 3179
rect 730 3179 736 3180
rect 730 3178 731 3179
rect 725 3176 731 3178
rect 642 3174 648 3175
rect 730 3175 731 3176
rect 735 3175 736 3179
rect 834 3179 840 3180
rect 834 3178 835 3179
rect 829 3176 835 3178
rect 730 3174 736 3175
rect 834 3175 835 3176
rect 839 3175 840 3179
rect 834 3174 840 3175
rect 842 3179 848 3180
rect 842 3175 843 3179
rect 847 3178 848 3179
rect 990 3179 996 3180
rect 847 3176 905 3178
rect 847 3175 848 3176
rect 842 3174 848 3175
rect 990 3175 991 3179
rect 995 3178 996 3179
rect 1106 3179 1112 3180
rect 995 3176 1041 3178
rect 995 3175 996 3176
rect 990 3174 996 3175
rect 1106 3175 1107 3179
rect 1111 3178 1112 3179
rect 1478 3179 1484 3180
rect 1478 3178 1479 3179
rect 1111 3176 1209 3178
rect 1437 3176 1479 3178
rect 1111 3175 1112 3176
rect 1106 3174 1112 3175
rect 1478 3175 1479 3176
rect 1483 3175 1484 3179
rect 1478 3174 1484 3175
rect 1486 3179 1492 3180
rect 1486 3175 1487 3179
rect 1491 3178 1492 3179
rect 1818 3179 1824 3180
rect 1818 3178 1819 3179
rect 1491 3176 1585 3178
rect 1805 3176 1819 3178
rect 1491 3175 1492 3176
rect 1486 3174 1492 3175
rect 1818 3175 1819 3176
rect 1823 3175 1824 3179
rect 1818 3174 1824 3175
rect 1894 3172 1900 3173
rect 1870 3169 1876 3170
rect 110 3168 116 3169
rect 110 3164 111 3168
rect 115 3164 116 3168
rect 110 3163 116 3164
rect 1830 3168 1836 3169
rect 1830 3164 1831 3168
rect 1835 3164 1836 3168
rect 1870 3165 1871 3169
rect 1875 3165 1876 3169
rect 1894 3168 1895 3172
rect 1899 3168 1900 3172
rect 1894 3167 1900 3168
rect 1990 3172 1996 3173
rect 1990 3168 1991 3172
rect 1995 3168 1996 3172
rect 1990 3167 1996 3168
rect 2118 3172 2124 3173
rect 2118 3168 2119 3172
rect 2123 3168 2124 3172
rect 2118 3167 2124 3168
rect 2246 3172 2252 3173
rect 2246 3168 2247 3172
rect 2251 3168 2252 3172
rect 2246 3167 2252 3168
rect 2382 3172 2388 3173
rect 2382 3168 2383 3172
rect 2387 3168 2388 3172
rect 2382 3167 2388 3168
rect 2510 3172 2516 3173
rect 2510 3168 2511 3172
rect 2515 3168 2516 3172
rect 2510 3167 2516 3168
rect 2638 3172 2644 3173
rect 2638 3168 2639 3172
rect 2643 3168 2644 3172
rect 2638 3167 2644 3168
rect 2766 3172 2772 3173
rect 2766 3168 2767 3172
rect 2771 3168 2772 3172
rect 2766 3167 2772 3168
rect 2894 3172 2900 3173
rect 2894 3168 2895 3172
rect 2899 3168 2900 3172
rect 2894 3167 2900 3168
rect 3030 3172 3036 3173
rect 3030 3168 3031 3172
rect 3035 3168 3036 3172
rect 3030 3167 3036 3168
rect 3174 3172 3180 3173
rect 3174 3168 3175 3172
rect 3179 3168 3180 3172
rect 3174 3167 3180 3168
rect 3326 3172 3332 3173
rect 3326 3168 3327 3172
rect 3331 3168 3332 3172
rect 3326 3167 3332 3168
rect 3486 3172 3492 3173
rect 3486 3168 3487 3172
rect 3491 3168 3492 3172
rect 3486 3167 3492 3168
rect 3590 3169 3596 3170
rect 1870 3164 1876 3165
rect 3590 3165 3591 3169
rect 3595 3165 3596 3169
rect 3590 3164 3596 3165
rect 1830 3163 1836 3164
rect 1962 3163 1968 3164
rect 1962 3162 1963 3163
rect 1957 3160 1963 3162
rect 1962 3159 1963 3160
rect 1967 3159 1968 3163
rect 2062 3163 2068 3164
rect 2062 3162 2063 3163
rect 2053 3160 2063 3162
rect 1962 3158 1968 3159
rect 2062 3159 2063 3160
rect 2067 3159 2068 3163
rect 2350 3163 2356 3164
rect 2062 3158 2068 3159
rect 2180 3156 2182 3161
rect 2256 3160 2265 3162
rect 2254 3159 2260 3160
rect 2178 3155 2184 3156
rect 1870 3152 1876 3153
rect 494 3150 500 3151
rect 494 3146 495 3150
rect 499 3146 500 3150
rect 494 3145 500 3146
rect 582 3150 588 3151
rect 582 3146 583 3150
rect 587 3146 588 3150
rect 582 3145 588 3146
rect 670 3150 676 3151
rect 670 3146 671 3150
rect 675 3146 676 3150
rect 670 3145 676 3146
rect 774 3150 780 3151
rect 774 3146 775 3150
rect 779 3146 780 3150
rect 774 3145 780 3146
rect 894 3150 900 3151
rect 894 3146 895 3150
rect 899 3146 900 3150
rect 894 3145 900 3146
rect 1030 3150 1036 3151
rect 1030 3146 1031 3150
rect 1035 3146 1036 3150
rect 1030 3145 1036 3146
rect 1198 3150 1204 3151
rect 1198 3146 1199 3150
rect 1203 3146 1204 3150
rect 1198 3145 1204 3146
rect 1382 3150 1388 3151
rect 1382 3146 1383 3150
rect 1387 3146 1388 3150
rect 1382 3145 1388 3146
rect 1574 3150 1580 3151
rect 1574 3146 1575 3150
rect 1579 3146 1580 3150
rect 1574 3145 1580 3146
rect 1750 3150 1756 3151
rect 1750 3146 1751 3150
rect 1755 3146 1756 3150
rect 1870 3148 1871 3152
rect 1875 3148 1876 3152
rect 2178 3151 2179 3155
rect 2183 3151 2184 3155
rect 2254 3155 2255 3159
rect 2259 3155 2260 3159
rect 2350 3159 2351 3163
rect 2355 3162 2356 3163
rect 2582 3163 2588 3164
rect 2582 3162 2583 3163
rect 2355 3160 2401 3162
rect 2573 3160 2583 3162
rect 2355 3159 2356 3160
rect 2350 3158 2356 3159
rect 2582 3159 2583 3160
rect 2587 3159 2588 3163
rect 2710 3163 2716 3164
rect 2710 3162 2711 3163
rect 2701 3160 2711 3162
rect 2582 3158 2588 3159
rect 2710 3159 2711 3160
rect 2715 3159 2716 3163
rect 2838 3163 2844 3164
rect 2838 3162 2839 3163
rect 2829 3160 2839 3162
rect 2710 3158 2716 3159
rect 2838 3159 2839 3160
rect 2843 3159 2844 3163
rect 2970 3163 2976 3164
rect 2970 3162 2971 3163
rect 2957 3160 2971 3162
rect 2838 3158 2844 3159
rect 2970 3159 2971 3160
rect 2975 3159 2976 3163
rect 3098 3163 3104 3164
rect 3098 3162 3099 3163
rect 3093 3160 3099 3162
rect 2970 3158 2976 3159
rect 3098 3159 3099 3160
rect 3103 3159 3104 3163
rect 3258 3163 3264 3164
rect 3258 3162 3259 3163
rect 3237 3160 3259 3162
rect 3098 3158 3104 3159
rect 3258 3159 3259 3160
rect 3263 3159 3264 3163
rect 3258 3158 3264 3159
rect 3266 3163 3272 3164
rect 3266 3159 3267 3163
rect 3271 3162 3272 3163
rect 3271 3160 3345 3162
rect 3271 3159 3272 3160
rect 3266 3158 3272 3159
rect 2254 3154 2260 3155
rect 3238 3155 3244 3156
rect 2178 3150 2184 3151
rect 3238 3151 3239 3155
rect 3243 3154 3244 3155
rect 3504 3154 3506 3161
rect 3243 3152 3506 3154
rect 3590 3152 3596 3153
rect 3243 3151 3244 3152
rect 3238 3150 3244 3151
rect 1870 3147 1876 3148
rect 3590 3148 3591 3152
rect 3595 3148 3596 3152
rect 3590 3147 3596 3148
rect 1750 3145 1756 3146
rect 487 3139 493 3140
rect 487 3135 488 3139
rect 492 3138 493 3139
rect 502 3139 508 3140
rect 502 3138 503 3139
rect 492 3136 503 3138
rect 492 3135 493 3136
rect 487 3134 493 3135
rect 502 3135 503 3136
rect 507 3135 508 3139
rect 502 3134 508 3135
rect 554 3139 560 3140
rect 554 3135 555 3139
rect 559 3138 560 3139
rect 575 3139 581 3140
rect 575 3138 576 3139
rect 559 3136 576 3138
rect 559 3135 560 3136
rect 554 3134 560 3135
rect 575 3135 576 3136
rect 580 3135 581 3139
rect 575 3134 581 3135
rect 642 3139 648 3140
rect 642 3135 643 3139
rect 647 3138 648 3139
rect 663 3139 669 3140
rect 663 3138 664 3139
rect 647 3136 664 3138
rect 647 3135 648 3136
rect 642 3134 648 3135
rect 663 3135 664 3136
rect 668 3135 669 3139
rect 663 3134 669 3135
rect 730 3139 736 3140
rect 730 3135 731 3139
rect 735 3138 736 3139
rect 767 3139 773 3140
rect 767 3138 768 3139
rect 735 3136 768 3138
rect 735 3135 736 3136
rect 730 3134 736 3135
rect 767 3135 768 3136
rect 772 3135 773 3139
rect 767 3134 773 3135
rect 834 3139 840 3140
rect 834 3135 835 3139
rect 839 3138 840 3139
rect 887 3139 893 3140
rect 887 3138 888 3139
rect 839 3136 888 3138
rect 839 3135 840 3136
rect 834 3134 840 3135
rect 887 3135 888 3136
rect 892 3135 893 3139
rect 887 3134 893 3135
rect 1023 3139 1029 3140
rect 1023 3135 1024 3139
rect 1028 3138 1029 3139
rect 1106 3139 1112 3140
rect 1106 3138 1107 3139
rect 1028 3136 1107 3138
rect 1028 3135 1029 3136
rect 1023 3134 1029 3135
rect 1106 3135 1107 3136
rect 1111 3135 1112 3139
rect 1106 3134 1112 3135
rect 1191 3139 1197 3140
rect 1191 3135 1192 3139
rect 1196 3138 1197 3139
rect 1206 3139 1212 3140
rect 1206 3138 1207 3139
rect 1196 3136 1207 3138
rect 1196 3135 1197 3136
rect 1191 3134 1197 3135
rect 1206 3135 1207 3136
rect 1211 3135 1212 3139
rect 1206 3134 1212 3135
rect 1375 3139 1381 3140
rect 1375 3135 1376 3139
rect 1380 3138 1381 3139
rect 1390 3139 1396 3140
rect 1390 3138 1391 3139
rect 1380 3136 1391 3138
rect 1380 3135 1381 3136
rect 1375 3134 1381 3135
rect 1390 3135 1391 3136
rect 1395 3135 1396 3139
rect 1390 3134 1396 3135
rect 1478 3139 1484 3140
rect 1478 3135 1479 3139
rect 1483 3138 1484 3139
rect 1567 3139 1573 3140
rect 1567 3138 1568 3139
rect 1483 3136 1568 3138
rect 1483 3135 1484 3136
rect 1478 3134 1484 3135
rect 1567 3135 1568 3136
rect 1572 3135 1573 3139
rect 1567 3134 1573 3135
rect 1743 3139 1749 3140
rect 1743 3135 1744 3139
rect 1748 3138 1749 3139
rect 1758 3139 1764 3140
rect 1758 3138 1759 3139
rect 1748 3136 1759 3138
rect 1748 3135 1749 3136
rect 1743 3134 1749 3135
rect 1758 3135 1759 3136
rect 1763 3135 1764 3139
rect 1758 3134 1764 3135
rect 1902 3134 1908 3135
rect 1902 3130 1903 3134
rect 1907 3130 1908 3134
rect 1902 3129 1908 3130
rect 1998 3134 2004 3135
rect 1998 3130 1999 3134
rect 2003 3130 2004 3134
rect 1998 3129 2004 3130
rect 2126 3134 2132 3135
rect 2126 3130 2127 3134
rect 2131 3130 2132 3134
rect 2126 3129 2132 3130
rect 2254 3134 2260 3135
rect 2254 3130 2255 3134
rect 2259 3130 2260 3134
rect 2254 3129 2260 3130
rect 2390 3134 2396 3135
rect 2390 3130 2391 3134
rect 2395 3130 2396 3134
rect 2390 3129 2396 3130
rect 2518 3134 2524 3135
rect 2518 3130 2519 3134
rect 2523 3130 2524 3134
rect 2518 3129 2524 3130
rect 2646 3134 2652 3135
rect 2646 3130 2647 3134
rect 2651 3130 2652 3134
rect 2646 3129 2652 3130
rect 2774 3134 2780 3135
rect 2774 3130 2775 3134
rect 2779 3130 2780 3134
rect 2774 3129 2780 3130
rect 2902 3134 2908 3135
rect 2902 3130 2903 3134
rect 2907 3130 2908 3134
rect 2902 3129 2908 3130
rect 3038 3134 3044 3135
rect 3038 3130 3039 3134
rect 3043 3130 3044 3134
rect 3038 3129 3044 3130
rect 3182 3134 3188 3135
rect 3182 3130 3183 3134
rect 3187 3130 3188 3134
rect 3182 3129 3188 3130
rect 3334 3134 3340 3135
rect 3334 3130 3335 3134
rect 3339 3130 3340 3134
rect 3334 3129 3340 3130
rect 3494 3134 3500 3135
rect 3494 3130 3495 3134
rect 3499 3130 3500 3134
rect 3494 3129 3500 3130
rect 583 3123 589 3124
rect 583 3119 584 3123
rect 588 3122 589 3123
rect 634 3123 640 3124
rect 634 3122 635 3123
rect 588 3120 635 3122
rect 588 3119 589 3120
rect 583 3118 589 3119
rect 634 3119 635 3120
rect 639 3119 640 3123
rect 634 3118 640 3119
rect 642 3123 648 3124
rect 642 3119 643 3123
rect 647 3122 648 3123
rect 663 3123 669 3124
rect 663 3122 664 3123
rect 647 3120 664 3122
rect 647 3119 648 3120
rect 642 3118 648 3119
rect 663 3119 664 3120
rect 668 3119 669 3123
rect 663 3118 669 3119
rect 722 3123 728 3124
rect 722 3119 723 3123
rect 727 3122 728 3123
rect 751 3123 757 3124
rect 751 3122 752 3123
rect 727 3120 752 3122
rect 727 3119 728 3120
rect 722 3118 728 3119
rect 751 3119 752 3120
rect 756 3119 757 3123
rect 751 3118 757 3119
rect 810 3123 816 3124
rect 810 3119 811 3123
rect 815 3122 816 3123
rect 839 3123 845 3124
rect 839 3122 840 3123
rect 815 3120 840 3122
rect 815 3119 816 3120
rect 810 3118 816 3119
rect 839 3119 840 3120
rect 844 3119 845 3123
rect 839 3118 845 3119
rect 926 3123 933 3124
rect 926 3119 927 3123
rect 932 3119 933 3123
rect 926 3118 933 3119
rect 1015 3123 1021 3124
rect 1015 3119 1016 3123
rect 1020 3122 1021 3123
rect 1066 3123 1072 3124
rect 1066 3122 1067 3123
rect 1020 3120 1067 3122
rect 1020 3119 1021 3120
rect 1015 3118 1021 3119
rect 1066 3119 1067 3120
rect 1071 3119 1072 3123
rect 1066 3118 1072 3119
rect 1074 3123 1080 3124
rect 1074 3119 1075 3123
rect 1079 3122 1080 3123
rect 1103 3123 1109 3124
rect 1103 3122 1104 3123
rect 1079 3120 1104 3122
rect 1079 3119 1080 3120
rect 1074 3118 1080 3119
rect 1103 3119 1104 3120
rect 1108 3119 1109 3123
rect 1103 3118 1109 3119
rect 1162 3123 1168 3124
rect 1162 3119 1163 3123
rect 1167 3122 1168 3123
rect 1191 3123 1197 3124
rect 1191 3122 1192 3123
rect 1167 3120 1192 3122
rect 1167 3119 1168 3120
rect 1162 3118 1168 3119
rect 1191 3119 1192 3120
rect 1196 3119 1197 3123
rect 1191 3118 1197 3119
rect 1250 3123 1256 3124
rect 1250 3119 1251 3123
rect 1255 3122 1256 3123
rect 1279 3123 1285 3124
rect 1279 3122 1280 3123
rect 1255 3120 1280 3122
rect 1255 3119 1256 3120
rect 1250 3118 1256 3119
rect 1279 3119 1280 3120
rect 1284 3119 1285 3123
rect 1279 3118 1285 3119
rect 1338 3123 1344 3124
rect 1338 3119 1339 3123
rect 1343 3122 1344 3123
rect 1367 3123 1373 3124
rect 1367 3122 1368 3123
rect 1343 3120 1368 3122
rect 1343 3119 1344 3120
rect 1338 3118 1344 3119
rect 1367 3119 1368 3120
rect 1372 3119 1373 3123
rect 1367 3118 1373 3119
rect 1818 3123 1824 3124
rect 1818 3119 1819 3123
rect 1823 3122 1824 3123
rect 1895 3123 1901 3124
rect 1895 3122 1896 3123
rect 1823 3120 1896 3122
rect 1823 3119 1824 3120
rect 1818 3118 1824 3119
rect 1895 3119 1896 3120
rect 1900 3119 1901 3123
rect 1895 3118 1901 3119
rect 1962 3123 1968 3124
rect 1962 3119 1963 3123
rect 1967 3122 1968 3123
rect 1991 3123 1997 3124
rect 1991 3122 1992 3123
rect 1967 3120 1992 3122
rect 1967 3119 1968 3120
rect 1962 3118 1968 3119
rect 1991 3119 1992 3120
rect 1996 3119 1997 3123
rect 1991 3118 1997 3119
rect 2062 3123 2068 3124
rect 2062 3119 2063 3123
rect 2067 3122 2068 3123
rect 2119 3123 2125 3124
rect 2119 3122 2120 3123
rect 2067 3120 2120 3122
rect 2067 3119 2068 3120
rect 2062 3118 2068 3119
rect 2119 3119 2120 3120
rect 2124 3119 2125 3123
rect 2119 3118 2125 3119
rect 2247 3123 2253 3124
rect 2247 3119 2248 3123
rect 2252 3122 2253 3123
rect 2350 3123 2356 3124
rect 2350 3122 2351 3123
rect 2252 3120 2351 3122
rect 2252 3119 2253 3120
rect 2247 3118 2253 3119
rect 2350 3119 2351 3120
rect 2355 3119 2356 3123
rect 2350 3118 2356 3119
rect 2383 3123 2389 3124
rect 2383 3119 2384 3123
rect 2388 3122 2389 3123
rect 2414 3123 2420 3124
rect 2414 3122 2415 3123
rect 2388 3120 2415 3122
rect 2388 3119 2389 3120
rect 2383 3118 2389 3119
rect 2414 3119 2415 3120
rect 2419 3119 2420 3123
rect 2414 3118 2420 3119
rect 2511 3123 2517 3124
rect 2511 3119 2512 3123
rect 2516 3122 2517 3123
rect 2550 3123 2556 3124
rect 2550 3122 2551 3123
rect 2516 3120 2551 3122
rect 2516 3119 2517 3120
rect 2511 3118 2517 3119
rect 2550 3119 2551 3120
rect 2555 3119 2556 3123
rect 2550 3118 2556 3119
rect 2582 3123 2588 3124
rect 2582 3119 2583 3123
rect 2587 3122 2588 3123
rect 2639 3123 2645 3124
rect 2639 3122 2640 3123
rect 2587 3120 2640 3122
rect 2587 3119 2588 3120
rect 2582 3118 2588 3119
rect 2639 3119 2640 3120
rect 2644 3119 2645 3123
rect 2639 3118 2645 3119
rect 2710 3123 2716 3124
rect 2710 3119 2711 3123
rect 2715 3122 2716 3123
rect 2767 3123 2773 3124
rect 2767 3122 2768 3123
rect 2715 3120 2768 3122
rect 2715 3119 2716 3120
rect 2710 3118 2716 3119
rect 2767 3119 2768 3120
rect 2772 3119 2773 3123
rect 2767 3118 2773 3119
rect 2838 3123 2844 3124
rect 2838 3119 2839 3123
rect 2843 3122 2844 3123
rect 2895 3123 2901 3124
rect 2895 3122 2896 3123
rect 2843 3120 2896 3122
rect 2843 3119 2844 3120
rect 2838 3118 2844 3119
rect 2895 3119 2896 3120
rect 2900 3119 2901 3123
rect 2895 3118 2901 3119
rect 2970 3123 2976 3124
rect 2970 3119 2971 3123
rect 2975 3122 2976 3123
rect 3031 3123 3037 3124
rect 3031 3122 3032 3123
rect 2975 3120 3032 3122
rect 2975 3119 2976 3120
rect 2970 3118 2976 3119
rect 3031 3119 3032 3120
rect 3036 3119 3037 3123
rect 3031 3118 3037 3119
rect 3098 3123 3104 3124
rect 3098 3119 3099 3123
rect 3103 3122 3104 3123
rect 3175 3123 3181 3124
rect 3175 3122 3176 3123
rect 3103 3120 3176 3122
rect 3103 3119 3104 3120
rect 3098 3118 3104 3119
rect 3175 3119 3176 3120
rect 3180 3119 3181 3123
rect 3175 3118 3181 3119
rect 3258 3123 3264 3124
rect 3258 3119 3259 3123
rect 3263 3122 3264 3123
rect 3327 3123 3333 3124
rect 3327 3122 3328 3123
rect 3263 3120 3328 3122
rect 3263 3119 3264 3120
rect 3258 3118 3264 3119
rect 3327 3119 3328 3120
rect 3332 3119 3333 3123
rect 3327 3118 3333 3119
rect 3426 3123 3432 3124
rect 3426 3119 3427 3123
rect 3431 3122 3432 3123
rect 3487 3123 3493 3124
rect 3487 3122 3488 3123
rect 3431 3120 3488 3122
rect 3431 3119 3432 3120
rect 3426 3118 3432 3119
rect 3487 3119 3488 3120
rect 3492 3119 3493 3123
rect 3487 3118 3493 3119
rect 590 3114 596 3115
rect 590 3110 591 3114
rect 595 3110 596 3114
rect 590 3109 596 3110
rect 670 3114 676 3115
rect 670 3110 671 3114
rect 675 3110 676 3114
rect 670 3109 676 3110
rect 758 3114 764 3115
rect 758 3110 759 3114
rect 763 3110 764 3114
rect 758 3109 764 3110
rect 846 3114 852 3115
rect 846 3110 847 3114
rect 851 3110 852 3114
rect 846 3109 852 3110
rect 934 3114 940 3115
rect 934 3110 935 3114
rect 939 3110 940 3114
rect 934 3109 940 3110
rect 1022 3114 1028 3115
rect 1022 3110 1023 3114
rect 1027 3110 1028 3114
rect 1022 3109 1028 3110
rect 1110 3114 1116 3115
rect 1110 3110 1111 3114
rect 1115 3110 1116 3114
rect 1110 3109 1116 3110
rect 1198 3114 1204 3115
rect 1198 3110 1199 3114
rect 1203 3110 1204 3114
rect 1198 3109 1204 3110
rect 1286 3114 1292 3115
rect 1286 3110 1287 3114
rect 1291 3110 1292 3114
rect 1286 3109 1292 3110
rect 1374 3114 1380 3115
rect 1374 3110 1375 3114
rect 1379 3110 1380 3114
rect 1374 3109 1380 3110
rect 110 3096 116 3097
rect 110 3092 111 3096
rect 115 3092 116 3096
rect 110 3091 116 3092
rect 1830 3096 1836 3097
rect 1830 3092 1831 3096
rect 1835 3092 1836 3096
rect 1830 3091 1836 3092
rect 1895 3095 1901 3096
rect 1895 3091 1896 3095
rect 1900 3094 1901 3095
rect 1910 3095 1916 3096
rect 1910 3094 1911 3095
rect 1900 3092 1911 3094
rect 1900 3091 1901 3092
rect 1895 3090 1901 3091
rect 1910 3091 1911 3092
rect 1915 3091 1916 3095
rect 1910 3090 1916 3091
rect 1954 3095 1960 3096
rect 1954 3091 1955 3095
rect 1959 3094 1960 3095
rect 2007 3095 2013 3096
rect 2007 3094 2008 3095
rect 1959 3092 2008 3094
rect 1959 3091 1960 3092
rect 1954 3090 1960 3091
rect 2007 3091 2008 3092
rect 2012 3091 2013 3095
rect 2007 3090 2013 3091
rect 2178 3095 2189 3096
rect 2178 3091 2179 3095
rect 2183 3091 2184 3095
rect 2188 3091 2189 3095
rect 2178 3090 2189 3091
rect 2346 3095 2352 3096
rect 2346 3091 2347 3095
rect 2351 3094 2352 3095
rect 2399 3095 2405 3096
rect 2399 3094 2400 3095
rect 2351 3092 2400 3094
rect 2351 3091 2352 3092
rect 2346 3090 2352 3091
rect 2399 3091 2400 3092
rect 2404 3091 2405 3095
rect 2399 3090 2405 3091
rect 2458 3095 2464 3096
rect 2458 3091 2459 3095
rect 2463 3094 2464 3095
rect 2647 3095 2653 3096
rect 2647 3094 2648 3095
rect 2463 3092 2648 3094
rect 2463 3091 2464 3092
rect 2458 3090 2464 3091
rect 2647 3091 2648 3092
rect 2652 3091 2653 3095
rect 2647 3090 2653 3091
rect 2706 3095 2712 3096
rect 2706 3091 2707 3095
rect 2711 3094 2712 3095
rect 2927 3095 2933 3096
rect 2927 3094 2928 3095
rect 2711 3092 2928 3094
rect 2711 3091 2712 3092
rect 2706 3090 2712 3091
rect 2927 3091 2928 3092
rect 2932 3091 2933 3095
rect 2927 3090 2933 3091
rect 3223 3095 3229 3096
rect 3223 3091 3224 3095
rect 3228 3094 3229 3095
rect 3238 3095 3244 3096
rect 3238 3094 3239 3095
rect 3228 3092 3239 3094
rect 3228 3091 3229 3092
rect 3223 3090 3229 3091
rect 3238 3091 3239 3092
rect 3243 3091 3244 3095
rect 3238 3090 3244 3091
rect 3282 3095 3288 3096
rect 3282 3091 3283 3095
rect 3287 3094 3288 3095
rect 3503 3095 3509 3096
rect 3503 3094 3504 3095
rect 3287 3092 3504 3094
rect 3287 3091 3288 3092
rect 3282 3090 3288 3091
rect 3503 3091 3504 3092
rect 3508 3091 3509 3095
rect 3503 3090 3509 3091
rect 642 3087 648 3088
rect 642 3083 643 3087
rect 647 3083 648 3087
rect 642 3082 648 3083
rect 722 3087 728 3088
rect 722 3083 723 3087
rect 727 3083 728 3087
rect 722 3082 728 3083
rect 810 3087 816 3088
rect 810 3083 811 3087
rect 815 3083 816 3087
rect 926 3087 932 3088
rect 926 3086 927 3087
rect 901 3084 927 3086
rect 810 3082 816 3083
rect 926 3083 927 3084
rect 931 3083 932 3087
rect 926 3082 932 3083
rect 986 3087 992 3088
rect 986 3083 987 3087
rect 991 3083 992 3087
rect 986 3082 992 3083
rect 1074 3087 1080 3088
rect 1074 3083 1075 3087
rect 1079 3083 1080 3087
rect 1074 3082 1080 3083
rect 1162 3087 1168 3088
rect 1162 3083 1163 3087
rect 1167 3083 1168 3087
rect 1162 3082 1168 3083
rect 1250 3087 1256 3088
rect 1250 3083 1251 3087
rect 1255 3083 1256 3087
rect 1250 3082 1256 3083
rect 1338 3087 1344 3088
rect 1338 3083 1339 3087
rect 1343 3083 1344 3087
rect 1338 3082 1344 3083
rect 1390 3087 1396 3088
rect 1390 3083 1391 3087
rect 1395 3083 1396 3087
rect 1390 3082 1396 3083
rect 1902 3086 1908 3087
rect 1902 3082 1903 3086
rect 1907 3082 1908 3086
rect 1902 3081 1908 3082
rect 2014 3086 2020 3087
rect 2014 3082 2015 3086
rect 2019 3082 2020 3086
rect 2014 3081 2020 3082
rect 2190 3086 2196 3087
rect 2190 3082 2191 3086
rect 2195 3082 2196 3086
rect 2190 3081 2196 3082
rect 2406 3086 2412 3087
rect 2406 3082 2407 3086
rect 2411 3082 2412 3086
rect 2406 3081 2412 3082
rect 2654 3086 2660 3087
rect 2654 3082 2655 3086
rect 2659 3082 2660 3086
rect 2654 3081 2660 3082
rect 2934 3086 2940 3087
rect 2934 3082 2935 3086
rect 2939 3082 2940 3086
rect 2934 3081 2940 3082
rect 3230 3086 3236 3087
rect 3230 3082 3231 3086
rect 3235 3082 3236 3086
rect 3230 3081 3236 3082
rect 3510 3086 3516 3087
rect 3510 3082 3511 3086
rect 3515 3082 3516 3086
rect 3510 3081 3516 3082
rect 110 3079 116 3080
rect 110 3075 111 3079
rect 115 3075 116 3079
rect 1830 3079 1836 3080
rect 110 3074 116 3075
rect 582 3076 588 3077
rect 582 3072 583 3076
rect 587 3072 588 3076
rect 582 3071 588 3072
rect 662 3076 668 3077
rect 662 3072 663 3076
rect 667 3072 668 3076
rect 662 3071 668 3072
rect 750 3076 756 3077
rect 750 3072 751 3076
rect 755 3072 756 3076
rect 750 3071 756 3072
rect 838 3076 844 3077
rect 838 3072 839 3076
rect 843 3072 844 3076
rect 838 3071 844 3072
rect 926 3076 932 3077
rect 926 3072 927 3076
rect 931 3072 932 3076
rect 926 3071 932 3072
rect 1014 3076 1020 3077
rect 1014 3072 1015 3076
rect 1019 3072 1020 3076
rect 1014 3071 1020 3072
rect 1102 3076 1108 3077
rect 1102 3072 1103 3076
rect 1107 3072 1108 3076
rect 1102 3071 1108 3072
rect 1190 3076 1196 3077
rect 1190 3072 1191 3076
rect 1195 3072 1196 3076
rect 1190 3071 1196 3072
rect 1278 3076 1284 3077
rect 1278 3072 1279 3076
rect 1283 3072 1284 3076
rect 1278 3071 1284 3072
rect 1366 3076 1372 3077
rect 1366 3072 1367 3076
rect 1371 3072 1372 3076
rect 1830 3075 1831 3079
rect 1835 3075 1836 3079
rect 1830 3074 1836 3075
rect 1366 3071 1372 3072
rect 1870 3068 1876 3069
rect 1870 3064 1871 3068
rect 1875 3064 1876 3068
rect 1870 3063 1876 3064
rect 3590 3068 3596 3069
rect 3590 3064 3591 3068
rect 3595 3064 3596 3068
rect 3590 3063 3596 3064
rect 1954 3059 1960 3060
rect 1954 3055 1955 3059
rect 1959 3055 1960 3059
rect 1954 3054 1960 3055
rect 2038 3059 2044 3060
rect 2038 3055 2039 3059
rect 2043 3055 2044 3059
rect 2038 3054 2044 3055
rect 2198 3059 2204 3060
rect 2198 3055 2199 3059
rect 2203 3055 2204 3059
rect 2198 3054 2204 3055
rect 2458 3059 2464 3060
rect 2458 3055 2459 3059
rect 2463 3055 2464 3059
rect 2458 3054 2464 3055
rect 2706 3059 2712 3060
rect 2706 3055 2707 3059
rect 2711 3055 2712 3059
rect 2706 3054 2712 3055
rect 2942 3059 2948 3060
rect 2942 3055 2943 3059
rect 2947 3055 2948 3059
rect 2942 3054 2948 3055
rect 3282 3059 3288 3060
rect 3282 3055 3283 3059
rect 3287 3055 3288 3059
rect 3282 3054 3288 3055
rect 1870 3051 1876 3052
rect 1870 3047 1871 3051
rect 1875 3047 1876 3051
rect 3590 3051 3596 3052
rect 1870 3046 1876 3047
rect 1894 3048 1900 3049
rect 1894 3044 1895 3048
rect 1899 3044 1900 3048
rect 1894 3043 1900 3044
rect 2006 3048 2012 3049
rect 2006 3044 2007 3048
rect 2011 3044 2012 3048
rect 2006 3043 2012 3044
rect 2182 3048 2188 3049
rect 2182 3044 2183 3048
rect 2187 3044 2188 3048
rect 2182 3043 2188 3044
rect 2398 3048 2404 3049
rect 2398 3044 2399 3048
rect 2403 3044 2404 3048
rect 2398 3043 2404 3044
rect 2646 3048 2652 3049
rect 2646 3044 2647 3048
rect 2651 3044 2652 3048
rect 2646 3043 2652 3044
rect 2926 3048 2932 3049
rect 2926 3044 2927 3048
rect 2931 3044 2932 3048
rect 2926 3043 2932 3044
rect 3222 3048 3228 3049
rect 3222 3044 3223 3048
rect 3227 3044 3228 3048
rect 3222 3043 3228 3044
rect 3502 3048 3508 3049
rect 3502 3044 3503 3048
rect 3507 3044 3508 3048
rect 3590 3047 3591 3051
rect 3595 3047 3596 3051
rect 3590 3046 3596 3047
rect 3502 3043 3508 3044
rect 3518 3031 3525 3032
rect 542 3028 548 3029
rect 110 3025 116 3026
rect 110 3021 111 3025
rect 115 3021 116 3025
rect 542 3024 543 3028
rect 547 3024 548 3028
rect 542 3023 548 3024
rect 622 3028 628 3029
rect 622 3024 623 3028
rect 627 3024 628 3028
rect 622 3023 628 3024
rect 710 3028 716 3029
rect 710 3024 711 3028
rect 715 3024 716 3028
rect 710 3023 716 3024
rect 806 3028 812 3029
rect 806 3024 807 3028
rect 811 3024 812 3028
rect 806 3023 812 3024
rect 902 3028 908 3029
rect 902 3024 903 3028
rect 907 3024 908 3028
rect 902 3023 908 3024
rect 998 3028 1004 3029
rect 998 3024 999 3028
rect 1003 3024 1004 3028
rect 998 3023 1004 3024
rect 1086 3028 1092 3029
rect 1086 3024 1087 3028
rect 1091 3024 1092 3028
rect 1086 3023 1092 3024
rect 1182 3028 1188 3029
rect 1182 3024 1183 3028
rect 1187 3024 1188 3028
rect 1182 3023 1188 3024
rect 1278 3028 1284 3029
rect 1278 3024 1279 3028
rect 1283 3024 1284 3028
rect 1278 3023 1284 3024
rect 1374 3028 1380 3029
rect 1374 3024 1375 3028
rect 1379 3024 1380 3028
rect 1374 3023 1380 3024
rect 1470 3028 1476 3029
rect 1470 3024 1471 3028
rect 1475 3024 1476 3028
rect 3518 3027 3519 3031
rect 3524 3027 3525 3031
rect 3518 3026 3525 3027
rect 1470 3023 1476 3024
rect 1830 3025 1836 3026
rect 110 3020 116 3021
rect 1830 3021 1831 3025
rect 1835 3021 1836 3025
rect 1830 3020 1836 3021
rect 610 3019 616 3020
rect 610 3018 611 3019
rect 605 3016 611 3018
rect 610 3015 611 3016
rect 615 3015 616 3019
rect 694 3019 700 3020
rect 694 3018 695 3019
rect 685 3016 695 3018
rect 610 3014 616 3015
rect 694 3015 695 3016
rect 699 3015 700 3019
rect 778 3019 784 3020
rect 694 3014 700 3015
rect 602 3011 608 3012
rect 110 3008 116 3009
rect 110 3004 111 3008
rect 115 3004 116 3008
rect 602 3007 603 3011
rect 607 3010 608 3011
rect 728 3010 730 3017
rect 778 3015 779 3019
rect 783 3018 784 3019
rect 874 3019 880 3020
rect 783 3016 825 3018
rect 783 3015 784 3016
rect 778 3014 784 3015
rect 874 3015 875 3019
rect 879 3018 880 3019
rect 970 3019 976 3020
rect 879 3016 921 3018
rect 879 3015 880 3016
rect 874 3014 880 3015
rect 970 3015 971 3019
rect 975 3018 976 3019
rect 1066 3019 1072 3020
rect 975 3016 1017 3018
rect 975 3015 976 3016
rect 970 3014 976 3015
rect 1066 3015 1067 3019
rect 1071 3018 1072 3019
rect 1154 3019 1160 3020
rect 1071 3016 1105 3018
rect 1071 3015 1072 3016
rect 1066 3014 1072 3015
rect 1154 3015 1155 3019
rect 1159 3018 1160 3019
rect 1254 3019 1260 3020
rect 1159 3016 1201 3018
rect 1159 3015 1160 3016
rect 1154 3014 1160 3015
rect 1254 3015 1255 3019
rect 1259 3018 1260 3019
rect 1346 3019 1352 3020
rect 1259 3016 1297 3018
rect 1259 3015 1260 3016
rect 1254 3014 1260 3015
rect 1346 3015 1347 3019
rect 1351 3018 1352 3019
rect 1442 3019 1448 3020
rect 1351 3016 1393 3018
rect 1351 3015 1352 3016
rect 1346 3014 1352 3015
rect 1442 3015 1443 3019
rect 1447 3018 1448 3019
rect 1447 3016 1489 3018
rect 1447 3015 1448 3016
rect 1442 3014 1448 3015
rect 607 3008 730 3010
rect 1830 3008 1836 3009
rect 607 3007 608 3008
rect 602 3006 608 3007
rect 110 3003 116 3004
rect 1830 3004 1831 3008
rect 1835 3004 1836 3008
rect 1830 3003 1836 3004
rect 1894 2996 1900 2997
rect 1870 2993 1876 2994
rect 550 2990 556 2991
rect 550 2986 551 2990
rect 555 2986 556 2990
rect 550 2985 556 2986
rect 630 2990 636 2991
rect 630 2986 631 2990
rect 635 2986 636 2990
rect 630 2985 636 2986
rect 718 2990 724 2991
rect 718 2986 719 2990
rect 723 2986 724 2990
rect 718 2985 724 2986
rect 814 2990 820 2991
rect 814 2986 815 2990
rect 819 2986 820 2990
rect 814 2985 820 2986
rect 910 2990 916 2991
rect 910 2986 911 2990
rect 915 2986 916 2990
rect 910 2985 916 2986
rect 1006 2990 1012 2991
rect 1006 2986 1007 2990
rect 1011 2986 1012 2990
rect 1006 2985 1012 2986
rect 1094 2990 1100 2991
rect 1094 2986 1095 2990
rect 1099 2986 1100 2990
rect 1094 2985 1100 2986
rect 1190 2990 1196 2991
rect 1190 2986 1191 2990
rect 1195 2986 1196 2990
rect 1190 2985 1196 2986
rect 1286 2990 1292 2991
rect 1286 2986 1287 2990
rect 1291 2986 1292 2990
rect 1286 2985 1292 2986
rect 1382 2990 1388 2991
rect 1382 2986 1383 2990
rect 1387 2986 1388 2990
rect 1382 2985 1388 2986
rect 1478 2990 1484 2991
rect 1478 2986 1479 2990
rect 1483 2986 1484 2990
rect 1870 2989 1871 2993
rect 1875 2989 1876 2993
rect 1894 2992 1895 2996
rect 1899 2992 1900 2996
rect 1894 2991 1900 2992
rect 2046 2996 2052 2997
rect 2046 2992 2047 2996
rect 2051 2992 2052 2996
rect 2046 2991 2052 2992
rect 2222 2996 2228 2997
rect 2222 2992 2223 2996
rect 2227 2992 2228 2996
rect 2222 2991 2228 2992
rect 2390 2996 2396 2997
rect 2390 2992 2391 2996
rect 2395 2992 2396 2996
rect 2390 2991 2396 2992
rect 2542 2996 2548 2997
rect 2542 2992 2543 2996
rect 2547 2992 2548 2996
rect 2542 2991 2548 2992
rect 2686 2996 2692 2997
rect 2686 2992 2687 2996
rect 2691 2992 2692 2996
rect 2686 2991 2692 2992
rect 2814 2996 2820 2997
rect 2814 2992 2815 2996
rect 2819 2992 2820 2996
rect 2814 2991 2820 2992
rect 2926 2996 2932 2997
rect 2926 2992 2927 2996
rect 2931 2992 2932 2996
rect 2926 2991 2932 2992
rect 3038 2996 3044 2997
rect 3038 2992 3039 2996
rect 3043 2992 3044 2996
rect 3038 2991 3044 2992
rect 3142 2996 3148 2997
rect 3142 2992 3143 2996
rect 3147 2992 3148 2996
rect 3142 2991 3148 2992
rect 3238 2996 3244 2997
rect 3238 2992 3239 2996
rect 3243 2992 3244 2996
rect 3238 2991 3244 2992
rect 3334 2996 3340 2997
rect 3334 2992 3335 2996
rect 3339 2992 3340 2996
rect 3334 2991 3340 2992
rect 3422 2996 3428 2997
rect 3422 2992 3423 2996
rect 3427 2992 3428 2996
rect 3422 2991 3428 2992
rect 3502 2996 3508 2997
rect 3502 2992 3503 2996
rect 3507 2992 3508 2996
rect 3502 2991 3508 2992
rect 3590 2993 3596 2994
rect 1870 2988 1876 2989
rect 3590 2989 3591 2993
rect 3595 2989 3596 2993
rect 3590 2988 3596 2989
rect 1962 2987 1968 2988
rect 1478 2985 1484 2986
rect 1896 2984 1913 2986
rect 1894 2983 1900 2984
rect 543 2979 549 2980
rect 543 2975 544 2979
rect 548 2978 549 2979
rect 602 2979 608 2980
rect 602 2978 603 2979
rect 548 2976 603 2978
rect 548 2975 549 2976
rect 543 2974 549 2975
rect 602 2975 603 2976
rect 607 2975 608 2979
rect 602 2974 608 2975
rect 610 2979 616 2980
rect 610 2975 611 2979
rect 615 2978 616 2979
rect 623 2979 629 2980
rect 623 2978 624 2979
rect 615 2976 624 2978
rect 615 2975 616 2976
rect 610 2974 616 2975
rect 623 2975 624 2976
rect 628 2975 629 2979
rect 623 2974 629 2975
rect 711 2979 717 2980
rect 711 2975 712 2979
rect 716 2978 717 2979
rect 778 2979 784 2980
rect 778 2978 779 2979
rect 716 2976 779 2978
rect 716 2975 717 2976
rect 711 2974 717 2975
rect 778 2975 779 2976
rect 783 2975 784 2979
rect 778 2974 784 2975
rect 807 2979 813 2980
rect 807 2975 808 2979
rect 812 2978 813 2979
rect 874 2979 880 2980
rect 874 2978 875 2979
rect 812 2976 875 2978
rect 812 2975 813 2976
rect 807 2974 813 2975
rect 874 2975 875 2976
rect 879 2975 880 2979
rect 874 2974 880 2975
rect 903 2979 909 2980
rect 903 2975 904 2979
rect 908 2978 909 2979
rect 970 2979 976 2980
rect 970 2978 971 2979
rect 908 2976 971 2978
rect 908 2975 909 2976
rect 903 2974 909 2975
rect 970 2975 971 2976
rect 975 2975 976 2979
rect 970 2974 976 2975
rect 986 2979 992 2980
rect 986 2975 987 2979
rect 991 2978 992 2979
rect 999 2979 1005 2980
rect 999 2978 1000 2979
rect 991 2976 1000 2978
rect 991 2975 992 2976
rect 986 2974 992 2975
rect 999 2975 1000 2976
rect 1004 2975 1005 2979
rect 999 2974 1005 2975
rect 1087 2979 1093 2980
rect 1087 2975 1088 2979
rect 1092 2978 1093 2979
rect 1154 2979 1160 2980
rect 1154 2978 1155 2979
rect 1092 2976 1155 2978
rect 1092 2975 1093 2976
rect 1087 2974 1093 2975
rect 1154 2975 1155 2976
rect 1159 2975 1160 2979
rect 1154 2974 1160 2975
rect 1183 2979 1189 2980
rect 1183 2975 1184 2979
rect 1188 2978 1189 2979
rect 1254 2979 1260 2980
rect 1254 2978 1255 2979
rect 1188 2976 1255 2978
rect 1188 2975 1189 2976
rect 1183 2974 1189 2975
rect 1254 2975 1255 2976
rect 1259 2975 1260 2979
rect 1254 2974 1260 2975
rect 1279 2979 1285 2980
rect 1279 2975 1280 2979
rect 1284 2978 1285 2979
rect 1346 2979 1352 2980
rect 1346 2978 1347 2979
rect 1284 2976 1347 2978
rect 1284 2975 1285 2976
rect 1279 2974 1285 2975
rect 1346 2975 1347 2976
rect 1351 2975 1352 2979
rect 1346 2974 1352 2975
rect 1375 2979 1381 2980
rect 1375 2975 1376 2979
rect 1380 2978 1381 2979
rect 1442 2979 1448 2980
rect 1442 2978 1443 2979
rect 1380 2976 1443 2978
rect 1380 2975 1381 2976
rect 1375 2974 1381 2975
rect 1442 2975 1443 2976
rect 1447 2975 1448 2979
rect 1442 2974 1448 2975
rect 1471 2979 1477 2980
rect 1471 2975 1472 2979
rect 1476 2978 1477 2979
rect 1598 2979 1604 2980
rect 1598 2978 1599 2979
rect 1476 2976 1599 2978
rect 1476 2975 1477 2976
rect 1471 2974 1477 2975
rect 1598 2975 1599 2976
rect 1603 2975 1604 2979
rect 1894 2979 1895 2983
rect 1899 2979 1900 2983
rect 1962 2983 1963 2987
rect 1967 2986 1968 2987
rect 2346 2987 2352 2988
rect 2346 2986 2347 2987
rect 1967 2984 2065 2986
rect 2285 2984 2347 2986
rect 1967 2983 1968 2984
rect 1962 2982 1968 2983
rect 2346 2983 2347 2984
rect 2351 2983 2352 2987
rect 2346 2982 2352 2983
rect 2354 2987 2360 2988
rect 2354 2983 2355 2987
rect 2359 2986 2360 2987
rect 2610 2987 2616 2988
rect 2610 2986 2611 2987
rect 2359 2984 2409 2986
rect 2605 2984 2611 2986
rect 2359 2983 2360 2984
rect 2354 2982 2360 2983
rect 2610 2983 2611 2984
rect 2615 2983 2616 2987
rect 2758 2987 2764 2988
rect 2758 2986 2759 2987
rect 2749 2984 2759 2986
rect 2610 2982 2616 2983
rect 2758 2983 2759 2984
rect 2763 2983 2764 2987
rect 2910 2987 2916 2988
rect 2910 2986 2911 2987
rect 2877 2984 2911 2986
rect 2758 2982 2764 2983
rect 2910 2983 2911 2984
rect 2915 2983 2916 2987
rect 2910 2982 2916 2983
rect 2918 2987 2924 2988
rect 2918 2983 2919 2987
rect 2923 2986 2924 2987
rect 2999 2987 3005 2988
rect 2923 2984 2945 2986
rect 2923 2983 2924 2984
rect 2918 2982 2924 2983
rect 2999 2983 3000 2987
rect 3004 2986 3005 2987
rect 3106 2987 3112 2988
rect 3004 2984 3057 2986
rect 3004 2983 3005 2984
rect 2999 2982 3005 2983
rect 3106 2983 3107 2987
rect 3111 2986 3112 2987
rect 3210 2987 3216 2988
rect 3111 2984 3161 2986
rect 3111 2983 3112 2984
rect 3106 2982 3112 2983
rect 3210 2983 3211 2987
rect 3215 2986 3216 2987
rect 3402 2987 3408 2988
rect 3402 2986 3403 2987
rect 3215 2984 3257 2986
rect 3397 2984 3403 2986
rect 3215 2983 3216 2984
rect 3210 2982 3216 2983
rect 3402 2983 3403 2984
rect 3407 2983 3408 2987
rect 3490 2987 3496 2988
rect 3424 2984 3441 2986
rect 3402 2982 3408 2983
rect 3422 2983 3428 2984
rect 1894 2978 1900 2979
rect 3422 2979 3423 2983
rect 3427 2979 3428 2983
rect 3490 2983 3491 2987
rect 3495 2986 3496 2987
rect 3495 2984 3521 2986
rect 3495 2983 3496 2984
rect 3490 2982 3496 2983
rect 3422 2978 3428 2979
rect 1598 2974 1604 2975
rect 1870 2976 1876 2977
rect 1870 2972 1871 2976
rect 1875 2972 1876 2976
rect 1870 2971 1876 2972
rect 3590 2976 3596 2977
rect 3590 2972 3591 2976
rect 3595 2972 3596 2976
rect 3590 2971 3596 2972
rect 463 2967 469 2968
rect 463 2963 464 2967
rect 468 2966 469 2967
rect 530 2967 536 2968
rect 530 2966 531 2967
rect 468 2964 531 2966
rect 468 2963 469 2964
rect 463 2962 469 2963
rect 530 2963 531 2964
rect 535 2963 536 2967
rect 530 2962 536 2963
rect 567 2967 573 2968
rect 567 2963 568 2967
rect 572 2966 573 2967
rect 654 2967 660 2968
rect 654 2966 655 2967
rect 572 2964 655 2966
rect 572 2963 573 2964
rect 567 2962 573 2963
rect 654 2963 655 2964
rect 659 2963 660 2967
rect 654 2962 660 2963
rect 679 2967 685 2968
rect 679 2963 680 2967
rect 684 2966 685 2967
rect 694 2967 700 2968
rect 694 2966 695 2967
rect 684 2964 695 2966
rect 684 2963 685 2964
rect 679 2962 685 2963
rect 694 2963 695 2964
rect 699 2963 700 2967
rect 694 2962 700 2963
rect 738 2967 744 2968
rect 738 2963 739 2967
rect 743 2966 744 2967
rect 799 2967 805 2968
rect 799 2966 800 2967
rect 743 2964 800 2966
rect 743 2963 744 2964
rect 738 2962 744 2963
rect 799 2963 800 2964
rect 804 2963 805 2967
rect 799 2962 805 2963
rect 858 2967 864 2968
rect 858 2963 859 2967
rect 863 2966 864 2967
rect 935 2967 941 2968
rect 935 2966 936 2967
rect 863 2964 936 2966
rect 863 2963 864 2964
rect 858 2962 864 2963
rect 935 2963 936 2964
rect 940 2963 941 2967
rect 935 2962 941 2963
rect 1079 2967 1085 2968
rect 1079 2963 1080 2967
rect 1084 2966 1085 2967
rect 1102 2967 1108 2968
rect 1102 2966 1103 2967
rect 1084 2964 1103 2966
rect 1084 2963 1085 2964
rect 1079 2962 1085 2963
rect 1102 2963 1103 2964
rect 1107 2963 1108 2967
rect 1102 2962 1108 2963
rect 1138 2967 1144 2968
rect 1138 2963 1139 2967
rect 1143 2966 1144 2967
rect 1239 2967 1245 2968
rect 1239 2966 1240 2967
rect 1143 2964 1240 2966
rect 1143 2963 1144 2964
rect 1138 2962 1144 2963
rect 1239 2963 1240 2964
rect 1244 2963 1245 2967
rect 1239 2962 1245 2963
rect 1298 2967 1304 2968
rect 1298 2963 1299 2967
rect 1303 2966 1304 2967
rect 1407 2967 1413 2968
rect 1407 2966 1408 2967
rect 1303 2964 1408 2966
rect 1303 2963 1304 2964
rect 1298 2962 1304 2963
rect 1407 2963 1408 2964
rect 1412 2963 1413 2967
rect 1407 2962 1413 2963
rect 1466 2967 1472 2968
rect 1466 2963 1467 2967
rect 1471 2966 1472 2967
rect 1583 2967 1589 2968
rect 1583 2966 1584 2967
rect 1471 2964 1584 2966
rect 1471 2963 1472 2964
rect 1466 2962 1472 2963
rect 1583 2963 1584 2964
rect 1588 2963 1589 2967
rect 1583 2962 1589 2963
rect 1743 2967 1749 2968
rect 1743 2963 1744 2967
rect 1748 2966 1749 2967
rect 1798 2967 1804 2968
rect 1798 2966 1799 2967
rect 1748 2964 1799 2966
rect 1748 2963 1749 2964
rect 1743 2962 1749 2963
rect 1798 2963 1799 2964
rect 1803 2963 1804 2967
rect 1798 2962 1804 2963
rect 3394 2967 3400 2968
rect 3394 2963 3395 2967
rect 3399 2966 3400 2967
rect 3490 2967 3496 2968
rect 3490 2966 3491 2967
rect 3399 2964 3491 2966
rect 3399 2963 3400 2964
rect 3394 2962 3400 2963
rect 3490 2963 3491 2964
rect 3495 2963 3496 2967
rect 3490 2962 3496 2963
rect 470 2958 476 2959
rect 470 2954 471 2958
rect 475 2954 476 2958
rect 470 2953 476 2954
rect 574 2958 580 2959
rect 574 2954 575 2958
rect 579 2954 580 2958
rect 574 2953 580 2954
rect 686 2958 692 2959
rect 686 2954 687 2958
rect 691 2954 692 2958
rect 686 2953 692 2954
rect 806 2958 812 2959
rect 806 2954 807 2958
rect 811 2954 812 2958
rect 806 2953 812 2954
rect 942 2958 948 2959
rect 942 2954 943 2958
rect 947 2954 948 2958
rect 942 2953 948 2954
rect 1086 2958 1092 2959
rect 1086 2954 1087 2958
rect 1091 2954 1092 2958
rect 1086 2953 1092 2954
rect 1246 2958 1252 2959
rect 1246 2954 1247 2958
rect 1251 2954 1252 2958
rect 1246 2953 1252 2954
rect 1414 2958 1420 2959
rect 1414 2954 1415 2958
rect 1419 2954 1420 2958
rect 1414 2953 1420 2954
rect 1590 2958 1596 2959
rect 1590 2954 1591 2958
rect 1595 2954 1596 2958
rect 1590 2953 1596 2954
rect 1750 2958 1756 2959
rect 1750 2954 1751 2958
rect 1755 2954 1756 2958
rect 1750 2953 1756 2954
rect 1902 2958 1908 2959
rect 1902 2954 1903 2958
rect 1907 2954 1908 2958
rect 1902 2953 1908 2954
rect 2054 2958 2060 2959
rect 2054 2954 2055 2958
rect 2059 2954 2060 2958
rect 2054 2953 2060 2954
rect 2230 2958 2236 2959
rect 2230 2954 2231 2958
rect 2235 2954 2236 2958
rect 2230 2953 2236 2954
rect 2398 2958 2404 2959
rect 2398 2954 2399 2958
rect 2403 2954 2404 2958
rect 2398 2953 2404 2954
rect 2550 2958 2556 2959
rect 2550 2954 2551 2958
rect 2555 2954 2556 2958
rect 2550 2953 2556 2954
rect 2694 2958 2700 2959
rect 2694 2954 2695 2958
rect 2699 2954 2700 2958
rect 2694 2953 2700 2954
rect 2822 2958 2828 2959
rect 2822 2954 2823 2958
rect 2827 2954 2828 2958
rect 2822 2953 2828 2954
rect 2934 2958 2940 2959
rect 2934 2954 2935 2958
rect 2939 2954 2940 2958
rect 2934 2953 2940 2954
rect 3046 2958 3052 2959
rect 3046 2954 3047 2958
rect 3051 2954 3052 2958
rect 3046 2953 3052 2954
rect 3150 2958 3156 2959
rect 3150 2954 3151 2958
rect 3155 2954 3156 2958
rect 3150 2953 3156 2954
rect 3246 2958 3252 2959
rect 3246 2954 3247 2958
rect 3251 2954 3252 2958
rect 3246 2953 3252 2954
rect 3342 2958 3348 2959
rect 3342 2954 3343 2958
rect 3347 2954 3348 2958
rect 3342 2953 3348 2954
rect 3430 2958 3436 2959
rect 3430 2954 3431 2958
rect 3435 2954 3436 2958
rect 3430 2953 3436 2954
rect 3510 2958 3516 2959
rect 3510 2954 3511 2958
rect 3515 2954 3516 2958
rect 3510 2953 3516 2954
rect 1895 2947 1901 2948
rect 1895 2943 1896 2947
rect 1900 2946 1901 2947
rect 1962 2947 1968 2948
rect 1962 2946 1963 2947
rect 1900 2944 1963 2946
rect 1900 2943 1901 2944
rect 1895 2942 1901 2943
rect 1962 2943 1963 2944
rect 1967 2943 1968 2947
rect 1962 2942 1968 2943
rect 2038 2947 2044 2948
rect 2038 2943 2039 2947
rect 2043 2946 2044 2947
rect 2047 2947 2053 2948
rect 2047 2946 2048 2947
rect 2043 2944 2048 2946
rect 2043 2943 2044 2944
rect 2038 2942 2044 2943
rect 2047 2943 2048 2944
rect 2052 2943 2053 2947
rect 2047 2942 2053 2943
rect 2223 2947 2229 2948
rect 2223 2943 2224 2947
rect 2228 2946 2229 2947
rect 2354 2947 2360 2948
rect 2354 2946 2355 2947
rect 2228 2944 2355 2946
rect 2228 2943 2229 2944
rect 2223 2942 2229 2943
rect 2354 2943 2355 2944
rect 2359 2943 2360 2947
rect 2354 2942 2360 2943
rect 2391 2947 2397 2948
rect 2391 2943 2392 2947
rect 2396 2946 2397 2947
rect 2494 2947 2500 2948
rect 2494 2946 2495 2947
rect 2396 2944 2495 2946
rect 2396 2943 2397 2944
rect 2391 2942 2397 2943
rect 2494 2943 2495 2944
rect 2499 2943 2500 2947
rect 2494 2942 2500 2943
rect 2543 2947 2549 2948
rect 2543 2943 2544 2947
rect 2548 2946 2549 2947
rect 2566 2947 2572 2948
rect 2566 2946 2567 2947
rect 2548 2944 2567 2946
rect 2548 2943 2549 2944
rect 2543 2942 2549 2943
rect 2566 2943 2567 2944
rect 2571 2943 2572 2947
rect 2566 2942 2572 2943
rect 2610 2947 2616 2948
rect 2610 2943 2611 2947
rect 2615 2946 2616 2947
rect 2687 2947 2693 2948
rect 2687 2946 2688 2947
rect 2615 2944 2688 2946
rect 2615 2943 2616 2944
rect 2610 2942 2616 2943
rect 2687 2943 2688 2944
rect 2692 2943 2693 2947
rect 2687 2942 2693 2943
rect 2758 2947 2764 2948
rect 2758 2943 2759 2947
rect 2763 2946 2764 2947
rect 2815 2947 2821 2948
rect 2815 2946 2816 2947
rect 2763 2944 2816 2946
rect 2763 2943 2764 2944
rect 2758 2942 2764 2943
rect 2815 2943 2816 2944
rect 2820 2943 2821 2947
rect 2815 2942 2821 2943
rect 2927 2947 2933 2948
rect 2927 2943 2928 2947
rect 2932 2946 2933 2947
rect 2999 2947 3005 2948
rect 2999 2946 3000 2947
rect 2932 2944 3000 2946
rect 2932 2943 2933 2944
rect 2927 2942 2933 2943
rect 2999 2943 3000 2944
rect 3004 2943 3005 2947
rect 2999 2942 3005 2943
rect 3039 2947 3045 2948
rect 3039 2943 3040 2947
rect 3044 2946 3045 2947
rect 3106 2947 3112 2948
rect 3106 2946 3107 2947
rect 3044 2944 3107 2946
rect 3044 2943 3045 2944
rect 3039 2942 3045 2943
rect 3106 2943 3107 2944
rect 3111 2943 3112 2947
rect 3106 2942 3112 2943
rect 3143 2947 3149 2948
rect 3143 2943 3144 2947
rect 3148 2946 3149 2947
rect 3210 2947 3216 2948
rect 3210 2946 3211 2947
rect 3148 2944 3211 2946
rect 3148 2943 3149 2944
rect 3143 2942 3149 2943
rect 3210 2943 3211 2944
rect 3215 2943 3216 2947
rect 3210 2942 3216 2943
rect 3239 2947 3245 2948
rect 3239 2943 3240 2947
rect 3244 2946 3245 2947
rect 3335 2947 3341 2948
rect 3244 2944 3330 2946
rect 3244 2943 3245 2944
rect 3239 2942 3245 2943
rect 110 2940 116 2941
rect 110 2936 111 2940
rect 115 2936 116 2940
rect 110 2935 116 2936
rect 1830 2940 1836 2941
rect 1830 2936 1831 2940
rect 1835 2936 1836 2940
rect 3328 2938 3330 2944
rect 3335 2943 3336 2947
rect 3340 2946 3341 2947
rect 3394 2947 3400 2948
rect 3394 2946 3395 2947
rect 3340 2944 3395 2946
rect 3340 2943 3341 2944
rect 3335 2942 3341 2943
rect 3394 2943 3395 2944
rect 3399 2943 3400 2947
rect 3394 2942 3400 2943
rect 3402 2947 3408 2948
rect 3402 2943 3403 2947
rect 3407 2946 3408 2947
rect 3423 2947 3429 2948
rect 3423 2946 3424 2947
rect 3407 2944 3424 2946
rect 3407 2943 3408 2944
rect 3402 2942 3408 2943
rect 3423 2943 3424 2944
rect 3428 2943 3429 2947
rect 3423 2942 3429 2943
rect 3503 2947 3509 2948
rect 3503 2943 3504 2947
rect 3508 2946 3509 2947
rect 3518 2947 3524 2948
rect 3518 2946 3519 2947
rect 3508 2944 3519 2946
rect 3508 2943 3509 2944
rect 3503 2942 3509 2943
rect 3518 2943 3519 2944
rect 3523 2943 3524 2947
rect 3518 2942 3524 2943
rect 3362 2939 3368 2940
rect 3362 2938 3363 2939
rect 3328 2936 3363 2938
rect 1830 2935 1836 2936
rect 1894 2935 1901 2936
rect 522 2931 528 2932
rect 522 2927 523 2931
rect 527 2927 528 2931
rect 522 2926 528 2927
rect 530 2931 536 2932
rect 530 2927 531 2931
rect 535 2930 536 2931
rect 738 2931 744 2932
rect 535 2928 585 2930
rect 535 2927 536 2928
rect 530 2926 536 2927
rect 738 2927 739 2931
rect 743 2927 744 2931
rect 738 2926 744 2927
rect 858 2931 864 2932
rect 858 2927 859 2931
rect 863 2927 864 2931
rect 858 2926 864 2927
rect 950 2931 956 2932
rect 950 2927 951 2931
rect 955 2927 956 2931
rect 950 2926 956 2927
rect 1138 2931 1144 2932
rect 1138 2927 1139 2931
rect 1143 2927 1144 2931
rect 1138 2926 1144 2927
rect 1298 2931 1304 2932
rect 1298 2927 1299 2931
rect 1303 2927 1304 2931
rect 1298 2926 1304 2927
rect 1466 2931 1472 2932
rect 1466 2927 1467 2931
rect 1471 2927 1472 2931
rect 1466 2926 1472 2927
rect 1598 2931 1604 2932
rect 1598 2927 1599 2931
rect 1603 2927 1604 2931
rect 1894 2931 1895 2935
rect 1900 2931 1901 2935
rect 1894 2930 1901 2931
rect 2079 2935 2085 2936
rect 2079 2931 2080 2935
rect 2084 2934 2085 2935
rect 2094 2935 2100 2936
rect 2094 2934 2095 2935
rect 2084 2932 2095 2934
rect 2084 2931 2085 2932
rect 2079 2930 2085 2931
rect 2094 2931 2095 2932
rect 2099 2931 2100 2935
rect 2094 2930 2100 2931
rect 2138 2935 2144 2936
rect 2138 2931 2139 2935
rect 2143 2934 2144 2935
rect 2287 2935 2293 2936
rect 2287 2934 2288 2935
rect 2143 2932 2288 2934
rect 2143 2931 2144 2932
rect 2138 2930 2144 2931
rect 2287 2931 2288 2932
rect 2292 2931 2293 2935
rect 2287 2930 2293 2931
rect 2346 2935 2352 2936
rect 2346 2931 2347 2935
rect 2351 2934 2352 2935
rect 2479 2935 2485 2936
rect 2479 2934 2480 2935
rect 2351 2932 2480 2934
rect 2351 2931 2352 2932
rect 2346 2930 2352 2931
rect 2479 2931 2480 2932
rect 2484 2931 2485 2935
rect 2479 2930 2485 2931
rect 2663 2935 2669 2936
rect 2663 2931 2664 2935
rect 2668 2934 2669 2935
rect 2714 2935 2720 2936
rect 2714 2934 2715 2935
rect 2668 2932 2715 2934
rect 2668 2931 2669 2932
rect 2663 2930 2669 2931
rect 2714 2931 2715 2932
rect 2719 2931 2720 2935
rect 2714 2930 2720 2931
rect 2722 2935 2728 2936
rect 2722 2931 2723 2935
rect 2727 2934 2728 2935
rect 2831 2935 2837 2936
rect 2831 2934 2832 2935
rect 2727 2932 2832 2934
rect 2727 2931 2728 2932
rect 2722 2930 2728 2931
rect 2831 2931 2832 2932
rect 2836 2931 2837 2935
rect 2831 2930 2837 2931
rect 2910 2935 2916 2936
rect 2910 2931 2911 2935
rect 2915 2934 2916 2935
rect 2991 2935 2997 2936
rect 2991 2934 2992 2935
rect 2915 2932 2992 2934
rect 2915 2931 2916 2932
rect 2910 2930 2916 2931
rect 2991 2931 2992 2932
rect 2996 2931 2997 2935
rect 2991 2930 2997 2931
rect 3098 2935 3104 2936
rect 3098 2931 3099 2935
rect 3103 2934 3104 2935
rect 3143 2935 3149 2936
rect 3143 2934 3144 2935
rect 3103 2932 3144 2934
rect 3103 2931 3104 2932
rect 3098 2930 3104 2931
rect 3143 2931 3144 2932
rect 3148 2931 3149 2935
rect 3143 2930 3149 2931
rect 3202 2935 3208 2936
rect 3202 2931 3203 2935
rect 3207 2934 3208 2935
rect 3295 2935 3301 2936
rect 3295 2934 3296 2935
rect 3207 2932 3296 2934
rect 3207 2931 3208 2932
rect 3202 2930 3208 2931
rect 3295 2931 3296 2932
rect 3300 2931 3301 2935
rect 3362 2935 3363 2936
rect 3367 2935 3368 2939
rect 3362 2934 3368 2935
rect 3422 2935 3428 2936
rect 3295 2930 3301 2931
rect 3422 2931 3423 2935
rect 3427 2934 3428 2935
rect 3447 2935 3453 2936
rect 3447 2934 3448 2935
rect 3427 2932 3448 2934
rect 3427 2931 3428 2932
rect 3422 2930 3428 2931
rect 3447 2931 3448 2932
rect 3452 2931 3453 2935
rect 3447 2930 3453 2931
rect 1598 2926 1604 2927
rect 1902 2926 1908 2927
rect 110 2923 116 2924
rect 110 2919 111 2923
rect 115 2919 116 2923
rect 1830 2923 1836 2924
rect 110 2918 116 2919
rect 462 2920 468 2921
rect 462 2916 463 2920
rect 467 2916 468 2920
rect 462 2915 468 2916
rect 566 2920 572 2921
rect 566 2916 567 2920
rect 571 2916 572 2920
rect 566 2915 572 2916
rect 678 2920 684 2921
rect 678 2916 679 2920
rect 683 2916 684 2920
rect 678 2915 684 2916
rect 798 2920 804 2921
rect 798 2916 799 2920
rect 803 2916 804 2920
rect 798 2915 804 2916
rect 934 2920 940 2921
rect 934 2916 935 2920
rect 939 2916 940 2920
rect 934 2915 940 2916
rect 1078 2920 1084 2921
rect 1078 2916 1079 2920
rect 1083 2916 1084 2920
rect 1078 2915 1084 2916
rect 1238 2920 1244 2921
rect 1238 2916 1239 2920
rect 1243 2916 1244 2920
rect 1238 2915 1244 2916
rect 1406 2920 1412 2921
rect 1406 2916 1407 2920
rect 1411 2916 1412 2920
rect 1406 2915 1412 2916
rect 1582 2920 1588 2921
rect 1582 2916 1583 2920
rect 1587 2916 1588 2920
rect 1582 2915 1588 2916
rect 1742 2920 1748 2921
rect 1742 2916 1743 2920
rect 1747 2916 1748 2920
rect 1830 2919 1831 2923
rect 1835 2919 1836 2923
rect 1902 2922 1903 2926
rect 1907 2922 1908 2926
rect 1902 2921 1908 2922
rect 2086 2926 2092 2927
rect 2086 2922 2087 2926
rect 2091 2922 2092 2926
rect 2086 2921 2092 2922
rect 2294 2926 2300 2927
rect 2294 2922 2295 2926
rect 2299 2922 2300 2926
rect 2294 2921 2300 2922
rect 2486 2926 2492 2927
rect 2486 2922 2487 2926
rect 2491 2922 2492 2926
rect 2486 2921 2492 2922
rect 2670 2926 2676 2927
rect 2670 2922 2671 2926
rect 2675 2922 2676 2926
rect 2670 2921 2676 2922
rect 2838 2926 2844 2927
rect 2838 2922 2839 2926
rect 2843 2922 2844 2926
rect 2838 2921 2844 2922
rect 2998 2926 3004 2927
rect 2998 2922 2999 2926
rect 3003 2922 3004 2926
rect 2998 2921 3004 2922
rect 3150 2926 3156 2927
rect 3150 2922 3151 2926
rect 3155 2922 3156 2926
rect 3150 2921 3156 2922
rect 3302 2926 3308 2927
rect 3302 2922 3303 2926
rect 3307 2922 3308 2926
rect 3302 2921 3308 2922
rect 3454 2926 3460 2927
rect 3454 2922 3455 2926
rect 3459 2922 3460 2926
rect 3454 2921 3460 2922
rect 1830 2918 1836 2919
rect 1742 2915 1748 2916
rect 1870 2908 1876 2909
rect 1870 2904 1871 2908
rect 1875 2904 1876 2908
rect 1758 2903 1765 2904
rect 1870 2903 1876 2904
rect 3590 2908 3596 2909
rect 3590 2904 3591 2908
rect 3595 2904 3596 2908
rect 3590 2903 3596 2904
rect 1758 2899 1759 2903
rect 1764 2899 1765 2903
rect 1758 2898 1765 2899
rect 1798 2899 1804 2900
rect 1798 2895 1799 2899
rect 1803 2898 1804 2899
rect 2138 2899 2144 2900
rect 1803 2896 1913 2898
rect 1803 2895 1804 2896
rect 1798 2894 1804 2895
rect 2138 2895 2139 2899
rect 2143 2895 2144 2899
rect 2138 2894 2144 2895
rect 2346 2899 2352 2900
rect 2346 2895 2347 2899
rect 2351 2895 2352 2899
rect 2346 2894 2352 2895
rect 2494 2899 2500 2900
rect 2494 2895 2495 2899
rect 2499 2895 2500 2899
rect 2494 2894 2500 2895
rect 2722 2899 2728 2900
rect 2722 2895 2723 2899
rect 2727 2895 2728 2899
rect 2722 2894 2728 2895
rect 2878 2899 2884 2900
rect 2878 2895 2879 2899
rect 2883 2895 2884 2899
rect 3098 2899 3104 2900
rect 3098 2898 3099 2899
rect 3053 2896 3099 2898
rect 2878 2894 2884 2895
rect 3098 2895 3099 2896
rect 3103 2895 3104 2899
rect 3098 2894 3104 2895
rect 3202 2899 3208 2900
rect 3202 2895 3203 2899
rect 3207 2895 3208 2899
rect 3202 2894 3208 2895
rect 3310 2899 3316 2900
rect 3310 2895 3311 2899
rect 3315 2895 3316 2899
rect 3310 2894 3316 2895
rect 3362 2899 3368 2900
rect 3362 2895 3363 2899
rect 3367 2898 3368 2899
rect 3367 2896 3465 2898
rect 3367 2895 3368 2896
rect 3362 2894 3368 2895
rect 1870 2891 1876 2892
rect 1870 2887 1871 2891
rect 1875 2887 1876 2891
rect 3590 2891 3596 2892
rect 1870 2886 1876 2887
rect 1894 2888 1900 2889
rect 1894 2884 1895 2888
rect 1899 2884 1900 2888
rect 1894 2883 1900 2884
rect 2078 2888 2084 2889
rect 2078 2884 2079 2888
rect 2083 2884 2084 2888
rect 2078 2883 2084 2884
rect 2286 2888 2292 2889
rect 2286 2884 2287 2888
rect 2291 2884 2292 2888
rect 2286 2883 2292 2884
rect 2478 2888 2484 2889
rect 2478 2884 2479 2888
rect 2483 2884 2484 2888
rect 2478 2883 2484 2884
rect 2662 2888 2668 2889
rect 2662 2884 2663 2888
rect 2667 2884 2668 2888
rect 2662 2883 2668 2884
rect 2830 2888 2836 2889
rect 2830 2884 2831 2888
rect 2835 2884 2836 2888
rect 2830 2883 2836 2884
rect 2990 2888 2996 2889
rect 2990 2884 2991 2888
rect 2995 2884 2996 2888
rect 2990 2883 2996 2884
rect 3142 2888 3148 2889
rect 3142 2884 3143 2888
rect 3147 2884 3148 2888
rect 3142 2883 3148 2884
rect 3294 2888 3300 2889
rect 3294 2884 3295 2888
rect 3299 2884 3300 2888
rect 3294 2883 3300 2884
rect 3446 2888 3452 2889
rect 3446 2884 3447 2888
rect 3451 2884 3452 2888
rect 3590 2887 3591 2891
rect 3595 2887 3596 2891
rect 3590 2886 3596 2887
rect 3446 2883 3452 2884
rect 310 2876 316 2877
rect 110 2873 116 2874
rect 110 2869 111 2873
rect 115 2869 116 2873
rect 310 2872 311 2876
rect 315 2872 316 2876
rect 310 2871 316 2872
rect 430 2876 436 2877
rect 430 2872 431 2876
rect 435 2872 436 2876
rect 430 2871 436 2872
rect 550 2876 556 2877
rect 550 2872 551 2876
rect 555 2872 556 2876
rect 550 2871 556 2872
rect 678 2876 684 2877
rect 678 2872 679 2876
rect 683 2872 684 2876
rect 678 2871 684 2872
rect 814 2876 820 2877
rect 814 2872 815 2876
rect 819 2872 820 2876
rect 814 2871 820 2872
rect 950 2876 956 2877
rect 950 2872 951 2876
rect 955 2872 956 2876
rect 950 2871 956 2872
rect 1086 2876 1092 2877
rect 1086 2872 1087 2876
rect 1091 2872 1092 2876
rect 1086 2871 1092 2872
rect 1222 2876 1228 2877
rect 1222 2872 1223 2876
rect 1227 2872 1228 2876
rect 1222 2871 1228 2872
rect 1358 2876 1364 2877
rect 1358 2872 1359 2876
rect 1363 2872 1364 2876
rect 1358 2871 1364 2872
rect 1494 2876 1500 2877
rect 1494 2872 1495 2876
rect 1499 2872 1500 2876
rect 1494 2871 1500 2872
rect 1630 2876 1636 2877
rect 1630 2872 1631 2876
rect 1635 2872 1636 2876
rect 1630 2871 1636 2872
rect 1742 2876 1748 2877
rect 1742 2872 1743 2876
rect 1747 2872 1748 2876
rect 1742 2871 1748 2872
rect 1830 2873 1836 2874
rect 110 2868 116 2869
rect 1830 2869 1831 2873
rect 1835 2869 1836 2873
rect 1830 2868 1836 2869
rect 378 2867 384 2868
rect 378 2866 379 2867
rect 373 2864 379 2866
rect 378 2863 379 2864
rect 383 2863 384 2867
rect 671 2867 677 2868
rect 671 2866 672 2867
rect 432 2864 449 2866
rect 613 2864 672 2866
rect 378 2862 384 2863
rect 430 2863 436 2864
rect 430 2859 431 2863
rect 435 2859 436 2863
rect 671 2863 672 2864
rect 676 2863 677 2867
rect 754 2867 760 2868
rect 754 2866 755 2867
rect 741 2864 755 2866
rect 671 2862 677 2863
rect 754 2863 755 2864
rect 759 2863 760 2867
rect 754 2862 760 2863
rect 762 2867 768 2868
rect 762 2863 763 2867
rect 767 2866 768 2867
rect 1026 2867 1032 2868
rect 1026 2866 1027 2867
rect 767 2864 833 2866
rect 1013 2864 1027 2866
rect 767 2863 768 2864
rect 762 2862 768 2863
rect 1026 2863 1027 2864
rect 1031 2863 1032 2867
rect 1162 2867 1168 2868
rect 1162 2866 1163 2867
rect 1149 2864 1163 2866
rect 1026 2862 1032 2863
rect 1162 2863 1163 2864
rect 1167 2863 1168 2867
rect 1298 2867 1304 2868
rect 1298 2866 1299 2867
rect 1285 2864 1299 2866
rect 1162 2862 1168 2863
rect 1298 2863 1299 2864
rect 1303 2863 1304 2867
rect 1298 2862 1304 2863
rect 1306 2867 1312 2868
rect 1306 2863 1307 2867
rect 1311 2866 1312 2867
rect 1562 2867 1568 2868
rect 1311 2864 1377 2866
rect 1311 2863 1312 2864
rect 1306 2862 1312 2863
rect 1556 2860 1558 2865
rect 1562 2863 1563 2867
rect 1567 2866 1568 2867
rect 1698 2867 1704 2868
rect 1567 2864 1649 2866
rect 1567 2863 1568 2864
rect 1562 2862 1568 2863
rect 1698 2863 1699 2867
rect 1703 2866 1704 2867
rect 1703 2864 1761 2866
rect 1703 2863 1704 2864
rect 1698 2862 1704 2863
rect 430 2858 436 2859
rect 1554 2859 1560 2860
rect 110 2856 116 2857
rect 110 2852 111 2856
rect 115 2852 116 2856
rect 1554 2855 1555 2859
rect 1559 2855 1560 2859
rect 1554 2854 1560 2855
rect 1830 2856 1836 2857
rect 110 2851 116 2852
rect 1830 2852 1831 2856
rect 1835 2852 1836 2856
rect 1830 2851 1836 2852
rect 318 2838 324 2839
rect 318 2834 319 2838
rect 323 2834 324 2838
rect 318 2833 324 2834
rect 438 2838 444 2839
rect 438 2834 439 2838
rect 443 2834 444 2838
rect 438 2833 444 2834
rect 558 2838 564 2839
rect 558 2834 559 2838
rect 563 2834 564 2838
rect 558 2833 564 2834
rect 686 2838 692 2839
rect 686 2834 687 2838
rect 691 2834 692 2838
rect 686 2833 692 2834
rect 822 2838 828 2839
rect 822 2834 823 2838
rect 827 2834 828 2838
rect 822 2833 828 2834
rect 958 2838 964 2839
rect 958 2834 959 2838
rect 963 2834 964 2838
rect 958 2833 964 2834
rect 1094 2838 1100 2839
rect 1094 2834 1095 2838
rect 1099 2834 1100 2838
rect 1094 2833 1100 2834
rect 1230 2838 1236 2839
rect 1230 2834 1231 2838
rect 1235 2834 1236 2838
rect 1230 2833 1236 2834
rect 1366 2838 1372 2839
rect 1366 2834 1367 2838
rect 1371 2834 1372 2838
rect 1366 2833 1372 2834
rect 1502 2838 1508 2839
rect 1502 2834 1503 2838
rect 1507 2834 1508 2838
rect 1502 2833 1508 2834
rect 1638 2838 1644 2839
rect 1638 2834 1639 2838
rect 1643 2834 1644 2838
rect 1638 2833 1644 2834
rect 1750 2838 1756 2839
rect 1750 2834 1751 2838
rect 1755 2834 1756 2838
rect 2134 2836 2140 2837
rect 1750 2833 1756 2834
rect 1870 2833 1876 2834
rect 1870 2829 1871 2833
rect 1875 2829 1876 2833
rect 2134 2832 2135 2836
rect 2139 2832 2140 2836
rect 2134 2831 2140 2832
rect 2262 2836 2268 2837
rect 2262 2832 2263 2836
rect 2267 2832 2268 2836
rect 2262 2831 2268 2832
rect 2390 2836 2396 2837
rect 2390 2832 2391 2836
rect 2395 2832 2396 2836
rect 2390 2831 2396 2832
rect 2518 2836 2524 2837
rect 2518 2832 2519 2836
rect 2523 2832 2524 2836
rect 2518 2831 2524 2832
rect 2646 2836 2652 2837
rect 2646 2832 2647 2836
rect 2651 2832 2652 2836
rect 2646 2831 2652 2832
rect 2766 2836 2772 2837
rect 2766 2832 2767 2836
rect 2771 2832 2772 2836
rect 2766 2831 2772 2832
rect 2886 2836 2892 2837
rect 2886 2832 2887 2836
rect 2891 2832 2892 2836
rect 2886 2831 2892 2832
rect 3006 2836 3012 2837
rect 3006 2832 3007 2836
rect 3011 2832 3012 2836
rect 3006 2831 3012 2832
rect 3134 2836 3140 2837
rect 3134 2832 3135 2836
rect 3139 2832 3140 2836
rect 3134 2831 3140 2832
rect 3590 2833 3596 2834
rect 1870 2828 1876 2829
rect 3590 2829 3591 2833
rect 3595 2829 3596 2833
rect 3590 2828 3596 2829
rect 311 2827 317 2828
rect 311 2823 312 2827
rect 316 2826 317 2827
rect 326 2827 332 2828
rect 326 2826 327 2827
rect 316 2824 327 2826
rect 316 2823 317 2824
rect 311 2822 317 2823
rect 326 2823 327 2824
rect 331 2823 332 2827
rect 326 2822 332 2823
rect 378 2827 384 2828
rect 378 2823 379 2827
rect 383 2826 384 2827
rect 431 2827 437 2828
rect 431 2826 432 2827
rect 383 2824 432 2826
rect 383 2823 384 2824
rect 378 2822 384 2823
rect 431 2823 432 2824
rect 436 2823 437 2827
rect 431 2822 437 2823
rect 522 2827 528 2828
rect 522 2823 523 2827
rect 527 2826 528 2827
rect 551 2827 557 2828
rect 551 2826 552 2827
rect 527 2824 552 2826
rect 527 2823 528 2824
rect 522 2822 528 2823
rect 551 2823 552 2824
rect 556 2823 557 2827
rect 551 2822 557 2823
rect 671 2827 677 2828
rect 671 2823 672 2827
rect 676 2826 677 2827
rect 679 2827 685 2828
rect 679 2826 680 2827
rect 676 2824 680 2826
rect 676 2823 677 2824
rect 671 2822 677 2823
rect 679 2823 680 2824
rect 684 2823 685 2827
rect 679 2822 685 2823
rect 754 2827 760 2828
rect 754 2823 755 2827
rect 759 2826 760 2827
rect 815 2827 821 2828
rect 815 2826 816 2827
rect 759 2824 816 2826
rect 759 2823 760 2824
rect 754 2822 760 2823
rect 815 2823 816 2824
rect 820 2823 821 2827
rect 815 2822 821 2823
rect 951 2827 957 2828
rect 951 2823 952 2827
rect 956 2826 957 2827
rect 966 2827 972 2828
rect 966 2826 967 2827
rect 956 2824 967 2826
rect 956 2823 957 2824
rect 951 2822 957 2823
rect 966 2823 967 2824
rect 971 2823 972 2827
rect 966 2822 972 2823
rect 1026 2827 1032 2828
rect 1026 2823 1027 2827
rect 1031 2826 1032 2827
rect 1087 2827 1093 2828
rect 1087 2826 1088 2827
rect 1031 2824 1088 2826
rect 1031 2823 1032 2824
rect 1026 2822 1032 2823
rect 1087 2823 1088 2824
rect 1092 2823 1093 2827
rect 1087 2822 1093 2823
rect 1162 2827 1168 2828
rect 1162 2823 1163 2827
rect 1167 2826 1168 2827
rect 1223 2827 1229 2828
rect 1223 2826 1224 2827
rect 1167 2824 1224 2826
rect 1167 2823 1168 2824
rect 1162 2822 1168 2823
rect 1223 2823 1224 2824
rect 1228 2823 1229 2827
rect 1223 2822 1229 2823
rect 1298 2827 1304 2828
rect 1298 2823 1299 2827
rect 1303 2826 1304 2827
rect 1359 2827 1365 2828
rect 1359 2826 1360 2827
rect 1303 2824 1360 2826
rect 1303 2823 1304 2824
rect 1298 2822 1304 2823
rect 1359 2823 1360 2824
rect 1364 2823 1365 2827
rect 1359 2822 1365 2823
rect 1495 2827 1501 2828
rect 1495 2823 1496 2827
rect 1500 2826 1501 2827
rect 1562 2827 1568 2828
rect 1562 2826 1563 2827
rect 1500 2824 1563 2826
rect 1500 2823 1501 2824
rect 1495 2822 1501 2823
rect 1562 2823 1563 2824
rect 1567 2823 1568 2827
rect 1562 2822 1568 2823
rect 1631 2827 1637 2828
rect 1631 2823 1632 2827
rect 1636 2826 1637 2827
rect 1698 2827 1704 2828
rect 1698 2826 1699 2827
rect 1636 2824 1699 2826
rect 1636 2823 1637 2824
rect 1631 2822 1637 2823
rect 1698 2823 1699 2824
rect 1703 2823 1704 2827
rect 1698 2822 1704 2823
rect 1743 2827 1749 2828
rect 1743 2823 1744 2827
rect 1748 2826 1749 2827
rect 1758 2827 1764 2828
rect 1758 2826 1759 2827
rect 1748 2824 1759 2826
rect 1748 2823 1749 2824
rect 1743 2822 1749 2823
rect 1758 2823 1759 2824
rect 1763 2823 1764 2827
rect 1758 2822 1764 2823
rect 2094 2827 2100 2828
rect 2094 2823 2095 2827
rect 2099 2826 2100 2827
rect 2202 2827 2208 2828
rect 2099 2824 2153 2826
rect 2099 2823 2100 2824
rect 2094 2822 2100 2823
rect 2202 2823 2203 2827
rect 2207 2826 2208 2827
rect 2351 2827 2357 2828
rect 2207 2824 2281 2826
rect 2207 2823 2208 2824
rect 2202 2822 2208 2823
rect 2351 2823 2352 2827
rect 2356 2826 2357 2827
rect 2463 2827 2469 2828
rect 2356 2824 2409 2826
rect 2356 2823 2357 2824
rect 2351 2822 2357 2823
rect 2463 2823 2464 2827
rect 2468 2826 2469 2827
rect 2714 2827 2720 2828
rect 2714 2826 2715 2827
rect 2468 2824 2537 2826
rect 2709 2824 2715 2826
rect 2468 2823 2469 2824
rect 2463 2822 2469 2823
rect 2714 2823 2715 2824
rect 2719 2823 2720 2827
rect 2954 2827 2960 2828
rect 2954 2826 2955 2827
rect 2714 2822 2720 2823
rect 2828 2820 2830 2825
rect 2949 2824 2955 2826
rect 2954 2823 2955 2824
rect 2959 2823 2960 2827
rect 3078 2827 3084 2828
rect 3078 2826 3079 2827
rect 3069 2824 3079 2826
rect 2954 2822 2960 2823
rect 3078 2823 3079 2824
rect 3083 2823 3084 2827
rect 3078 2822 3084 2823
rect 3086 2827 3092 2828
rect 3086 2823 3087 2827
rect 3091 2826 3092 2827
rect 3091 2824 3153 2826
rect 3091 2823 3092 2824
rect 3086 2822 3092 2823
rect 2826 2819 2832 2820
rect 1870 2816 1876 2817
rect 159 2815 165 2816
rect 159 2811 160 2815
rect 164 2814 165 2815
rect 210 2815 216 2816
rect 210 2814 211 2815
rect 164 2812 211 2814
rect 164 2811 165 2812
rect 159 2810 165 2811
rect 210 2811 211 2812
rect 215 2811 216 2815
rect 210 2810 216 2811
rect 218 2815 224 2816
rect 218 2811 219 2815
rect 223 2814 224 2815
rect 295 2815 301 2816
rect 295 2814 296 2815
rect 223 2812 296 2814
rect 223 2811 224 2812
rect 218 2810 224 2811
rect 295 2811 296 2812
rect 300 2811 301 2815
rect 295 2810 301 2811
rect 430 2815 436 2816
rect 430 2811 431 2815
rect 435 2814 436 2815
rect 439 2815 445 2816
rect 439 2814 440 2815
rect 435 2812 440 2814
rect 435 2811 436 2812
rect 430 2810 436 2811
rect 439 2811 440 2812
rect 444 2811 445 2815
rect 439 2810 445 2811
rect 498 2815 504 2816
rect 498 2811 499 2815
rect 503 2814 504 2815
rect 599 2815 605 2816
rect 599 2814 600 2815
rect 503 2812 600 2814
rect 503 2811 504 2812
rect 498 2810 504 2811
rect 599 2811 600 2812
rect 604 2811 605 2815
rect 599 2810 605 2811
rect 658 2815 664 2816
rect 658 2811 659 2815
rect 663 2814 664 2815
rect 775 2815 781 2816
rect 775 2814 776 2815
rect 663 2812 776 2814
rect 663 2811 664 2812
rect 658 2810 664 2811
rect 775 2811 776 2812
rect 780 2811 781 2815
rect 775 2810 781 2811
rect 951 2815 957 2816
rect 951 2811 952 2815
rect 956 2814 957 2815
rect 1018 2815 1024 2816
rect 1018 2814 1019 2815
rect 956 2812 1019 2814
rect 956 2811 957 2812
rect 951 2810 957 2811
rect 1018 2811 1019 2812
rect 1023 2811 1024 2815
rect 1018 2810 1024 2811
rect 1135 2815 1141 2816
rect 1135 2811 1136 2815
rect 1140 2814 1141 2815
rect 1202 2815 1208 2816
rect 1202 2814 1203 2815
rect 1140 2812 1203 2814
rect 1140 2811 1141 2812
rect 1135 2810 1141 2811
rect 1202 2811 1203 2812
rect 1207 2811 1208 2815
rect 1202 2810 1208 2811
rect 1266 2815 1272 2816
rect 1266 2811 1267 2815
rect 1271 2814 1272 2815
rect 1327 2815 1333 2816
rect 1327 2814 1328 2815
rect 1271 2812 1328 2814
rect 1271 2811 1272 2812
rect 1266 2810 1272 2811
rect 1327 2811 1328 2812
rect 1332 2811 1333 2815
rect 1327 2810 1333 2811
rect 1527 2815 1533 2816
rect 1527 2811 1528 2815
rect 1532 2814 1533 2815
rect 1554 2815 1560 2816
rect 1554 2814 1555 2815
rect 1532 2812 1555 2814
rect 1532 2811 1533 2812
rect 1527 2810 1533 2811
rect 1554 2811 1555 2812
rect 1559 2811 1560 2815
rect 1554 2810 1560 2811
rect 1586 2815 1592 2816
rect 1586 2811 1587 2815
rect 1591 2814 1592 2815
rect 1727 2815 1733 2816
rect 1727 2814 1728 2815
rect 1591 2812 1728 2814
rect 1591 2811 1592 2812
rect 1586 2810 1592 2811
rect 1727 2811 1728 2812
rect 1732 2811 1733 2815
rect 1870 2812 1871 2816
rect 1875 2812 1876 2816
rect 2826 2815 2827 2819
rect 2831 2815 2832 2819
rect 2826 2814 2832 2815
rect 3590 2816 3596 2817
rect 1870 2811 1876 2812
rect 3590 2812 3591 2816
rect 3595 2812 3596 2816
rect 3590 2811 3596 2812
rect 1727 2810 1733 2811
rect 166 2806 172 2807
rect 166 2802 167 2806
rect 171 2802 172 2806
rect 166 2801 172 2802
rect 302 2806 308 2807
rect 302 2802 303 2806
rect 307 2802 308 2806
rect 302 2801 308 2802
rect 446 2806 452 2807
rect 446 2802 447 2806
rect 451 2802 452 2806
rect 446 2801 452 2802
rect 606 2806 612 2807
rect 606 2802 607 2806
rect 611 2802 612 2806
rect 606 2801 612 2802
rect 782 2806 788 2807
rect 782 2802 783 2806
rect 787 2802 788 2806
rect 782 2801 788 2802
rect 958 2806 964 2807
rect 958 2802 959 2806
rect 963 2802 964 2806
rect 958 2801 964 2802
rect 1142 2806 1148 2807
rect 1142 2802 1143 2806
rect 1147 2802 1148 2806
rect 1142 2801 1148 2802
rect 1334 2806 1340 2807
rect 1334 2802 1335 2806
rect 1339 2802 1340 2806
rect 1334 2801 1340 2802
rect 1534 2806 1540 2807
rect 1534 2802 1535 2806
rect 1539 2802 1540 2806
rect 1534 2801 1540 2802
rect 1734 2806 1740 2807
rect 1734 2802 1735 2806
rect 1739 2802 1740 2806
rect 1734 2801 1740 2802
rect 2142 2798 2148 2799
rect 2142 2794 2143 2798
rect 2147 2794 2148 2798
rect 2142 2793 2148 2794
rect 2270 2798 2276 2799
rect 2270 2794 2271 2798
rect 2275 2794 2276 2798
rect 2270 2793 2276 2794
rect 2398 2798 2404 2799
rect 2398 2794 2399 2798
rect 2403 2794 2404 2798
rect 2398 2793 2404 2794
rect 2526 2798 2532 2799
rect 2526 2794 2527 2798
rect 2531 2794 2532 2798
rect 2526 2793 2532 2794
rect 2654 2798 2660 2799
rect 2654 2794 2655 2798
rect 2659 2794 2660 2798
rect 2654 2793 2660 2794
rect 2774 2798 2780 2799
rect 2774 2794 2775 2798
rect 2779 2794 2780 2798
rect 2774 2793 2780 2794
rect 2894 2798 2900 2799
rect 2894 2794 2895 2798
rect 2899 2794 2900 2798
rect 2894 2793 2900 2794
rect 3014 2798 3020 2799
rect 3014 2794 3015 2798
rect 3019 2794 3020 2798
rect 3014 2793 3020 2794
rect 3142 2798 3148 2799
rect 3142 2794 3143 2798
rect 3147 2794 3148 2798
rect 3142 2793 3148 2794
rect 110 2788 116 2789
rect 110 2784 111 2788
rect 115 2784 116 2788
rect 110 2783 116 2784
rect 1830 2788 1836 2789
rect 1830 2784 1831 2788
rect 1835 2784 1836 2788
rect 1830 2783 1836 2784
rect 2135 2787 2141 2788
rect 2135 2783 2136 2787
rect 2140 2786 2141 2787
rect 2202 2787 2208 2788
rect 2202 2786 2203 2787
rect 2140 2784 2203 2786
rect 2140 2783 2141 2784
rect 2135 2782 2141 2783
rect 2202 2783 2203 2784
rect 2207 2783 2208 2787
rect 2202 2782 2208 2783
rect 2263 2787 2269 2788
rect 2263 2783 2264 2787
rect 2268 2786 2269 2787
rect 2351 2787 2357 2788
rect 2351 2786 2352 2787
rect 2268 2784 2352 2786
rect 2268 2783 2269 2784
rect 2263 2782 2269 2783
rect 2351 2783 2352 2784
rect 2356 2783 2357 2787
rect 2351 2782 2357 2783
rect 2391 2787 2397 2788
rect 2391 2783 2392 2787
rect 2396 2786 2397 2787
rect 2463 2787 2469 2788
rect 2463 2786 2464 2787
rect 2396 2784 2464 2786
rect 2396 2783 2397 2784
rect 2391 2782 2397 2783
rect 2463 2783 2464 2784
rect 2468 2783 2469 2787
rect 2463 2782 2469 2783
rect 2519 2787 2525 2788
rect 2519 2783 2520 2787
rect 2524 2786 2525 2787
rect 2558 2787 2564 2788
rect 2558 2786 2559 2787
rect 2524 2784 2559 2786
rect 2524 2783 2525 2784
rect 2519 2782 2525 2783
rect 2558 2783 2559 2784
rect 2563 2783 2564 2787
rect 2558 2782 2564 2783
rect 2647 2787 2653 2788
rect 2647 2783 2648 2787
rect 2652 2786 2653 2787
rect 2662 2787 2668 2788
rect 2662 2786 2663 2787
rect 2652 2784 2663 2786
rect 2652 2783 2653 2784
rect 2647 2782 2653 2783
rect 2662 2783 2663 2784
rect 2667 2783 2668 2787
rect 2662 2782 2668 2783
rect 2714 2787 2720 2788
rect 2714 2783 2715 2787
rect 2719 2786 2720 2787
rect 2767 2787 2773 2788
rect 2767 2786 2768 2787
rect 2719 2784 2768 2786
rect 2719 2783 2720 2784
rect 2714 2782 2720 2783
rect 2767 2783 2768 2784
rect 2772 2783 2773 2787
rect 2767 2782 2773 2783
rect 2878 2787 2884 2788
rect 2878 2783 2879 2787
rect 2883 2786 2884 2787
rect 2887 2787 2893 2788
rect 2887 2786 2888 2787
rect 2883 2784 2888 2786
rect 2883 2783 2884 2784
rect 2878 2782 2884 2783
rect 2887 2783 2888 2784
rect 2892 2783 2893 2787
rect 2887 2782 2893 2783
rect 2954 2787 2960 2788
rect 2954 2783 2955 2787
rect 2959 2786 2960 2787
rect 3007 2787 3013 2788
rect 3007 2786 3008 2787
rect 2959 2784 3008 2786
rect 2959 2783 2960 2784
rect 2954 2782 2960 2783
rect 3007 2783 3008 2784
rect 3012 2783 3013 2787
rect 3007 2782 3013 2783
rect 3078 2787 3084 2788
rect 3078 2783 3079 2787
rect 3083 2786 3084 2787
rect 3135 2787 3141 2788
rect 3135 2786 3136 2787
rect 3083 2784 3136 2786
rect 3083 2783 3084 2784
rect 3078 2782 3084 2783
rect 3135 2783 3136 2784
rect 3140 2783 3141 2787
rect 3135 2782 3141 2783
rect 218 2779 224 2780
rect 218 2775 219 2779
rect 223 2775 224 2779
rect 218 2774 224 2775
rect 354 2779 360 2780
rect 354 2775 355 2779
rect 359 2775 360 2779
rect 354 2774 360 2775
rect 498 2779 504 2780
rect 498 2775 499 2779
rect 503 2775 504 2779
rect 498 2774 504 2775
rect 658 2779 664 2780
rect 658 2775 659 2779
rect 663 2775 664 2779
rect 658 2774 664 2775
rect 966 2779 972 2780
rect 966 2775 967 2779
rect 971 2775 972 2779
rect 966 2774 972 2775
rect 1018 2779 1024 2780
rect 1018 2775 1019 2779
rect 1023 2778 1024 2779
rect 1202 2779 1208 2780
rect 1023 2776 1153 2778
rect 1023 2775 1024 2776
rect 1018 2774 1024 2775
rect 1202 2775 1203 2779
rect 1207 2778 1208 2779
rect 1586 2779 1592 2780
rect 1207 2776 1345 2778
rect 1207 2775 1208 2776
rect 1202 2774 1208 2775
rect 1586 2775 1587 2779
rect 1591 2775 1592 2779
rect 1586 2774 1592 2775
rect 110 2771 116 2772
rect 110 2767 111 2771
rect 115 2767 116 2771
rect 1830 2771 1836 2772
rect 110 2766 116 2767
rect 158 2768 164 2769
rect 158 2764 159 2768
rect 163 2764 164 2768
rect 158 2763 164 2764
rect 294 2768 300 2769
rect 294 2764 295 2768
rect 299 2764 300 2768
rect 294 2763 300 2764
rect 438 2768 444 2769
rect 438 2764 439 2768
rect 443 2764 444 2768
rect 438 2763 444 2764
rect 598 2768 604 2769
rect 598 2764 599 2768
rect 603 2764 604 2768
rect 598 2763 604 2764
rect 774 2768 780 2769
rect 774 2764 775 2768
rect 779 2764 780 2768
rect 774 2763 780 2764
rect 950 2768 956 2769
rect 950 2764 951 2768
rect 955 2764 956 2768
rect 950 2763 956 2764
rect 1134 2768 1140 2769
rect 1134 2764 1135 2768
rect 1139 2764 1140 2768
rect 1134 2763 1140 2764
rect 1326 2768 1332 2769
rect 1326 2764 1327 2768
rect 1331 2764 1332 2768
rect 1326 2763 1332 2764
rect 1526 2768 1532 2769
rect 1526 2764 1527 2768
rect 1531 2764 1532 2768
rect 1526 2763 1532 2764
rect 1726 2768 1732 2769
rect 1726 2764 1727 2768
rect 1731 2764 1732 2768
rect 1830 2767 1831 2771
rect 1835 2767 1836 2771
rect 1830 2766 1836 2767
rect 2215 2767 2221 2768
rect 1726 2763 1732 2764
rect 2215 2763 2216 2767
rect 2220 2766 2221 2767
rect 2223 2767 2229 2768
rect 2223 2766 2224 2767
rect 2220 2764 2224 2766
rect 2220 2763 2221 2764
rect 2215 2762 2221 2763
rect 2223 2763 2224 2764
rect 2228 2763 2229 2767
rect 2223 2762 2229 2763
rect 2282 2767 2288 2768
rect 2282 2763 2283 2767
rect 2287 2766 2288 2767
rect 2303 2767 2309 2768
rect 2303 2766 2304 2767
rect 2287 2764 2304 2766
rect 2287 2763 2288 2764
rect 2282 2762 2288 2763
rect 2303 2763 2304 2764
rect 2308 2763 2309 2767
rect 2303 2762 2309 2763
rect 2362 2767 2368 2768
rect 2362 2763 2363 2767
rect 2367 2766 2368 2767
rect 2383 2767 2389 2768
rect 2383 2766 2384 2767
rect 2367 2764 2384 2766
rect 2367 2763 2368 2764
rect 2362 2762 2368 2763
rect 2383 2763 2384 2764
rect 2388 2763 2389 2767
rect 2383 2762 2389 2763
rect 2442 2767 2448 2768
rect 2442 2763 2443 2767
rect 2447 2766 2448 2767
rect 2463 2767 2469 2768
rect 2463 2766 2464 2767
rect 2447 2764 2464 2766
rect 2447 2763 2448 2764
rect 2442 2762 2448 2763
rect 2463 2763 2464 2764
rect 2468 2763 2469 2767
rect 2463 2762 2469 2763
rect 2542 2767 2549 2768
rect 2542 2763 2543 2767
rect 2548 2763 2549 2767
rect 2542 2762 2549 2763
rect 2631 2767 2637 2768
rect 2631 2763 2632 2767
rect 2636 2766 2637 2767
rect 2646 2767 2652 2768
rect 2646 2766 2647 2767
rect 2636 2764 2647 2766
rect 2636 2763 2637 2764
rect 2631 2762 2637 2763
rect 2646 2763 2647 2764
rect 2651 2763 2652 2767
rect 2646 2762 2652 2763
rect 2690 2767 2696 2768
rect 2690 2763 2691 2767
rect 2695 2766 2696 2767
rect 2719 2767 2725 2768
rect 2719 2766 2720 2767
rect 2695 2764 2720 2766
rect 2695 2763 2696 2764
rect 2690 2762 2696 2763
rect 2719 2763 2720 2764
rect 2724 2763 2725 2767
rect 2719 2762 2725 2763
rect 2807 2767 2813 2768
rect 2807 2763 2808 2767
rect 2812 2766 2813 2767
rect 2826 2767 2832 2768
rect 2826 2766 2827 2767
rect 2812 2764 2827 2766
rect 2812 2763 2813 2764
rect 2807 2762 2813 2763
rect 2826 2763 2827 2764
rect 2831 2763 2832 2767
rect 2826 2762 2832 2763
rect 2866 2767 2872 2768
rect 2866 2763 2867 2767
rect 2871 2766 2872 2767
rect 2895 2767 2901 2768
rect 2895 2766 2896 2767
rect 2871 2764 2896 2766
rect 2871 2763 2872 2764
rect 2866 2762 2872 2763
rect 2895 2763 2896 2764
rect 2900 2763 2901 2767
rect 2895 2762 2901 2763
rect 2954 2767 2960 2768
rect 2954 2763 2955 2767
rect 2959 2766 2960 2767
rect 2983 2767 2989 2768
rect 2983 2766 2984 2767
rect 2959 2764 2984 2766
rect 2959 2763 2960 2764
rect 2954 2762 2960 2763
rect 2983 2763 2984 2764
rect 2988 2763 2989 2767
rect 2983 2762 2989 2763
rect 2230 2758 2236 2759
rect 2230 2754 2231 2758
rect 2235 2754 2236 2758
rect 2230 2753 2236 2754
rect 2310 2758 2316 2759
rect 2310 2754 2311 2758
rect 2315 2754 2316 2758
rect 2310 2753 2316 2754
rect 2390 2758 2396 2759
rect 2390 2754 2391 2758
rect 2395 2754 2396 2758
rect 2390 2753 2396 2754
rect 2470 2758 2476 2759
rect 2470 2754 2471 2758
rect 2475 2754 2476 2758
rect 2470 2753 2476 2754
rect 2550 2758 2556 2759
rect 2550 2754 2551 2758
rect 2555 2754 2556 2758
rect 2550 2753 2556 2754
rect 2638 2758 2644 2759
rect 2638 2754 2639 2758
rect 2643 2754 2644 2758
rect 2638 2753 2644 2754
rect 2726 2758 2732 2759
rect 2726 2754 2727 2758
rect 2731 2754 2732 2758
rect 2726 2753 2732 2754
rect 2814 2758 2820 2759
rect 2814 2754 2815 2758
rect 2819 2754 2820 2758
rect 2814 2753 2820 2754
rect 2902 2758 2908 2759
rect 2902 2754 2903 2758
rect 2907 2754 2908 2758
rect 2902 2753 2908 2754
rect 2990 2758 2996 2759
rect 2990 2754 2991 2758
rect 2995 2754 2996 2758
rect 2990 2753 2996 2754
rect 210 2751 216 2752
rect 210 2747 211 2751
rect 215 2750 216 2751
rect 791 2751 797 2752
rect 791 2750 792 2751
rect 215 2748 792 2750
rect 215 2747 216 2748
rect 210 2746 216 2747
rect 791 2747 792 2748
rect 796 2747 797 2751
rect 791 2746 797 2747
rect 1702 2751 1708 2752
rect 1702 2747 1703 2751
rect 1707 2750 1708 2751
rect 1743 2751 1749 2752
rect 1743 2750 1744 2751
rect 1707 2748 1744 2750
rect 1707 2747 1708 2748
rect 1702 2746 1708 2747
rect 1743 2747 1744 2748
rect 1748 2747 1749 2751
rect 1743 2746 1749 2747
rect 1870 2740 1876 2741
rect 1870 2736 1871 2740
rect 1875 2736 1876 2740
rect 1870 2735 1876 2736
rect 3590 2740 3596 2741
rect 3590 2736 3591 2740
rect 3595 2736 3596 2740
rect 3590 2735 3596 2736
rect 2282 2731 2288 2732
rect 2282 2727 2283 2731
rect 2287 2727 2288 2731
rect 2282 2726 2288 2727
rect 2362 2731 2368 2732
rect 2362 2727 2363 2731
rect 2367 2727 2368 2731
rect 2362 2726 2368 2727
rect 2442 2731 2448 2732
rect 2442 2727 2443 2731
rect 2447 2727 2448 2731
rect 2542 2731 2548 2732
rect 2542 2730 2543 2731
rect 2525 2728 2543 2730
rect 2442 2726 2448 2727
rect 2542 2727 2543 2728
rect 2547 2727 2548 2731
rect 2542 2726 2548 2727
rect 2558 2731 2564 2732
rect 2558 2727 2559 2731
rect 2563 2727 2564 2731
rect 2558 2726 2564 2727
rect 2690 2731 2696 2732
rect 2690 2727 2691 2731
rect 2695 2727 2696 2731
rect 2690 2726 2696 2727
rect 2778 2731 2784 2732
rect 2778 2727 2779 2731
rect 2783 2727 2784 2731
rect 2778 2726 2784 2727
rect 2866 2731 2872 2732
rect 2866 2727 2867 2731
rect 2871 2727 2872 2731
rect 2866 2726 2872 2727
rect 2954 2731 2960 2732
rect 2954 2727 2955 2731
rect 2959 2727 2960 2731
rect 2954 2726 2960 2727
rect 2998 2731 3004 2732
rect 2998 2727 2999 2731
rect 3003 2727 3004 2731
rect 2998 2726 3004 2727
rect 1870 2723 1876 2724
rect 134 2720 140 2721
rect 110 2717 116 2718
rect 110 2713 111 2717
rect 115 2713 116 2717
rect 134 2716 135 2720
rect 139 2716 140 2720
rect 134 2715 140 2716
rect 246 2720 252 2721
rect 246 2716 247 2720
rect 251 2716 252 2720
rect 246 2715 252 2716
rect 390 2720 396 2721
rect 390 2716 391 2720
rect 395 2716 396 2720
rect 390 2715 396 2716
rect 550 2720 556 2721
rect 550 2716 551 2720
rect 555 2716 556 2720
rect 550 2715 556 2716
rect 710 2720 716 2721
rect 710 2716 711 2720
rect 715 2716 716 2720
rect 710 2715 716 2716
rect 878 2720 884 2721
rect 878 2716 879 2720
rect 883 2716 884 2720
rect 878 2715 884 2716
rect 1038 2720 1044 2721
rect 1038 2716 1039 2720
rect 1043 2716 1044 2720
rect 1038 2715 1044 2716
rect 1198 2720 1204 2721
rect 1198 2716 1199 2720
rect 1203 2716 1204 2720
rect 1198 2715 1204 2716
rect 1358 2720 1364 2721
rect 1358 2716 1359 2720
rect 1363 2716 1364 2720
rect 1358 2715 1364 2716
rect 1518 2720 1524 2721
rect 1518 2716 1519 2720
rect 1523 2716 1524 2720
rect 1518 2715 1524 2716
rect 1686 2720 1692 2721
rect 1686 2716 1687 2720
rect 1691 2716 1692 2720
rect 1870 2719 1871 2723
rect 1875 2719 1876 2723
rect 3590 2723 3596 2724
rect 1870 2718 1876 2719
rect 2222 2720 2228 2721
rect 1686 2715 1692 2716
rect 1830 2717 1836 2718
rect 110 2712 116 2713
rect 1830 2713 1831 2717
rect 1835 2713 1836 2717
rect 2222 2716 2223 2720
rect 2227 2716 2228 2720
rect 2222 2715 2228 2716
rect 2302 2720 2308 2721
rect 2302 2716 2303 2720
rect 2307 2716 2308 2720
rect 2302 2715 2308 2716
rect 2382 2720 2388 2721
rect 2382 2716 2383 2720
rect 2387 2716 2388 2720
rect 2382 2715 2388 2716
rect 2462 2720 2468 2721
rect 2462 2716 2463 2720
rect 2467 2716 2468 2720
rect 2462 2715 2468 2716
rect 2542 2720 2548 2721
rect 2542 2716 2543 2720
rect 2547 2716 2548 2720
rect 2542 2715 2548 2716
rect 2630 2720 2636 2721
rect 2630 2716 2631 2720
rect 2635 2716 2636 2720
rect 2630 2715 2636 2716
rect 2718 2720 2724 2721
rect 2718 2716 2719 2720
rect 2723 2716 2724 2720
rect 2718 2715 2724 2716
rect 2806 2720 2812 2721
rect 2806 2716 2807 2720
rect 2811 2716 2812 2720
rect 2806 2715 2812 2716
rect 2894 2720 2900 2721
rect 2894 2716 2895 2720
rect 2899 2716 2900 2720
rect 2894 2715 2900 2716
rect 2982 2720 2988 2721
rect 2982 2716 2983 2720
rect 2987 2716 2988 2720
rect 3590 2719 3591 2723
rect 3595 2719 3596 2723
rect 3590 2718 3596 2719
rect 2982 2715 2988 2716
rect 1830 2712 1836 2713
rect 202 2711 208 2712
rect 136 2708 153 2710
rect 134 2707 140 2708
rect 134 2703 135 2707
rect 139 2703 140 2707
rect 202 2707 203 2711
rect 207 2710 208 2711
rect 478 2711 484 2712
rect 478 2710 479 2711
rect 207 2708 265 2710
rect 453 2708 479 2710
rect 207 2707 208 2708
rect 202 2706 208 2707
rect 478 2707 479 2708
rect 483 2707 484 2711
rect 703 2711 709 2712
rect 703 2710 704 2711
rect 613 2708 704 2710
rect 478 2706 484 2707
rect 703 2707 704 2708
rect 708 2707 709 2711
rect 962 2711 968 2712
rect 962 2710 963 2711
rect 703 2706 709 2707
rect 134 2702 140 2703
rect 650 2703 656 2704
rect 110 2700 116 2701
rect 110 2696 111 2700
rect 115 2696 116 2700
rect 650 2699 651 2703
rect 655 2702 656 2703
rect 728 2702 730 2709
rect 941 2708 963 2710
rect 962 2707 963 2708
rect 967 2707 968 2711
rect 1110 2711 1116 2712
rect 1110 2710 1111 2711
rect 1101 2708 1111 2710
rect 962 2706 968 2707
rect 1110 2707 1111 2708
rect 1115 2707 1116 2711
rect 1266 2711 1272 2712
rect 1266 2710 1267 2711
rect 1261 2708 1267 2710
rect 1110 2706 1116 2707
rect 1266 2707 1267 2708
rect 1271 2707 1272 2711
rect 1426 2711 1432 2712
rect 1360 2708 1377 2710
rect 1266 2706 1272 2707
rect 1358 2707 1364 2708
rect 1358 2703 1359 2707
rect 1363 2703 1364 2707
rect 1426 2707 1427 2711
rect 1431 2710 1432 2711
rect 1586 2711 1592 2712
rect 1431 2708 1537 2710
rect 1431 2707 1432 2708
rect 1426 2706 1432 2707
rect 1586 2707 1587 2711
rect 1591 2710 1592 2711
rect 1591 2708 1705 2710
rect 1591 2707 1592 2708
rect 1586 2706 1592 2707
rect 1358 2702 1364 2703
rect 655 2700 730 2702
rect 1830 2700 1836 2701
rect 655 2699 656 2700
rect 650 2698 656 2699
rect 110 2695 116 2696
rect 1830 2696 1831 2700
rect 1835 2696 1836 2700
rect 1830 2695 1836 2696
rect 142 2682 148 2683
rect 142 2678 143 2682
rect 147 2678 148 2682
rect 142 2677 148 2678
rect 254 2682 260 2683
rect 254 2678 255 2682
rect 259 2678 260 2682
rect 254 2677 260 2678
rect 398 2682 404 2683
rect 398 2678 399 2682
rect 403 2678 404 2682
rect 398 2677 404 2678
rect 558 2682 564 2683
rect 558 2678 559 2682
rect 563 2678 564 2682
rect 558 2677 564 2678
rect 718 2682 724 2683
rect 718 2678 719 2682
rect 723 2678 724 2682
rect 718 2677 724 2678
rect 886 2682 892 2683
rect 886 2678 887 2682
rect 891 2678 892 2682
rect 886 2677 892 2678
rect 1046 2682 1052 2683
rect 1046 2678 1047 2682
rect 1051 2678 1052 2682
rect 1046 2677 1052 2678
rect 1206 2682 1212 2683
rect 1206 2678 1207 2682
rect 1211 2678 1212 2682
rect 1206 2677 1212 2678
rect 1366 2682 1372 2683
rect 1366 2678 1367 2682
rect 1371 2678 1372 2682
rect 1366 2677 1372 2678
rect 1526 2682 1532 2683
rect 1526 2678 1527 2682
rect 1531 2678 1532 2682
rect 1526 2677 1532 2678
rect 1694 2682 1700 2683
rect 1694 2678 1695 2682
rect 1699 2678 1700 2682
rect 1694 2677 1700 2678
rect 2238 2676 2244 2677
rect 1870 2673 1876 2674
rect 135 2671 141 2672
rect 135 2667 136 2671
rect 140 2670 141 2671
rect 202 2671 208 2672
rect 202 2670 203 2671
rect 140 2668 203 2670
rect 140 2667 141 2668
rect 135 2666 141 2667
rect 202 2667 203 2668
rect 207 2667 208 2671
rect 202 2666 208 2667
rect 247 2671 253 2672
rect 247 2667 248 2671
rect 252 2670 253 2671
rect 262 2671 268 2672
rect 262 2670 263 2671
rect 252 2668 263 2670
rect 252 2667 253 2668
rect 247 2666 253 2667
rect 262 2667 263 2668
rect 267 2667 268 2671
rect 262 2666 268 2667
rect 354 2671 360 2672
rect 354 2667 355 2671
rect 359 2670 360 2671
rect 391 2671 397 2672
rect 391 2670 392 2671
rect 359 2668 392 2670
rect 359 2667 360 2668
rect 354 2666 360 2667
rect 391 2667 392 2668
rect 396 2667 397 2671
rect 391 2666 397 2667
rect 478 2671 484 2672
rect 478 2667 479 2671
rect 483 2670 484 2671
rect 551 2671 557 2672
rect 551 2670 552 2671
rect 483 2668 552 2670
rect 483 2667 484 2668
rect 478 2666 484 2667
rect 551 2667 552 2668
rect 556 2667 557 2671
rect 551 2666 557 2667
rect 703 2671 709 2672
rect 703 2667 704 2671
rect 708 2670 709 2671
rect 711 2671 717 2672
rect 711 2670 712 2671
rect 708 2668 712 2670
rect 708 2667 709 2668
rect 703 2666 709 2667
rect 711 2667 712 2668
rect 716 2667 717 2671
rect 711 2666 717 2667
rect 879 2671 885 2672
rect 879 2667 880 2671
rect 884 2670 885 2671
rect 894 2671 900 2672
rect 894 2670 895 2671
rect 884 2668 895 2670
rect 884 2667 885 2668
rect 879 2666 885 2667
rect 894 2667 895 2668
rect 899 2667 900 2671
rect 894 2666 900 2667
rect 962 2671 968 2672
rect 962 2667 963 2671
rect 967 2670 968 2671
rect 1039 2671 1045 2672
rect 1039 2670 1040 2671
rect 967 2668 1040 2670
rect 967 2667 968 2668
rect 962 2666 968 2667
rect 1039 2667 1040 2668
rect 1044 2667 1045 2671
rect 1039 2666 1045 2667
rect 1110 2671 1116 2672
rect 1110 2667 1111 2671
rect 1115 2670 1116 2671
rect 1199 2671 1205 2672
rect 1199 2670 1200 2671
rect 1115 2668 1200 2670
rect 1115 2667 1116 2668
rect 1110 2666 1116 2667
rect 1199 2667 1200 2668
rect 1204 2667 1205 2671
rect 1199 2666 1205 2667
rect 1359 2671 1365 2672
rect 1359 2667 1360 2671
rect 1364 2670 1365 2671
rect 1426 2671 1432 2672
rect 1426 2670 1427 2671
rect 1364 2668 1427 2670
rect 1364 2667 1365 2668
rect 1359 2666 1365 2667
rect 1426 2667 1427 2668
rect 1431 2667 1432 2671
rect 1426 2666 1432 2667
rect 1519 2671 1525 2672
rect 1519 2667 1520 2671
rect 1524 2670 1525 2671
rect 1586 2671 1592 2672
rect 1586 2670 1587 2671
rect 1524 2668 1587 2670
rect 1524 2667 1525 2668
rect 1519 2666 1525 2667
rect 1586 2667 1587 2668
rect 1591 2667 1592 2671
rect 1586 2666 1592 2667
rect 1687 2671 1693 2672
rect 1687 2667 1688 2671
rect 1692 2670 1693 2671
rect 1702 2671 1708 2672
rect 1702 2670 1703 2671
rect 1692 2668 1703 2670
rect 1692 2667 1693 2668
rect 1687 2666 1693 2667
rect 1702 2667 1703 2668
rect 1707 2667 1708 2671
rect 1870 2669 1871 2673
rect 1875 2669 1876 2673
rect 2238 2672 2239 2676
rect 2243 2672 2244 2676
rect 2238 2671 2244 2672
rect 2318 2676 2324 2677
rect 2318 2672 2319 2676
rect 2323 2672 2324 2676
rect 2318 2671 2324 2672
rect 2398 2676 2404 2677
rect 2398 2672 2399 2676
rect 2403 2672 2404 2676
rect 2398 2671 2404 2672
rect 2478 2676 2484 2677
rect 2478 2672 2479 2676
rect 2483 2672 2484 2676
rect 2478 2671 2484 2672
rect 2558 2676 2564 2677
rect 2558 2672 2559 2676
rect 2563 2672 2564 2676
rect 2558 2671 2564 2672
rect 2638 2676 2644 2677
rect 2638 2672 2639 2676
rect 2643 2672 2644 2676
rect 2638 2671 2644 2672
rect 2718 2676 2724 2677
rect 2718 2672 2719 2676
rect 2723 2672 2724 2676
rect 2718 2671 2724 2672
rect 2798 2676 2804 2677
rect 2798 2672 2799 2676
rect 2803 2672 2804 2676
rect 2798 2671 2804 2672
rect 2878 2676 2884 2677
rect 2878 2672 2879 2676
rect 2883 2672 2884 2676
rect 2878 2671 2884 2672
rect 2958 2676 2964 2677
rect 2958 2672 2959 2676
rect 2963 2672 2964 2676
rect 2958 2671 2964 2672
rect 3590 2673 3596 2674
rect 1870 2668 1876 2669
rect 3590 2669 3591 2673
rect 3595 2669 3596 2673
rect 3590 2668 3596 2669
rect 1702 2666 1708 2667
rect 2215 2667 2221 2668
rect 2215 2663 2216 2667
rect 2220 2666 2221 2667
rect 2311 2667 2317 2668
rect 2220 2664 2257 2666
rect 2220 2663 2221 2664
rect 2215 2662 2221 2663
rect 2311 2663 2312 2667
rect 2316 2666 2317 2667
rect 2386 2667 2392 2668
rect 2316 2664 2337 2666
rect 2316 2663 2317 2664
rect 2311 2662 2317 2663
rect 2386 2663 2387 2667
rect 2391 2666 2392 2667
rect 2466 2667 2472 2668
rect 2391 2664 2417 2666
rect 2391 2663 2392 2664
rect 2386 2662 2392 2663
rect 2466 2663 2467 2667
rect 2471 2666 2472 2667
rect 2546 2667 2552 2668
rect 2471 2664 2497 2666
rect 2471 2663 2472 2664
rect 2466 2662 2472 2663
rect 2546 2663 2547 2667
rect 2551 2666 2552 2667
rect 2706 2667 2712 2668
rect 2551 2664 2577 2666
rect 2640 2664 2657 2666
rect 2551 2663 2552 2664
rect 2546 2662 2552 2663
rect 2638 2663 2644 2664
rect 134 2659 141 2660
rect 134 2655 135 2659
rect 140 2655 141 2659
rect 134 2654 141 2655
rect 194 2659 200 2660
rect 194 2655 195 2659
rect 199 2658 200 2659
rect 247 2659 253 2660
rect 247 2658 248 2659
rect 199 2656 248 2658
rect 199 2655 200 2656
rect 194 2654 200 2655
rect 247 2655 248 2656
rect 252 2655 253 2659
rect 247 2654 253 2655
rect 306 2659 312 2660
rect 306 2655 307 2659
rect 311 2658 312 2659
rect 391 2659 397 2660
rect 391 2658 392 2659
rect 311 2656 392 2658
rect 311 2655 312 2656
rect 306 2654 312 2655
rect 391 2655 392 2656
rect 396 2655 397 2659
rect 391 2654 397 2655
rect 450 2659 456 2660
rect 450 2655 451 2659
rect 455 2658 456 2659
rect 543 2659 549 2660
rect 543 2658 544 2659
rect 455 2656 544 2658
rect 455 2655 456 2656
rect 450 2654 456 2655
rect 543 2655 544 2656
rect 548 2655 549 2659
rect 543 2654 549 2655
rect 602 2659 608 2660
rect 602 2655 603 2659
rect 607 2658 608 2659
rect 703 2659 709 2660
rect 703 2658 704 2659
rect 607 2656 704 2658
rect 607 2655 608 2656
rect 602 2654 608 2655
rect 703 2655 704 2656
rect 708 2655 709 2659
rect 703 2654 709 2655
rect 871 2659 877 2660
rect 871 2655 872 2659
rect 876 2658 877 2659
rect 938 2659 944 2660
rect 938 2658 939 2659
rect 876 2656 939 2658
rect 876 2655 877 2656
rect 871 2654 877 2655
rect 938 2655 939 2656
rect 943 2655 944 2659
rect 938 2654 944 2655
rect 1039 2659 1045 2660
rect 1039 2655 1040 2659
rect 1044 2658 1045 2659
rect 1134 2659 1140 2660
rect 1134 2658 1135 2659
rect 1044 2656 1135 2658
rect 1044 2655 1045 2656
rect 1039 2654 1045 2655
rect 1134 2655 1135 2656
rect 1139 2655 1140 2659
rect 1134 2654 1140 2655
rect 1186 2659 1192 2660
rect 1186 2655 1187 2659
rect 1191 2658 1192 2659
rect 1207 2659 1213 2660
rect 1207 2658 1208 2659
rect 1191 2656 1208 2658
rect 1191 2655 1192 2656
rect 1186 2654 1192 2655
rect 1207 2655 1208 2656
rect 1212 2655 1213 2659
rect 1207 2654 1213 2655
rect 1358 2659 1364 2660
rect 1358 2655 1359 2659
rect 1363 2658 1364 2659
rect 1383 2659 1389 2660
rect 1383 2658 1384 2659
rect 1363 2656 1384 2658
rect 1363 2655 1364 2656
rect 1358 2654 1364 2655
rect 1383 2655 1384 2656
rect 1388 2655 1389 2659
rect 1383 2654 1389 2655
rect 1442 2659 1448 2660
rect 1442 2655 1443 2659
rect 1447 2658 1448 2659
rect 1559 2659 1565 2660
rect 1559 2658 1560 2659
rect 1447 2656 1560 2658
rect 1447 2655 1448 2656
rect 1442 2654 1448 2655
rect 1559 2655 1560 2656
rect 1564 2655 1565 2659
rect 2638 2659 2639 2663
rect 2643 2659 2644 2663
rect 2706 2663 2707 2667
rect 2711 2666 2712 2667
rect 2866 2667 2872 2668
rect 2866 2666 2867 2667
rect 2711 2664 2737 2666
rect 2861 2664 2867 2666
rect 2711 2663 2712 2664
rect 2706 2662 2712 2663
rect 2866 2663 2867 2664
rect 2871 2663 2872 2667
rect 2946 2667 2952 2668
rect 2946 2666 2947 2667
rect 2941 2664 2947 2666
rect 2866 2662 2872 2663
rect 2946 2663 2947 2664
rect 2951 2663 2952 2667
rect 2946 2662 2952 2663
rect 2638 2658 2644 2659
rect 2786 2659 2792 2660
rect 1559 2654 1565 2655
rect 1870 2656 1876 2657
rect 1870 2652 1871 2656
rect 1875 2652 1876 2656
rect 2786 2655 2787 2659
rect 2791 2658 2792 2659
rect 2976 2658 2978 2665
rect 2791 2656 2978 2658
rect 3590 2656 3596 2657
rect 2791 2655 2792 2656
rect 2786 2654 2792 2655
rect 1870 2651 1876 2652
rect 3590 2652 3591 2656
rect 3595 2652 3596 2656
rect 3590 2651 3596 2652
rect 142 2650 148 2651
rect 142 2646 143 2650
rect 147 2646 148 2650
rect 142 2645 148 2646
rect 254 2650 260 2651
rect 254 2646 255 2650
rect 259 2646 260 2650
rect 254 2645 260 2646
rect 398 2650 404 2651
rect 398 2646 399 2650
rect 403 2646 404 2650
rect 398 2645 404 2646
rect 550 2650 556 2651
rect 550 2646 551 2650
rect 555 2646 556 2650
rect 550 2645 556 2646
rect 710 2650 716 2651
rect 710 2646 711 2650
rect 715 2646 716 2650
rect 710 2645 716 2646
rect 878 2650 884 2651
rect 878 2646 879 2650
rect 883 2646 884 2650
rect 878 2645 884 2646
rect 1046 2650 1052 2651
rect 1046 2646 1047 2650
rect 1051 2646 1052 2650
rect 1046 2645 1052 2646
rect 1214 2650 1220 2651
rect 1214 2646 1215 2650
rect 1219 2646 1220 2650
rect 1214 2645 1220 2646
rect 1390 2650 1396 2651
rect 1390 2646 1391 2650
rect 1395 2646 1396 2650
rect 1390 2645 1396 2646
rect 1566 2650 1572 2651
rect 1566 2646 1567 2650
rect 1571 2646 1572 2650
rect 1566 2645 1572 2646
rect 2246 2638 2252 2639
rect 2246 2634 2247 2638
rect 2251 2634 2252 2638
rect 2246 2633 2252 2634
rect 2326 2638 2332 2639
rect 2326 2634 2327 2638
rect 2331 2634 2332 2638
rect 2326 2633 2332 2634
rect 2406 2638 2412 2639
rect 2406 2634 2407 2638
rect 2411 2634 2412 2638
rect 2406 2633 2412 2634
rect 2486 2638 2492 2639
rect 2486 2634 2487 2638
rect 2491 2634 2492 2638
rect 2486 2633 2492 2634
rect 2566 2638 2572 2639
rect 2566 2634 2567 2638
rect 2571 2634 2572 2638
rect 2566 2633 2572 2634
rect 2646 2638 2652 2639
rect 2646 2634 2647 2638
rect 2651 2634 2652 2638
rect 2646 2633 2652 2634
rect 2726 2638 2732 2639
rect 2726 2634 2727 2638
rect 2731 2634 2732 2638
rect 2806 2638 2812 2639
rect 2786 2635 2792 2636
rect 2786 2634 2787 2635
rect 2726 2633 2732 2634
rect 110 2632 116 2633
rect 110 2628 111 2632
rect 115 2628 116 2632
rect 110 2627 116 2628
rect 1830 2632 1836 2633
rect 1830 2628 1831 2632
rect 1835 2628 1836 2632
rect 2772 2632 2787 2634
rect 1830 2627 1836 2628
rect 2239 2627 2245 2628
rect 194 2623 200 2624
rect 194 2619 195 2623
rect 199 2619 200 2623
rect 194 2618 200 2619
rect 306 2623 312 2624
rect 306 2619 307 2623
rect 311 2619 312 2623
rect 306 2618 312 2619
rect 450 2623 456 2624
rect 450 2619 451 2623
rect 455 2619 456 2623
rect 450 2618 456 2619
rect 602 2623 608 2624
rect 602 2619 603 2623
rect 607 2619 608 2623
rect 602 2618 608 2619
rect 894 2623 900 2624
rect 894 2619 895 2623
rect 899 2619 900 2623
rect 894 2618 900 2619
rect 938 2623 944 2624
rect 938 2619 939 2623
rect 943 2622 944 2623
rect 1134 2623 1140 2624
rect 943 2620 1057 2622
rect 943 2619 944 2620
rect 938 2618 944 2619
rect 1134 2619 1135 2623
rect 1139 2622 1140 2623
rect 1442 2623 1448 2624
rect 1139 2620 1225 2622
rect 1139 2619 1140 2620
rect 1134 2618 1140 2619
rect 1442 2619 1443 2623
rect 1447 2619 1448 2623
rect 2239 2623 2240 2627
rect 2244 2626 2245 2627
rect 2311 2627 2317 2628
rect 2311 2626 2312 2627
rect 2244 2624 2312 2626
rect 2244 2623 2245 2624
rect 2239 2622 2245 2623
rect 2311 2623 2312 2624
rect 2316 2623 2317 2627
rect 2311 2622 2317 2623
rect 2319 2627 2325 2628
rect 2319 2623 2320 2627
rect 2324 2626 2325 2627
rect 2386 2627 2392 2628
rect 2386 2626 2387 2627
rect 2324 2624 2387 2626
rect 2324 2623 2325 2624
rect 2319 2622 2325 2623
rect 2386 2623 2387 2624
rect 2391 2623 2392 2627
rect 2386 2622 2392 2623
rect 2399 2627 2405 2628
rect 2399 2623 2400 2627
rect 2404 2626 2405 2627
rect 2466 2627 2472 2628
rect 2466 2626 2467 2627
rect 2404 2624 2467 2626
rect 2404 2623 2405 2624
rect 2399 2622 2405 2623
rect 2466 2623 2467 2624
rect 2471 2623 2472 2627
rect 2466 2622 2472 2623
rect 2479 2627 2485 2628
rect 2479 2623 2480 2627
rect 2484 2626 2485 2627
rect 2546 2627 2552 2628
rect 2546 2626 2547 2627
rect 2484 2624 2547 2626
rect 2484 2623 2485 2624
rect 2479 2622 2485 2623
rect 2546 2623 2547 2624
rect 2551 2623 2552 2627
rect 2546 2622 2552 2623
rect 2559 2627 2565 2628
rect 2559 2623 2560 2627
rect 2564 2626 2565 2627
rect 2598 2627 2604 2628
rect 2598 2626 2599 2627
rect 2564 2624 2599 2626
rect 2564 2623 2565 2624
rect 2559 2622 2565 2623
rect 2598 2623 2599 2624
rect 2603 2623 2604 2627
rect 2598 2622 2604 2623
rect 2639 2627 2645 2628
rect 2639 2623 2640 2627
rect 2644 2626 2645 2627
rect 2706 2627 2712 2628
rect 2706 2626 2707 2627
rect 2644 2624 2707 2626
rect 2644 2623 2645 2624
rect 2639 2622 2645 2623
rect 2706 2623 2707 2624
rect 2711 2623 2712 2627
rect 2706 2622 2712 2623
rect 2719 2627 2725 2628
rect 2719 2623 2720 2627
rect 2724 2626 2725 2627
rect 2772 2626 2774 2632
rect 2786 2631 2787 2632
rect 2791 2631 2792 2635
rect 2806 2634 2807 2638
rect 2811 2634 2812 2638
rect 2806 2633 2812 2634
rect 2886 2638 2892 2639
rect 2886 2634 2887 2638
rect 2891 2634 2892 2638
rect 2886 2633 2892 2634
rect 2966 2638 2972 2639
rect 2966 2634 2967 2638
rect 2971 2634 2972 2638
rect 2966 2633 2972 2634
rect 2786 2630 2792 2631
rect 2724 2624 2774 2626
rect 2778 2627 2784 2628
rect 2724 2623 2725 2624
rect 2719 2622 2725 2623
rect 2778 2623 2779 2627
rect 2783 2626 2784 2627
rect 2799 2627 2805 2628
rect 2799 2626 2800 2627
rect 2783 2624 2800 2626
rect 2783 2623 2784 2624
rect 2778 2622 2784 2623
rect 2799 2623 2800 2624
rect 2804 2623 2805 2627
rect 2799 2622 2805 2623
rect 2866 2627 2872 2628
rect 2866 2623 2867 2627
rect 2871 2626 2872 2627
rect 2879 2627 2885 2628
rect 2879 2626 2880 2627
rect 2871 2624 2880 2626
rect 2871 2623 2872 2624
rect 2866 2622 2872 2623
rect 2879 2623 2880 2624
rect 2884 2623 2885 2627
rect 2879 2622 2885 2623
rect 2946 2627 2952 2628
rect 2946 2623 2947 2627
rect 2951 2626 2952 2627
rect 2959 2627 2965 2628
rect 2959 2626 2960 2627
rect 2951 2624 2960 2626
rect 2951 2623 2952 2624
rect 2946 2622 2952 2623
rect 2959 2623 2960 2624
rect 2964 2623 2965 2627
rect 2959 2622 2965 2623
rect 1442 2618 1448 2619
rect 110 2615 116 2616
rect 110 2611 111 2615
rect 115 2611 116 2615
rect 1830 2615 1836 2616
rect 110 2610 116 2611
rect 134 2612 140 2613
rect 134 2608 135 2612
rect 139 2608 140 2612
rect 134 2607 140 2608
rect 246 2612 252 2613
rect 246 2608 247 2612
rect 251 2608 252 2612
rect 246 2607 252 2608
rect 390 2612 396 2613
rect 390 2608 391 2612
rect 395 2608 396 2612
rect 390 2607 396 2608
rect 542 2612 548 2613
rect 542 2608 543 2612
rect 547 2608 548 2612
rect 542 2607 548 2608
rect 702 2612 708 2613
rect 702 2608 703 2612
rect 707 2608 708 2612
rect 702 2607 708 2608
rect 870 2612 876 2613
rect 870 2608 871 2612
rect 875 2608 876 2612
rect 870 2607 876 2608
rect 1038 2612 1044 2613
rect 1038 2608 1039 2612
rect 1043 2608 1044 2612
rect 1038 2607 1044 2608
rect 1206 2612 1212 2613
rect 1206 2608 1207 2612
rect 1211 2608 1212 2612
rect 1206 2607 1212 2608
rect 1382 2612 1388 2613
rect 1382 2608 1383 2612
rect 1387 2608 1388 2612
rect 1382 2607 1388 2608
rect 1558 2612 1564 2613
rect 1558 2608 1559 2612
rect 1563 2608 1564 2612
rect 1830 2611 1831 2615
rect 1835 2611 1836 2615
rect 2474 2615 2480 2616
rect 2474 2614 2475 2615
rect 1830 2610 1836 2611
rect 2244 2612 2475 2614
rect 1558 2607 1564 2608
rect 2183 2607 2189 2608
rect 2183 2603 2184 2607
rect 2188 2606 2189 2607
rect 2244 2606 2246 2612
rect 2474 2611 2475 2612
rect 2479 2611 2480 2615
rect 2474 2610 2480 2611
rect 2188 2604 2246 2606
rect 2254 2607 2260 2608
rect 2188 2603 2189 2604
rect 2183 2602 2189 2603
rect 2254 2603 2255 2607
rect 2259 2606 2260 2607
rect 2263 2607 2269 2608
rect 2263 2606 2264 2607
rect 2259 2604 2264 2606
rect 2259 2603 2260 2604
rect 2254 2602 2260 2603
rect 2263 2603 2264 2604
rect 2268 2603 2269 2607
rect 2263 2602 2269 2603
rect 2334 2607 2340 2608
rect 2334 2603 2335 2607
rect 2339 2606 2340 2607
rect 2343 2607 2349 2608
rect 2343 2606 2344 2607
rect 2339 2604 2344 2606
rect 2339 2603 2340 2604
rect 2334 2602 2340 2603
rect 2343 2603 2344 2604
rect 2348 2603 2349 2607
rect 2343 2602 2349 2603
rect 2414 2607 2420 2608
rect 2414 2603 2415 2607
rect 2419 2606 2420 2607
rect 2423 2607 2429 2608
rect 2423 2606 2424 2607
rect 2419 2604 2424 2606
rect 2419 2603 2420 2604
rect 2414 2602 2420 2603
rect 2423 2603 2424 2604
rect 2428 2603 2429 2607
rect 2423 2602 2429 2603
rect 2494 2607 2500 2608
rect 2494 2603 2495 2607
rect 2499 2606 2500 2607
rect 2503 2607 2509 2608
rect 2503 2606 2504 2607
rect 2499 2604 2504 2606
rect 2499 2603 2500 2604
rect 2494 2602 2500 2603
rect 2503 2603 2504 2604
rect 2508 2603 2509 2607
rect 2503 2602 2509 2603
rect 2582 2607 2589 2608
rect 2582 2603 2583 2607
rect 2588 2603 2589 2607
rect 2582 2602 2589 2603
rect 2638 2607 2644 2608
rect 2638 2603 2639 2607
rect 2643 2606 2644 2607
rect 2663 2607 2669 2608
rect 2663 2606 2664 2607
rect 2643 2604 2664 2606
rect 2643 2603 2644 2604
rect 2638 2602 2644 2603
rect 2663 2603 2664 2604
rect 2668 2603 2669 2607
rect 2663 2602 2669 2603
rect 2734 2607 2740 2608
rect 2734 2603 2735 2607
rect 2739 2606 2740 2607
rect 2743 2607 2749 2608
rect 2743 2606 2744 2607
rect 2739 2604 2744 2606
rect 2739 2603 2740 2604
rect 2734 2602 2740 2603
rect 2743 2603 2744 2604
rect 2748 2603 2749 2607
rect 2743 2602 2749 2603
rect 2814 2607 2820 2608
rect 2814 2603 2815 2607
rect 2819 2606 2820 2607
rect 2823 2607 2829 2608
rect 2823 2606 2824 2607
rect 2819 2604 2824 2606
rect 2819 2603 2820 2604
rect 2814 2602 2820 2603
rect 2823 2603 2824 2604
rect 2828 2603 2829 2607
rect 2823 2602 2829 2603
rect 2894 2607 2900 2608
rect 2894 2603 2895 2607
rect 2899 2606 2900 2607
rect 2903 2607 2909 2608
rect 2903 2606 2904 2607
rect 2899 2604 2904 2606
rect 2899 2603 2900 2604
rect 2894 2602 2900 2603
rect 2903 2603 2904 2604
rect 2908 2603 2909 2607
rect 2903 2602 2909 2603
rect 2974 2607 2980 2608
rect 2974 2603 2975 2607
rect 2979 2606 2980 2607
rect 2983 2607 2989 2608
rect 2983 2606 2984 2607
rect 2979 2604 2984 2606
rect 2979 2603 2980 2604
rect 2974 2602 2980 2603
rect 2983 2603 2984 2604
rect 2988 2603 2989 2607
rect 2983 2602 2989 2603
rect 2190 2598 2196 2599
rect 642 2595 648 2596
rect 642 2591 643 2595
rect 647 2594 648 2595
rect 719 2595 725 2596
rect 719 2594 720 2595
rect 647 2592 720 2594
rect 647 2591 648 2592
rect 642 2590 648 2591
rect 719 2591 720 2592
rect 724 2591 725 2595
rect 719 2590 725 2591
rect 1542 2595 1548 2596
rect 1542 2591 1543 2595
rect 1547 2594 1548 2595
rect 1575 2595 1581 2596
rect 1575 2594 1576 2595
rect 1547 2592 1576 2594
rect 1547 2591 1548 2592
rect 1542 2590 1548 2591
rect 1575 2591 1576 2592
rect 1580 2591 1581 2595
rect 2190 2594 2191 2598
rect 2195 2594 2196 2598
rect 2190 2593 2196 2594
rect 2270 2598 2276 2599
rect 2270 2594 2271 2598
rect 2275 2594 2276 2598
rect 2270 2593 2276 2594
rect 2350 2598 2356 2599
rect 2350 2594 2351 2598
rect 2355 2594 2356 2598
rect 2350 2593 2356 2594
rect 2430 2598 2436 2599
rect 2430 2594 2431 2598
rect 2435 2594 2436 2598
rect 2430 2593 2436 2594
rect 2510 2598 2516 2599
rect 2510 2594 2511 2598
rect 2515 2594 2516 2598
rect 2510 2593 2516 2594
rect 2590 2598 2596 2599
rect 2590 2594 2591 2598
rect 2595 2594 2596 2598
rect 2590 2593 2596 2594
rect 2670 2598 2676 2599
rect 2670 2594 2671 2598
rect 2675 2594 2676 2598
rect 2670 2593 2676 2594
rect 2750 2598 2756 2599
rect 2750 2594 2751 2598
rect 2755 2594 2756 2598
rect 2750 2593 2756 2594
rect 2830 2598 2836 2599
rect 2830 2594 2831 2598
rect 2835 2594 2836 2598
rect 2830 2593 2836 2594
rect 2910 2598 2916 2599
rect 2910 2594 2911 2598
rect 2915 2594 2916 2598
rect 2910 2593 2916 2594
rect 2990 2598 2996 2599
rect 2990 2594 2991 2598
rect 2995 2594 2996 2598
rect 2990 2593 2996 2594
rect 1575 2590 1581 2591
rect 1870 2580 1876 2581
rect 1870 2576 1871 2580
rect 1875 2576 1876 2580
rect 1870 2575 1876 2576
rect 3590 2580 3596 2581
rect 3590 2576 3591 2580
rect 3595 2576 3596 2580
rect 3590 2575 3596 2576
rect 2254 2571 2260 2572
rect 2254 2570 2255 2571
rect 2245 2568 2255 2570
rect 2254 2567 2255 2568
rect 2259 2567 2260 2571
rect 2334 2571 2340 2572
rect 2334 2570 2335 2571
rect 2325 2568 2335 2570
rect 2254 2566 2260 2567
rect 2334 2567 2335 2568
rect 2339 2567 2340 2571
rect 2414 2571 2420 2572
rect 2414 2570 2415 2571
rect 2405 2568 2415 2570
rect 2334 2566 2340 2567
rect 2414 2567 2415 2568
rect 2419 2567 2420 2571
rect 2494 2571 2500 2572
rect 2494 2570 2495 2571
rect 2485 2568 2495 2570
rect 2414 2566 2420 2567
rect 2494 2567 2495 2568
rect 2499 2567 2500 2571
rect 2582 2571 2588 2572
rect 2582 2570 2583 2571
rect 2565 2568 2583 2570
rect 2494 2566 2500 2567
rect 2582 2567 2583 2568
rect 2587 2567 2588 2571
rect 2582 2566 2588 2567
rect 2598 2571 2604 2572
rect 2598 2567 2599 2571
rect 2603 2567 2604 2571
rect 2734 2571 2740 2572
rect 2734 2570 2735 2571
rect 2725 2568 2735 2570
rect 2598 2566 2604 2567
rect 2734 2567 2735 2568
rect 2739 2567 2740 2571
rect 2814 2571 2820 2572
rect 2814 2570 2815 2571
rect 2805 2568 2815 2570
rect 2734 2566 2740 2567
rect 2814 2567 2815 2568
rect 2819 2567 2820 2571
rect 2894 2571 2900 2572
rect 2894 2570 2895 2571
rect 2885 2568 2895 2570
rect 2814 2566 2820 2567
rect 2894 2567 2895 2568
rect 2899 2567 2900 2571
rect 2974 2571 2980 2572
rect 2974 2570 2975 2571
rect 2965 2568 2975 2570
rect 2894 2566 2900 2567
rect 2974 2567 2975 2568
rect 2979 2567 2980 2571
rect 2974 2566 2980 2567
rect 158 2564 164 2565
rect 110 2561 116 2562
rect 110 2557 111 2561
rect 115 2557 116 2561
rect 158 2560 159 2564
rect 163 2560 164 2564
rect 158 2559 164 2560
rect 278 2564 284 2565
rect 278 2560 279 2564
rect 283 2560 284 2564
rect 278 2559 284 2560
rect 414 2564 420 2565
rect 414 2560 415 2564
rect 419 2560 420 2564
rect 414 2559 420 2560
rect 558 2564 564 2565
rect 558 2560 559 2564
rect 563 2560 564 2564
rect 558 2559 564 2560
rect 702 2564 708 2565
rect 702 2560 703 2564
rect 707 2560 708 2564
rect 702 2559 708 2560
rect 846 2564 852 2565
rect 846 2560 847 2564
rect 851 2560 852 2564
rect 846 2559 852 2560
rect 982 2564 988 2565
rect 982 2560 983 2564
rect 987 2560 988 2564
rect 982 2559 988 2560
rect 1118 2564 1124 2565
rect 1118 2560 1119 2564
rect 1123 2560 1124 2564
rect 1118 2559 1124 2560
rect 1254 2564 1260 2565
rect 1254 2560 1255 2564
rect 1259 2560 1260 2564
rect 1254 2559 1260 2560
rect 1390 2564 1396 2565
rect 1390 2560 1391 2564
rect 1395 2560 1396 2564
rect 1390 2559 1396 2560
rect 1526 2564 1532 2565
rect 1526 2560 1527 2564
rect 1531 2560 1532 2564
rect 1870 2563 1876 2564
rect 1526 2559 1532 2560
rect 1830 2561 1836 2562
rect 110 2556 116 2557
rect 1830 2557 1831 2561
rect 1835 2557 1836 2561
rect 1870 2559 1871 2563
rect 1875 2559 1876 2563
rect 3590 2563 3596 2564
rect 1870 2558 1876 2559
rect 2182 2560 2188 2561
rect 1830 2556 1836 2557
rect 2182 2556 2183 2560
rect 2187 2556 2188 2560
rect 226 2555 232 2556
rect 226 2554 227 2555
rect 221 2552 227 2554
rect 226 2551 227 2552
rect 231 2551 232 2555
rect 346 2555 352 2556
rect 346 2554 347 2555
rect 341 2552 347 2554
rect 226 2550 232 2551
rect 346 2551 347 2552
rect 351 2551 352 2555
rect 482 2555 488 2556
rect 482 2554 483 2555
rect 477 2552 483 2554
rect 346 2550 352 2551
rect 482 2551 483 2552
rect 487 2551 488 2555
rect 634 2555 640 2556
rect 634 2554 635 2555
rect 621 2552 635 2554
rect 482 2550 488 2551
rect 634 2551 635 2552
rect 639 2551 640 2555
rect 634 2550 640 2551
rect 666 2555 672 2556
rect 666 2551 667 2555
rect 671 2554 672 2555
rect 914 2555 920 2556
rect 914 2554 915 2555
rect 671 2552 721 2554
rect 909 2552 915 2554
rect 671 2551 672 2552
rect 666 2550 672 2551
rect 914 2551 915 2552
rect 919 2551 920 2555
rect 1050 2555 1056 2556
rect 1050 2554 1051 2555
rect 1045 2552 1051 2554
rect 914 2550 920 2551
rect 1050 2551 1051 2552
rect 1055 2551 1056 2555
rect 1186 2555 1192 2556
rect 1186 2554 1187 2555
rect 1181 2552 1187 2554
rect 1050 2550 1056 2551
rect 1186 2551 1187 2552
rect 1191 2551 1192 2555
rect 1330 2555 1336 2556
rect 1186 2550 1192 2551
rect 1316 2548 1318 2553
rect 1330 2551 1331 2555
rect 1335 2554 1336 2555
rect 1478 2555 1484 2556
rect 2182 2555 2188 2556
rect 2262 2560 2268 2561
rect 2262 2556 2263 2560
rect 2267 2556 2268 2560
rect 2262 2555 2268 2556
rect 2342 2560 2348 2561
rect 2342 2556 2343 2560
rect 2347 2556 2348 2560
rect 2342 2555 2348 2556
rect 2422 2560 2428 2561
rect 2422 2556 2423 2560
rect 2427 2556 2428 2560
rect 2422 2555 2428 2556
rect 2502 2560 2508 2561
rect 2502 2556 2503 2560
rect 2507 2556 2508 2560
rect 2502 2555 2508 2556
rect 2582 2560 2588 2561
rect 2582 2556 2583 2560
rect 2587 2556 2588 2560
rect 2582 2555 2588 2556
rect 2662 2560 2668 2561
rect 2662 2556 2663 2560
rect 2667 2556 2668 2560
rect 2662 2555 2668 2556
rect 2742 2560 2748 2561
rect 2742 2556 2743 2560
rect 2747 2556 2748 2560
rect 2742 2555 2748 2556
rect 2822 2560 2828 2561
rect 2822 2556 2823 2560
rect 2827 2556 2828 2560
rect 2822 2555 2828 2556
rect 2902 2560 2908 2561
rect 2902 2556 2903 2560
rect 2907 2556 2908 2560
rect 2902 2555 2908 2556
rect 2982 2560 2988 2561
rect 2982 2556 2983 2560
rect 2987 2556 2988 2560
rect 3590 2559 3591 2563
rect 3595 2559 3596 2563
rect 3590 2558 3596 2559
rect 2982 2555 2988 2556
rect 1335 2552 1409 2554
rect 1335 2551 1336 2552
rect 1330 2550 1336 2551
rect 1478 2551 1479 2555
rect 1483 2554 1484 2555
rect 1483 2552 1545 2554
rect 1483 2551 1484 2552
rect 1478 2550 1484 2551
rect 1314 2547 1320 2548
rect 110 2544 116 2545
rect 110 2540 111 2544
rect 115 2540 116 2544
rect 1314 2543 1315 2547
rect 1319 2543 1320 2547
rect 1314 2542 1320 2543
rect 1830 2544 1836 2545
rect 110 2539 116 2540
rect 1830 2540 1831 2544
rect 1835 2540 1836 2544
rect 1830 2539 1836 2540
rect 2606 2543 2612 2544
rect 2606 2539 2607 2543
rect 2611 2542 2612 2543
rect 2999 2543 3005 2544
rect 2999 2542 3000 2543
rect 2611 2540 3000 2542
rect 2611 2539 2612 2540
rect 2606 2538 2612 2539
rect 2999 2539 3000 2540
rect 3004 2539 3005 2543
rect 2999 2538 3005 2539
rect 166 2526 172 2527
rect 166 2522 167 2526
rect 171 2522 172 2526
rect 166 2521 172 2522
rect 286 2526 292 2527
rect 286 2522 287 2526
rect 291 2522 292 2526
rect 286 2521 292 2522
rect 422 2526 428 2527
rect 422 2522 423 2526
rect 427 2522 428 2526
rect 422 2521 428 2522
rect 566 2526 572 2527
rect 566 2522 567 2526
rect 571 2522 572 2526
rect 566 2521 572 2522
rect 710 2526 716 2527
rect 710 2522 711 2526
rect 715 2522 716 2526
rect 710 2521 716 2522
rect 854 2526 860 2527
rect 854 2522 855 2526
rect 859 2522 860 2526
rect 854 2521 860 2522
rect 990 2526 996 2527
rect 990 2522 991 2526
rect 995 2522 996 2526
rect 990 2521 996 2522
rect 1126 2526 1132 2527
rect 1126 2522 1127 2526
rect 1131 2522 1132 2526
rect 1126 2521 1132 2522
rect 1262 2526 1268 2527
rect 1262 2522 1263 2526
rect 1267 2522 1268 2526
rect 1262 2521 1268 2522
rect 1398 2526 1404 2527
rect 1398 2522 1399 2526
rect 1403 2522 1404 2526
rect 1398 2521 1404 2522
rect 1534 2526 1540 2527
rect 1534 2522 1535 2526
rect 1539 2522 1540 2526
rect 1534 2521 1540 2522
rect 159 2515 165 2516
rect 159 2511 160 2515
rect 164 2514 165 2515
rect 174 2515 180 2516
rect 174 2514 175 2515
rect 164 2512 175 2514
rect 164 2511 165 2512
rect 159 2510 165 2511
rect 174 2511 175 2512
rect 179 2511 180 2515
rect 174 2510 180 2511
rect 226 2515 232 2516
rect 226 2511 227 2515
rect 231 2514 232 2515
rect 279 2515 285 2516
rect 279 2514 280 2515
rect 231 2512 280 2514
rect 231 2511 232 2512
rect 226 2510 232 2511
rect 279 2511 280 2512
rect 284 2511 285 2515
rect 279 2510 285 2511
rect 346 2515 352 2516
rect 346 2511 347 2515
rect 351 2514 352 2515
rect 415 2515 421 2516
rect 415 2514 416 2515
rect 351 2512 416 2514
rect 351 2511 352 2512
rect 346 2510 352 2511
rect 415 2511 416 2512
rect 420 2511 421 2515
rect 415 2510 421 2511
rect 482 2515 488 2516
rect 482 2511 483 2515
rect 487 2514 488 2515
rect 559 2515 565 2516
rect 559 2514 560 2515
rect 487 2512 560 2514
rect 487 2511 488 2512
rect 482 2510 488 2511
rect 559 2511 560 2512
rect 564 2511 565 2515
rect 559 2510 565 2511
rect 634 2515 640 2516
rect 634 2511 635 2515
rect 639 2514 640 2515
rect 703 2515 709 2516
rect 703 2514 704 2515
rect 639 2512 704 2514
rect 639 2511 640 2512
rect 634 2510 640 2511
rect 703 2511 704 2512
rect 708 2511 709 2515
rect 703 2510 709 2511
rect 847 2515 853 2516
rect 847 2511 848 2515
rect 852 2514 853 2515
rect 886 2515 892 2516
rect 886 2514 887 2515
rect 852 2512 887 2514
rect 852 2511 853 2512
rect 847 2510 853 2511
rect 886 2511 887 2512
rect 891 2511 892 2515
rect 886 2510 892 2511
rect 914 2515 920 2516
rect 914 2511 915 2515
rect 919 2514 920 2515
rect 983 2515 989 2516
rect 983 2514 984 2515
rect 919 2512 984 2514
rect 919 2511 920 2512
rect 914 2510 920 2511
rect 983 2511 984 2512
rect 988 2511 989 2515
rect 983 2510 989 2511
rect 1050 2515 1056 2516
rect 1050 2511 1051 2515
rect 1055 2514 1056 2515
rect 1119 2515 1125 2516
rect 1119 2514 1120 2515
rect 1055 2512 1120 2514
rect 1055 2511 1056 2512
rect 1050 2510 1056 2511
rect 1119 2511 1120 2512
rect 1124 2511 1125 2515
rect 1119 2510 1125 2511
rect 1255 2515 1261 2516
rect 1255 2511 1256 2515
rect 1260 2514 1261 2515
rect 1330 2515 1336 2516
rect 1330 2514 1331 2515
rect 1260 2512 1331 2514
rect 1260 2511 1261 2512
rect 1255 2510 1261 2511
rect 1330 2511 1331 2512
rect 1335 2511 1336 2515
rect 1330 2510 1336 2511
rect 1391 2515 1397 2516
rect 1391 2511 1392 2515
rect 1396 2514 1397 2515
rect 1478 2515 1484 2516
rect 1478 2514 1479 2515
rect 1396 2512 1479 2514
rect 1396 2511 1397 2512
rect 1391 2510 1397 2511
rect 1478 2511 1479 2512
rect 1483 2511 1484 2515
rect 1478 2510 1484 2511
rect 1527 2515 1533 2516
rect 1527 2511 1528 2515
rect 1532 2514 1533 2515
rect 1542 2515 1548 2516
rect 1542 2514 1543 2515
rect 1532 2512 1543 2514
rect 1532 2511 1533 2512
rect 1527 2510 1533 2511
rect 1542 2511 1543 2512
rect 1547 2511 1548 2515
rect 1542 2510 1548 2511
rect 2118 2508 2124 2509
rect 1870 2505 1876 2506
rect 1870 2501 1871 2505
rect 1875 2501 1876 2505
rect 2118 2504 2119 2508
rect 2123 2504 2124 2508
rect 2118 2503 2124 2504
rect 2206 2508 2212 2509
rect 2206 2504 2207 2508
rect 2211 2504 2212 2508
rect 2206 2503 2212 2504
rect 2302 2508 2308 2509
rect 2302 2504 2303 2508
rect 2307 2504 2308 2508
rect 2302 2503 2308 2504
rect 2398 2508 2404 2509
rect 2398 2504 2399 2508
rect 2403 2504 2404 2508
rect 2398 2503 2404 2504
rect 2494 2508 2500 2509
rect 2494 2504 2495 2508
rect 2499 2504 2500 2508
rect 2494 2503 2500 2504
rect 2590 2508 2596 2509
rect 2590 2504 2591 2508
rect 2595 2504 2596 2508
rect 2590 2503 2596 2504
rect 2686 2508 2692 2509
rect 2686 2504 2687 2508
rect 2691 2504 2692 2508
rect 2686 2503 2692 2504
rect 2782 2508 2788 2509
rect 2782 2504 2783 2508
rect 2787 2504 2788 2508
rect 2782 2503 2788 2504
rect 2878 2508 2884 2509
rect 2878 2504 2879 2508
rect 2883 2504 2884 2508
rect 2878 2503 2884 2504
rect 2974 2508 2980 2509
rect 2974 2504 2975 2508
rect 2979 2504 2980 2508
rect 2974 2503 2980 2504
rect 3078 2508 3084 2509
rect 3078 2504 3079 2508
rect 3083 2504 3084 2508
rect 3078 2503 3084 2504
rect 3590 2505 3596 2506
rect 1870 2500 1876 2501
rect 3590 2501 3591 2505
rect 3595 2501 3596 2505
rect 3590 2500 3596 2501
rect 327 2499 333 2500
rect 327 2495 328 2499
rect 332 2498 333 2499
rect 354 2499 360 2500
rect 354 2498 355 2499
rect 332 2496 355 2498
rect 332 2495 333 2496
rect 327 2494 333 2495
rect 354 2495 355 2496
rect 359 2495 360 2499
rect 354 2494 360 2495
rect 386 2499 392 2500
rect 386 2495 387 2499
rect 391 2498 392 2499
rect 407 2499 413 2500
rect 407 2498 408 2499
rect 391 2496 408 2498
rect 391 2495 392 2496
rect 386 2494 392 2495
rect 407 2495 408 2496
rect 412 2495 413 2499
rect 407 2494 413 2495
rect 466 2499 472 2500
rect 466 2495 467 2499
rect 471 2498 472 2499
rect 495 2499 501 2500
rect 495 2498 496 2499
rect 471 2496 496 2498
rect 471 2495 472 2496
rect 466 2494 472 2495
rect 495 2495 496 2496
rect 500 2495 501 2499
rect 495 2494 501 2495
rect 554 2499 560 2500
rect 554 2495 555 2499
rect 559 2498 560 2499
rect 591 2499 597 2500
rect 591 2498 592 2499
rect 559 2496 592 2498
rect 559 2495 560 2496
rect 554 2494 560 2495
rect 591 2495 592 2496
rect 596 2495 597 2499
rect 591 2494 597 2495
rect 650 2499 656 2500
rect 650 2495 651 2499
rect 655 2498 656 2499
rect 695 2499 701 2500
rect 695 2498 696 2499
rect 655 2496 696 2498
rect 655 2495 656 2496
rect 650 2494 656 2495
rect 695 2495 696 2496
rect 700 2495 701 2499
rect 695 2494 701 2495
rect 754 2499 760 2500
rect 754 2495 755 2499
rect 759 2498 760 2499
rect 807 2499 813 2500
rect 807 2498 808 2499
rect 759 2496 808 2498
rect 759 2495 760 2496
rect 754 2494 760 2495
rect 807 2495 808 2496
rect 812 2495 813 2499
rect 807 2494 813 2495
rect 927 2499 933 2500
rect 927 2495 928 2499
rect 932 2498 933 2499
rect 998 2499 1004 2500
rect 998 2498 999 2499
rect 932 2496 999 2498
rect 932 2495 933 2496
rect 927 2494 933 2495
rect 998 2495 999 2496
rect 1003 2495 1004 2499
rect 998 2494 1004 2495
rect 1055 2499 1061 2500
rect 1055 2495 1056 2499
rect 1060 2498 1061 2499
rect 1127 2499 1133 2500
rect 1127 2498 1128 2499
rect 1060 2496 1128 2498
rect 1060 2495 1061 2496
rect 1055 2494 1061 2495
rect 1127 2495 1128 2496
rect 1132 2495 1133 2499
rect 1127 2494 1133 2495
rect 1183 2499 1189 2500
rect 1183 2495 1184 2499
rect 1188 2498 1189 2499
rect 1270 2499 1276 2500
rect 1270 2498 1271 2499
rect 1188 2496 1271 2498
rect 1188 2495 1189 2496
rect 1183 2494 1189 2495
rect 1270 2495 1271 2496
rect 1275 2495 1276 2499
rect 1270 2494 1276 2495
rect 1314 2499 1325 2500
rect 1314 2495 1315 2499
rect 1319 2495 1320 2499
rect 1324 2495 1325 2499
rect 1314 2494 1325 2495
rect 1378 2499 1384 2500
rect 1378 2495 1379 2499
rect 1383 2498 1384 2499
rect 1463 2499 1469 2500
rect 1463 2498 1464 2499
rect 1383 2496 1464 2498
rect 1383 2495 1384 2496
rect 1378 2494 1384 2495
rect 1463 2495 1464 2496
rect 1468 2495 1469 2499
rect 2186 2499 2192 2500
rect 2186 2498 2187 2499
rect 2181 2496 2187 2498
rect 1463 2494 1469 2495
rect 2186 2495 2187 2496
rect 2191 2495 2192 2499
rect 2274 2499 2280 2500
rect 2274 2498 2275 2499
rect 2269 2496 2275 2498
rect 2186 2494 2192 2495
rect 2274 2495 2275 2496
rect 2279 2495 2280 2499
rect 2370 2499 2376 2500
rect 2370 2498 2371 2499
rect 2365 2496 2371 2498
rect 2274 2494 2280 2495
rect 2370 2495 2371 2496
rect 2375 2495 2376 2499
rect 2466 2499 2472 2500
rect 2466 2498 2467 2499
rect 2461 2496 2467 2498
rect 2370 2494 2376 2495
rect 2466 2495 2467 2496
rect 2471 2495 2472 2499
rect 2466 2494 2472 2495
rect 2474 2499 2480 2500
rect 2474 2495 2475 2499
rect 2479 2498 2480 2499
rect 2658 2499 2664 2500
rect 2658 2498 2659 2499
rect 2479 2496 2513 2498
rect 2653 2496 2659 2498
rect 2479 2495 2480 2496
rect 2474 2494 2480 2495
rect 2658 2495 2659 2496
rect 2663 2495 2664 2499
rect 2754 2499 2760 2500
rect 2754 2498 2755 2499
rect 2749 2496 2755 2498
rect 2658 2494 2664 2495
rect 2754 2495 2755 2496
rect 2759 2495 2760 2499
rect 2850 2499 2856 2500
rect 2850 2498 2851 2499
rect 2845 2496 2851 2498
rect 2754 2494 2760 2495
rect 2850 2495 2851 2496
rect 2855 2495 2856 2499
rect 2946 2499 2952 2500
rect 2946 2498 2947 2499
rect 2941 2496 2947 2498
rect 2850 2494 2856 2495
rect 2946 2495 2947 2496
rect 2951 2495 2952 2499
rect 3042 2499 3048 2500
rect 3042 2498 3043 2499
rect 3037 2496 3043 2498
rect 2946 2494 2952 2495
rect 3042 2495 3043 2496
rect 3047 2495 3048 2499
rect 3042 2494 3048 2495
rect 3050 2499 3056 2500
rect 3050 2495 3051 2499
rect 3055 2498 3056 2499
rect 3055 2496 3097 2498
rect 3055 2495 3056 2496
rect 3050 2494 3056 2495
rect 334 2490 340 2491
rect 334 2486 335 2490
rect 339 2486 340 2490
rect 334 2485 340 2486
rect 414 2490 420 2491
rect 414 2486 415 2490
rect 419 2486 420 2490
rect 414 2485 420 2486
rect 502 2490 508 2491
rect 502 2486 503 2490
rect 507 2486 508 2490
rect 502 2485 508 2486
rect 598 2490 604 2491
rect 598 2486 599 2490
rect 603 2486 604 2490
rect 598 2485 604 2486
rect 702 2490 708 2491
rect 702 2486 703 2490
rect 707 2486 708 2490
rect 702 2485 708 2486
rect 814 2490 820 2491
rect 814 2486 815 2490
rect 819 2486 820 2490
rect 814 2485 820 2486
rect 934 2490 940 2491
rect 934 2486 935 2490
rect 939 2486 940 2490
rect 934 2485 940 2486
rect 1062 2490 1068 2491
rect 1062 2486 1063 2490
rect 1067 2486 1068 2490
rect 1062 2485 1068 2486
rect 1190 2490 1196 2491
rect 1190 2486 1191 2490
rect 1195 2486 1196 2490
rect 1190 2485 1196 2486
rect 1326 2490 1332 2491
rect 1326 2486 1327 2490
rect 1331 2486 1332 2490
rect 1326 2485 1332 2486
rect 1470 2490 1476 2491
rect 1470 2486 1471 2490
rect 1475 2486 1476 2490
rect 1470 2485 1476 2486
rect 1870 2488 1876 2489
rect 1870 2484 1871 2488
rect 1875 2484 1876 2488
rect 1870 2483 1876 2484
rect 3590 2488 3596 2489
rect 3590 2484 3591 2488
rect 3595 2484 3596 2488
rect 3590 2483 3596 2484
rect 110 2472 116 2473
rect 110 2468 111 2472
rect 115 2468 116 2472
rect 110 2467 116 2468
rect 1830 2472 1836 2473
rect 1830 2468 1831 2472
rect 1835 2468 1836 2472
rect 1830 2467 1836 2468
rect 2126 2470 2132 2471
rect 2126 2466 2127 2470
rect 2131 2466 2132 2470
rect 2126 2465 2132 2466
rect 2214 2470 2220 2471
rect 2214 2466 2215 2470
rect 2219 2466 2220 2470
rect 2214 2465 2220 2466
rect 2310 2470 2316 2471
rect 2310 2466 2311 2470
rect 2315 2466 2316 2470
rect 2310 2465 2316 2466
rect 2406 2470 2412 2471
rect 2406 2466 2407 2470
rect 2411 2466 2412 2470
rect 2406 2465 2412 2466
rect 2502 2470 2508 2471
rect 2502 2466 2503 2470
rect 2507 2466 2508 2470
rect 2502 2465 2508 2466
rect 2598 2470 2604 2471
rect 2598 2466 2599 2470
rect 2603 2466 2604 2470
rect 2598 2465 2604 2466
rect 2694 2470 2700 2471
rect 2694 2466 2695 2470
rect 2699 2466 2700 2470
rect 2694 2465 2700 2466
rect 2790 2470 2796 2471
rect 2790 2466 2791 2470
rect 2795 2466 2796 2470
rect 2790 2465 2796 2466
rect 2886 2470 2892 2471
rect 2886 2466 2887 2470
rect 2891 2466 2892 2470
rect 2886 2465 2892 2466
rect 2982 2470 2988 2471
rect 2982 2466 2983 2470
rect 2987 2466 2988 2470
rect 2982 2465 2988 2466
rect 3086 2470 3092 2471
rect 3086 2466 3087 2470
rect 3091 2466 3092 2470
rect 3086 2465 3092 2466
rect 386 2463 392 2464
rect 386 2459 387 2463
rect 391 2459 392 2463
rect 386 2458 392 2459
rect 466 2463 472 2464
rect 466 2459 467 2463
rect 471 2459 472 2463
rect 466 2458 472 2459
rect 554 2463 560 2464
rect 554 2459 555 2463
rect 559 2459 560 2463
rect 554 2458 560 2459
rect 650 2463 656 2464
rect 650 2459 651 2463
rect 655 2459 656 2463
rect 650 2458 656 2459
rect 754 2463 760 2464
rect 754 2459 755 2463
rect 759 2459 760 2463
rect 754 2458 760 2459
rect 886 2463 892 2464
rect 886 2459 887 2463
rect 891 2462 892 2463
rect 998 2463 1004 2464
rect 891 2460 945 2462
rect 891 2459 892 2460
rect 886 2458 892 2459
rect 998 2459 999 2463
rect 1003 2462 1004 2463
rect 1127 2463 1133 2464
rect 1003 2460 1073 2462
rect 1003 2459 1004 2460
rect 998 2458 1004 2459
rect 1127 2459 1128 2463
rect 1132 2462 1133 2463
rect 1378 2463 1384 2464
rect 1132 2460 1201 2462
rect 1132 2459 1133 2460
rect 1127 2458 1133 2459
rect 1378 2459 1379 2463
rect 1383 2459 1384 2463
rect 1378 2458 1384 2459
rect 1518 2463 1524 2464
rect 1518 2459 1519 2463
rect 1523 2459 1524 2463
rect 1518 2458 1524 2459
rect 2119 2459 2125 2460
rect 110 2455 116 2456
rect 110 2451 111 2455
rect 115 2451 116 2455
rect 1830 2455 1836 2456
rect 110 2450 116 2451
rect 326 2452 332 2453
rect 326 2448 327 2452
rect 331 2448 332 2452
rect 326 2447 332 2448
rect 406 2452 412 2453
rect 406 2448 407 2452
rect 411 2448 412 2452
rect 406 2447 412 2448
rect 494 2452 500 2453
rect 494 2448 495 2452
rect 499 2448 500 2452
rect 494 2447 500 2448
rect 590 2452 596 2453
rect 590 2448 591 2452
rect 595 2448 596 2452
rect 590 2447 596 2448
rect 694 2452 700 2453
rect 694 2448 695 2452
rect 699 2448 700 2452
rect 694 2447 700 2448
rect 806 2452 812 2453
rect 806 2448 807 2452
rect 811 2448 812 2452
rect 806 2447 812 2448
rect 926 2452 932 2453
rect 926 2448 927 2452
rect 931 2448 932 2452
rect 926 2447 932 2448
rect 1054 2452 1060 2453
rect 1054 2448 1055 2452
rect 1059 2448 1060 2452
rect 1054 2447 1060 2448
rect 1182 2452 1188 2453
rect 1182 2448 1183 2452
rect 1187 2448 1188 2452
rect 1182 2447 1188 2448
rect 1318 2452 1324 2453
rect 1318 2448 1319 2452
rect 1323 2448 1324 2452
rect 1318 2447 1324 2448
rect 1462 2452 1468 2453
rect 1462 2448 1463 2452
rect 1467 2448 1468 2452
rect 1830 2451 1831 2455
rect 1835 2451 1836 2455
rect 2119 2455 2120 2459
rect 2124 2458 2125 2459
rect 2178 2459 2184 2460
rect 2178 2458 2179 2459
rect 2124 2456 2179 2458
rect 2124 2455 2125 2456
rect 2119 2454 2125 2455
rect 2178 2455 2179 2456
rect 2183 2455 2184 2459
rect 2178 2454 2184 2455
rect 2186 2459 2192 2460
rect 2186 2455 2187 2459
rect 2191 2458 2192 2459
rect 2207 2459 2213 2460
rect 2207 2458 2208 2459
rect 2191 2456 2208 2458
rect 2191 2455 2192 2456
rect 2186 2454 2192 2455
rect 2207 2455 2208 2456
rect 2212 2455 2213 2459
rect 2207 2454 2213 2455
rect 2274 2459 2280 2460
rect 2274 2455 2275 2459
rect 2279 2458 2280 2459
rect 2303 2459 2309 2460
rect 2303 2458 2304 2459
rect 2279 2456 2304 2458
rect 2279 2455 2280 2456
rect 2274 2454 2280 2455
rect 2303 2455 2304 2456
rect 2308 2455 2309 2459
rect 2303 2454 2309 2455
rect 2370 2459 2376 2460
rect 2370 2455 2371 2459
rect 2375 2458 2376 2459
rect 2399 2459 2405 2460
rect 2399 2458 2400 2459
rect 2375 2456 2400 2458
rect 2375 2455 2376 2456
rect 2370 2454 2376 2455
rect 2399 2455 2400 2456
rect 2404 2455 2405 2459
rect 2399 2454 2405 2455
rect 2466 2459 2472 2460
rect 2466 2455 2467 2459
rect 2471 2458 2472 2459
rect 2495 2459 2501 2460
rect 2495 2458 2496 2459
rect 2471 2456 2496 2458
rect 2471 2455 2472 2456
rect 2466 2454 2472 2455
rect 2495 2455 2496 2456
rect 2500 2455 2501 2459
rect 2495 2454 2501 2455
rect 2591 2459 2597 2460
rect 2591 2455 2592 2459
rect 2596 2458 2597 2459
rect 2606 2459 2612 2460
rect 2606 2458 2607 2459
rect 2596 2456 2607 2458
rect 2596 2455 2597 2456
rect 2591 2454 2597 2455
rect 2606 2455 2607 2456
rect 2611 2455 2612 2459
rect 2606 2454 2612 2455
rect 2658 2459 2664 2460
rect 2658 2455 2659 2459
rect 2663 2458 2664 2459
rect 2687 2459 2693 2460
rect 2687 2458 2688 2459
rect 2663 2456 2688 2458
rect 2663 2455 2664 2456
rect 2658 2454 2664 2455
rect 2687 2455 2688 2456
rect 2692 2455 2693 2459
rect 2687 2454 2693 2455
rect 2754 2459 2760 2460
rect 2754 2455 2755 2459
rect 2759 2458 2760 2459
rect 2783 2459 2789 2460
rect 2783 2458 2784 2459
rect 2759 2456 2784 2458
rect 2759 2455 2760 2456
rect 2754 2454 2760 2455
rect 2783 2455 2784 2456
rect 2788 2455 2789 2459
rect 2783 2454 2789 2455
rect 2850 2459 2856 2460
rect 2850 2455 2851 2459
rect 2855 2458 2856 2459
rect 2879 2459 2885 2460
rect 2879 2458 2880 2459
rect 2855 2456 2880 2458
rect 2855 2455 2856 2456
rect 2850 2454 2856 2455
rect 2879 2455 2880 2456
rect 2884 2455 2885 2459
rect 2879 2454 2885 2455
rect 2946 2459 2952 2460
rect 2946 2455 2947 2459
rect 2951 2458 2952 2459
rect 2975 2459 2981 2460
rect 2975 2458 2976 2459
rect 2951 2456 2976 2458
rect 2951 2455 2952 2456
rect 2946 2454 2952 2455
rect 2975 2455 2976 2456
rect 2980 2455 2981 2459
rect 2975 2454 2981 2455
rect 3042 2459 3048 2460
rect 3042 2455 3043 2459
rect 3047 2458 3048 2459
rect 3079 2459 3085 2460
rect 3079 2458 3080 2459
rect 3047 2456 3080 2458
rect 3047 2455 3048 2456
rect 3042 2454 3048 2455
rect 3079 2455 3080 2456
rect 3084 2455 3085 2459
rect 3079 2454 3085 2455
rect 1830 2450 1836 2451
rect 1462 2447 1468 2448
rect 1895 2443 1901 2444
rect 1895 2439 1896 2443
rect 1900 2442 1901 2443
rect 1946 2443 1952 2444
rect 1946 2442 1947 2443
rect 1900 2440 1947 2442
rect 1900 2439 1901 2440
rect 1895 2438 1901 2439
rect 1946 2439 1947 2440
rect 1951 2439 1952 2443
rect 1946 2438 1952 2439
rect 1954 2443 1960 2444
rect 1954 2439 1955 2443
rect 1959 2442 1960 2443
rect 1983 2443 1989 2444
rect 1983 2442 1984 2443
rect 1959 2440 1984 2442
rect 1959 2439 1960 2440
rect 1954 2438 1960 2439
rect 1983 2439 1984 2440
rect 1988 2439 1989 2443
rect 1983 2438 1989 2439
rect 2042 2443 2048 2444
rect 2042 2439 2043 2443
rect 2047 2442 2048 2443
rect 2103 2443 2109 2444
rect 2103 2442 2104 2443
rect 2047 2440 2104 2442
rect 2047 2439 2048 2440
rect 2042 2438 2048 2439
rect 2103 2439 2104 2440
rect 2108 2439 2109 2443
rect 2103 2438 2109 2439
rect 2162 2443 2168 2444
rect 2162 2439 2163 2443
rect 2167 2442 2168 2443
rect 2239 2443 2245 2444
rect 2239 2442 2240 2443
rect 2167 2440 2240 2442
rect 2167 2439 2168 2440
rect 2162 2438 2168 2439
rect 2239 2439 2240 2440
rect 2244 2439 2245 2443
rect 2239 2438 2245 2439
rect 2298 2443 2304 2444
rect 2298 2439 2299 2443
rect 2303 2442 2304 2443
rect 2383 2443 2389 2444
rect 2383 2442 2384 2443
rect 2303 2440 2384 2442
rect 2303 2439 2304 2440
rect 2298 2438 2304 2439
rect 2383 2439 2384 2440
rect 2388 2439 2389 2443
rect 2383 2438 2389 2439
rect 2442 2443 2448 2444
rect 2442 2439 2443 2443
rect 2447 2442 2448 2443
rect 2527 2443 2533 2444
rect 2527 2442 2528 2443
rect 2447 2440 2528 2442
rect 2447 2439 2448 2440
rect 2442 2438 2448 2439
rect 2527 2439 2528 2440
rect 2532 2439 2533 2443
rect 2527 2438 2533 2439
rect 2663 2443 2669 2444
rect 2663 2439 2664 2443
rect 2668 2442 2669 2443
rect 2702 2443 2708 2444
rect 2702 2442 2703 2443
rect 2668 2440 2703 2442
rect 2668 2439 2669 2440
rect 2663 2438 2669 2439
rect 2702 2439 2703 2440
rect 2707 2439 2708 2443
rect 2702 2438 2708 2439
rect 2722 2443 2728 2444
rect 2722 2439 2723 2443
rect 2727 2442 2728 2443
rect 2799 2443 2805 2444
rect 2799 2442 2800 2443
rect 2727 2440 2800 2442
rect 2727 2439 2728 2440
rect 2722 2438 2728 2439
rect 2799 2439 2800 2440
rect 2804 2439 2805 2443
rect 2799 2438 2805 2439
rect 2858 2443 2864 2444
rect 2858 2439 2859 2443
rect 2863 2442 2864 2443
rect 2935 2443 2941 2444
rect 2935 2442 2936 2443
rect 2863 2440 2936 2442
rect 2863 2439 2864 2440
rect 2858 2438 2864 2439
rect 2935 2439 2936 2440
rect 2940 2439 2941 2443
rect 2935 2438 2941 2439
rect 2994 2443 3000 2444
rect 2994 2439 2995 2443
rect 2999 2442 3000 2443
rect 3071 2443 3077 2444
rect 3071 2442 3072 2443
rect 2999 2440 3072 2442
rect 2999 2439 3000 2440
rect 2994 2438 3000 2439
rect 3071 2439 3072 2440
rect 3076 2439 3077 2443
rect 3071 2438 3077 2439
rect 3130 2443 3136 2444
rect 3130 2439 3131 2443
rect 3135 2442 3136 2443
rect 3207 2443 3213 2444
rect 3207 2442 3208 2443
rect 3135 2440 3208 2442
rect 3135 2439 3136 2440
rect 3130 2438 3136 2439
rect 3207 2439 3208 2440
rect 3212 2439 3213 2443
rect 3207 2438 3213 2439
rect 798 2435 804 2436
rect 798 2431 799 2435
rect 803 2434 804 2435
rect 823 2435 829 2436
rect 823 2434 824 2435
rect 803 2432 824 2434
rect 803 2431 804 2432
rect 798 2430 804 2431
rect 823 2431 824 2432
rect 828 2431 829 2435
rect 823 2430 829 2431
rect 1902 2434 1908 2435
rect 1902 2430 1903 2434
rect 1907 2430 1908 2434
rect 1902 2429 1908 2430
rect 1990 2434 1996 2435
rect 1990 2430 1991 2434
rect 1995 2430 1996 2434
rect 1990 2429 1996 2430
rect 2110 2434 2116 2435
rect 2110 2430 2111 2434
rect 2115 2430 2116 2434
rect 2110 2429 2116 2430
rect 2246 2434 2252 2435
rect 2246 2430 2247 2434
rect 2251 2430 2252 2434
rect 2246 2429 2252 2430
rect 2390 2434 2396 2435
rect 2390 2430 2391 2434
rect 2395 2430 2396 2434
rect 2390 2429 2396 2430
rect 2534 2434 2540 2435
rect 2534 2430 2535 2434
rect 2539 2430 2540 2434
rect 2534 2429 2540 2430
rect 2670 2434 2676 2435
rect 2670 2430 2671 2434
rect 2675 2430 2676 2434
rect 2670 2429 2676 2430
rect 2806 2434 2812 2435
rect 2806 2430 2807 2434
rect 2811 2430 2812 2434
rect 2806 2429 2812 2430
rect 2942 2434 2948 2435
rect 2942 2430 2943 2434
rect 2947 2430 2948 2434
rect 2942 2429 2948 2430
rect 3078 2434 3084 2435
rect 3078 2430 3079 2434
rect 3083 2430 3084 2434
rect 3078 2429 3084 2430
rect 3214 2434 3220 2435
rect 3214 2430 3215 2434
rect 3219 2430 3220 2434
rect 3214 2429 3220 2430
rect 1870 2416 1876 2417
rect 1870 2412 1871 2416
rect 1875 2412 1876 2416
rect 1870 2411 1876 2412
rect 3590 2416 3596 2417
rect 3590 2412 3591 2416
rect 3595 2412 3596 2416
rect 3590 2411 3596 2412
rect 1954 2407 1960 2408
rect 1954 2403 1955 2407
rect 1959 2403 1960 2407
rect 1954 2402 1960 2403
rect 2042 2407 2048 2408
rect 2042 2403 2043 2407
rect 2047 2403 2048 2407
rect 2042 2402 2048 2403
rect 2162 2407 2168 2408
rect 2162 2403 2163 2407
rect 2167 2403 2168 2407
rect 2162 2402 2168 2403
rect 2298 2407 2304 2408
rect 2298 2403 2299 2407
rect 2303 2403 2304 2407
rect 2298 2402 2304 2403
rect 2442 2407 2448 2408
rect 2442 2403 2443 2407
rect 2447 2403 2448 2407
rect 2442 2402 2448 2403
rect 2542 2407 2548 2408
rect 2542 2403 2543 2407
rect 2547 2403 2548 2407
rect 2542 2402 2548 2403
rect 2722 2407 2728 2408
rect 2722 2403 2723 2407
rect 2727 2403 2728 2407
rect 2722 2402 2728 2403
rect 2858 2407 2864 2408
rect 2858 2403 2859 2407
rect 2863 2403 2864 2407
rect 2858 2402 2864 2403
rect 2994 2407 3000 2408
rect 2994 2403 2995 2407
rect 2999 2403 3000 2407
rect 2994 2402 3000 2403
rect 3130 2407 3136 2408
rect 3130 2403 3131 2407
rect 3135 2403 3136 2407
rect 3130 2402 3136 2403
rect 382 2400 388 2401
rect 110 2397 116 2398
rect 110 2393 111 2397
rect 115 2393 116 2397
rect 382 2396 383 2400
rect 387 2396 388 2400
rect 382 2395 388 2396
rect 462 2400 468 2401
rect 462 2396 463 2400
rect 467 2396 468 2400
rect 462 2395 468 2396
rect 542 2400 548 2401
rect 542 2396 543 2400
rect 547 2396 548 2400
rect 542 2395 548 2396
rect 622 2400 628 2401
rect 622 2396 623 2400
rect 627 2396 628 2400
rect 622 2395 628 2396
rect 702 2400 708 2401
rect 702 2396 703 2400
rect 707 2396 708 2400
rect 702 2395 708 2396
rect 782 2400 788 2401
rect 782 2396 783 2400
rect 787 2396 788 2400
rect 782 2395 788 2396
rect 862 2400 868 2401
rect 862 2396 863 2400
rect 867 2396 868 2400
rect 862 2395 868 2396
rect 942 2400 948 2401
rect 942 2396 943 2400
rect 947 2396 948 2400
rect 942 2395 948 2396
rect 1022 2400 1028 2401
rect 1022 2396 1023 2400
rect 1027 2396 1028 2400
rect 1022 2395 1028 2396
rect 1102 2400 1108 2401
rect 1102 2396 1103 2400
rect 1107 2396 1108 2400
rect 1102 2395 1108 2396
rect 1182 2400 1188 2401
rect 1182 2396 1183 2400
rect 1187 2396 1188 2400
rect 1182 2395 1188 2396
rect 1262 2400 1268 2401
rect 1262 2396 1263 2400
rect 1267 2396 1268 2400
rect 1262 2395 1268 2396
rect 1350 2400 1356 2401
rect 1350 2396 1351 2400
rect 1355 2396 1356 2400
rect 1350 2395 1356 2396
rect 1438 2400 1444 2401
rect 1438 2396 1439 2400
rect 1443 2396 1444 2400
rect 1438 2395 1444 2396
rect 1526 2400 1532 2401
rect 1526 2396 1527 2400
rect 1531 2396 1532 2400
rect 1870 2399 1876 2400
rect 1526 2395 1532 2396
rect 1830 2397 1836 2398
rect 110 2392 116 2393
rect 1830 2393 1831 2397
rect 1835 2393 1836 2397
rect 1870 2395 1871 2399
rect 1875 2395 1876 2399
rect 3590 2399 3596 2400
rect 1870 2394 1876 2395
rect 1894 2396 1900 2397
rect 1830 2392 1836 2393
rect 1894 2392 1895 2396
rect 1899 2392 1900 2396
rect 450 2391 456 2392
rect 450 2390 451 2391
rect 445 2388 451 2390
rect 450 2387 451 2388
rect 455 2387 456 2391
rect 530 2391 536 2392
rect 530 2390 531 2391
rect 525 2388 531 2390
rect 450 2386 456 2387
rect 530 2387 531 2388
rect 535 2387 536 2391
rect 610 2391 616 2392
rect 610 2390 611 2391
rect 605 2388 611 2390
rect 530 2386 536 2387
rect 610 2387 611 2388
rect 615 2387 616 2391
rect 690 2391 696 2392
rect 690 2390 691 2391
rect 685 2388 691 2390
rect 610 2386 616 2387
rect 690 2387 691 2388
rect 695 2387 696 2391
rect 770 2391 776 2392
rect 770 2390 771 2391
rect 765 2388 771 2390
rect 690 2386 696 2387
rect 770 2387 771 2388
rect 775 2387 776 2391
rect 930 2391 936 2392
rect 930 2390 931 2391
rect 845 2388 866 2390
rect 925 2388 931 2390
rect 770 2386 776 2387
rect 862 2387 868 2388
rect 862 2383 863 2387
rect 867 2383 868 2387
rect 930 2387 931 2388
rect 935 2387 936 2391
rect 1010 2391 1016 2392
rect 1010 2390 1011 2391
rect 1005 2388 1011 2390
rect 930 2386 936 2387
rect 1010 2387 1011 2388
rect 1015 2387 1016 2391
rect 1090 2391 1096 2392
rect 1090 2390 1091 2391
rect 1085 2388 1091 2390
rect 1010 2386 1016 2387
rect 1090 2387 1091 2388
rect 1095 2387 1096 2391
rect 1170 2391 1176 2392
rect 1170 2390 1171 2391
rect 1165 2388 1171 2390
rect 1090 2386 1096 2387
rect 1170 2387 1171 2388
rect 1175 2387 1176 2391
rect 1250 2391 1256 2392
rect 1250 2390 1251 2391
rect 1245 2388 1251 2390
rect 1170 2386 1176 2387
rect 1250 2387 1251 2388
rect 1255 2387 1256 2391
rect 1418 2391 1424 2392
rect 1418 2390 1419 2391
rect 1250 2386 1256 2387
rect 1270 2387 1276 2388
rect 862 2382 868 2383
rect 1270 2383 1271 2387
rect 1275 2386 1276 2387
rect 1280 2386 1282 2389
rect 1413 2388 1419 2390
rect 1418 2387 1419 2388
rect 1423 2387 1424 2391
rect 1418 2386 1424 2387
rect 1426 2391 1432 2392
rect 1426 2387 1427 2391
rect 1431 2390 1432 2391
rect 1506 2391 1512 2392
rect 1894 2391 1900 2392
rect 1982 2396 1988 2397
rect 1982 2392 1983 2396
rect 1987 2392 1988 2396
rect 1982 2391 1988 2392
rect 2102 2396 2108 2397
rect 2102 2392 2103 2396
rect 2107 2392 2108 2396
rect 2102 2391 2108 2392
rect 2238 2396 2244 2397
rect 2238 2392 2239 2396
rect 2243 2392 2244 2396
rect 2238 2391 2244 2392
rect 2382 2396 2388 2397
rect 2382 2392 2383 2396
rect 2387 2392 2388 2396
rect 2382 2391 2388 2392
rect 2526 2396 2532 2397
rect 2526 2392 2527 2396
rect 2531 2392 2532 2396
rect 2526 2391 2532 2392
rect 2662 2396 2668 2397
rect 2662 2392 2663 2396
rect 2667 2392 2668 2396
rect 2662 2391 2668 2392
rect 2798 2396 2804 2397
rect 2798 2392 2799 2396
rect 2803 2392 2804 2396
rect 2798 2391 2804 2392
rect 2934 2396 2940 2397
rect 2934 2392 2935 2396
rect 2939 2392 2940 2396
rect 2934 2391 2940 2392
rect 3070 2396 3076 2397
rect 3070 2392 3071 2396
rect 3075 2392 3076 2396
rect 3070 2391 3076 2392
rect 3206 2396 3212 2397
rect 3206 2392 3207 2396
rect 3211 2392 3212 2396
rect 3590 2395 3591 2399
rect 3595 2395 3596 2399
rect 3590 2394 3596 2395
rect 3206 2391 3212 2392
rect 1431 2388 1457 2390
rect 1431 2387 1432 2388
rect 1426 2386 1432 2387
rect 1506 2387 1507 2391
rect 1511 2390 1512 2391
rect 1511 2388 1545 2390
rect 1511 2387 1512 2388
rect 1506 2386 1512 2387
rect 1275 2384 1282 2386
rect 1275 2383 1276 2384
rect 1270 2382 1276 2383
rect 110 2380 116 2381
rect 110 2376 111 2380
rect 115 2376 116 2380
rect 110 2375 116 2376
rect 1830 2380 1836 2381
rect 1830 2376 1831 2380
rect 1835 2376 1836 2380
rect 1830 2375 1836 2376
rect 3138 2379 3144 2380
rect 3138 2375 3139 2379
rect 3143 2378 3144 2379
rect 3223 2379 3229 2380
rect 3223 2378 3224 2379
rect 3143 2376 3224 2378
rect 3143 2375 3144 2376
rect 3138 2374 3144 2375
rect 3223 2375 3224 2376
rect 3228 2375 3229 2379
rect 3223 2374 3229 2375
rect 390 2362 396 2363
rect 390 2358 391 2362
rect 395 2358 396 2362
rect 390 2357 396 2358
rect 470 2362 476 2363
rect 470 2358 471 2362
rect 475 2358 476 2362
rect 470 2357 476 2358
rect 550 2362 556 2363
rect 550 2358 551 2362
rect 555 2358 556 2362
rect 550 2357 556 2358
rect 630 2362 636 2363
rect 630 2358 631 2362
rect 635 2358 636 2362
rect 630 2357 636 2358
rect 710 2362 716 2363
rect 710 2358 711 2362
rect 715 2358 716 2362
rect 710 2357 716 2358
rect 790 2362 796 2363
rect 790 2358 791 2362
rect 795 2358 796 2362
rect 790 2357 796 2358
rect 870 2362 876 2363
rect 870 2358 871 2362
rect 875 2358 876 2362
rect 870 2357 876 2358
rect 950 2362 956 2363
rect 950 2358 951 2362
rect 955 2358 956 2362
rect 950 2357 956 2358
rect 1030 2362 1036 2363
rect 1030 2358 1031 2362
rect 1035 2358 1036 2362
rect 1030 2357 1036 2358
rect 1110 2362 1116 2363
rect 1110 2358 1111 2362
rect 1115 2358 1116 2362
rect 1110 2357 1116 2358
rect 1190 2362 1196 2363
rect 1190 2358 1191 2362
rect 1195 2358 1196 2362
rect 1190 2357 1196 2358
rect 1270 2362 1276 2363
rect 1270 2358 1271 2362
rect 1275 2358 1276 2362
rect 1270 2357 1276 2358
rect 1358 2362 1364 2363
rect 1358 2358 1359 2362
rect 1363 2358 1364 2362
rect 1358 2357 1364 2358
rect 1446 2362 1452 2363
rect 1446 2358 1447 2362
rect 1451 2358 1452 2362
rect 1446 2357 1452 2358
rect 1534 2362 1540 2363
rect 1534 2358 1535 2362
rect 1539 2358 1540 2362
rect 1534 2357 1540 2358
rect 383 2351 389 2352
rect 383 2347 384 2351
rect 388 2350 389 2351
rect 450 2351 456 2352
rect 388 2348 446 2350
rect 388 2347 389 2348
rect 383 2346 389 2347
rect 444 2342 446 2348
rect 450 2347 451 2351
rect 455 2350 456 2351
rect 463 2351 469 2352
rect 463 2350 464 2351
rect 455 2348 464 2350
rect 455 2347 456 2348
rect 450 2346 456 2347
rect 463 2347 464 2348
rect 468 2347 469 2351
rect 463 2346 469 2347
rect 530 2351 536 2352
rect 530 2347 531 2351
rect 535 2350 536 2351
rect 543 2351 549 2352
rect 543 2350 544 2351
rect 535 2348 544 2350
rect 535 2347 536 2348
rect 530 2346 536 2347
rect 543 2347 544 2348
rect 548 2347 549 2351
rect 543 2346 549 2347
rect 610 2351 616 2352
rect 610 2347 611 2351
rect 615 2350 616 2351
rect 623 2351 629 2352
rect 623 2350 624 2351
rect 615 2348 624 2350
rect 615 2347 616 2348
rect 610 2346 616 2347
rect 623 2347 624 2348
rect 628 2347 629 2351
rect 623 2346 629 2347
rect 690 2351 696 2352
rect 690 2347 691 2351
rect 695 2350 696 2351
rect 703 2351 709 2352
rect 703 2350 704 2351
rect 695 2348 704 2350
rect 695 2347 696 2348
rect 690 2346 696 2347
rect 703 2347 704 2348
rect 708 2347 709 2351
rect 703 2346 709 2347
rect 770 2351 776 2352
rect 770 2347 771 2351
rect 775 2350 776 2351
rect 783 2351 789 2352
rect 783 2350 784 2351
rect 775 2348 784 2350
rect 775 2347 776 2348
rect 770 2346 776 2347
rect 783 2347 784 2348
rect 788 2347 789 2351
rect 783 2346 789 2347
rect 862 2351 869 2352
rect 862 2347 863 2351
rect 868 2347 869 2351
rect 862 2346 869 2347
rect 930 2351 936 2352
rect 930 2347 931 2351
rect 935 2350 936 2351
rect 943 2351 949 2352
rect 943 2350 944 2351
rect 935 2348 944 2350
rect 935 2347 936 2348
rect 930 2346 936 2347
rect 943 2347 944 2348
rect 948 2347 949 2351
rect 943 2346 949 2347
rect 1010 2351 1016 2352
rect 1010 2347 1011 2351
rect 1015 2350 1016 2351
rect 1023 2351 1029 2352
rect 1023 2350 1024 2351
rect 1015 2348 1024 2350
rect 1015 2347 1016 2348
rect 1010 2346 1016 2347
rect 1023 2347 1024 2348
rect 1028 2347 1029 2351
rect 1023 2346 1029 2347
rect 1090 2351 1096 2352
rect 1090 2347 1091 2351
rect 1095 2350 1096 2351
rect 1103 2351 1109 2352
rect 1103 2350 1104 2351
rect 1095 2348 1104 2350
rect 1095 2347 1096 2348
rect 1090 2346 1096 2347
rect 1103 2347 1104 2348
rect 1108 2347 1109 2351
rect 1103 2346 1109 2347
rect 1170 2351 1176 2352
rect 1170 2347 1171 2351
rect 1175 2350 1176 2351
rect 1183 2351 1189 2352
rect 1183 2350 1184 2351
rect 1175 2348 1184 2350
rect 1175 2347 1176 2348
rect 1170 2346 1176 2347
rect 1183 2347 1184 2348
rect 1188 2347 1189 2351
rect 1183 2346 1189 2347
rect 1250 2351 1256 2352
rect 1250 2347 1251 2351
rect 1255 2350 1256 2351
rect 1263 2351 1269 2352
rect 1263 2350 1264 2351
rect 1255 2348 1264 2350
rect 1255 2347 1256 2348
rect 1250 2346 1256 2347
rect 1263 2347 1264 2348
rect 1268 2347 1269 2351
rect 1263 2346 1269 2347
rect 1351 2351 1357 2352
rect 1351 2347 1352 2351
rect 1356 2350 1357 2351
rect 1426 2351 1432 2352
rect 1426 2350 1427 2351
rect 1356 2348 1427 2350
rect 1356 2347 1357 2348
rect 1351 2346 1357 2347
rect 1426 2347 1427 2348
rect 1431 2347 1432 2351
rect 1426 2346 1432 2347
rect 1439 2351 1445 2352
rect 1439 2347 1440 2351
rect 1444 2350 1445 2351
rect 1506 2351 1512 2352
rect 1506 2350 1507 2351
rect 1444 2348 1507 2350
rect 1444 2347 1445 2348
rect 1439 2346 1445 2347
rect 1506 2347 1507 2348
rect 1511 2347 1512 2351
rect 1506 2346 1512 2347
rect 1518 2351 1524 2352
rect 1518 2347 1519 2351
rect 1523 2350 1524 2351
rect 1527 2351 1533 2352
rect 1527 2350 1528 2351
rect 1523 2348 1528 2350
rect 1523 2347 1524 2348
rect 1518 2346 1524 2347
rect 1527 2347 1528 2348
rect 1532 2347 1533 2351
rect 1527 2346 1533 2347
rect 1894 2344 1900 2345
rect 798 2343 804 2344
rect 798 2342 799 2343
rect 444 2340 799 2342
rect 798 2339 799 2340
rect 803 2339 804 2343
rect 1870 2341 1876 2342
rect 798 2338 804 2339
rect 1399 2339 1405 2340
rect 1399 2335 1400 2339
rect 1404 2338 1405 2339
rect 1418 2339 1424 2340
rect 1418 2338 1419 2339
rect 1404 2336 1419 2338
rect 1404 2335 1405 2336
rect 1399 2334 1405 2335
rect 1418 2335 1419 2336
rect 1423 2335 1424 2339
rect 1418 2334 1424 2335
rect 1458 2339 1464 2340
rect 1458 2335 1459 2339
rect 1463 2338 1464 2339
rect 1479 2339 1485 2340
rect 1479 2338 1480 2339
rect 1463 2336 1480 2338
rect 1463 2335 1464 2336
rect 1458 2334 1464 2335
rect 1479 2335 1480 2336
rect 1484 2335 1485 2339
rect 1479 2334 1485 2335
rect 1558 2339 1565 2340
rect 1558 2335 1559 2339
rect 1564 2335 1565 2339
rect 1558 2334 1565 2335
rect 1618 2339 1624 2340
rect 1618 2335 1619 2339
rect 1623 2338 1624 2339
rect 1639 2339 1645 2340
rect 1639 2338 1640 2339
rect 1623 2336 1640 2338
rect 1623 2335 1624 2336
rect 1618 2334 1624 2335
rect 1639 2335 1640 2336
rect 1644 2335 1645 2339
rect 1870 2337 1871 2341
rect 1875 2337 1876 2341
rect 1894 2340 1895 2344
rect 1899 2340 1900 2344
rect 1894 2339 1900 2340
rect 2014 2344 2020 2345
rect 2014 2340 2015 2344
rect 2019 2340 2020 2344
rect 2014 2339 2020 2340
rect 2174 2344 2180 2345
rect 2174 2340 2175 2344
rect 2179 2340 2180 2344
rect 2174 2339 2180 2340
rect 2342 2344 2348 2345
rect 2342 2340 2343 2344
rect 2347 2340 2348 2344
rect 2342 2339 2348 2340
rect 2510 2344 2516 2345
rect 2510 2340 2511 2344
rect 2515 2340 2516 2344
rect 2510 2339 2516 2340
rect 2670 2344 2676 2345
rect 2670 2340 2671 2344
rect 2675 2340 2676 2344
rect 2670 2339 2676 2340
rect 2822 2344 2828 2345
rect 2822 2340 2823 2344
rect 2827 2340 2828 2344
rect 2822 2339 2828 2340
rect 2958 2344 2964 2345
rect 2958 2340 2959 2344
rect 2963 2340 2964 2344
rect 2958 2339 2964 2340
rect 3078 2344 3084 2345
rect 3078 2340 3079 2344
rect 3083 2340 3084 2344
rect 3078 2339 3084 2340
rect 3190 2344 3196 2345
rect 3190 2340 3191 2344
rect 3195 2340 3196 2344
rect 3190 2339 3196 2340
rect 3302 2344 3308 2345
rect 3302 2340 3303 2344
rect 3307 2340 3308 2344
rect 3302 2339 3308 2340
rect 3414 2344 3420 2345
rect 3414 2340 3415 2344
rect 3419 2340 3420 2344
rect 3414 2339 3420 2340
rect 3502 2344 3508 2345
rect 3502 2340 3503 2344
rect 3507 2340 3508 2344
rect 3502 2339 3508 2340
rect 3590 2341 3596 2342
rect 1870 2336 1876 2337
rect 3590 2337 3591 2341
rect 3595 2337 3596 2341
rect 3590 2336 3596 2337
rect 1639 2334 1645 2335
rect 1962 2335 1968 2336
rect 1962 2334 1963 2335
rect 1957 2332 1963 2334
rect 1962 2331 1963 2332
rect 1967 2331 1968 2335
rect 2098 2335 2104 2336
rect 2098 2334 2099 2335
rect 2077 2332 2099 2334
rect 1406 2330 1412 2331
rect 1406 2326 1407 2330
rect 1411 2326 1412 2330
rect 1406 2325 1412 2326
rect 1486 2330 1492 2331
rect 1486 2326 1487 2330
rect 1491 2326 1492 2330
rect 1486 2325 1492 2326
rect 1566 2330 1572 2331
rect 1566 2326 1567 2330
rect 1571 2326 1572 2330
rect 1566 2325 1572 2326
rect 1646 2330 1652 2331
rect 1962 2330 1968 2331
rect 2098 2331 2099 2332
rect 2103 2331 2104 2335
rect 2242 2335 2248 2336
rect 2242 2334 2243 2335
rect 2237 2332 2243 2334
rect 2098 2330 2104 2331
rect 2242 2331 2243 2332
rect 2247 2331 2248 2335
rect 2434 2335 2440 2336
rect 2434 2334 2435 2335
rect 2405 2332 2435 2334
rect 2242 2330 2248 2331
rect 2434 2331 2435 2332
rect 2439 2331 2440 2335
rect 2434 2330 2440 2331
rect 2458 2335 2464 2336
rect 2458 2331 2459 2335
rect 2463 2334 2464 2335
rect 2754 2335 2760 2336
rect 2754 2334 2755 2335
rect 2463 2332 2529 2334
rect 2733 2332 2755 2334
rect 2463 2331 2464 2332
rect 2458 2330 2464 2331
rect 2754 2331 2755 2332
rect 2759 2331 2760 2335
rect 2890 2335 2896 2336
rect 2890 2334 2891 2335
rect 2885 2332 2891 2334
rect 2754 2330 2760 2331
rect 2890 2331 2891 2332
rect 2895 2331 2896 2335
rect 3030 2335 3036 2336
rect 3030 2334 3031 2335
rect 3021 2332 3031 2334
rect 2890 2330 2896 2331
rect 3030 2331 3031 2332
rect 3035 2331 3036 2335
rect 3146 2335 3152 2336
rect 3146 2334 3147 2335
rect 3141 2332 3147 2334
rect 3030 2330 3036 2331
rect 3146 2331 3147 2332
rect 3151 2331 3152 2335
rect 3262 2335 3268 2336
rect 3262 2334 3263 2335
rect 3253 2332 3263 2334
rect 3146 2330 3152 2331
rect 3262 2331 3263 2332
rect 3267 2331 3268 2335
rect 3370 2335 3376 2336
rect 3370 2334 3371 2335
rect 3365 2332 3371 2334
rect 3262 2330 3268 2331
rect 3370 2331 3371 2332
rect 3375 2331 3376 2335
rect 3482 2335 3488 2336
rect 3482 2334 3483 2335
rect 3477 2332 3483 2334
rect 3370 2330 3376 2331
rect 3482 2331 3483 2332
rect 3487 2331 3488 2335
rect 3482 2330 3488 2331
rect 3495 2335 3501 2336
rect 3495 2331 3496 2335
rect 3500 2334 3501 2335
rect 3500 2332 3521 2334
rect 3500 2331 3501 2332
rect 3495 2330 3501 2331
rect 1646 2326 1647 2330
rect 1651 2326 1652 2330
rect 1646 2325 1652 2326
rect 1870 2324 1876 2325
rect 1870 2320 1871 2324
rect 1875 2320 1876 2324
rect 1870 2319 1876 2320
rect 3590 2324 3596 2325
rect 3590 2320 3591 2324
rect 3595 2320 3596 2324
rect 3590 2319 3596 2320
rect 110 2312 116 2313
rect 110 2308 111 2312
rect 115 2308 116 2312
rect 110 2307 116 2308
rect 1830 2312 1836 2313
rect 1830 2308 1831 2312
rect 1835 2308 1836 2312
rect 1830 2307 1836 2308
rect 1902 2306 1908 2307
rect 1458 2303 1464 2304
rect 1458 2299 1459 2303
rect 1463 2299 1464 2303
rect 1558 2303 1564 2304
rect 1558 2302 1559 2303
rect 1541 2300 1559 2302
rect 1458 2298 1464 2299
rect 1558 2299 1559 2300
rect 1563 2299 1564 2303
rect 1558 2298 1564 2299
rect 1618 2303 1624 2304
rect 1618 2299 1619 2303
rect 1623 2299 1624 2303
rect 1902 2302 1903 2306
rect 1907 2302 1908 2306
rect 1902 2301 1908 2302
rect 2022 2306 2028 2307
rect 2022 2302 2023 2306
rect 2027 2302 2028 2306
rect 2022 2301 2028 2302
rect 2182 2306 2188 2307
rect 2182 2302 2183 2306
rect 2187 2302 2188 2306
rect 2182 2301 2188 2302
rect 2350 2306 2356 2307
rect 2350 2302 2351 2306
rect 2355 2302 2356 2306
rect 2350 2301 2356 2302
rect 2518 2306 2524 2307
rect 2518 2302 2519 2306
rect 2523 2302 2524 2306
rect 2518 2301 2524 2302
rect 2678 2306 2684 2307
rect 2678 2302 2679 2306
rect 2683 2302 2684 2306
rect 2678 2301 2684 2302
rect 2830 2306 2836 2307
rect 2830 2302 2831 2306
rect 2835 2302 2836 2306
rect 2830 2301 2836 2302
rect 2966 2306 2972 2307
rect 2966 2302 2967 2306
rect 2971 2302 2972 2306
rect 2966 2301 2972 2302
rect 3086 2306 3092 2307
rect 3086 2302 3087 2306
rect 3091 2302 3092 2306
rect 3086 2301 3092 2302
rect 3198 2306 3204 2307
rect 3198 2302 3199 2306
rect 3203 2302 3204 2306
rect 3198 2301 3204 2302
rect 3310 2306 3316 2307
rect 3310 2302 3311 2306
rect 3315 2302 3316 2306
rect 3310 2301 3316 2302
rect 3422 2306 3428 2307
rect 3422 2302 3423 2306
rect 3427 2302 3428 2306
rect 3422 2301 3428 2302
rect 3510 2306 3516 2307
rect 3510 2302 3511 2306
rect 3515 2302 3516 2306
rect 3510 2301 3516 2302
rect 1618 2298 1624 2299
rect 110 2295 116 2296
rect 110 2291 111 2295
rect 115 2291 116 2295
rect 1830 2295 1836 2296
rect 110 2290 116 2291
rect 1398 2292 1404 2293
rect 1398 2288 1399 2292
rect 1403 2288 1404 2292
rect 1398 2287 1404 2288
rect 1478 2292 1484 2293
rect 1478 2288 1479 2292
rect 1483 2288 1484 2292
rect 1478 2287 1484 2288
rect 1558 2292 1564 2293
rect 1558 2288 1559 2292
rect 1563 2288 1564 2292
rect 1558 2287 1564 2288
rect 1638 2292 1644 2293
rect 1638 2288 1639 2292
rect 1643 2288 1644 2292
rect 1830 2291 1831 2295
rect 1835 2291 1836 2295
rect 1830 2290 1836 2291
rect 1895 2295 1901 2296
rect 1895 2291 1896 2295
rect 1900 2294 1901 2295
rect 1910 2295 1916 2296
rect 1910 2294 1911 2295
rect 1900 2292 1911 2294
rect 1900 2291 1901 2292
rect 1895 2290 1901 2291
rect 1910 2291 1911 2292
rect 1915 2291 1916 2295
rect 1910 2290 1916 2291
rect 1962 2295 1968 2296
rect 1962 2291 1963 2295
rect 1967 2294 1968 2295
rect 2015 2295 2021 2296
rect 2015 2294 2016 2295
rect 1967 2292 2016 2294
rect 1967 2291 1968 2292
rect 1962 2290 1968 2291
rect 2015 2291 2016 2292
rect 2020 2291 2021 2295
rect 2015 2290 2021 2291
rect 2098 2295 2104 2296
rect 2098 2291 2099 2295
rect 2103 2294 2104 2295
rect 2175 2295 2181 2296
rect 2175 2294 2176 2295
rect 2103 2292 2176 2294
rect 2103 2291 2104 2292
rect 2098 2290 2104 2291
rect 2175 2291 2176 2292
rect 2180 2291 2181 2295
rect 2175 2290 2181 2291
rect 2242 2295 2248 2296
rect 2242 2291 2243 2295
rect 2247 2294 2248 2295
rect 2343 2295 2349 2296
rect 2343 2294 2344 2295
rect 2247 2292 2344 2294
rect 2247 2291 2248 2292
rect 2242 2290 2248 2291
rect 2343 2291 2344 2292
rect 2348 2291 2349 2295
rect 2343 2290 2349 2291
rect 2434 2295 2440 2296
rect 2434 2291 2435 2295
rect 2439 2294 2440 2295
rect 2511 2295 2517 2296
rect 2511 2294 2512 2295
rect 2439 2292 2512 2294
rect 2439 2291 2440 2292
rect 2434 2290 2440 2291
rect 2511 2291 2512 2292
rect 2516 2291 2517 2295
rect 2511 2290 2517 2291
rect 2671 2295 2677 2296
rect 2671 2291 2672 2295
rect 2676 2294 2677 2295
rect 2686 2295 2692 2296
rect 2686 2294 2687 2295
rect 2676 2292 2687 2294
rect 2676 2291 2677 2292
rect 2671 2290 2677 2291
rect 2686 2291 2687 2292
rect 2691 2291 2692 2295
rect 2686 2290 2692 2291
rect 2754 2295 2760 2296
rect 2754 2291 2755 2295
rect 2759 2294 2760 2295
rect 2823 2295 2829 2296
rect 2823 2294 2824 2295
rect 2759 2292 2824 2294
rect 2759 2291 2760 2292
rect 2754 2290 2760 2291
rect 2823 2291 2824 2292
rect 2828 2291 2829 2295
rect 2823 2290 2829 2291
rect 2890 2295 2896 2296
rect 2890 2291 2891 2295
rect 2895 2294 2896 2295
rect 2959 2295 2965 2296
rect 2959 2294 2960 2295
rect 2895 2292 2960 2294
rect 2895 2291 2896 2292
rect 2890 2290 2896 2291
rect 2959 2291 2960 2292
rect 2964 2291 2965 2295
rect 2959 2290 2965 2291
rect 3030 2295 3036 2296
rect 3030 2291 3031 2295
rect 3035 2294 3036 2295
rect 3079 2295 3085 2296
rect 3079 2294 3080 2295
rect 3035 2292 3080 2294
rect 3035 2291 3036 2292
rect 3030 2290 3036 2291
rect 3079 2291 3080 2292
rect 3084 2291 3085 2295
rect 3146 2295 3152 2296
rect 3079 2290 3085 2291
rect 3087 2291 3093 2292
rect 1638 2287 1644 2288
rect 3087 2287 3088 2291
rect 3092 2290 3093 2291
rect 3146 2291 3147 2295
rect 3151 2294 3152 2295
rect 3191 2295 3197 2296
rect 3191 2294 3192 2295
rect 3151 2292 3192 2294
rect 3151 2291 3152 2292
rect 3146 2290 3152 2291
rect 3191 2291 3192 2292
rect 3196 2291 3197 2295
rect 3191 2290 3197 2291
rect 3262 2295 3268 2296
rect 3262 2291 3263 2295
rect 3267 2294 3268 2295
rect 3303 2295 3309 2296
rect 3303 2294 3304 2295
rect 3267 2292 3304 2294
rect 3267 2291 3268 2292
rect 3262 2290 3268 2291
rect 3303 2291 3304 2292
rect 3308 2291 3309 2295
rect 3303 2290 3309 2291
rect 3370 2295 3376 2296
rect 3370 2291 3371 2295
rect 3375 2294 3376 2295
rect 3415 2295 3421 2296
rect 3415 2294 3416 2295
rect 3375 2292 3416 2294
rect 3375 2291 3376 2292
rect 3370 2290 3376 2291
rect 3415 2291 3416 2292
rect 3420 2291 3421 2295
rect 3415 2290 3421 2291
rect 3482 2295 3488 2296
rect 3482 2291 3483 2295
rect 3487 2294 3488 2295
rect 3503 2295 3509 2296
rect 3503 2294 3504 2295
rect 3487 2292 3504 2294
rect 3487 2291 3488 2292
rect 3482 2290 3488 2291
rect 3503 2291 3504 2292
rect 3508 2291 3509 2295
rect 3503 2290 3509 2291
rect 3092 2288 3141 2290
rect 3092 2287 3093 2288
rect 3087 2286 3093 2287
rect 3139 2286 3141 2288
rect 3240 2288 3258 2290
rect 3240 2286 3242 2288
rect 3139 2284 3242 2286
rect 3256 2286 3258 2288
rect 3342 2287 3348 2288
rect 3342 2286 3343 2287
rect 3256 2284 3343 2286
rect 1895 2283 1901 2284
rect 1895 2279 1896 2283
rect 1900 2282 1901 2283
rect 1962 2283 1968 2284
rect 1962 2282 1963 2283
rect 1900 2280 1963 2282
rect 1900 2279 1901 2280
rect 1895 2278 1901 2279
rect 1962 2279 1963 2280
rect 1967 2279 1968 2283
rect 1962 2278 1968 2279
rect 2023 2283 2029 2284
rect 2023 2279 2024 2283
rect 2028 2282 2029 2283
rect 2103 2283 2109 2284
rect 2103 2282 2104 2283
rect 2028 2280 2104 2282
rect 2028 2279 2029 2280
rect 2023 2278 2029 2279
rect 2103 2279 2104 2280
rect 2108 2279 2109 2283
rect 2103 2278 2109 2279
rect 2175 2283 2181 2284
rect 2175 2279 2176 2283
rect 2180 2282 2181 2283
rect 2247 2283 2253 2284
rect 2247 2282 2248 2283
rect 2180 2280 2248 2282
rect 2180 2279 2181 2280
rect 2175 2278 2181 2279
rect 2247 2279 2248 2280
rect 2252 2279 2253 2283
rect 2247 2278 2253 2279
rect 2359 2283 2365 2284
rect 2359 2279 2360 2283
rect 2364 2282 2365 2283
rect 2374 2283 2380 2284
rect 2374 2282 2375 2283
rect 2364 2280 2375 2282
rect 2364 2279 2365 2280
rect 2359 2278 2365 2279
rect 2374 2279 2375 2280
rect 2379 2279 2380 2283
rect 2374 2278 2380 2279
rect 2478 2283 2484 2284
rect 2478 2279 2479 2283
rect 2483 2282 2484 2283
rect 2567 2283 2573 2284
rect 2567 2282 2568 2283
rect 2483 2280 2568 2282
rect 2483 2279 2484 2280
rect 2478 2278 2484 2279
rect 2567 2279 2568 2280
rect 2572 2279 2573 2283
rect 2567 2278 2573 2279
rect 2626 2283 2632 2284
rect 2626 2279 2627 2283
rect 2631 2282 2632 2283
rect 2783 2283 2789 2284
rect 2783 2282 2784 2283
rect 2631 2280 2784 2282
rect 2631 2279 2632 2280
rect 2626 2278 2632 2279
rect 2783 2279 2784 2280
rect 2788 2279 2789 2283
rect 2783 2278 2789 2279
rect 3015 2283 3021 2284
rect 3015 2279 3016 2283
rect 3020 2282 3021 2283
rect 3074 2283 3080 2284
rect 3020 2280 3070 2282
rect 3020 2279 3021 2280
rect 3015 2278 3021 2279
rect 1578 2275 1584 2276
rect 1578 2271 1579 2275
rect 1583 2274 1584 2275
rect 1655 2275 1661 2276
rect 1655 2274 1656 2275
rect 1583 2272 1656 2274
rect 1583 2271 1584 2272
rect 1578 2270 1584 2271
rect 1655 2271 1656 2272
rect 1660 2271 1661 2275
rect 1655 2270 1661 2271
rect 1902 2274 1908 2275
rect 1902 2270 1903 2274
rect 1907 2270 1908 2274
rect 1902 2269 1908 2270
rect 2030 2274 2036 2275
rect 2030 2270 2031 2274
rect 2035 2270 2036 2274
rect 2030 2269 2036 2270
rect 2182 2274 2188 2275
rect 2182 2270 2183 2274
rect 2187 2270 2188 2274
rect 2182 2269 2188 2270
rect 2366 2274 2372 2275
rect 2366 2270 2367 2274
rect 2371 2270 2372 2274
rect 2366 2269 2372 2270
rect 2574 2274 2580 2275
rect 2574 2270 2575 2274
rect 2579 2270 2580 2274
rect 2574 2269 2580 2270
rect 2790 2274 2796 2275
rect 2790 2270 2791 2274
rect 2795 2270 2796 2274
rect 2790 2269 2796 2270
rect 3022 2274 3028 2275
rect 3022 2270 3023 2274
rect 3027 2270 3028 2274
rect 3068 2274 3070 2280
rect 3074 2279 3075 2283
rect 3079 2282 3080 2283
rect 3247 2283 3253 2284
rect 3247 2282 3248 2283
rect 3079 2280 3248 2282
rect 3079 2279 3080 2280
rect 3074 2278 3080 2279
rect 3247 2279 3248 2280
rect 3252 2279 3253 2283
rect 3342 2283 3343 2284
rect 3347 2283 3348 2287
rect 3342 2282 3348 2283
rect 3487 2283 3493 2284
rect 3247 2278 3253 2279
rect 3487 2279 3488 2283
rect 3492 2282 3493 2283
rect 3495 2283 3501 2284
rect 3495 2282 3496 2283
rect 3492 2280 3496 2282
rect 3492 2279 3493 2280
rect 3487 2278 3493 2279
rect 3495 2279 3496 2280
rect 3500 2279 3501 2283
rect 3495 2278 3501 2279
rect 3087 2275 3093 2276
rect 3087 2274 3088 2275
rect 3068 2272 3088 2274
rect 3087 2271 3088 2272
rect 3092 2271 3093 2275
rect 3087 2270 3093 2271
rect 3254 2274 3260 2275
rect 3254 2270 3255 2274
rect 3259 2270 3260 2274
rect 3022 2269 3028 2270
rect 3254 2269 3260 2270
rect 3494 2274 3500 2275
rect 3494 2270 3495 2274
rect 3499 2270 3500 2274
rect 3494 2269 3500 2270
rect 1870 2256 1876 2257
rect 1870 2252 1871 2256
rect 1875 2252 1876 2256
rect 1870 2251 1876 2252
rect 3590 2256 3596 2257
rect 3590 2252 3591 2256
rect 3595 2252 3596 2256
rect 3590 2251 3596 2252
rect 1910 2247 1916 2248
rect 1910 2243 1911 2247
rect 1915 2243 1916 2247
rect 1910 2242 1916 2243
rect 1962 2247 1968 2248
rect 1962 2243 1963 2247
rect 1967 2246 1968 2247
rect 2103 2247 2109 2248
rect 1967 2244 2041 2246
rect 1967 2243 1968 2244
rect 1962 2242 1968 2243
rect 2103 2243 2104 2247
rect 2108 2246 2109 2247
rect 2247 2247 2253 2248
rect 2108 2244 2193 2246
rect 2108 2243 2109 2244
rect 2103 2242 2109 2243
rect 2247 2243 2248 2247
rect 2252 2246 2253 2247
rect 2626 2247 2632 2248
rect 2252 2244 2377 2246
rect 2252 2243 2253 2244
rect 2247 2242 2253 2243
rect 2626 2243 2627 2247
rect 2631 2243 2632 2247
rect 2626 2242 2632 2243
rect 3074 2247 3080 2248
rect 3074 2243 3075 2247
rect 3079 2243 3080 2247
rect 3334 2247 3340 2248
rect 3334 2246 3335 2247
rect 3309 2244 3335 2246
rect 3074 2242 3080 2243
rect 3334 2243 3335 2244
rect 3339 2243 3340 2247
rect 3334 2242 3340 2243
rect 3342 2247 3348 2248
rect 3342 2243 3343 2247
rect 3347 2246 3348 2247
rect 3347 2244 3505 2246
rect 3347 2243 3348 2244
rect 3342 2242 3348 2243
rect 134 2240 140 2241
rect 110 2237 116 2238
rect 110 2233 111 2237
rect 115 2233 116 2237
rect 134 2236 135 2240
rect 139 2236 140 2240
rect 134 2235 140 2236
rect 214 2240 220 2241
rect 214 2236 215 2240
rect 219 2236 220 2240
rect 214 2235 220 2236
rect 294 2240 300 2241
rect 294 2236 295 2240
rect 299 2236 300 2240
rect 294 2235 300 2236
rect 382 2240 388 2241
rect 382 2236 383 2240
rect 387 2236 388 2240
rect 382 2235 388 2236
rect 518 2240 524 2241
rect 518 2236 519 2240
rect 523 2236 524 2240
rect 518 2235 524 2236
rect 670 2240 676 2241
rect 670 2236 671 2240
rect 675 2236 676 2240
rect 670 2235 676 2236
rect 830 2240 836 2241
rect 830 2236 831 2240
rect 835 2236 836 2240
rect 830 2235 836 2236
rect 998 2240 1004 2241
rect 998 2236 999 2240
rect 1003 2236 1004 2240
rect 998 2235 1004 2236
rect 1158 2240 1164 2241
rect 1158 2236 1159 2240
rect 1163 2236 1164 2240
rect 1158 2235 1164 2236
rect 1310 2240 1316 2241
rect 1310 2236 1311 2240
rect 1315 2236 1316 2240
rect 1310 2235 1316 2236
rect 1454 2240 1460 2241
rect 1454 2236 1455 2240
rect 1459 2236 1460 2240
rect 1454 2235 1460 2236
rect 1606 2240 1612 2241
rect 1606 2236 1607 2240
rect 1611 2236 1612 2240
rect 1606 2235 1612 2236
rect 1742 2240 1748 2241
rect 1742 2236 1743 2240
rect 1747 2236 1748 2240
rect 1870 2239 1876 2240
rect 1742 2235 1748 2236
rect 1830 2237 1836 2238
rect 110 2232 116 2233
rect 1830 2233 1831 2237
rect 1835 2233 1836 2237
rect 1870 2235 1871 2239
rect 1875 2235 1876 2239
rect 3590 2239 3596 2240
rect 1870 2234 1876 2235
rect 1894 2236 1900 2237
rect 1830 2232 1836 2233
rect 1894 2232 1895 2236
rect 1899 2232 1900 2236
rect 202 2231 208 2232
rect 202 2230 203 2231
rect 197 2228 203 2230
rect 202 2227 203 2228
rect 207 2227 208 2231
rect 282 2231 288 2232
rect 282 2230 283 2231
rect 277 2228 283 2230
rect 202 2226 208 2227
rect 282 2227 283 2228
rect 287 2227 288 2231
rect 362 2231 368 2232
rect 362 2230 363 2231
rect 357 2228 363 2230
rect 282 2226 288 2227
rect 362 2227 363 2228
rect 367 2227 368 2231
rect 458 2231 464 2232
rect 458 2230 459 2231
rect 445 2228 459 2230
rect 362 2226 368 2227
rect 458 2227 459 2228
rect 463 2227 464 2231
rect 586 2231 592 2232
rect 586 2230 587 2231
rect 581 2228 587 2230
rect 458 2226 464 2227
rect 586 2227 587 2228
rect 591 2227 592 2231
rect 754 2231 760 2232
rect 754 2230 755 2231
rect 733 2228 755 2230
rect 586 2226 592 2227
rect 754 2227 755 2228
rect 759 2227 760 2231
rect 922 2231 928 2232
rect 922 2230 923 2231
rect 893 2228 923 2230
rect 754 2226 760 2227
rect 922 2227 923 2228
rect 927 2227 928 2231
rect 1234 2231 1240 2232
rect 1234 2230 1235 2231
rect 1000 2228 1017 2230
rect 1221 2228 1235 2230
rect 922 2226 928 2227
rect 998 2227 1004 2228
rect 998 2223 999 2227
rect 1003 2223 1004 2227
rect 1234 2227 1235 2228
rect 1239 2227 1240 2231
rect 1378 2231 1384 2232
rect 1378 2230 1379 2231
rect 1373 2228 1379 2230
rect 1234 2226 1240 2227
rect 1378 2227 1379 2228
rect 1383 2227 1384 2231
rect 1530 2231 1536 2232
rect 1530 2230 1531 2231
rect 1517 2228 1531 2230
rect 1378 2226 1384 2227
rect 1530 2227 1531 2228
rect 1535 2227 1536 2231
rect 1682 2231 1688 2232
rect 1682 2230 1683 2231
rect 1669 2228 1683 2230
rect 1530 2226 1536 2227
rect 1682 2227 1683 2228
rect 1687 2227 1688 2231
rect 1682 2226 1688 2227
rect 1690 2231 1696 2232
rect 1894 2231 1900 2232
rect 2022 2236 2028 2237
rect 2022 2232 2023 2236
rect 2027 2232 2028 2236
rect 2022 2231 2028 2232
rect 2174 2236 2180 2237
rect 2174 2232 2175 2236
rect 2179 2232 2180 2236
rect 2174 2231 2180 2232
rect 2358 2236 2364 2237
rect 2358 2232 2359 2236
rect 2363 2232 2364 2236
rect 2358 2231 2364 2232
rect 2566 2236 2572 2237
rect 2566 2232 2567 2236
rect 2571 2232 2572 2236
rect 2566 2231 2572 2232
rect 2782 2236 2788 2237
rect 2782 2232 2783 2236
rect 2787 2232 2788 2236
rect 2782 2231 2788 2232
rect 3014 2236 3020 2237
rect 3014 2232 3015 2236
rect 3019 2232 3020 2236
rect 3014 2231 3020 2232
rect 3246 2236 3252 2237
rect 3246 2232 3247 2236
rect 3251 2232 3252 2236
rect 3246 2231 3252 2232
rect 3486 2236 3492 2237
rect 3486 2232 3487 2236
rect 3491 2232 3492 2236
rect 3590 2235 3591 2239
rect 3595 2235 3596 2239
rect 3590 2234 3596 2235
rect 3486 2231 3492 2232
rect 1690 2227 1691 2231
rect 1695 2230 1696 2231
rect 1695 2228 1761 2230
rect 1695 2227 1696 2228
rect 1690 2226 1696 2227
rect 998 2222 1004 2223
rect 110 2220 116 2221
rect 110 2216 111 2220
rect 115 2216 116 2220
rect 110 2215 116 2216
rect 1830 2220 1836 2221
rect 1830 2216 1831 2220
rect 1835 2216 1836 2220
rect 1830 2215 1836 2216
rect 2374 2219 2380 2220
rect 2374 2215 2375 2219
rect 2379 2218 2380 2219
rect 2799 2219 2805 2220
rect 2799 2218 2800 2219
rect 2379 2216 2800 2218
rect 2379 2215 2380 2216
rect 2374 2214 2380 2215
rect 2799 2215 2800 2216
rect 2804 2215 2805 2219
rect 2799 2214 2805 2215
rect 142 2202 148 2203
rect 142 2198 143 2202
rect 147 2198 148 2202
rect 142 2197 148 2198
rect 222 2202 228 2203
rect 222 2198 223 2202
rect 227 2198 228 2202
rect 222 2197 228 2198
rect 302 2202 308 2203
rect 302 2198 303 2202
rect 307 2198 308 2202
rect 302 2197 308 2198
rect 390 2202 396 2203
rect 390 2198 391 2202
rect 395 2198 396 2202
rect 390 2197 396 2198
rect 526 2202 532 2203
rect 526 2198 527 2202
rect 531 2198 532 2202
rect 526 2197 532 2198
rect 678 2202 684 2203
rect 678 2198 679 2202
rect 683 2198 684 2202
rect 678 2197 684 2198
rect 838 2202 844 2203
rect 838 2198 839 2202
rect 843 2198 844 2202
rect 838 2197 844 2198
rect 1006 2202 1012 2203
rect 1006 2198 1007 2202
rect 1011 2198 1012 2202
rect 1006 2197 1012 2198
rect 1166 2202 1172 2203
rect 1166 2198 1167 2202
rect 1171 2198 1172 2202
rect 1166 2197 1172 2198
rect 1318 2202 1324 2203
rect 1318 2198 1319 2202
rect 1323 2198 1324 2202
rect 1318 2197 1324 2198
rect 1462 2202 1468 2203
rect 1462 2198 1463 2202
rect 1467 2198 1468 2202
rect 1462 2197 1468 2198
rect 1614 2202 1620 2203
rect 1614 2198 1615 2202
rect 1619 2198 1620 2202
rect 1614 2197 1620 2198
rect 1750 2202 1756 2203
rect 1750 2198 1751 2202
rect 1755 2198 1756 2202
rect 1750 2197 1756 2198
rect 135 2191 141 2192
rect 135 2187 136 2191
rect 140 2190 141 2191
rect 143 2191 149 2192
rect 143 2190 144 2191
rect 140 2188 144 2190
rect 140 2187 141 2188
rect 135 2186 141 2187
rect 143 2187 144 2188
rect 148 2187 149 2191
rect 143 2186 149 2187
rect 202 2191 208 2192
rect 202 2187 203 2191
rect 207 2190 208 2191
rect 215 2191 221 2192
rect 215 2190 216 2191
rect 207 2188 216 2190
rect 207 2187 208 2188
rect 202 2186 208 2187
rect 215 2187 216 2188
rect 220 2187 221 2191
rect 215 2186 221 2187
rect 282 2191 288 2192
rect 282 2187 283 2191
rect 287 2190 288 2191
rect 295 2191 301 2192
rect 295 2190 296 2191
rect 287 2188 296 2190
rect 287 2187 288 2188
rect 282 2186 288 2187
rect 295 2187 296 2188
rect 300 2187 301 2191
rect 295 2186 301 2187
rect 362 2191 368 2192
rect 362 2187 363 2191
rect 367 2190 368 2191
rect 383 2191 389 2192
rect 383 2190 384 2191
rect 367 2188 384 2190
rect 367 2187 368 2188
rect 362 2186 368 2187
rect 383 2187 384 2188
rect 388 2187 389 2191
rect 383 2186 389 2187
rect 458 2191 464 2192
rect 458 2187 459 2191
rect 463 2190 464 2191
rect 519 2191 525 2192
rect 519 2190 520 2191
rect 463 2188 520 2190
rect 463 2187 464 2188
rect 458 2186 464 2187
rect 519 2187 520 2188
rect 524 2187 525 2191
rect 519 2186 525 2187
rect 586 2191 592 2192
rect 586 2187 587 2191
rect 591 2190 592 2191
rect 671 2191 677 2192
rect 671 2190 672 2191
rect 591 2188 672 2190
rect 591 2187 592 2188
rect 586 2186 592 2187
rect 671 2187 672 2188
rect 676 2187 677 2191
rect 671 2186 677 2187
rect 754 2191 760 2192
rect 754 2187 755 2191
rect 759 2190 760 2191
rect 831 2191 837 2192
rect 831 2190 832 2191
rect 759 2188 832 2190
rect 759 2187 760 2188
rect 754 2186 760 2187
rect 831 2187 832 2188
rect 836 2187 837 2191
rect 831 2186 837 2187
rect 922 2191 928 2192
rect 922 2187 923 2191
rect 927 2190 928 2191
rect 999 2191 1005 2192
rect 999 2190 1000 2191
rect 927 2188 1000 2190
rect 927 2187 928 2188
rect 922 2186 928 2187
rect 999 2187 1000 2188
rect 1004 2187 1005 2191
rect 999 2186 1005 2187
rect 1159 2191 1165 2192
rect 1159 2187 1160 2191
rect 1164 2190 1165 2191
rect 1174 2191 1180 2192
rect 1174 2190 1175 2191
rect 1164 2188 1175 2190
rect 1164 2187 1165 2188
rect 1159 2186 1165 2187
rect 1174 2187 1175 2188
rect 1179 2187 1180 2191
rect 1174 2186 1180 2187
rect 1234 2191 1240 2192
rect 1234 2187 1235 2191
rect 1239 2190 1240 2191
rect 1311 2191 1317 2192
rect 1311 2190 1312 2191
rect 1239 2188 1312 2190
rect 1239 2187 1240 2188
rect 1234 2186 1240 2187
rect 1311 2187 1312 2188
rect 1316 2187 1317 2191
rect 1311 2186 1317 2187
rect 1378 2191 1384 2192
rect 1378 2187 1379 2191
rect 1383 2190 1384 2191
rect 1455 2191 1461 2192
rect 1455 2190 1456 2191
rect 1383 2188 1456 2190
rect 1383 2187 1384 2188
rect 1378 2186 1384 2187
rect 1455 2187 1456 2188
rect 1460 2187 1461 2191
rect 1455 2186 1461 2187
rect 1530 2191 1536 2192
rect 1530 2187 1531 2191
rect 1535 2190 1536 2191
rect 1607 2191 1613 2192
rect 1607 2190 1608 2191
rect 1535 2188 1608 2190
rect 1535 2187 1536 2188
rect 1530 2186 1536 2187
rect 1607 2187 1608 2188
rect 1612 2187 1613 2191
rect 1607 2186 1613 2187
rect 1682 2191 1688 2192
rect 1682 2187 1683 2191
rect 1687 2190 1688 2191
rect 1743 2191 1749 2192
rect 1743 2190 1744 2191
rect 1687 2188 1744 2190
rect 1687 2187 1688 2188
rect 1682 2186 1688 2187
rect 1743 2187 1744 2188
rect 1748 2187 1749 2191
rect 1743 2186 1749 2187
rect 183 2175 189 2176
rect 183 2171 184 2175
rect 188 2174 189 2175
rect 198 2175 204 2176
rect 198 2174 199 2175
rect 188 2172 199 2174
rect 188 2171 189 2172
rect 183 2170 189 2171
rect 198 2171 199 2172
rect 203 2171 204 2175
rect 198 2170 204 2171
rect 282 2175 288 2176
rect 282 2171 283 2175
rect 287 2174 288 2175
rect 303 2175 309 2176
rect 303 2174 304 2175
rect 287 2172 304 2174
rect 287 2171 288 2172
rect 282 2170 288 2171
rect 303 2171 304 2172
rect 308 2171 309 2175
rect 303 2170 309 2171
rect 362 2175 368 2176
rect 362 2171 363 2175
rect 367 2174 368 2175
rect 455 2175 461 2176
rect 455 2174 456 2175
rect 367 2172 456 2174
rect 367 2171 368 2172
rect 362 2170 368 2171
rect 455 2171 456 2172
rect 460 2171 461 2175
rect 455 2170 461 2171
rect 631 2175 637 2176
rect 631 2171 632 2175
rect 636 2174 637 2175
rect 646 2175 652 2176
rect 646 2174 647 2175
rect 636 2172 647 2174
rect 636 2171 637 2172
rect 631 2170 637 2171
rect 646 2171 647 2172
rect 651 2171 652 2175
rect 646 2170 652 2171
rect 690 2175 696 2176
rect 690 2171 691 2175
rect 695 2174 696 2175
rect 815 2175 821 2176
rect 815 2174 816 2175
rect 695 2172 816 2174
rect 695 2171 696 2172
rect 690 2170 696 2171
rect 815 2171 816 2172
rect 820 2171 821 2175
rect 815 2170 821 2171
rect 998 2175 1004 2176
rect 998 2171 999 2175
rect 1003 2174 1004 2175
rect 1007 2175 1013 2176
rect 1007 2174 1008 2175
rect 1003 2172 1008 2174
rect 1003 2171 1004 2172
rect 998 2170 1004 2171
rect 1007 2171 1008 2172
rect 1012 2171 1013 2175
rect 1007 2170 1013 2171
rect 1191 2175 1197 2176
rect 1191 2171 1192 2175
rect 1196 2174 1197 2175
rect 1206 2175 1212 2176
rect 1206 2174 1207 2175
rect 1196 2172 1207 2174
rect 1196 2171 1197 2172
rect 1191 2170 1197 2171
rect 1206 2171 1207 2172
rect 1211 2171 1212 2175
rect 1206 2170 1212 2171
rect 1250 2175 1256 2176
rect 1250 2171 1251 2175
rect 1255 2174 1256 2175
rect 1383 2175 1389 2176
rect 1383 2174 1384 2175
rect 1255 2172 1384 2174
rect 1255 2171 1256 2172
rect 1250 2170 1256 2171
rect 1383 2171 1384 2172
rect 1388 2171 1389 2175
rect 1383 2170 1389 2171
rect 1442 2175 1448 2176
rect 1442 2171 1443 2175
rect 1447 2174 1448 2175
rect 1575 2175 1581 2176
rect 1575 2174 1576 2175
rect 1447 2172 1576 2174
rect 1447 2171 1448 2172
rect 1442 2170 1448 2171
rect 1575 2171 1576 2172
rect 1580 2171 1581 2175
rect 1575 2170 1581 2171
rect 1634 2175 1640 2176
rect 1634 2171 1635 2175
rect 1639 2174 1640 2175
rect 1743 2175 1749 2176
rect 1743 2174 1744 2175
rect 1639 2172 1744 2174
rect 1639 2171 1640 2172
rect 1634 2170 1640 2171
rect 1743 2171 1744 2172
rect 1748 2171 1749 2175
rect 1743 2170 1749 2171
rect 2198 2172 2204 2173
rect 1870 2169 1876 2170
rect 190 2166 196 2167
rect 190 2162 191 2166
rect 195 2162 196 2166
rect 190 2161 196 2162
rect 310 2166 316 2167
rect 310 2162 311 2166
rect 315 2162 316 2166
rect 310 2161 316 2162
rect 462 2166 468 2167
rect 462 2162 463 2166
rect 467 2162 468 2166
rect 462 2161 468 2162
rect 638 2166 644 2167
rect 638 2162 639 2166
rect 643 2162 644 2166
rect 638 2161 644 2162
rect 822 2166 828 2167
rect 822 2162 823 2166
rect 827 2162 828 2166
rect 822 2161 828 2162
rect 1014 2166 1020 2167
rect 1014 2162 1015 2166
rect 1019 2162 1020 2166
rect 1014 2161 1020 2162
rect 1198 2166 1204 2167
rect 1198 2162 1199 2166
rect 1203 2162 1204 2166
rect 1198 2161 1204 2162
rect 1390 2166 1396 2167
rect 1390 2162 1391 2166
rect 1395 2162 1396 2166
rect 1390 2161 1396 2162
rect 1582 2166 1588 2167
rect 1582 2162 1583 2166
rect 1587 2162 1588 2166
rect 1582 2161 1588 2162
rect 1750 2166 1756 2167
rect 1750 2162 1751 2166
rect 1755 2162 1756 2166
rect 1870 2165 1871 2169
rect 1875 2165 1876 2169
rect 2198 2168 2199 2172
rect 2203 2168 2204 2172
rect 2198 2167 2204 2168
rect 2294 2172 2300 2173
rect 2294 2168 2295 2172
rect 2299 2168 2300 2172
rect 2294 2167 2300 2168
rect 2398 2172 2404 2173
rect 2398 2168 2399 2172
rect 2403 2168 2404 2172
rect 2398 2167 2404 2168
rect 2518 2172 2524 2173
rect 2518 2168 2519 2172
rect 2523 2168 2524 2172
rect 2518 2167 2524 2168
rect 2638 2172 2644 2173
rect 2638 2168 2639 2172
rect 2643 2168 2644 2172
rect 2638 2167 2644 2168
rect 2758 2172 2764 2173
rect 2758 2168 2759 2172
rect 2763 2168 2764 2172
rect 2758 2167 2764 2168
rect 2878 2172 2884 2173
rect 2878 2168 2879 2172
rect 2883 2168 2884 2172
rect 2878 2167 2884 2168
rect 2990 2172 2996 2173
rect 2990 2168 2991 2172
rect 2995 2168 2996 2172
rect 2990 2167 2996 2168
rect 3094 2172 3100 2173
rect 3094 2168 3095 2172
rect 3099 2168 3100 2172
rect 3094 2167 3100 2168
rect 3198 2172 3204 2173
rect 3198 2168 3199 2172
rect 3203 2168 3204 2172
rect 3198 2167 3204 2168
rect 3302 2172 3308 2173
rect 3302 2168 3303 2172
rect 3307 2168 3308 2172
rect 3302 2167 3308 2168
rect 3406 2172 3412 2173
rect 3406 2168 3407 2172
rect 3411 2168 3412 2172
rect 3406 2167 3412 2168
rect 3502 2172 3508 2173
rect 3502 2168 3503 2172
rect 3507 2168 3508 2172
rect 3502 2167 3508 2168
rect 3590 2169 3596 2170
rect 1870 2164 1876 2165
rect 3590 2165 3591 2169
rect 3595 2165 3596 2169
rect 3590 2164 3596 2165
rect 2266 2163 2272 2164
rect 2266 2162 2267 2163
rect 1750 2161 1756 2162
rect 2261 2160 2267 2162
rect 2266 2159 2267 2160
rect 2271 2159 2272 2163
rect 2362 2163 2368 2164
rect 2362 2162 2363 2163
rect 2357 2160 2363 2162
rect 2266 2158 2272 2159
rect 2362 2159 2363 2160
rect 2367 2159 2368 2163
rect 2478 2163 2484 2164
rect 2478 2162 2479 2163
rect 2461 2160 2479 2162
rect 2362 2158 2368 2159
rect 2478 2159 2479 2160
rect 2483 2159 2484 2163
rect 2478 2158 2484 2159
rect 2486 2163 2492 2164
rect 2486 2159 2487 2163
rect 2491 2162 2492 2163
rect 2586 2163 2592 2164
rect 2491 2160 2537 2162
rect 2491 2159 2492 2160
rect 2486 2158 2492 2159
rect 2586 2159 2587 2163
rect 2591 2162 2592 2163
rect 2706 2163 2712 2164
rect 2591 2160 2657 2162
rect 2591 2159 2592 2160
rect 2586 2158 2592 2159
rect 2706 2159 2707 2163
rect 2711 2162 2712 2163
rect 2847 2163 2853 2164
rect 2711 2160 2777 2162
rect 2711 2159 2712 2160
rect 2706 2158 2712 2159
rect 2847 2159 2848 2163
rect 2852 2162 2853 2163
rect 2946 2163 2952 2164
rect 2852 2160 2897 2162
rect 2852 2159 2853 2160
rect 2847 2158 2853 2159
rect 2946 2159 2947 2163
rect 2951 2162 2952 2163
rect 3058 2163 3064 2164
rect 2951 2160 3009 2162
rect 2951 2159 2952 2160
rect 2946 2158 2952 2159
rect 3058 2159 3059 2163
rect 3063 2162 3064 2163
rect 3174 2163 3180 2164
rect 3063 2160 3113 2162
rect 3063 2159 3064 2160
rect 3058 2158 3064 2159
rect 3174 2159 3175 2163
rect 3179 2162 3180 2163
rect 3266 2163 3272 2164
rect 3179 2160 3217 2162
rect 3179 2159 3180 2160
rect 3174 2158 3180 2159
rect 3266 2159 3267 2163
rect 3271 2162 3272 2163
rect 3474 2163 3480 2164
rect 3474 2162 3475 2163
rect 3271 2160 3321 2162
rect 3469 2160 3475 2162
rect 3271 2159 3272 2160
rect 3266 2158 3272 2159
rect 3474 2159 3475 2160
rect 3479 2159 3480 2163
rect 3504 2160 3521 2162
rect 3474 2158 3480 2159
rect 3502 2159 3508 2160
rect 3502 2155 3503 2159
rect 3507 2155 3508 2159
rect 3502 2154 3508 2155
rect 1870 2152 1876 2153
rect 110 2148 116 2149
rect 110 2144 111 2148
rect 115 2144 116 2148
rect 110 2143 116 2144
rect 1830 2148 1836 2149
rect 1830 2144 1831 2148
rect 1835 2144 1836 2148
rect 1870 2148 1871 2152
rect 1875 2148 1876 2152
rect 1870 2147 1876 2148
rect 3590 2152 3596 2153
rect 3590 2148 3591 2152
rect 3595 2148 3596 2152
rect 3590 2147 3596 2148
rect 1830 2143 1836 2144
rect 143 2139 149 2140
rect 143 2135 144 2139
rect 148 2138 149 2139
rect 362 2139 368 2140
rect 148 2136 201 2138
rect 148 2135 149 2136
rect 143 2134 149 2135
rect 362 2135 363 2139
rect 367 2135 368 2139
rect 362 2134 368 2135
rect 470 2139 476 2140
rect 470 2135 471 2139
rect 475 2135 476 2139
rect 470 2134 476 2135
rect 690 2139 696 2140
rect 690 2135 691 2139
rect 695 2135 696 2139
rect 690 2134 696 2135
rect 874 2139 880 2140
rect 874 2135 875 2139
rect 879 2135 880 2139
rect 874 2134 880 2135
rect 1022 2139 1028 2140
rect 1022 2135 1023 2139
rect 1027 2135 1028 2139
rect 1022 2134 1028 2135
rect 1250 2139 1256 2140
rect 1250 2135 1251 2139
rect 1255 2135 1256 2139
rect 1250 2134 1256 2135
rect 1442 2139 1448 2140
rect 1442 2135 1443 2139
rect 1447 2135 1448 2139
rect 1442 2134 1448 2135
rect 1634 2139 1640 2140
rect 1634 2135 1635 2139
rect 1639 2135 1640 2139
rect 1634 2134 1640 2135
rect 2206 2134 2212 2135
rect 110 2131 116 2132
rect 110 2127 111 2131
rect 115 2127 116 2131
rect 1830 2131 1836 2132
rect 110 2126 116 2127
rect 182 2128 188 2129
rect 182 2124 183 2128
rect 187 2124 188 2128
rect 182 2123 188 2124
rect 302 2128 308 2129
rect 302 2124 303 2128
rect 307 2124 308 2128
rect 302 2123 308 2124
rect 454 2128 460 2129
rect 454 2124 455 2128
rect 459 2124 460 2128
rect 454 2123 460 2124
rect 630 2128 636 2129
rect 630 2124 631 2128
rect 635 2124 636 2128
rect 630 2123 636 2124
rect 814 2128 820 2129
rect 814 2124 815 2128
rect 819 2124 820 2128
rect 814 2123 820 2124
rect 1006 2128 1012 2129
rect 1006 2124 1007 2128
rect 1011 2124 1012 2128
rect 1006 2123 1012 2124
rect 1190 2128 1196 2129
rect 1190 2124 1191 2128
rect 1195 2124 1196 2128
rect 1190 2123 1196 2124
rect 1382 2128 1388 2129
rect 1382 2124 1383 2128
rect 1387 2124 1388 2128
rect 1382 2123 1388 2124
rect 1574 2128 1580 2129
rect 1574 2124 1575 2128
rect 1579 2124 1580 2128
rect 1574 2123 1580 2124
rect 1742 2128 1748 2129
rect 1742 2124 1743 2128
rect 1747 2124 1748 2128
rect 1830 2127 1831 2131
rect 1835 2127 1836 2131
rect 2206 2130 2207 2134
rect 2211 2130 2212 2134
rect 2206 2129 2212 2130
rect 2302 2134 2308 2135
rect 2302 2130 2303 2134
rect 2307 2130 2308 2134
rect 2302 2129 2308 2130
rect 2406 2134 2412 2135
rect 2406 2130 2407 2134
rect 2411 2130 2412 2134
rect 2406 2129 2412 2130
rect 2526 2134 2532 2135
rect 2526 2130 2527 2134
rect 2531 2130 2532 2134
rect 2526 2129 2532 2130
rect 2646 2134 2652 2135
rect 2646 2130 2647 2134
rect 2651 2130 2652 2134
rect 2646 2129 2652 2130
rect 2766 2134 2772 2135
rect 2766 2130 2767 2134
rect 2771 2130 2772 2134
rect 2766 2129 2772 2130
rect 2886 2134 2892 2135
rect 2886 2130 2887 2134
rect 2891 2130 2892 2134
rect 2886 2129 2892 2130
rect 2998 2134 3004 2135
rect 2998 2130 2999 2134
rect 3003 2130 3004 2134
rect 2998 2129 3004 2130
rect 3102 2134 3108 2135
rect 3102 2130 3103 2134
rect 3107 2130 3108 2134
rect 3102 2129 3108 2130
rect 3206 2134 3212 2135
rect 3206 2130 3207 2134
rect 3211 2130 3212 2134
rect 3206 2129 3212 2130
rect 3310 2134 3316 2135
rect 3310 2130 3311 2134
rect 3315 2130 3316 2134
rect 3310 2129 3316 2130
rect 3414 2134 3420 2135
rect 3414 2130 3415 2134
rect 3419 2130 3420 2134
rect 3414 2129 3420 2130
rect 3510 2134 3516 2135
rect 3510 2130 3511 2134
rect 3515 2130 3516 2134
rect 3510 2129 3516 2130
rect 1830 2126 1836 2127
rect 1742 2123 1748 2124
rect 2199 2123 2205 2124
rect 2199 2119 2200 2123
rect 2204 2122 2205 2123
rect 2214 2123 2220 2124
rect 2214 2122 2215 2123
rect 2204 2120 2215 2122
rect 2204 2119 2205 2120
rect 2199 2118 2205 2119
rect 2214 2119 2215 2120
rect 2219 2119 2220 2123
rect 2214 2118 2220 2119
rect 2266 2123 2272 2124
rect 2266 2119 2267 2123
rect 2271 2122 2272 2123
rect 2295 2123 2301 2124
rect 2295 2122 2296 2123
rect 2271 2120 2296 2122
rect 2271 2119 2272 2120
rect 2266 2118 2272 2119
rect 2295 2119 2296 2120
rect 2300 2119 2301 2123
rect 2295 2118 2301 2119
rect 2362 2123 2368 2124
rect 2362 2119 2363 2123
rect 2367 2122 2368 2123
rect 2399 2123 2405 2124
rect 2399 2122 2400 2123
rect 2367 2120 2400 2122
rect 2367 2119 2368 2120
rect 2362 2118 2368 2119
rect 2399 2119 2400 2120
rect 2404 2119 2405 2123
rect 2399 2118 2405 2119
rect 2519 2123 2525 2124
rect 2519 2119 2520 2123
rect 2524 2122 2525 2123
rect 2586 2123 2592 2124
rect 2586 2122 2587 2123
rect 2524 2120 2587 2122
rect 2524 2119 2525 2120
rect 2519 2118 2525 2119
rect 2586 2119 2587 2120
rect 2591 2119 2592 2123
rect 2586 2118 2592 2119
rect 2639 2123 2645 2124
rect 2639 2119 2640 2123
rect 2644 2122 2645 2123
rect 2706 2123 2712 2124
rect 2706 2122 2707 2123
rect 2644 2120 2707 2122
rect 2644 2119 2645 2120
rect 2639 2118 2645 2119
rect 2706 2119 2707 2120
rect 2711 2119 2712 2123
rect 2706 2118 2712 2119
rect 2758 2123 2765 2124
rect 2758 2119 2759 2123
rect 2764 2119 2765 2123
rect 2758 2118 2765 2119
rect 2879 2123 2885 2124
rect 2879 2119 2880 2123
rect 2884 2122 2885 2123
rect 2946 2123 2952 2124
rect 2946 2122 2947 2123
rect 2884 2120 2947 2122
rect 2884 2119 2885 2120
rect 2879 2118 2885 2119
rect 2946 2119 2947 2120
rect 2951 2119 2952 2123
rect 2946 2118 2952 2119
rect 2991 2123 2997 2124
rect 2991 2119 2992 2123
rect 2996 2122 2997 2123
rect 3058 2123 3064 2124
rect 3058 2122 3059 2123
rect 2996 2120 3059 2122
rect 2996 2119 2997 2120
rect 2991 2118 2997 2119
rect 3058 2119 3059 2120
rect 3063 2119 3064 2123
rect 3058 2118 3064 2119
rect 3095 2123 3101 2124
rect 3095 2119 3096 2123
rect 3100 2122 3101 2123
rect 3174 2123 3180 2124
rect 3174 2122 3175 2123
rect 3100 2120 3175 2122
rect 3100 2119 3101 2120
rect 3095 2118 3101 2119
rect 3174 2119 3175 2120
rect 3179 2119 3180 2123
rect 3174 2118 3180 2119
rect 3199 2123 3205 2124
rect 3199 2119 3200 2123
rect 3204 2122 3205 2123
rect 3266 2123 3272 2124
rect 3266 2122 3267 2123
rect 3204 2120 3267 2122
rect 3204 2119 3205 2120
rect 3199 2118 3205 2119
rect 3266 2119 3267 2120
rect 3271 2119 3272 2123
rect 3266 2118 3272 2119
rect 3303 2123 3309 2124
rect 3303 2119 3304 2123
rect 3308 2122 3309 2123
rect 3318 2123 3324 2124
rect 3318 2122 3319 2123
rect 3308 2120 3319 2122
rect 3308 2119 3309 2120
rect 3303 2118 3309 2119
rect 3318 2119 3319 2120
rect 3323 2119 3324 2123
rect 3318 2118 3324 2119
rect 3334 2123 3340 2124
rect 3334 2119 3335 2123
rect 3339 2122 3340 2123
rect 3407 2123 3413 2124
rect 3407 2122 3408 2123
rect 3339 2120 3408 2122
rect 3339 2119 3340 2120
rect 3334 2118 3340 2119
rect 3407 2119 3408 2120
rect 3412 2119 3413 2123
rect 3407 2118 3413 2119
rect 3474 2123 3480 2124
rect 3474 2119 3475 2123
rect 3479 2122 3480 2123
rect 3503 2123 3509 2124
rect 3503 2122 3504 2123
rect 3479 2120 3504 2122
rect 3479 2119 3480 2120
rect 3474 2118 3480 2119
rect 3503 2119 3504 2120
rect 3508 2119 3509 2123
rect 3503 2118 3509 2119
rect 1758 2111 1765 2112
rect 1758 2107 1759 2111
rect 1764 2107 1765 2111
rect 1758 2106 1765 2107
rect 2454 2107 2460 2108
rect 2454 2106 2455 2107
rect 2220 2104 2455 2106
rect 2167 2099 2173 2100
rect 2167 2095 2168 2099
rect 2172 2098 2173 2099
rect 2220 2098 2222 2104
rect 2454 2103 2455 2104
rect 2459 2103 2460 2107
rect 3422 2107 3428 2108
rect 3422 2106 3423 2107
rect 2454 2102 2460 2103
rect 3236 2104 3423 2106
rect 2172 2096 2222 2098
rect 2226 2099 2232 2100
rect 2172 2095 2173 2096
rect 2167 2094 2173 2095
rect 2226 2095 2227 2099
rect 2231 2098 2232 2099
rect 2263 2099 2269 2100
rect 2263 2098 2264 2099
rect 2231 2096 2264 2098
rect 2231 2095 2232 2096
rect 2226 2094 2232 2095
rect 2263 2095 2264 2096
rect 2268 2095 2269 2099
rect 2263 2094 2269 2095
rect 2322 2099 2328 2100
rect 2322 2095 2323 2099
rect 2327 2098 2328 2099
rect 2367 2099 2373 2100
rect 2367 2098 2368 2099
rect 2327 2096 2368 2098
rect 2327 2095 2328 2096
rect 2322 2094 2328 2095
rect 2367 2095 2368 2096
rect 2372 2095 2373 2099
rect 2367 2094 2373 2095
rect 2426 2099 2432 2100
rect 2426 2095 2427 2099
rect 2431 2098 2432 2099
rect 2479 2099 2485 2100
rect 2479 2098 2480 2099
rect 2431 2096 2480 2098
rect 2431 2095 2432 2096
rect 2426 2094 2432 2095
rect 2479 2095 2480 2096
rect 2484 2095 2485 2099
rect 2479 2094 2485 2095
rect 2538 2099 2544 2100
rect 2538 2095 2539 2099
rect 2543 2098 2544 2099
rect 2599 2099 2605 2100
rect 2599 2098 2600 2099
rect 2543 2096 2600 2098
rect 2543 2095 2544 2096
rect 2538 2094 2544 2095
rect 2599 2095 2600 2096
rect 2604 2095 2605 2099
rect 2599 2094 2605 2095
rect 2658 2099 2664 2100
rect 2658 2095 2659 2099
rect 2663 2098 2664 2099
rect 2719 2099 2725 2100
rect 2719 2098 2720 2099
rect 2663 2096 2720 2098
rect 2663 2095 2664 2096
rect 2658 2094 2664 2095
rect 2719 2095 2720 2096
rect 2724 2095 2725 2099
rect 2719 2094 2725 2095
rect 2839 2099 2845 2100
rect 2839 2095 2840 2099
rect 2844 2098 2845 2099
rect 2847 2099 2853 2100
rect 2847 2098 2848 2099
rect 2844 2096 2848 2098
rect 2844 2095 2845 2096
rect 2839 2094 2845 2095
rect 2847 2095 2848 2096
rect 2852 2095 2853 2099
rect 2847 2094 2853 2095
rect 2898 2099 2904 2100
rect 2898 2095 2899 2099
rect 2903 2098 2904 2099
rect 2959 2099 2965 2100
rect 2959 2098 2960 2099
rect 2903 2096 2960 2098
rect 2903 2095 2904 2096
rect 2898 2094 2904 2095
rect 2959 2095 2960 2096
rect 2964 2095 2965 2099
rect 2959 2094 2965 2095
rect 3018 2099 3024 2100
rect 3018 2095 3019 2099
rect 3023 2098 3024 2099
rect 3071 2099 3077 2100
rect 3071 2098 3072 2099
rect 3023 2096 3072 2098
rect 3023 2095 3024 2096
rect 3018 2094 3024 2095
rect 3071 2095 3072 2096
rect 3076 2095 3077 2099
rect 3071 2094 3077 2095
rect 3183 2099 3189 2100
rect 3183 2095 3184 2099
rect 3188 2098 3189 2099
rect 3236 2098 3238 2104
rect 3422 2103 3423 2104
rect 3427 2103 3428 2107
rect 3422 2102 3428 2103
rect 3188 2096 3238 2098
rect 3242 2099 3248 2100
rect 3188 2095 3189 2096
rect 3183 2094 3189 2095
rect 3242 2095 3243 2099
rect 3247 2098 3248 2099
rect 3295 2099 3301 2100
rect 3295 2098 3296 2099
rect 3247 2096 3296 2098
rect 3247 2095 3248 2096
rect 3242 2094 3248 2095
rect 3295 2095 3296 2096
rect 3300 2095 3301 2099
rect 3295 2094 3301 2095
rect 3407 2099 3413 2100
rect 3407 2095 3408 2099
rect 3412 2098 3413 2099
rect 3430 2099 3436 2100
rect 3430 2098 3431 2099
rect 3412 2096 3431 2098
rect 3412 2095 3413 2096
rect 3407 2094 3413 2095
rect 3430 2095 3431 2096
rect 3435 2095 3436 2099
rect 3430 2094 3436 2095
rect 3502 2099 3509 2100
rect 3502 2095 3503 2099
rect 3508 2095 3509 2099
rect 3502 2094 3509 2095
rect 2174 2090 2180 2091
rect 2174 2086 2175 2090
rect 2179 2086 2180 2090
rect 2174 2085 2180 2086
rect 2270 2090 2276 2091
rect 2270 2086 2271 2090
rect 2275 2086 2276 2090
rect 2270 2085 2276 2086
rect 2374 2090 2380 2091
rect 2374 2086 2375 2090
rect 2379 2086 2380 2090
rect 2374 2085 2380 2086
rect 2486 2090 2492 2091
rect 2486 2086 2487 2090
rect 2491 2086 2492 2090
rect 2486 2085 2492 2086
rect 2606 2090 2612 2091
rect 2606 2086 2607 2090
rect 2611 2086 2612 2090
rect 2606 2085 2612 2086
rect 2726 2090 2732 2091
rect 2726 2086 2727 2090
rect 2731 2086 2732 2090
rect 2726 2085 2732 2086
rect 2846 2090 2852 2091
rect 2846 2086 2847 2090
rect 2851 2086 2852 2090
rect 2846 2085 2852 2086
rect 2966 2090 2972 2091
rect 2966 2086 2967 2090
rect 2971 2086 2972 2090
rect 2966 2085 2972 2086
rect 3078 2090 3084 2091
rect 3078 2086 3079 2090
rect 3083 2086 3084 2090
rect 3078 2085 3084 2086
rect 3190 2090 3196 2091
rect 3190 2086 3191 2090
rect 3195 2086 3196 2090
rect 3190 2085 3196 2086
rect 3302 2090 3308 2091
rect 3302 2086 3303 2090
rect 3307 2086 3308 2090
rect 3302 2085 3308 2086
rect 3414 2090 3420 2091
rect 3414 2086 3415 2090
rect 3419 2086 3420 2090
rect 3414 2085 3420 2086
rect 3510 2090 3516 2091
rect 3510 2086 3511 2090
rect 3515 2086 3516 2090
rect 3510 2085 3516 2086
rect 214 2080 220 2081
rect 110 2077 116 2078
rect 110 2073 111 2077
rect 115 2073 116 2077
rect 214 2076 215 2080
rect 219 2076 220 2080
rect 214 2075 220 2076
rect 358 2080 364 2081
rect 358 2076 359 2080
rect 363 2076 364 2080
rect 358 2075 364 2076
rect 518 2080 524 2081
rect 518 2076 519 2080
rect 523 2076 524 2080
rect 518 2075 524 2076
rect 702 2080 708 2081
rect 702 2076 703 2080
rect 707 2076 708 2080
rect 702 2075 708 2076
rect 894 2080 900 2081
rect 894 2076 895 2080
rect 899 2076 900 2080
rect 894 2075 900 2076
rect 1102 2080 1108 2081
rect 1102 2076 1103 2080
rect 1107 2076 1108 2080
rect 1102 2075 1108 2076
rect 1310 2080 1316 2081
rect 1310 2076 1311 2080
rect 1315 2076 1316 2080
rect 1310 2075 1316 2076
rect 1526 2080 1532 2081
rect 1526 2076 1527 2080
rect 1531 2076 1532 2080
rect 1526 2075 1532 2076
rect 1742 2080 1748 2081
rect 1742 2076 1743 2080
rect 1747 2076 1748 2080
rect 1742 2075 1748 2076
rect 1830 2077 1836 2078
rect 110 2072 116 2073
rect 1830 2073 1831 2077
rect 1835 2073 1836 2077
rect 1830 2072 1836 2073
rect 1870 2072 1876 2073
rect 282 2071 288 2072
rect 282 2070 283 2071
rect 277 2068 283 2070
rect 282 2067 283 2068
rect 287 2067 288 2071
rect 282 2066 288 2067
rect 290 2071 296 2072
rect 290 2067 291 2071
rect 295 2070 296 2071
rect 495 2071 501 2072
rect 295 2068 377 2070
rect 295 2067 296 2068
rect 290 2066 296 2067
rect 495 2067 496 2071
rect 500 2070 501 2071
rect 586 2071 592 2072
rect 500 2068 537 2070
rect 500 2067 501 2068
rect 495 2066 501 2067
rect 586 2067 587 2071
rect 591 2070 592 2071
rect 770 2071 776 2072
rect 591 2068 721 2070
rect 591 2067 592 2068
rect 586 2066 592 2067
rect 770 2067 771 2071
rect 775 2070 776 2071
rect 1214 2071 1220 2072
rect 1214 2070 1215 2071
rect 775 2068 913 2070
rect 1165 2068 1215 2070
rect 775 2067 776 2068
rect 770 2066 776 2067
rect 1214 2067 1215 2068
rect 1219 2067 1220 2071
rect 1594 2071 1600 2072
rect 1594 2070 1595 2071
rect 1214 2066 1220 2067
rect 1095 2063 1101 2064
rect 110 2060 116 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 1095 2059 1096 2063
rect 1100 2062 1101 2063
rect 1328 2062 1330 2069
rect 1589 2068 1595 2070
rect 1594 2067 1595 2068
rect 1599 2067 1600 2071
rect 1594 2066 1600 2067
rect 1602 2071 1608 2072
rect 1602 2067 1603 2071
rect 1607 2070 1608 2071
rect 1607 2068 1761 2070
rect 1870 2068 1871 2072
rect 1875 2068 1876 2072
rect 1607 2067 1608 2068
rect 1870 2067 1876 2068
rect 3590 2072 3596 2073
rect 3590 2068 3591 2072
rect 3595 2068 3596 2072
rect 3590 2067 3596 2068
rect 1602 2066 1608 2067
rect 1100 2060 1330 2062
rect 2226 2063 2232 2064
rect 1830 2060 1836 2061
rect 1100 2059 1101 2060
rect 1095 2058 1101 2059
rect 110 2055 116 2056
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 2226 2059 2227 2063
rect 2231 2059 2232 2063
rect 2226 2058 2232 2059
rect 2322 2063 2328 2064
rect 2322 2059 2323 2063
rect 2327 2059 2328 2063
rect 2322 2058 2328 2059
rect 2426 2063 2432 2064
rect 2426 2059 2427 2063
rect 2431 2059 2432 2063
rect 2426 2058 2432 2059
rect 2538 2063 2544 2064
rect 2538 2059 2539 2063
rect 2543 2059 2544 2063
rect 2538 2058 2544 2059
rect 2658 2063 2664 2064
rect 2658 2059 2659 2063
rect 2663 2059 2664 2063
rect 2658 2058 2664 2059
rect 2758 2063 2764 2064
rect 2758 2059 2759 2063
rect 2763 2059 2764 2063
rect 2758 2058 2764 2059
rect 2898 2063 2904 2064
rect 2898 2059 2899 2063
rect 2903 2059 2904 2063
rect 2898 2058 2904 2059
rect 3018 2063 3024 2064
rect 3018 2059 3019 2063
rect 3023 2059 3024 2063
rect 3018 2058 3024 2059
rect 3242 2063 3248 2064
rect 3242 2059 3243 2063
rect 3247 2059 3248 2063
rect 3242 2058 3248 2059
rect 3318 2063 3324 2064
rect 3318 2059 3319 2063
rect 3323 2059 3324 2063
rect 3318 2058 3324 2059
rect 3422 2063 3428 2064
rect 3422 2059 3423 2063
rect 3427 2059 3428 2063
rect 3422 2058 3428 2059
rect 1830 2055 1836 2056
rect 1870 2055 1876 2056
rect 1870 2051 1871 2055
rect 1875 2051 1876 2055
rect 3590 2055 3596 2056
rect 1870 2050 1876 2051
rect 2166 2052 2172 2053
rect 2166 2048 2167 2052
rect 2171 2048 2172 2052
rect 2166 2047 2172 2048
rect 2262 2052 2268 2053
rect 2262 2048 2263 2052
rect 2267 2048 2268 2052
rect 2262 2047 2268 2048
rect 2366 2052 2372 2053
rect 2366 2048 2367 2052
rect 2371 2048 2372 2052
rect 2366 2047 2372 2048
rect 2478 2052 2484 2053
rect 2478 2048 2479 2052
rect 2483 2048 2484 2052
rect 2478 2047 2484 2048
rect 2598 2052 2604 2053
rect 2598 2048 2599 2052
rect 2603 2048 2604 2052
rect 2598 2047 2604 2048
rect 2718 2052 2724 2053
rect 2718 2048 2719 2052
rect 2723 2048 2724 2052
rect 2718 2047 2724 2048
rect 2838 2052 2844 2053
rect 2838 2048 2839 2052
rect 2843 2048 2844 2052
rect 2838 2047 2844 2048
rect 2958 2052 2964 2053
rect 2958 2048 2959 2052
rect 2963 2048 2964 2052
rect 2958 2047 2964 2048
rect 3070 2052 3076 2053
rect 3070 2048 3071 2052
rect 3075 2048 3076 2052
rect 3070 2047 3076 2048
rect 3182 2052 3188 2053
rect 3182 2048 3183 2052
rect 3187 2048 3188 2052
rect 3182 2047 3188 2048
rect 3294 2052 3300 2053
rect 3294 2048 3295 2052
rect 3299 2048 3300 2052
rect 3294 2047 3300 2048
rect 3406 2052 3412 2053
rect 3406 2048 3407 2052
rect 3411 2048 3412 2052
rect 3406 2047 3412 2048
rect 3502 2052 3508 2053
rect 3502 2048 3503 2052
rect 3507 2048 3508 2052
rect 3590 2051 3591 2055
rect 3595 2051 3596 2055
rect 3590 2050 3596 2051
rect 3502 2047 3508 2048
rect 222 2042 228 2043
rect 222 2038 223 2042
rect 227 2038 228 2042
rect 222 2037 228 2038
rect 366 2042 372 2043
rect 366 2038 367 2042
rect 371 2038 372 2042
rect 366 2037 372 2038
rect 526 2042 532 2043
rect 526 2038 527 2042
rect 531 2038 532 2042
rect 526 2037 532 2038
rect 710 2042 716 2043
rect 710 2038 711 2042
rect 715 2038 716 2042
rect 710 2037 716 2038
rect 902 2042 908 2043
rect 902 2038 903 2042
rect 907 2038 908 2042
rect 902 2037 908 2038
rect 1110 2042 1116 2043
rect 1110 2038 1111 2042
rect 1115 2038 1116 2042
rect 1110 2037 1116 2038
rect 1318 2042 1324 2043
rect 1318 2038 1319 2042
rect 1323 2038 1324 2042
rect 1318 2037 1324 2038
rect 1534 2042 1540 2043
rect 1534 2038 1535 2042
rect 1539 2038 1540 2042
rect 1534 2037 1540 2038
rect 1750 2042 1756 2043
rect 1750 2038 1751 2042
rect 1755 2038 1756 2042
rect 1750 2037 1756 2038
rect 3030 2035 3036 2036
rect 215 2031 221 2032
rect 215 2027 216 2031
rect 220 2030 221 2031
rect 290 2031 296 2032
rect 290 2030 291 2031
rect 220 2028 291 2030
rect 220 2027 221 2028
rect 215 2026 221 2027
rect 290 2027 291 2028
rect 295 2027 296 2031
rect 290 2026 296 2027
rect 359 2031 365 2032
rect 359 2027 360 2031
rect 364 2030 365 2031
rect 390 2031 396 2032
rect 390 2030 391 2031
rect 364 2028 391 2030
rect 364 2027 365 2028
rect 359 2026 365 2027
rect 390 2027 391 2028
rect 395 2027 396 2031
rect 390 2026 396 2027
rect 519 2031 525 2032
rect 519 2027 520 2031
rect 524 2030 525 2031
rect 586 2031 592 2032
rect 586 2030 587 2031
rect 524 2028 587 2030
rect 524 2027 525 2028
rect 519 2026 525 2027
rect 586 2027 587 2028
rect 591 2027 592 2031
rect 586 2026 592 2027
rect 703 2031 709 2032
rect 703 2027 704 2031
rect 708 2030 709 2031
rect 770 2031 776 2032
rect 770 2030 771 2031
rect 708 2028 771 2030
rect 708 2027 709 2028
rect 703 2026 709 2027
rect 770 2027 771 2028
rect 775 2027 776 2031
rect 770 2026 776 2027
rect 874 2031 880 2032
rect 874 2027 875 2031
rect 879 2030 880 2031
rect 895 2031 901 2032
rect 895 2030 896 2031
rect 879 2028 896 2030
rect 879 2027 880 2028
rect 874 2026 880 2027
rect 895 2027 896 2028
rect 900 2027 901 2031
rect 895 2026 901 2027
rect 1074 2031 1080 2032
rect 1074 2027 1075 2031
rect 1079 2030 1080 2031
rect 1103 2031 1109 2032
rect 1103 2030 1104 2031
rect 1079 2028 1104 2030
rect 1079 2027 1080 2028
rect 1074 2026 1080 2027
rect 1103 2027 1104 2028
rect 1108 2027 1109 2031
rect 1103 2026 1109 2027
rect 1214 2031 1220 2032
rect 1214 2027 1215 2031
rect 1219 2030 1220 2031
rect 1311 2031 1317 2032
rect 1311 2030 1312 2031
rect 1219 2028 1312 2030
rect 1219 2027 1220 2028
rect 1214 2026 1220 2027
rect 1311 2027 1312 2028
rect 1316 2027 1317 2031
rect 1311 2026 1317 2027
rect 1527 2031 1533 2032
rect 1527 2027 1528 2031
rect 1532 2030 1533 2031
rect 1602 2031 1608 2032
rect 1602 2030 1603 2031
rect 1532 2028 1603 2030
rect 1532 2027 1533 2028
rect 1527 2026 1533 2027
rect 1602 2027 1603 2028
rect 1607 2027 1608 2031
rect 1602 2026 1608 2027
rect 1743 2031 1749 2032
rect 1743 2027 1744 2031
rect 1748 2030 1749 2031
rect 1758 2031 1764 2032
rect 1758 2030 1759 2031
rect 1748 2028 1759 2030
rect 1748 2027 1749 2028
rect 1743 2026 1749 2027
rect 1758 2027 1759 2028
rect 1763 2027 1764 2031
rect 3030 2031 3031 2035
rect 3035 2034 3036 2035
rect 3087 2035 3093 2036
rect 3087 2034 3088 2035
rect 3035 2032 3088 2034
rect 3035 2031 3036 2032
rect 3030 2030 3036 2031
rect 3087 2031 3088 2032
rect 3092 2031 3093 2035
rect 3087 2030 3093 2031
rect 3518 2035 3525 2036
rect 3518 2031 3519 2035
rect 3524 2031 3525 2035
rect 3518 2030 3525 2031
rect 1758 2026 1764 2027
rect 135 2019 141 2020
rect 135 2015 136 2019
rect 140 2018 141 2019
rect 150 2019 156 2020
rect 150 2018 151 2019
rect 140 2016 151 2018
rect 140 2015 141 2016
rect 135 2014 141 2015
rect 150 2015 151 2016
rect 155 2015 156 2019
rect 150 2014 156 2015
rect 194 2019 200 2020
rect 194 2015 195 2019
rect 199 2018 200 2019
rect 255 2019 261 2020
rect 255 2018 256 2019
rect 199 2016 256 2018
rect 199 2015 200 2016
rect 194 2014 200 2015
rect 255 2015 256 2016
rect 260 2015 261 2019
rect 255 2014 261 2015
rect 314 2019 320 2020
rect 314 2015 315 2019
rect 319 2018 320 2019
rect 375 2019 381 2020
rect 375 2018 376 2019
rect 319 2016 376 2018
rect 319 2015 320 2016
rect 314 2014 320 2015
rect 375 2015 376 2016
rect 380 2015 381 2019
rect 375 2014 381 2015
rect 487 2019 493 2020
rect 487 2015 488 2019
rect 492 2018 493 2019
rect 495 2019 501 2020
rect 495 2018 496 2019
rect 492 2016 496 2018
rect 492 2015 493 2016
rect 487 2014 493 2015
rect 495 2015 496 2016
rect 500 2015 501 2019
rect 495 2014 501 2015
rect 546 2019 552 2020
rect 546 2015 547 2019
rect 551 2018 552 2019
rect 599 2019 605 2020
rect 599 2018 600 2019
rect 551 2016 600 2018
rect 551 2015 552 2016
rect 546 2014 552 2015
rect 599 2015 600 2016
rect 604 2015 605 2019
rect 599 2014 605 2015
rect 658 2019 664 2020
rect 658 2015 659 2019
rect 663 2018 664 2019
rect 711 2019 717 2020
rect 711 2018 712 2019
rect 663 2016 712 2018
rect 663 2015 664 2016
rect 658 2014 664 2015
rect 711 2015 712 2016
rect 716 2015 717 2019
rect 711 2014 717 2015
rect 815 2019 821 2020
rect 815 2015 816 2019
rect 820 2018 821 2019
rect 866 2019 872 2020
rect 866 2018 867 2019
rect 820 2016 867 2018
rect 820 2015 821 2016
rect 815 2014 821 2015
rect 866 2015 867 2016
rect 871 2015 872 2019
rect 866 2014 872 2015
rect 874 2019 880 2020
rect 874 2015 875 2019
rect 879 2018 880 2019
rect 919 2019 925 2020
rect 919 2018 920 2019
rect 879 2016 920 2018
rect 879 2015 880 2016
rect 874 2014 880 2015
rect 919 2015 920 2016
rect 924 2015 925 2019
rect 919 2014 925 2015
rect 978 2019 984 2020
rect 978 2015 979 2019
rect 983 2018 984 2019
rect 1015 2019 1021 2020
rect 1015 2018 1016 2019
rect 983 2016 1016 2018
rect 983 2015 984 2016
rect 978 2014 984 2015
rect 1015 2015 1016 2016
rect 1020 2015 1021 2019
rect 1015 2014 1021 2015
rect 1095 2019 1101 2020
rect 1095 2015 1096 2019
rect 1100 2018 1101 2019
rect 1103 2019 1109 2020
rect 1103 2018 1104 2019
rect 1100 2016 1104 2018
rect 1100 2015 1101 2016
rect 1095 2014 1101 2015
rect 1103 2015 1104 2016
rect 1108 2015 1109 2019
rect 1103 2014 1109 2015
rect 1162 2019 1168 2020
rect 1162 2015 1163 2019
rect 1167 2018 1168 2019
rect 1199 2019 1205 2020
rect 1199 2018 1200 2019
rect 1167 2016 1200 2018
rect 1167 2015 1168 2016
rect 1162 2014 1168 2015
rect 1199 2015 1200 2016
rect 1204 2015 1205 2019
rect 1199 2014 1205 2015
rect 1258 2019 1264 2020
rect 1258 2015 1259 2019
rect 1263 2018 1264 2019
rect 1287 2019 1293 2020
rect 1287 2018 1288 2019
rect 1263 2016 1288 2018
rect 1263 2015 1264 2016
rect 1258 2014 1264 2015
rect 1287 2015 1288 2016
rect 1292 2015 1293 2019
rect 1287 2014 1293 2015
rect 1346 2019 1352 2020
rect 1346 2015 1347 2019
rect 1351 2018 1352 2019
rect 1383 2019 1389 2020
rect 1383 2018 1384 2019
rect 1351 2016 1384 2018
rect 1351 2015 1352 2016
rect 1346 2014 1352 2015
rect 1383 2015 1384 2016
rect 1388 2015 1389 2019
rect 1383 2014 1389 2015
rect 1442 2019 1448 2020
rect 1442 2015 1443 2019
rect 1447 2018 1448 2019
rect 1479 2019 1485 2020
rect 1479 2018 1480 2019
rect 1447 2016 1480 2018
rect 1447 2015 1448 2016
rect 1442 2014 1448 2015
rect 1479 2015 1480 2016
rect 1484 2015 1485 2019
rect 1479 2014 1485 2015
rect 1575 2019 1581 2020
rect 1575 2015 1576 2019
rect 1580 2018 1581 2019
rect 1594 2019 1600 2020
rect 1594 2018 1595 2019
rect 1580 2016 1595 2018
rect 1580 2015 1581 2016
rect 1575 2014 1581 2015
rect 1594 2015 1595 2016
rect 1599 2015 1600 2019
rect 1594 2014 1600 2015
rect 1634 2019 1640 2020
rect 1634 2015 1635 2019
rect 1639 2018 1640 2019
rect 1663 2019 1669 2020
rect 1663 2018 1664 2019
rect 1639 2016 1664 2018
rect 1639 2015 1640 2016
rect 1634 2014 1640 2015
rect 1663 2015 1664 2016
rect 1668 2015 1669 2019
rect 1663 2014 1669 2015
rect 1722 2019 1728 2020
rect 1722 2015 1723 2019
rect 1727 2018 1728 2019
rect 1743 2019 1749 2020
rect 1743 2018 1744 2019
rect 1727 2016 1744 2018
rect 1727 2015 1728 2016
rect 1722 2014 1728 2015
rect 1743 2015 1744 2016
rect 1748 2015 1749 2019
rect 1743 2014 1749 2015
rect 142 2010 148 2011
rect 142 2006 143 2010
rect 147 2006 148 2010
rect 142 2005 148 2006
rect 262 2010 268 2011
rect 262 2006 263 2010
rect 267 2006 268 2010
rect 262 2005 268 2006
rect 382 2010 388 2011
rect 382 2006 383 2010
rect 387 2006 388 2010
rect 382 2005 388 2006
rect 494 2010 500 2011
rect 494 2006 495 2010
rect 499 2006 500 2010
rect 494 2005 500 2006
rect 606 2010 612 2011
rect 606 2006 607 2010
rect 611 2006 612 2010
rect 606 2005 612 2006
rect 718 2010 724 2011
rect 718 2006 719 2010
rect 723 2006 724 2010
rect 718 2005 724 2006
rect 822 2010 828 2011
rect 822 2006 823 2010
rect 827 2006 828 2010
rect 822 2005 828 2006
rect 926 2010 932 2011
rect 926 2006 927 2010
rect 931 2006 932 2010
rect 926 2005 932 2006
rect 1022 2010 1028 2011
rect 1022 2006 1023 2010
rect 1027 2006 1028 2010
rect 1022 2005 1028 2006
rect 1110 2010 1116 2011
rect 1110 2006 1111 2010
rect 1115 2006 1116 2010
rect 1110 2005 1116 2006
rect 1206 2010 1212 2011
rect 1206 2006 1207 2010
rect 1211 2006 1212 2010
rect 1206 2005 1212 2006
rect 1294 2010 1300 2011
rect 1294 2006 1295 2010
rect 1299 2006 1300 2010
rect 1294 2005 1300 2006
rect 1390 2010 1396 2011
rect 1390 2006 1391 2010
rect 1395 2006 1396 2010
rect 1390 2005 1396 2006
rect 1486 2010 1492 2011
rect 1486 2006 1487 2010
rect 1491 2006 1492 2010
rect 1486 2005 1492 2006
rect 1582 2010 1588 2011
rect 1582 2006 1583 2010
rect 1587 2006 1588 2010
rect 1582 2005 1588 2006
rect 1670 2010 1676 2011
rect 1670 2006 1671 2010
rect 1675 2006 1676 2010
rect 1670 2005 1676 2006
rect 1750 2010 1756 2011
rect 1750 2006 1751 2010
rect 1755 2006 1756 2010
rect 1750 2005 1756 2006
rect 2070 2004 2076 2005
rect 1870 2001 1876 2002
rect 1870 1997 1871 2001
rect 1875 1997 1876 2001
rect 2070 2000 2071 2004
rect 2075 2000 2076 2004
rect 2070 1999 2076 2000
rect 2206 2004 2212 2005
rect 2206 2000 2207 2004
rect 2211 2000 2212 2004
rect 2206 1999 2212 2000
rect 2358 2004 2364 2005
rect 2358 2000 2359 2004
rect 2363 2000 2364 2004
rect 2358 1999 2364 2000
rect 2518 2004 2524 2005
rect 2518 2000 2519 2004
rect 2523 2000 2524 2004
rect 2518 1999 2524 2000
rect 2678 2004 2684 2005
rect 2678 2000 2679 2004
rect 2683 2000 2684 2004
rect 2678 1999 2684 2000
rect 2846 2004 2852 2005
rect 2846 2000 2847 2004
rect 2851 2000 2852 2004
rect 2846 1999 2852 2000
rect 3014 2004 3020 2005
rect 3014 2000 3015 2004
rect 3019 2000 3020 2004
rect 3014 1999 3020 2000
rect 3182 2004 3188 2005
rect 3182 2000 3183 2004
rect 3187 2000 3188 2004
rect 3182 1999 3188 2000
rect 3350 2004 3356 2005
rect 3350 2000 3351 2004
rect 3355 2000 3356 2004
rect 3350 1999 3356 2000
rect 3502 2004 3508 2005
rect 3502 2000 3503 2004
rect 3507 2000 3508 2004
rect 3502 1999 3508 2000
rect 3590 2001 3596 2002
rect 1870 1996 1876 1997
rect 3590 1997 3591 2001
rect 3595 1997 3596 2001
rect 3590 1996 3596 1997
rect 2146 1995 2152 1996
rect 2146 1994 2147 1995
rect 110 1992 116 1993
rect 110 1988 111 1992
rect 115 1988 116 1992
rect 110 1987 116 1988
rect 1830 1992 1836 1993
rect 2133 1992 2147 1994
rect 1830 1988 1831 1992
rect 1835 1988 1836 1992
rect 2146 1991 2147 1992
rect 2151 1991 2152 1995
rect 2274 1995 2280 1996
rect 2274 1994 2275 1995
rect 2269 1992 2275 1994
rect 2146 1990 2152 1991
rect 2274 1991 2275 1992
rect 2279 1991 2280 1995
rect 2446 1995 2452 1996
rect 2446 1994 2447 1995
rect 2421 1992 2447 1994
rect 2274 1990 2280 1991
rect 2446 1991 2447 1992
rect 2451 1991 2452 1995
rect 2446 1990 2452 1991
rect 2454 1995 2460 1996
rect 2454 1991 2455 1995
rect 2459 1994 2460 1995
rect 2598 1995 2604 1996
rect 2459 1992 2537 1994
rect 2459 1991 2460 1992
rect 2454 1990 2460 1991
rect 2598 1991 2599 1995
rect 2603 1994 2604 1995
rect 2746 1995 2752 1996
rect 2603 1992 2697 1994
rect 2603 1991 2604 1992
rect 2598 1990 2604 1991
rect 2746 1991 2747 1995
rect 2751 1994 2752 1995
rect 2914 1995 2920 1996
rect 2751 1992 2865 1994
rect 2751 1991 2752 1992
rect 2746 1990 2752 1991
rect 2914 1991 2915 1995
rect 2919 1994 2920 1995
rect 3274 1995 3280 1996
rect 3274 1994 3275 1995
rect 2919 1992 3033 1994
rect 3245 1992 3275 1994
rect 2919 1991 2920 1992
rect 2914 1990 2920 1991
rect 3274 1991 3275 1992
rect 3279 1991 3280 1995
rect 3430 1995 3436 1996
rect 3430 1994 3431 1995
rect 3413 1992 3431 1994
rect 3274 1990 3280 1991
rect 3430 1991 3431 1992
rect 3435 1991 3436 1995
rect 3430 1990 3436 1991
rect 1830 1987 1836 1988
rect 3262 1987 3268 1988
rect 1870 1984 1876 1985
rect 194 1983 200 1984
rect 194 1979 195 1983
rect 199 1979 200 1983
rect 194 1978 200 1979
rect 314 1983 320 1984
rect 314 1979 315 1983
rect 319 1979 320 1983
rect 314 1978 320 1979
rect 390 1983 396 1984
rect 390 1979 391 1983
rect 395 1979 396 1983
rect 390 1978 396 1979
rect 546 1983 552 1984
rect 546 1979 547 1983
rect 551 1979 552 1983
rect 546 1978 552 1979
rect 658 1983 664 1984
rect 658 1979 659 1983
rect 663 1979 664 1983
rect 658 1978 664 1979
rect 770 1983 776 1984
rect 770 1979 771 1983
rect 775 1979 776 1983
rect 770 1978 776 1979
rect 874 1983 880 1984
rect 874 1979 875 1983
rect 879 1979 880 1983
rect 874 1978 880 1979
rect 978 1983 984 1984
rect 978 1979 979 1983
rect 983 1979 984 1983
rect 978 1978 984 1979
rect 1074 1983 1080 1984
rect 1074 1979 1075 1983
rect 1079 1979 1080 1983
rect 1074 1978 1080 1979
rect 1162 1983 1168 1984
rect 1162 1979 1163 1983
rect 1167 1979 1168 1983
rect 1162 1978 1168 1979
rect 1258 1983 1264 1984
rect 1258 1979 1259 1983
rect 1263 1979 1264 1983
rect 1258 1978 1264 1979
rect 1346 1983 1352 1984
rect 1346 1979 1347 1983
rect 1351 1979 1352 1983
rect 1346 1978 1352 1979
rect 1442 1983 1448 1984
rect 1442 1979 1443 1983
rect 1447 1979 1448 1983
rect 1442 1978 1448 1979
rect 1634 1983 1640 1984
rect 1634 1979 1635 1983
rect 1639 1979 1640 1983
rect 1634 1978 1640 1979
rect 1722 1983 1728 1984
rect 1722 1979 1723 1983
rect 1727 1979 1728 1983
rect 1870 1980 1871 1984
rect 1875 1980 1876 1984
rect 3262 1983 3263 1987
rect 3267 1986 3268 1987
rect 3520 1986 3522 1993
rect 3267 1984 3522 1986
rect 3590 1984 3596 1985
rect 3267 1983 3268 1984
rect 3262 1982 3268 1983
rect 1870 1979 1876 1980
rect 3590 1980 3591 1984
rect 3595 1980 3596 1984
rect 3590 1979 3596 1980
rect 1722 1978 1728 1979
rect 110 1975 116 1976
rect 110 1971 111 1975
rect 115 1971 116 1975
rect 1830 1975 1836 1976
rect 110 1970 116 1971
rect 134 1972 140 1973
rect 134 1968 135 1972
rect 139 1968 140 1972
rect 134 1967 140 1968
rect 254 1972 260 1973
rect 254 1968 255 1972
rect 259 1968 260 1972
rect 254 1967 260 1968
rect 374 1972 380 1973
rect 374 1968 375 1972
rect 379 1968 380 1972
rect 374 1967 380 1968
rect 486 1972 492 1973
rect 486 1968 487 1972
rect 491 1968 492 1972
rect 486 1967 492 1968
rect 598 1972 604 1973
rect 598 1968 599 1972
rect 603 1968 604 1972
rect 598 1967 604 1968
rect 710 1972 716 1973
rect 710 1968 711 1972
rect 715 1968 716 1972
rect 710 1967 716 1968
rect 814 1972 820 1973
rect 814 1968 815 1972
rect 819 1968 820 1972
rect 814 1967 820 1968
rect 918 1972 924 1973
rect 918 1968 919 1972
rect 923 1968 924 1972
rect 918 1967 924 1968
rect 1014 1972 1020 1973
rect 1014 1968 1015 1972
rect 1019 1968 1020 1972
rect 1014 1967 1020 1968
rect 1102 1972 1108 1973
rect 1102 1968 1103 1972
rect 1107 1968 1108 1972
rect 1102 1967 1108 1968
rect 1198 1972 1204 1973
rect 1198 1968 1199 1972
rect 1203 1968 1204 1972
rect 1198 1967 1204 1968
rect 1286 1972 1292 1973
rect 1286 1968 1287 1972
rect 1291 1968 1292 1972
rect 1286 1967 1292 1968
rect 1382 1972 1388 1973
rect 1382 1968 1383 1972
rect 1387 1968 1388 1972
rect 1382 1967 1388 1968
rect 1478 1972 1484 1973
rect 1478 1968 1479 1972
rect 1483 1968 1484 1972
rect 1478 1967 1484 1968
rect 1574 1972 1580 1973
rect 1574 1968 1575 1972
rect 1579 1968 1580 1972
rect 1574 1967 1580 1968
rect 1662 1972 1668 1973
rect 1662 1968 1663 1972
rect 1667 1968 1668 1972
rect 1662 1967 1668 1968
rect 1742 1972 1748 1973
rect 1742 1968 1743 1972
rect 1747 1968 1748 1972
rect 1830 1971 1831 1975
rect 1835 1971 1836 1975
rect 1830 1970 1836 1971
rect 1742 1967 1748 1968
rect 2078 1966 2084 1967
rect 2078 1962 2079 1966
rect 2083 1962 2084 1966
rect 2078 1961 2084 1962
rect 2214 1966 2220 1967
rect 2214 1962 2215 1966
rect 2219 1962 2220 1966
rect 2214 1961 2220 1962
rect 2366 1966 2372 1967
rect 2366 1962 2367 1966
rect 2371 1962 2372 1966
rect 2366 1961 2372 1962
rect 2526 1966 2532 1967
rect 2526 1962 2527 1966
rect 2531 1962 2532 1966
rect 2526 1961 2532 1962
rect 2686 1966 2692 1967
rect 2686 1962 2687 1966
rect 2691 1962 2692 1966
rect 2686 1961 2692 1962
rect 2854 1966 2860 1967
rect 2854 1962 2855 1966
rect 2859 1962 2860 1966
rect 2854 1961 2860 1962
rect 3022 1966 3028 1967
rect 3022 1962 3023 1966
rect 3027 1962 3028 1966
rect 3022 1961 3028 1962
rect 3190 1966 3196 1967
rect 3190 1962 3191 1966
rect 3195 1962 3196 1966
rect 3190 1961 3196 1962
rect 3358 1966 3364 1967
rect 3358 1962 3359 1966
rect 3363 1962 3364 1966
rect 3358 1961 3364 1962
rect 3510 1966 3516 1967
rect 3510 1962 3511 1966
rect 3515 1962 3516 1966
rect 3510 1961 3516 1962
rect 1230 1955 1236 1956
rect 1230 1951 1231 1955
rect 1235 1954 1236 1955
rect 1495 1955 1501 1956
rect 1495 1954 1496 1955
rect 1235 1952 1496 1954
rect 1235 1951 1236 1952
rect 1230 1950 1236 1951
rect 1495 1951 1496 1952
rect 1500 1951 1501 1955
rect 1495 1950 1501 1951
rect 1758 1955 1765 1956
rect 1758 1951 1759 1955
rect 1764 1951 1765 1955
rect 1758 1950 1765 1951
rect 2058 1955 2064 1956
rect 2058 1951 2059 1955
rect 2063 1954 2064 1955
rect 2071 1955 2077 1956
rect 2071 1954 2072 1955
rect 2063 1952 2072 1954
rect 2063 1951 2064 1952
rect 2058 1950 2064 1951
rect 2071 1951 2072 1952
rect 2076 1951 2077 1955
rect 2071 1950 2077 1951
rect 2146 1955 2152 1956
rect 2146 1951 2147 1955
rect 2151 1954 2152 1955
rect 2207 1955 2213 1956
rect 2207 1954 2208 1955
rect 2151 1952 2208 1954
rect 2151 1951 2152 1952
rect 2146 1950 2152 1951
rect 2207 1951 2208 1952
rect 2212 1951 2213 1955
rect 2207 1950 2213 1951
rect 2274 1955 2280 1956
rect 2274 1951 2275 1955
rect 2279 1954 2280 1955
rect 2359 1955 2365 1956
rect 2359 1954 2360 1955
rect 2279 1952 2360 1954
rect 2279 1951 2280 1952
rect 2274 1950 2280 1951
rect 2359 1951 2360 1952
rect 2364 1951 2365 1955
rect 2359 1950 2365 1951
rect 2446 1955 2452 1956
rect 2446 1951 2447 1955
rect 2451 1954 2452 1955
rect 2519 1955 2525 1956
rect 2519 1954 2520 1955
rect 2451 1952 2520 1954
rect 2451 1951 2452 1952
rect 2446 1950 2452 1951
rect 2519 1951 2520 1952
rect 2524 1951 2525 1955
rect 2519 1950 2525 1951
rect 2679 1955 2685 1956
rect 2679 1951 2680 1955
rect 2684 1954 2685 1955
rect 2746 1955 2752 1956
rect 2746 1954 2747 1955
rect 2684 1952 2747 1954
rect 2684 1951 2685 1952
rect 2679 1950 2685 1951
rect 2746 1951 2747 1952
rect 2751 1951 2752 1955
rect 2746 1950 2752 1951
rect 2847 1955 2853 1956
rect 2847 1951 2848 1955
rect 2852 1954 2853 1955
rect 2914 1955 2920 1956
rect 2914 1954 2915 1955
rect 2852 1952 2915 1954
rect 2852 1951 2853 1952
rect 2847 1950 2853 1951
rect 2914 1951 2915 1952
rect 2919 1951 2920 1955
rect 2914 1950 2920 1951
rect 3015 1955 3021 1956
rect 3015 1951 3016 1955
rect 3020 1954 3021 1955
rect 3030 1955 3036 1956
rect 3030 1954 3031 1955
rect 3020 1952 3031 1954
rect 3020 1951 3021 1952
rect 3015 1950 3021 1951
rect 3030 1951 3031 1952
rect 3035 1951 3036 1955
rect 3030 1950 3036 1951
rect 3183 1955 3189 1956
rect 3183 1951 3184 1955
rect 3188 1954 3189 1955
rect 3262 1955 3268 1956
rect 3262 1954 3263 1955
rect 3188 1952 3263 1954
rect 3188 1951 3189 1952
rect 3183 1950 3189 1951
rect 3262 1951 3263 1952
rect 3267 1951 3268 1955
rect 3262 1950 3268 1951
rect 3274 1955 3280 1956
rect 3274 1951 3275 1955
rect 3279 1954 3280 1955
rect 3351 1955 3357 1956
rect 3351 1954 3352 1955
rect 3279 1952 3352 1954
rect 3279 1951 3280 1952
rect 3274 1950 3280 1951
rect 3351 1951 3352 1952
rect 3356 1951 3357 1955
rect 3351 1950 3357 1951
rect 3503 1955 3509 1956
rect 3503 1951 3504 1955
rect 3508 1954 3509 1955
rect 3518 1955 3524 1956
rect 3518 1954 3519 1955
rect 3508 1952 3519 1954
rect 3508 1951 3509 1952
rect 3503 1950 3509 1951
rect 3518 1951 3519 1952
rect 3523 1951 3524 1955
rect 3518 1950 3524 1951
rect 1810 1943 1816 1944
rect 1810 1939 1811 1943
rect 1815 1942 1816 1943
rect 1895 1943 1901 1944
rect 1895 1942 1896 1943
rect 1815 1940 1896 1942
rect 1815 1939 1816 1940
rect 1810 1938 1816 1939
rect 1895 1939 1896 1940
rect 1900 1939 1901 1943
rect 1895 1938 1901 1939
rect 1999 1943 2005 1944
rect 1999 1939 2000 1943
rect 2004 1942 2005 1943
rect 2066 1943 2072 1944
rect 2066 1942 2067 1943
rect 2004 1940 2067 1942
rect 2004 1939 2005 1940
rect 1999 1938 2005 1939
rect 2066 1939 2067 1940
rect 2071 1939 2072 1943
rect 2066 1938 2072 1939
rect 2127 1943 2133 1944
rect 2127 1939 2128 1943
rect 2132 1942 2133 1943
rect 2194 1943 2200 1944
rect 2194 1942 2195 1943
rect 2132 1940 2195 1942
rect 2132 1939 2133 1940
rect 2127 1938 2133 1939
rect 2194 1939 2195 1940
rect 2199 1939 2200 1943
rect 2194 1938 2200 1939
rect 2247 1943 2253 1944
rect 2247 1939 2248 1943
rect 2252 1942 2253 1943
rect 2350 1943 2356 1944
rect 2350 1942 2351 1943
rect 2252 1940 2351 1942
rect 2252 1939 2253 1940
rect 2247 1938 2253 1939
rect 2350 1939 2351 1940
rect 2355 1939 2356 1943
rect 2350 1938 2356 1939
rect 2367 1943 2373 1944
rect 2367 1939 2368 1943
rect 2372 1942 2373 1943
rect 2382 1943 2388 1944
rect 2382 1942 2383 1943
rect 2372 1940 2383 1942
rect 2372 1939 2373 1940
rect 2367 1938 2373 1939
rect 2382 1939 2383 1940
rect 2387 1939 2388 1943
rect 2382 1938 2388 1939
rect 2426 1943 2432 1944
rect 2426 1939 2427 1943
rect 2431 1942 2432 1943
rect 2479 1943 2485 1944
rect 2479 1942 2480 1943
rect 2431 1940 2480 1942
rect 2431 1939 2432 1940
rect 2426 1938 2432 1939
rect 2479 1939 2480 1940
rect 2484 1939 2485 1943
rect 2479 1938 2485 1939
rect 2538 1943 2544 1944
rect 2538 1939 2539 1943
rect 2543 1942 2544 1943
rect 2591 1943 2597 1944
rect 2591 1942 2592 1943
rect 2543 1940 2592 1942
rect 2543 1939 2544 1940
rect 2538 1938 2544 1939
rect 2591 1939 2592 1940
rect 2596 1939 2597 1943
rect 2591 1938 2597 1939
rect 2650 1943 2656 1944
rect 2650 1939 2651 1943
rect 2655 1942 2656 1943
rect 2711 1943 2717 1944
rect 2711 1942 2712 1943
rect 2655 1940 2712 1942
rect 2655 1939 2656 1940
rect 2650 1938 2656 1939
rect 2711 1939 2712 1940
rect 2716 1939 2717 1943
rect 2711 1938 2717 1939
rect 2770 1943 2776 1944
rect 2770 1939 2771 1943
rect 2775 1942 2776 1943
rect 2831 1943 2837 1944
rect 2831 1942 2832 1943
rect 2775 1940 2832 1942
rect 2775 1939 2776 1940
rect 2770 1938 2776 1939
rect 2831 1939 2832 1940
rect 2836 1939 2837 1943
rect 2831 1938 2837 1939
rect 1902 1934 1908 1935
rect 1902 1930 1903 1934
rect 1907 1930 1908 1934
rect 1902 1929 1908 1930
rect 2006 1934 2012 1935
rect 2006 1930 2007 1934
rect 2011 1930 2012 1934
rect 2006 1929 2012 1930
rect 2134 1934 2140 1935
rect 2134 1930 2135 1934
rect 2139 1930 2140 1934
rect 2134 1929 2140 1930
rect 2254 1934 2260 1935
rect 2254 1930 2255 1934
rect 2259 1930 2260 1934
rect 2254 1929 2260 1930
rect 2374 1934 2380 1935
rect 2374 1930 2375 1934
rect 2379 1930 2380 1934
rect 2374 1929 2380 1930
rect 2486 1934 2492 1935
rect 2486 1930 2487 1934
rect 2491 1930 2492 1934
rect 2486 1929 2492 1930
rect 2598 1934 2604 1935
rect 2598 1930 2599 1934
rect 2603 1930 2604 1934
rect 2598 1929 2604 1930
rect 2718 1934 2724 1935
rect 2718 1930 2719 1934
rect 2723 1930 2724 1934
rect 2718 1929 2724 1930
rect 2838 1934 2844 1935
rect 2838 1930 2839 1934
rect 2843 1930 2844 1934
rect 2838 1929 2844 1930
rect 166 1920 172 1921
rect 110 1917 116 1918
rect 110 1913 111 1917
rect 115 1913 116 1917
rect 166 1916 167 1920
rect 171 1916 172 1920
rect 166 1915 172 1916
rect 326 1920 332 1921
rect 326 1916 327 1920
rect 331 1916 332 1920
rect 326 1915 332 1916
rect 486 1920 492 1921
rect 486 1916 487 1920
rect 491 1916 492 1920
rect 486 1915 492 1916
rect 646 1920 652 1921
rect 646 1916 647 1920
rect 651 1916 652 1920
rect 646 1915 652 1916
rect 798 1920 804 1921
rect 798 1916 799 1920
rect 803 1916 804 1920
rect 798 1915 804 1916
rect 942 1920 948 1921
rect 942 1916 943 1920
rect 947 1916 948 1920
rect 942 1915 948 1916
rect 1078 1920 1084 1921
rect 1078 1916 1079 1920
rect 1083 1916 1084 1920
rect 1078 1915 1084 1916
rect 1214 1920 1220 1921
rect 1214 1916 1215 1920
rect 1219 1916 1220 1920
rect 1214 1915 1220 1916
rect 1350 1920 1356 1921
rect 1350 1916 1351 1920
rect 1355 1916 1356 1920
rect 1350 1915 1356 1916
rect 1486 1920 1492 1921
rect 1486 1916 1487 1920
rect 1491 1916 1492 1920
rect 1486 1915 1492 1916
rect 1622 1920 1628 1921
rect 1622 1916 1623 1920
rect 1627 1916 1628 1920
rect 1622 1915 1628 1916
rect 1742 1920 1748 1921
rect 1742 1916 1743 1920
rect 1747 1916 1748 1920
rect 1742 1915 1748 1916
rect 1830 1917 1836 1918
rect 110 1912 116 1913
rect 1830 1913 1831 1917
rect 1835 1913 1836 1917
rect 1830 1912 1836 1913
rect 1870 1916 1876 1917
rect 1870 1912 1871 1916
rect 1875 1912 1876 1916
rect 150 1911 156 1912
rect 150 1907 151 1911
rect 155 1910 156 1911
rect 234 1911 240 1912
rect 155 1908 185 1910
rect 155 1907 156 1908
rect 150 1906 156 1907
rect 234 1907 235 1911
rect 239 1910 240 1911
rect 554 1911 560 1912
rect 554 1910 555 1911
rect 239 1908 345 1910
rect 549 1908 555 1910
rect 239 1907 240 1908
rect 234 1906 240 1907
rect 554 1907 555 1908
rect 559 1907 560 1911
rect 554 1906 560 1907
rect 562 1911 568 1912
rect 562 1907 563 1911
rect 567 1910 568 1911
rect 714 1911 720 1912
rect 567 1908 665 1910
rect 567 1907 568 1908
rect 562 1906 568 1907
rect 714 1907 715 1911
rect 719 1910 720 1911
rect 866 1911 872 1912
rect 719 1908 817 1910
rect 719 1907 720 1908
rect 714 1906 720 1907
rect 866 1907 867 1911
rect 871 1910 872 1911
rect 1010 1911 1016 1912
rect 871 1908 961 1910
rect 871 1907 872 1908
rect 866 1906 872 1907
rect 1010 1907 1011 1911
rect 1015 1910 1016 1911
rect 1290 1911 1296 1912
rect 1290 1910 1291 1911
rect 1015 1908 1097 1910
rect 1277 1908 1291 1910
rect 1015 1907 1016 1908
rect 1010 1906 1016 1907
rect 1290 1907 1291 1908
rect 1295 1907 1296 1911
rect 1418 1911 1424 1912
rect 1418 1910 1419 1911
rect 1413 1908 1419 1910
rect 1290 1906 1296 1907
rect 1418 1907 1419 1908
rect 1423 1907 1424 1911
rect 1554 1911 1560 1912
rect 1554 1910 1555 1911
rect 1549 1908 1555 1910
rect 1418 1906 1424 1907
rect 1554 1907 1555 1908
rect 1559 1907 1560 1911
rect 1810 1911 1816 1912
rect 1870 1911 1876 1912
rect 3590 1916 3596 1917
rect 3590 1912 3591 1916
rect 3595 1912 3596 1916
rect 3590 1911 3596 1912
rect 1810 1910 1811 1911
rect 1554 1906 1560 1907
rect 1342 1903 1348 1904
rect 110 1900 116 1901
rect 110 1896 111 1900
rect 115 1896 116 1900
rect 1342 1899 1343 1903
rect 1347 1902 1348 1903
rect 1640 1902 1642 1909
rect 1805 1908 1811 1910
rect 1810 1907 1811 1908
rect 1815 1907 1816 1911
rect 1810 1906 1816 1907
rect 2058 1907 2064 1908
rect 2058 1903 2059 1907
rect 2063 1903 2064 1907
rect 2058 1902 2064 1903
rect 2066 1907 2072 1908
rect 2066 1903 2067 1907
rect 2071 1906 2072 1907
rect 2194 1907 2200 1908
rect 2071 1904 2145 1906
rect 2071 1903 2072 1904
rect 2066 1902 2072 1903
rect 2194 1903 2195 1907
rect 2199 1906 2200 1907
rect 2426 1907 2432 1908
rect 2199 1904 2265 1906
rect 2199 1903 2200 1904
rect 2194 1902 2200 1903
rect 2426 1903 2427 1907
rect 2431 1903 2432 1907
rect 2426 1902 2432 1903
rect 2538 1907 2544 1908
rect 2538 1903 2539 1907
rect 2543 1903 2544 1907
rect 2538 1902 2544 1903
rect 2650 1907 2656 1908
rect 2650 1903 2651 1907
rect 2655 1903 2656 1907
rect 2650 1902 2656 1903
rect 2770 1907 2776 1908
rect 2770 1903 2771 1907
rect 2775 1903 2776 1907
rect 2770 1902 2776 1903
rect 1347 1900 1642 1902
rect 1830 1900 1836 1901
rect 1347 1899 1348 1900
rect 1342 1898 1348 1899
rect 110 1895 116 1896
rect 1830 1896 1831 1900
rect 1835 1896 1836 1900
rect 1830 1895 1836 1896
rect 1870 1899 1876 1900
rect 1870 1895 1871 1899
rect 1875 1895 1876 1899
rect 3590 1899 3596 1900
rect 1870 1894 1876 1895
rect 1894 1896 1900 1897
rect 1894 1892 1895 1896
rect 1899 1892 1900 1896
rect 1894 1891 1900 1892
rect 1998 1896 2004 1897
rect 1998 1892 1999 1896
rect 2003 1892 2004 1896
rect 1998 1891 2004 1892
rect 2126 1896 2132 1897
rect 2126 1892 2127 1896
rect 2131 1892 2132 1896
rect 2126 1891 2132 1892
rect 2246 1896 2252 1897
rect 2246 1892 2247 1896
rect 2251 1892 2252 1896
rect 2246 1891 2252 1892
rect 2366 1896 2372 1897
rect 2366 1892 2367 1896
rect 2371 1892 2372 1896
rect 2366 1891 2372 1892
rect 2478 1896 2484 1897
rect 2478 1892 2479 1896
rect 2483 1892 2484 1896
rect 2478 1891 2484 1892
rect 2590 1896 2596 1897
rect 2590 1892 2591 1896
rect 2595 1892 2596 1896
rect 2590 1891 2596 1892
rect 2710 1896 2716 1897
rect 2710 1892 2711 1896
rect 2715 1892 2716 1896
rect 2710 1891 2716 1892
rect 2830 1896 2836 1897
rect 2830 1892 2831 1896
rect 2835 1892 2836 1896
rect 3590 1895 3591 1899
rect 3595 1895 3596 1899
rect 3590 1894 3596 1895
rect 2830 1891 2836 1892
rect 174 1882 180 1883
rect 174 1878 175 1882
rect 179 1878 180 1882
rect 174 1877 180 1878
rect 334 1882 340 1883
rect 334 1878 335 1882
rect 339 1878 340 1882
rect 334 1877 340 1878
rect 494 1882 500 1883
rect 494 1878 495 1882
rect 499 1878 500 1882
rect 494 1877 500 1878
rect 654 1882 660 1883
rect 654 1878 655 1882
rect 659 1878 660 1882
rect 654 1877 660 1878
rect 806 1882 812 1883
rect 806 1878 807 1882
rect 811 1878 812 1882
rect 806 1877 812 1878
rect 950 1882 956 1883
rect 950 1878 951 1882
rect 955 1878 956 1882
rect 950 1877 956 1878
rect 1086 1882 1092 1883
rect 1086 1878 1087 1882
rect 1091 1878 1092 1882
rect 1086 1877 1092 1878
rect 1222 1882 1228 1883
rect 1222 1878 1223 1882
rect 1227 1878 1228 1882
rect 1222 1877 1228 1878
rect 1358 1882 1364 1883
rect 1358 1878 1359 1882
rect 1363 1878 1364 1882
rect 1358 1877 1364 1878
rect 1494 1882 1500 1883
rect 1494 1878 1495 1882
rect 1499 1878 1500 1882
rect 1494 1877 1500 1878
rect 1630 1882 1636 1883
rect 1630 1878 1631 1882
rect 1635 1878 1636 1882
rect 1630 1877 1636 1878
rect 1750 1882 1756 1883
rect 1750 1878 1751 1882
rect 1755 1878 1756 1882
rect 1750 1877 1756 1878
rect 1910 1879 1917 1880
rect 1910 1875 1911 1879
rect 1916 1875 1917 1879
rect 1910 1874 1917 1875
rect 2534 1879 2540 1880
rect 2534 1875 2535 1879
rect 2539 1878 2540 1879
rect 2847 1879 2853 1880
rect 2847 1878 2848 1879
rect 2539 1876 2848 1878
rect 2539 1875 2540 1876
rect 2534 1874 2540 1875
rect 2847 1875 2848 1876
rect 2852 1875 2853 1879
rect 2847 1874 2853 1875
rect 167 1871 173 1872
rect 167 1867 168 1871
rect 172 1870 173 1871
rect 234 1871 240 1872
rect 234 1870 235 1871
rect 172 1868 235 1870
rect 172 1867 173 1868
rect 167 1866 173 1867
rect 234 1867 235 1868
rect 239 1867 240 1871
rect 234 1866 240 1867
rect 326 1871 333 1872
rect 326 1867 327 1871
rect 332 1867 333 1871
rect 326 1866 333 1867
rect 487 1871 493 1872
rect 487 1867 488 1871
rect 492 1870 493 1871
rect 562 1871 568 1872
rect 562 1870 563 1871
rect 492 1868 563 1870
rect 492 1867 493 1868
rect 487 1866 493 1867
rect 562 1867 563 1868
rect 567 1867 568 1871
rect 562 1866 568 1867
rect 647 1871 653 1872
rect 647 1867 648 1871
rect 652 1870 653 1871
rect 714 1871 720 1872
rect 714 1870 715 1871
rect 652 1868 715 1870
rect 652 1867 653 1868
rect 647 1866 653 1867
rect 714 1867 715 1868
rect 719 1867 720 1871
rect 714 1866 720 1867
rect 770 1871 776 1872
rect 770 1867 771 1871
rect 775 1870 776 1871
rect 799 1871 805 1872
rect 799 1870 800 1871
rect 775 1868 800 1870
rect 775 1867 776 1868
rect 770 1866 776 1867
rect 799 1867 800 1868
rect 804 1867 805 1871
rect 799 1866 805 1867
rect 943 1871 949 1872
rect 943 1867 944 1871
rect 948 1870 949 1871
rect 1010 1871 1016 1872
rect 1010 1870 1011 1871
rect 948 1868 1011 1870
rect 948 1867 949 1868
rect 943 1866 949 1867
rect 1010 1867 1011 1868
rect 1015 1867 1016 1871
rect 1010 1866 1016 1867
rect 1078 1871 1085 1872
rect 1078 1867 1079 1871
rect 1084 1867 1085 1871
rect 1078 1866 1085 1867
rect 1215 1871 1221 1872
rect 1215 1867 1216 1871
rect 1220 1870 1221 1871
rect 1230 1871 1236 1872
rect 1230 1870 1231 1871
rect 1220 1868 1231 1870
rect 1220 1867 1221 1868
rect 1215 1866 1221 1867
rect 1230 1867 1231 1868
rect 1235 1867 1236 1871
rect 1230 1866 1236 1867
rect 1290 1871 1296 1872
rect 1290 1867 1291 1871
rect 1295 1870 1296 1871
rect 1351 1871 1357 1872
rect 1351 1870 1352 1871
rect 1295 1868 1352 1870
rect 1295 1867 1296 1868
rect 1290 1866 1296 1867
rect 1351 1867 1352 1868
rect 1356 1867 1357 1871
rect 1351 1866 1357 1867
rect 1418 1871 1424 1872
rect 1418 1867 1419 1871
rect 1423 1870 1424 1871
rect 1487 1871 1493 1872
rect 1487 1870 1488 1871
rect 1423 1868 1488 1870
rect 1423 1867 1424 1868
rect 1418 1866 1424 1867
rect 1487 1867 1488 1868
rect 1492 1867 1493 1871
rect 1487 1866 1493 1867
rect 1554 1871 1560 1872
rect 1554 1867 1555 1871
rect 1559 1870 1560 1871
rect 1623 1871 1629 1872
rect 1623 1870 1624 1871
rect 1559 1868 1624 1870
rect 1559 1867 1560 1868
rect 1554 1866 1560 1867
rect 1623 1867 1624 1868
rect 1628 1867 1629 1871
rect 1623 1866 1629 1867
rect 1743 1871 1749 1872
rect 1743 1867 1744 1871
rect 1748 1870 1749 1871
rect 1758 1871 1764 1872
rect 1758 1870 1759 1871
rect 1748 1868 1759 1870
rect 1748 1867 1749 1868
rect 1743 1866 1749 1867
rect 1758 1867 1759 1868
rect 1763 1867 1764 1871
rect 1758 1866 1764 1867
rect 151 1859 157 1860
rect 151 1855 152 1859
rect 156 1858 157 1859
rect 182 1859 188 1860
rect 182 1858 183 1859
rect 156 1856 183 1858
rect 156 1855 157 1856
rect 151 1854 157 1855
rect 182 1855 183 1856
rect 187 1855 188 1859
rect 182 1854 188 1855
rect 210 1859 216 1860
rect 210 1855 211 1859
rect 215 1858 216 1859
rect 295 1859 301 1860
rect 295 1858 296 1859
rect 215 1856 296 1858
rect 215 1855 216 1856
rect 210 1854 216 1855
rect 295 1855 296 1856
rect 300 1855 301 1859
rect 295 1854 301 1855
rect 430 1859 436 1860
rect 430 1855 431 1859
rect 435 1858 436 1859
rect 439 1859 445 1860
rect 439 1858 440 1859
rect 435 1856 440 1858
rect 435 1855 436 1856
rect 430 1854 436 1855
rect 439 1855 440 1856
rect 444 1855 445 1859
rect 439 1854 445 1855
rect 554 1859 560 1860
rect 554 1855 555 1859
rect 559 1858 560 1859
rect 591 1859 597 1860
rect 591 1858 592 1859
rect 559 1856 592 1858
rect 559 1855 560 1856
rect 554 1854 560 1855
rect 591 1855 592 1856
rect 596 1855 597 1859
rect 591 1854 597 1855
rect 679 1859 685 1860
rect 679 1855 680 1859
rect 684 1858 685 1859
rect 743 1859 749 1860
rect 743 1858 744 1859
rect 684 1856 744 1858
rect 684 1855 685 1856
rect 679 1854 685 1855
rect 743 1855 744 1856
rect 748 1855 749 1859
rect 743 1854 749 1855
rect 838 1859 844 1860
rect 838 1855 839 1859
rect 843 1858 844 1859
rect 895 1859 901 1860
rect 895 1858 896 1859
rect 843 1856 896 1858
rect 843 1855 844 1856
rect 838 1854 844 1855
rect 895 1855 896 1856
rect 900 1855 901 1859
rect 895 1854 901 1855
rect 1047 1859 1053 1860
rect 1047 1855 1048 1859
rect 1052 1858 1053 1859
rect 1127 1859 1133 1860
rect 1127 1858 1128 1859
rect 1052 1856 1128 1858
rect 1052 1855 1053 1856
rect 1047 1854 1053 1855
rect 1127 1855 1128 1856
rect 1132 1855 1133 1859
rect 1127 1854 1133 1855
rect 1198 1859 1205 1860
rect 1198 1855 1199 1859
rect 1204 1855 1205 1859
rect 1198 1854 1205 1855
rect 1342 1859 1349 1860
rect 1342 1855 1343 1859
rect 1348 1855 1349 1859
rect 1342 1854 1349 1855
rect 1402 1859 1408 1860
rect 1402 1855 1403 1859
rect 1407 1858 1408 1859
rect 1479 1859 1485 1860
rect 1479 1858 1480 1859
rect 1407 1856 1480 1858
rect 1407 1855 1408 1856
rect 1402 1854 1408 1855
rect 1479 1855 1480 1856
rect 1484 1855 1485 1859
rect 1479 1854 1485 1855
rect 1538 1859 1544 1860
rect 1538 1855 1539 1859
rect 1543 1858 1544 1859
rect 1623 1859 1629 1860
rect 1623 1858 1624 1859
rect 1543 1856 1624 1858
rect 1543 1855 1544 1856
rect 1538 1854 1544 1855
rect 1623 1855 1624 1856
rect 1628 1855 1629 1859
rect 1623 1854 1629 1855
rect 1682 1859 1688 1860
rect 1682 1855 1683 1859
rect 1687 1858 1688 1859
rect 1743 1859 1749 1860
rect 1743 1858 1744 1859
rect 1687 1856 1744 1858
rect 1687 1855 1688 1856
rect 1682 1854 1688 1855
rect 1743 1855 1744 1856
rect 1748 1855 1749 1859
rect 1743 1854 1749 1855
rect 1894 1852 1900 1853
rect 158 1850 164 1851
rect 158 1846 159 1850
rect 163 1846 164 1850
rect 158 1845 164 1846
rect 302 1850 308 1851
rect 302 1846 303 1850
rect 307 1846 308 1850
rect 302 1845 308 1846
rect 446 1850 452 1851
rect 446 1846 447 1850
rect 451 1846 452 1850
rect 446 1845 452 1846
rect 598 1850 604 1851
rect 598 1846 599 1850
rect 603 1846 604 1850
rect 598 1845 604 1846
rect 750 1850 756 1851
rect 750 1846 751 1850
rect 755 1846 756 1850
rect 750 1845 756 1846
rect 902 1850 908 1851
rect 902 1846 903 1850
rect 907 1846 908 1850
rect 902 1845 908 1846
rect 1054 1850 1060 1851
rect 1054 1846 1055 1850
rect 1059 1846 1060 1850
rect 1054 1845 1060 1846
rect 1206 1850 1212 1851
rect 1206 1846 1207 1850
rect 1211 1846 1212 1850
rect 1206 1845 1212 1846
rect 1350 1850 1356 1851
rect 1350 1846 1351 1850
rect 1355 1846 1356 1850
rect 1350 1845 1356 1846
rect 1486 1850 1492 1851
rect 1486 1846 1487 1850
rect 1491 1846 1492 1850
rect 1486 1845 1492 1846
rect 1630 1850 1636 1851
rect 1630 1846 1631 1850
rect 1635 1846 1636 1850
rect 1630 1845 1636 1846
rect 1750 1850 1756 1851
rect 1750 1846 1751 1850
rect 1755 1846 1756 1850
rect 1750 1845 1756 1846
rect 1870 1849 1876 1850
rect 1870 1845 1871 1849
rect 1875 1845 1876 1849
rect 1894 1848 1895 1852
rect 1899 1848 1900 1852
rect 1894 1847 1900 1848
rect 1990 1852 1996 1853
rect 1990 1848 1991 1852
rect 1995 1848 1996 1852
rect 1990 1847 1996 1848
rect 2118 1852 2124 1853
rect 2118 1848 2119 1852
rect 2123 1848 2124 1852
rect 2118 1847 2124 1848
rect 2246 1852 2252 1853
rect 2246 1848 2247 1852
rect 2251 1848 2252 1852
rect 2246 1847 2252 1848
rect 2382 1852 2388 1853
rect 2382 1848 2383 1852
rect 2387 1848 2388 1852
rect 2382 1847 2388 1848
rect 2518 1852 2524 1853
rect 2518 1848 2519 1852
rect 2523 1848 2524 1852
rect 2518 1847 2524 1848
rect 2654 1852 2660 1853
rect 2654 1848 2655 1852
rect 2659 1848 2660 1852
rect 2654 1847 2660 1848
rect 2806 1852 2812 1853
rect 2806 1848 2807 1852
rect 2811 1848 2812 1852
rect 2806 1847 2812 1848
rect 2974 1852 2980 1853
rect 2974 1848 2975 1852
rect 2979 1848 2980 1852
rect 2974 1847 2980 1848
rect 3150 1852 3156 1853
rect 3150 1848 3151 1852
rect 3155 1848 3156 1852
rect 3150 1847 3156 1848
rect 3334 1852 3340 1853
rect 3334 1848 3335 1852
rect 3339 1848 3340 1852
rect 3334 1847 3340 1848
rect 3502 1852 3508 1853
rect 3502 1848 3503 1852
rect 3507 1848 3508 1852
rect 3502 1847 3508 1848
rect 3590 1849 3596 1850
rect 1870 1844 1876 1845
rect 3590 1845 3591 1849
rect 3595 1845 3596 1849
rect 3590 1844 3596 1845
rect 1962 1843 1968 1844
rect 1962 1842 1963 1843
rect 1957 1840 1963 1842
rect 1962 1839 1963 1840
rect 1967 1839 1968 1843
rect 1962 1838 1968 1839
rect 1970 1843 1976 1844
rect 1970 1839 1971 1843
rect 1975 1842 1976 1843
rect 2190 1843 2196 1844
rect 2190 1842 2191 1843
rect 1975 1840 2009 1842
rect 2181 1840 2191 1842
rect 1975 1839 1976 1840
rect 1970 1838 1976 1839
rect 2190 1839 2191 1840
rect 2195 1839 2196 1843
rect 2342 1843 2348 1844
rect 2342 1842 2343 1843
rect 2309 1840 2343 1842
rect 2190 1838 2196 1839
rect 2342 1839 2343 1840
rect 2347 1839 2348 1843
rect 2342 1838 2348 1839
rect 2350 1843 2356 1844
rect 2350 1839 2351 1843
rect 2355 1842 2356 1843
rect 2594 1843 2600 1844
rect 2594 1842 2595 1843
rect 2355 1840 2401 1842
rect 2581 1840 2595 1842
rect 2355 1839 2356 1840
rect 2350 1838 2356 1839
rect 2594 1839 2595 1840
rect 2599 1839 2600 1843
rect 2730 1843 2736 1844
rect 2730 1842 2731 1843
rect 2717 1840 2731 1842
rect 2594 1838 2600 1839
rect 2730 1839 2731 1840
rect 2735 1839 2736 1843
rect 2898 1843 2904 1844
rect 2898 1842 2899 1843
rect 2869 1840 2899 1842
rect 2730 1838 2736 1839
rect 2898 1839 2899 1840
rect 2903 1839 2904 1843
rect 3050 1843 3056 1844
rect 3050 1842 3051 1843
rect 3037 1840 3051 1842
rect 2898 1838 2904 1839
rect 3050 1839 3051 1840
rect 3055 1839 3056 1843
rect 3250 1843 3256 1844
rect 3250 1842 3251 1843
rect 3213 1840 3251 1842
rect 3050 1838 3056 1839
rect 3250 1839 3251 1840
rect 3255 1839 3256 1843
rect 3250 1838 3256 1839
rect 3258 1843 3264 1844
rect 3258 1839 3259 1843
rect 3263 1842 3264 1843
rect 3263 1840 3353 1842
rect 3504 1840 3521 1842
rect 3263 1839 3264 1840
rect 3258 1838 3264 1839
rect 3502 1839 3508 1840
rect 3502 1835 3503 1839
rect 3507 1835 3508 1839
rect 3502 1834 3508 1835
rect 110 1832 116 1833
rect 110 1828 111 1832
rect 115 1828 116 1832
rect 110 1827 116 1828
rect 1830 1832 1836 1833
rect 1830 1828 1831 1832
rect 1835 1828 1836 1832
rect 1830 1827 1836 1828
rect 1870 1832 1876 1833
rect 1870 1828 1871 1832
rect 1875 1828 1876 1832
rect 1870 1827 1876 1828
rect 3590 1832 3596 1833
rect 3590 1828 3591 1832
rect 3595 1828 3596 1832
rect 3590 1827 3596 1828
rect 210 1823 216 1824
rect 210 1819 211 1823
rect 215 1819 216 1823
rect 210 1818 216 1819
rect 326 1823 332 1824
rect 326 1819 327 1823
rect 331 1819 332 1823
rect 326 1818 332 1819
rect 454 1823 460 1824
rect 454 1819 455 1823
rect 459 1819 460 1823
rect 679 1823 685 1824
rect 679 1822 680 1823
rect 653 1820 680 1822
rect 454 1818 460 1819
rect 679 1819 680 1820
rect 684 1819 685 1823
rect 838 1823 844 1824
rect 838 1822 839 1823
rect 805 1820 839 1822
rect 679 1818 685 1819
rect 838 1819 839 1820
rect 843 1819 844 1823
rect 838 1818 844 1819
rect 1078 1823 1084 1824
rect 1078 1819 1079 1823
rect 1083 1819 1084 1823
rect 1078 1818 1084 1819
rect 1127 1823 1133 1824
rect 1127 1819 1128 1823
rect 1132 1822 1133 1823
rect 1402 1823 1408 1824
rect 1132 1820 1217 1822
rect 1132 1819 1133 1820
rect 1127 1818 1133 1819
rect 1402 1819 1403 1823
rect 1407 1819 1408 1823
rect 1402 1818 1408 1819
rect 1538 1823 1544 1824
rect 1538 1819 1539 1823
rect 1543 1819 1544 1823
rect 1538 1818 1544 1819
rect 1682 1823 1688 1824
rect 1682 1819 1683 1823
rect 1687 1819 1688 1823
rect 2111 1823 2117 1824
rect 2111 1822 2112 1823
rect 1805 1820 2112 1822
rect 1682 1818 1688 1819
rect 2111 1819 2112 1820
rect 2116 1819 2117 1823
rect 2111 1818 2117 1819
rect 110 1815 116 1816
rect 110 1811 111 1815
rect 115 1811 116 1815
rect 1830 1815 1836 1816
rect 110 1810 116 1811
rect 150 1812 156 1813
rect 150 1808 151 1812
rect 155 1808 156 1812
rect 150 1807 156 1808
rect 294 1812 300 1813
rect 294 1808 295 1812
rect 299 1808 300 1812
rect 294 1807 300 1808
rect 438 1812 444 1813
rect 438 1808 439 1812
rect 443 1808 444 1812
rect 438 1807 444 1808
rect 590 1812 596 1813
rect 590 1808 591 1812
rect 595 1808 596 1812
rect 590 1807 596 1808
rect 742 1812 748 1813
rect 742 1808 743 1812
rect 747 1808 748 1812
rect 742 1807 748 1808
rect 894 1812 900 1813
rect 894 1808 895 1812
rect 899 1808 900 1812
rect 894 1807 900 1808
rect 1046 1812 1052 1813
rect 1046 1808 1047 1812
rect 1051 1808 1052 1812
rect 1046 1807 1052 1808
rect 1198 1812 1204 1813
rect 1198 1808 1199 1812
rect 1203 1808 1204 1812
rect 1198 1807 1204 1808
rect 1342 1812 1348 1813
rect 1342 1808 1343 1812
rect 1347 1808 1348 1812
rect 1342 1807 1348 1808
rect 1478 1812 1484 1813
rect 1478 1808 1479 1812
rect 1483 1808 1484 1812
rect 1478 1807 1484 1808
rect 1622 1812 1628 1813
rect 1622 1808 1623 1812
rect 1627 1808 1628 1812
rect 1622 1807 1628 1808
rect 1742 1812 1748 1813
rect 1742 1808 1743 1812
rect 1747 1808 1748 1812
rect 1830 1811 1831 1815
rect 1835 1811 1836 1815
rect 1830 1810 1836 1811
rect 1902 1814 1908 1815
rect 1902 1810 1903 1814
rect 1907 1810 1908 1814
rect 1902 1809 1908 1810
rect 1998 1814 2004 1815
rect 1998 1810 1999 1814
rect 2003 1810 2004 1814
rect 1998 1809 2004 1810
rect 2126 1814 2132 1815
rect 2126 1810 2127 1814
rect 2131 1810 2132 1814
rect 2126 1809 2132 1810
rect 2254 1814 2260 1815
rect 2254 1810 2255 1814
rect 2259 1810 2260 1814
rect 2254 1809 2260 1810
rect 2390 1814 2396 1815
rect 2390 1810 2391 1814
rect 2395 1810 2396 1814
rect 2390 1809 2396 1810
rect 2526 1814 2532 1815
rect 2526 1810 2527 1814
rect 2531 1810 2532 1814
rect 2526 1809 2532 1810
rect 2662 1814 2668 1815
rect 2662 1810 2663 1814
rect 2667 1810 2668 1814
rect 2662 1809 2668 1810
rect 2814 1814 2820 1815
rect 2814 1810 2815 1814
rect 2819 1810 2820 1814
rect 2814 1809 2820 1810
rect 2982 1814 2988 1815
rect 2982 1810 2983 1814
rect 2987 1810 2988 1814
rect 2982 1809 2988 1810
rect 3158 1814 3164 1815
rect 3158 1810 3159 1814
rect 3163 1810 3164 1814
rect 3158 1809 3164 1810
rect 3342 1814 3348 1815
rect 3342 1810 3343 1814
rect 3347 1810 3348 1814
rect 3342 1809 3348 1810
rect 3510 1814 3516 1815
rect 3510 1810 3511 1814
rect 3515 1810 3516 1814
rect 3510 1809 3516 1810
rect 1742 1807 1748 1808
rect 1895 1803 1901 1804
rect 1895 1799 1896 1803
rect 1900 1802 1901 1803
rect 1910 1803 1916 1804
rect 1910 1802 1911 1803
rect 1900 1800 1911 1802
rect 1900 1799 1901 1800
rect 1895 1798 1901 1799
rect 1910 1799 1911 1800
rect 1915 1799 1916 1803
rect 1910 1798 1916 1799
rect 1962 1803 1968 1804
rect 1962 1799 1963 1803
rect 1967 1802 1968 1803
rect 1991 1803 1997 1804
rect 1991 1802 1992 1803
rect 1967 1800 1992 1802
rect 1967 1799 1968 1800
rect 1962 1798 1968 1799
rect 1991 1799 1992 1800
rect 1996 1799 1997 1803
rect 1991 1798 1997 1799
rect 2111 1803 2117 1804
rect 2111 1799 2112 1803
rect 2116 1802 2117 1803
rect 2119 1803 2125 1804
rect 2119 1802 2120 1803
rect 2116 1800 2120 1802
rect 2116 1799 2117 1800
rect 2111 1798 2117 1799
rect 2119 1799 2120 1800
rect 2124 1799 2125 1803
rect 2119 1798 2125 1799
rect 2190 1803 2196 1804
rect 2190 1799 2191 1803
rect 2195 1802 2196 1803
rect 2247 1803 2253 1804
rect 2247 1802 2248 1803
rect 2195 1800 2248 1802
rect 2195 1799 2196 1800
rect 2190 1798 2196 1799
rect 2247 1799 2248 1800
rect 2252 1799 2253 1803
rect 2247 1798 2253 1799
rect 2342 1803 2348 1804
rect 2342 1799 2343 1803
rect 2347 1802 2348 1803
rect 2383 1803 2389 1804
rect 2383 1802 2384 1803
rect 2347 1800 2384 1802
rect 2347 1799 2348 1800
rect 2342 1798 2348 1799
rect 2383 1799 2384 1800
rect 2388 1799 2389 1803
rect 2383 1798 2389 1799
rect 2519 1803 2525 1804
rect 2519 1799 2520 1803
rect 2524 1802 2525 1803
rect 2534 1803 2540 1804
rect 2534 1802 2535 1803
rect 2524 1800 2535 1802
rect 2524 1799 2525 1800
rect 2519 1798 2525 1799
rect 2534 1799 2535 1800
rect 2539 1799 2540 1803
rect 2534 1798 2540 1799
rect 2594 1803 2600 1804
rect 2594 1799 2595 1803
rect 2599 1802 2600 1803
rect 2655 1803 2661 1804
rect 2655 1802 2656 1803
rect 2599 1800 2656 1802
rect 2599 1799 2600 1800
rect 2594 1798 2600 1799
rect 2655 1799 2656 1800
rect 2660 1799 2661 1803
rect 2655 1798 2661 1799
rect 2730 1803 2736 1804
rect 2730 1799 2731 1803
rect 2735 1802 2736 1803
rect 2807 1803 2813 1804
rect 2807 1802 2808 1803
rect 2735 1800 2808 1802
rect 2735 1799 2736 1800
rect 2730 1798 2736 1799
rect 2807 1799 2808 1800
rect 2812 1799 2813 1803
rect 2807 1798 2813 1799
rect 2898 1803 2904 1804
rect 2898 1799 2899 1803
rect 2903 1802 2904 1803
rect 2975 1803 2981 1804
rect 2975 1802 2976 1803
rect 2903 1800 2976 1802
rect 2903 1799 2904 1800
rect 2898 1798 2904 1799
rect 2975 1799 2976 1800
rect 2980 1799 2981 1803
rect 2975 1798 2981 1799
rect 3050 1803 3056 1804
rect 3050 1799 3051 1803
rect 3055 1802 3056 1803
rect 3151 1803 3157 1804
rect 3151 1802 3152 1803
rect 3055 1800 3152 1802
rect 3055 1799 3056 1800
rect 3050 1798 3056 1799
rect 3151 1799 3152 1800
rect 3156 1799 3157 1803
rect 3151 1798 3157 1799
rect 3250 1803 3256 1804
rect 3250 1799 3251 1803
rect 3255 1802 3256 1803
rect 3335 1803 3341 1804
rect 3335 1802 3336 1803
rect 3255 1800 3336 1802
rect 3255 1799 3256 1800
rect 3250 1798 3256 1799
rect 3335 1799 3336 1800
rect 3340 1799 3341 1803
rect 3335 1798 3341 1799
rect 3503 1803 3509 1804
rect 3503 1799 3504 1803
rect 3508 1802 3509 1803
rect 3526 1803 3532 1804
rect 3526 1802 3527 1803
rect 3508 1800 3527 1802
rect 3508 1799 3509 1800
rect 3503 1798 3509 1799
rect 3526 1799 3527 1800
rect 3531 1799 3532 1803
rect 3526 1798 3532 1799
rect 766 1795 772 1796
rect 766 1791 767 1795
rect 771 1794 772 1795
rect 911 1795 917 1796
rect 911 1794 912 1795
rect 771 1792 912 1794
rect 771 1791 772 1792
rect 766 1790 772 1791
rect 911 1791 912 1792
rect 916 1791 917 1795
rect 911 1790 917 1791
rect 1970 1787 1976 1788
rect 1970 1786 1971 1787
rect 1944 1784 1971 1786
rect 1895 1779 1901 1780
rect 1895 1775 1896 1779
rect 1900 1778 1901 1779
rect 1944 1778 1946 1784
rect 1970 1783 1971 1784
rect 1975 1783 1976 1787
rect 1970 1782 1976 1783
rect 1900 1776 1946 1778
rect 1954 1779 1960 1780
rect 1900 1775 1901 1776
rect 1895 1774 1901 1775
rect 1954 1775 1955 1779
rect 1959 1778 1960 1779
rect 2023 1779 2029 1780
rect 2023 1778 2024 1779
rect 1959 1776 2024 1778
rect 1959 1775 1960 1776
rect 1954 1774 1960 1775
rect 2023 1775 2024 1776
rect 2028 1775 2029 1779
rect 2023 1774 2029 1775
rect 2082 1779 2088 1780
rect 2082 1775 2083 1779
rect 2087 1778 2088 1779
rect 2183 1779 2189 1780
rect 2183 1778 2184 1779
rect 2087 1776 2184 1778
rect 2087 1775 2088 1776
rect 2082 1774 2088 1775
rect 2183 1775 2184 1776
rect 2188 1775 2189 1779
rect 2183 1774 2189 1775
rect 2242 1779 2248 1780
rect 2242 1775 2243 1779
rect 2247 1778 2248 1779
rect 2351 1779 2357 1780
rect 2351 1778 2352 1779
rect 2247 1776 2352 1778
rect 2247 1775 2248 1776
rect 2242 1774 2248 1775
rect 2351 1775 2352 1776
rect 2356 1775 2357 1779
rect 2351 1774 2357 1775
rect 2410 1779 2416 1780
rect 2410 1775 2411 1779
rect 2415 1778 2416 1779
rect 2519 1779 2525 1780
rect 2519 1778 2520 1779
rect 2415 1776 2520 1778
rect 2415 1775 2416 1776
rect 2410 1774 2416 1775
rect 2519 1775 2520 1776
rect 2524 1775 2525 1779
rect 2519 1774 2525 1775
rect 2679 1779 2685 1780
rect 2679 1775 2680 1779
rect 2684 1778 2685 1779
rect 2694 1779 2700 1780
rect 2694 1778 2695 1779
rect 2684 1776 2695 1778
rect 2684 1775 2685 1776
rect 2679 1774 2685 1775
rect 2694 1775 2695 1776
rect 2699 1775 2700 1779
rect 2694 1774 2700 1775
rect 2738 1779 2744 1780
rect 2738 1775 2739 1779
rect 2743 1778 2744 1779
rect 2831 1779 2837 1780
rect 2831 1778 2832 1779
rect 2743 1776 2832 1778
rect 2743 1775 2744 1776
rect 2738 1774 2744 1775
rect 2831 1775 2832 1776
rect 2836 1775 2837 1779
rect 2831 1774 2837 1775
rect 2890 1779 2896 1780
rect 2890 1775 2891 1779
rect 2895 1778 2896 1779
rect 2975 1779 2981 1780
rect 2975 1778 2976 1779
rect 2895 1776 2976 1778
rect 2895 1775 2896 1776
rect 2890 1774 2896 1775
rect 2975 1775 2976 1776
rect 2980 1775 2981 1779
rect 2975 1774 2981 1775
rect 3034 1779 3040 1780
rect 3034 1775 3035 1779
rect 3039 1778 3040 1779
rect 3111 1779 3117 1780
rect 3111 1778 3112 1779
rect 3039 1776 3112 1778
rect 3039 1775 3040 1776
rect 3034 1774 3040 1775
rect 3111 1775 3112 1776
rect 3116 1775 3117 1779
rect 3111 1774 3117 1775
rect 3170 1779 3176 1780
rect 3170 1775 3171 1779
rect 3175 1778 3176 1779
rect 3247 1779 3253 1780
rect 3247 1778 3248 1779
rect 3175 1776 3248 1778
rect 3175 1775 3176 1776
rect 3170 1774 3176 1775
rect 3247 1775 3248 1776
rect 3252 1775 3253 1779
rect 3247 1774 3253 1775
rect 3306 1779 3312 1780
rect 3306 1775 3307 1779
rect 3311 1778 3312 1779
rect 3383 1779 3389 1780
rect 3383 1778 3384 1779
rect 3311 1776 3384 1778
rect 3311 1775 3312 1776
rect 3306 1774 3312 1775
rect 3383 1775 3384 1776
rect 3388 1775 3389 1779
rect 3383 1774 3389 1775
rect 3502 1779 3509 1780
rect 3502 1775 3503 1779
rect 3508 1775 3509 1779
rect 3502 1774 3509 1775
rect 1902 1770 1908 1771
rect 1902 1766 1903 1770
rect 1907 1766 1908 1770
rect 1902 1765 1908 1766
rect 2030 1770 2036 1771
rect 2030 1766 2031 1770
rect 2035 1766 2036 1770
rect 2030 1765 2036 1766
rect 2190 1770 2196 1771
rect 2190 1766 2191 1770
rect 2195 1766 2196 1770
rect 2190 1765 2196 1766
rect 2358 1770 2364 1771
rect 2358 1766 2359 1770
rect 2363 1766 2364 1770
rect 2358 1765 2364 1766
rect 2526 1770 2532 1771
rect 2526 1766 2527 1770
rect 2531 1766 2532 1770
rect 2526 1765 2532 1766
rect 2686 1770 2692 1771
rect 2686 1766 2687 1770
rect 2691 1766 2692 1770
rect 2686 1765 2692 1766
rect 2838 1770 2844 1771
rect 2838 1766 2839 1770
rect 2843 1766 2844 1770
rect 2838 1765 2844 1766
rect 2982 1770 2988 1771
rect 2982 1766 2983 1770
rect 2987 1766 2988 1770
rect 2982 1765 2988 1766
rect 3118 1770 3124 1771
rect 3118 1766 3119 1770
rect 3123 1766 3124 1770
rect 3118 1765 3124 1766
rect 3254 1770 3260 1771
rect 3254 1766 3255 1770
rect 3259 1766 3260 1770
rect 3254 1765 3260 1766
rect 3390 1770 3396 1771
rect 3390 1766 3391 1770
rect 3395 1766 3396 1770
rect 3390 1765 3396 1766
rect 3510 1770 3516 1771
rect 3510 1766 3511 1770
rect 3515 1766 3516 1770
rect 3510 1765 3516 1766
rect 246 1764 252 1765
rect 110 1761 116 1762
rect 110 1757 111 1761
rect 115 1757 116 1761
rect 246 1760 247 1764
rect 251 1760 252 1764
rect 246 1759 252 1760
rect 422 1764 428 1765
rect 422 1760 423 1764
rect 427 1760 428 1764
rect 422 1759 428 1760
rect 590 1764 596 1765
rect 590 1760 591 1764
rect 595 1760 596 1764
rect 590 1759 596 1760
rect 750 1764 756 1765
rect 750 1760 751 1764
rect 755 1760 756 1764
rect 750 1759 756 1760
rect 894 1764 900 1765
rect 894 1760 895 1764
rect 899 1760 900 1764
rect 894 1759 900 1760
rect 1022 1764 1028 1765
rect 1022 1760 1023 1764
rect 1027 1760 1028 1764
rect 1022 1759 1028 1760
rect 1142 1764 1148 1765
rect 1142 1760 1143 1764
rect 1147 1760 1148 1764
rect 1142 1759 1148 1760
rect 1262 1764 1268 1765
rect 1262 1760 1263 1764
rect 1267 1760 1268 1764
rect 1262 1759 1268 1760
rect 1390 1764 1396 1765
rect 1390 1760 1391 1764
rect 1395 1760 1396 1764
rect 1390 1759 1396 1760
rect 1830 1761 1836 1762
rect 110 1756 116 1757
rect 1830 1757 1831 1761
rect 1835 1757 1836 1761
rect 1830 1756 1836 1757
rect 342 1755 348 1756
rect 342 1754 343 1755
rect 309 1752 343 1754
rect 342 1751 343 1752
rect 347 1751 348 1755
rect 582 1755 588 1756
rect 342 1750 348 1751
rect 430 1751 436 1752
rect 430 1747 431 1751
rect 435 1750 436 1751
rect 440 1750 442 1753
rect 582 1751 583 1755
rect 587 1754 588 1755
rect 678 1755 684 1756
rect 587 1752 609 1754
rect 587 1751 588 1752
rect 582 1750 588 1751
rect 678 1751 679 1755
rect 683 1754 684 1755
rect 966 1755 972 1756
rect 966 1754 967 1755
rect 683 1752 769 1754
rect 957 1752 967 1754
rect 683 1751 684 1752
rect 678 1750 684 1751
rect 966 1751 967 1752
rect 971 1751 972 1755
rect 1090 1755 1096 1756
rect 1090 1754 1091 1755
rect 1085 1752 1091 1754
rect 966 1750 972 1751
rect 1090 1751 1091 1752
rect 1095 1751 1096 1755
rect 1210 1755 1216 1756
rect 1210 1754 1211 1755
rect 1205 1752 1211 1754
rect 1090 1750 1096 1751
rect 1210 1751 1211 1752
rect 1215 1751 1216 1755
rect 1334 1755 1340 1756
rect 1334 1754 1335 1755
rect 1325 1752 1335 1754
rect 1210 1750 1216 1751
rect 1334 1751 1335 1752
rect 1339 1751 1340 1755
rect 1334 1750 1340 1751
rect 1342 1755 1348 1756
rect 1342 1751 1343 1755
rect 1347 1754 1348 1755
rect 1347 1752 1409 1754
rect 1870 1752 1876 1753
rect 1347 1751 1348 1752
rect 1342 1750 1348 1751
rect 435 1748 442 1750
rect 1870 1748 1871 1752
rect 1875 1748 1876 1752
rect 435 1747 436 1748
rect 1870 1747 1876 1748
rect 3590 1752 3596 1753
rect 3590 1748 3591 1752
rect 3595 1748 3596 1752
rect 3590 1747 3596 1748
rect 430 1746 436 1747
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 110 1739 116 1740
rect 1830 1744 1836 1745
rect 1830 1740 1831 1744
rect 1835 1740 1836 1744
rect 1830 1739 1836 1740
rect 1954 1743 1960 1744
rect 1954 1739 1955 1743
rect 1959 1739 1960 1743
rect 1954 1738 1960 1739
rect 2082 1743 2088 1744
rect 2082 1739 2083 1743
rect 2087 1739 2088 1743
rect 2082 1738 2088 1739
rect 2242 1743 2248 1744
rect 2242 1739 2243 1743
rect 2247 1739 2248 1743
rect 2242 1738 2248 1739
rect 2410 1743 2416 1744
rect 2410 1739 2411 1743
rect 2415 1739 2416 1743
rect 2410 1738 2416 1739
rect 2738 1743 2744 1744
rect 2738 1739 2739 1743
rect 2743 1739 2744 1743
rect 2738 1738 2744 1739
rect 2890 1743 2896 1744
rect 2890 1739 2891 1743
rect 2895 1739 2896 1743
rect 2890 1738 2896 1739
rect 3034 1743 3040 1744
rect 3034 1739 3035 1743
rect 3039 1739 3040 1743
rect 3034 1738 3040 1739
rect 3170 1743 3176 1744
rect 3170 1739 3171 1743
rect 3175 1739 3176 1743
rect 3170 1738 3176 1739
rect 3306 1743 3312 1744
rect 3306 1739 3307 1743
rect 3311 1739 3312 1743
rect 3306 1738 3312 1739
rect 1870 1735 1876 1736
rect 1870 1731 1871 1735
rect 1875 1731 1876 1735
rect 3590 1735 3596 1736
rect 1870 1730 1876 1731
rect 1894 1732 1900 1733
rect 1894 1728 1895 1732
rect 1899 1728 1900 1732
rect 1894 1727 1900 1728
rect 2022 1732 2028 1733
rect 2022 1728 2023 1732
rect 2027 1728 2028 1732
rect 2022 1727 2028 1728
rect 2182 1732 2188 1733
rect 2182 1728 2183 1732
rect 2187 1728 2188 1732
rect 2182 1727 2188 1728
rect 2350 1732 2356 1733
rect 2350 1728 2351 1732
rect 2355 1728 2356 1732
rect 2350 1727 2356 1728
rect 2518 1732 2524 1733
rect 2518 1728 2519 1732
rect 2523 1728 2524 1732
rect 2518 1727 2524 1728
rect 2678 1732 2684 1733
rect 2678 1728 2679 1732
rect 2683 1728 2684 1732
rect 2678 1727 2684 1728
rect 2830 1732 2836 1733
rect 2830 1728 2831 1732
rect 2835 1728 2836 1732
rect 2830 1727 2836 1728
rect 2974 1732 2980 1733
rect 2974 1728 2975 1732
rect 2979 1728 2980 1732
rect 2974 1727 2980 1728
rect 3110 1732 3116 1733
rect 3110 1728 3111 1732
rect 3115 1728 3116 1732
rect 3110 1727 3116 1728
rect 3246 1732 3252 1733
rect 3246 1728 3247 1732
rect 3251 1728 3252 1732
rect 3246 1727 3252 1728
rect 3382 1732 3388 1733
rect 3382 1728 3383 1732
rect 3387 1728 3388 1732
rect 3382 1727 3388 1728
rect 3502 1732 3508 1733
rect 3502 1728 3503 1732
rect 3507 1728 3508 1732
rect 3590 1731 3591 1735
rect 3595 1731 3596 1735
rect 3590 1730 3596 1731
rect 3502 1727 3508 1728
rect 254 1726 260 1727
rect 254 1722 255 1726
rect 259 1722 260 1726
rect 254 1721 260 1722
rect 430 1726 436 1727
rect 430 1722 431 1726
rect 435 1722 436 1726
rect 430 1721 436 1722
rect 598 1726 604 1727
rect 598 1722 599 1726
rect 603 1722 604 1726
rect 598 1721 604 1722
rect 758 1726 764 1727
rect 758 1722 759 1726
rect 763 1722 764 1726
rect 758 1721 764 1722
rect 902 1726 908 1727
rect 902 1722 903 1726
rect 907 1722 908 1726
rect 902 1721 908 1722
rect 1030 1726 1036 1727
rect 1030 1722 1031 1726
rect 1035 1722 1036 1726
rect 1030 1721 1036 1722
rect 1150 1726 1156 1727
rect 1150 1722 1151 1726
rect 1155 1722 1156 1726
rect 1150 1721 1156 1722
rect 1270 1726 1276 1727
rect 1270 1722 1271 1726
rect 1275 1722 1276 1726
rect 1270 1721 1276 1722
rect 1398 1726 1404 1727
rect 1398 1722 1399 1726
rect 1403 1722 1404 1726
rect 1398 1721 1404 1722
rect 247 1715 253 1716
rect 247 1711 248 1715
rect 252 1714 253 1715
rect 342 1715 348 1716
rect 252 1712 338 1714
rect 252 1711 253 1712
rect 247 1710 253 1711
rect 336 1706 338 1712
rect 342 1711 343 1715
rect 347 1714 348 1715
rect 423 1715 429 1716
rect 423 1714 424 1715
rect 347 1712 424 1714
rect 347 1711 348 1712
rect 342 1710 348 1711
rect 423 1711 424 1712
rect 428 1711 429 1715
rect 423 1710 429 1711
rect 591 1715 597 1716
rect 591 1711 592 1715
rect 596 1714 597 1715
rect 678 1715 684 1716
rect 678 1714 679 1715
rect 596 1712 679 1714
rect 596 1711 597 1712
rect 591 1710 597 1711
rect 678 1711 679 1712
rect 683 1711 684 1715
rect 678 1710 684 1711
rect 751 1715 757 1716
rect 751 1711 752 1715
rect 756 1714 757 1715
rect 766 1715 772 1716
rect 766 1714 767 1715
rect 756 1712 767 1714
rect 756 1711 757 1712
rect 751 1710 757 1711
rect 766 1711 767 1712
rect 771 1711 772 1715
rect 766 1710 772 1711
rect 895 1715 901 1716
rect 895 1711 896 1715
rect 900 1714 901 1715
rect 910 1715 916 1716
rect 910 1714 911 1715
rect 900 1712 911 1714
rect 900 1711 901 1712
rect 895 1710 901 1711
rect 910 1711 911 1712
rect 915 1711 916 1715
rect 910 1710 916 1711
rect 966 1715 972 1716
rect 966 1711 967 1715
rect 971 1714 972 1715
rect 1023 1715 1029 1716
rect 1023 1714 1024 1715
rect 971 1712 1024 1714
rect 971 1711 972 1712
rect 966 1710 972 1711
rect 1023 1711 1024 1712
rect 1028 1711 1029 1715
rect 1023 1710 1029 1711
rect 1090 1715 1096 1716
rect 1090 1711 1091 1715
rect 1095 1714 1096 1715
rect 1143 1715 1149 1716
rect 1143 1714 1144 1715
rect 1095 1712 1144 1714
rect 1095 1711 1096 1712
rect 1090 1710 1096 1711
rect 1143 1711 1144 1712
rect 1148 1711 1149 1715
rect 1143 1710 1149 1711
rect 1234 1715 1240 1716
rect 1234 1711 1235 1715
rect 1239 1714 1240 1715
rect 1263 1715 1269 1716
rect 1263 1714 1264 1715
rect 1239 1712 1264 1714
rect 1239 1711 1240 1712
rect 1234 1710 1240 1711
rect 1263 1711 1264 1712
rect 1268 1711 1269 1715
rect 1263 1710 1269 1711
rect 1334 1715 1340 1716
rect 1334 1711 1335 1715
rect 1339 1714 1340 1715
rect 1391 1715 1397 1716
rect 1391 1714 1392 1715
rect 1339 1712 1392 1714
rect 1339 1711 1340 1712
rect 1334 1710 1340 1711
rect 1391 1711 1392 1712
rect 1396 1711 1397 1715
rect 1391 1710 1397 1711
rect 2418 1715 2424 1716
rect 2418 1711 2419 1715
rect 2423 1714 2424 1715
rect 2535 1715 2541 1716
rect 2535 1714 2536 1715
rect 2423 1712 2536 1714
rect 2423 1711 2424 1712
rect 2418 1710 2424 1711
rect 2535 1711 2536 1712
rect 2540 1711 2541 1715
rect 2535 1710 2541 1711
rect 3398 1715 3405 1716
rect 3398 1711 3399 1715
rect 3404 1711 3405 1715
rect 3398 1710 3405 1711
rect 3518 1715 3525 1716
rect 3518 1711 3519 1715
rect 3524 1711 3525 1715
rect 3518 1710 3525 1711
rect 454 1707 460 1708
rect 454 1706 455 1707
rect 336 1704 455 1706
rect 454 1703 455 1704
rect 459 1703 460 1707
rect 454 1702 460 1703
rect 174 1699 180 1700
rect 174 1695 175 1699
rect 179 1698 180 1699
rect 183 1699 189 1700
rect 183 1698 184 1699
rect 179 1696 184 1698
rect 179 1695 180 1696
rect 174 1694 180 1695
rect 183 1695 184 1696
rect 188 1695 189 1699
rect 183 1694 189 1695
rect 242 1699 248 1700
rect 242 1695 243 1699
rect 247 1698 248 1699
rect 303 1699 309 1700
rect 303 1698 304 1699
rect 247 1696 304 1698
rect 247 1695 248 1696
rect 242 1694 248 1695
rect 303 1695 304 1696
rect 308 1695 309 1699
rect 303 1694 309 1695
rect 362 1699 368 1700
rect 362 1695 363 1699
rect 367 1698 368 1699
rect 439 1699 445 1700
rect 439 1698 440 1699
rect 367 1696 440 1698
rect 367 1695 368 1696
rect 362 1694 368 1695
rect 439 1695 440 1696
rect 444 1695 445 1699
rect 439 1694 445 1695
rect 582 1699 589 1700
rect 582 1695 583 1699
rect 588 1695 589 1699
rect 582 1694 589 1695
rect 642 1699 648 1700
rect 642 1695 643 1699
rect 647 1698 648 1699
rect 735 1699 741 1700
rect 735 1698 736 1699
rect 647 1696 736 1698
rect 647 1695 648 1696
rect 642 1694 648 1695
rect 735 1695 736 1696
rect 740 1695 741 1699
rect 735 1694 741 1695
rect 794 1699 800 1700
rect 794 1695 795 1699
rect 799 1698 800 1699
rect 887 1699 893 1700
rect 887 1698 888 1699
rect 799 1696 888 1698
rect 799 1695 800 1696
rect 794 1694 800 1695
rect 887 1695 888 1696
rect 892 1695 893 1699
rect 887 1694 893 1695
rect 946 1699 952 1700
rect 946 1695 947 1699
rect 951 1698 952 1699
rect 1031 1699 1037 1700
rect 1031 1698 1032 1699
rect 951 1696 1032 1698
rect 951 1695 952 1696
rect 946 1694 952 1695
rect 1031 1695 1032 1696
rect 1036 1695 1037 1699
rect 1031 1694 1037 1695
rect 1175 1699 1181 1700
rect 1175 1695 1176 1699
rect 1180 1698 1181 1699
rect 1242 1699 1248 1700
rect 1242 1698 1243 1699
rect 1180 1696 1243 1698
rect 1180 1695 1181 1696
rect 1175 1694 1181 1695
rect 1242 1695 1243 1696
rect 1247 1695 1248 1699
rect 1242 1694 1248 1695
rect 1311 1699 1317 1700
rect 1311 1695 1312 1699
rect 1316 1698 1317 1699
rect 1378 1699 1384 1700
rect 1378 1698 1379 1699
rect 1316 1696 1379 1698
rect 1316 1695 1317 1696
rect 1311 1694 1317 1695
rect 1378 1695 1379 1696
rect 1383 1695 1384 1699
rect 1378 1694 1384 1695
rect 1439 1699 1445 1700
rect 1439 1695 1440 1699
rect 1444 1698 1445 1699
rect 1519 1699 1525 1700
rect 1519 1698 1520 1699
rect 1444 1696 1520 1698
rect 1444 1695 1445 1696
rect 1439 1694 1445 1695
rect 1519 1695 1520 1696
rect 1524 1695 1525 1699
rect 1519 1694 1525 1695
rect 1567 1699 1573 1700
rect 1567 1695 1568 1699
rect 1572 1698 1573 1699
rect 1634 1699 1640 1700
rect 1634 1698 1635 1699
rect 1572 1696 1635 1698
rect 1572 1695 1573 1696
rect 1567 1694 1573 1695
rect 1634 1695 1635 1696
rect 1639 1695 1640 1699
rect 1634 1694 1640 1695
rect 1703 1699 1709 1700
rect 1703 1695 1704 1699
rect 1708 1698 1709 1699
rect 1726 1699 1732 1700
rect 1726 1698 1727 1699
rect 1708 1696 1727 1698
rect 1708 1695 1709 1696
rect 1703 1694 1709 1695
rect 1726 1695 1727 1696
rect 1731 1695 1732 1699
rect 1726 1694 1732 1695
rect 190 1690 196 1691
rect 190 1686 191 1690
rect 195 1686 196 1690
rect 190 1685 196 1686
rect 310 1690 316 1691
rect 310 1686 311 1690
rect 315 1686 316 1690
rect 310 1685 316 1686
rect 446 1690 452 1691
rect 446 1686 447 1690
rect 451 1686 452 1690
rect 446 1685 452 1686
rect 590 1690 596 1691
rect 590 1686 591 1690
rect 595 1686 596 1690
rect 590 1685 596 1686
rect 742 1690 748 1691
rect 742 1686 743 1690
rect 747 1686 748 1690
rect 742 1685 748 1686
rect 894 1690 900 1691
rect 894 1686 895 1690
rect 899 1686 900 1690
rect 894 1685 900 1686
rect 1038 1690 1044 1691
rect 1038 1686 1039 1690
rect 1043 1686 1044 1690
rect 1038 1685 1044 1686
rect 1182 1690 1188 1691
rect 1182 1686 1183 1690
rect 1187 1686 1188 1690
rect 1182 1685 1188 1686
rect 1318 1690 1324 1691
rect 1318 1686 1319 1690
rect 1323 1686 1324 1690
rect 1318 1685 1324 1686
rect 1446 1690 1452 1691
rect 1446 1686 1447 1690
rect 1451 1686 1452 1690
rect 1446 1685 1452 1686
rect 1574 1690 1580 1691
rect 1574 1686 1575 1690
rect 1579 1686 1580 1690
rect 1574 1685 1580 1686
rect 1710 1690 1716 1691
rect 1710 1686 1711 1690
rect 1715 1686 1716 1690
rect 1710 1685 1716 1686
rect 1894 1684 1900 1685
rect 1870 1681 1876 1682
rect 1870 1677 1871 1681
rect 1875 1677 1876 1681
rect 1894 1680 1895 1684
rect 1899 1680 1900 1684
rect 1894 1679 1900 1680
rect 1990 1684 1996 1685
rect 1990 1680 1991 1684
rect 1995 1680 1996 1684
rect 1990 1679 1996 1680
rect 2134 1684 2140 1685
rect 2134 1680 2135 1684
rect 2139 1680 2140 1684
rect 2134 1679 2140 1680
rect 2294 1684 2300 1685
rect 2294 1680 2295 1684
rect 2299 1680 2300 1684
rect 2294 1679 2300 1680
rect 2470 1684 2476 1685
rect 2470 1680 2471 1684
rect 2475 1680 2476 1684
rect 2470 1679 2476 1680
rect 2646 1684 2652 1685
rect 2646 1680 2647 1684
rect 2651 1680 2652 1684
rect 2646 1679 2652 1680
rect 2814 1684 2820 1685
rect 2814 1680 2815 1684
rect 2819 1680 2820 1684
rect 2814 1679 2820 1680
rect 2966 1684 2972 1685
rect 2966 1680 2967 1684
rect 2971 1680 2972 1684
rect 2966 1679 2972 1680
rect 3110 1684 3116 1685
rect 3110 1680 3111 1684
rect 3115 1680 3116 1684
rect 3110 1679 3116 1680
rect 3246 1684 3252 1685
rect 3246 1680 3247 1684
rect 3251 1680 3252 1684
rect 3246 1679 3252 1680
rect 3382 1684 3388 1685
rect 3382 1680 3383 1684
rect 3387 1680 3388 1684
rect 3382 1679 3388 1680
rect 3502 1684 3508 1685
rect 3502 1680 3503 1684
rect 3507 1680 3508 1684
rect 3502 1679 3508 1680
rect 3590 1681 3596 1682
rect 1870 1676 1876 1677
rect 3590 1677 3591 1681
rect 3595 1677 3596 1681
rect 3590 1676 3596 1677
rect 1962 1675 1968 1676
rect 1962 1674 1963 1675
rect 110 1672 116 1673
rect 110 1668 111 1672
rect 115 1668 116 1672
rect 110 1667 116 1668
rect 1830 1672 1836 1673
rect 1957 1672 1963 1674
rect 1830 1668 1831 1672
rect 1835 1668 1836 1672
rect 1962 1671 1963 1672
rect 1967 1671 1968 1675
rect 2070 1675 2076 1676
rect 2070 1674 2071 1675
rect 2053 1672 2071 1674
rect 1962 1670 1968 1671
rect 2070 1671 2071 1672
rect 2075 1671 2076 1675
rect 2222 1675 2228 1676
rect 2222 1674 2223 1675
rect 2197 1672 2223 1674
rect 2070 1670 2076 1671
rect 2222 1671 2223 1672
rect 2227 1671 2228 1675
rect 2390 1675 2396 1676
rect 2390 1674 2391 1675
rect 2357 1672 2391 1674
rect 2222 1670 2228 1671
rect 2390 1671 2391 1672
rect 2395 1671 2396 1675
rect 2566 1675 2572 1676
rect 2566 1674 2567 1675
rect 2533 1672 2567 1674
rect 2390 1670 2396 1671
rect 2566 1671 2567 1672
rect 2571 1671 2572 1675
rect 2566 1670 2572 1671
rect 2574 1675 2580 1676
rect 2574 1671 2575 1675
rect 2579 1674 2580 1675
rect 2890 1675 2896 1676
rect 2890 1674 2891 1675
rect 2579 1672 2665 1674
rect 2877 1672 2891 1674
rect 2579 1671 2580 1672
rect 2574 1670 2580 1671
rect 2890 1671 2891 1672
rect 2895 1671 2896 1675
rect 3046 1675 3052 1676
rect 3046 1674 3047 1675
rect 3029 1672 3047 1674
rect 2890 1670 2896 1671
rect 3046 1671 3047 1672
rect 3051 1671 3052 1675
rect 3178 1675 3184 1676
rect 3178 1674 3179 1675
rect 3173 1672 3179 1674
rect 3046 1670 3052 1671
rect 3178 1671 3179 1672
rect 3183 1671 3184 1675
rect 3178 1670 3184 1671
rect 3186 1675 3192 1676
rect 3186 1671 3187 1675
rect 3191 1674 3192 1675
rect 3322 1675 3328 1676
rect 3191 1672 3265 1674
rect 3191 1671 3192 1672
rect 3186 1670 3192 1671
rect 3322 1671 3323 1675
rect 3327 1674 3328 1675
rect 3487 1675 3493 1676
rect 3327 1672 3401 1674
rect 3327 1671 3328 1672
rect 3322 1670 3328 1671
rect 3487 1671 3488 1675
rect 3492 1674 3493 1675
rect 3492 1672 3521 1674
rect 3492 1671 3493 1672
rect 3487 1670 3493 1671
rect 1830 1667 1836 1668
rect 1870 1664 1876 1665
rect 242 1663 248 1664
rect 242 1659 243 1663
rect 247 1659 248 1663
rect 242 1658 248 1659
rect 362 1663 368 1664
rect 362 1659 363 1663
rect 367 1659 368 1663
rect 362 1658 368 1659
rect 454 1663 460 1664
rect 454 1659 455 1663
rect 459 1659 460 1663
rect 454 1658 460 1659
rect 642 1663 648 1664
rect 642 1659 643 1663
rect 647 1659 648 1663
rect 642 1658 648 1659
rect 794 1663 800 1664
rect 794 1659 795 1663
rect 799 1659 800 1663
rect 794 1658 800 1659
rect 946 1663 952 1664
rect 946 1659 947 1663
rect 951 1659 952 1663
rect 946 1658 952 1659
rect 1234 1663 1240 1664
rect 1234 1659 1235 1663
rect 1239 1659 1240 1663
rect 1234 1658 1240 1659
rect 1242 1663 1248 1664
rect 1242 1659 1243 1663
rect 1247 1662 1248 1663
rect 1378 1663 1384 1664
rect 1247 1660 1329 1662
rect 1247 1659 1248 1660
rect 1242 1658 1248 1659
rect 1378 1659 1379 1663
rect 1383 1662 1384 1663
rect 1519 1663 1525 1664
rect 1383 1660 1457 1662
rect 1383 1659 1384 1660
rect 1378 1658 1384 1659
rect 1519 1659 1520 1663
rect 1524 1662 1525 1663
rect 1634 1663 1640 1664
rect 1524 1660 1585 1662
rect 1524 1659 1525 1660
rect 1519 1658 1525 1659
rect 1634 1659 1635 1663
rect 1639 1662 1640 1663
rect 1639 1660 1721 1662
rect 1870 1660 1871 1664
rect 1875 1660 1876 1664
rect 1639 1659 1640 1660
rect 1870 1659 1876 1660
rect 3590 1664 3596 1665
rect 3590 1660 3591 1664
rect 3595 1660 3596 1664
rect 3590 1659 3596 1660
rect 1634 1658 1640 1659
rect 110 1655 116 1656
rect 110 1651 111 1655
rect 115 1651 116 1655
rect 1830 1655 1836 1656
rect 110 1650 116 1651
rect 182 1652 188 1653
rect 182 1648 183 1652
rect 187 1648 188 1652
rect 182 1647 188 1648
rect 302 1652 308 1653
rect 302 1648 303 1652
rect 307 1648 308 1652
rect 302 1647 308 1648
rect 438 1652 444 1653
rect 438 1648 439 1652
rect 443 1648 444 1652
rect 438 1647 444 1648
rect 582 1652 588 1653
rect 582 1648 583 1652
rect 587 1648 588 1652
rect 582 1647 588 1648
rect 734 1652 740 1653
rect 734 1648 735 1652
rect 739 1648 740 1652
rect 734 1647 740 1648
rect 886 1652 892 1653
rect 886 1648 887 1652
rect 891 1648 892 1652
rect 886 1647 892 1648
rect 1030 1652 1036 1653
rect 1030 1648 1031 1652
rect 1035 1648 1036 1652
rect 1030 1647 1036 1648
rect 1174 1652 1180 1653
rect 1174 1648 1175 1652
rect 1179 1648 1180 1652
rect 1174 1647 1180 1648
rect 1310 1652 1316 1653
rect 1310 1648 1311 1652
rect 1315 1648 1316 1652
rect 1310 1647 1316 1648
rect 1438 1652 1444 1653
rect 1438 1648 1439 1652
rect 1443 1648 1444 1652
rect 1438 1647 1444 1648
rect 1566 1652 1572 1653
rect 1566 1648 1567 1652
rect 1571 1648 1572 1652
rect 1566 1647 1572 1648
rect 1702 1652 1708 1653
rect 1702 1648 1703 1652
rect 1707 1648 1708 1652
rect 1830 1651 1831 1655
rect 1835 1651 1836 1655
rect 1830 1650 1836 1651
rect 1702 1647 1708 1648
rect 1902 1646 1908 1647
rect 1902 1642 1903 1646
rect 1907 1642 1908 1646
rect 1902 1641 1908 1642
rect 1998 1646 2004 1647
rect 1998 1642 1999 1646
rect 2003 1642 2004 1646
rect 1998 1641 2004 1642
rect 2142 1646 2148 1647
rect 2142 1642 2143 1646
rect 2147 1642 2148 1646
rect 2142 1641 2148 1642
rect 2302 1646 2308 1647
rect 2302 1642 2303 1646
rect 2307 1642 2308 1646
rect 2302 1641 2308 1642
rect 2478 1646 2484 1647
rect 2478 1642 2479 1646
rect 2483 1642 2484 1646
rect 2478 1641 2484 1642
rect 2654 1646 2660 1647
rect 2654 1642 2655 1646
rect 2659 1642 2660 1646
rect 2654 1641 2660 1642
rect 2822 1646 2828 1647
rect 2822 1642 2823 1646
rect 2827 1642 2828 1646
rect 2822 1641 2828 1642
rect 2974 1646 2980 1647
rect 2974 1642 2975 1646
rect 2979 1642 2980 1646
rect 2974 1641 2980 1642
rect 3118 1646 3124 1647
rect 3118 1642 3119 1646
rect 3123 1642 3124 1646
rect 3118 1641 3124 1642
rect 3254 1646 3260 1647
rect 3254 1642 3255 1646
rect 3259 1642 3260 1646
rect 3254 1641 3260 1642
rect 3390 1646 3396 1647
rect 3390 1642 3391 1646
rect 3395 1642 3396 1646
rect 3390 1641 3396 1642
rect 3510 1646 3516 1647
rect 3510 1642 3511 1646
rect 3515 1642 3516 1646
rect 3510 1641 3516 1642
rect 918 1635 924 1636
rect 918 1631 919 1635
rect 923 1634 924 1635
rect 1047 1635 1053 1636
rect 1047 1634 1048 1635
rect 923 1632 1048 1634
rect 923 1631 924 1632
rect 918 1630 924 1631
rect 1047 1631 1048 1632
rect 1052 1631 1053 1635
rect 1047 1630 1053 1631
rect 1895 1635 1901 1636
rect 1895 1631 1896 1635
rect 1900 1634 1901 1635
rect 1910 1635 1916 1636
rect 1910 1634 1911 1635
rect 1900 1632 1911 1634
rect 1900 1631 1901 1632
rect 1895 1630 1901 1631
rect 1910 1631 1911 1632
rect 1915 1631 1916 1635
rect 1910 1630 1916 1631
rect 1962 1635 1968 1636
rect 1962 1631 1963 1635
rect 1967 1634 1968 1635
rect 1991 1635 1997 1636
rect 1991 1634 1992 1635
rect 1967 1632 1992 1634
rect 1967 1631 1968 1632
rect 1962 1630 1968 1631
rect 1991 1631 1992 1632
rect 1996 1631 1997 1635
rect 1991 1630 1997 1631
rect 2070 1635 2076 1636
rect 2070 1631 2071 1635
rect 2075 1634 2076 1635
rect 2135 1635 2141 1636
rect 2135 1634 2136 1635
rect 2075 1632 2136 1634
rect 2075 1631 2076 1632
rect 2070 1630 2076 1631
rect 2135 1631 2136 1632
rect 2140 1631 2141 1635
rect 2135 1630 2141 1631
rect 2222 1635 2228 1636
rect 2222 1631 2223 1635
rect 2227 1634 2228 1635
rect 2295 1635 2301 1636
rect 2295 1634 2296 1635
rect 2227 1632 2296 1634
rect 2227 1631 2228 1632
rect 2222 1630 2228 1631
rect 2295 1631 2296 1632
rect 2300 1631 2301 1635
rect 2295 1630 2301 1631
rect 2390 1635 2396 1636
rect 2390 1631 2391 1635
rect 2395 1634 2396 1635
rect 2471 1635 2477 1636
rect 2471 1634 2472 1635
rect 2395 1632 2472 1634
rect 2395 1631 2396 1632
rect 2390 1630 2396 1631
rect 2471 1631 2472 1632
rect 2476 1631 2477 1635
rect 2471 1630 2477 1631
rect 2566 1635 2572 1636
rect 2566 1631 2567 1635
rect 2571 1634 2572 1635
rect 2647 1635 2653 1636
rect 2647 1634 2648 1635
rect 2571 1632 2648 1634
rect 2571 1631 2572 1632
rect 2566 1630 2572 1631
rect 2647 1631 2648 1632
rect 2652 1631 2653 1635
rect 2647 1630 2653 1631
rect 2815 1635 2821 1636
rect 2815 1631 2816 1635
rect 2820 1634 2821 1635
rect 2830 1635 2836 1636
rect 2830 1634 2831 1635
rect 2820 1632 2831 1634
rect 2820 1631 2821 1632
rect 2815 1630 2821 1631
rect 2830 1631 2831 1632
rect 2835 1631 2836 1635
rect 2830 1630 2836 1631
rect 2890 1635 2896 1636
rect 2890 1631 2891 1635
rect 2895 1634 2896 1635
rect 2967 1635 2973 1636
rect 2967 1634 2968 1635
rect 2895 1632 2968 1634
rect 2895 1631 2896 1632
rect 2890 1630 2896 1631
rect 2967 1631 2968 1632
rect 2972 1631 2973 1635
rect 2967 1630 2973 1631
rect 3046 1635 3052 1636
rect 3046 1631 3047 1635
rect 3051 1634 3052 1635
rect 3111 1635 3117 1636
rect 3111 1634 3112 1635
rect 3051 1632 3112 1634
rect 3051 1631 3052 1632
rect 3046 1630 3052 1631
rect 3111 1631 3112 1632
rect 3116 1631 3117 1635
rect 3111 1630 3117 1631
rect 3247 1635 3253 1636
rect 3247 1631 3248 1635
rect 3252 1634 3253 1635
rect 3322 1635 3328 1636
rect 3322 1634 3323 1635
rect 3252 1632 3323 1634
rect 3252 1631 3253 1632
rect 3247 1630 3253 1631
rect 3322 1631 3323 1632
rect 3327 1631 3328 1635
rect 3322 1630 3328 1631
rect 3383 1635 3389 1636
rect 3383 1631 3384 1635
rect 3388 1634 3389 1635
rect 3398 1635 3404 1636
rect 3398 1634 3399 1635
rect 3388 1632 3399 1634
rect 3388 1631 3389 1632
rect 3383 1630 3389 1631
rect 3398 1631 3399 1632
rect 3403 1631 3404 1635
rect 3398 1630 3404 1631
rect 3503 1635 3509 1636
rect 3503 1631 3504 1635
rect 3508 1634 3509 1635
rect 3518 1635 3524 1636
rect 3518 1634 3519 1635
rect 3508 1632 3519 1634
rect 3508 1631 3509 1632
rect 3503 1630 3509 1631
rect 3518 1631 3519 1632
rect 3523 1631 3524 1635
rect 3518 1630 3524 1631
rect 2574 1627 2580 1628
rect 2574 1626 2575 1627
rect 2020 1624 2575 1626
rect 1967 1619 1973 1620
rect 1967 1615 1968 1619
rect 1972 1618 1973 1619
rect 2020 1618 2022 1624
rect 2574 1623 2575 1624
rect 2579 1623 2580 1627
rect 3062 1627 3068 1628
rect 3062 1626 3063 1627
rect 2574 1622 2580 1623
rect 2684 1624 3063 1626
rect 1972 1616 2022 1618
rect 2026 1619 2032 1620
rect 1972 1615 1973 1616
rect 1967 1614 1973 1615
rect 2026 1615 2027 1619
rect 2031 1618 2032 1619
rect 2087 1619 2093 1620
rect 2087 1618 2088 1619
rect 2031 1616 2088 1618
rect 2031 1615 2032 1616
rect 2026 1614 2032 1615
rect 2087 1615 2088 1616
rect 2092 1615 2093 1619
rect 2087 1614 2093 1615
rect 2198 1619 2204 1620
rect 2198 1615 2199 1619
rect 2203 1618 2204 1619
rect 2223 1619 2229 1620
rect 2223 1618 2224 1619
rect 2203 1616 2224 1618
rect 2203 1615 2204 1616
rect 2198 1614 2204 1615
rect 2223 1615 2224 1616
rect 2228 1615 2229 1619
rect 2223 1614 2229 1615
rect 2282 1619 2288 1620
rect 2282 1615 2283 1619
rect 2287 1618 2288 1619
rect 2359 1619 2365 1620
rect 2359 1618 2360 1619
rect 2287 1616 2360 1618
rect 2287 1615 2288 1616
rect 2282 1614 2288 1615
rect 2359 1615 2360 1616
rect 2364 1615 2365 1619
rect 2359 1614 2365 1615
rect 2418 1619 2424 1620
rect 2418 1615 2419 1619
rect 2423 1618 2424 1619
rect 2495 1619 2501 1620
rect 2495 1618 2496 1619
rect 2423 1616 2496 1618
rect 2423 1615 2424 1616
rect 2418 1614 2424 1615
rect 2495 1615 2496 1616
rect 2500 1615 2501 1619
rect 2495 1614 2501 1615
rect 2631 1619 2637 1620
rect 2631 1615 2632 1619
rect 2636 1618 2637 1619
rect 2684 1618 2686 1624
rect 3062 1623 3063 1624
rect 3067 1623 3068 1627
rect 3374 1627 3380 1628
rect 3374 1626 3375 1627
rect 3062 1622 3068 1623
rect 3139 1624 3375 1626
rect 2636 1616 2686 1618
rect 2690 1619 2696 1620
rect 2636 1615 2637 1616
rect 2631 1614 2637 1615
rect 2690 1615 2691 1619
rect 2695 1618 2696 1619
rect 2767 1619 2773 1620
rect 2767 1618 2768 1619
rect 2695 1616 2768 1618
rect 2695 1615 2696 1616
rect 2690 1614 2696 1615
rect 2767 1615 2768 1616
rect 2772 1615 2773 1619
rect 2767 1614 2773 1615
rect 2866 1619 2872 1620
rect 2866 1615 2867 1619
rect 2871 1618 2872 1619
rect 2903 1619 2909 1620
rect 2903 1618 2904 1619
rect 2871 1616 2904 1618
rect 2871 1615 2872 1616
rect 2866 1614 2872 1615
rect 2903 1615 2904 1616
rect 2908 1615 2909 1619
rect 2903 1614 2909 1615
rect 3047 1619 3053 1620
rect 3047 1615 3048 1619
rect 3052 1618 3053 1619
rect 3139 1618 3141 1624
rect 3374 1623 3375 1624
rect 3379 1623 3380 1627
rect 3374 1622 3380 1623
rect 3052 1616 3141 1618
rect 3178 1619 3184 1620
rect 3052 1615 3053 1616
rect 3047 1614 3053 1615
rect 3178 1615 3179 1619
rect 3183 1618 3184 1619
rect 3199 1619 3205 1620
rect 3199 1618 3200 1619
rect 3183 1616 3200 1618
rect 3183 1615 3184 1616
rect 3178 1614 3184 1615
rect 3199 1615 3200 1616
rect 3204 1615 3205 1619
rect 3199 1614 3205 1615
rect 3290 1619 3296 1620
rect 3290 1615 3291 1619
rect 3295 1618 3296 1619
rect 3359 1619 3365 1620
rect 3359 1618 3360 1619
rect 3295 1616 3360 1618
rect 3295 1615 3296 1616
rect 3290 1614 3296 1615
rect 3359 1615 3360 1616
rect 3364 1615 3365 1619
rect 3359 1614 3365 1615
rect 3486 1619 3492 1620
rect 3486 1615 3487 1619
rect 3491 1618 3492 1619
rect 3503 1619 3509 1620
rect 3503 1618 3504 1619
rect 3491 1616 3504 1618
rect 3491 1615 3492 1616
rect 3486 1614 3492 1615
rect 3503 1615 3504 1616
rect 3508 1615 3509 1619
rect 3503 1614 3509 1615
rect 1974 1610 1980 1611
rect 1974 1606 1975 1610
rect 1979 1606 1980 1610
rect 1974 1605 1980 1606
rect 2094 1610 2100 1611
rect 2094 1606 2095 1610
rect 2099 1606 2100 1610
rect 2094 1605 2100 1606
rect 2230 1610 2236 1611
rect 2230 1606 2231 1610
rect 2235 1606 2236 1610
rect 2230 1605 2236 1606
rect 2366 1610 2372 1611
rect 2366 1606 2367 1610
rect 2371 1606 2372 1610
rect 2366 1605 2372 1606
rect 2502 1610 2508 1611
rect 2502 1606 2503 1610
rect 2507 1606 2508 1610
rect 2502 1605 2508 1606
rect 2638 1610 2644 1611
rect 2638 1606 2639 1610
rect 2643 1606 2644 1610
rect 2638 1605 2644 1606
rect 2774 1610 2780 1611
rect 2774 1606 2775 1610
rect 2779 1606 2780 1610
rect 2774 1605 2780 1606
rect 2910 1610 2916 1611
rect 2910 1606 2911 1610
rect 2915 1606 2916 1610
rect 2910 1605 2916 1606
rect 3054 1610 3060 1611
rect 3054 1606 3055 1610
rect 3059 1606 3060 1610
rect 3054 1605 3060 1606
rect 3206 1610 3212 1611
rect 3206 1606 3207 1610
rect 3211 1606 3212 1610
rect 3206 1605 3212 1606
rect 3366 1610 3372 1611
rect 3366 1606 3367 1610
rect 3371 1606 3372 1610
rect 3366 1605 3372 1606
rect 3510 1610 3516 1611
rect 3510 1606 3511 1610
rect 3515 1606 3516 1610
rect 3510 1605 3516 1606
rect 166 1600 172 1601
rect 110 1597 116 1598
rect 110 1593 111 1597
rect 115 1593 116 1597
rect 166 1596 167 1600
rect 171 1596 172 1600
rect 166 1595 172 1596
rect 350 1600 356 1601
rect 350 1596 351 1600
rect 355 1596 356 1600
rect 350 1595 356 1596
rect 542 1600 548 1601
rect 542 1596 543 1600
rect 547 1596 548 1600
rect 542 1595 548 1596
rect 726 1600 732 1601
rect 726 1596 727 1600
rect 731 1596 732 1600
rect 726 1595 732 1596
rect 902 1600 908 1601
rect 902 1596 903 1600
rect 907 1596 908 1600
rect 902 1595 908 1596
rect 1070 1600 1076 1601
rect 1070 1596 1071 1600
rect 1075 1596 1076 1600
rect 1070 1595 1076 1596
rect 1222 1600 1228 1601
rect 1222 1596 1223 1600
rect 1227 1596 1228 1600
rect 1222 1595 1228 1596
rect 1358 1600 1364 1601
rect 1358 1596 1359 1600
rect 1363 1596 1364 1600
rect 1358 1595 1364 1596
rect 1494 1600 1500 1601
rect 1494 1596 1495 1600
rect 1499 1596 1500 1600
rect 1494 1595 1500 1596
rect 1622 1600 1628 1601
rect 1622 1596 1623 1600
rect 1627 1596 1628 1600
rect 1622 1595 1628 1596
rect 1742 1600 1748 1601
rect 1742 1596 1743 1600
rect 1747 1596 1748 1600
rect 1742 1595 1748 1596
rect 1830 1597 1836 1598
rect 110 1592 116 1593
rect 1830 1593 1831 1597
rect 1835 1593 1836 1597
rect 1830 1592 1836 1593
rect 1870 1592 1876 1593
rect 234 1591 240 1592
rect 174 1587 180 1588
rect 174 1583 175 1587
rect 179 1586 180 1587
rect 184 1586 186 1589
rect 234 1587 235 1591
rect 239 1590 240 1591
rect 418 1591 424 1592
rect 239 1588 369 1590
rect 239 1587 240 1588
rect 234 1586 240 1587
rect 418 1587 419 1591
rect 423 1590 424 1591
rect 610 1591 616 1592
rect 423 1588 561 1590
rect 423 1587 424 1588
rect 418 1586 424 1587
rect 610 1587 611 1591
rect 615 1590 616 1591
rect 794 1591 800 1592
rect 615 1588 745 1590
rect 615 1587 616 1588
rect 610 1586 616 1587
rect 794 1587 795 1591
rect 799 1590 800 1591
rect 1154 1591 1160 1592
rect 1154 1590 1155 1591
rect 799 1588 921 1590
rect 1133 1588 1155 1590
rect 799 1587 800 1588
rect 794 1586 800 1587
rect 1154 1587 1155 1588
rect 1159 1587 1160 1591
rect 1290 1591 1296 1592
rect 1290 1590 1291 1591
rect 1285 1588 1291 1590
rect 1154 1586 1160 1587
rect 1290 1587 1291 1588
rect 1295 1587 1296 1591
rect 1426 1591 1432 1592
rect 1426 1590 1427 1591
rect 1421 1588 1427 1590
rect 1290 1586 1296 1587
rect 1426 1587 1427 1588
rect 1431 1587 1432 1591
rect 1566 1591 1572 1592
rect 1566 1590 1567 1591
rect 1557 1588 1567 1590
rect 1426 1586 1432 1587
rect 1566 1587 1567 1588
rect 1571 1587 1572 1591
rect 1690 1591 1696 1592
rect 1690 1590 1691 1591
rect 1685 1588 1691 1590
rect 1566 1586 1572 1587
rect 1690 1587 1691 1588
rect 1695 1587 1696 1591
rect 1690 1586 1696 1587
rect 1726 1591 1732 1592
rect 1726 1587 1727 1591
rect 1731 1590 1732 1591
rect 1731 1588 1761 1590
rect 1870 1588 1871 1592
rect 1875 1588 1876 1592
rect 1731 1587 1732 1588
rect 1870 1587 1876 1588
rect 3590 1592 3596 1593
rect 3590 1588 3591 1592
rect 3595 1588 3596 1592
rect 3590 1587 3596 1588
rect 1726 1586 1732 1587
rect 179 1584 186 1586
rect 179 1583 180 1584
rect 174 1582 180 1583
rect 2026 1583 2032 1584
rect 110 1580 116 1581
rect 110 1576 111 1580
rect 115 1576 116 1580
rect 110 1575 116 1576
rect 1830 1580 1836 1581
rect 1830 1576 1831 1580
rect 1835 1576 1836 1580
rect 2026 1579 2027 1583
rect 2031 1579 2032 1583
rect 2198 1583 2204 1584
rect 2198 1582 2199 1583
rect 2149 1580 2199 1582
rect 2026 1578 2032 1579
rect 2198 1579 2199 1580
rect 2203 1579 2204 1583
rect 2198 1578 2204 1579
rect 2282 1583 2288 1584
rect 2282 1579 2283 1583
rect 2287 1579 2288 1583
rect 2282 1578 2288 1579
rect 2418 1583 2424 1584
rect 2418 1579 2419 1583
rect 2423 1579 2424 1583
rect 2418 1578 2424 1579
rect 2690 1583 2696 1584
rect 2690 1579 2691 1583
rect 2695 1579 2696 1583
rect 2866 1583 2872 1584
rect 2866 1582 2867 1583
rect 2829 1580 2867 1582
rect 2690 1578 2696 1579
rect 2866 1579 2867 1580
rect 2871 1579 2872 1583
rect 2866 1578 2872 1579
rect 2934 1583 2940 1584
rect 2934 1579 2935 1583
rect 2939 1579 2940 1583
rect 2934 1578 2940 1579
rect 3062 1583 3068 1584
rect 3062 1579 3063 1583
rect 3067 1579 3068 1583
rect 3290 1583 3296 1584
rect 3290 1582 3291 1583
rect 3261 1580 3291 1582
rect 3062 1578 3068 1579
rect 3290 1579 3291 1580
rect 3295 1579 3296 1583
rect 3290 1578 3296 1579
rect 3374 1583 3380 1584
rect 3374 1579 3375 1583
rect 3379 1579 3380 1583
rect 3374 1578 3380 1579
rect 3526 1583 3532 1584
rect 3526 1579 3527 1583
rect 3531 1579 3532 1583
rect 3526 1578 3532 1579
rect 1830 1575 1836 1576
rect 1870 1575 1876 1576
rect 1870 1571 1871 1575
rect 1875 1571 1876 1575
rect 3590 1575 3596 1576
rect 1870 1570 1876 1571
rect 1966 1572 1972 1573
rect 1966 1568 1967 1572
rect 1971 1568 1972 1572
rect 1966 1567 1972 1568
rect 2086 1572 2092 1573
rect 2086 1568 2087 1572
rect 2091 1568 2092 1572
rect 2086 1567 2092 1568
rect 2222 1572 2228 1573
rect 2222 1568 2223 1572
rect 2227 1568 2228 1572
rect 2222 1567 2228 1568
rect 2358 1572 2364 1573
rect 2358 1568 2359 1572
rect 2363 1568 2364 1572
rect 2358 1567 2364 1568
rect 2494 1572 2500 1573
rect 2494 1568 2495 1572
rect 2499 1568 2500 1572
rect 2494 1567 2500 1568
rect 2630 1572 2636 1573
rect 2630 1568 2631 1572
rect 2635 1568 2636 1572
rect 2630 1567 2636 1568
rect 2766 1572 2772 1573
rect 2766 1568 2767 1572
rect 2771 1568 2772 1572
rect 2766 1567 2772 1568
rect 2902 1572 2908 1573
rect 2902 1568 2903 1572
rect 2907 1568 2908 1572
rect 2902 1567 2908 1568
rect 3046 1572 3052 1573
rect 3046 1568 3047 1572
rect 3051 1568 3052 1572
rect 3046 1567 3052 1568
rect 3198 1572 3204 1573
rect 3198 1568 3199 1572
rect 3203 1568 3204 1572
rect 3198 1567 3204 1568
rect 3358 1572 3364 1573
rect 3358 1568 3359 1572
rect 3363 1568 3364 1572
rect 3358 1567 3364 1568
rect 3502 1572 3508 1573
rect 3502 1568 3503 1572
rect 3507 1568 3508 1572
rect 3590 1571 3591 1575
rect 3595 1571 3596 1575
rect 3590 1570 3596 1571
rect 3502 1567 3508 1568
rect 174 1562 180 1563
rect 174 1558 175 1562
rect 179 1558 180 1562
rect 174 1557 180 1558
rect 358 1562 364 1563
rect 358 1558 359 1562
rect 363 1558 364 1562
rect 358 1557 364 1558
rect 550 1562 556 1563
rect 550 1558 551 1562
rect 555 1558 556 1562
rect 550 1557 556 1558
rect 734 1562 740 1563
rect 734 1558 735 1562
rect 739 1558 740 1562
rect 734 1557 740 1558
rect 910 1562 916 1563
rect 910 1558 911 1562
rect 915 1558 916 1562
rect 910 1557 916 1558
rect 1078 1562 1084 1563
rect 1078 1558 1079 1562
rect 1083 1558 1084 1562
rect 1078 1557 1084 1558
rect 1230 1562 1236 1563
rect 1230 1558 1231 1562
rect 1235 1558 1236 1562
rect 1230 1557 1236 1558
rect 1366 1562 1372 1563
rect 1366 1558 1367 1562
rect 1371 1558 1372 1562
rect 1366 1557 1372 1558
rect 1502 1562 1508 1563
rect 1502 1558 1503 1562
rect 1507 1558 1508 1562
rect 1502 1557 1508 1558
rect 1630 1562 1636 1563
rect 1630 1558 1631 1562
rect 1635 1558 1636 1562
rect 1630 1557 1636 1558
rect 1750 1562 1756 1563
rect 1750 1558 1751 1562
rect 1755 1558 1756 1562
rect 1750 1557 1756 1558
rect 2418 1555 2424 1556
rect 167 1551 173 1552
rect 167 1547 168 1551
rect 172 1550 173 1551
rect 234 1551 240 1552
rect 234 1550 235 1551
rect 172 1548 235 1550
rect 172 1547 173 1548
rect 167 1546 173 1547
rect 234 1547 235 1548
rect 239 1547 240 1551
rect 234 1546 240 1547
rect 298 1551 304 1552
rect 298 1547 299 1551
rect 303 1550 304 1551
rect 351 1551 357 1552
rect 351 1550 352 1551
rect 303 1548 352 1550
rect 303 1547 304 1548
rect 298 1546 304 1547
rect 351 1547 352 1548
rect 356 1547 357 1551
rect 351 1546 357 1547
rect 543 1551 549 1552
rect 543 1547 544 1551
rect 548 1550 549 1551
rect 610 1551 616 1552
rect 610 1550 611 1551
rect 548 1548 611 1550
rect 548 1547 549 1548
rect 543 1546 549 1547
rect 610 1547 611 1548
rect 615 1547 616 1551
rect 610 1546 616 1547
rect 727 1551 733 1552
rect 727 1547 728 1551
rect 732 1550 733 1551
rect 794 1551 800 1552
rect 794 1550 795 1551
rect 732 1548 795 1550
rect 732 1547 733 1548
rect 727 1546 733 1547
rect 794 1547 795 1548
rect 799 1547 800 1551
rect 794 1546 800 1547
rect 903 1551 909 1552
rect 903 1547 904 1551
rect 908 1550 909 1551
rect 918 1551 924 1552
rect 918 1550 919 1551
rect 908 1548 919 1550
rect 908 1547 909 1548
rect 903 1546 909 1547
rect 918 1547 919 1548
rect 923 1547 924 1551
rect 918 1546 924 1547
rect 1071 1551 1077 1552
rect 1071 1547 1072 1551
rect 1076 1550 1077 1551
rect 1154 1551 1160 1552
rect 1076 1548 1150 1550
rect 1076 1547 1077 1548
rect 1071 1546 1077 1547
rect 1148 1542 1150 1548
rect 1154 1547 1155 1551
rect 1159 1550 1160 1551
rect 1223 1551 1229 1552
rect 1223 1550 1224 1551
rect 1159 1548 1224 1550
rect 1159 1547 1160 1548
rect 1154 1546 1160 1547
rect 1223 1547 1224 1548
rect 1228 1547 1229 1551
rect 1223 1546 1229 1547
rect 1290 1551 1296 1552
rect 1290 1547 1291 1551
rect 1295 1550 1296 1551
rect 1359 1551 1365 1552
rect 1359 1550 1360 1551
rect 1295 1548 1360 1550
rect 1295 1547 1296 1548
rect 1290 1546 1296 1547
rect 1359 1547 1360 1548
rect 1364 1547 1365 1551
rect 1359 1546 1365 1547
rect 1426 1551 1432 1552
rect 1426 1547 1427 1551
rect 1431 1550 1432 1551
rect 1495 1551 1501 1552
rect 1495 1550 1496 1551
rect 1431 1548 1496 1550
rect 1431 1547 1432 1548
rect 1426 1546 1432 1547
rect 1495 1547 1496 1548
rect 1500 1547 1501 1551
rect 1495 1546 1501 1547
rect 1566 1551 1572 1552
rect 1566 1547 1567 1551
rect 1571 1550 1572 1551
rect 1623 1551 1629 1552
rect 1623 1550 1624 1551
rect 1571 1548 1624 1550
rect 1571 1547 1572 1548
rect 1566 1546 1572 1547
rect 1623 1547 1624 1548
rect 1628 1547 1629 1551
rect 1623 1546 1629 1547
rect 1690 1551 1696 1552
rect 1690 1547 1691 1551
rect 1695 1550 1696 1551
rect 1743 1551 1749 1552
rect 1743 1550 1744 1551
rect 1695 1548 1744 1550
rect 1695 1547 1696 1548
rect 1690 1546 1696 1547
rect 1743 1547 1744 1548
rect 1748 1547 1749 1551
rect 2418 1551 2419 1555
rect 2423 1554 2424 1555
rect 2511 1555 2517 1556
rect 2511 1554 2512 1555
rect 2423 1552 2512 1554
rect 2423 1551 2424 1552
rect 2418 1550 2424 1551
rect 2511 1551 2512 1552
rect 2516 1551 2517 1555
rect 2511 1550 2517 1551
rect 1743 1546 1749 1547
rect 1478 1543 1484 1544
rect 1478 1542 1479 1543
rect 1148 1540 1479 1542
rect 1478 1539 1479 1540
rect 1483 1539 1484 1543
rect 1478 1538 1484 1539
rect 127 1535 133 1536
rect 127 1531 128 1535
rect 132 1534 133 1535
rect 135 1535 141 1536
rect 135 1534 136 1535
rect 132 1532 136 1534
rect 132 1531 133 1532
rect 127 1530 133 1531
rect 135 1531 136 1532
rect 140 1531 141 1535
rect 135 1530 141 1531
rect 194 1535 200 1536
rect 194 1531 195 1535
rect 199 1534 200 1535
rect 239 1535 245 1536
rect 239 1534 240 1535
rect 199 1532 240 1534
rect 199 1531 200 1532
rect 194 1530 200 1531
rect 239 1531 240 1532
rect 244 1531 245 1535
rect 239 1530 245 1531
rect 375 1535 381 1536
rect 375 1531 376 1535
rect 380 1534 381 1535
rect 418 1535 424 1536
rect 418 1534 419 1535
rect 380 1532 419 1534
rect 380 1531 381 1532
rect 375 1530 381 1531
rect 418 1531 419 1532
rect 423 1531 424 1535
rect 418 1530 424 1531
rect 434 1535 440 1536
rect 434 1531 435 1535
rect 439 1534 440 1535
rect 519 1535 525 1536
rect 519 1534 520 1535
rect 439 1532 520 1534
rect 439 1531 440 1532
rect 434 1530 440 1531
rect 519 1531 520 1532
rect 524 1531 525 1535
rect 519 1530 525 1531
rect 578 1535 584 1536
rect 578 1531 579 1535
rect 583 1534 584 1535
rect 663 1535 669 1536
rect 663 1534 664 1535
rect 583 1532 664 1534
rect 583 1531 584 1532
rect 578 1530 584 1531
rect 663 1531 664 1532
rect 668 1531 669 1535
rect 663 1530 669 1531
rect 722 1535 728 1536
rect 722 1531 723 1535
rect 727 1534 728 1535
rect 807 1535 813 1536
rect 807 1534 808 1535
rect 727 1532 808 1534
rect 727 1531 728 1532
rect 722 1530 728 1531
rect 807 1531 808 1532
rect 812 1531 813 1535
rect 807 1530 813 1531
rect 943 1535 949 1536
rect 943 1531 944 1535
rect 948 1534 949 1535
rect 958 1535 964 1536
rect 958 1534 959 1535
rect 948 1532 959 1534
rect 948 1531 949 1532
rect 943 1530 949 1531
rect 958 1531 959 1532
rect 963 1531 964 1535
rect 958 1530 964 1531
rect 1002 1535 1008 1536
rect 1002 1531 1003 1535
rect 1007 1534 1008 1535
rect 1071 1535 1077 1536
rect 1071 1534 1072 1535
rect 1007 1532 1072 1534
rect 1007 1531 1008 1532
rect 1002 1530 1008 1531
rect 1071 1531 1072 1532
rect 1076 1531 1077 1535
rect 1071 1530 1077 1531
rect 1130 1535 1136 1536
rect 1130 1531 1131 1535
rect 1135 1534 1136 1535
rect 1199 1535 1205 1536
rect 1199 1534 1200 1535
rect 1135 1532 1200 1534
rect 1135 1531 1136 1532
rect 1130 1530 1136 1531
rect 1199 1531 1200 1532
rect 1204 1531 1205 1535
rect 1199 1530 1205 1531
rect 1258 1535 1264 1536
rect 1258 1531 1259 1535
rect 1263 1534 1264 1535
rect 1327 1535 1333 1536
rect 1327 1534 1328 1535
rect 1263 1532 1328 1534
rect 1263 1531 1264 1532
rect 1258 1530 1264 1531
rect 1327 1531 1328 1532
rect 1332 1531 1333 1535
rect 1327 1530 1333 1531
rect 1386 1535 1392 1536
rect 1386 1531 1387 1535
rect 1391 1534 1392 1535
rect 1463 1535 1469 1536
rect 1463 1534 1464 1535
rect 1391 1532 1464 1534
rect 1391 1531 1392 1532
rect 1386 1530 1392 1531
rect 1463 1531 1464 1532
rect 1468 1531 1469 1535
rect 1463 1530 1469 1531
rect 142 1526 148 1527
rect 142 1522 143 1526
rect 147 1522 148 1526
rect 142 1521 148 1522
rect 246 1526 252 1527
rect 246 1522 247 1526
rect 251 1522 252 1526
rect 246 1521 252 1522
rect 382 1526 388 1527
rect 382 1522 383 1526
rect 387 1522 388 1526
rect 382 1521 388 1522
rect 526 1526 532 1527
rect 526 1522 527 1526
rect 531 1522 532 1526
rect 526 1521 532 1522
rect 670 1526 676 1527
rect 670 1522 671 1526
rect 675 1522 676 1526
rect 670 1521 676 1522
rect 814 1526 820 1527
rect 814 1522 815 1526
rect 819 1522 820 1526
rect 814 1521 820 1522
rect 950 1526 956 1527
rect 950 1522 951 1526
rect 955 1522 956 1526
rect 950 1521 956 1522
rect 1078 1526 1084 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1206 1526 1212 1527
rect 1206 1522 1207 1526
rect 1211 1522 1212 1526
rect 1206 1521 1212 1522
rect 1334 1526 1340 1527
rect 1334 1522 1335 1526
rect 1339 1522 1340 1526
rect 1334 1521 1340 1522
rect 1470 1526 1476 1527
rect 1470 1522 1471 1526
rect 1475 1522 1476 1526
rect 2086 1524 2092 1525
rect 1470 1521 1476 1522
rect 1870 1521 1876 1522
rect 1870 1517 1871 1521
rect 1875 1517 1876 1521
rect 2086 1520 2087 1524
rect 2091 1520 2092 1524
rect 2086 1519 2092 1520
rect 2166 1524 2172 1525
rect 2166 1520 2167 1524
rect 2171 1520 2172 1524
rect 2166 1519 2172 1520
rect 2254 1524 2260 1525
rect 2254 1520 2255 1524
rect 2259 1520 2260 1524
rect 2254 1519 2260 1520
rect 2342 1524 2348 1525
rect 2342 1520 2343 1524
rect 2347 1520 2348 1524
rect 2342 1519 2348 1520
rect 2438 1524 2444 1525
rect 2438 1520 2439 1524
rect 2443 1520 2444 1524
rect 2438 1519 2444 1520
rect 2534 1524 2540 1525
rect 2534 1520 2535 1524
rect 2539 1520 2540 1524
rect 2534 1519 2540 1520
rect 2646 1524 2652 1525
rect 2646 1520 2647 1524
rect 2651 1520 2652 1524
rect 2646 1519 2652 1520
rect 2782 1524 2788 1525
rect 2782 1520 2783 1524
rect 2787 1520 2788 1524
rect 2782 1519 2788 1520
rect 2942 1524 2948 1525
rect 2942 1520 2943 1524
rect 2947 1520 2948 1524
rect 2942 1519 2948 1520
rect 3118 1524 3124 1525
rect 3118 1520 3119 1524
rect 3123 1520 3124 1524
rect 3118 1519 3124 1520
rect 3302 1524 3308 1525
rect 3302 1520 3303 1524
rect 3307 1520 3308 1524
rect 3302 1519 3308 1520
rect 3494 1524 3500 1525
rect 3494 1520 3495 1524
rect 3499 1520 3500 1524
rect 3494 1519 3500 1520
rect 3590 1521 3596 1522
rect 1870 1516 1876 1517
rect 3590 1517 3591 1521
rect 3595 1517 3596 1521
rect 3590 1516 3596 1517
rect 2154 1515 2160 1516
rect 2154 1514 2155 1515
rect 2149 1512 2155 1514
rect 2154 1511 2155 1512
rect 2159 1511 2160 1515
rect 2234 1515 2240 1516
rect 2234 1514 2235 1515
rect 2229 1512 2235 1514
rect 2154 1510 2160 1511
rect 2234 1511 2235 1512
rect 2239 1511 2240 1515
rect 2322 1515 2328 1516
rect 2322 1514 2323 1515
rect 2317 1512 2323 1514
rect 2234 1510 2240 1511
rect 2322 1511 2323 1512
rect 2327 1511 2328 1515
rect 2410 1515 2416 1516
rect 2410 1514 2411 1515
rect 2405 1512 2411 1514
rect 2322 1510 2328 1511
rect 2410 1511 2411 1512
rect 2415 1511 2416 1515
rect 2506 1515 2512 1516
rect 2506 1514 2507 1515
rect 2501 1512 2507 1514
rect 2410 1510 2416 1511
rect 2506 1511 2507 1512
rect 2511 1511 2512 1515
rect 2722 1515 2728 1516
rect 2722 1514 2723 1515
rect 2539 1512 2553 1514
rect 2709 1512 2723 1514
rect 2506 1510 2512 1511
rect 2514 1511 2520 1512
rect 110 1508 116 1509
rect 110 1504 111 1508
rect 115 1504 116 1508
rect 110 1503 116 1504
rect 1830 1508 1836 1509
rect 1830 1504 1831 1508
rect 1835 1504 1836 1508
rect 2514 1507 2515 1511
rect 2519 1510 2520 1511
rect 2539 1510 2541 1512
rect 2722 1511 2723 1512
rect 2727 1511 2728 1515
rect 2850 1515 2856 1516
rect 2850 1514 2851 1515
rect 2845 1512 2851 1514
rect 2722 1510 2728 1511
rect 2850 1511 2851 1512
rect 2855 1511 2856 1515
rect 3038 1515 3044 1516
rect 3038 1514 3039 1515
rect 3005 1512 3039 1514
rect 2850 1510 2856 1511
rect 3038 1511 3039 1512
rect 3043 1511 3044 1515
rect 3194 1515 3200 1516
rect 3194 1514 3195 1515
rect 3181 1512 3195 1514
rect 3038 1510 3044 1511
rect 3194 1511 3195 1512
rect 3199 1511 3200 1515
rect 3194 1510 3200 1511
rect 3202 1515 3208 1516
rect 3202 1511 3203 1515
rect 3207 1514 3208 1515
rect 3479 1515 3485 1516
rect 3207 1512 3321 1514
rect 3207 1511 3208 1512
rect 3202 1510 3208 1511
rect 3479 1511 3480 1515
rect 3484 1514 3485 1515
rect 3484 1512 3513 1514
rect 3484 1511 3485 1512
rect 3479 1510 3485 1511
rect 2519 1508 2541 1510
rect 2519 1507 2520 1508
rect 2514 1506 2520 1507
rect 1830 1503 1836 1504
rect 1870 1504 1876 1505
rect 1870 1500 1871 1504
rect 1875 1500 1876 1504
rect 194 1499 200 1500
rect 194 1495 195 1499
rect 199 1495 200 1499
rect 194 1494 200 1495
rect 298 1499 304 1500
rect 298 1495 299 1499
rect 303 1495 304 1499
rect 298 1494 304 1495
rect 434 1499 440 1500
rect 434 1495 435 1499
rect 439 1495 440 1499
rect 434 1494 440 1495
rect 578 1499 584 1500
rect 578 1495 579 1499
rect 583 1495 584 1499
rect 578 1494 584 1495
rect 722 1499 728 1500
rect 722 1495 723 1499
rect 727 1495 728 1499
rect 722 1494 728 1495
rect 1002 1499 1008 1500
rect 1002 1495 1003 1499
rect 1007 1495 1008 1499
rect 1002 1494 1008 1495
rect 1130 1499 1136 1500
rect 1130 1495 1131 1499
rect 1135 1495 1136 1499
rect 1130 1494 1136 1495
rect 1258 1499 1264 1500
rect 1258 1495 1259 1499
rect 1263 1495 1264 1499
rect 1258 1494 1264 1495
rect 1386 1499 1392 1500
rect 1386 1495 1387 1499
rect 1391 1495 1392 1499
rect 1386 1494 1392 1495
rect 1478 1499 1484 1500
rect 1870 1499 1876 1500
rect 3590 1504 3596 1505
rect 3590 1500 3591 1504
rect 3595 1500 3596 1504
rect 3590 1499 3596 1500
rect 1478 1495 1479 1499
rect 1483 1495 1484 1499
rect 1478 1494 1484 1495
rect 110 1491 116 1492
rect 110 1487 111 1491
rect 115 1487 116 1491
rect 1830 1491 1836 1492
rect 110 1486 116 1487
rect 134 1488 140 1489
rect 134 1484 135 1488
rect 139 1484 140 1488
rect 134 1483 140 1484
rect 238 1488 244 1489
rect 238 1484 239 1488
rect 243 1484 244 1488
rect 238 1483 244 1484
rect 374 1488 380 1489
rect 374 1484 375 1488
rect 379 1484 380 1488
rect 374 1483 380 1484
rect 518 1488 524 1489
rect 518 1484 519 1488
rect 523 1484 524 1488
rect 518 1483 524 1484
rect 662 1488 668 1489
rect 662 1484 663 1488
rect 667 1484 668 1488
rect 662 1483 668 1484
rect 806 1488 812 1489
rect 806 1484 807 1488
rect 811 1484 812 1488
rect 806 1483 812 1484
rect 942 1488 948 1489
rect 942 1484 943 1488
rect 947 1484 948 1488
rect 942 1483 948 1484
rect 1070 1488 1076 1489
rect 1070 1484 1071 1488
rect 1075 1484 1076 1488
rect 1070 1483 1076 1484
rect 1198 1488 1204 1489
rect 1198 1484 1199 1488
rect 1203 1484 1204 1488
rect 1198 1483 1204 1484
rect 1326 1488 1332 1489
rect 1326 1484 1327 1488
rect 1331 1484 1332 1488
rect 1326 1483 1332 1484
rect 1462 1488 1468 1489
rect 1462 1484 1463 1488
rect 1467 1484 1468 1488
rect 1830 1487 1831 1491
rect 1835 1487 1836 1491
rect 1830 1486 1836 1487
rect 2094 1486 2100 1487
rect 1462 1483 1468 1484
rect 2094 1482 2095 1486
rect 2099 1482 2100 1486
rect 2094 1481 2100 1482
rect 2174 1486 2180 1487
rect 2174 1482 2175 1486
rect 2179 1482 2180 1486
rect 2174 1481 2180 1482
rect 2262 1486 2268 1487
rect 2262 1482 2263 1486
rect 2267 1482 2268 1486
rect 2262 1481 2268 1482
rect 2350 1486 2356 1487
rect 2350 1482 2351 1486
rect 2355 1482 2356 1486
rect 2350 1481 2356 1482
rect 2446 1486 2452 1487
rect 2446 1482 2447 1486
rect 2451 1482 2452 1486
rect 2446 1481 2452 1482
rect 2542 1486 2548 1487
rect 2542 1482 2543 1486
rect 2547 1482 2548 1486
rect 2542 1481 2548 1482
rect 2654 1486 2660 1487
rect 2654 1482 2655 1486
rect 2659 1482 2660 1486
rect 2654 1481 2660 1482
rect 2790 1486 2796 1487
rect 2790 1482 2791 1486
rect 2795 1482 2796 1486
rect 2790 1481 2796 1482
rect 2950 1486 2956 1487
rect 2950 1482 2951 1486
rect 2955 1482 2956 1486
rect 2950 1481 2956 1482
rect 3126 1486 3132 1487
rect 3126 1482 3127 1486
rect 3131 1482 3132 1486
rect 3126 1481 3132 1482
rect 3310 1486 3316 1487
rect 3310 1482 3311 1486
rect 3315 1482 3316 1486
rect 3310 1481 3316 1482
rect 3502 1486 3508 1487
rect 3502 1482 3503 1486
rect 3507 1482 3508 1486
rect 3502 1481 3508 1482
rect 2087 1475 2093 1476
rect 614 1471 620 1472
rect 614 1467 615 1471
rect 619 1470 620 1471
rect 823 1471 829 1472
rect 823 1470 824 1471
rect 619 1468 824 1470
rect 619 1467 620 1468
rect 614 1466 620 1467
rect 823 1467 824 1468
rect 828 1467 829 1471
rect 2087 1471 2088 1475
rect 2092 1474 2093 1475
rect 2102 1475 2108 1476
rect 2102 1474 2103 1475
rect 2092 1472 2103 1474
rect 2092 1471 2093 1472
rect 2087 1470 2093 1471
rect 2102 1471 2103 1472
rect 2107 1471 2108 1475
rect 2102 1470 2108 1471
rect 2154 1475 2160 1476
rect 2154 1471 2155 1475
rect 2159 1474 2160 1475
rect 2167 1475 2173 1476
rect 2167 1474 2168 1475
rect 2159 1472 2168 1474
rect 2159 1471 2160 1472
rect 2154 1470 2160 1471
rect 2167 1471 2168 1472
rect 2172 1471 2173 1475
rect 2167 1470 2173 1471
rect 2234 1475 2240 1476
rect 2234 1471 2235 1475
rect 2239 1474 2240 1475
rect 2255 1475 2261 1476
rect 2255 1474 2256 1475
rect 2239 1472 2256 1474
rect 2239 1471 2240 1472
rect 2234 1470 2240 1471
rect 2255 1471 2256 1472
rect 2260 1471 2261 1475
rect 2255 1470 2261 1471
rect 2322 1475 2328 1476
rect 2322 1471 2323 1475
rect 2327 1474 2328 1475
rect 2343 1475 2349 1476
rect 2343 1474 2344 1475
rect 2327 1472 2344 1474
rect 2327 1471 2328 1472
rect 2322 1470 2328 1471
rect 2343 1471 2344 1472
rect 2348 1471 2349 1475
rect 2343 1470 2349 1471
rect 2410 1475 2416 1476
rect 2410 1471 2411 1475
rect 2415 1474 2416 1475
rect 2439 1475 2445 1476
rect 2439 1474 2440 1475
rect 2415 1472 2440 1474
rect 2415 1471 2416 1472
rect 2410 1470 2416 1471
rect 2439 1471 2440 1472
rect 2444 1471 2445 1475
rect 2439 1470 2445 1471
rect 2506 1475 2512 1476
rect 2506 1471 2507 1475
rect 2511 1474 2512 1475
rect 2535 1475 2541 1476
rect 2535 1474 2536 1475
rect 2511 1472 2536 1474
rect 2511 1471 2512 1472
rect 2506 1470 2512 1471
rect 2535 1471 2536 1472
rect 2540 1471 2541 1475
rect 2535 1470 2541 1471
rect 2647 1475 2653 1476
rect 2647 1471 2648 1475
rect 2652 1474 2653 1475
rect 2662 1475 2668 1476
rect 2662 1474 2663 1475
rect 2652 1472 2663 1474
rect 2652 1471 2653 1472
rect 2647 1470 2653 1471
rect 2662 1471 2663 1472
rect 2667 1471 2668 1475
rect 2662 1470 2668 1471
rect 2722 1475 2728 1476
rect 2722 1471 2723 1475
rect 2727 1474 2728 1475
rect 2783 1475 2789 1476
rect 2783 1474 2784 1475
rect 2727 1472 2784 1474
rect 2727 1471 2728 1472
rect 2722 1470 2728 1471
rect 2783 1471 2784 1472
rect 2788 1471 2789 1475
rect 2783 1470 2789 1471
rect 2934 1475 2940 1476
rect 2934 1471 2935 1475
rect 2939 1474 2940 1475
rect 2943 1475 2949 1476
rect 2943 1474 2944 1475
rect 2939 1472 2944 1474
rect 2939 1471 2940 1472
rect 2934 1470 2940 1471
rect 2943 1471 2944 1472
rect 2948 1471 2949 1475
rect 2943 1470 2949 1471
rect 3038 1475 3044 1476
rect 3038 1471 3039 1475
rect 3043 1474 3044 1475
rect 3119 1475 3125 1476
rect 3119 1474 3120 1475
rect 3043 1472 3120 1474
rect 3043 1471 3044 1472
rect 3038 1470 3044 1471
rect 3119 1471 3120 1472
rect 3124 1471 3125 1475
rect 3119 1470 3125 1471
rect 3194 1475 3200 1476
rect 3194 1471 3195 1475
rect 3199 1474 3200 1475
rect 3303 1475 3309 1476
rect 3303 1474 3304 1475
rect 3199 1472 3304 1474
rect 3199 1471 3200 1472
rect 3194 1470 3200 1471
rect 3303 1471 3304 1472
rect 3308 1471 3309 1475
rect 3303 1470 3309 1471
rect 3487 1475 3493 1476
rect 3487 1471 3488 1475
rect 3492 1474 3493 1475
rect 3495 1475 3501 1476
rect 3495 1474 3496 1475
rect 3492 1472 3496 1474
rect 3492 1471 3493 1472
rect 3487 1470 3493 1471
rect 3495 1471 3496 1472
rect 3500 1471 3501 1475
rect 3495 1470 3501 1471
rect 823 1466 829 1467
rect 2255 1459 2261 1460
rect 2255 1455 2256 1459
rect 2260 1458 2261 1459
rect 2270 1459 2276 1460
rect 2270 1458 2271 1459
rect 2260 1456 2271 1458
rect 2260 1455 2261 1456
rect 2255 1454 2261 1455
rect 2270 1455 2271 1456
rect 2275 1455 2276 1459
rect 2270 1454 2276 1455
rect 2314 1459 2320 1460
rect 2314 1455 2315 1459
rect 2319 1458 2320 1459
rect 2335 1459 2341 1460
rect 2335 1458 2336 1459
rect 2319 1456 2336 1458
rect 2319 1455 2320 1456
rect 2314 1454 2320 1455
rect 2335 1455 2336 1456
rect 2340 1455 2341 1459
rect 2335 1454 2341 1455
rect 2394 1459 2400 1460
rect 2394 1455 2395 1459
rect 2399 1458 2400 1459
rect 2415 1459 2421 1460
rect 2415 1458 2416 1459
rect 2399 1456 2416 1458
rect 2399 1455 2400 1456
rect 2394 1454 2400 1455
rect 2415 1455 2416 1456
rect 2420 1455 2421 1459
rect 2415 1454 2421 1455
rect 2474 1459 2480 1460
rect 2474 1455 2475 1459
rect 2479 1458 2480 1459
rect 2495 1459 2501 1460
rect 2495 1458 2496 1459
rect 2479 1456 2496 1458
rect 2479 1455 2480 1456
rect 2474 1454 2480 1455
rect 2495 1455 2496 1456
rect 2500 1455 2501 1459
rect 2495 1454 2501 1455
rect 2599 1459 2605 1460
rect 2599 1455 2600 1459
rect 2604 1458 2605 1459
rect 2666 1459 2672 1460
rect 2666 1458 2667 1459
rect 2604 1456 2667 1458
rect 2604 1455 2605 1456
rect 2599 1454 2605 1455
rect 2666 1455 2667 1456
rect 2671 1455 2672 1459
rect 2666 1454 2672 1455
rect 2727 1459 2733 1460
rect 2727 1455 2728 1459
rect 2732 1458 2733 1459
rect 2842 1459 2848 1460
rect 2842 1458 2843 1459
rect 2732 1456 2843 1458
rect 2732 1455 2733 1456
rect 2727 1454 2733 1455
rect 2842 1455 2843 1456
rect 2847 1455 2848 1459
rect 2842 1454 2848 1455
rect 2850 1459 2856 1460
rect 2850 1455 2851 1459
rect 2855 1458 2856 1459
rect 2887 1459 2893 1460
rect 2887 1458 2888 1459
rect 2855 1456 2888 1458
rect 2855 1455 2856 1456
rect 2850 1454 2856 1455
rect 2887 1455 2888 1456
rect 2892 1455 2893 1459
rect 2887 1454 2893 1455
rect 3070 1459 3077 1460
rect 3070 1455 3071 1459
rect 3076 1455 3077 1459
rect 3070 1454 3077 1455
rect 3190 1459 3196 1460
rect 3190 1455 3191 1459
rect 3195 1458 3196 1459
rect 3271 1459 3277 1460
rect 3271 1458 3272 1459
rect 3195 1456 3272 1458
rect 3195 1455 3196 1456
rect 3190 1454 3196 1455
rect 3271 1455 3272 1456
rect 3276 1455 3277 1459
rect 3271 1454 3277 1455
rect 3471 1459 3477 1460
rect 3471 1455 3472 1459
rect 3476 1458 3477 1459
rect 3479 1459 3485 1460
rect 3479 1458 3480 1459
rect 3476 1456 3480 1458
rect 3476 1455 3477 1456
rect 3471 1454 3477 1455
rect 3479 1455 3480 1456
rect 3484 1455 3485 1459
rect 3479 1454 3485 1455
rect 2262 1450 2268 1451
rect 2262 1446 2263 1450
rect 2267 1446 2268 1450
rect 2262 1445 2268 1446
rect 2342 1450 2348 1451
rect 2342 1446 2343 1450
rect 2347 1446 2348 1450
rect 2342 1445 2348 1446
rect 2422 1450 2428 1451
rect 2422 1446 2423 1450
rect 2427 1446 2428 1450
rect 2422 1445 2428 1446
rect 2502 1450 2508 1451
rect 2502 1446 2503 1450
rect 2507 1446 2508 1450
rect 2502 1445 2508 1446
rect 2606 1450 2612 1451
rect 2606 1446 2607 1450
rect 2611 1446 2612 1450
rect 2606 1445 2612 1446
rect 2734 1450 2740 1451
rect 2734 1446 2735 1450
rect 2739 1446 2740 1450
rect 2734 1445 2740 1446
rect 2894 1450 2900 1451
rect 2894 1446 2895 1450
rect 2899 1446 2900 1450
rect 2894 1445 2900 1446
rect 3078 1450 3084 1451
rect 3078 1446 3079 1450
rect 3083 1446 3084 1450
rect 3078 1445 3084 1446
rect 3278 1450 3284 1451
rect 3278 1446 3279 1450
rect 3283 1446 3284 1450
rect 3278 1445 3284 1446
rect 3478 1450 3484 1451
rect 3478 1446 3479 1450
rect 3483 1446 3484 1450
rect 3478 1445 3484 1446
rect 134 1440 140 1441
rect 110 1437 116 1438
rect 110 1433 111 1437
rect 115 1433 116 1437
rect 134 1436 135 1440
rect 139 1436 140 1440
rect 134 1435 140 1436
rect 230 1440 236 1441
rect 230 1436 231 1440
rect 235 1436 236 1440
rect 230 1435 236 1436
rect 358 1440 364 1441
rect 358 1436 359 1440
rect 363 1436 364 1440
rect 358 1435 364 1436
rect 478 1440 484 1441
rect 478 1436 479 1440
rect 483 1436 484 1440
rect 478 1435 484 1436
rect 598 1440 604 1441
rect 598 1436 599 1440
rect 603 1436 604 1440
rect 598 1435 604 1436
rect 718 1440 724 1441
rect 718 1436 719 1440
rect 723 1436 724 1440
rect 718 1435 724 1436
rect 830 1440 836 1441
rect 830 1436 831 1440
rect 835 1436 836 1440
rect 830 1435 836 1436
rect 934 1440 940 1441
rect 934 1436 935 1440
rect 939 1436 940 1440
rect 934 1435 940 1436
rect 1038 1440 1044 1441
rect 1038 1436 1039 1440
rect 1043 1436 1044 1440
rect 1038 1435 1044 1436
rect 1142 1440 1148 1441
rect 1142 1436 1143 1440
rect 1147 1436 1148 1440
rect 1142 1435 1148 1436
rect 1254 1440 1260 1441
rect 1254 1436 1255 1440
rect 1259 1436 1260 1440
rect 1254 1435 1260 1436
rect 1830 1437 1836 1438
rect 110 1432 116 1433
rect 1830 1433 1831 1437
rect 1835 1433 1836 1437
rect 1830 1432 1836 1433
rect 1870 1432 1876 1433
rect 127 1431 133 1432
rect 127 1427 128 1431
rect 132 1430 133 1431
rect 202 1431 208 1432
rect 132 1428 153 1430
rect 132 1427 133 1428
rect 127 1426 133 1427
rect 202 1427 203 1431
rect 207 1430 208 1431
rect 298 1431 304 1432
rect 207 1428 249 1430
rect 207 1427 208 1428
rect 202 1426 208 1427
rect 298 1427 299 1431
rect 303 1430 304 1431
rect 426 1431 432 1432
rect 303 1428 377 1430
rect 303 1427 304 1428
rect 298 1426 304 1427
rect 426 1427 427 1431
rect 431 1430 432 1431
rect 546 1431 552 1432
rect 431 1428 497 1430
rect 431 1427 432 1428
rect 426 1426 432 1427
rect 546 1427 547 1431
rect 551 1430 552 1431
rect 786 1431 792 1432
rect 786 1430 787 1431
rect 551 1428 617 1430
rect 781 1428 787 1430
rect 551 1427 552 1428
rect 546 1426 552 1427
rect 786 1427 787 1428
rect 791 1427 792 1431
rect 898 1431 904 1432
rect 898 1430 899 1431
rect 893 1428 899 1430
rect 786 1426 792 1427
rect 898 1427 899 1428
rect 903 1427 904 1431
rect 1002 1431 1008 1432
rect 1002 1430 1003 1431
rect 997 1428 1003 1430
rect 898 1426 904 1427
rect 1002 1427 1003 1428
rect 1007 1427 1008 1431
rect 1106 1431 1112 1432
rect 1106 1430 1107 1431
rect 1101 1428 1107 1430
rect 1002 1426 1008 1427
rect 1106 1427 1107 1428
rect 1111 1427 1112 1431
rect 1210 1431 1216 1432
rect 1210 1430 1211 1431
rect 1205 1428 1211 1430
rect 1106 1426 1112 1427
rect 1210 1427 1211 1428
rect 1215 1427 1216 1431
rect 1210 1426 1216 1427
rect 1218 1431 1224 1432
rect 1218 1427 1219 1431
rect 1223 1430 1224 1431
rect 1223 1428 1273 1430
rect 1870 1428 1871 1432
rect 1875 1428 1876 1432
rect 1223 1427 1224 1428
rect 1870 1427 1876 1428
rect 3590 1432 3596 1433
rect 3590 1428 3591 1432
rect 3595 1428 3596 1432
rect 3590 1427 3596 1428
rect 1218 1426 1224 1427
rect 2314 1423 2320 1424
rect 110 1420 116 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 110 1415 116 1416
rect 1830 1420 1836 1421
rect 1830 1416 1831 1420
rect 1835 1416 1836 1420
rect 2314 1419 2315 1423
rect 2319 1419 2320 1423
rect 2314 1418 2320 1419
rect 2394 1423 2400 1424
rect 2394 1419 2395 1423
rect 2399 1419 2400 1423
rect 2394 1418 2400 1419
rect 2474 1423 2480 1424
rect 2474 1419 2475 1423
rect 2479 1419 2480 1423
rect 2474 1418 2480 1419
rect 2666 1423 2672 1424
rect 2666 1419 2667 1423
rect 2671 1422 2672 1423
rect 3070 1423 3076 1424
rect 3070 1422 3071 1423
rect 2671 1420 2745 1422
rect 2949 1420 3071 1422
rect 2671 1419 2672 1420
rect 2666 1418 2672 1419
rect 3070 1419 3071 1420
rect 3075 1419 3076 1423
rect 3190 1423 3196 1424
rect 3190 1422 3191 1423
rect 3133 1420 3191 1422
rect 3070 1418 3076 1419
rect 3190 1419 3191 1420
rect 3195 1419 3196 1423
rect 3190 1418 3196 1419
rect 3286 1423 3292 1424
rect 3286 1419 3287 1423
rect 3291 1419 3292 1423
rect 3286 1418 3292 1419
rect 1830 1415 1836 1416
rect 1870 1415 1876 1416
rect 1870 1411 1871 1415
rect 1875 1411 1876 1415
rect 3590 1415 3596 1416
rect 1870 1410 1876 1411
rect 2254 1412 2260 1413
rect 2254 1408 2255 1412
rect 2259 1408 2260 1412
rect 2254 1407 2260 1408
rect 2334 1412 2340 1413
rect 2334 1408 2335 1412
rect 2339 1408 2340 1412
rect 2334 1407 2340 1408
rect 2414 1412 2420 1413
rect 2414 1408 2415 1412
rect 2419 1408 2420 1412
rect 2414 1407 2420 1408
rect 2494 1412 2500 1413
rect 2494 1408 2495 1412
rect 2499 1408 2500 1412
rect 2494 1407 2500 1408
rect 2598 1412 2604 1413
rect 2598 1408 2599 1412
rect 2603 1408 2604 1412
rect 2598 1407 2604 1408
rect 2726 1412 2732 1413
rect 2726 1408 2727 1412
rect 2731 1408 2732 1412
rect 2726 1407 2732 1408
rect 2886 1412 2892 1413
rect 2886 1408 2887 1412
rect 2891 1408 2892 1412
rect 2886 1407 2892 1408
rect 3070 1412 3076 1413
rect 3070 1408 3071 1412
rect 3075 1408 3076 1412
rect 3070 1407 3076 1408
rect 3270 1412 3276 1413
rect 3270 1408 3271 1412
rect 3275 1408 3276 1412
rect 3270 1407 3276 1408
rect 3470 1412 3476 1413
rect 3470 1408 3471 1412
rect 3475 1408 3476 1412
rect 3590 1411 3591 1415
rect 3595 1411 3596 1415
rect 3590 1410 3596 1411
rect 3470 1407 3476 1408
rect 142 1402 148 1403
rect 142 1398 143 1402
rect 147 1398 148 1402
rect 238 1402 244 1403
rect 202 1399 208 1400
rect 202 1398 203 1399
rect 142 1397 148 1398
rect 188 1396 203 1398
rect 135 1391 141 1392
rect 135 1387 136 1391
rect 140 1390 141 1391
rect 188 1390 190 1396
rect 202 1395 203 1396
rect 207 1395 208 1399
rect 238 1398 239 1402
rect 243 1398 244 1402
rect 238 1397 244 1398
rect 366 1402 372 1403
rect 366 1398 367 1402
rect 371 1398 372 1402
rect 366 1397 372 1398
rect 486 1402 492 1403
rect 486 1398 487 1402
rect 491 1398 492 1402
rect 486 1397 492 1398
rect 606 1402 612 1403
rect 606 1398 607 1402
rect 611 1398 612 1402
rect 606 1397 612 1398
rect 726 1402 732 1403
rect 726 1398 727 1402
rect 731 1398 732 1402
rect 726 1397 732 1398
rect 838 1402 844 1403
rect 838 1398 839 1402
rect 843 1398 844 1402
rect 838 1397 844 1398
rect 942 1402 948 1403
rect 942 1398 943 1402
rect 947 1398 948 1402
rect 942 1397 948 1398
rect 1046 1402 1052 1403
rect 1046 1398 1047 1402
rect 1051 1398 1052 1402
rect 1046 1397 1052 1398
rect 1150 1402 1156 1403
rect 1150 1398 1151 1402
rect 1155 1398 1156 1402
rect 1150 1397 1156 1398
rect 1262 1402 1268 1403
rect 1262 1398 1263 1402
rect 1267 1398 1268 1402
rect 1262 1397 1268 1398
rect 202 1394 208 1395
rect 2415 1395 2421 1396
rect 140 1388 190 1390
rect 194 1391 200 1392
rect 140 1387 141 1388
rect 135 1386 141 1387
rect 194 1387 195 1391
rect 199 1390 200 1391
rect 231 1391 237 1392
rect 231 1390 232 1391
rect 199 1388 232 1390
rect 199 1387 200 1388
rect 194 1386 200 1387
rect 231 1387 232 1388
rect 236 1387 237 1391
rect 231 1386 237 1387
rect 359 1391 365 1392
rect 359 1387 360 1391
rect 364 1390 365 1391
rect 426 1391 432 1392
rect 426 1390 427 1391
rect 364 1388 427 1390
rect 364 1387 365 1388
rect 359 1386 365 1387
rect 426 1387 427 1388
rect 431 1387 432 1391
rect 426 1386 432 1387
rect 479 1391 485 1392
rect 479 1387 480 1391
rect 484 1390 485 1391
rect 546 1391 552 1392
rect 546 1390 547 1391
rect 484 1388 547 1390
rect 484 1387 485 1388
rect 479 1386 485 1387
rect 546 1387 547 1388
rect 551 1387 552 1391
rect 546 1386 552 1387
rect 599 1391 605 1392
rect 599 1387 600 1391
rect 604 1390 605 1391
rect 614 1391 620 1392
rect 614 1390 615 1391
rect 604 1388 615 1390
rect 604 1387 605 1388
rect 599 1386 605 1387
rect 614 1387 615 1388
rect 619 1387 620 1391
rect 614 1386 620 1387
rect 719 1391 725 1392
rect 719 1387 720 1391
rect 724 1390 725 1391
rect 786 1391 792 1392
rect 724 1388 782 1390
rect 724 1387 725 1388
rect 719 1386 725 1387
rect 780 1382 782 1388
rect 786 1387 787 1391
rect 791 1390 792 1391
rect 831 1391 837 1392
rect 831 1390 832 1391
rect 791 1388 832 1390
rect 791 1387 792 1388
rect 786 1386 792 1387
rect 831 1387 832 1388
rect 836 1387 837 1391
rect 831 1386 837 1387
rect 898 1391 904 1392
rect 898 1387 899 1391
rect 903 1390 904 1391
rect 935 1391 941 1392
rect 935 1390 936 1391
rect 903 1388 936 1390
rect 903 1387 904 1388
rect 898 1386 904 1387
rect 935 1387 936 1388
rect 940 1387 941 1391
rect 935 1386 941 1387
rect 1002 1391 1008 1392
rect 1002 1387 1003 1391
rect 1007 1390 1008 1391
rect 1039 1391 1045 1392
rect 1039 1390 1040 1391
rect 1007 1388 1040 1390
rect 1007 1387 1008 1388
rect 1002 1386 1008 1387
rect 1039 1387 1040 1388
rect 1044 1387 1045 1391
rect 1039 1386 1045 1387
rect 1106 1391 1112 1392
rect 1106 1387 1107 1391
rect 1111 1390 1112 1391
rect 1143 1391 1149 1392
rect 1143 1390 1144 1391
rect 1111 1388 1144 1390
rect 1111 1387 1112 1388
rect 1106 1386 1112 1387
rect 1143 1387 1144 1388
rect 1148 1387 1149 1391
rect 1143 1386 1149 1387
rect 1210 1391 1216 1392
rect 1210 1387 1211 1391
rect 1215 1390 1216 1391
rect 1255 1391 1261 1392
rect 1255 1390 1256 1391
rect 1215 1388 1256 1390
rect 1215 1387 1216 1388
rect 1210 1386 1216 1387
rect 1255 1387 1256 1388
rect 1260 1387 1261 1391
rect 2415 1391 2416 1395
rect 2420 1394 2421 1395
rect 2511 1395 2517 1396
rect 2511 1394 2512 1395
rect 2420 1392 2512 1394
rect 2420 1391 2421 1392
rect 2415 1390 2421 1391
rect 2511 1391 2512 1392
rect 2516 1391 2517 1395
rect 2511 1390 2517 1391
rect 2606 1395 2612 1396
rect 2606 1391 2607 1395
rect 2611 1394 2612 1395
rect 2615 1395 2621 1396
rect 2615 1394 2616 1395
rect 2611 1392 2616 1394
rect 2611 1391 2612 1392
rect 2606 1390 2612 1391
rect 2615 1391 2616 1392
rect 2620 1391 2621 1395
rect 2615 1390 2621 1391
rect 3414 1395 3420 1396
rect 3414 1391 3415 1395
rect 3419 1394 3420 1395
rect 3487 1395 3493 1396
rect 3487 1394 3488 1395
rect 3419 1392 3488 1394
rect 3419 1391 3420 1392
rect 3414 1390 3420 1391
rect 3487 1391 3488 1392
rect 3492 1391 3493 1395
rect 3487 1390 3493 1391
rect 1255 1386 1261 1387
rect 1174 1383 1180 1384
rect 1174 1382 1175 1383
rect 780 1380 1175 1382
rect 1174 1379 1175 1380
rect 1179 1379 1180 1383
rect 1174 1378 1180 1379
rect 2262 1368 2268 1369
rect 1870 1365 1876 1366
rect 127 1363 133 1364
rect 127 1359 128 1363
rect 132 1362 133 1363
rect 135 1363 141 1364
rect 135 1362 136 1363
rect 132 1360 136 1362
rect 132 1359 133 1360
rect 127 1358 133 1359
rect 135 1359 136 1360
rect 140 1359 141 1363
rect 135 1358 141 1359
rect 279 1363 285 1364
rect 279 1359 280 1363
rect 284 1362 285 1363
rect 298 1363 304 1364
rect 298 1362 299 1363
rect 284 1360 299 1362
rect 284 1359 285 1360
rect 279 1358 285 1359
rect 298 1359 299 1360
rect 303 1359 304 1363
rect 298 1358 304 1359
rect 338 1363 344 1364
rect 338 1359 339 1363
rect 343 1362 344 1363
rect 423 1363 429 1364
rect 423 1362 424 1363
rect 343 1360 424 1362
rect 343 1359 344 1360
rect 338 1358 344 1359
rect 423 1359 424 1360
rect 428 1359 429 1363
rect 423 1358 429 1359
rect 575 1363 581 1364
rect 575 1359 576 1363
rect 580 1362 581 1363
rect 634 1363 640 1364
rect 580 1360 630 1362
rect 580 1359 581 1360
rect 575 1358 581 1359
rect 142 1354 148 1355
rect 142 1350 143 1354
rect 147 1350 148 1354
rect 142 1349 148 1350
rect 286 1354 292 1355
rect 286 1350 287 1354
rect 291 1350 292 1354
rect 286 1349 292 1350
rect 430 1354 436 1355
rect 430 1350 431 1354
rect 435 1350 436 1354
rect 430 1349 436 1350
rect 582 1354 588 1355
rect 582 1350 583 1354
rect 587 1350 588 1354
rect 628 1354 630 1360
rect 634 1359 635 1363
rect 639 1362 640 1363
rect 727 1363 733 1364
rect 727 1362 728 1363
rect 639 1360 728 1362
rect 639 1359 640 1360
rect 634 1358 640 1359
rect 727 1359 728 1360
rect 732 1359 733 1363
rect 727 1358 733 1359
rect 786 1363 792 1364
rect 786 1359 787 1363
rect 791 1362 792 1363
rect 871 1363 877 1364
rect 871 1362 872 1363
rect 791 1360 872 1362
rect 791 1359 792 1360
rect 786 1358 792 1359
rect 871 1359 872 1360
rect 876 1359 877 1363
rect 871 1358 877 1359
rect 930 1363 936 1364
rect 930 1359 931 1363
rect 935 1362 936 1363
rect 1015 1363 1021 1364
rect 1015 1362 1016 1363
rect 935 1360 1016 1362
rect 935 1359 936 1360
rect 930 1358 936 1359
rect 1015 1359 1016 1360
rect 1020 1359 1021 1363
rect 1015 1358 1021 1359
rect 1074 1363 1080 1364
rect 1074 1359 1075 1363
rect 1079 1362 1080 1363
rect 1159 1363 1165 1364
rect 1159 1362 1160 1363
rect 1079 1360 1160 1362
rect 1079 1359 1080 1360
rect 1074 1358 1080 1359
rect 1159 1359 1160 1360
rect 1164 1359 1165 1363
rect 1159 1358 1165 1359
rect 1311 1363 1317 1364
rect 1311 1359 1312 1363
rect 1316 1362 1317 1363
rect 1383 1363 1389 1364
rect 1383 1362 1384 1363
rect 1316 1360 1384 1362
rect 1316 1359 1317 1360
rect 1311 1358 1317 1359
rect 1383 1359 1384 1360
rect 1388 1359 1389 1363
rect 1383 1358 1389 1359
rect 1463 1363 1469 1364
rect 1463 1359 1464 1363
rect 1468 1362 1469 1363
rect 1550 1363 1556 1364
rect 1550 1362 1551 1363
rect 1468 1360 1551 1362
rect 1468 1359 1469 1360
rect 1463 1358 1469 1359
rect 1550 1359 1551 1360
rect 1555 1359 1556 1363
rect 1550 1358 1556 1359
rect 1599 1363 1605 1364
rect 1599 1359 1600 1363
rect 1604 1362 1605 1363
rect 1615 1363 1621 1364
rect 1615 1362 1616 1363
rect 1604 1360 1616 1362
rect 1604 1359 1605 1360
rect 1599 1358 1605 1359
rect 1615 1359 1616 1360
rect 1620 1359 1621 1363
rect 1870 1361 1871 1365
rect 1875 1361 1876 1365
rect 2262 1364 2263 1368
rect 2267 1364 2268 1368
rect 2262 1363 2268 1364
rect 2342 1368 2348 1369
rect 2342 1364 2343 1368
rect 2347 1364 2348 1368
rect 2342 1363 2348 1364
rect 2422 1368 2428 1369
rect 2422 1364 2423 1368
rect 2427 1364 2428 1368
rect 2422 1363 2428 1364
rect 2502 1368 2508 1369
rect 2502 1364 2503 1368
rect 2507 1364 2508 1368
rect 2502 1363 2508 1364
rect 2590 1368 2596 1369
rect 2590 1364 2591 1368
rect 2595 1364 2596 1368
rect 2590 1363 2596 1364
rect 2694 1368 2700 1369
rect 2694 1364 2695 1368
rect 2699 1364 2700 1368
rect 2694 1363 2700 1364
rect 2806 1368 2812 1369
rect 2806 1364 2807 1368
rect 2811 1364 2812 1368
rect 2806 1363 2812 1364
rect 2918 1368 2924 1369
rect 2918 1364 2919 1368
rect 2923 1364 2924 1368
rect 2918 1363 2924 1364
rect 3038 1368 3044 1369
rect 3038 1364 3039 1368
rect 3043 1364 3044 1368
rect 3038 1363 3044 1364
rect 3158 1368 3164 1369
rect 3158 1364 3159 1368
rect 3163 1364 3164 1368
rect 3158 1363 3164 1364
rect 3278 1368 3284 1369
rect 3278 1364 3279 1368
rect 3283 1364 3284 1368
rect 3278 1363 3284 1364
rect 3398 1368 3404 1369
rect 3398 1364 3399 1368
rect 3403 1364 3404 1368
rect 3398 1363 3404 1364
rect 3502 1368 3508 1369
rect 3502 1364 3503 1368
rect 3507 1364 3508 1368
rect 3502 1363 3508 1364
rect 3590 1365 3596 1366
rect 1870 1360 1876 1361
rect 3590 1361 3591 1365
rect 3595 1361 3596 1365
rect 3590 1360 3596 1361
rect 1615 1358 1621 1359
rect 2330 1359 2336 1360
rect 2330 1358 2331 1359
rect 2325 1356 2331 1358
rect 662 1355 668 1356
rect 2330 1355 2331 1356
rect 2335 1355 2336 1359
rect 2414 1359 2420 1360
rect 2414 1358 2415 1359
rect 2405 1356 2415 1358
rect 662 1354 663 1355
rect 628 1352 663 1354
rect 662 1351 663 1352
rect 667 1351 668 1355
rect 662 1350 668 1351
rect 734 1354 740 1355
rect 734 1350 735 1354
rect 739 1350 740 1354
rect 582 1349 588 1350
rect 734 1349 740 1350
rect 878 1354 884 1355
rect 878 1350 879 1354
rect 883 1350 884 1354
rect 878 1349 884 1350
rect 1022 1354 1028 1355
rect 1022 1350 1023 1354
rect 1027 1350 1028 1354
rect 1022 1349 1028 1350
rect 1166 1354 1172 1355
rect 1166 1350 1167 1354
rect 1171 1350 1172 1354
rect 1166 1349 1172 1350
rect 1318 1354 1324 1355
rect 1318 1350 1319 1354
rect 1323 1350 1324 1354
rect 1318 1349 1324 1350
rect 1470 1354 1476 1355
rect 1470 1350 1471 1354
rect 1475 1350 1476 1354
rect 1470 1349 1476 1350
rect 1622 1354 1628 1355
rect 2330 1354 2336 1355
rect 2414 1355 2415 1356
rect 2419 1355 2420 1359
rect 2582 1359 2588 1360
rect 2582 1358 2583 1359
rect 2424 1356 2441 1358
rect 2565 1356 2583 1358
rect 2414 1354 2420 1355
rect 2422 1355 2428 1356
rect 1622 1350 1623 1354
rect 1627 1350 1628 1354
rect 2422 1351 2423 1355
rect 2427 1351 2428 1355
rect 2582 1355 2583 1356
rect 2587 1355 2588 1359
rect 2658 1359 2664 1360
rect 2658 1358 2659 1359
rect 2653 1356 2659 1358
rect 2582 1354 2588 1355
rect 2658 1355 2659 1356
rect 2663 1355 2664 1359
rect 2762 1359 2768 1360
rect 2762 1358 2763 1359
rect 2757 1356 2763 1358
rect 2658 1354 2664 1355
rect 2762 1355 2763 1356
rect 2767 1355 2768 1359
rect 2762 1354 2768 1355
rect 2770 1359 2776 1360
rect 2770 1355 2771 1359
rect 2775 1358 2776 1359
rect 2986 1359 2992 1360
rect 2986 1358 2987 1359
rect 2775 1356 2825 1358
rect 2981 1356 2987 1358
rect 2775 1355 2776 1356
rect 2770 1354 2776 1355
rect 2986 1355 2987 1356
rect 2991 1355 2992 1359
rect 3226 1359 3232 1360
rect 3226 1358 3227 1359
rect 3040 1356 3057 1358
rect 3221 1356 3227 1358
rect 2986 1354 2992 1355
rect 3038 1355 3044 1356
rect 2422 1350 2428 1351
rect 3038 1351 3039 1355
rect 3043 1351 3044 1355
rect 3226 1355 3227 1356
rect 3231 1355 3232 1359
rect 3226 1354 3232 1355
rect 3234 1359 3240 1360
rect 3234 1355 3235 1359
rect 3239 1358 3240 1359
rect 3346 1359 3352 1360
rect 3239 1356 3297 1358
rect 3239 1355 3240 1356
rect 3234 1354 3240 1355
rect 3346 1355 3347 1359
rect 3351 1358 3352 1359
rect 3486 1359 3492 1360
rect 3351 1356 3417 1358
rect 3351 1355 3352 1356
rect 3346 1354 3352 1355
rect 3486 1355 3487 1359
rect 3491 1358 3492 1359
rect 3491 1356 3521 1358
rect 3491 1355 3492 1356
rect 3486 1354 3492 1355
rect 3038 1350 3044 1351
rect 1622 1349 1628 1350
rect 1870 1348 1876 1349
rect 1870 1344 1871 1348
rect 1875 1344 1876 1348
rect 1870 1343 1876 1344
rect 3590 1348 3596 1349
rect 3590 1344 3591 1348
rect 3595 1344 3596 1348
rect 3590 1343 3596 1344
rect 2322 1339 2328 1340
rect 110 1336 116 1337
rect 110 1332 111 1336
rect 115 1332 116 1336
rect 110 1331 116 1332
rect 1830 1336 1836 1337
rect 1830 1332 1831 1336
rect 1835 1332 1836 1336
rect 2322 1335 2323 1339
rect 2327 1338 2328 1339
rect 2770 1339 2776 1340
rect 2770 1338 2771 1339
rect 2327 1336 2771 1338
rect 2327 1335 2328 1336
rect 2322 1334 2328 1335
rect 2770 1335 2771 1336
rect 2775 1335 2776 1339
rect 2770 1334 2776 1335
rect 1830 1331 1836 1332
rect 2270 1330 2276 1331
rect 194 1327 200 1328
rect 194 1323 195 1327
rect 199 1323 200 1327
rect 194 1322 200 1323
rect 338 1327 344 1328
rect 338 1323 339 1327
rect 343 1323 344 1327
rect 338 1322 344 1323
rect 634 1327 640 1328
rect 634 1323 635 1327
rect 639 1323 640 1327
rect 634 1322 640 1323
rect 786 1327 792 1328
rect 786 1323 787 1327
rect 791 1323 792 1327
rect 786 1322 792 1323
rect 930 1327 936 1328
rect 930 1323 931 1327
rect 935 1323 936 1327
rect 930 1322 936 1323
rect 1074 1327 1080 1328
rect 1074 1323 1075 1327
rect 1079 1323 1080 1327
rect 1074 1322 1080 1323
rect 1174 1327 1180 1328
rect 1174 1323 1175 1327
rect 1179 1323 1180 1327
rect 1174 1322 1180 1323
rect 1342 1327 1348 1328
rect 1342 1323 1343 1327
rect 1347 1323 1348 1327
rect 1342 1322 1348 1323
rect 1383 1327 1389 1328
rect 1383 1323 1384 1327
rect 1388 1326 1389 1327
rect 1550 1327 1556 1328
rect 1388 1324 1481 1326
rect 1388 1323 1389 1324
rect 1383 1322 1389 1323
rect 1550 1323 1551 1327
rect 1555 1326 1556 1327
rect 2270 1326 2271 1330
rect 2275 1326 2276 1330
rect 1555 1324 1633 1326
rect 2270 1325 2276 1326
rect 2350 1330 2356 1331
rect 2350 1326 2351 1330
rect 2355 1326 2356 1330
rect 2350 1325 2356 1326
rect 2430 1330 2436 1331
rect 2430 1326 2431 1330
rect 2435 1326 2436 1330
rect 2430 1325 2436 1326
rect 2510 1330 2516 1331
rect 2510 1326 2511 1330
rect 2515 1326 2516 1330
rect 2510 1325 2516 1326
rect 2598 1330 2604 1331
rect 2598 1326 2599 1330
rect 2603 1326 2604 1330
rect 2598 1325 2604 1326
rect 2702 1330 2708 1331
rect 2702 1326 2703 1330
rect 2707 1326 2708 1330
rect 2702 1325 2708 1326
rect 2814 1330 2820 1331
rect 2814 1326 2815 1330
rect 2819 1326 2820 1330
rect 2814 1325 2820 1326
rect 2926 1330 2932 1331
rect 2926 1326 2927 1330
rect 2931 1326 2932 1330
rect 2926 1325 2932 1326
rect 3046 1330 3052 1331
rect 3046 1326 3047 1330
rect 3051 1326 3052 1330
rect 3046 1325 3052 1326
rect 3166 1330 3172 1331
rect 3166 1326 3167 1330
rect 3171 1326 3172 1330
rect 3166 1325 3172 1326
rect 3286 1330 3292 1331
rect 3286 1326 3287 1330
rect 3291 1326 3292 1330
rect 3286 1325 3292 1326
rect 3406 1330 3412 1331
rect 3406 1326 3407 1330
rect 3411 1326 3412 1330
rect 3406 1325 3412 1326
rect 3510 1330 3516 1331
rect 3510 1326 3511 1330
rect 3515 1326 3516 1330
rect 3510 1325 3516 1326
rect 1555 1323 1556 1324
rect 1550 1322 1556 1323
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 1830 1319 1836 1320
rect 110 1314 116 1315
rect 134 1316 140 1317
rect 134 1312 135 1316
rect 139 1312 140 1316
rect 134 1311 140 1312
rect 278 1316 284 1317
rect 278 1312 279 1316
rect 283 1312 284 1316
rect 278 1311 284 1312
rect 422 1316 428 1317
rect 422 1312 423 1316
rect 427 1312 428 1316
rect 422 1311 428 1312
rect 574 1316 580 1317
rect 574 1312 575 1316
rect 579 1312 580 1316
rect 574 1311 580 1312
rect 726 1316 732 1317
rect 726 1312 727 1316
rect 731 1312 732 1316
rect 726 1311 732 1312
rect 870 1316 876 1317
rect 870 1312 871 1316
rect 875 1312 876 1316
rect 870 1311 876 1312
rect 1014 1316 1020 1317
rect 1014 1312 1015 1316
rect 1019 1312 1020 1316
rect 1014 1311 1020 1312
rect 1158 1316 1164 1317
rect 1158 1312 1159 1316
rect 1163 1312 1164 1316
rect 1158 1311 1164 1312
rect 1310 1316 1316 1317
rect 1310 1312 1311 1316
rect 1315 1312 1316 1316
rect 1310 1311 1316 1312
rect 1462 1316 1468 1317
rect 1462 1312 1463 1316
rect 1467 1312 1468 1316
rect 1462 1311 1468 1312
rect 1614 1316 1620 1317
rect 1614 1312 1615 1316
rect 1619 1312 1620 1316
rect 1830 1315 1831 1319
rect 1835 1315 1836 1319
rect 1830 1314 1836 1315
rect 2263 1319 2269 1320
rect 2263 1315 2264 1319
rect 2268 1318 2269 1319
rect 2322 1319 2328 1320
rect 2322 1318 2323 1319
rect 2268 1316 2323 1318
rect 2268 1315 2269 1316
rect 2263 1314 2269 1315
rect 2322 1315 2323 1316
rect 2327 1315 2328 1319
rect 2322 1314 2328 1315
rect 2330 1319 2336 1320
rect 2330 1315 2331 1319
rect 2335 1318 2336 1319
rect 2343 1319 2349 1320
rect 2343 1318 2344 1319
rect 2335 1316 2344 1318
rect 2335 1315 2336 1316
rect 2330 1314 2336 1315
rect 2343 1315 2344 1316
rect 2348 1315 2349 1319
rect 2343 1314 2349 1315
rect 2415 1319 2421 1320
rect 2415 1315 2416 1319
rect 2420 1318 2421 1319
rect 2423 1319 2429 1320
rect 2423 1318 2424 1319
rect 2420 1316 2424 1318
rect 2420 1315 2421 1316
rect 2415 1314 2421 1315
rect 2423 1315 2424 1316
rect 2428 1315 2429 1319
rect 2503 1319 2509 1320
rect 2503 1318 2504 1319
rect 2423 1314 2429 1315
rect 2436 1316 2504 1318
rect 1614 1311 1620 1312
rect 2414 1311 2420 1312
rect 2414 1307 2415 1311
rect 2419 1310 2420 1311
rect 2436 1310 2438 1316
rect 2503 1315 2504 1316
rect 2508 1315 2509 1319
rect 2503 1314 2509 1315
rect 2591 1319 2597 1320
rect 2591 1315 2592 1319
rect 2596 1318 2597 1319
rect 2606 1319 2612 1320
rect 2606 1318 2607 1319
rect 2596 1316 2607 1318
rect 2596 1315 2597 1316
rect 2591 1314 2597 1315
rect 2606 1315 2607 1316
rect 2611 1315 2612 1319
rect 2606 1314 2612 1315
rect 2658 1319 2664 1320
rect 2658 1315 2659 1319
rect 2663 1318 2664 1319
rect 2695 1319 2701 1320
rect 2695 1318 2696 1319
rect 2663 1316 2696 1318
rect 2663 1315 2664 1316
rect 2658 1314 2664 1315
rect 2695 1315 2696 1316
rect 2700 1315 2701 1319
rect 2695 1314 2701 1315
rect 2762 1319 2768 1320
rect 2762 1315 2763 1319
rect 2767 1318 2768 1319
rect 2807 1319 2813 1320
rect 2807 1318 2808 1319
rect 2767 1316 2808 1318
rect 2767 1315 2768 1316
rect 2762 1314 2768 1315
rect 2807 1315 2808 1316
rect 2812 1315 2813 1319
rect 2807 1314 2813 1315
rect 2838 1319 2844 1320
rect 2838 1315 2839 1319
rect 2843 1318 2844 1319
rect 2919 1319 2925 1320
rect 2919 1318 2920 1319
rect 2843 1316 2920 1318
rect 2843 1315 2844 1316
rect 2838 1314 2844 1315
rect 2919 1315 2920 1316
rect 2924 1315 2925 1319
rect 2919 1314 2925 1315
rect 2986 1319 2992 1320
rect 2986 1315 2987 1319
rect 2991 1318 2992 1319
rect 3039 1319 3045 1320
rect 3039 1318 3040 1319
rect 2991 1316 3040 1318
rect 2991 1315 2992 1316
rect 2986 1314 2992 1315
rect 3039 1315 3040 1316
rect 3044 1315 3045 1319
rect 3039 1314 3045 1315
rect 3159 1319 3165 1320
rect 3159 1315 3160 1319
rect 3164 1318 3165 1319
rect 3234 1319 3240 1320
rect 3234 1318 3235 1319
rect 3164 1316 3235 1318
rect 3164 1315 3165 1316
rect 3159 1314 3165 1315
rect 3234 1315 3235 1316
rect 3239 1315 3240 1319
rect 3234 1314 3240 1315
rect 3279 1319 3285 1320
rect 3279 1315 3280 1319
rect 3284 1318 3285 1319
rect 3346 1319 3352 1320
rect 3346 1318 3347 1319
rect 3284 1316 3347 1318
rect 3284 1315 3285 1316
rect 3279 1314 3285 1315
rect 3346 1315 3347 1316
rect 3351 1315 3352 1319
rect 3346 1314 3352 1315
rect 3399 1319 3405 1320
rect 3399 1315 3400 1319
rect 3404 1318 3405 1319
rect 3414 1319 3420 1320
rect 3414 1318 3415 1319
rect 3404 1316 3415 1318
rect 3404 1315 3405 1316
rect 3399 1314 3405 1315
rect 3414 1315 3415 1316
rect 3419 1315 3420 1319
rect 3414 1314 3420 1315
rect 3503 1319 3509 1320
rect 3503 1315 3504 1319
rect 3508 1318 3509 1319
rect 3518 1319 3524 1320
rect 3518 1318 3519 1319
rect 3508 1316 3519 1318
rect 3508 1315 3509 1316
rect 3503 1314 3509 1315
rect 3518 1315 3519 1316
rect 3523 1315 3524 1319
rect 3518 1314 3524 1315
rect 2419 1308 2438 1310
rect 2419 1307 2420 1308
rect 2414 1306 2420 1307
rect 2670 1303 2676 1304
rect 2670 1302 2671 1303
rect 2369 1300 2671 1302
rect 438 1299 445 1300
rect 438 1295 439 1299
rect 444 1295 445 1299
rect 2369 1296 2371 1300
rect 2670 1299 2671 1300
rect 2675 1299 2676 1303
rect 2670 1298 2676 1299
rect 438 1294 445 1295
rect 2207 1295 2213 1296
rect 2207 1291 2208 1295
rect 2212 1294 2213 1295
rect 2278 1295 2284 1296
rect 2278 1294 2279 1295
rect 2212 1292 2279 1294
rect 2212 1291 2213 1292
rect 2207 1290 2213 1291
rect 2278 1291 2279 1292
rect 2283 1291 2284 1295
rect 2278 1290 2284 1291
rect 2287 1295 2293 1296
rect 2287 1291 2288 1295
rect 2292 1294 2293 1295
rect 2358 1295 2364 1296
rect 2358 1294 2359 1295
rect 2292 1292 2359 1294
rect 2292 1291 2293 1292
rect 2287 1290 2293 1291
rect 2358 1291 2359 1292
rect 2363 1291 2364 1295
rect 2358 1290 2364 1291
rect 2367 1295 2373 1296
rect 2367 1291 2368 1295
rect 2372 1291 2373 1295
rect 2367 1290 2373 1291
rect 2422 1295 2428 1296
rect 2422 1291 2423 1295
rect 2427 1294 2428 1295
rect 2447 1295 2453 1296
rect 2447 1294 2448 1295
rect 2427 1292 2448 1294
rect 2427 1291 2428 1292
rect 2422 1290 2428 1291
rect 2447 1291 2448 1292
rect 2452 1291 2453 1295
rect 2447 1290 2453 1291
rect 2519 1295 2525 1296
rect 2519 1291 2520 1295
rect 2524 1294 2525 1295
rect 2543 1295 2549 1296
rect 2543 1294 2544 1295
rect 2524 1292 2544 1294
rect 2524 1291 2525 1292
rect 2519 1290 2525 1291
rect 2543 1291 2544 1292
rect 2548 1291 2549 1295
rect 2543 1290 2549 1291
rect 2654 1295 2661 1296
rect 2654 1291 2655 1295
rect 2660 1291 2661 1295
rect 2654 1290 2661 1291
rect 2783 1295 2789 1296
rect 2783 1291 2784 1295
rect 2788 1294 2789 1295
rect 2850 1295 2856 1296
rect 2850 1294 2851 1295
rect 2788 1292 2851 1294
rect 2788 1291 2789 1292
rect 2783 1290 2789 1291
rect 2850 1291 2851 1292
rect 2855 1291 2856 1295
rect 2850 1290 2856 1291
rect 2919 1295 2925 1296
rect 2919 1291 2920 1295
rect 2924 1294 2925 1295
rect 2998 1295 3004 1296
rect 2998 1294 2999 1295
rect 2924 1292 2999 1294
rect 2924 1291 2925 1292
rect 2919 1290 2925 1291
rect 2998 1291 2999 1292
rect 3003 1291 3004 1295
rect 2998 1290 3004 1291
rect 3038 1295 3044 1296
rect 3038 1291 3039 1295
rect 3043 1294 3044 1295
rect 3063 1295 3069 1296
rect 3063 1294 3064 1295
rect 3043 1292 3064 1294
rect 3043 1291 3044 1292
rect 3038 1290 3044 1291
rect 3063 1291 3064 1292
rect 3068 1291 3069 1295
rect 3063 1290 3069 1291
rect 3207 1295 3213 1296
rect 3207 1291 3208 1295
rect 3212 1294 3213 1295
rect 3226 1295 3232 1296
rect 3226 1294 3227 1295
rect 3212 1292 3227 1294
rect 3212 1291 3213 1292
rect 3207 1290 3213 1291
rect 3226 1291 3227 1292
rect 3231 1291 3232 1295
rect 3226 1290 3232 1291
rect 3266 1295 3272 1296
rect 3266 1291 3267 1295
rect 3271 1294 3272 1295
rect 3359 1295 3365 1296
rect 3359 1294 3360 1295
rect 3271 1292 3360 1294
rect 3271 1291 3272 1292
rect 3266 1290 3272 1291
rect 3359 1291 3360 1292
rect 3364 1291 3365 1295
rect 3359 1290 3365 1291
rect 3487 1295 3493 1296
rect 3487 1291 3488 1295
rect 3492 1294 3493 1295
rect 3503 1295 3509 1296
rect 3503 1294 3504 1295
rect 3492 1292 3504 1294
rect 3492 1291 3493 1292
rect 3487 1290 3493 1291
rect 3503 1291 3504 1292
rect 3508 1291 3509 1295
rect 3503 1290 3509 1291
rect 2214 1286 2220 1287
rect 2214 1282 2215 1286
rect 2219 1282 2220 1286
rect 2214 1281 2220 1282
rect 2294 1286 2300 1287
rect 2294 1282 2295 1286
rect 2299 1282 2300 1286
rect 2294 1281 2300 1282
rect 2374 1286 2380 1287
rect 2374 1282 2375 1286
rect 2379 1282 2380 1286
rect 2374 1281 2380 1282
rect 2454 1286 2460 1287
rect 2454 1282 2455 1286
rect 2459 1282 2460 1286
rect 2454 1281 2460 1282
rect 2550 1286 2556 1287
rect 2550 1282 2551 1286
rect 2555 1282 2556 1286
rect 2550 1281 2556 1282
rect 2662 1286 2668 1287
rect 2662 1282 2663 1286
rect 2667 1282 2668 1286
rect 2662 1281 2668 1282
rect 2790 1286 2796 1287
rect 2790 1282 2791 1286
rect 2795 1282 2796 1286
rect 2790 1281 2796 1282
rect 2926 1286 2932 1287
rect 2926 1282 2927 1286
rect 2931 1282 2932 1286
rect 2926 1281 2932 1282
rect 3070 1286 3076 1287
rect 3070 1282 3071 1286
rect 3075 1282 3076 1286
rect 3070 1281 3076 1282
rect 3214 1286 3220 1287
rect 3214 1282 3215 1286
rect 3219 1282 3220 1286
rect 3214 1281 3220 1282
rect 3366 1286 3372 1287
rect 3366 1282 3367 1286
rect 3371 1282 3372 1286
rect 3366 1281 3372 1282
rect 3510 1286 3516 1287
rect 3510 1282 3511 1286
rect 3515 1282 3516 1286
rect 3510 1281 3516 1282
rect 134 1268 140 1269
rect 110 1265 116 1266
rect 110 1261 111 1265
rect 115 1261 116 1265
rect 134 1264 135 1268
rect 139 1264 140 1268
rect 134 1263 140 1264
rect 262 1268 268 1269
rect 262 1264 263 1268
rect 267 1264 268 1268
rect 262 1263 268 1264
rect 422 1268 428 1269
rect 422 1264 423 1268
rect 427 1264 428 1268
rect 422 1263 428 1264
rect 590 1268 596 1269
rect 590 1264 591 1268
rect 595 1264 596 1268
rect 590 1263 596 1264
rect 758 1268 764 1269
rect 758 1264 759 1268
rect 763 1264 764 1268
rect 758 1263 764 1264
rect 926 1268 932 1269
rect 926 1264 927 1268
rect 931 1264 932 1268
rect 926 1263 932 1264
rect 1078 1268 1084 1269
rect 1078 1264 1079 1268
rect 1083 1264 1084 1268
rect 1078 1263 1084 1264
rect 1222 1268 1228 1269
rect 1222 1264 1223 1268
rect 1227 1264 1228 1268
rect 1222 1263 1228 1264
rect 1350 1268 1356 1269
rect 1350 1264 1351 1268
rect 1355 1264 1356 1268
rect 1350 1263 1356 1264
rect 1478 1268 1484 1269
rect 1478 1264 1479 1268
rect 1483 1264 1484 1268
rect 1478 1263 1484 1264
rect 1606 1268 1612 1269
rect 1606 1264 1607 1268
rect 1611 1264 1612 1268
rect 1606 1263 1612 1264
rect 1734 1268 1740 1269
rect 1734 1264 1735 1268
rect 1739 1264 1740 1268
rect 1870 1268 1876 1269
rect 1734 1263 1740 1264
rect 1830 1265 1836 1266
rect 110 1260 116 1261
rect 1830 1261 1831 1265
rect 1835 1261 1836 1265
rect 1870 1264 1871 1268
rect 1875 1264 1876 1268
rect 1870 1263 1876 1264
rect 3590 1268 3596 1269
rect 3590 1264 3591 1268
rect 3595 1264 3596 1268
rect 3590 1263 3596 1264
rect 1830 1260 1836 1261
rect 127 1259 133 1260
rect 127 1255 128 1259
rect 132 1258 133 1259
rect 207 1259 213 1260
rect 132 1256 153 1258
rect 132 1255 133 1256
rect 127 1254 133 1255
rect 207 1255 208 1259
rect 212 1258 213 1259
rect 498 1259 504 1260
rect 498 1258 499 1259
rect 212 1256 281 1258
rect 485 1256 499 1258
rect 212 1255 213 1256
rect 207 1254 213 1255
rect 498 1255 499 1256
rect 503 1255 504 1259
rect 498 1254 504 1255
rect 506 1259 512 1260
rect 506 1255 507 1259
rect 511 1258 512 1259
rect 662 1259 668 1260
rect 511 1256 609 1258
rect 511 1255 512 1256
rect 506 1254 512 1255
rect 662 1255 663 1259
rect 667 1258 668 1259
rect 826 1259 832 1260
rect 667 1256 777 1258
rect 667 1255 668 1256
rect 662 1254 668 1255
rect 826 1255 827 1259
rect 831 1258 832 1259
rect 1158 1259 1164 1260
rect 1158 1258 1159 1259
rect 831 1256 945 1258
rect 1141 1256 1159 1258
rect 831 1255 832 1256
rect 826 1254 832 1255
rect 1158 1255 1159 1256
rect 1163 1255 1164 1259
rect 1290 1259 1296 1260
rect 1158 1254 1164 1255
rect 1284 1252 1286 1257
rect 1290 1255 1291 1259
rect 1295 1258 1296 1259
rect 1550 1259 1556 1260
rect 1550 1258 1551 1259
rect 1295 1256 1369 1258
rect 1541 1256 1551 1258
rect 1295 1255 1296 1256
rect 1290 1254 1296 1255
rect 1550 1255 1551 1256
rect 1555 1255 1556 1259
rect 1550 1254 1556 1255
rect 1599 1259 1605 1260
rect 1599 1255 1600 1259
rect 1604 1258 1605 1259
rect 2278 1259 2284 1260
rect 1604 1256 1625 1258
rect 1604 1255 1605 1256
rect 1599 1254 1605 1255
rect 1282 1251 1288 1252
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 1282 1247 1283 1251
rect 1287 1247 1288 1251
rect 1282 1246 1288 1247
rect 1538 1251 1544 1252
rect 1538 1247 1539 1251
rect 1543 1250 1544 1251
rect 1752 1250 1754 1257
rect 2278 1255 2279 1259
rect 2283 1258 2284 1259
rect 2358 1259 2364 1260
rect 2283 1256 2305 1258
rect 2283 1255 2284 1256
rect 2278 1254 2284 1255
rect 2358 1255 2359 1259
rect 2363 1258 2364 1259
rect 2519 1259 2525 1260
rect 2519 1258 2520 1259
rect 2363 1256 2385 1258
rect 2509 1256 2520 1258
rect 2363 1255 2364 1256
rect 2358 1254 2364 1255
rect 2519 1255 2520 1256
rect 2524 1255 2525 1259
rect 2654 1259 2660 1260
rect 2654 1258 2655 1259
rect 2605 1256 2655 1258
rect 2519 1254 2525 1255
rect 2654 1255 2655 1256
rect 2659 1255 2660 1259
rect 2654 1254 2660 1255
rect 2670 1259 2676 1260
rect 2670 1255 2671 1259
rect 2675 1255 2676 1259
rect 2670 1254 2676 1255
rect 2850 1259 2856 1260
rect 2850 1255 2851 1259
rect 2855 1258 2856 1259
rect 2998 1259 3004 1260
rect 2855 1256 2937 1258
rect 2855 1255 2856 1256
rect 2850 1254 2856 1255
rect 2998 1255 2999 1259
rect 3003 1258 3004 1259
rect 3266 1259 3272 1260
rect 3003 1256 3081 1258
rect 3003 1255 3004 1256
rect 2998 1254 3004 1255
rect 3266 1255 3267 1259
rect 3271 1255 3272 1259
rect 3266 1254 3272 1255
rect 3518 1259 3524 1260
rect 3518 1255 3519 1259
rect 3523 1255 3524 1259
rect 3518 1254 3524 1255
rect 1543 1248 1754 1250
rect 1870 1251 1876 1252
rect 1830 1248 1836 1249
rect 1543 1247 1544 1248
rect 1538 1246 1544 1247
rect 110 1243 116 1244
rect 1830 1244 1831 1248
rect 1835 1244 1836 1248
rect 1870 1247 1871 1251
rect 1875 1247 1876 1251
rect 3590 1251 3596 1252
rect 1870 1246 1876 1247
rect 2206 1248 2212 1249
rect 1830 1243 1836 1244
rect 2206 1244 2207 1248
rect 2211 1244 2212 1248
rect 2206 1243 2212 1244
rect 2286 1248 2292 1249
rect 2286 1244 2287 1248
rect 2291 1244 2292 1248
rect 2286 1243 2292 1244
rect 2366 1248 2372 1249
rect 2366 1244 2367 1248
rect 2371 1244 2372 1248
rect 2366 1243 2372 1244
rect 2446 1248 2452 1249
rect 2446 1244 2447 1248
rect 2451 1244 2452 1248
rect 2446 1243 2452 1244
rect 2542 1248 2548 1249
rect 2542 1244 2543 1248
rect 2547 1244 2548 1248
rect 2542 1243 2548 1244
rect 2654 1248 2660 1249
rect 2654 1244 2655 1248
rect 2659 1244 2660 1248
rect 2654 1243 2660 1244
rect 2782 1248 2788 1249
rect 2782 1244 2783 1248
rect 2787 1244 2788 1248
rect 2782 1243 2788 1244
rect 2918 1248 2924 1249
rect 2918 1244 2919 1248
rect 2923 1244 2924 1248
rect 2918 1243 2924 1244
rect 3062 1248 3068 1249
rect 3062 1244 3063 1248
rect 3067 1244 3068 1248
rect 3062 1243 3068 1244
rect 3206 1248 3212 1249
rect 3206 1244 3207 1248
rect 3211 1244 3212 1248
rect 3206 1243 3212 1244
rect 3358 1248 3364 1249
rect 3358 1244 3359 1248
rect 3363 1244 3364 1248
rect 3358 1243 3364 1244
rect 3502 1248 3508 1249
rect 3502 1244 3503 1248
rect 3507 1244 3508 1248
rect 3590 1247 3591 1251
rect 3595 1247 3596 1251
rect 3590 1246 3596 1247
rect 3502 1243 3508 1244
rect 2126 1231 2132 1232
rect 142 1230 148 1231
rect 142 1226 143 1230
rect 147 1226 148 1230
rect 270 1230 276 1231
rect 207 1227 213 1228
rect 207 1226 208 1227
rect 142 1225 148 1226
rect 188 1224 208 1226
rect 135 1219 141 1220
rect 135 1215 136 1219
rect 140 1218 141 1219
rect 188 1218 190 1224
rect 207 1223 208 1224
rect 212 1223 213 1227
rect 270 1226 271 1230
rect 275 1226 276 1230
rect 270 1225 276 1226
rect 430 1230 436 1231
rect 430 1226 431 1230
rect 435 1226 436 1230
rect 430 1225 436 1226
rect 598 1230 604 1231
rect 598 1226 599 1230
rect 603 1226 604 1230
rect 598 1225 604 1226
rect 766 1230 772 1231
rect 766 1226 767 1230
rect 771 1226 772 1230
rect 766 1225 772 1226
rect 934 1230 940 1231
rect 934 1226 935 1230
rect 939 1226 940 1230
rect 934 1225 940 1226
rect 1086 1230 1092 1231
rect 1086 1226 1087 1230
rect 1091 1226 1092 1230
rect 1086 1225 1092 1226
rect 1230 1230 1236 1231
rect 1230 1226 1231 1230
rect 1235 1226 1236 1230
rect 1230 1225 1236 1226
rect 1358 1230 1364 1231
rect 1358 1226 1359 1230
rect 1363 1226 1364 1230
rect 1358 1225 1364 1226
rect 1486 1230 1492 1231
rect 1486 1226 1487 1230
rect 1491 1226 1492 1230
rect 1486 1225 1492 1226
rect 1614 1230 1620 1231
rect 1614 1226 1615 1230
rect 1619 1226 1620 1230
rect 1614 1225 1620 1226
rect 1742 1230 1748 1231
rect 1742 1226 1743 1230
rect 1747 1226 1748 1230
rect 2126 1227 2127 1231
rect 2131 1230 2132 1231
rect 2223 1231 2229 1232
rect 2223 1230 2224 1231
rect 2131 1228 2224 1230
rect 2131 1227 2132 1228
rect 2126 1226 2132 1227
rect 2223 1227 2224 1228
rect 2228 1227 2229 1231
rect 2223 1226 2229 1227
rect 2662 1231 2668 1232
rect 2662 1227 2663 1231
rect 2667 1230 2668 1231
rect 2799 1231 2805 1232
rect 2799 1230 2800 1231
rect 2667 1228 2800 1230
rect 2667 1227 2668 1228
rect 2662 1226 2668 1227
rect 2799 1227 2800 1228
rect 2804 1227 2805 1231
rect 2799 1226 2805 1227
rect 3366 1231 3372 1232
rect 3366 1227 3367 1231
rect 3371 1230 3372 1231
rect 3375 1231 3381 1232
rect 3375 1230 3376 1231
rect 3371 1228 3376 1230
rect 3371 1227 3372 1228
rect 3366 1226 3372 1227
rect 3375 1227 3376 1228
rect 3380 1227 3381 1231
rect 3375 1226 3381 1227
rect 1742 1225 1748 1226
rect 207 1222 213 1223
rect 140 1216 190 1218
rect 194 1219 200 1220
rect 140 1215 141 1216
rect 135 1214 141 1215
rect 194 1215 195 1219
rect 199 1218 200 1219
rect 263 1219 269 1220
rect 263 1218 264 1219
rect 199 1216 264 1218
rect 199 1215 200 1216
rect 194 1214 200 1215
rect 263 1215 264 1216
rect 268 1215 269 1219
rect 263 1214 269 1215
rect 423 1219 429 1220
rect 423 1215 424 1219
rect 428 1218 429 1219
rect 438 1219 444 1220
rect 438 1218 439 1219
rect 428 1216 439 1218
rect 428 1215 429 1216
rect 423 1214 429 1215
rect 438 1215 439 1216
rect 443 1215 444 1219
rect 438 1214 444 1215
rect 498 1219 504 1220
rect 498 1215 499 1219
rect 503 1218 504 1219
rect 591 1219 597 1220
rect 591 1218 592 1219
rect 503 1216 592 1218
rect 503 1215 504 1216
rect 498 1214 504 1215
rect 591 1215 592 1216
rect 596 1215 597 1219
rect 591 1214 597 1215
rect 759 1219 765 1220
rect 759 1215 760 1219
rect 764 1218 765 1219
rect 826 1219 832 1220
rect 826 1218 827 1219
rect 764 1216 827 1218
rect 764 1215 765 1216
rect 759 1214 765 1215
rect 826 1215 827 1216
rect 831 1215 832 1219
rect 826 1214 832 1215
rect 898 1219 904 1220
rect 898 1215 899 1219
rect 903 1218 904 1219
rect 927 1219 933 1220
rect 927 1218 928 1219
rect 903 1216 928 1218
rect 903 1215 904 1216
rect 898 1214 904 1215
rect 927 1215 928 1216
rect 932 1215 933 1219
rect 927 1214 933 1215
rect 1079 1219 1085 1220
rect 1079 1215 1080 1219
rect 1084 1218 1085 1219
rect 1094 1219 1100 1220
rect 1094 1218 1095 1219
rect 1084 1216 1095 1218
rect 1084 1215 1085 1216
rect 1079 1214 1085 1215
rect 1094 1215 1095 1216
rect 1099 1215 1100 1219
rect 1094 1214 1100 1215
rect 1158 1219 1164 1220
rect 1158 1215 1159 1219
rect 1163 1218 1164 1219
rect 1223 1219 1229 1220
rect 1223 1218 1224 1219
rect 1163 1216 1224 1218
rect 1163 1215 1164 1216
rect 1158 1214 1164 1215
rect 1223 1215 1224 1216
rect 1228 1215 1229 1219
rect 1223 1214 1229 1215
rect 1342 1219 1348 1220
rect 1342 1215 1343 1219
rect 1347 1218 1348 1219
rect 1351 1219 1357 1220
rect 1351 1218 1352 1219
rect 1347 1216 1352 1218
rect 1347 1215 1348 1216
rect 1342 1214 1348 1215
rect 1351 1215 1352 1216
rect 1356 1215 1357 1219
rect 1351 1214 1357 1215
rect 1479 1219 1485 1220
rect 1479 1215 1480 1219
rect 1484 1218 1485 1219
rect 1538 1219 1544 1220
rect 1538 1218 1539 1219
rect 1484 1216 1539 1218
rect 1484 1215 1485 1216
rect 1479 1214 1485 1215
rect 1538 1215 1539 1216
rect 1543 1215 1544 1219
rect 1538 1214 1544 1215
rect 1550 1219 1556 1220
rect 1550 1215 1551 1219
rect 1555 1218 1556 1219
rect 1607 1219 1613 1220
rect 1607 1218 1608 1219
rect 1555 1216 1608 1218
rect 1555 1215 1556 1216
rect 1550 1214 1556 1215
rect 1607 1215 1608 1216
rect 1612 1215 1613 1219
rect 1607 1214 1613 1215
rect 1735 1219 1741 1220
rect 1735 1215 1736 1219
rect 1740 1218 1741 1219
rect 1758 1219 1764 1220
rect 1758 1218 1759 1219
rect 1740 1216 1759 1218
rect 1740 1215 1741 1216
rect 1735 1214 1741 1215
rect 1758 1215 1759 1216
rect 1763 1215 1764 1219
rect 1758 1214 1764 1215
rect 1302 1207 1308 1208
rect 1302 1206 1303 1207
rect 1052 1204 1303 1206
rect 127 1199 133 1200
rect 127 1195 128 1199
rect 132 1198 133 1199
rect 135 1199 141 1200
rect 135 1198 136 1199
rect 132 1196 136 1198
rect 132 1195 133 1196
rect 127 1194 133 1195
rect 135 1195 136 1196
rect 140 1195 141 1199
rect 135 1194 141 1195
rect 303 1199 309 1200
rect 303 1195 304 1199
rect 308 1198 309 1199
rect 422 1199 428 1200
rect 422 1198 423 1199
rect 308 1196 423 1198
rect 308 1195 309 1196
rect 303 1194 309 1195
rect 422 1195 423 1196
rect 427 1195 428 1199
rect 422 1194 428 1195
rect 479 1199 485 1200
rect 479 1195 480 1199
rect 484 1198 485 1199
rect 506 1199 512 1200
rect 506 1198 507 1199
rect 484 1196 507 1198
rect 484 1195 485 1196
rect 479 1194 485 1195
rect 506 1195 507 1196
rect 511 1195 512 1199
rect 506 1194 512 1195
rect 538 1199 544 1200
rect 538 1195 539 1199
rect 543 1198 544 1199
rect 663 1199 669 1200
rect 663 1198 664 1199
rect 543 1196 664 1198
rect 543 1195 544 1196
rect 538 1194 544 1195
rect 663 1195 664 1196
rect 668 1195 669 1199
rect 663 1194 669 1195
rect 839 1199 845 1200
rect 839 1195 840 1199
rect 844 1198 845 1199
rect 854 1199 860 1200
rect 854 1198 855 1199
rect 844 1196 855 1198
rect 844 1195 845 1196
rect 839 1194 845 1195
rect 854 1195 855 1196
rect 859 1195 860 1199
rect 854 1194 860 1195
rect 999 1199 1005 1200
rect 999 1195 1000 1199
rect 1004 1198 1005 1199
rect 1052 1198 1054 1204
rect 1302 1203 1303 1204
rect 1307 1203 1308 1207
rect 1570 1207 1576 1208
rect 1570 1206 1571 1207
rect 1302 1202 1308 1203
rect 1459 1204 1571 1206
rect 1004 1196 1054 1198
rect 1058 1199 1064 1200
rect 1004 1195 1005 1196
rect 999 1194 1005 1195
rect 1058 1195 1059 1199
rect 1063 1198 1064 1199
rect 1151 1199 1157 1200
rect 1151 1198 1152 1199
rect 1063 1196 1152 1198
rect 1063 1195 1064 1196
rect 1058 1194 1064 1195
rect 1151 1195 1152 1196
rect 1156 1195 1157 1199
rect 1151 1194 1157 1195
rect 1282 1199 1293 1200
rect 1282 1195 1283 1199
rect 1287 1195 1288 1199
rect 1292 1195 1293 1199
rect 1282 1194 1293 1195
rect 1407 1199 1413 1200
rect 1407 1195 1408 1199
rect 1412 1198 1413 1199
rect 1459 1198 1461 1204
rect 1570 1203 1571 1204
rect 1575 1203 1576 1207
rect 1570 1202 1576 1203
rect 2110 1200 2116 1201
rect 1412 1196 1461 1198
rect 1466 1199 1472 1200
rect 1412 1195 1413 1196
rect 1407 1194 1413 1195
rect 1466 1195 1467 1199
rect 1471 1198 1472 1199
rect 1527 1199 1533 1200
rect 1527 1198 1528 1199
rect 1471 1196 1528 1198
rect 1471 1195 1472 1196
rect 1466 1194 1472 1195
rect 1527 1195 1528 1196
rect 1532 1195 1533 1199
rect 1527 1194 1533 1195
rect 1586 1199 1592 1200
rect 1586 1195 1587 1199
rect 1591 1198 1592 1199
rect 1647 1199 1653 1200
rect 1647 1198 1648 1199
rect 1591 1196 1648 1198
rect 1591 1195 1592 1196
rect 1586 1194 1592 1195
rect 1647 1195 1648 1196
rect 1652 1195 1653 1199
rect 1647 1194 1653 1195
rect 1706 1199 1712 1200
rect 1706 1195 1707 1199
rect 1711 1198 1712 1199
rect 1743 1199 1749 1200
rect 1743 1198 1744 1199
rect 1711 1196 1744 1198
rect 1711 1195 1712 1196
rect 1706 1194 1712 1195
rect 1743 1195 1744 1196
rect 1748 1195 1749 1199
rect 1743 1194 1749 1195
rect 1870 1197 1876 1198
rect 1870 1193 1871 1197
rect 1875 1193 1876 1197
rect 2110 1196 2111 1200
rect 2115 1196 2116 1200
rect 2110 1195 2116 1196
rect 2206 1200 2212 1201
rect 2206 1196 2207 1200
rect 2211 1196 2212 1200
rect 2206 1195 2212 1196
rect 2302 1200 2308 1201
rect 2302 1196 2303 1200
rect 2307 1196 2308 1200
rect 2302 1195 2308 1196
rect 2406 1200 2412 1201
rect 2406 1196 2407 1200
rect 2411 1196 2412 1200
rect 2406 1195 2412 1196
rect 2526 1200 2532 1201
rect 2526 1196 2527 1200
rect 2531 1196 2532 1200
rect 2526 1195 2532 1196
rect 2646 1200 2652 1201
rect 2646 1196 2647 1200
rect 2651 1196 2652 1200
rect 2646 1195 2652 1196
rect 2774 1200 2780 1201
rect 2774 1196 2775 1200
rect 2779 1196 2780 1200
rect 2774 1195 2780 1196
rect 2910 1200 2916 1201
rect 2910 1196 2911 1200
rect 2915 1196 2916 1200
rect 2910 1195 2916 1196
rect 3054 1200 3060 1201
rect 3054 1196 3055 1200
rect 3059 1196 3060 1200
rect 3054 1195 3060 1196
rect 3198 1200 3204 1201
rect 3198 1196 3199 1200
rect 3203 1196 3204 1200
rect 3198 1195 3204 1196
rect 3342 1200 3348 1201
rect 3342 1196 3343 1200
rect 3347 1196 3348 1200
rect 3342 1195 3348 1196
rect 3494 1200 3500 1201
rect 3494 1196 3495 1200
rect 3499 1196 3500 1200
rect 3494 1195 3500 1196
rect 3590 1197 3596 1198
rect 1870 1192 1876 1193
rect 3590 1193 3591 1197
rect 3595 1193 3596 1197
rect 3590 1192 3596 1193
rect 2178 1191 2184 1192
rect 142 1190 148 1191
rect 142 1186 143 1190
rect 147 1186 148 1190
rect 142 1185 148 1186
rect 310 1190 316 1191
rect 310 1186 311 1190
rect 315 1186 316 1190
rect 310 1185 316 1186
rect 486 1190 492 1191
rect 486 1186 487 1190
rect 491 1186 492 1190
rect 486 1185 492 1186
rect 670 1190 676 1191
rect 670 1186 671 1190
rect 675 1186 676 1190
rect 670 1185 676 1186
rect 846 1190 852 1191
rect 846 1186 847 1190
rect 851 1186 852 1190
rect 846 1185 852 1186
rect 1006 1190 1012 1191
rect 1006 1186 1007 1190
rect 1011 1186 1012 1190
rect 1006 1185 1012 1186
rect 1158 1190 1164 1191
rect 1158 1186 1159 1190
rect 1163 1186 1164 1190
rect 1158 1185 1164 1186
rect 1294 1190 1300 1191
rect 1294 1186 1295 1190
rect 1299 1186 1300 1190
rect 1294 1185 1300 1186
rect 1414 1190 1420 1191
rect 1414 1186 1415 1190
rect 1419 1186 1420 1190
rect 1414 1185 1420 1186
rect 1534 1190 1540 1191
rect 1534 1186 1535 1190
rect 1539 1186 1540 1190
rect 1534 1185 1540 1186
rect 1654 1190 1660 1191
rect 1654 1186 1655 1190
rect 1659 1186 1660 1190
rect 1654 1185 1660 1186
rect 1750 1190 1756 1191
rect 2178 1190 2179 1191
rect 1750 1186 1751 1190
rect 1755 1186 1756 1190
rect 2173 1188 2179 1190
rect 2178 1187 2179 1188
rect 2183 1187 2184 1191
rect 2274 1191 2280 1192
rect 2274 1190 2275 1191
rect 2269 1188 2275 1190
rect 2178 1186 2184 1187
rect 2274 1187 2275 1188
rect 2279 1187 2280 1191
rect 2370 1191 2376 1192
rect 2370 1190 2371 1191
rect 2365 1188 2371 1190
rect 2274 1186 2280 1187
rect 2370 1187 2371 1188
rect 2375 1187 2376 1191
rect 2474 1191 2480 1192
rect 2474 1190 2475 1191
rect 2469 1188 2475 1190
rect 2370 1186 2376 1187
rect 2474 1187 2475 1188
rect 2479 1187 2480 1191
rect 2474 1186 2480 1187
rect 2482 1191 2488 1192
rect 2482 1187 2483 1191
rect 2487 1190 2488 1191
rect 2718 1191 2724 1192
rect 2718 1190 2719 1191
rect 2487 1188 2545 1190
rect 2709 1188 2719 1190
rect 2487 1187 2488 1188
rect 2482 1186 2488 1187
rect 2718 1187 2719 1188
rect 2723 1187 2724 1191
rect 2850 1191 2856 1192
rect 2850 1190 2851 1191
rect 2837 1188 2851 1190
rect 2718 1186 2724 1187
rect 2850 1187 2851 1188
rect 2855 1187 2856 1191
rect 2990 1191 2996 1192
rect 2990 1190 2991 1191
rect 2973 1188 2991 1190
rect 2850 1186 2856 1187
rect 2990 1187 2991 1188
rect 2995 1187 2996 1191
rect 2990 1186 2996 1187
rect 2998 1191 3004 1192
rect 2998 1187 2999 1191
rect 3003 1190 3004 1191
rect 3274 1191 3280 1192
rect 3274 1190 3275 1191
rect 3003 1188 3073 1190
rect 3261 1188 3275 1190
rect 3003 1187 3004 1188
rect 2998 1186 3004 1187
rect 3274 1187 3275 1188
rect 3279 1187 3280 1191
rect 3274 1186 3280 1187
rect 3282 1191 3288 1192
rect 3282 1187 3283 1191
rect 3287 1190 3288 1191
rect 3487 1191 3493 1192
rect 3287 1188 3361 1190
rect 3287 1187 3288 1188
rect 3282 1186 3288 1187
rect 3487 1187 3488 1191
rect 3492 1190 3493 1191
rect 3492 1188 3513 1190
rect 3492 1187 3493 1188
rect 3487 1186 3493 1187
rect 1750 1185 1756 1186
rect 1870 1180 1876 1181
rect 1870 1176 1871 1180
rect 1875 1176 1876 1180
rect 1870 1175 1876 1176
rect 3590 1180 3596 1181
rect 3590 1176 3591 1180
rect 3595 1176 3596 1180
rect 3590 1175 3596 1176
rect 110 1172 116 1173
rect 110 1168 111 1172
rect 115 1168 116 1172
rect 110 1167 116 1168
rect 1830 1172 1836 1173
rect 1830 1168 1831 1172
rect 1835 1168 1836 1172
rect 1830 1167 1836 1168
rect 194 1163 200 1164
rect 194 1159 195 1163
rect 199 1159 200 1163
rect 194 1158 200 1159
rect 538 1163 544 1164
rect 538 1159 539 1163
rect 543 1159 544 1163
rect 538 1158 544 1159
rect 678 1163 684 1164
rect 678 1159 679 1163
rect 683 1159 684 1163
rect 678 1158 684 1159
rect 898 1163 904 1164
rect 898 1159 899 1163
rect 903 1159 904 1163
rect 898 1158 904 1159
rect 1058 1163 1064 1164
rect 1058 1159 1059 1163
rect 1063 1159 1064 1163
rect 1058 1158 1064 1159
rect 1210 1163 1216 1164
rect 1210 1159 1211 1163
rect 1215 1159 1216 1163
rect 1210 1158 1216 1159
rect 1302 1163 1308 1164
rect 1302 1159 1303 1163
rect 1307 1159 1308 1163
rect 1302 1158 1308 1159
rect 1466 1163 1472 1164
rect 1466 1159 1467 1163
rect 1471 1159 1472 1163
rect 1466 1158 1472 1159
rect 1586 1163 1592 1164
rect 1586 1159 1587 1163
rect 1591 1159 1592 1163
rect 1586 1158 1592 1159
rect 1706 1163 1712 1164
rect 1706 1159 1707 1163
rect 1711 1159 1712 1163
rect 1706 1158 1712 1159
rect 1758 1163 1764 1164
rect 1758 1159 1759 1163
rect 1763 1159 1764 1163
rect 1758 1158 1764 1159
rect 2118 1162 2124 1163
rect 2118 1158 2119 1162
rect 2123 1158 2124 1162
rect 2118 1157 2124 1158
rect 2214 1162 2220 1163
rect 2214 1158 2215 1162
rect 2219 1158 2220 1162
rect 2214 1157 2220 1158
rect 2310 1162 2316 1163
rect 2310 1158 2311 1162
rect 2315 1158 2316 1162
rect 2310 1157 2316 1158
rect 2414 1162 2420 1163
rect 2414 1158 2415 1162
rect 2419 1158 2420 1162
rect 2414 1157 2420 1158
rect 2534 1162 2540 1163
rect 2534 1158 2535 1162
rect 2539 1158 2540 1162
rect 2534 1157 2540 1158
rect 2654 1162 2660 1163
rect 2654 1158 2655 1162
rect 2659 1158 2660 1162
rect 2654 1157 2660 1158
rect 2782 1162 2788 1163
rect 2782 1158 2783 1162
rect 2787 1158 2788 1162
rect 2782 1157 2788 1158
rect 2918 1162 2924 1163
rect 2918 1158 2919 1162
rect 2923 1158 2924 1162
rect 2918 1157 2924 1158
rect 3062 1162 3068 1163
rect 3062 1158 3063 1162
rect 3067 1158 3068 1162
rect 3062 1157 3068 1158
rect 3206 1162 3212 1163
rect 3206 1158 3207 1162
rect 3211 1158 3212 1162
rect 3206 1157 3212 1158
rect 3350 1162 3356 1163
rect 3350 1158 3351 1162
rect 3355 1158 3356 1162
rect 3350 1157 3356 1158
rect 3502 1162 3508 1163
rect 3502 1158 3503 1162
rect 3507 1158 3508 1162
rect 3502 1157 3508 1158
rect 110 1155 116 1156
rect 110 1151 111 1155
rect 115 1151 116 1155
rect 1830 1155 1836 1156
rect 110 1150 116 1151
rect 134 1152 140 1153
rect 134 1148 135 1152
rect 139 1148 140 1152
rect 134 1147 140 1148
rect 302 1152 308 1153
rect 302 1148 303 1152
rect 307 1148 308 1152
rect 302 1147 308 1148
rect 478 1152 484 1153
rect 478 1148 479 1152
rect 483 1148 484 1152
rect 478 1147 484 1148
rect 662 1152 668 1153
rect 662 1148 663 1152
rect 667 1148 668 1152
rect 662 1147 668 1148
rect 838 1152 844 1153
rect 838 1148 839 1152
rect 843 1148 844 1152
rect 838 1147 844 1148
rect 998 1152 1004 1153
rect 998 1148 999 1152
rect 1003 1148 1004 1152
rect 998 1147 1004 1148
rect 1150 1152 1156 1153
rect 1150 1148 1151 1152
rect 1155 1148 1156 1152
rect 1150 1147 1156 1148
rect 1286 1152 1292 1153
rect 1286 1148 1287 1152
rect 1291 1148 1292 1152
rect 1286 1147 1292 1148
rect 1406 1152 1412 1153
rect 1406 1148 1407 1152
rect 1411 1148 1412 1152
rect 1406 1147 1412 1148
rect 1526 1152 1532 1153
rect 1526 1148 1527 1152
rect 1531 1148 1532 1152
rect 1526 1147 1532 1148
rect 1646 1152 1652 1153
rect 1646 1148 1647 1152
rect 1651 1148 1652 1152
rect 1646 1147 1652 1148
rect 1742 1152 1748 1153
rect 1742 1148 1743 1152
rect 1747 1148 1748 1152
rect 1830 1151 1831 1155
rect 1835 1151 1836 1155
rect 1830 1150 1836 1151
rect 2111 1151 2117 1152
rect 1742 1147 1748 1148
rect 2111 1147 2112 1151
rect 2116 1150 2117 1151
rect 2126 1151 2132 1152
rect 2126 1150 2127 1151
rect 2116 1148 2127 1150
rect 2116 1147 2117 1148
rect 2111 1146 2117 1147
rect 2126 1147 2127 1148
rect 2131 1147 2132 1151
rect 2126 1146 2132 1147
rect 2178 1151 2184 1152
rect 2178 1147 2179 1151
rect 2183 1150 2184 1151
rect 2207 1151 2213 1152
rect 2207 1150 2208 1151
rect 2183 1148 2208 1150
rect 2183 1147 2184 1148
rect 2178 1146 2184 1147
rect 2207 1147 2208 1148
rect 2212 1147 2213 1151
rect 2207 1146 2213 1147
rect 2274 1151 2280 1152
rect 2274 1147 2275 1151
rect 2279 1150 2280 1151
rect 2303 1151 2309 1152
rect 2303 1150 2304 1151
rect 2279 1148 2304 1150
rect 2279 1147 2280 1148
rect 2274 1146 2280 1147
rect 2303 1147 2304 1148
rect 2308 1147 2309 1151
rect 2303 1146 2309 1147
rect 2370 1151 2376 1152
rect 2370 1147 2371 1151
rect 2375 1150 2376 1151
rect 2407 1151 2413 1152
rect 2407 1150 2408 1151
rect 2375 1148 2408 1150
rect 2375 1147 2376 1148
rect 2370 1146 2376 1147
rect 2407 1147 2408 1148
rect 2412 1147 2413 1151
rect 2407 1146 2413 1147
rect 2474 1151 2480 1152
rect 2474 1147 2475 1151
rect 2479 1150 2480 1151
rect 2527 1151 2533 1152
rect 2527 1150 2528 1151
rect 2479 1148 2528 1150
rect 2479 1147 2480 1148
rect 2474 1146 2480 1147
rect 2527 1147 2528 1148
rect 2532 1147 2533 1151
rect 2527 1146 2533 1147
rect 2647 1151 2653 1152
rect 2647 1147 2648 1151
rect 2652 1150 2653 1151
rect 2662 1151 2668 1152
rect 2662 1150 2663 1151
rect 2652 1148 2663 1150
rect 2652 1147 2653 1148
rect 2647 1146 2653 1147
rect 2662 1147 2663 1148
rect 2667 1147 2668 1151
rect 2662 1146 2668 1147
rect 2718 1151 2724 1152
rect 2718 1147 2719 1151
rect 2723 1150 2724 1151
rect 2775 1151 2781 1152
rect 2775 1150 2776 1151
rect 2723 1148 2776 1150
rect 2723 1147 2724 1148
rect 2718 1146 2724 1147
rect 2775 1147 2776 1148
rect 2780 1147 2781 1151
rect 2775 1146 2781 1147
rect 2850 1151 2856 1152
rect 2850 1147 2851 1151
rect 2855 1150 2856 1151
rect 2911 1151 2917 1152
rect 2911 1150 2912 1151
rect 2855 1148 2912 1150
rect 2855 1147 2856 1148
rect 2850 1146 2856 1147
rect 2911 1147 2912 1148
rect 2916 1147 2917 1151
rect 2911 1146 2917 1147
rect 2990 1151 2996 1152
rect 2990 1147 2991 1151
rect 2995 1150 2996 1151
rect 3055 1151 3061 1152
rect 3055 1150 3056 1151
rect 2995 1148 3056 1150
rect 2995 1147 2996 1148
rect 2990 1146 2996 1147
rect 3055 1147 3056 1148
rect 3060 1147 3061 1151
rect 3055 1146 3061 1147
rect 3199 1151 3205 1152
rect 3199 1147 3200 1151
rect 3204 1150 3205 1151
rect 3282 1151 3288 1152
rect 3282 1150 3283 1151
rect 3204 1148 3283 1150
rect 3204 1147 3205 1148
rect 3199 1146 3205 1147
rect 3282 1147 3283 1148
rect 3287 1147 3288 1151
rect 3282 1146 3288 1147
rect 3343 1151 3349 1152
rect 3343 1147 3344 1151
rect 3348 1150 3349 1151
rect 3366 1151 3372 1152
rect 3366 1150 3367 1151
rect 3348 1148 3367 1150
rect 3348 1147 3349 1148
rect 3343 1146 3349 1147
rect 3366 1147 3367 1148
rect 3371 1147 3372 1151
rect 3366 1146 3372 1147
rect 3495 1151 3501 1152
rect 3495 1147 3496 1151
rect 3500 1150 3501 1151
rect 3518 1151 3524 1152
rect 3518 1150 3519 1151
rect 3500 1148 3519 1150
rect 3500 1147 3501 1148
rect 3495 1146 3501 1147
rect 3518 1147 3519 1148
rect 3523 1147 3524 1151
rect 3518 1146 3524 1147
rect 262 1135 268 1136
rect 262 1131 263 1135
rect 267 1134 268 1135
rect 319 1135 325 1136
rect 319 1134 320 1135
rect 267 1132 320 1134
rect 267 1131 268 1132
rect 262 1130 268 1131
rect 319 1131 320 1132
rect 324 1131 325 1135
rect 319 1130 325 1131
rect 1887 1131 1893 1132
rect 1887 1127 1888 1131
rect 1892 1130 1893 1131
rect 1895 1131 1901 1132
rect 1895 1130 1896 1131
rect 1892 1128 1896 1130
rect 1892 1127 1893 1128
rect 1887 1126 1893 1127
rect 1895 1127 1896 1128
rect 1900 1127 1901 1131
rect 1895 1126 1901 1127
rect 2119 1131 2125 1132
rect 2119 1127 2120 1131
rect 2124 1130 2125 1131
rect 2263 1131 2269 1132
rect 2263 1130 2264 1131
rect 2124 1128 2264 1130
rect 2124 1127 2125 1128
rect 2119 1126 2125 1127
rect 2263 1127 2264 1128
rect 2268 1127 2269 1131
rect 2263 1126 2269 1127
rect 2351 1131 2357 1132
rect 2351 1127 2352 1131
rect 2356 1130 2357 1131
rect 2482 1131 2488 1132
rect 2482 1130 2483 1131
rect 2356 1128 2483 1130
rect 2356 1127 2357 1128
rect 2351 1126 2357 1127
rect 2482 1127 2483 1128
rect 2487 1127 2488 1131
rect 2482 1126 2488 1127
rect 2567 1131 2573 1132
rect 2567 1127 2568 1131
rect 2572 1130 2573 1131
rect 2582 1131 2588 1132
rect 2582 1130 2583 1131
rect 2572 1128 2583 1130
rect 2572 1127 2573 1128
rect 2567 1126 2573 1127
rect 2582 1127 2583 1128
rect 2587 1127 2588 1131
rect 2582 1126 2588 1127
rect 2626 1131 2632 1132
rect 2626 1127 2627 1131
rect 2631 1130 2632 1131
rect 2767 1131 2773 1132
rect 2767 1130 2768 1131
rect 2631 1128 2768 1130
rect 2631 1127 2632 1128
rect 2626 1126 2632 1127
rect 2767 1127 2768 1128
rect 2772 1127 2773 1131
rect 2767 1126 2773 1127
rect 2826 1131 2832 1132
rect 2826 1127 2827 1131
rect 2831 1130 2832 1131
rect 2959 1131 2965 1132
rect 2959 1130 2960 1131
rect 2831 1128 2960 1130
rect 2831 1127 2832 1128
rect 2826 1126 2832 1127
rect 2959 1127 2960 1128
rect 2964 1127 2965 1131
rect 2959 1126 2965 1127
rect 3151 1131 3157 1132
rect 3151 1127 3152 1131
rect 3156 1130 3157 1131
rect 3254 1131 3260 1132
rect 3254 1130 3255 1131
rect 3156 1128 3255 1130
rect 3156 1127 3157 1128
rect 3151 1126 3157 1127
rect 3254 1127 3255 1128
rect 3259 1127 3260 1131
rect 3254 1126 3260 1127
rect 3274 1131 3280 1132
rect 3274 1127 3275 1131
rect 3279 1130 3280 1131
rect 3335 1131 3341 1132
rect 3335 1130 3336 1131
rect 3279 1128 3336 1130
rect 3279 1127 3280 1128
rect 3274 1126 3280 1127
rect 3335 1127 3336 1128
rect 3340 1127 3341 1131
rect 3335 1126 3341 1127
rect 3495 1131 3501 1132
rect 3495 1127 3496 1131
rect 3500 1130 3501 1131
rect 3503 1131 3509 1132
rect 3503 1130 3504 1131
rect 3500 1128 3504 1130
rect 3500 1127 3501 1128
rect 3495 1126 3501 1127
rect 3503 1127 3504 1128
rect 3508 1127 3509 1131
rect 3503 1126 3509 1127
rect 1902 1122 1908 1123
rect 1902 1118 1903 1122
rect 1907 1118 1908 1122
rect 1902 1117 1908 1118
rect 2126 1122 2132 1123
rect 2126 1118 2127 1122
rect 2131 1118 2132 1122
rect 2126 1117 2132 1118
rect 2358 1122 2364 1123
rect 2358 1118 2359 1122
rect 2363 1118 2364 1122
rect 2358 1117 2364 1118
rect 2574 1122 2580 1123
rect 2574 1118 2575 1122
rect 2579 1118 2580 1122
rect 2574 1117 2580 1118
rect 2774 1122 2780 1123
rect 2774 1118 2775 1122
rect 2779 1118 2780 1122
rect 2774 1117 2780 1118
rect 2966 1122 2972 1123
rect 2966 1118 2967 1122
rect 2971 1118 2972 1122
rect 2966 1117 2972 1118
rect 3158 1122 3164 1123
rect 3158 1118 3159 1122
rect 3163 1118 3164 1122
rect 3158 1117 3164 1118
rect 3342 1122 3348 1123
rect 3342 1118 3343 1122
rect 3347 1118 3348 1122
rect 3342 1117 3348 1118
rect 3510 1122 3516 1123
rect 3510 1118 3511 1122
rect 3515 1118 3516 1122
rect 3510 1117 3516 1118
rect 134 1108 140 1109
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 134 1104 135 1108
rect 139 1104 140 1108
rect 134 1103 140 1104
rect 246 1108 252 1109
rect 246 1104 247 1108
rect 251 1104 252 1108
rect 246 1103 252 1104
rect 382 1108 388 1109
rect 382 1104 383 1108
rect 387 1104 388 1108
rect 382 1103 388 1104
rect 518 1108 524 1109
rect 518 1104 519 1108
rect 523 1104 524 1108
rect 518 1103 524 1104
rect 646 1108 652 1109
rect 646 1104 647 1108
rect 651 1104 652 1108
rect 646 1103 652 1104
rect 774 1108 780 1109
rect 774 1104 775 1108
rect 779 1104 780 1108
rect 774 1103 780 1104
rect 894 1108 900 1109
rect 894 1104 895 1108
rect 899 1104 900 1108
rect 894 1103 900 1104
rect 1014 1108 1020 1109
rect 1014 1104 1015 1108
rect 1019 1104 1020 1108
rect 1014 1103 1020 1104
rect 1134 1108 1140 1109
rect 1134 1104 1135 1108
rect 1139 1104 1140 1108
rect 1134 1103 1140 1104
rect 1254 1108 1260 1109
rect 1254 1104 1255 1108
rect 1259 1104 1260 1108
rect 1254 1103 1260 1104
rect 1374 1108 1380 1109
rect 1374 1104 1375 1108
rect 1379 1104 1380 1108
rect 1374 1103 1380 1104
rect 1502 1108 1508 1109
rect 1502 1104 1503 1108
rect 1507 1104 1508 1108
rect 1502 1103 1508 1104
rect 1630 1108 1636 1109
rect 1630 1104 1631 1108
rect 1635 1104 1636 1108
rect 1630 1103 1636 1104
rect 1742 1108 1748 1109
rect 1742 1104 1743 1108
rect 1747 1104 1748 1108
rect 1742 1103 1748 1104
rect 1830 1105 1836 1106
rect 110 1100 116 1101
rect 1830 1101 1831 1105
rect 1835 1101 1836 1105
rect 1830 1100 1836 1101
rect 1870 1104 1876 1105
rect 1870 1100 1871 1104
rect 1875 1100 1876 1104
rect 127 1099 133 1100
rect 127 1095 128 1099
rect 132 1098 133 1099
rect 314 1099 320 1100
rect 314 1098 315 1099
rect 132 1096 153 1098
rect 309 1096 315 1098
rect 132 1095 133 1096
rect 127 1094 133 1095
rect 314 1095 315 1096
rect 319 1095 320 1099
rect 458 1099 464 1100
rect 458 1098 459 1099
rect 445 1096 459 1098
rect 314 1094 320 1095
rect 458 1095 459 1096
rect 463 1095 464 1099
rect 718 1099 724 1100
rect 718 1098 719 1099
rect 458 1094 464 1095
rect 359 1091 365 1092
rect 110 1088 116 1089
rect 110 1084 111 1088
rect 115 1084 116 1088
rect 359 1087 360 1091
rect 364 1090 365 1091
rect 536 1090 538 1097
rect 709 1096 719 1098
rect 718 1095 719 1096
rect 723 1095 724 1099
rect 854 1099 860 1100
rect 854 1098 855 1099
rect 837 1096 855 1098
rect 718 1094 724 1095
rect 854 1095 855 1096
rect 859 1095 860 1099
rect 962 1099 968 1100
rect 854 1094 860 1095
rect 364 1088 538 1090
rect 767 1091 773 1092
rect 364 1087 365 1088
rect 359 1086 365 1087
rect 767 1087 768 1091
rect 772 1090 773 1091
rect 912 1090 914 1097
rect 962 1095 963 1099
rect 967 1098 968 1099
rect 1082 1099 1088 1100
rect 967 1096 1033 1098
rect 967 1095 968 1096
rect 962 1094 968 1095
rect 1082 1095 1083 1099
rect 1087 1098 1088 1099
rect 1322 1099 1328 1100
rect 1322 1098 1323 1099
rect 1087 1096 1153 1098
rect 1317 1096 1323 1098
rect 1087 1095 1088 1096
rect 1082 1094 1088 1095
rect 1322 1095 1323 1096
rect 1327 1095 1328 1099
rect 1442 1099 1448 1100
rect 1442 1098 1443 1099
rect 1437 1096 1443 1098
rect 1322 1094 1328 1095
rect 1442 1095 1443 1096
rect 1447 1095 1448 1099
rect 1570 1099 1576 1100
rect 1442 1094 1448 1095
rect 1459 1096 1521 1098
rect 772 1088 914 1090
rect 1194 1091 1200 1092
rect 772 1087 773 1088
rect 767 1086 773 1087
rect 1194 1087 1195 1091
rect 1199 1090 1200 1091
rect 1459 1090 1461 1096
rect 1570 1095 1571 1099
rect 1575 1098 1576 1099
rect 1698 1099 1704 1100
rect 1870 1099 1876 1100
rect 3590 1104 3596 1105
rect 3590 1100 3591 1104
rect 3595 1100 3596 1104
rect 3590 1099 3596 1100
rect 1575 1096 1649 1098
rect 1575 1095 1576 1096
rect 1570 1094 1576 1095
rect 1698 1095 1699 1099
rect 1703 1098 1704 1099
rect 1703 1096 1761 1098
rect 1703 1095 1704 1096
rect 1698 1094 1704 1095
rect 2214 1095 2220 1096
rect 2214 1094 2215 1095
rect 2181 1092 2215 1094
rect 2214 1091 2215 1092
rect 2219 1091 2220 1095
rect 2214 1090 2220 1091
rect 2263 1095 2269 1096
rect 2263 1091 2264 1095
rect 2268 1094 2269 1095
rect 2626 1095 2632 1096
rect 2268 1092 2369 1094
rect 2268 1091 2269 1092
rect 2263 1090 2269 1091
rect 2626 1091 2627 1095
rect 2631 1091 2632 1095
rect 2626 1090 2632 1091
rect 2826 1095 2832 1096
rect 2826 1091 2827 1095
rect 2831 1091 2832 1095
rect 2826 1090 2832 1091
rect 3018 1095 3024 1096
rect 3018 1091 3019 1095
rect 3023 1091 3024 1095
rect 3018 1090 3024 1091
rect 3210 1095 3216 1096
rect 3210 1091 3211 1095
rect 3215 1091 3216 1095
rect 3210 1090 3216 1091
rect 3254 1095 3260 1096
rect 3254 1091 3255 1095
rect 3259 1094 3260 1095
rect 3518 1095 3524 1096
rect 3259 1092 3353 1094
rect 3259 1091 3260 1092
rect 3254 1090 3260 1091
rect 3518 1091 3519 1095
rect 3523 1091 3524 1095
rect 3518 1090 3524 1091
rect 1199 1088 1461 1090
rect 1830 1088 1836 1089
rect 1199 1087 1200 1088
rect 1194 1086 1200 1087
rect 110 1083 116 1084
rect 1830 1084 1831 1088
rect 1835 1084 1836 1088
rect 1830 1083 1836 1084
rect 1870 1087 1876 1088
rect 1870 1083 1871 1087
rect 1875 1083 1876 1087
rect 3590 1087 3596 1088
rect 1870 1082 1876 1083
rect 1894 1084 1900 1085
rect 1894 1080 1895 1084
rect 1899 1080 1900 1084
rect 1894 1079 1900 1080
rect 2118 1084 2124 1085
rect 2118 1080 2119 1084
rect 2123 1080 2124 1084
rect 2118 1079 2124 1080
rect 2350 1084 2356 1085
rect 2350 1080 2351 1084
rect 2355 1080 2356 1084
rect 2350 1079 2356 1080
rect 2566 1084 2572 1085
rect 2566 1080 2567 1084
rect 2571 1080 2572 1084
rect 2566 1079 2572 1080
rect 2766 1084 2772 1085
rect 2766 1080 2767 1084
rect 2771 1080 2772 1084
rect 2766 1079 2772 1080
rect 2958 1084 2964 1085
rect 2958 1080 2959 1084
rect 2963 1080 2964 1084
rect 2958 1079 2964 1080
rect 3150 1084 3156 1085
rect 3150 1080 3151 1084
rect 3155 1080 3156 1084
rect 3150 1079 3156 1080
rect 3334 1084 3340 1085
rect 3334 1080 3335 1084
rect 3339 1080 3340 1084
rect 3334 1079 3340 1080
rect 3502 1084 3508 1085
rect 3502 1080 3503 1084
rect 3507 1080 3508 1084
rect 3590 1083 3591 1087
rect 3595 1083 3596 1087
rect 3590 1082 3596 1083
rect 3502 1079 3508 1080
rect 142 1070 148 1071
rect 142 1066 143 1070
rect 147 1066 148 1070
rect 142 1065 148 1066
rect 254 1070 260 1071
rect 254 1066 255 1070
rect 259 1066 260 1070
rect 254 1065 260 1066
rect 390 1070 396 1071
rect 390 1066 391 1070
rect 395 1066 396 1070
rect 390 1065 396 1066
rect 526 1070 532 1071
rect 526 1066 527 1070
rect 531 1066 532 1070
rect 526 1065 532 1066
rect 654 1070 660 1071
rect 654 1066 655 1070
rect 659 1066 660 1070
rect 654 1065 660 1066
rect 782 1070 788 1071
rect 782 1066 783 1070
rect 787 1066 788 1070
rect 782 1065 788 1066
rect 902 1070 908 1071
rect 902 1066 903 1070
rect 907 1066 908 1070
rect 902 1065 908 1066
rect 1022 1070 1028 1071
rect 1022 1066 1023 1070
rect 1027 1066 1028 1070
rect 1022 1065 1028 1066
rect 1142 1070 1148 1071
rect 1142 1066 1143 1070
rect 1147 1066 1148 1070
rect 1142 1065 1148 1066
rect 1262 1070 1268 1071
rect 1262 1066 1263 1070
rect 1267 1066 1268 1070
rect 1262 1065 1268 1066
rect 1382 1070 1388 1071
rect 1382 1066 1383 1070
rect 1387 1066 1388 1070
rect 1382 1065 1388 1066
rect 1510 1070 1516 1071
rect 1510 1066 1511 1070
rect 1515 1066 1516 1070
rect 1510 1065 1516 1066
rect 1638 1070 1644 1071
rect 1638 1066 1639 1070
rect 1643 1066 1644 1070
rect 1638 1065 1644 1066
rect 1750 1070 1756 1071
rect 1750 1066 1751 1070
rect 1755 1066 1756 1070
rect 1911 1067 1917 1068
rect 1911 1066 1912 1067
rect 1750 1065 1756 1066
rect 1828 1064 1912 1066
rect 135 1059 141 1060
rect 135 1055 136 1059
rect 140 1058 141 1059
rect 150 1059 156 1060
rect 150 1058 151 1059
rect 140 1056 151 1058
rect 140 1055 141 1056
rect 135 1054 141 1055
rect 150 1055 151 1056
rect 155 1055 156 1059
rect 150 1054 156 1055
rect 247 1059 253 1060
rect 247 1055 248 1059
rect 252 1058 253 1059
rect 262 1059 268 1060
rect 262 1058 263 1059
rect 252 1056 263 1058
rect 252 1055 253 1056
rect 247 1054 253 1055
rect 262 1055 263 1056
rect 267 1055 268 1059
rect 262 1054 268 1055
rect 314 1059 320 1060
rect 314 1055 315 1059
rect 319 1058 320 1059
rect 383 1059 389 1060
rect 383 1058 384 1059
rect 319 1056 384 1058
rect 319 1055 320 1056
rect 314 1054 320 1055
rect 383 1055 384 1056
rect 388 1055 389 1059
rect 383 1054 389 1055
rect 458 1059 464 1060
rect 458 1055 459 1059
rect 463 1058 464 1059
rect 519 1059 525 1060
rect 519 1058 520 1059
rect 463 1056 520 1058
rect 463 1055 464 1056
rect 458 1054 464 1055
rect 519 1055 520 1056
rect 524 1055 525 1059
rect 519 1054 525 1055
rect 626 1059 632 1060
rect 626 1055 627 1059
rect 631 1058 632 1059
rect 647 1059 653 1060
rect 647 1058 648 1059
rect 631 1056 648 1058
rect 631 1055 632 1056
rect 626 1054 632 1055
rect 647 1055 648 1056
rect 652 1055 653 1059
rect 647 1054 653 1055
rect 718 1059 724 1060
rect 718 1055 719 1059
rect 723 1058 724 1059
rect 775 1059 781 1060
rect 775 1058 776 1059
rect 723 1056 776 1058
rect 723 1055 724 1056
rect 718 1054 724 1055
rect 775 1055 776 1056
rect 780 1055 781 1059
rect 775 1054 781 1055
rect 895 1059 901 1060
rect 895 1055 896 1059
rect 900 1058 901 1059
rect 962 1059 968 1060
rect 962 1058 963 1059
rect 900 1056 963 1058
rect 900 1055 901 1056
rect 895 1054 901 1055
rect 962 1055 963 1056
rect 967 1055 968 1059
rect 962 1054 968 1055
rect 1015 1059 1021 1060
rect 1015 1055 1016 1059
rect 1020 1058 1021 1059
rect 1082 1059 1088 1060
rect 1082 1058 1083 1059
rect 1020 1056 1083 1058
rect 1020 1055 1021 1056
rect 1015 1054 1021 1055
rect 1082 1055 1083 1056
rect 1087 1055 1088 1059
rect 1082 1054 1088 1055
rect 1135 1059 1141 1060
rect 1135 1055 1136 1059
rect 1140 1058 1141 1059
rect 1194 1059 1200 1060
rect 1194 1058 1195 1059
rect 1140 1056 1195 1058
rect 1140 1055 1141 1056
rect 1135 1054 1141 1055
rect 1194 1055 1195 1056
rect 1199 1055 1200 1059
rect 1194 1054 1200 1055
rect 1210 1059 1216 1060
rect 1210 1055 1211 1059
rect 1215 1058 1216 1059
rect 1255 1059 1261 1060
rect 1255 1058 1256 1059
rect 1215 1056 1256 1058
rect 1215 1055 1216 1056
rect 1210 1054 1216 1055
rect 1255 1055 1256 1056
rect 1260 1055 1261 1059
rect 1255 1054 1261 1055
rect 1322 1059 1328 1060
rect 1322 1055 1323 1059
rect 1327 1058 1328 1059
rect 1375 1059 1381 1060
rect 1375 1058 1376 1059
rect 1327 1056 1376 1058
rect 1327 1055 1328 1056
rect 1322 1054 1328 1055
rect 1375 1055 1376 1056
rect 1380 1055 1381 1059
rect 1375 1054 1381 1055
rect 1442 1059 1448 1060
rect 1442 1055 1443 1059
rect 1447 1058 1448 1059
rect 1503 1059 1509 1060
rect 1503 1058 1504 1059
rect 1447 1056 1504 1058
rect 1447 1055 1448 1056
rect 1442 1054 1448 1055
rect 1503 1055 1504 1056
rect 1508 1055 1509 1059
rect 1503 1054 1509 1055
rect 1631 1059 1637 1060
rect 1631 1055 1632 1059
rect 1636 1058 1637 1059
rect 1698 1059 1704 1060
rect 1698 1058 1699 1059
rect 1636 1056 1699 1058
rect 1636 1055 1637 1056
rect 1631 1054 1637 1055
rect 1698 1055 1699 1056
rect 1703 1055 1704 1059
rect 1698 1054 1704 1055
rect 1743 1059 1749 1060
rect 1743 1055 1744 1059
rect 1748 1058 1749 1059
rect 1828 1058 1830 1064
rect 1911 1063 1912 1064
rect 1916 1063 1917 1067
rect 1911 1062 1917 1063
rect 1748 1056 1830 1058
rect 1748 1055 1749 1056
rect 1743 1054 1749 1055
rect 678 1043 684 1044
rect 678 1042 679 1043
rect 528 1040 679 1042
rect 127 1035 133 1036
rect 127 1031 128 1035
rect 132 1034 133 1035
rect 135 1035 141 1036
rect 135 1034 136 1035
rect 132 1032 136 1034
rect 132 1031 133 1032
rect 127 1030 133 1031
rect 135 1031 136 1032
rect 140 1031 141 1035
rect 135 1030 141 1031
rect 231 1035 237 1036
rect 231 1031 232 1035
rect 236 1034 237 1035
rect 298 1035 304 1036
rect 298 1034 299 1035
rect 236 1032 299 1034
rect 236 1031 237 1032
rect 231 1030 237 1031
rect 298 1031 299 1032
rect 303 1031 304 1035
rect 298 1030 304 1031
rect 351 1035 357 1036
rect 351 1031 352 1035
rect 356 1034 357 1035
rect 359 1035 365 1036
rect 359 1034 360 1035
rect 356 1032 360 1034
rect 356 1031 357 1032
rect 351 1030 357 1031
rect 359 1031 360 1032
rect 364 1031 365 1035
rect 359 1030 365 1031
rect 463 1035 469 1036
rect 463 1031 464 1035
rect 468 1034 469 1035
rect 528 1034 530 1040
rect 678 1039 679 1040
rect 683 1039 684 1043
rect 678 1038 684 1039
rect 1894 1040 1900 1041
rect 1870 1037 1876 1038
rect 468 1032 530 1034
rect 534 1035 540 1036
rect 468 1031 469 1032
rect 463 1030 469 1031
rect 534 1031 535 1035
rect 539 1034 540 1035
rect 567 1035 573 1036
rect 567 1034 568 1035
rect 539 1032 568 1034
rect 539 1031 540 1032
rect 534 1030 540 1031
rect 567 1031 568 1032
rect 572 1031 573 1035
rect 567 1030 573 1031
rect 663 1035 669 1036
rect 663 1031 664 1035
rect 668 1034 669 1035
rect 686 1035 692 1036
rect 686 1034 687 1035
rect 668 1032 687 1034
rect 668 1031 669 1032
rect 663 1030 669 1031
rect 686 1031 687 1032
rect 691 1031 692 1035
rect 686 1030 692 1031
rect 759 1035 765 1036
rect 759 1031 760 1035
rect 764 1034 765 1035
rect 767 1035 773 1036
rect 767 1034 768 1035
rect 764 1032 768 1034
rect 764 1031 765 1032
rect 759 1030 765 1031
rect 767 1031 768 1032
rect 772 1031 773 1035
rect 767 1030 773 1031
rect 818 1035 824 1036
rect 818 1031 819 1035
rect 823 1034 824 1035
rect 847 1035 853 1036
rect 847 1034 848 1035
rect 823 1032 848 1034
rect 823 1031 824 1032
rect 818 1030 824 1031
rect 847 1031 848 1032
rect 852 1031 853 1035
rect 847 1030 853 1031
rect 934 1035 941 1036
rect 934 1031 935 1035
rect 940 1031 941 1035
rect 934 1030 941 1031
rect 994 1035 1000 1036
rect 994 1031 995 1035
rect 999 1034 1000 1035
rect 1023 1035 1029 1036
rect 1023 1034 1024 1035
rect 999 1032 1024 1034
rect 999 1031 1000 1032
rect 994 1030 1000 1031
rect 1023 1031 1024 1032
rect 1028 1031 1029 1035
rect 1023 1030 1029 1031
rect 1082 1035 1088 1036
rect 1082 1031 1083 1035
rect 1087 1034 1088 1035
rect 1119 1035 1125 1036
rect 1119 1034 1120 1035
rect 1087 1032 1120 1034
rect 1087 1031 1088 1032
rect 1082 1030 1088 1031
rect 1119 1031 1120 1032
rect 1124 1031 1125 1035
rect 1119 1030 1125 1031
rect 1178 1035 1184 1036
rect 1178 1031 1179 1035
rect 1183 1034 1184 1035
rect 1215 1035 1221 1036
rect 1215 1034 1216 1035
rect 1183 1032 1216 1034
rect 1183 1031 1184 1032
rect 1178 1030 1184 1031
rect 1215 1031 1216 1032
rect 1220 1031 1221 1035
rect 1870 1033 1871 1037
rect 1875 1033 1876 1037
rect 1894 1036 1895 1040
rect 1899 1036 1900 1040
rect 1894 1035 1900 1036
rect 2014 1040 2020 1041
rect 2014 1036 2015 1040
rect 2019 1036 2020 1040
rect 2014 1035 2020 1036
rect 2166 1040 2172 1041
rect 2166 1036 2167 1040
rect 2171 1036 2172 1040
rect 2166 1035 2172 1036
rect 2326 1040 2332 1041
rect 2326 1036 2327 1040
rect 2331 1036 2332 1040
rect 2326 1035 2332 1036
rect 2486 1040 2492 1041
rect 2486 1036 2487 1040
rect 2491 1036 2492 1040
rect 2486 1035 2492 1036
rect 2638 1040 2644 1041
rect 2638 1036 2639 1040
rect 2643 1036 2644 1040
rect 2638 1035 2644 1036
rect 2790 1040 2796 1041
rect 2790 1036 2791 1040
rect 2795 1036 2796 1040
rect 2790 1035 2796 1036
rect 2934 1040 2940 1041
rect 2934 1036 2935 1040
rect 2939 1036 2940 1040
rect 2934 1035 2940 1036
rect 3078 1040 3084 1041
rect 3078 1036 3079 1040
rect 3083 1036 3084 1040
rect 3078 1035 3084 1036
rect 3222 1040 3228 1041
rect 3222 1036 3223 1040
rect 3227 1036 3228 1040
rect 3222 1035 3228 1036
rect 3374 1040 3380 1041
rect 3374 1036 3375 1040
rect 3379 1036 3380 1040
rect 3374 1035 3380 1036
rect 3502 1040 3508 1041
rect 3502 1036 3503 1040
rect 3507 1036 3508 1040
rect 3502 1035 3508 1036
rect 3590 1037 3596 1038
rect 1870 1032 1876 1033
rect 3590 1033 3591 1037
rect 3595 1033 3596 1037
rect 3590 1032 3596 1033
rect 1215 1030 1221 1031
rect 1887 1031 1893 1032
rect 1887 1027 1888 1031
rect 1892 1030 1893 1031
rect 1962 1031 1968 1032
rect 1892 1028 1913 1030
rect 1892 1027 1893 1028
rect 142 1026 148 1027
rect 142 1022 143 1026
rect 147 1022 148 1026
rect 142 1021 148 1022
rect 238 1026 244 1027
rect 238 1022 239 1026
rect 243 1022 244 1026
rect 238 1021 244 1022
rect 358 1026 364 1027
rect 358 1022 359 1026
rect 363 1022 364 1026
rect 358 1021 364 1022
rect 470 1026 476 1027
rect 470 1022 471 1026
rect 475 1022 476 1026
rect 470 1021 476 1022
rect 574 1026 580 1027
rect 574 1022 575 1026
rect 579 1022 580 1026
rect 574 1021 580 1022
rect 670 1026 676 1027
rect 670 1022 671 1026
rect 675 1022 676 1026
rect 670 1021 676 1022
rect 766 1026 772 1027
rect 766 1022 767 1026
rect 771 1022 772 1026
rect 766 1021 772 1022
rect 854 1026 860 1027
rect 854 1022 855 1026
rect 859 1022 860 1026
rect 854 1021 860 1022
rect 942 1026 948 1027
rect 942 1022 943 1026
rect 947 1022 948 1026
rect 942 1021 948 1022
rect 1030 1026 1036 1027
rect 1030 1022 1031 1026
rect 1035 1022 1036 1026
rect 1030 1021 1036 1022
rect 1126 1026 1132 1027
rect 1126 1022 1127 1026
rect 1131 1022 1132 1026
rect 1126 1021 1132 1022
rect 1222 1026 1228 1027
rect 1887 1026 1893 1027
rect 1962 1027 1963 1031
rect 1967 1030 1968 1031
rect 2082 1031 2088 1032
rect 1967 1028 2033 1030
rect 1967 1027 1968 1028
rect 1962 1026 1968 1027
rect 2082 1027 2083 1031
rect 2087 1030 2088 1031
rect 2414 1031 2420 1032
rect 2414 1030 2415 1031
rect 2087 1028 2185 1030
rect 2389 1028 2415 1030
rect 2087 1027 2088 1028
rect 2082 1026 2088 1027
rect 2414 1027 2415 1028
rect 2419 1027 2420 1031
rect 2414 1026 2420 1027
rect 2479 1031 2485 1032
rect 2479 1027 2480 1031
rect 2484 1030 2485 1031
rect 2631 1031 2637 1032
rect 2484 1028 2505 1030
rect 2484 1027 2485 1028
rect 2479 1026 2485 1027
rect 2631 1027 2632 1031
rect 2636 1030 2637 1031
rect 2706 1031 2712 1032
rect 2636 1028 2657 1030
rect 2636 1027 2637 1028
rect 2631 1026 2637 1027
rect 2706 1027 2707 1031
rect 2711 1030 2712 1031
rect 2858 1031 2864 1032
rect 2711 1028 2809 1030
rect 2711 1027 2712 1028
rect 2706 1026 2712 1027
rect 2858 1027 2859 1031
rect 2863 1030 2864 1031
rect 3002 1031 3008 1032
rect 2863 1028 2953 1030
rect 2863 1027 2864 1028
rect 2858 1026 2864 1027
rect 3002 1027 3003 1031
rect 3007 1030 3008 1031
rect 3306 1031 3312 1032
rect 3306 1030 3307 1031
rect 3007 1028 3097 1030
rect 3285 1028 3307 1030
rect 3007 1027 3008 1028
rect 3002 1026 3008 1027
rect 3306 1027 3307 1028
rect 3311 1027 3312 1031
rect 3306 1026 3312 1027
rect 3343 1031 3349 1032
rect 3343 1027 3344 1031
rect 3348 1030 3349 1031
rect 3495 1031 3501 1032
rect 3348 1028 3393 1030
rect 3348 1027 3349 1028
rect 3343 1026 3349 1027
rect 3495 1027 3496 1031
rect 3500 1030 3501 1031
rect 3500 1028 3521 1030
rect 3500 1027 3501 1028
rect 3495 1026 3501 1027
rect 1222 1022 1223 1026
rect 1227 1022 1228 1026
rect 1222 1021 1228 1022
rect 1870 1020 1876 1021
rect 1870 1016 1871 1020
rect 1875 1016 1876 1020
rect 1870 1015 1876 1016
rect 3590 1020 3596 1021
rect 3590 1016 3591 1020
rect 3595 1016 3596 1020
rect 3590 1015 3596 1016
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 1830 1008 1836 1009
rect 1830 1004 1831 1008
rect 1835 1004 1836 1008
rect 1830 1003 1836 1004
rect 1902 1002 1908 1003
rect 150 999 156 1000
rect 150 995 151 999
rect 155 995 156 999
rect 150 994 156 995
rect 298 999 304 1000
rect 298 995 299 999
rect 303 998 304 999
rect 534 999 540 1000
rect 534 998 535 999
rect 303 996 369 998
rect 525 996 535 998
rect 303 995 304 996
rect 298 994 304 995
rect 534 995 535 996
rect 539 995 540 999
rect 534 994 540 995
rect 626 999 632 1000
rect 626 995 627 999
rect 631 995 632 999
rect 626 994 632 995
rect 678 999 684 1000
rect 678 995 679 999
rect 683 995 684 999
rect 678 994 684 995
rect 818 999 824 1000
rect 818 995 819 999
rect 823 995 824 999
rect 934 999 940 1000
rect 934 998 935 999
rect 909 996 935 998
rect 818 994 824 995
rect 934 995 935 996
rect 939 995 940 999
rect 934 994 940 995
rect 994 999 1000 1000
rect 994 995 995 999
rect 999 995 1000 999
rect 994 994 1000 995
rect 1082 999 1088 1000
rect 1082 995 1083 999
rect 1087 995 1088 999
rect 1082 994 1088 995
rect 1178 999 1184 1000
rect 1178 995 1179 999
rect 1183 995 1184 999
rect 1902 998 1903 1002
rect 1907 998 1908 1002
rect 1902 997 1908 998
rect 2022 1002 2028 1003
rect 2022 998 2023 1002
rect 2027 998 2028 1002
rect 2022 997 2028 998
rect 2174 1002 2180 1003
rect 2174 998 2175 1002
rect 2179 998 2180 1002
rect 2174 997 2180 998
rect 2334 1002 2340 1003
rect 2334 998 2335 1002
rect 2339 998 2340 1002
rect 2334 997 2340 998
rect 2494 1002 2500 1003
rect 2494 998 2495 1002
rect 2499 998 2500 1002
rect 2494 997 2500 998
rect 2646 1002 2652 1003
rect 2646 998 2647 1002
rect 2651 998 2652 1002
rect 2646 997 2652 998
rect 2798 1002 2804 1003
rect 2798 998 2799 1002
rect 2803 998 2804 1002
rect 2798 997 2804 998
rect 2942 1002 2948 1003
rect 2942 998 2943 1002
rect 2947 998 2948 1002
rect 2942 997 2948 998
rect 3086 1002 3092 1003
rect 3086 998 3087 1002
rect 3091 998 3092 1002
rect 3086 997 3092 998
rect 3230 1002 3236 1003
rect 3230 998 3231 1002
rect 3235 998 3236 1002
rect 3230 997 3236 998
rect 3382 1002 3388 1003
rect 3382 998 3383 1002
rect 3387 998 3388 1002
rect 3382 997 3388 998
rect 3510 1002 3516 1003
rect 3510 998 3511 1002
rect 3515 998 3516 1002
rect 3510 997 3516 998
rect 1178 994 1184 995
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1830 991 1836 992
rect 110 986 116 987
rect 134 988 140 989
rect 134 984 135 988
rect 139 984 140 988
rect 134 983 140 984
rect 230 988 236 989
rect 230 984 231 988
rect 235 984 236 988
rect 230 983 236 984
rect 350 988 356 989
rect 350 984 351 988
rect 355 984 356 988
rect 350 983 356 984
rect 462 988 468 989
rect 462 984 463 988
rect 467 984 468 988
rect 462 983 468 984
rect 566 988 572 989
rect 566 984 567 988
rect 571 984 572 988
rect 566 983 572 984
rect 662 988 668 989
rect 662 984 663 988
rect 667 984 668 988
rect 662 983 668 984
rect 758 988 764 989
rect 758 984 759 988
rect 763 984 764 988
rect 758 983 764 984
rect 846 988 852 989
rect 846 984 847 988
rect 851 984 852 988
rect 846 983 852 984
rect 934 988 940 989
rect 934 984 935 988
rect 939 984 940 988
rect 934 983 940 984
rect 1022 988 1028 989
rect 1022 984 1023 988
rect 1027 984 1028 988
rect 1022 983 1028 984
rect 1118 988 1124 989
rect 1118 984 1119 988
rect 1123 984 1124 988
rect 1118 983 1124 984
rect 1214 988 1220 989
rect 1214 984 1215 988
rect 1219 984 1220 988
rect 1830 987 1831 991
rect 1835 987 1836 991
rect 1830 986 1836 987
rect 1895 991 1901 992
rect 1895 987 1896 991
rect 1900 990 1901 991
rect 1962 991 1968 992
rect 1962 990 1963 991
rect 1900 988 1963 990
rect 1900 987 1901 988
rect 1895 986 1901 987
rect 1962 987 1963 988
rect 1967 987 1968 991
rect 1962 986 1968 987
rect 2015 991 2021 992
rect 2015 987 2016 991
rect 2020 990 2021 991
rect 2082 991 2088 992
rect 2082 990 2083 991
rect 2020 988 2083 990
rect 2020 987 2021 988
rect 2015 986 2021 987
rect 2082 987 2083 988
rect 2087 987 2088 991
rect 2082 986 2088 987
rect 2167 991 2173 992
rect 2167 987 2168 991
rect 2172 990 2173 991
rect 2206 991 2212 992
rect 2206 990 2207 991
rect 2172 988 2207 990
rect 2172 987 2173 988
rect 2167 986 2173 987
rect 2206 987 2207 988
rect 2211 987 2212 991
rect 2206 986 2212 987
rect 2214 991 2220 992
rect 2214 987 2215 991
rect 2219 990 2220 991
rect 2327 991 2333 992
rect 2327 990 2328 991
rect 2219 988 2328 990
rect 2219 987 2220 988
rect 2214 986 2220 987
rect 2327 987 2328 988
rect 2332 987 2333 991
rect 2327 986 2333 987
rect 2414 991 2420 992
rect 2414 987 2415 991
rect 2419 990 2420 991
rect 2487 991 2493 992
rect 2487 990 2488 991
rect 2419 988 2488 990
rect 2419 987 2420 988
rect 2414 986 2420 987
rect 2487 987 2488 988
rect 2492 987 2493 991
rect 2487 986 2493 987
rect 2639 991 2645 992
rect 2639 987 2640 991
rect 2644 990 2645 991
rect 2706 991 2712 992
rect 2706 990 2707 991
rect 2644 988 2707 990
rect 2644 987 2645 988
rect 2639 986 2645 987
rect 2706 987 2707 988
rect 2711 987 2712 991
rect 2706 986 2712 987
rect 2791 991 2797 992
rect 2791 987 2792 991
rect 2796 990 2797 991
rect 2858 991 2864 992
rect 2858 990 2859 991
rect 2796 988 2859 990
rect 2796 987 2797 988
rect 2791 986 2797 987
rect 2858 987 2859 988
rect 2863 987 2864 991
rect 2858 986 2864 987
rect 2935 991 2941 992
rect 2935 987 2936 991
rect 2940 990 2941 991
rect 3002 991 3008 992
rect 3002 990 3003 991
rect 2940 988 3003 990
rect 2940 987 2941 988
rect 2935 986 2941 987
rect 3002 987 3003 988
rect 3007 987 3008 991
rect 3002 986 3008 987
rect 3018 991 3024 992
rect 3018 987 3019 991
rect 3023 990 3024 991
rect 3079 991 3085 992
rect 3079 990 3080 991
rect 3023 988 3080 990
rect 3023 987 3024 988
rect 3018 986 3024 987
rect 3079 987 3080 988
rect 3084 987 3085 991
rect 3079 986 3085 987
rect 3210 991 3216 992
rect 3210 987 3211 991
rect 3215 990 3216 991
rect 3223 991 3229 992
rect 3223 990 3224 991
rect 3215 988 3224 990
rect 3215 987 3216 988
rect 3210 986 3216 987
rect 3223 987 3224 988
rect 3228 987 3229 991
rect 3223 986 3229 987
rect 3306 991 3312 992
rect 3306 987 3307 991
rect 3311 990 3312 991
rect 3375 991 3381 992
rect 3375 990 3376 991
rect 3311 988 3376 990
rect 3311 987 3312 988
rect 3306 986 3312 987
rect 3375 987 3376 988
rect 3380 987 3381 991
rect 3375 986 3381 987
rect 3503 991 3509 992
rect 3503 987 3504 991
rect 3508 990 3509 991
rect 3518 991 3524 992
rect 3518 990 3519 991
rect 3508 988 3519 990
rect 3508 987 3509 988
rect 3503 986 3509 987
rect 3518 987 3519 988
rect 3523 987 3524 991
rect 3518 986 3524 987
rect 1214 983 1220 984
rect 1887 975 1893 976
rect 247 971 253 972
rect 247 967 248 971
rect 252 970 253 971
rect 255 971 261 972
rect 255 970 256 971
rect 252 968 256 970
rect 252 967 253 968
rect 247 966 253 967
rect 255 967 256 968
rect 260 967 261 971
rect 255 966 261 967
rect 1215 971 1221 972
rect 1215 967 1216 971
rect 1220 970 1221 971
rect 1231 971 1237 972
rect 1231 970 1232 971
rect 1220 968 1232 970
rect 1220 967 1221 968
rect 1215 966 1221 967
rect 1231 967 1232 968
rect 1236 967 1237 971
rect 1887 971 1888 975
rect 1892 974 1893 975
rect 1895 975 1901 976
rect 1895 974 1896 975
rect 1892 972 1896 974
rect 1892 971 1893 972
rect 1887 970 1893 971
rect 1895 971 1896 972
rect 1900 971 1901 975
rect 1895 970 1901 971
rect 1954 975 1960 976
rect 1954 971 1955 975
rect 1959 974 1960 975
rect 1975 975 1981 976
rect 1975 974 1976 975
rect 1959 972 1976 974
rect 1959 971 1960 972
rect 1954 970 1960 971
rect 1975 971 1976 972
rect 1980 971 1981 975
rect 1975 970 1981 971
rect 2034 975 2040 976
rect 2034 971 2035 975
rect 2039 974 2040 975
rect 2071 975 2077 976
rect 2071 974 2072 975
rect 2039 972 2072 974
rect 2039 971 2040 972
rect 2034 970 2040 971
rect 2071 971 2072 972
rect 2076 971 2077 975
rect 2071 970 2077 971
rect 2130 975 2136 976
rect 2130 971 2131 975
rect 2135 974 2136 975
rect 2191 975 2197 976
rect 2191 974 2192 975
rect 2135 972 2192 974
rect 2135 971 2136 972
rect 2130 970 2136 971
rect 2191 971 2192 972
rect 2196 971 2197 975
rect 2191 970 2197 971
rect 2327 975 2333 976
rect 2327 971 2328 975
rect 2332 974 2333 975
rect 2406 975 2412 976
rect 2406 974 2407 975
rect 2332 972 2407 974
rect 2332 971 2333 972
rect 2327 970 2333 971
rect 2406 971 2407 972
rect 2411 971 2412 975
rect 2406 970 2412 971
rect 2471 975 2477 976
rect 2471 971 2472 975
rect 2476 974 2477 975
rect 2479 975 2485 976
rect 2479 974 2480 975
rect 2476 972 2480 974
rect 2476 971 2477 972
rect 2471 970 2477 971
rect 2479 971 2480 972
rect 2484 971 2485 975
rect 2479 970 2485 971
rect 2623 975 2629 976
rect 2623 971 2624 975
rect 2628 974 2629 975
rect 2631 975 2637 976
rect 2631 974 2632 975
rect 2628 972 2632 974
rect 2628 971 2629 972
rect 2623 970 2629 971
rect 2631 971 2632 972
rect 2636 971 2637 975
rect 2631 970 2637 971
rect 2682 975 2688 976
rect 2682 971 2683 975
rect 2687 974 2688 975
rect 2783 975 2789 976
rect 2783 974 2784 975
rect 2687 972 2784 974
rect 2687 971 2688 972
rect 2682 970 2688 971
rect 2783 971 2784 972
rect 2788 971 2789 975
rect 2783 970 2789 971
rect 2842 975 2848 976
rect 2842 971 2843 975
rect 2847 974 2848 975
rect 2959 975 2965 976
rect 2959 974 2960 975
rect 2847 972 2960 974
rect 2847 971 2848 972
rect 2842 970 2848 971
rect 2959 971 2960 972
rect 2964 971 2965 975
rect 2959 970 2965 971
rect 3143 975 3149 976
rect 3143 971 3144 975
rect 3148 974 3149 975
rect 3210 975 3216 976
rect 3210 974 3211 975
rect 3148 972 3211 974
rect 3148 971 3149 972
rect 3143 970 3149 971
rect 3210 971 3211 972
rect 3215 971 3216 975
rect 3210 970 3216 971
rect 3335 975 3341 976
rect 3335 971 3336 975
rect 3340 974 3341 975
rect 3343 975 3349 976
rect 3343 974 3344 975
rect 3340 972 3344 974
rect 3340 971 3341 972
rect 3335 970 3341 971
rect 3343 971 3344 972
rect 3348 971 3349 975
rect 3343 970 3349 971
rect 3495 975 3501 976
rect 3495 971 3496 975
rect 3500 974 3501 975
rect 3503 975 3509 976
rect 3503 974 3504 975
rect 3500 972 3504 974
rect 3500 971 3501 972
rect 3495 970 3501 971
rect 3503 971 3504 972
rect 3508 971 3509 975
rect 3503 970 3509 971
rect 1231 966 1237 967
rect 1902 966 1908 967
rect 1902 962 1903 966
rect 1907 962 1908 966
rect 1902 961 1908 962
rect 1982 966 1988 967
rect 1982 962 1983 966
rect 1987 962 1988 966
rect 1982 961 1988 962
rect 2078 966 2084 967
rect 2078 962 2079 966
rect 2083 962 2084 966
rect 2078 961 2084 962
rect 2198 966 2204 967
rect 2198 962 2199 966
rect 2203 962 2204 966
rect 2198 961 2204 962
rect 2334 966 2340 967
rect 2334 962 2335 966
rect 2339 962 2340 966
rect 2334 961 2340 962
rect 2478 966 2484 967
rect 2478 962 2479 966
rect 2483 962 2484 966
rect 2478 961 2484 962
rect 2630 966 2636 967
rect 2630 962 2631 966
rect 2635 962 2636 966
rect 2630 961 2636 962
rect 2790 966 2796 967
rect 2790 962 2791 966
rect 2795 962 2796 966
rect 2790 961 2796 962
rect 2966 966 2972 967
rect 2966 962 2967 966
rect 2971 962 2972 966
rect 2966 961 2972 962
rect 3150 966 3156 967
rect 3150 962 3151 966
rect 3155 962 3156 966
rect 3150 961 3156 962
rect 3342 966 3348 967
rect 3342 962 3343 966
rect 3347 962 3348 966
rect 3342 961 3348 962
rect 3510 966 3516 967
rect 3510 962 3511 966
rect 3515 962 3516 966
rect 3510 961 3516 962
rect 1870 948 1876 949
rect 1870 944 1871 948
rect 1875 944 1876 948
rect 1870 943 1876 944
rect 3590 948 3596 949
rect 3590 944 3591 948
rect 3595 944 3596 948
rect 3590 943 3596 944
rect 1954 939 1960 940
rect 1954 935 1955 939
rect 1959 935 1960 939
rect 1954 934 1960 935
rect 2034 939 2040 940
rect 2034 935 2035 939
rect 2039 935 2040 939
rect 2034 934 2040 935
rect 2130 939 2136 940
rect 2130 935 2131 939
rect 2135 935 2136 939
rect 2130 934 2136 935
rect 2206 939 2212 940
rect 2206 935 2207 939
rect 2211 935 2212 939
rect 2206 934 2212 935
rect 2406 939 2412 940
rect 2406 935 2407 939
rect 2411 938 2412 939
rect 2682 939 2688 940
rect 2411 936 2489 938
rect 2411 935 2412 936
rect 2406 934 2412 935
rect 2682 935 2683 939
rect 2687 935 2688 939
rect 2682 934 2688 935
rect 2842 939 2848 940
rect 2842 935 2843 939
rect 2847 935 2848 939
rect 2842 934 2848 935
rect 3202 939 3208 940
rect 3202 935 3203 939
rect 3207 935 3208 939
rect 3202 934 3208 935
rect 3210 939 3216 940
rect 3210 935 3211 939
rect 3215 938 3216 939
rect 3518 939 3524 940
rect 3215 936 3353 938
rect 3215 935 3216 936
rect 3210 934 3216 935
rect 3518 935 3519 939
rect 3523 935 3524 939
rect 3518 934 3524 935
rect 134 932 140 933
rect 110 929 116 930
rect 110 925 111 929
rect 115 925 116 929
rect 134 928 135 932
rect 139 928 140 932
rect 134 927 140 928
rect 262 932 268 933
rect 262 928 263 932
rect 267 928 268 932
rect 262 927 268 928
rect 414 932 420 933
rect 414 928 415 932
rect 419 928 420 932
rect 414 927 420 928
rect 558 932 564 933
rect 558 928 559 932
rect 563 928 564 932
rect 558 927 564 928
rect 702 932 708 933
rect 702 928 703 932
rect 707 928 708 932
rect 702 927 708 928
rect 838 932 844 933
rect 838 928 839 932
rect 843 928 844 932
rect 838 927 844 928
rect 974 932 980 933
rect 974 928 975 932
rect 979 928 980 932
rect 974 927 980 928
rect 1102 932 1108 933
rect 1102 928 1103 932
rect 1107 928 1108 932
rect 1102 927 1108 928
rect 1222 932 1228 933
rect 1222 928 1223 932
rect 1227 928 1228 932
rect 1222 927 1228 928
rect 1334 932 1340 933
rect 1334 928 1335 932
rect 1339 928 1340 932
rect 1334 927 1340 928
rect 1438 932 1444 933
rect 1438 928 1439 932
rect 1443 928 1444 932
rect 1438 927 1444 928
rect 1542 932 1548 933
rect 1542 928 1543 932
rect 1547 928 1548 932
rect 1542 927 1548 928
rect 1654 932 1660 933
rect 1654 928 1655 932
rect 1659 928 1660 932
rect 1654 927 1660 928
rect 1742 932 1748 933
rect 1742 928 1743 932
rect 1747 928 1748 932
rect 1870 931 1876 932
rect 1742 927 1748 928
rect 1830 929 1836 930
rect 110 924 116 925
rect 1830 925 1831 929
rect 1835 925 1836 929
rect 1870 927 1871 931
rect 1875 927 1876 931
rect 3590 931 3596 932
rect 1870 926 1876 927
rect 1894 928 1900 929
rect 1830 924 1836 925
rect 1894 924 1895 928
rect 1899 924 1900 928
rect 127 923 133 924
rect 127 919 128 923
rect 132 922 133 923
rect 338 923 344 924
rect 338 922 339 923
rect 132 920 153 922
rect 325 920 339 922
rect 132 919 133 920
rect 127 918 133 919
rect 338 919 339 920
rect 343 919 344 923
rect 494 923 500 924
rect 494 922 495 923
rect 477 920 495 922
rect 338 918 344 919
rect 494 919 495 920
rect 499 919 500 923
rect 634 923 640 924
rect 634 922 635 923
rect 621 920 635 922
rect 494 918 500 919
rect 634 919 635 920
rect 639 919 640 923
rect 634 918 640 919
rect 686 923 692 924
rect 686 919 687 923
rect 691 922 692 923
rect 778 923 784 924
rect 691 920 721 922
rect 691 919 692 920
rect 686 918 692 919
rect 778 919 779 923
rect 783 922 784 923
rect 959 923 965 924
rect 783 920 857 922
rect 783 919 784 920
rect 778 918 784 919
rect 959 919 960 923
rect 964 922 965 923
rect 1042 923 1048 924
rect 964 920 993 922
rect 964 919 965 920
rect 959 918 965 919
rect 1042 919 1043 923
rect 1047 922 1048 923
rect 1170 923 1176 924
rect 1047 920 1121 922
rect 1047 919 1048 920
rect 1042 918 1048 919
rect 1170 919 1171 923
rect 1175 922 1176 923
rect 1402 923 1408 924
rect 1402 922 1403 923
rect 1175 920 1241 922
rect 1397 920 1403 922
rect 1175 919 1176 920
rect 1170 918 1176 919
rect 1402 919 1403 920
rect 1407 919 1408 923
rect 1506 923 1512 924
rect 1506 922 1507 923
rect 1501 920 1507 922
rect 1402 918 1408 919
rect 1506 919 1507 920
rect 1511 919 1512 923
rect 1610 923 1616 924
rect 1610 922 1611 923
rect 1605 920 1611 922
rect 1506 918 1512 919
rect 1610 919 1611 920
rect 1615 919 1616 923
rect 1722 923 1728 924
rect 1894 923 1900 924
rect 1974 928 1980 929
rect 1974 924 1975 928
rect 1979 924 1980 928
rect 1974 923 1980 924
rect 2070 928 2076 929
rect 2070 924 2071 928
rect 2075 924 2076 928
rect 2070 923 2076 924
rect 2190 928 2196 929
rect 2190 924 2191 928
rect 2195 924 2196 928
rect 2190 923 2196 924
rect 2326 928 2332 929
rect 2326 924 2327 928
rect 2331 924 2332 928
rect 2326 923 2332 924
rect 2470 928 2476 929
rect 2470 924 2471 928
rect 2475 924 2476 928
rect 2470 923 2476 924
rect 2622 928 2628 929
rect 2622 924 2623 928
rect 2627 924 2628 928
rect 2622 923 2628 924
rect 2782 928 2788 929
rect 2782 924 2783 928
rect 2787 924 2788 928
rect 2782 923 2788 924
rect 2958 928 2964 929
rect 2958 924 2959 928
rect 2963 924 2964 928
rect 2958 923 2964 924
rect 3142 928 3148 929
rect 3142 924 3143 928
rect 3147 924 3148 928
rect 3142 923 3148 924
rect 3334 928 3340 929
rect 3334 924 3335 928
rect 3339 924 3340 928
rect 3334 923 3340 924
rect 3502 928 3508 929
rect 3502 924 3503 928
rect 3507 924 3508 928
rect 3590 927 3591 931
rect 3595 927 3596 931
rect 3590 926 3596 927
rect 3502 923 3508 924
rect 1722 922 1723 923
rect 1717 920 1723 922
rect 1610 918 1616 919
rect 1722 919 1723 920
rect 1727 919 1728 923
rect 1744 920 1761 922
rect 1722 918 1728 919
rect 1742 919 1748 920
rect 1742 915 1743 919
rect 1747 915 1748 919
rect 1742 914 1748 915
rect 110 912 116 913
rect 110 908 111 912
rect 115 908 116 912
rect 110 907 116 908
rect 1830 912 1836 913
rect 1830 908 1831 912
rect 1835 908 1836 912
rect 1830 907 1836 908
rect 2310 911 2316 912
rect 2310 907 2311 911
rect 2315 910 2316 911
rect 2343 911 2349 912
rect 2343 910 2344 911
rect 2315 908 2344 910
rect 2315 907 2316 908
rect 2310 906 2316 907
rect 2343 907 2344 908
rect 2348 907 2349 911
rect 2343 906 2349 907
rect 2878 911 2884 912
rect 2878 907 2879 911
rect 2883 910 2884 911
rect 2975 911 2981 912
rect 2975 910 2976 911
rect 2883 908 2976 910
rect 2883 907 2884 908
rect 2878 906 2884 907
rect 2975 907 2976 908
rect 2980 907 2981 911
rect 2975 906 2981 907
rect 142 894 148 895
rect 142 890 143 894
rect 147 890 148 894
rect 142 889 148 890
rect 270 894 276 895
rect 270 890 271 894
rect 275 890 276 894
rect 270 889 276 890
rect 422 894 428 895
rect 422 890 423 894
rect 427 890 428 894
rect 422 889 428 890
rect 566 894 572 895
rect 566 890 567 894
rect 571 890 572 894
rect 566 889 572 890
rect 710 894 716 895
rect 710 890 711 894
rect 715 890 716 894
rect 710 889 716 890
rect 846 894 852 895
rect 846 890 847 894
rect 851 890 852 894
rect 846 889 852 890
rect 982 894 988 895
rect 982 890 983 894
rect 987 890 988 894
rect 982 889 988 890
rect 1110 894 1116 895
rect 1110 890 1111 894
rect 1115 890 1116 894
rect 1110 889 1116 890
rect 1230 894 1236 895
rect 1230 890 1231 894
rect 1235 890 1236 894
rect 1230 889 1236 890
rect 1342 894 1348 895
rect 1342 890 1343 894
rect 1347 890 1348 894
rect 1342 889 1348 890
rect 1446 894 1452 895
rect 1446 890 1447 894
rect 1451 890 1452 894
rect 1446 889 1452 890
rect 1550 894 1556 895
rect 1550 890 1551 894
rect 1555 890 1556 894
rect 1550 889 1556 890
rect 1662 894 1668 895
rect 1662 890 1663 894
rect 1667 890 1668 894
rect 1662 889 1668 890
rect 1750 894 1756 895
rect 1750 890 1751 894
rect 1755 890 1756 894
rect 1750 889 1756 890
rect 135 883 141 884
rect 135 879 136 883
rect 140 882 141 883
rect 150 883 156 884
rect 150 882 151 883
rect 140 880 151 882
rect 140 879 141 880
rect 135 878 141 879
rect 150 879 151 880
rect 155 879 156 883
rect 150 878 156 879
rect 255 883 261 884
rect 255 879 256 883
rect 260 882 261 883
rect 263 883 269 884
rect 263 882 264 883
rect 260 880 264 882
rect 260 879 261 880
rect 255 878 261 879
rect 263 879 264 880
rect 268 879 269 883
rect 263 878 269 879
rect 338 883 344 884
rect 338 879 339 883
rect 343 882 344 883
rect 415 883 421 884
rect 415 882 416 883
rect 343 880 416 882
rect 343 879 344 880
rect 338 878 344 879
rect 415 879 416 880
rect 420 879 421 883
rect 415 878 421 879
rect 494 883 500 884
rect 494 879 495 883
rect 499 882 500 883
rect 559 883 565 884
rect 559 882 560 883
rect 499 880 560 882
rect 499 879 500 880
rect 494 878 500 879
rect 559 879 560 880
rect 564 879 565 883
rect 559 878 565 879
rect 703 883 709 884
rect 703 879 704 883
rect 708 882 709 883
rect 778 883 784 884
rect 778 882 779 883
rect 708 880 779 882
rect 708 879 709 880
rect 703 878 709 879
rect 778 879 779 880
rect 783 879 784 883
rect 778 878 784 879
rect 838 883 845 884
rect 838 879 839 883
rect 844 879 845 883
rect 838 878 845 879
rect 975 883 981 884
rect 975 879 976 883
rect 980 882 981 883
rect 1042 883 1048 884
rect 1042 882 1043 883
rect 980 880 1043 882
rect 980 879 981 880
rect 975 878 981 879
rect 1042 879 1043 880
rect 1047 879 1048 883
rect 1042 878 1048 879
rect 1103 883 1109 884
rect 1103 879 1104 883
rect 1108 882 1109 883
rect 1170 883 1176 884
rect 1170 882 1171 883
rect 1108 880 1171 882
rect 1108 879 1109 880
rect 1103 878 1109 879
rect 1170 879 1171 880
rect 1175 879 1176 883
rect 1170 878 1176 879
rect 1215 883 1221 884
rect 1215 879 1216 883
rect 1220 882 1221 883
rect 1223 883 1229 884
rect 1223 882 1224 883
rect 1220 880 1224 882
rect 1220 879 1221 880
rect 1215 878 1221 879
rect 1223 879 1224 880
rect 1228 879 1229 883
rect 1223 878 1229 879
rect 1335 883 1341 884
rect 1335 879 1336 883
rect 1340 882 1341 883
rect 1390 883 1396 884
rect 1390 882 1391 883
rect 1340 880 1391 882
rect 1340 879 1341 880
rect 1335 878 1341 879
rect 1390 879 1391 880
rect 1395 879 1396 883
rect 1390 878 1396 879
rect 1402 883 1408 884
rect 1402 879 1403 883
rect 1407 882 1408 883
rect 1439 883 1445 884
rect 1439 882 1440 883
rect 1407 880 1440 882
rect 1407 879 1408 880
rect 1402 878 1408 879
rect 1439 879 1440 880
rect 1444 879 1445 883
rect 1439 878 1445 879
rect 1506 883 1512 884
rect 1506 879 1507 883
rect 1511 882 1512 883
rect 1543 883 1549 884
rect 1543 882 1544 883
rect 1511 880 1544 882
rect 1511 879 1512 880
rect 1506 878 1512 879
rect 1543 879 1544 880
rect 1548 879 1549 883
rect 1543 878 1549 879
rect 1610 883 1616 884
rect 1610 879 1611 883
rect 1615 882 1616 883
rect 1655 883 1661 884
rect 1655 882 1656 883
rect 1615 880 1656 882
rect 1615 879 1616 880
rect 1610 878 1616 879
rect 1655 879 1656 880
rect 1660 879 1661 883
rect 1655 878 1661 879
rect 1722 883 1728 884
rect 1722 879 1723 883
rect 1727 882 1728 883
rect 1743 883 1749 884
rect 1743 882 1744 883
rect 1727 880 1744 882
rect 1727 879 1728 880
rect 1722 878 1728 879
rect 1743 879 1744 880
rect 1748 879 1749 883
rect 1743 878 1749 879
rect 1646 875 1652 876
rect 1646 874 1647 875
rect 1459 872 1647 874
rect 135 867 141 868
rect 135 863 136 867
rect 140 866 141 867
rect 202 867 208 868
rect 202 866 203 867
rect 140 864 203 866
rect 140 863 141 864
rect 135 862 141 863
rect 202 863 203 864
rect 207 863 208 867
rect 202 862 208 863
rect 239 867 245 868
rect 239 863 240 867
rect 244 866 245 867
rect 258 867 264 868
rect 258 866 259 867
rect 244 864 259 866
rect 244 863 245 864
rect 239 862 245 863
rect 258 863 259 864
rect 263 863 264 867
rect 258 862 264 863
rect 366 867 372 868
rect 366 863 367 867
rect 371 866 372 867
rect 375 867 381 868
rect 375 866 376 867
rect 371 864 376 866
rect 371 863 372 864
rect 366 862 372 863
rect 375 863 376 864
rect 380 863 381 867
rect 375 862 381 863
rect 434 867 440 868
rect 434 863 435 867
rect 439 866 440 867
rect 511 867 517 868
rect 511 866 512 867
rect 439 864 512 866
rect 439 863 440 864
rect 434 862 440 863
rect 511 863 512 864
rect 516 863 517 867
rect 511 862 517 863
rect 634 867 640 868
rect 634 863 635 867
rect 639 866 640 867
rect 655 867 661 868
rect 655 866 656 867
rect 639 864 656 866
rect 639 863 640 864
rect 634 862 640 863
rect 655 863 656 864
rect 660 863 661 867
rect 655 862 661 863
rect 751 867 757 868
rect 751 863 752 867
rect 756 866 757 867
rect 807 867 813 868
rect 807 866 808 867
rect 756 864 808 866
rect 756 863 757 864
rect 751 862 757 863
rect 807 863 808 864
rect 812 863 813 867
rect 807 862 813 863
rect 951 867 957 868
rect 951 863 952 867
rect 956 866 957 867
rect 959 867 965 868
rect 959 866 960 867
rect 956 864 960 866
rect 956 863 957 864
rect 951 862 957 863
rect 959 863 960 864
rect 964 863 965 867
rect 959 862 965 863
rect 1010 867 1016 868
rect 1010 863 1011 867
rect 1015 866 1016 867
rect 1095 867 1101 868
rect 1095 866 1096 867
rect 1015 864 1096 866
rect 1015 863 1016 864
rect 1010 862 1016 863
rect 1095 863 1096 864
rect 1100 863 1101 867
rect 1095 862 1101 863
rect 1154 867 1160 868
rect 1154 863 1155 867
rect 1159 866 1160 867
rect 1239 867 1245 868
rect 1239 866 1240 867
rect 1159 864 1240 866
rect 1159 863 1160 864
rect 1154 862 1160 863
rect 1239 863 1240 864
rect 1244 863 1245 867
rect 1239 862 1245 863
rect 1375 867 1381 868
rect 1375 863 1376 867
rect 1380 866 1381 867
rect 1459 866 1461 872
rect 1646 871 1647 872
rect 1651 871 1652 875
rect 1646 870 1652 871
rect 1918 872 1924 873
rect 1870 869 1876 870
rect 1380 864 1461 866
rect 1503 867 1509 868
rect 1380 863 1381 864
rect 1375 862 1381 863
rect 1503 863 1504 867
rect 1508 866 1509 867
rect 1518 867 1524 868
rect 1518 866 1519 867
rect 1508 864 1519 866
rect 1508 863 1509 864
rect 1503 862 1509 863
rect 1518 863 1519 864
rect 1523 863 1524 867
rect 1518 862 1524 863
rect 1562 867 1568 868
rect 1562 863 1563 867
rect 1567 866 1568 867
rect 1631 867 1637 868
rect 1631 866 1632 867
rect 1567 864 1632 866
rect 1567 863 1568 864
rect 1562 862 1568 863
rect 1631 863 1632 864
rect 1636 863 1637 867
rect 1631 862 1637 863
rect 1742 867 1749 868
rect 1742 863 1743 867
rect 1748 863 1749 867
rect 1870 865 1871 869
rect 1875 865 1876 869
rect 1918 868 1919 872
rect 1923 868 1924 872
rect 1918 867 1924 868
rect 2094 872 2100 873
rect 2094 868 2095 872
rect 2099 868 2100 872
rect 2094 867 2100 868
rect 2270 872 2276 873
rect 2270 868 2271 872
rect 2275 868 2276 872
rect 2270 867 2276 868
rect 2454 872 2460 873
rect 2454 868 2455 872
rect 2459 868 2460 872
rect 2454 867 2460 868
rect 2654 872 2660 873
rect 2654 868 2655 872
rect 2659 868 2660 872
rect 2654 867 2660 868
rect 2862 872 2868 873
rect 2862 868 2863 872
rect 2867 868 2868 872
rect 2862 867 2868 868
rect 3078 872 3084 873
rect 3078 868 3079 872
rect 3083 868 3084 872
rect 3078 867 3084 868
rect 3302 872 3308 873
rect 3302 868 3303 872
rect 3307 868 3308 872
rect 3302 867 3308 868
rect 3502 872 3508 873
rect 3502 868 3503 872
rect 3507 868 3508 872
rect 3502 867 3508 868
rect 3590 869 3596 870
rect 1870 864 1876 865
rect 3590 865 3591 869
rect 3595 865 3596 869
rect 3590 864 3596 865
rect 1742 862 1749 863
rect 1903 863 1909 864
rect 1903 859 1904 863
rect 1908 862 1909 863
rect 1986 863 1992 864
rect 1908 860 1937 862
rect 1908 859 1909 860
rect 142 858 148 859
rect 142 854 143 858
rect 147 854 148 858
rect 142 853 148 854
rect 246 858 252 859
rect 246 854 247 858
rect 251 854 252 858
rect 246 853 252 854
rect 382 858 388 859
rect 382 854 383 858
rect 387 854 388 858
rect 382 853 388 854
rect 518 858 524 859
rect 518 854 519 858
rect 523 854 524 858
rect 518 853 524 854
rect 662 858 668 859
rect 662 854 663 858
rect 667 854 668 858
rect 662 853 668 854
rect 814 858 820 859
rect 814 854 815 858
rect 819 854 820 858
rect 814 853 820 854
rect 958 858 964 859
rect 958 854 959 858
rect 963 854 964 858
rect 958 853 964 854
rect 1102 858 1108 859
rect 1102 854 1103 858
rect 1107 854 1108 858
rect 1102 853 1108 854
rect 1246 858 1252 859
rect 1246 854 1247 858
rect 1251 854 1252 858
rect 1246 853 1252 854
rect 1382 858 1388 859
rect 1382 854 1383 858
rect 1387 854 1388 858
rect 1382 853 1388 854
rect 1510 858 1516 859
rect 1510 854 1511 858
rect 1515 854 1516 858
rect 1510 853 1516 854
rect 1638 858 1644 859
rect 1638 854 1639 858
rect 1643 854 1644 858
rect 1638 853 1644 854
rect 1750 858 1756 859
rect 1903 858 1909 859
rect 1986 859 1987 863
rect 1991 862 1992 863
rect 2167 863 2173 864
rect 1991 860 2113 862
rect 1991 859 1992 860
rect 1986 858 1992 859
rect 2167 859 2168 863
rect 2172 862 2173 863
rect 2551 863 2557 864
rect 2551 862 2552 863
rect 2172 860 2289 862
rect 2517 860 2552 862
rect 2172 859 2173 860
rect 2167 858 2173 859
rect 2551 859 2552 860
rect 2556 859 2557 863
rect 2551 858 2557 859
rect 2559 863 2565 864
rect 2559 859 2560 863
rect 2564 862 2565 863
rect 2722 863 2728 864
rect 2564 860 2673 862
rect 2564 859 2565 860
rect 2559 858 2565 859
rect 2722 859 2723 863
rect 2727 862 2728 863
rect 2930 863 2936 864
rect 2727 860 2881 862
rect 2727 859 2728 860
rect 2722 858 2728 859
rect 2930 859 2931 863
rect 2935 862 2936 863
rect 3194 863 3200 864
rect 2935 860 3097 862
rect 2935 859 2936 860
rect 2930 858 2936 859
rect 3194 859 3195 863
rect 3199 862 3200 863
rect 3495 863 3501 864
rect 3199 860 3321 862
rect 3199 859 3200 860
rect 3194 858 3200 859
rect 3495 859 3496 863
rect 3500 862 3501 863
rect 3500 860 3521 862
rect 3500 859 3501 860
rect 3495 858 3501 859
rect 1750 854 1751 858
rect 1755 854 1756 858
rect 1750 853 1756 854
rect 1870 852 1876 853
rect 1870 848 1871 852
rect 1875 848 1876 852
rect 1870 847 1876 848
rect 3590 852 3596 853
rect 3590 848 3591 852
rect 3595 848 3596 852
rect 3590 847 3596 848
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 1830 840 1836 841
rect 1830 836 1831 840
rect 1835 836 1836 840
rect 1830 835 1836 836
rect 1926 834 1932 835
rect 150 831 156 832
rect 150 827 151 831
rect 155 827 156 831
rect 150 826 156 827
rect 202 831 208 832
rect 202 827 203 831
rect 207 830 208 831
rect 434 831 440 832
rect 207 828 257 830
rect 207 827 208 828
rect 202 826 208 827
rect 434 827 435 831
rect 439 827 440 831
rect 434 826 440 827
rect 526 831 532 832
rect 526 827 527 831
rect 531 827 532 831
rect 751 831 757 832
rect 751 830 752 831
rect 717 828 752 830
rect 526 826 532 827
rect 751 827 752 828
rect 756 827 757 831
rect 751 826 757 827
rect 838 831 844 832
rect 838 827 839 831
rect 843 827 844 831
rect 838 826 844 827
rect 1010 831 1016 832
rect 1010 827 1011 831
rect 1015 827 1016 831
rect 1010 826 1016 827
rect 1154 831 1160 832
rect 1154 827 1155 831
rect 1159 827 1160 831
rect 1154 826 1160 827
rect 1390 831 1396 832
rect 1390 827 1391 831
rect 1395 827 1396 831
rect 1390 826 1396 827
rect 1562 831 1568 832
rect 1562 827 1563 831
rect 1567 827 1568 831
rect 1562 826 1568 827
rect 1646 831 1652 832
rect 1646 827 1647 831
rect 1651 827 1652 831
rect 1887 831 1893 832
rect 1887 830 1888 831
rect 1805 828 1888 830
rect 1646 826 1652 827
rect 1887 827 1888 828
rect 1892 827 1893 831
rect 1926 830 1927 834
rect 1931 830 1932 834
rect 1926 829 1932 830
rect 2102 834 2108 835
rect 2102 830 2103 834
rect 2107 830 2108 834
rect 2102 829 2108 830
rect 2278 834 2284 835
rect 2278 830 2279 834
rect 2283 830 2284 834
rect 2278 829 2284 830
rect 2462 834 2468 835
rect 2462 830 2463 834
rect 2467 830 2468 834
rect 2462 829 2468 830
rect 2662 834 2668 835
rect 2662 830 2663 834
rect 2667 830 2668 834
rect 2662 829 2668 830
rect 2870 834 2876 835
rect 2870 830 2871 834
rect 2875 830 2876 834
rect 2870 829 2876 830
rect 3086 834 3092 835
rect 3086 830 3087 834
rect 3091 830 3092 834
rect 3086 829 3092 830
rect 3310 834 3316 835
rect 3310 830 3311 834
rect 3315 830 3316 834
rect 3310 829 3316 830
rect 3510 834 3516 835
rect 3510 830 3511 834
rect 3515 830 3516 834
rect 3510 829 3516 830
rect 1887 826 1893 827
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 1830 823 1836 824
rect 110 818 116 819
rect 134 820 140 821
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 238 820 244 821
rect 238 816 239 820
rect 243 816 244 820
rect 238 815 244 816
rect 374 820 380 821
rect 374 816 375 820
rect 379 816 380 820
rect 374 815 380 816
rect 510 820 516 821
rect 510 816 511 820
rect 515 816 516 820
rect 510 815 516 816
rect 654 820 660 821
rect 654 816 655 820
rect 659 816 660 820
rect 654 815 660 816
rect 806 820 812 821
rect 806 816 807 820
rect 811 816 812 820
rect 806 815 812 816
rect 950 820 956 821
rect 950 816 951 820
rect 955 816 956 820
rect 950 815 956 816
rect 1094 820 1100 821
rect 1094 816 1095 820
rect 1099 816 1100 820
rect 1094 815 1100 816
rect 1238 820 1244 821
rect 1238 816 1239 820
rect 1243 816 1244 820
rect 1238 815 1244 816
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1502 820 1508 821
rect 1502 816 1503 820
rect 1507 816 1508 820
rect 1502 815 1508 816
rect 1630 820 1636 821
rect 1630 816 1631 820
rect 1635 816 1636 820
rect 1630 815 1636 816
rect 1742 820 1748 821
rect 1742 816 1743 820
rect 1747 816 1748 820
rect 1830 819 1831 823
rect 1835 819 1836 823
rect 1830 818 1836 819
rect 1919 823 1925 824
rect 1919 819 1920 823
rect 1924 822 1925 823
rect 1986 823 1992 824
rect 1986 822 1987 823
rect 1924 820 1987 822
rect 1924 819 1925 820
rect 1919 818 1925 819
rect 1986 819 1987 820
rect 1991 819 1992 823
rect 1986 818 1992 819
rect 2095 823 2101 824
rect 2095 819 2096 823
rect 2100 822 2101 823
rect 2167 823 2173 824
rect 2167 822 2168 823
rect 2100 820 2168 822
rect 2100 819 2101 820
rect 2095 818 2101 819
rect 2167 819 2168 820
rect 2172 819 2173 823
rect 2167 818 2173 819
rect 2271 823 2277 824
rect 2271 819 2272 823
rect 2276 822 2277 823
rect 2310 823 2316 824
rect 2310 822 2311 823
rect 2276 820 2311 822
rect 2276 819 2277 820
rect 2271 818 2277 819
rect 2310 819 2311 820
rect 2315 819 2316 823
rect 2310 818 2316 819
rect 2455 823 2461 824
rect 2455 819 2456 823
rect 2460 822 2461 823
rect 2559 823 2565 824
rect 2559 822 2560 823
rect 2460 820 2560 822
rect 2460 819 2461 820
rect 2455 818 2461 819
rect 2559 819 2560 820
rect 2564 819 2565 823
rect 2559 818 2565 819
rect 2655 823 2661 824
rect 2655 819 2656 823
rect 2660 822 2661 823
rect 2722 823 2728 824
rect 2722 822 2723 823
rect 2660 820 2723 822
rect 2660 819 2661 820
rect 2655 818 2661 819
rect 2722 819 2723 820
rect 2727 819 2728 823
rect 2722 818 2728 819
rect 2863 823 2869 824
rect 2863 819 2864 823
rect 2868 822 2869 823
rect 2878 823 2884 824
rect 2878 822 2879 823
rect 2868 820 2879 822
rect 2868 819 2869 820
rect 2863 818 2869 819
rect 2878 819 2879 820
rect 2883 819 2884 823
rect 2878 818 2884 819
rect 3079 823 3085 824
rect 3079 819 3080 823
rect 3084 822 3085 823
rect 3194 823 3200 824
rect 3194 822 3195 823
rect 3084 820 3195 822
rect 3084 819 3085 820
rect 3079 818 3085 819
rect 3194 819 3195 820
rect 3199 819 3200 823
rect 3194 818 3200 819
rect 3202 823 3208 824
rect 3202 819 3203 823
rect 3207 822 3208 823
rect 3303 823 3309 824
rect 3303 822 3304 823
rect 3207 820 3304 822
rect 3207 819 3208 820
rect 3202 818 3208 819
rect 3303 819 3304 820
rect 3308 819 3309 823
rect 3303 818 3309 819
rect 3503 823 3509 824
rect 3503 819 3504 823
rect 3508 822 3509 823
rect 3518 823 3524 824
rect 3518 822 3519 823
rect 3508 820 3519 822
rect 3508 819 3509 820
rect 3503 818 3509 819
rect 3518 819 3519 820
rect 3523 819 3524 823
rect 3518 818 3524 819
rect 1742 815 1748 816
rect 1895 811 1901 812
rect 1895 807 1896 811
rect 1900 810 1901 811
rect 1903 811 1909 812
rect 1903 810 1904 811
rect 1900 808 1904 810
rect 1900 807 1901 808
rect 1895 806 1901 807
rect 1903 807 1904 808
rect 1908 807 1909 811
rect 1903 806 1909 807
rect 1954 811 1960 812
rect 1954 807 1955 811
rect 1959 810 1960 811
rect 2007 811 2013 812
rect 2007 810 2008 811
rect 1959 808 2008 810
rect 1959 807 1960 808
rect 1954 806 1960 807
rect 2007 807 2008 808
rect 2012 807 2013 811
rect 2007 806 2013 807
rect 2066 811 2072 812
rect 2066 807 2067 811
rect 2071 810 2072 811
rect 2159 811 2165 812
rect 2159 810 2160 811
rect 2071 808 2160 810
rect 2071 807 2072 808
rect 2066 806 2072 807
rect 2159 807 2160 808
rect 2164 807 2165 811
rect 2159 806 2165 807
rect 2218 811 2224 812
rect 2218 807 2219 811
rect 2223 810 2224 811
rect 2319 811 2325 812
rect 2319 810 2320 811
rect 2223 808 2320 810
rect 2223 807 2224 808
rect 2218 806 2224 807
rect 2319 807 2320 808
rect 2324 807 2325 811
rect 2319 806 2325 807
rect 2378 811 2384 812
rect 2378 807 2379 811
rect 2383 810 2384 811
rect 2479 811 2485 812
rect 2479 810 2480 811
rect 2383 808 2480 810
rect 2383 807 2384 808
rect 2378 806 2384 807
rect 2479 807 2480 808
rect 2484 807 2485 811
rect 2479 806 2485 807
rect 2551 811 2557 812
rect 2551 807 2552 811
rect 2556 810 2557 811
rect 2639 811 2645 812
rect 2639 810 2640 811
rect 2556 808 2640 810
rect 2556 807 2557 808
rect 2551 806 2557 807
rect 2639 807 2640 808
rect 2644 807 2645 811
rect 2639 806 2645 807
rect 2799 811 2805 812
rect 2799 807 2800 811
rect 2804 810 2805 811
rect 2930 811 2936 812
rect 2930 810 2931 811
rect 2804 808 2931 810
rect 2804 807 2805 808
rect 2799 806 2805 807
rect 2930 807 2931 808
rect 2935 807 2936 811
rect 2930 806 2936 807
rect 2951 811 2957 812
rect 2951 807 2952 811
rect 2956 810 2957 811
rect 2978 811 2984 812
rect 2978 810 2979 811
rect 2956 808 2979 810
rect 2956 807 2957 808
rect 2951 806 2957 807
rect 2978 807 2979 808
rect 2983 807 2984 811
rect 2978 806 2984 807
rect 3010 811 3016 812
rect 3010 807 3011 811
rect 3015 810 3016 811
rect 3095 811 3101 812
rect 3095 810 3096 811
rect 3015 808 3096 810
rect 3015 807 3016 808
rect 3010 806 3016 807
rect 3095 807 3096 808
rect 3100 807 3101 811
rect 3095 806 3101 807
rect 3154 811 3160 812
rect 3154 807 3155 811
rect 3159 810 3160 811
rect 3239 811 3245 812
rect 3239 810 3240 811
rect 3159 808 3240 810
rect 3159 807 3160 808
rect 3154 806 3160 807
rect 3239 807 3240 808
rect 3244 807 3245 811
rect 3239 806 3245 807
rect 3298 811 3304 812
rect 3298 807 3299 811
rect 3303 810 3304 811
rect 3383 811 3389 812
rect 3383 810 3384 811
rect 3303 808 3384 810
rect 3303 807 3304 808
rect 3298 806 3304 807
rect 3383 807 3384 808
rect 3388 807 3389 811
rect 3383 806 3389 807
rect 3495 811 3501 812
rect 3495 807 3496 811
rect 3500 810 3501 811
rect 3503 811 3509 812
rect 3503 810 3504 811
rect 3500 808 3504 810
rect 3500 807 3501 808
rect 3495 806 3501 807
rect 3503 807 3504 808
rect 3508 807 3509 811
rect 3503 806 3509 807
rect 1158 803 1164 804
rect 1158 799 1159 803
rect 1163 802 1164 803
rect 1255 803 1261 804
rect 1255 802 1256 803
rect 1163 800 1256 802
rect 1163 799 1164 800
rect 1158 798 1164 799
rect 1255 799 1256 800
rect 1260 799 1261 803
rect 1255 798 1261 799
rect 1902 802 1908 803
rect 1902 798 1903 802
rect 1907 798 1908 802
rect 1902 797 1908 798
rect 2014 802 2020 803
rect 2014 798 2015 802
rect 2019 798 2020 802
rect 2014 797 2020 798
rect 2166 802 2172 803
rect 2166 798 2167 802
rect 2171 798 2172 802
rect 2166 797 2172 798
rect 2326 802 2332 803
rect 2326 798 2327 802
rect 2331 798 2332 802
rect 2326 797 2332 798
rect 2486 802 2492 803
rect 2486 798 2487 802
rect 2491 798 2492 802
rect 2486 797 2492 798
rect 2646 802 2652 803
rect 2646 798 2647 802
rect 2651 798 2652 802
rect 2646 797 2652 798
rect 2806 802 2812 803
rect 2806 798 2807 802
rect 2811 798 2812 802
rect 2806 797 2812 798
rect 2958 802 2964 803
rect 2958 798 2959 802
rect 2963 798 2964 802
rect 2958 797 2964 798
rect 3102 802 3108 803
rect 3102 798 3103 802
rect 3107 798 3108 802
rect 3102 797 3108 798
rect 3246 802 3252 803
rect 3246 798 3247 802
rect 3251 798 3252 802
rect 3246 797 3252 798
rect 3390 802 3396 803
rect 3390 798 3391 802
rect 3395 798 3396 802
rect 3390 797 3396 798
rect 3510 802 3516 803
rect 3510 798 3511 802
rect 3515 798 3516 802
rect 3510 797 3516 798
rect 1870 784 1876 785
rect 1870 780 1871 784
rect 1875 780 1876 784
rect 1870 779 1876 780
rect 3590 784 3596 785
rect 3590 780 3591 784
rect 3595 780 3596 784
rect 3590 779 3596 780
rect 1954 775 1960 776
rect 1954 771 1955 775
rect 1959 771 1960 775
rect 1954 770 1960 771
rect 2066 775 2072 776
rect 2066 771 2067 775
rect 2071 771 2072 775
rect 2066 770 2072 771
rect 2218 775 2224 776
rect 2218 771 2219 775
rect 2223 771 2224 775
rect 2218 770 2224 771
rect 2378 775 2384 776
rect 2378 771 2379 775
rect 2383 771 2384 775
rect 2378 770 2384 771
rect 2698 775 2704 776
rect 2698 771 2699 775
rect 2703 771 2704 775
rect 2870 775 2876 776
rect 2870 774 2871 775
rect 2861 772 2871 774
rect 2698 770 2704 771
rect 2870 771 2871 772
rect 2875 771 2876 775
rect 2870 770 2876 771
rect 3010 775 3016 776
rect 3010 771 3011 775
rect 3015 771 3016 775
rect 3010 770 3016 771
rect 3154 775 3160 776
rect 3154 771 3155 775
rect 3159 771 3160 775
rect 3154 770 3160 771
rect 3298 775 3304 776
rect 3298 771 3299 775
rect 3303 771 3304 775
rect 3298 770 3304 771
rect 3518 775 3524 776
rect 3518 771 3519 775
rect 3523 771 3524 775
rect 3518 770 3524 771
rect 1870 767 1876 768
rect 134 764 140 765
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 134 760 135 764
rect 139 760 140 764
rect 134 759 140 760
rect 214 764 220 765
rect 214 760 215 764
rect 219 760 220 764
rect 214 759 220 760
rect 302 764 308 765
rect 302 760 303 764
rect 307 760 308 764
rect 302 759 308 760
rect 414 764 420 765
rect 414 760 415 764
rect 419 760 420 764
rect 414 759 420 760
rect 542 764 548 765
rect 542 760 543 764
rect 547 760 548 764
rect 542 759 548 760
rect 686 764 692 765
rect 686 760 687 764
rect 691 760 692 764
rect 686 759 692 760
rect 838 764 844 765
rect 838 760 839 764
rect 843 760 844 764
rect 838 759 844 760
rect 990 764 996 765
rect 990 760 991 764
rect 995 760 996 764
rect 990 759 996 760
rect 1142 764 1148 765
rect 1142 760 1143 764
rect 1147 760 1148 764
rect 1142 759 1148 760
rect 1294 764 1300 765
rect 1294 760 1295 764
rect 1299 760 1300 764
rect 1294 759 1300 760
rect 1446 764 1452 765
rect 1446 760 1447 764
rect 1451 760 1452 764
rect 1446 759 1452 760
rect 1606 764 1612 765
rect 1606 760 1607 764
rect 1611 760 1612 764
rect 1870 763 1871 767
rect 1875 763 1876 767
rect 3590 767 3596 768
rect 1870 762 1876 763
rect 1894 764 1900 765
rect 1606 759 1612 760
rect 1830 761 1836 762
rect 110 756 116 757
rect 1830 757 1831 761
rect 1835 757 1836 761
rect 1894 760 1895 764
rect 1899 760 1900 764
rect 1894 759 1900 760
rect 2006 764 2012 765
rect 2006 760 2007 764
rect 2011 760 2012 764
rect 2006 759 2012 760
rect 2158 764 2164 765
rect 2158 760 2159 764
rect 2163 760 2164 764
rect 2158 759 2164 760
rect 2318 764 2324 765
rect 2318 760 2319 764
rect 2323 760 2324 764
rect 2318 759 2324 760
rect 2478 764 2484 765
rect 2478 760 2479 764
rect 2483 760 2484 764
rect 2478 759 2484 760
rect 2638 764 2644 765
rect 2638 760 2639 764
rect 2643 760 2644 764
rect 2638 759 2644 760
rect 2798 764 2804 765
rect 2798 760 2799 764
rect 2803 760 2804 764
rect 2798 759 2804 760
rect 2950 764 2956 765
rect 2950 760 2951 764
rect 2955 760 2956 764
rect 2950 759 2956 760
rect 3094 764 3100 765
rect 3094 760 3095 764
rect 3099 760 3100 764
rect 3094 759 3100 760
rect 3238 764 3244 765
rect 3238 760 3239 764
rect 3243 760 3244 764
rect 3238 759 3244 760
rect 3382 764 3388 765
rect 3382 760 3383 764
rect 3387 760 3388 764
rect 3382 759 3388 760
rect 3502 764 3508 765
rect 3502 760 3503 764
rect 3507 760 3508 764
rect 3590 763 3591 767
rect 3595 763 3596 767
rect 3590 762 3596 763
rect 3502 759 3508 760
rect 1830 756 1836 757
rect 202 755 208 756
rect 202 754 203 755
rect 197 752 203 754
rect 202 751 203 752
rect 207 751 208 755
rect 282 755 288 756
rect 282 754 283 755
rect 277 752 283 754
rect 202 750 208 751
rect 282 751 283 752
rect 287 751 288 755
rect 370 755 376 756
rect 370 754 371 755
rect 365 752 371 754
rect 282 750 288 751
rect 370 751 371 752
rect 375 751 376 755
rect 486 755 492 756
rect 486 754 487 755
rect 477 752 487 754
rect 370 750 376 751
rect 486 751 487 752
rect 491 751 492 755
rect 610 755 616 756
rect 610 754 611 755
rect 605 752 611 754
rect 486 750 492 751
rect 610 751 611 752
rect 615 751 616 755
rect 610 750 616 751
rect 654 755 660 756
rect 654 751 655 755
rect 659 754 660 755
rect 906 755 912 756
rect 906 754 907 755
rect 659 752 705 754
rect 901 752 907 754
rect 659 751 660 752
rect 654 750 660 751
rect 906 751 907 752
rect 911 751 912 755
rect 906 750 912 751
rect 914 755 920 756
rect 914 751 915 755
rect 919 754 920 755
rect 1058 755 1064 756
rect 919 752 1009 754
rect 919 751 920 752
rect 914 750 920 751
rect 1058 751 1059 755
rect 1063 754 1064 755
rect 1378 755 1384 756
rect 1378 754 1379 755
rect 1063 752 1161 754
rect 1357 752 1379 754
rect 1063 751 1064 752
rect 1058 750 1064 751
rect 1378 751 1379 752
rect 1383 751 1384 755
rect 1518 755 1524 756
rect 1518 754 1519 755
rect 1509 752 1519 754
rect 1378 750 1384 751
rect 1518 751 1519 752
rect 1523 751 1524 755
rect 1518 750 1524 751
rect 1530 755 1536 756
rect 1530 751 1531 755
rect 1535 754 1536 755
rect 1535 752 1625 754
rect 1535 751 1536 752
rect 1530 750 1536 751
rect 2418 747 2424 748
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 2418 743 2419 747
rect 2423 746 2424 747
rect 2495 747 2501 748
rect 2495 746 2496 747
rect 2423 744 2496 746
rect 2423 743 2424 744
rect 2418 742 2424 743
rect 2495 743 2496 744
rect 2500 743 2501 747
rect 2495 742 2501 743
rect 3374 747 3380 748
rect 3374 743 3375 747
rect 3379 746 3380 747
rect 3399 747 3405 748
rect 3399 746 3400 747
rect 3379 744 3400 746
rect 3379 743 3380 744
rect 3374 742 3380 743
rect 3399 743 3400 744
rect 3404 743 3405 747
rect 3399 742 3405 743
rect 1830 739 1836 740
rect 142 726 148 727
rect 142 722 143 726
rect 147 722 148 726
rect 142 721 148 722
rect 222 726 228 727
rect 222 722 223 726
rect 227 722 228 726
rect 222 721 228 722
rect 310 726 316 727
rect 310 722 311 726
rect 315 722 316 726
rect 310 721 316 722
rect 422 726 428 727
rect 422 722 423 726
rect 427 722 428 726
rect 422 721 428 722
rect 550 726 556 727
rect 550 722 551 726
rect 555 722 556 726
rect 550 721 556 722
rect 694 726 700 727
rect 694 722 695 726
rect 699 722 700 726
rect 694 721 700 722
rect 846 726 852 727
rect 846 722 847 726
rect 851 722 852 726
rect 846 721 852 722
rect 998 726 1004 727
rect 998 722 999 726
rect 1003 722 1004 726
rect 998 721 1004 722
rect 1150 726 1156 727
rect 1150 722 1151 726
rect 1155 722 1156 726
rect 1150 721 1156 722
rect 1302 726 1308 727
rect 1302 722 1303 726
rect 1307 722 1308 726
rect 1302 721 1308 722
rect 1454 726 1460 727
rect 1454 722 1455 726
rect 1459 722 1460 726
rect 1454 721 1460 722
rect 1614 726 1620 727
rect 1614 722 1615 726
rect 1619 722 1620 726
rect 1614 721 1620 722
rect 1966 720 1972 721
rect 1870 717 1876 718
rect 135 715 141 716
rect 135 711 136 715
rect 140 714 141 715
rect 150 715 156 716
rect 150 714 151 715
rect 140 712 151 714
rect 140 711 141 712
rect 135 710 141 711
rect 150 711 151 712
rect 155 711 156 715
rect 150 710 156 711
rect 202 715 208 716
rect 202 711 203 715
rect 207 714 208 715
rect 215 715 221 716
rect 215 714 216 715
rect 207 712 216 714
rect 207 711 208 712
rect 202 710 208 711
rect 215 711 216 712
rect 220 711 221 715
rect 215 710 221 711
rect 282 715 288 716
rect 282 711 283 715
rect 287 714 288 715
rect 303 715 309 716
rect 303 714 304 715
rect 287 712 304 714
rect 287 711 288 712
rect 282 710 288 711
rect 303 711 304 712
rect 308 711 309 715
rect 303 710 309 711
rect 415 715 421 716
rect 415 711 416 715
rect 420 714 421 715
rect 430 715 436 716
rect 430 714 431 715
rect 420 712 431 714
rect 420 711 421 712
rect 415 710 421 711
rect 430 711 431 712
rect 435 711 436 715
rect 430 710 436 711
rect 486 715 492 716
rect 486 711 487 715
rect 491 714 492 715
rect 543 715 549 716
rect 543 714 544 715
rect 491 712 544 714
rect 491 711 492 712
rect 486 710 492 711
rect 543 711 544 712
rect 548 711 549 715
rect 543 710 549 711
rect 610 715 616 716
rect 610 711 611 715
rect 615 714 616 715
rect 687 715 693 716
rect 687 714 688 715
rect 615 712 688 714
rect 615 711 616 712
rect 610 710 616 711
rect 687 711 688 712
rect 692 711 693 715
rect 687 710 693 711
rect 839 715 845 716
rect 839 711 840 715
rect 844 714 845 715
rect 914 715 920 716
rect 914 714 915 715
rect 844 712 915 714
rect 844 711 845 712
rect 839 710 845 711
rect 914 711 915 712
rect 919 711 920 715
rect 914 710 920 711
rect 991 715 997 716
rect 991 711 992 715
rect 996 714 997 715
rect 1058 715 1064 716
rect 1058 714 1059 715
rect 996 712 1059 714
rect 996 711 997 712
rect 991 710 997 711
rect 1058 711 1059 712
rect 1063 711 1064 715
rect 1058 710 1064 711
rect 1143 715 1149 716
rect 1143 711 1144 715
rect 1148 714 1149 715
rect 1158 715 1164 716
rect 1158 714 1159 715
rect 1148 712 1159 714
rect 1148 711 1149 712
rect 1143 710 1149 711
rect 1158 711 1159 712
rect 1163 711 1164 715
rect 1158 710 1164 711
rect 1295 715 1301 716
rect 1295 711 1296 715
rect 1300 714 1301 715
rect 1310 715 1316 716
rect 1310 714 1311 715
rect 1300 712 1311 714
rect 1300 711 1301 712
rect 1295 710 1301 711
rect 1310 711 1311 712
rect 1315 711 1316 715
rect 1310 710 1316 711
rect 1378 715 1384 716
rect 1378 711 1379 715
rect 1383 714 1384 715
rect 1447 715 1453 716
rect 1447 714 1448 715
rect 1383 712 1448 714
rect 1383 711 1384 712
rect 1378 710 1384 711
rect 1447 711 1448 712
rect 1452 711 1453 715
rect 1447 710 1453 711
rect 1606 715 1613 716
rect 1606 711 1607 715
rect 1612 711 1613 715
rect 1870 713 1871 717
rect 1875 713 1876 717
rect 1966 716 1967 720
rect 1971 716 1972 720
rect 1966 715 1972 716
rect 2062 720 2068 721
rect 2062 716 2063 720
rect 2067 716 2068 720
rect 2062 715 2068 716
rect 2174 720 2180 721
rect 2174 716 2175 720
rect 2179 716 2180 720
rect 2174 715 2180 716
rect 2302 720 2308 721
rect 2302 716 2303 720
rect 2307 716 2308 720
rect 2302 715 2308 716
rect 2446 720 2452 721
rect 2446 716 2447 720
rect 2451 716 2452 720
rect 2446 715 2452 716
rect 2598 720 2604 721
rect 2598 716 2599 720
rect 2603 716 2604 720
rect 2598 715 2604 716
rect 2750 720 2756 721
rect 2750 716 2751 720
rect 2755 716 2756 720
rect 2750 715 2756 716
rect 2902 720 2908 721
rect 2902 716 2903 720
rect 2907 716 2908 720
rect 2902 715 2908 716
rect 3054 720 3060 721
rect 3054 716 3055 720
rect 3059 716 3060 720
rect 3054 715 3060 716
rect 3206 720 3212 721
rect 3206 716 3207 720
rect 3211 716 3212 720
rect 3206 715 3212 716
rect 3358 720 3364 721
rect 3358 716 3359 720
rect 3363 716 3364 720
rect 3358 715 3364 716
rect 3502 720 3508 721
rect 3502 716 3503 720
rect 3507 716 3508 720
rect 3502 715 3508 716
rect 3590 717 3596 718
rect 1870 712 1876 713
rect 3590 713 3591 717
rect 3595 713 3596 717
rect 3590 712 3596 713
rect 1606 710 1613 711
rect 2034 711 2040 712
rect 2034 710 2035 711
rect 2029 708 2035 710
rect 2034 707 2035 708
rect 2039 707 2040 711
rect 2130 711 2136 712
rect 2130 710 2131 711
rect 2125 708 2131 710
rect 2034 706 2040 707
rect 2130 707 2131 708
rect 2135 707 2136 711
rect 2246 711 2252 712
rect 2246 710 2247 711
rect 2237 708 2247 710
rect 2130 706 2136 707
rect 2246 707 2247 708
rect 2251 707 2252 711
rect 2382 711 2388 712
rect 2382 710 2383 711
rect 2365 708 2383 710
rect 2246 706 2252 707
rect 2382 707 2383 708
rect 2387 707 2388 711
rect 2591 711 2597 712
rect 2591 710 2592 711
rect 2509 708 2592 710
rect 2382 706 2388 707
rect 2591 707 2592 708
rect 2596 707 2597 711
rect 2818 711 2824 712
rect 2818 710 2819 711
rect 2591 706 2597 707
rect 2606 707 2612 708
rect 2606 703 2607 707
rect 2611 706 2612 707
rect 2616 706 2618 709
rect 2813 708 2819 710
rect 2818 707 2819 708
rect 2823 707 2824 711
rect 2978 711 2984 712
rect 2818 706 2824 707
rect 2611 704 2618 706
rect 2611 703 2612 704
rect 2606 702 2612 703
rect 2735 703 2741 704
rect 1870 700 1876 701
rect 1870 696 1871 700
rect 1875 696 1876 700
rect 2735 699 2736 703
rect 2740 702 2741 703
rect 2920 702 2922 709
rect 2978 707 2979 711
rect 2983 710 2984 711
rect 3274 711 3280 712
rect 2983 708 3073 710
rect 2983 707 2984 708
rect 2978 706 2984 707
rect 3268 704 3270 709
rect 3274 707 3275 711
rect 3279 710 3280 711
rect 3495 711 3501 712
rect 3279 708 3377 710
rect 3279 707 3280 708
rect 3274 706 3280 707
rect 3495 707 3496 711
rect 3500 710 3501 711
rect 3500 708 3521 710
rect 3500 707 3501 708
rect 3495 706 3501 707
rect 2740 700 2922 702
rect 3266 703 3272 704
rect 2740 699 2741 700
rect 2735 698 2741 699
rect 3266 699 3267 703
rect 3271 699 3272 703
rect 3266 698 3272 699
rect 3590 700 3596 701
rect 223 695 229 696
rect 223 691 224 695
rect 228 694 229 695
rect 274 695 280 696
rect 274 694 275 695
rect 228 692 275 694
rect 228 691 229 692
rect 223 690 229 691
rect 274 691 275 692
rect 279 691 280 695
rect 274 690 280 691
rect 282 695 288 696
rect 282 691 283 695
rect 287 694 288 695
rect 311 695 317 696
rect 311 694 312 695
rect 287 692 312 694
rect 287 691 288 692
rect 282 690 288 691
rect 311 691 312 692
rect 316 691 317 695
rect 311 690 317 691
rect 370 695 376 696
rect 370 691 371 695
rect 375 694 376 695
rect 415 695 421 696
rect 415 694 416 695
rect 375 692 416 694
rect 375 691 376 692
rect 370 690 376 691
rect 415 691 416 692
rect 420 691 421 695
rect 415 690 421 691
rect 535 695 541 696
rect 535 691 536 695
rect 540 694 541 695
rect 602 695 608 696
rect 602 694 603 695
rect 540 692 603 694
rect 540 691 541 692
rect 535 690 541 691
rect 602 691 603 692
rect 607 691 608 695
rect 602 690 608 691
rect 671 695 677 696
rect 671 691 672 695
rect 676 694 677 695
rect 738 695 744 696
rect 738 694 739 695
rect 676 692 739 694
rect 676 691 677 692
rect 671 690 677 691
rect 738 691 739 692
rect 743 691 744 695
rect 738 690 744 691
rect 807 695 813 696
rect 807 691 808 695
rect 812 694 813 695
rect 854 695 860 696
rect 854 694 855 695
rect 812 692 855 694
rect 812 691 813 692
rect 807 690 813 691
rect 854 691 855 692
rect 859 691 860 695
rect 854 690 860 691
rect 906 695 912 696
rect 906 691 907 695
rect 911 694 912 695
rect 943 695 949 696
rect 943 694 944 695
rect 911 692 944 694
rect 911 691 912 692
rect 906 690 912 691
rect 943 691 944 692
rect 948 691 949 695
rect 943 690 949 691
rect 1079 695 1085 696
rect 1079 691 1080 695
rect 1084 694 1085 695
rect 1094 695 1100 696
rect 1094 694 1095 695
rect 1084 692 1095 694
rect 1084 691 1085 692
rect 1079 690 1085 691
rect 1094 691 1095 692
rect 1099 691 1100 695
rect 1094 690 1100 691
rect 1138 695 1144 696
rect 1138 691 1139 695
rect 1143 694 1144 695
rect 1207 695 1213 696
rect 1207 694 1208 695
rect 1143 692 1208 694
rect 1143 691 1144 692
rect 1138 690 1144 691
rect 1207 691 1208 692
rect 1212 691 1213 695
rect 1207 690 1213 691
rect 1266 695 1272 696
rect 1266 691 1267 695
rect 1271 694 1272 695
rect 1327 695 1333 696
rect 1327 694 1328 695
rect 1271 692 1328 694
rect 1271 691 1272 692
rect 1266 690 1272 691
rect 1327 691 1328 692
rect 1332 691 1333 695
rect 1327 690 1333 691
rect 1386 695 1392 696
rect 1386 691 1387 695
rect 1391 694 1392 695
rect 1447 695 1453 696
rect 1447 694 1448 695
rect 1391 692 1448 694
rect 1391 691 1392 692
rect 1386 690 1392 691
rect 1447 691 1448 692
rect 1452 691 1453 695
rect 1447 690 1453 691
rect 1506 695 1512 696
rect 1506 691 1507 695
rect 1511 694 1512 695
rect 1575 695 1581 696
rect 1870 695 1876 696
rect 3590 696 3591 700
rect 3595 696 3596 700
rect 3590 695 3596 696
rect 1575 694 1576 695
rect 1511 692 1576 694
rect 1511 691 1512 692
rect 1506 690 1512 691
rect 1575 691 1576 692
rect 1580 691 1581 695
rect 1575 690 1581 691
rect 230 686 236 687
rect 230 682 231 686
rect 235 682 236 686
rect 230 681 236 682
rect 318 686 324 687
rect 318 682 319 686
rect 323 682 324 686
rect 318 681 324 682
rect 422 686 428 687
rect 422 682 423 686
rect 427 682 428 686
rect 422 681 428 682
rect 542 686 548 687
rect 542 682 543 686
rect 547 682 548 686
rect 542 681 548 682
rect 678 686 684 687
rect 678 682 679 686
rect 683 682 684 686
rect 678 681 684 682
rect 814 686 820 687
rect 814 682 815 686
rect 819 682 820 686
rect 814 681 820 682
rect 950 686 956 687
rect 950 682 951 686
rect 955 682 956 686
rect 950 681 956 682
rect 1086 686 1092 687
rect 1086 682 1087 686
rect 1091 682 1092 686
rect 1086 681 1092 682
rect 1214 686 1220 687
rect 1214 682 1215 686
rect 1219 682 1220 686
rect 1214 681 1220 682
rect 1334 686 1340 687
rect 1334 682 1335 686
rect 1339 682 1340 686
rect 1334 681 1340 682
rect 1454 686 1460 687
rect 1454 682 1455 686
rect 1459 682 1460 686
rect 1454 681 1460 682
rect 1582 686 1588 687
rect 1582 682 1583 686
rect 1587 682 1588 686
rect 1582 681 1588 682
rect 1974 682 1980 683
rect 1974 678 1975 682
rect 1979 678 1980 682
rect 1974 677 1980 678
rect 2070 682 2076 683
rect 2070 678 2071 682
rect 2075 678 2076 682
rect 2070 677 2076 678
rect 2182 682 2188 683
rect 2182 678 2183 682
rect 2187 678 2188 682
rect 2182 677 2188 678
rect 2310 682 2316 683
rect 2310 678 2311 682
rect 2315 678 2316 682
rect 2310 677 2316 678
rect 2454 682 2460 683
rect 2454 678 2455 682
rect 2459 678 2460 682
rect 2454 677 2460 678
rect 2606 682 2612 683
rect 2606 678 2607 682
rect 2611 678 2612 682
rect 2606 677 2612 678
rect 2758 682 2764 683
rect 2758 678 2759 682
rect 2763 678 2764 682
rect 2758 677 2764 678
rect 2910 682 2916 683
rect 2910 678 2911 682
rect 2915 678 2916 682
rect 2910 677 2916 678
rect 3062 682 3068 683
rect 3062 678 3063 682
rect 3067 678 3068 682
rect 3062 677 3068 678
rect 3214 682 3220 683
rect 3214 678 3215 682
rect 3219 678 3220 682
rect 3214 677 3220 678
rect 3366 682 3372 683
rect 3366 678 3367 682
rect 3371 678 3372 682
rect 3366 677 3372 678
rect 3510 682 3516 683
rect 3510 678 3511 682
rect 3515 678 3516 682
rect 3510 677 3516 678
rect 3374 675 3380 676
rect 3374 674 3375 675
rect 3368 672 3375 674
rect 1967 671 1973 672
rect 110 668 116 669
rect 110 664 111 668
rect 115 664 116 668
rect 110 663 116 664
rect 1830 668 1836 669
rect 1830 664 1831 668
rect 1835 664 1836 668
rect 1967 667 1968 671
rect 1972 670 1973 671
rect 1982 671 1988 672
rect 1982 670 1983 671
rect 1972 668 1983 670
rect 1972 667 1973 668
rect 1967 666 1973 667
rect 1982 667 1983 668
rect 1987 667 1988 671
rect 1982 666 1988 667
rect 2034 671 2040 672
rect 2034 667 2035 671
rect 2039 670 2040 671
rect 2063 671 2069 672
rect 2063 670 2064 671
rect 2039 668 2064 670
rect 2039 667 2040 668
rect 2034 666 2040 667
rect 2063 667 2064 668
rect 2068 667 2069 671
rect 2063 666 2069 667
rect 2130 671 2136 672
rect 2130 667 2131 671
rect 2135 670 2136 671
rect 2175 671 2181 672
rect 2175 670 2176 671
rect 2135 668 2176 670
rect 2135 667 2136 668
rect 2130 666 2136 667
rect 2175 667 2176 668
rect 2180 667 2181 671
rect 2175 666 2181 667
rect 2246 671 2252 672
rect 2246 667 2247 671
rect 2251 670 2252 671
rect 2303 671 2309 672
rect 2303 670 2304 671
rect 2251 668 2304 670
rect 2251 667 2252 668
rect 2246 666 2252 667
rect 2303 667 2304 668
rect 2308 667 2309 671
rect 2303 666 2309 667
rect 2382 671 2388 672
rect 2382 667 2383 671
rect 2387 670 2388 671
rect 2447 671 2453 672
rect 2447 670 2448 671
rect 2387 668 2448 670
rect 2387 667 2388 668
rect 2382 666 2388 667
rect 2447 667 2448 668
rect 2452 667 2453 671
rect 2447 666 2453 667
rect 2591 671 2597 672
rect 2591 667 2592 671
rect 2596 670 2597 671
rect 2599 671 2605 672
rect 2599 670 2600 671
rect 2596 668 2600 670
rect 2596 667 2597 668
rect 2591 666 2597 667
rect 2599 667 2600 668
rect 2604 667 2605 671
rect 2599 666 2605 667
rect 2698 671 2704 672
rect 2698 667 2699 671
rect 2703 670 2704 671
rect 2751 671 2757 672
rect 2751 670 2752 671
rect 2703 668 2752 670
rect 2703 667 2704 668
rect 2698 666 2704 667
rect 2751 667 2752 668
rect 2756 667 2757 671
rect 2751 666 2757 667
rect 2870 671 2876 672
rect 2870 667 2871 671
rect 2875 670 2876 671
rect 2903 671 2909 672
rect 2903 670 2904 671
rect 2875 668 2904 670
rect 2875 667 2876 668
rect 2870 666 2876 667
rect 2903 667 2904 668
rect 2908 667 2909 671
rect 2903 666 2909 667
rect 3055 671 3061 672
rect 3055 667 3056 671
rect 3060 670 3061 671
rect 3126 671 3132 672
rect 3126 670 3127 671
rect 3060 668 3127 670
rect 3060 667 3061 668
rect 3055 666 3061 667
rect 3126 667 3127 668
rect 3131 667 3132 671
rect 3126 666 3132 667
rect 3207 671 3213 672
rect 3207 667 3208 671
rect 3212 670 3213 671
rect 3274 671 3280 672
rect 3274 670 3275 671
rect 3212 668 3275 670
rect 3212 667 3213 668
rect 3207 666 3213 667
rect 3274 667 3275 668
rect 3279 667 3280 671
rect 3274 666 3280 667
rect 3359 671 3365 672
rect 3359 667 3360 671
rect 3364 670 3365 671
rect 3368 670 3370 672
rect 3374 671 3375 672
rect 3379 671 3380 675
rect 3374 670 3380 671
rect 3503 671 3509 672
rect 3364 668 3370 670
rect 3364 667 3365 668
rect 3359 666 3365 667
rect 3503 667 3504 671
rect 3508 670 3509 671
rect 3518 671 3524 672
rect 3518 670 3519 671
rect 3508 668 3519 670
rect 3508 667 3509 668
rect 3503 666 3509 667
rect 3518 667 3519 668
rect 3523 667 3524 671
rect 3518 666 3524 667
rect 1830 663 1836 664
rect 282 659 288 660
rect 282 655 283 659
rect 287 655 288 659
rect 282 654 288 655
rect 370 659 376 660
rect 370 655 371 659
rect 375 655 376 659
rect 370 654 376 655
rect 430 659 436 660
rect 430 655 431 659
rect 435 655 436 659
rect 430 654 436 655
rect 550 659 556 660
rect 550 655 551 659
rect 555 655 556 659
rect 550 654 556 655
rect 602 659 608 660
rect 602 655 603 659
rect 607 658 608 659
rect 738 659 744 660
rect 607 656 689 658
rect 607 655 608 656
rect 602 654 608 655
rect 738 655 739 659
rect 743 658 744 659
rect 1138 659 1144 660
rect 743 656 825 658
rect 743 655 744 656
rect 738 654 744 655
rect 1138 655 1139 659
rect 1143 655 1144 659
rect 1138 654 1144 655
rect 1266 659 1272 660
rect 1266 655 1267 659
rect 1271 655 1272 659
rect 1266 654 1272 655
rect 1386 659 1392 660
rect 1386 655 1387 659
rect 1391 655 1392 659
rect 1386 654 1392 655
rect 1506 659 1512 660
rect 1506 655 1507 659
rect 1511 655 1512 659
rect 1506 654 1512 655
rect 1606 659 1612 660
rect 1606 655 1607 659
rect 1611 655 1612 659
rect 1606 654 1612 655
rect 2167 659 2173 660
rect 2167 655 2168 659
rect 2172 658 2173 659
rect 2190 659 2196 660
rect 2190 658 2191 659
rect 2172 656 2191 658
rect 2172 655 2173 656
rect 2167 654 2173 655
rect 2190 655 2191 656
rect 2195 655 2196 659
rect 2190 654 2196 655
rect 2226 659 2232 660
rect 2226 655 2227 659
rect 2231 658 2232 659
rect 2263 659 2269 660
rect 2263 658 2264 659
rect 2231 656 2264 658
rect 2231 655 2232 656
rect 2226 654 2232 655
rect 2263 655 2264 656
rect 2268 655 2269 659
rect 2263 654 2269 655
rect 2322 659 2328 660
rect 2322 655 2323 659
rect 2327 658 2328 659
rect 2367 659 2373 660
rect 2367 658 2368 659
rect 2327 656 2368 658
rect 2327 655 2328 656
rect 2322 654 2328 655
rect 2367 655 2368 656
rect 2372 655 2373 659
rect 2367 654 2373 655
rect 2426 659 2432 660
rect 2426 655 2427 659
rect 2431 658 2432 659
rect 2479 659 2485 660
rect 2479 658 2480 659
rect 2431 656 2480 658
rect 2431 655 2432 656
rect 2426 654 2432 655
rect 2479 655 2480 656
rect 2484 655 2485 659
rect 2479 654 2485 655
rect 2538 659 2544 660
rect 2538 655 2539 659
rect 2543 658 2544 659
rect 2599 659 2605 660
rect 2599 658 2600 659
rect 2543 656 2600 658
rect 2543 655 2544 656
rect 2538 654 2544 655
rect 2599 655 2600 656
rect 2604 655 2605 659
rect 2599 654 2605 655
rect 2727 659 2733 660
rect 2727 655 2728 659
rect 2732 658 2733 659
rect 2735 659 2741 660
rect 2735 658 2736 659
rect 2732 656 2736 658
rect 2732 655 2733 656
rect 2727 654 2733 655
rect 2735 655 2736 656
rect 2740 655 2741 659
rect 2735 654 2741 655
rect 2818 659 2824 660
rect 2818 655 2819 659
rect 2823 658 2824 659
rect 2855 659 2861 660
rect 2855 658 2856 659
rect 2823 656 2856 658
rect 2823 655 2824 656
rect 2818 654 2824 655
rect 2855 655 2856 656
rect 2860 655 2861 659
rect 2855 654 2861 655
rect 2982 659 2989 660
rect 2982 655 2983 659
rect 2988 655 2989 659
rect 2982 654 2989 655
rect 3111 659 3117 660
rect 3111 655 3112 659
rect 3116 658 3117 659
rect 3183 659 3189 660
rect 3183 658 3184 659
rect 3116 656 3184 658
rect 3116 655 3117 656
rect 3111 654 3117 655
rect 3183 655 3184 656
rect 3188 655 3189 659
rect 3183 654 3189 655
rect 3239 659 3245 660
rect 3239 655 3240 659
rect 3244 658 3245 659
rect 3266 659 3272 660
rect 3266 658 3267 659
rect 3244 656 3267 658
rect 3244 655 3245 656
rect 3239 654 3245 655
rect 3266 655 3267 656
rect 3271 655 3272 659
rect 3266 654 3272 655
rect 3298 659 3304 660
rect 3298 655 3299 659
rect 3303 658 3304 659
rect 3367 659 3373 660
rect 3367 658 3368 659
rect 3303 656 3368 658
rect 3303 655 3304 656
rect 3298 654 3304 655
rect 3367 655 3368 656
rect 3372 655 3373 659
rect 3367 654 3373 655
rect 3503 659 3509 660
rect 3503 655 3504 659
rect 3508 658 3509 659
rect 3526 659 3532 660
rect 3526 658 3527 659
rect 3508 656 3527 658
rect 3508 655 3509 656
rect 3503 654 3509 655
rect 3526 655 3527 656
rect 3531 655 3532 659
rect 3526 654 3532 655
rect 110 651 116 652
rect 110 647 111 651
rect 115 647 116 651
rect 1830 651 1836 652
rect 110 646 116 647
rect 222 648 228 649
rect 222 644 223 648
rect 227 644 228 648
rect 222 643 228 644
rect 310 648 316 649
rect 310 644 311 648
rect 315 644 316 648
rect 310 643 316 644
rect 414 648 420 649
rect 414 644 415 648
rect 419 644 420 648
rect 414 643 420 644
rect 534 648 540 649
rect 534 644 535 648
rect 539 644 540 648
rect 534 643 540 644
rect 670 648 676 649
rect 670 644 671 648
rect 675 644 676 648
rect 670 643 676 644
rect 806 648 812 649
rect 806 644 807 648
rect 811 644 812 648
rect 806 643 812 644
rect 942 648 948 649
rect 942 644 943 648
rect 947 644 948 648
rect 942 643 948 644
rect 1078 648 1084 649
rect 1078 644 1079 648
rect 1083 644 1084 648
rect 1078 643 1084 644
rect 1206 648 1212 649
rect 1206 644 1207 648
rect 1211 644 1212 648
rect 1206 643 1212 644
rect 1326 648 1332 649
rect 1326 644 1327 648
rect 1331 644 1332 648
rect 1326 643 1332 644
rect 1446 648 1452 649
rect 1446 644 1447 648
rect 1451 644 1452 648
rect 1446 643 1452 644
rect 1574 648 1580 649
rect 1574 644 1575 648
rect 1579 644 1580 648
rect 1830 647 1831 651
rect 1835 647 1836 651
rect 1830 646 1836 647
rect 2174 650 2180 651
rect 2174 646 2175 650
rect 2179 646 2180 650
rect 2174 645 2180 646
rect 2270 650 2276 651
rect 2270 646 2271 650
rect 2275 646 2276 650
rect 2270 645 2276 646
rect 2374 650 2380 651
rect 2374 646 2375 650
rect 2379 646 2380 650
rect 2374 645 2380 646
rect 2486 650 2492 651
rect 2486 646 2487 650
rect 2491 646 2492 650
rect 2486 645 2492 646
rect 2606 650 2612 651
rect 2606 646 2607 650
rect 2611 646 2612 650
rect 2606 645 2612 646
rect 2734 650 2740 651
rect 2734 646 2735 650
rect 2739 646 2740 650
rect 2734 645 2740 646
rect 2862 650 2868 651
rect 2862 646 2863 650
rect 2867 646 2868 650
rect 2862 645 2868 646
rect 2990 650 2996 651
rect 2990 646 2991 650
rect 2995 646 2996 650
rect 2990 645 2996 646
rect 3118 650 3124 651
rect 3118 646 3119 650
rect 3123 646 3124 650
rect 3118 645 3124 646
rect 3246 650 3252 651
rect 3246 646 3247 650
rect 3251 646 3252 650
rect 3246 645 3252 646
rect 3374 650 3380 651
rect 3374 646 3375 650
rect 3379 646 3380 650
rect 3374 645 3380 646
rect 3510 650 3516 651
rect 3510 646 3511 650
rect 3515 646 3516 650
rect 3510 645 3516 646
rect 1574 643 1580 644
rect 1870 632 1876 633
rect 951 631 957 632
rect 951 627 952 631
rect 956 630 957 631
rect 959 631 965 632
rect 959 630 960 631
rect 956 628 960 630
rect 956 627 957 628
rect 951 626 957 627
rect 959 627 960 628
rect 964 627 965 631
rect 1870 628 1871 632
rect 1875 628 1876 632
rect 1870 627 1876 628
rect 3590 632 3596 633
rect 3590 628 3591 632
rect 3595 628 3596 632
rect 3590 627 3596 628
rect 959 626 965 627
rect 2226 623 2232 624
rect 2226 619 2227 623
rect 2231 619 2232 623
rect 2226 618 2232 619
rect 2322 623 2328 624
rect 2322 619 2323 623
rect 2327 619 2328 623
rect 2322 618 2328 619
rect 2426 623 2432 624
rect 2426 619 2427 623
rect 2431 619 2432 623
rect 2426 618 2432 619
rect 2538 623 2544 624
rect 2538 619 2539 623
rect 2543 619 2544 623
rect 2538 618 2544 619
rect 2786 623 2792 624
rect 2786 619 2787 623
rect 2791 619 2792 623
rect 2982 623 2988 624
rect 2982 622 2983 623
rect 2917 620 2983 622
rect 2786 618 2792 619
rect 2982 619 2983 620
rect 2987 619 2988 623
rect 2982 618 2988 619
rect 3042 623 3048 624
rect 3042 619 3043 623
rect 3047 619 3048 623
rect 3042 618 3048 619
rect 3126 623 3132 624
rect 3126 619 3127 623
rect 3131 619 3132 623
rect 3126 618 3132 619
rect 3298 623 3304 624
rect 3298 619 3299 623
rect 3303 619 3304 623
rect 3298 618 3304 619
rect 3426 623 3432 624
rect 3426 619 3427 623
rect 3431 619 3432 623
rect 3426 618 3432 619
rect 3518 623 3524 624
rect 3518 619 3519 623
rect 3523 619 3524 623
rect 3518 618 3524 619
rect 1870 615 1876 616
rect 1870 611 1871 615
rect 1875 611 1876 615
rect 3590 615 3596 616
rect 1870 610 1876 611
rect 2166 612 2172 613
rect 2166 608 2167 612
rect 2171 608 2172 612
rect 2166 607 2172 608
rect 2262 612 2268 613
rect 2262 608 2263 612
rect 2267 608 2268 612
rect 2262 607 2268 608
rect 2366 612 2372 613
rect 2366 608 2367 612
rect 2371 608 2372 612
rect 2366 607 2372 608
rect 2478 612 2484 613
rect 2478 608 2479 612
rect 2483 608 2484 612
rect 2478 607 2484 608
rect 2598 612 2604 613
rect 2598 608 2599 612
rect 2603 608 2604 612
rect 2598 607 2604 608
rect 2726 612 2732 613
rect 2726 608 2727 612
rect 2731 608 2732 612
rect 2726 607 2732 608
rect 2854 612 2860 613
rect 2854 608 2855 612
rect 2859 608 2860 612
rect 2854 607 2860 608
rect 2982 612 2988 613
rect 2982 608 2983 612
rect 2987 608 2988 612
rect 2982 607 2988 608
rect 3110 612 3116 613
rect 3110 608 3111 612
rect 3115 608 3116 612
rect 3110 607 3116 608
rect 3238 612 3244 613
rect 3238 608 3239 612
rect 3243 608 3244 612
rect 3238 607 3244 608
rect 3366 612 3372 613
rect 3366 608 3367 612
rect 3371 608 3372 612
rect 3366 607 3372 608
rect 3502 612 3508 613
rect 3502 608 3503 612
rect 3507 608 3508 612
rect 3590 611 3591 615
rect 3595 611 3596 615
rect 3590 610 3596 611
rect 3502 607 3508 608
rect 446 596 452 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 446 592 447 596
rect 451 592 452 596
rect 446 591 452 592
rect 526 596 532 597
rect 526 592 527 596
rect 531 592 532 596
rect 526 591 532 592
rect 606 596 612 597
rect 606 592 607 596
rect 611 592 612 596
rect 606 591 612 592
rect 686 596 692 597
rect 686 592 687 596
rect 691 592 692 596
rect 686 591 692 592
rect 774 596 780 597
rect 774 592 775 596
rect 779 592 780 596
rect 774 591 780 592
rect 870 596 876 597
rect 870 592 871 596
rect 875 592 876 596
rect 870 591 876 592
rect 958 596 964 597
rect 958 592 959 596
rect 963 592 964 596
rect 958 591 964 592
rect 1046 596 1052 597
rect 1046 592 1047 596
rect 1051 592 1052 596
rect 1046 591 1052 592
rect 1142 596 1148 597
rect 1142 592 1143 596
rect 1147 592 1148 596
rect 1142 591 1148 592
rect 1238 596 1244 597
rect 1238 592 1239 596
rect 1243 592 1244 596
rect 1238 591 1244 592
rect 1334 596 1340 597
rect 1334 592 1335 596
rect 1339 592 1340 596
rect 1334 591 1340 592
rect 1430 596 1436 597
rect 1430 592 1431 596
rect 1435 592 1436 596
rect 2538 595 2544 596
rect 1430 591 1436 592
rect 1830 593 1836 594
rect 110 588 116 589
rect 1830 589 1831 593
rect 1835 589 1836 593
rect 2538 591 2539 595
rect 2543 594 2544 595
rect 2615 595 2621 596
rect 2615 594 2616 595
rect 2543 592 2616 594
rect 2543 591 2544 592
rect 2538 590 2544 591
rect 2615 591 2616 592
rect 2620 591 2621 595
rect 2615 590 2621 591
rect 1830 588 1836 589
rect 514 587 520 588
rect 514 586 515 587
rect 509 584 515 586
rect 514 583 515 584
rect 519 583 520 587
rect 594 587 600 588
rect 594 586 595 587
rect 589 584 595 586
rect 514 582 520 583
rect 594 583 595 584
rect 599 583 600 587
rect 674 587 680 588
rect 674 586 675 587
rect 669 584 675 586
rect 594 582 600 583
rect 674 583 675 584
rect 679 583 680 587
rect 754 587 760 588
rect 754 586 755 587
rect 749 584 755 586
rect 674 582 680 583
rect 754 583 755 584
rect 759 583 760 587
rect 854 587 860 588
rect 854 586 855 587
rect 837 584 855 586
rect 754 582 760 583
rect 854 583 855 584
rect 859 583 860 587
rect 854 582 860 583
rect 862 587 868 588
rect 862 583 863 587
rect 867 586 868 587
rect 938 587 944 588
rect 867 584 889 586
rect 867 583 868 584
rect 862 582 868 583
rect 938 583 939 587
rect 943 586 944 587
rect 1114 587 1120 588
rect 1114 586 1115 587
rect 943 584 977 586
rect 1109 584 1115 586
rect 943 583 944 584
rect 938 582 944 583
rect 1114 583 1115 584
rect 1119 583 1120 587
rect 1210 587 1216 588
rect 1210 586 1211 587
rect 1205 584 1211 586
rect 1114 582 1120 583
rect 1210 583 1211 584
rect 1215 583 1216 587
rect 1306 587 1312 588
rect 1306 586 1307 587
rect 1301 584 1307 586
rect 1210 582 1216 583
rect 1306 583 1307 584
rect 1311 583 1312 587
rect 1402 587 1408 588
rect 1402 586 1403 587
rect 1397 584 1403 586
rect 1306 582 1312 583
rect 1402 583 1403 584
rect 1407 583 1408 587
rect 1402 582 1408 583
rect 1410 587 1416 588
rect 1410 583 1411 587
rect 1415 586 1416 587
rect 1415 584 1449 586
rect 1415 583 1416 584
rect 1410 582 1416 583
rect 110 576 116 577
rect 110 572 111 576
rect 115 572 116 576
rect 110 571 116 572
rect 1830 576 1836 577
rect 1830 572 1831 576
rect 1835 572 1836 576
rect 1830 571 1836 572
rect 2262 568 2268 569
rect 1870 565 1876 566
rect 1870 561 1871 565
rect 1875 561 1876 565
rect 2262 564 2263 568
rect 2267 564 2268 568
rect 2262 563 2268 564
rect 2342 568 2348 569
rect 2342 564 2343 568
rect 2347 564 2348 568
rect 2342 563 2348 564
rect 2422 568 2428 569
rect 2422 564 2423 568
rect 2427 564 2428 568
rect 2422 563 2428 564
rect 2502 568 2508 569
rect 2502 564 2503 568
rect 2507 564 2508 568
rect 2502 563 2508 564
rect 2590 568 2596 569
rect 2590 564 2591 568
rect 2595 564 2596 568
rect 2590 563 2596 564
rect 2694 568 2700 569
rect 2694 564 2695 568
rect 2699 564 2700 568
rect 2694 563 2700 564
rect 2814 568 2820 569
rect 2814 564 2815 568
rect 2819 564 2820 568
rect 2814 563 2820 564
rect 2958 568 2964 569
rect 2958 564 2959 568
rect 2963 564 2964 568
rect 2958 563 2964 564
rect 3110 568 3116 569
rect 3110 564 3111 568
rect 3115 564 3116 568
rect 3110 563 3116 564
rect 3278 568 3284 569
rect 3278 564 3279 568
rect 3283 564 3284 568
rect 3278 563 3284 564
rect 3446 568 3452 569
rect 3446 564 3447 568
rect 3451 564 3452 568
rect 3446 563 3452 564
rect 3590 565 3596 566
rect 1870 560 1876 561
rect 3590 561 3591 565
rect 3595 561 3596 565
rect 3590 560 3596 561
rect 2330 559 2336 560
rect 454 558 460 559
rect 454 554 455 558
rect 459 554 460 558
rect 454 553 460 554
rect 534 558 540 559
rect 534 554 535 558
rect 539 554 540 558
rect 534 553 540 554
rect 614 558 620 559
rect 614 554 615 558
rect 619 554 620 558
rect 614 553 620 554
rect 694 558 700 559
rect 694 554 695 558
rect 699 554 700 558
rect 694 553 700 554
rect 782 558 788 559
rect 782 554 783 558
rect 787 554 788 558
rect 782 553 788 554
rect 878 558 884 559
rect 878 554 879 558
rect 883 554 884 558
rect 878 553 884 554
rect 966 558 972 559
rect 966 554 967 558
rect 971 554 972 558
rect 966 553 972 554
rect 1054 558 1060 559
rect 1054 554 1055 558
rect 1059 554 1060 558
rect 1054 553 1060 554
rect 1150 558 1156 559
rect 1150 554 1151 558
rect 1155 554 1156 558
rect 1150 553 1156 554
rect 1246 558 1252 559
rect 1246 554 1247 558
rect 1251 554 1252 558
rect 1246 553 1252 554
rect 1342 558 1348 559
rect 1342 554 1343 558
rect 1347 554 1348 558
rect 1342 553 1348 554
rect 1438 558 1444 559
rect 2330 558 2331 559
rect 1438 554 1439 558
rect 1443 554 1444 558
rect 2325 556 2331 558
rect 2330 555 2331 556
rect 2335 555 2336 559
rect 2410 559 2416 560
rect 2410 558 2411 559
rect 2405 556 2411 558
rect 2330 554 2336 555
rect 2410 555 2411 556
rect 2415 555 2416 559
rect 2490 559 2496 560
rect 2490 558 2491 559
rect 2485 556 2491 558
rect 2410 554 2416 555
rect 2490 555 2491 556
rect 2495 555 2496 559
rect 2570 559 2576 560
rect 2570 558 2571 559
rect 2565 556 2571 558
rect 2490 554 2496 555
rect 2570 555 2571 556
rect 2575 555 2576 559
rect 2658 559 2664 560
rect 2658 558 2659 559
rect 2653 556 2659 558
rect 2570 554 2576 555
rect 2658 555 2659 556
rect 2663 555 2664 559
rect 2894 559 2900 560
rect 2894 558 2895 559
rect 2658 554 2664 555
rect 1438 553 1444 554
rect 2562 551 2568 552
rect 1870 548 1876 549
rect 447 547 453 548
rect 447 543 448 547
rect 452 546 453 547
rect 514 547 520 548
rect 452 544 510 546
rect 452 543 453 544
rect 447 542 453 543
rect 508 538 510 544
rect 514 543 515 547
rect 519 546 520 547
rect 527 547 533 548
rect 527 546 528 547
rect 519 544 528 546
rect 519 543 520 544
rect 514 542 520 543
rect 527 543 528 544
rect 532 543 533 547
rect 527 542 533 543
rect 594 547 600 548
rect 594 543 595 547
rect 599 546 600 547
rect 607 547 613 548
rect 607 546 608 547
rect 599 544 608 546
rect 599 543 600 544
rect 594 542 600 543
rect 607 543 608 544
rect 612 543 613 547
rect 607 542 613 543
rect 674 547 680 548
rect 674 543 675 547
rect 679 546 680 547
rect 687 547 693 548
rect 687 546 688 547
rect 679 544 688 546
rect 679 543 680 544
rect 674 542 680 543
rect 687 543 688 544
rect 692 543 693 547
rect 687 542 693 543
rect 754 547 760 548
rect 754 543 755 547
rect 759 546 760 547
rect 775 547 781 548
rect 775 546 776 547
rect 759 544 776 546
rect 759 543 760 544
rect 754 542 760 543
rect 775 543 776 544
rect 780 543 781 547
rect 775 542 781 543
rect 871 547 877 548
rect 871 543 872 547
rect 876 546 877 547
rect 938 547 944 548
rect 938 546 939 547
rect 876 544 939 546
rect 876 543 877 544
rect 871 542 877 543
rect 938 543 939 544
rect 943 543 944 547
rect 938 542 944 543
rect 951 547 957 548
rect 951 543 952 547
rect 956 546 957 547
rect 959 547 965 548
rect 959 546 960 547
rect 956 544 960 546
rect 956 543 957 544
rect 951 542 957 543
rect 959 543 960 544
rect 964 543 965 547
rect 959 542 965 543
rect 1047 547 1053 548
rect 1047 543 1048 547
rect 1052 546 1053 547
rect 1114 547 1120 548
rect 1052 544 1110 546
rect 1052 543 1053 544
rect 1047 542 1053 543
rect 598 539 604 540
rect 598 538 599 539
rect 508 536 599 538
rect 598 535 599 536
rect 603 535 604 539
rect 1108 538 1110 544
rect 1114 543 1115 547
rect 1119 546 1120 547
rect 1143 547 1149 548
rect 1143 546 1144 547
rect 1119 544 1144 546
rect 1119 543 1120 544
rect 1114 542 1120 543
rect 1143 543 1144 544
rect 1148 543 1149 547
rect 1143 542 1149 543
rect 1210 547 1216 548
rect 1210 543 1211 547
rect 1215 546 1216 547
rect 1239 547 1245 548
rect 1239 546 1240 547
rect 1215 544 1240 546
rect 1215 543 1216 544
rect 1210 542 1216 543
rect 1239 543 1240 544
rect 1244 543 1245 547
rect 1239 542 1245 543
rect 1306 547 1312 548
rect 1306 543 1307 547
rect 1311 546 1312 547
rect 1335 547 1341 548
rect 1335 546 1336 547
rect 1311 544 1336 546
rect 1311 543 1312 544
rect 1306 542 1312 543
rect 1335 543 1336 544
rect 1340 543 1341 547
rect 1335 542 1341 543
rect 1402 547 1408 548
rect 1402 543 1403 547
rect 1407 546 1408 547
rect 1431 547 1437 548
rect 1431 546 1432 547
rect 1407 544 1432 546
rect 1407 543 1408 544
rect 1402 542 1408 543
rect 1431 543 1432 544
rect 1436 543 1437 547
rect 1870 544 1871 548
rect 1875 544 1876 548
rect 2562 547 2563 551
rect 2567 550 2568 551
rect 2712 550 2714 557
rect 2877 556 2895 558
rect 2894 555 2895 556
rect 2899 555 2900 559
rect 3026 559 3032 560
rect 2894 554 2900 555
rect 2567 548 2714 550
rect 2754 551 2760 552
rect 2567 547 2568 548
rect 2562 546 2568 547
rect 2754 547 2755 551
rect 2759 550 2760 551
rect 2976 550 2978 557
rect 3026 555 3027 559
rect 3031 558 3032 559
rect 3183 559 3189 560
rect 3031 556 3129 558
rect 3031 555 3032 556
rect 3026 554 3032 555
rect 3183 555 3184 559
rect 3188 558 3189 559
rect 3526 559 3532 560
rect 3526 558 3527 559
rect 3188 556 3297 558
rect 3509 556 3527 558
rect 3188 555 3189 556
rect 3183 554 3189 555
rect 3526 555 3527 556
rect 3531 555 3532 559
rect 3526 554 3532 555
rect 2759 548 2978 550
rect 3590 548 3596 549
rect 2759 547 2760 548
rect 2754 546 2760 547
rect 1870 543 1876 544
rect 3590 544 3591 548
rect 3595 544 3596 548
rect 3590 543 3596 544
rect 1431 542 1437 543
rect 1286 539 1292 540
rect 1286 538 1287 539
rect 1108 536 1287 538
rect 598 534 604 535
rect 1286 535 1287 536
rect 1291 535 1292 539
rect 1286 534 1292 535
rect 862 531 868 532
rect 862 530 863 531
rect 716 528 863 530
rect 290 523 296 524
rect 290 519 291 523
rect 295 522 296 523
rect 327 523 333 524
rect 327 522 328 523
rect 295 520 328 522
rect 295 519 296 520
rect 290 518 296 519
rect 327 519 328 520
rect 332 519 333 523
rect 327 518 333 519
rect 386 523 392 524
rect 386 519 387 523
rect 391 522 392 523
rect 415 523 421 524
rect 415 522 416 523
rect 391 520 416 522
rect 391 519 392 520
rect 386 518 392 519
rect 415 519 416 520
rect 420 519 421 523
rect 415 518 421 519
rect 474 523 480 524
rect 474 519 475 523
rect 479 522 480 523
rect 503 523 509 524
rect 503 522 504 523
rect 479 520 504 522
rect 479 519 480 520
rect 474 518 480 519
rect 503 519 504 520
rect 508 519 509 523
rect 503 518 509 519
rect 562 523 568 524
rect 562 519 563 523
rect 567 522 568 523
rect 583 523 589 524
rect 583 522 584 523
rect 567 520 584 522
rect 567 519 568 520
rect 562 518 568 519
rect 583 519 584 520
rect 588 519 589 523
rect 583 518 589 519
rect 663 523 669 524
rect 663 519 664 523
rect 668 522 669 523
rect 716 522 718 528
rect 862 527 863 528
rect 867 527 868 531
rect 862 526 868 527
rect 2270 530 2276 531
rect 2270 526 2271 530
rect 2275 526 2276 530
rect 2270 525 2276 526
rect 2350 530 2356 531
rect 2350 526 2351 530
rect 2355 526 2356 530
rect 2350 525 2356 526
rect 2430 530 2436 531
rect 2430 526 2431 530
rect 2435 526 2436 530
rect 2430 525 2436 526
rect 2510 530 2516 531
rect 2510 526 2511 530
rect 2515 526 2516 530
rect 2510 525 2516 526
rect 2598 530 2604 531
rect 2598 526 2599 530
rect 2603 526 2604 530
rect 2598 525 2604 526
rect 2702 530 2708 531
rect 2702 526 2703 530
rect 2707 526 2708 530
rect 2702 525 2708 526
rect 2822 530 2828 531
rect 2822 526 2823 530
rect 2827 526 2828 530
rect 2822 525 2828 526
rect 2966 530 2972 531
rect 2966 526 2967 530
rect 2971 526 2972 530
rect 2966 525 2972 526
rect 3118 530 3124 531
rect 3118 526 3119 530
rect 3123 526 3124 530
rect 3118 525 3124 526
rect 3286 530 3292 531
rect 3286 526 3287 530
rect 3291 526 3292 530
rect 3286 525 3292 526
rect 3454 530 3460 531
rect 3454 526 3455 530
rect 3459 526 3460 530
rect 3454 525 3460 526
rect 668 520 718 522
rect 722 523 728 524
rect 668 519 669 520
rect 663 518 669 519
rect 722 519 723 523
rect 727 522 728 523
rect 743 523 749 524
rect 743 522 744 523
rect 727 520 744 522
rect 727 519 728 520
rect 722 518 728 519
rect 743 519 744 520
rect 748 519 749 523
rect 743 518 749 519
rect 831 523 837 524
rect 831 519 832 523
rect 836 522 837 523
rect 854 523 860 524
rect 854 522 855 523
rect 836 520 855 522
rect 836 519 837 520
rect 831 518 837 519
rect 854 519 855 520
rect 859 519 860 523
rect 854 518 860 519
rect 890 523 896 524
rect 890 519 891 523
rect 895 522 896 523
rect 919 523 925 524
rect 919 522 920 523
rect 895 520 920 522
rect 895 519 896 520
rect 890 518 896 519
rect 919 519 920 520
rect 924 519 925 523
rect 919 518 925 519
rect 978 523 984 524
rect 978 519 979 523
rect 983 522 984 523
rect 1007 523 1013 524
rect 1007 522 1008 523
rect 983 520 1008 522
rect 983 519 984 520
rect 978 518 984 519
rect 1007 519 1008 520
rect 1012 519 1013 523
rect 1007 518 1013 519
rect 1066 523 1072 524
rect 1066 519 1067 523
rect 1071 522 1072 523
rect 1095 523 1101 524
rect 1095 522 1096 523
rect 1071 520 1096 522
rect 1071 519 1072 520
rect 1066 518 1072 519
rect 1095 519 1096 520
rect 1100 519 1101 523
rect 1095 518 1101 519
rect 1182 523 1189 524
rect 1182 519 1183 523
rect 1188 519 1189 523
rect 1182 518 1189 519
rect 1270 523 1277 524
rect 1270 519 1271 523
rect 1276 519 1277 523
rect 1270 518 1277 519
rect 2263 519 2269 520
rect 2263 515 2264 519
rect 2268 518 2269 519
rect 2282 519 2288 520
rect 2282 518 2283 519
rect 2268 516 2283 518
rect 2268 515 2269 516
rect 334 514 340 515
rect 334 510 335 514
rect 339 510 340 514
rect 334 509 340 510
rect 422 514 428 515
rect 422 510 423 514
rect 427 510 428 514
rect 422 509 428 510
rect 510 514 516 515
rect 510 510 511 514
rect 515 510 516 514
rect 510 509 516 510
rect 590 514 596 515
rect 590 510 591 514
rect 595 510 596 514
rect 590 509 596 510
rect 670 514 676 515
rect 670 510 671 514
rect 675 510 676 514
rect 670 509 676 510
rect 750 514 756 515
rect 750 510 751 514
rect 755 510 756 514
rect 750 509 756 510
rect 838 514 844 515
rect 838 510 839 514
rect 843 510 844 514
rect 838 509 844 510
rect 926 514 932 515
rect 926 510 927 514
rect 931 510 932 514
rect 926 509 932 510
rect 1014 514 1020 515
rect 1014 510 1015 514
rect 1019 510 1020 514
rect 1014 509 1020 510
rect 1102 514 1108 515
rect 1102 510 1103 514
rect 1107 510 1108 514
rect 1102 509 1108 510
rect 1190 514 1196 515
rect 1190 510 1191 514
rect 1195 510 1196 514
rect 1190 509 1196 510
rect 1278 514 1284 515
rect 2263 514 2269 515
rect 2282 515 2283 516
rect 2287 515 2288 519
rect 2282 514 2288 515
rect 2330 519 2336 520
rect 2330 515 2331 519
rect 2335 518 2336 519
rect 2343 519 2349 520
rect 2343 518 2344 519
rect 2335 516 2344 518
rect 2335 515 2336 516
rect 2330 514 2336 515
rect 2343 515 2344 516
rect 2348 515 2349 519
rect 2343 514 2349 515
rect 2410 519 2416 520
rect 2410 515 2411 519
rect 2415 518 2416 519
rect 2423 519 2429 520
rect 2423 518 2424 519
rect 2415 516 2424 518
rect 2415 515 2416 516
rect 2410 514 2416 515
rect 2423 515 2424 516
rect 2428 515 2429 519
rect 2423 514 2429 515
rect 2490 519 2496 520
rect 2490 515 2491 519
rect 2495 518 2496 519
rect 2503 519 2509 520
rect 2503 518 2504 519
rect 2495 516 2504 518
rect 2495 515 2496 516
rect 2490 514 2496 515
rect 2503 515 2504 516
rect 2508 515 2509 519
rect 2503 514 2509 515
rect 2570 519 2576 520
rect 2570 515 2571 519
rect 2575 518 2576 519
rect 2591 519 2597 520
rect 2591 518 2592 519
rect 2575 516 2592 518
rect 2575 515 2576 516
rect 2570 514 2576 515
rect 2591 515 2592 516
rect 2596 515 2597 519
rect 2591 514 2597 515
rect 2658 519 2664 520
rect 2658 515 2659 519
rect 2663 518 2664 519
rect 2695 519 2701 520
rect 2695 518 2696 519
rect 2663 516 2696 518
rect 2663 515 2664 516
rect 2658 514 2664 515
rect 2695 515 2696 516
rect 2700 515 2701 519
rect 2695 514 2701 515
rect 2786 519 2792 520
rect 2786 515 2787 519
rect 2791 518 2792 519
rect 2815 519 2821 520
rect 2815 518 2816 519
rect 2791 516 2816 518
rect 2791 515 2792 516
rect 2786 514 2792 515
rect 2815 515 2816 516
rect 2820 515 2821 519
rect 2815 514 2821 515
rect 2894 519 2900 520
rect 2894 515 2895 519
rect 2899 518 2900 519
rect 2959 519 2965 520
rect 2959 518 2960 519
rect 2899 516 2960 518
rect 2899 515 2900 516
rect 2894 514 2900 515
rect 2959 515 2960 516
rect 2964 515 2965 519
rect 2959 514 2965 515
rect 3042 519 3048 520
rect 3042 515 3043 519
rect 3047 518 3048 519
rect 3111 519 3117 520
rect 3111 518 3112 519
rect 3047 516 3112 518
rect 3047 515 3048 516
rect 3042 514 3048 515
rect 3111 515 3112 516
rect 3116 515 3117 519
rect 3111 514 3117 515
rect 3279 519 3285 520
rect 3279 515 3280 519
rect 3284 518 3285 519
rect 3326 519 3332 520
rect 3326 518 3327 519
rect 3284 516 3327 518
rect 3284 515 3285 516
rect 3279 514 3285 515
rect 3326 515 3327 516
rect 3331 515 3332 519
rect 3326 514 3332 515
rect 3426 519 3432 520
rect 3426 515 3427 519
rect 3431 518 3432 519
rect 3447 519 3453 520
rect 3447 518 3448 519
rect 3431 516 3448 518
rect 3431 515 3432 516
rect 3426 514 3432 515
rect 3447 515 3448 516
rect 3452 515 3453 519
rect 3447 514 3453 515
rect 1278 510 1279 514
rect 1283 510 1284 514
rect 1278 509 1284 510
rect 3026 507 3032 508
rect 3026 506 3027 507
rect 2836 504 3027 506
rect 2183 499 2189 500
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 1830 496 1836 497
rect 1830 492 1831 496
rect 1835 492 1836 496
rect 2183 495 2184 499
rect 2188 498 2189 499
rect 2250 499 2256 500
rect 2250 498 2251 499
rect 2188 496 2251 498
rect 2188 495 2189 496
rect 2183 494 2189 495
rect 2250 495 2251 496
rect 2255 495 2256 499
rect 2250 494 2256 495
rect 2279 499 2285 500
rect 2279 495 2280 499
rect 2284 498 2285 499
rect 2351 499 2357 500
rect 2351 498 2352 499
rect 2284 496 2352 498
rect 2284 495 2285 496
rect 2279 494 2285 495
rect 2351 495 2352 496
rect 2356 495 2357 499
rect 2351 494 2357 495
rect 2375 499 2381 500
rect 2375 495 2376 499
rect 2380 498 2381 499
rect 2442 499 2448 500
rect 2442 498 2443 499
rect 2380 496 2443 498
rect 2380 495 2381 496
rect 2375 494 2381 495
rect 2442 495 2443 496
rect 2447 495 2448 499
rect 2442 494 2448 495
rect 2479 499 2485 500
rect 2479 495 2480 499
rect 2484 498 2485 499
rect 2562 499 2568 500
rect 2562 498 2563 499
rect 2484 496 2563 498
rect 2484 495 2485 496
rect 2479 494 2485 495
rect 2562 495 2563 496
rect 2567 495 2568 499
rect 2562 494 2568 495
rect 2575 499 2581 500
rect 2575 495 2576 499
rect 2580 498 2581 499
rect 2642 499 2648 500
rect 2642 498 2643 499
rect 2580 496 2643 498
rect 2580 495 2581 496
rect 2575 494 2581 495
rect 2642 495 2643 496
rect 2647 495 2648 499
rect 2642 494 2648 495
rect 2679 499 2685 500
rect 2679 495 2680 499
rect 2684 498 2685 499
rect 2754 499 2760 500
rect 2754 498 2755 499
rect 2684 496 2755 498
rect 2684 495 2685 496
rect 2679 494 2685 495
rect 2754 495 2755 496
rect 2759 495 2760 499
rect 2754 494 2760 495
rect 2783 499 2789 500
rect 2783 495 2784 499
rect 2788 498 2789 499
rect 2836 498 2838 504
rect 3026 503 3027 504
rect 3031 503 3032 507
rect 3026 502 3032 503
rect 2788 496 2838 498
rect 2842 499 2848 500
rect 2788 495 2789 496
rect 2783 494 2789 495
rect 2842 495 2843 499
rect 2847 498 2848 499
rect 2903 499 2909 500
rect 2903 498 2904 499
rect 2847 496 2904 498
rect 2847 495 2848 496
rect 2842 494 2848 495
rect 2903 495 2904 496
rect 2908 495 2909 499
rect 2903 494 2909 495
rect 3030 499 3037 500
rect 3030 495 3031 499
rect 3036 495 3037 499
rect 3030 494 3037 495
rect 3090 499 3096 500
rect 3090 495 3091 499
rect 3095 498 3096 499
rect 3167 499 3173 500
rect 3167 498 3168 499
rect 3095 496 3168 498
rect 3095 495 3096 496
rect 3090 494 3096 495
rect 3167 495 3168 496
rect 3172 495 3173 499
rect 3167 494 3173 495
rect 3226 499 3232 500
rect 3226 495 3227 499
rect 3231 498 3232 499
rect 3311 499 3317 500
rect 3311 498 3312 499
rect 3231 496 3312 498
rect 3231 495 3232 496
rect 3226 494 3232 495
rect 3311 495 3312 496
rect 3316 495 3317 499
rect 3311 494 3317 495
rect 3390 499 3396 500
rect 3390 495 3391 499
rect 3395 498 3396 499
rect 3463 499 3469 500
rect 3463 498 3464 499
rect 3395 496 3464 498
rect 3395 495 3396 496
rect 3390 494 3396 495
rect 3463 495 3464 496
rect 3468 495 3469 499
rect 3463 494 3469 495
rect 1830 491 1836 492
rect 2190 490 2196 491
rect 386 487 392 488
rect 386 483 387 487
rect 391 483 392 487
rect 386 482 392 483
rect 474 487 480 488
rect 474 483 475 487
rect 479 483 480 487
rect 474 482 480 483
rect 562 487 568 488
rect 562 483 563 487
rect 567 483 568 487
rect 562 482 568 483
rect 598 487 604 488
rect 598 483 599 487
rect 603 483 604 487
rect 598 482 604 483
rect 722 487 728 488
rect 722 483 723 487
rect 727 483 728 487
rect 722 482 728 483
rect 890 487 896 488
rect 890 483 891 487
rect 895 483 896 487
rect 890 482 896 483
rect 978 487 984 488
rect 978 483 979 487
rect 983 483 984 487
rect 978 482 984 483
rect 1066 487 1072 488
rect 1066 483 1067 487
rect 1071 483 1072 487
rect 1182 487 1188 488
rect 1182 486 1183 487
rect 1157 484 1183 486
rect 1066 482 1072 483
rect 1182 483 1183 484
rect 1187 483 1188 487
rect 1270 487 1276 488
rect 1270 486 1271 487
rect 1245 484 1271 486
rect 1182 482 1188 483
rect 1270 483 1271 484
rect 1275 483 1276 487
rect 1270 482 1276 483
rect 1286 487 1292 488
rect 1286 483 1287 487
rect 1291 483 1292 487
rect 2190 486 2191 490
rect 2195 486 2196 490
rect 2190 485 2196 486
rect 2286 490 2292 491
rect 2286 486 2287 490
rect 2291 486 2292 490
rect 2286 485 2292 486
rect 2382 490 2388 491
rect 2382 486 2383 490
rect 2387 486 2388 490
rect 2382 485 2388 486
rect 2486 490 2492 491
rect 2486 486 2487 490
rect 2491 486 2492 490
rect 2486 485 2492 486
rect 2582 490 2588 491
rect 2582 486 2583 490
rect 2587 486 2588 490
rect 2582 485 2588 486
rect 2686 490 2692 491
rect 2686 486 2687 490
rect 2691 486 2692 490
rect 2686 485 2692 486
rect 2790 490 2796 491
rect 2790 486 2791 490
rect 2795 486 2796 490
rect 2790 485 2796 486
rect 2910 490 2916 491
rect 2910 486 2911 490
rect 2915 486 2916 490
rect 2910 485 2916 486
rect 3038 490 3044 491
rect 3038 486 3039 490
rect 3043 486 3044 490
rect 3038 485 3044 486
rect 3174 490 3180 491
rect 3174 486 3175 490
rect 3179 486 3180 490
rect 3174 485 3180 486
rect 3318 490 3324 491
rect 3318 486 3319 490
rect 3323 486 3324 490
rect 3318 485 3324 486
rect 3470 490 3476 491
rect 3470 486 3471 490
rect 3475 486 3476 490
rect 3470 485 3476 486
rect 1286 482 1292 483
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 1830 479 1836 480
rect 110 474 116 475
rect 326 476 332 477
rect 326 472 327 476
rect 331 472 332 476
rect 326 471 332 472
rect 414 476 420 477
rect 414 472 415 476
rect 419 472 420 476
rect 414 471 420 472
rect 502 476 508 477
rect 502 472 503 476
rect 507 472 508 476
rect 502 471 508 472
rect 582 476 588 477
rect 582 472 583 476
rect 587 472 588 476
rect 582 471 588 472
rect 662 476 668 477
rect 662 472 663 476
rect 667 472 668 476
rect 662 471 668 472
rect 742 476 748 477
rect 742 472 743 476
rect 747 472 748 476
rect 742 471 748 472
rect 830 476 836 477
rect 830 472 831 476
rect 835 472 836 476
rect 830 471 836 472
rect 918 476 924 477
rect 918 472 919 476
rect 923 472 924 476
rect 918 471 924 472
rect 1006 476 1012 477
rect 1006 472 1007 476
rect 1011 472 1012 476
rect 1006 471 1012 472
rect 1094 476 1100 477
rect 1094 472 1095 476
rect 1099 472 1100 476
rect 1094 471 1100 472
rect 1182 476 1188 477
rect 1182 472 1183 476
rect 1187 472 1188 476
rect 1182 471 1188 472
rect 1270 476 1276 477
rect 1270 472 1271 476
rect 1275 472 1276 476
rect 1830 475 1831 479
rect 1835 475 1836 479
rect 1830 474 1836 475
rect 1270 471 1276 472
rect 1870 472 1876 473
rect 1870 468 1871 472
rect 1875 468 1876 472
rect 1870 467 1876 468
rect 3590 472 3596 473
rect 3590 468 3591 472
rect 3595 468 3596 472
rect 3590 467 3596 468
rect 2250 463 2256 464
rect 751 459 757 460
rect 751 455 752 459
rect 756 458 757 459
rect 759 459 765 460
rect 759 458 760 459
rect 756 456 760 458
rect 756 455 757 456
rect 751 454 757 455
rect 759 455 760 456
rect 764 455 765 459
rect 2250 459 2251 463
rect 2255 462 2256 463
rect 2351 463 2357 464
rect 2255 460 2297 462
rect 2255 459 2256 460
rect 2250 458 2256 459
rect 2351 459 2352 463
rect 2356 462 2357 463
rect 2442 463 2448 464
rect 2356 460 2393 462
rect 2356 459 2357 460
rect 2351 458 2357 459
rect 2442 459 2443 463
rect 2447 462 2448 463
rect 2642 463 2648 464
rect 2447 460 2497 462
rect 2447 459 2448 460
rect 2442 458 2448 459
rect 2642 459 2643 463
rect 2647 462 2648 463
rect 2842 463 2848 464
rect 2647 460 2697 462
rect 2647 459 2648 460
rect 2642 458 2648 459
rect 2842 459 2843 463
rect 2847 459 2848 463
rect 3030 463 3036 464
rect 3030 462 3031 463
rect 2965 460 3031 462
rect 2842 458 2848 459
rect 3030 459 3031 460
rect 3035 459 3036 463
rect 3030 458 3036 459
rect 3090 463 3096 464
rect 3090 459 3091 463
rect 3095 459 3096 463
rect 3090 458 3096 459
rect 3226 463 3232 464
rect 3226 459 3227 463
rect 3231 459 3232 463
rect 3226 458 3232 459
rect 3326 463 3332 464
rect 3326 459 3327 463
rect 3331 459 3332 463
rect 3326 458 3332 459
rect 759 454 765 455
rect 1870 455 1876 456
rect 1870 451 1871 455
rect 1875 451 1876 455
rect 3590 455 3596 456
rect 1870 450 1876 451
rect 2182 452 2188 453
rect 2182 448 2183 452
rect 2187 448 2188 452
rect 2182 447 2188 448
rect 2278 452 2284 453
rect 2278 448 2279 452
rect 2283 448 2284 452
rect 2278 447 2284 448
rect 2374 452 2380 453
rect 2374 448 2375 452
rect 2379 448 2380 452
rect 2374 447 2380 448
rect 2478 452 2484 453
rect 2478 448 2479 452
rect 2483 448 2484 452
rect 2478 447 2484 448
rect 2574 452 2580 453
rect 2574 448 2575 452
rect 2579 448 2580 452
rect 2574 447 2580 448
rect 2678 452 2684 453
rect 2678 448 2679 452
rect 2683 448 2684 452
rect 2678 447 2684 448
rect 2782 452 2788 453
rect 2782 448 2783 452
rect 2787 448 2788 452
rect 2782 447 2788 448
rect 2902 452 2908 453
rect 2902 448 2903 452
rect 2907 448 2908 452
rect 2902 447 2908 448
rect 3030 452 3036 453
rect 3030 448 3031 452
rect 3035 448 3036 452
rect 3030 447 3036 448
rect 3166 452 3172 453
rect 3166 448 3167 452
rect 3171 448 3172 452
rect 3166 447 3172 448
rect 3310 452 3316 453
rect 3310 448 3311 452
rect 3315 448 3316 452
rect 3310 447 3316 448
rect 3462 452 3468 453
rect 3462 448 3463 452
rect 3467 448 3468 452
rect 3590 451 3591 455
rect 3595 451 3596 455
rect 3590 450 3596 451
rect 3462 447 3468 448
rect 1990 435 1996 436
rect 1990 431 1991 435
rect 1995 434 1996 435
rect 2199 435 2205 436
rect 2199 434 2200 435
rect 1995 432 2200 434
rect 1995 431 1996 432
rect 1990 430 1996 431
rect 2199 431 2200 432
rect 2204 431 2205 435
rect 2199 430 2205 431
rect 2486 435 2492 436
rect 2486 431 2487 435
rect 2491 434 2492 435
rect 2591 435 2597 436
rect 2591 434 2592 435
rect 2491 432 2592 434
rect 2491 431 2492 432
rect 2486 430 2492 431
rect 2591 431 2592 432
rect 2596 431 2597 435
rect 2591 430 2597 431
rect 3479 435 3485 436
rect 3479 431 3480 435
rect 3484 434 3485 435
rect 3487 435 3493 436
rect 3487 434 3488 435
rect 3484 432 3488 434
rect 3484 431 3485 432
rect 3479 430 3485 431
rect 3487 431 3488 432
rect 3492 431 3493 435
rect 3487 430 3493 431
rect 222 424 228 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 222 420 223 424
rect 227 420 228 424
rect 222 419 228 420
rect 334 424 340 425
rect 334 420 335 424
rect 339 420 340 424
rect 334 419 340 420
rect 446 424 452 425
rect 446 420 447 424
rect 451 420 452 424
rect 446 419 452 420
rect 558 424 564 425
rect 558 420 559 424
rect 563 420 564 424
rect 558 419 564 420
rect 662 424 668 425
rect 662 420 663 424
rect 667 420 668 424
rect 662 419 668 420
rect 758 424 764 425
rect 758 420 759 424
rect 763 420 764 424
rect 758 419 764 420
rect 846 424 852 425
rect 846 420 847 424
rect 851 420 852 424
rect 846 419 852 420
rect 934 424 940 425
rect 934 420 935 424
rect 939 420 940 424
rect 934 419 940 420
rect 1022 424 1028 425
rect 1022 420 1023 424
rect 1027 420 1028 424
rect 1022 419 1028 420
rect 1110 424 1116 425
rect 1110 420 1111 424
rect 1115 420 1116 424
rect 1110 419 1116 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1294 424 1300 425
rect 1294 420 1295 424
rect 1299 420 1300 424
rect 1294 419 1300 420
rect 1830 421 1836 422
rect 110 416 116 417
rect 1830 417 1831 421
rect 1835 417 1836 421
rect 1830 416 1836 417
rect 290 415 296 416
rect 290 414 291 415
rect 285 412 291 414
rect 290 411 291 412
rect 295 411 296 415
rect 290 410 296 411
rect 298 415 304 416
rect 298 411 299 415
rect 303 414 304 415
rect 402 415 408 416
rect 303 412 353 414
rect 303 411 304 412
rect 298 410 304 411
rect 402 411 403 415
rect 407 414 408 415
rect 535 415 541 416
rect 407 412 465 414
rect 407 411 408 412
rect 402 410 408 411
rect 535 411 536 415
rect 540 414 541 415
rect 647 415 653 416
rect 540 412 577 414
rect 540 411 541 412
rect 535 410 541 411
rect 647 411 648 415
rect 652 414 653 415
rect 730 415 736 416
rect 652 412 681 414
rect 652 411 653 412
rect 647 410 653 411
rect 730 411 731 415
rect 735 414 736 415
rect 914 415 920 416
rect 735 412 777 414
rect 735 411 736 412
rect 730 410 736 411
rect 854 411 860 412
rect 854 407 855 411
rect 859 410 860 411
rect 864 410 866 413
rect 914 411 915 415
rect 919 414 920 415
rect 1002 415 1008 416
rect 919 412 953 414
rect 919 411 920 412
rect 914 410 920 411
rect 1002 411 1003 415
rect 1007 414 1008 415
rect 1090 415 1096 416
rect 1007 412 1041 414
rect 1007 411 1008 412
rect 1002 410 1008 411
rect 1090 411 1091 415
rect 1095 414 1096 415
rect 1266 415 1272 416
rect 1266 414 1267 415
rect 1095 412 1129 414
rect 1261 412 1267 414
rect 1095 411 1096 412
rect 1090 410 1096 411
rect 1266 411 1267 412
rect 1271 411 1272 415
rect 1266 410 1272 411
rect 859 408 866 410
rect 859 407 860 408
rect 854 406 860 407
rect 1170 407 1176 408
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 1170 403 1171 407
rect 1175 406 1176 407
rect 1312 406 1314 413
rect 1175 404 1314 406
rect 1830 404 1836 405
rect 1175 403 1176 404
rect 1170 402 1176 403
rect 110 399 116 400
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1974 404 1980 405
rect 1830 399 1836 400
rect 1870 401 1876 402
rect 1870 397 1871 401
rect 1875 397 1876 401
rect 1974 400 1975 404
rect 1979 400 1980 404
rect 1974 399 1980 400
rect 2062 404 2068 405
rect 2062 400 2063 404
rect 2067 400 2068 404
rect 2062 399 2068 400
rect 2158 404 2164 405
rect 2158 400 2159 404
rect 2163 400 2164 404
rect 2158 399 2164 400
rect 2254 404 2260 405
rect 2254 400 2255 404
rect 2259 400 2260 404
rect 2254 399 2260 400
rect 2358 404 2364 405
rect 2358 400 2359 404
rect 2363 400 2364 404
rect 2358 399 2364 400
rect 2470 404 2476 405
rect 2470 400 2471 404
rect 2475 400 2476 404
rect 2470 399 2476 400
rect 2606 404 2612 405
rect 2606 400 2607 404
rect 2611 400 2612 404
rect 2606 399 2612 400
rect 2758 404 2764 405
rect 2758 400 2759 404
rect 2763 400 2764 404
rect 2758 399 2764 400
rect 2926 404 2932 405
rect 2926 400 2927 404
rect 2931 400 2932 404
rect 2926 399 2932 400
rect 3110 404 3116 405
rect 3110 400 3111 404
rect 3115 400 3116 404
rect 3110 399 3116 400
rect 3302 404 3308 405
rect 3302 400 3303 404
rect 3307 400 3308 404
rect 3302 399 3308 400
rect 3494 404 3500 405
rect 3494 400 3495 404
rect 3499 400 3500 404
rect 3494 399 3500 400
rect 3590 401 3596 402
rect 1870 396 1876 397
rect 3590 397 3591 401
rect 3595 397 3596 401
rect 3590 396 3596 397
rect 2042 395 2048 396
rect 2042 394 2043 395
rect 2037 392 2043 394
rect 2042 391 2043 392
rect 2047 391 2048 395
rect 2130 395 2136 396
rect 2130 394 2131 395
rect 2125 392 2131 394
rect 2042 390 2048 391
rect 2130 391 2131 392
rect 2135 391 2136 395
rect 2226 395 2232 396
rect 2226 394 2227 395
rect 2221 392 2227 394
rect 2130 390 2136 391
rect 2226 391 2227 392
rect 2231 391 2232 395
rect 2327 395 2333 396
rect 2327 394 2328 395
rect 2317 392 2328 394
rect 2226 390 2232 391
rect 2327 391 2328 392
rect 2332 391 2333 395
rect 2538 395 2544 396
rect 2538 394 2539 395
rect 2327 390 2333 391
rect 2231 387 2237 388
rect 230 386 236 387
rect 230 382 231 386
rect 235 382 236 386
rect 230 381 236 382
rect 342 386 348 387
rect 342 382 343 386
rect 347 382 348 386
rect 342 381 348 382
rect 454 386 460 387
rect 454 382 455 386
rect 459 382 460 386
rect 454 381 460 382
rect 566 386 572 387
rect 566 382 567 386
rect 571 382 572 386
rect 566 381 572 382
rect 670 386 676 387
rect 670 382 671 386
rect 675 382 676 386
rect 670 381 676 382
rect 766 386 772 387
rect 766 382 767 386
rect 771 382 772 386
rect 766 381 772 382
rect 854 386 860 387
rect 854 382 855 386
rect 859 382 860 386
rect 854 381 860 382
rect 942 386 948 387
rect 942 382 943 386
rect 947 382 948 386
rect 942 381 948 382
rect 1030 386 1036 387
rect 1030 382 1031 386
rect 1035 382 1036 386
rect 1030 381 1036 382
rect 1118 386 1124 387
rect 1118 382 1119 386
rect 1123 382 1124 386
rect 1118 381 1124 382
rect 1206 386 1212 387
rect 1206 382 1207 386
rect 1211 382 1212 386
rect 1206 381 1212 382
rect 1302 386 1308 387
rect 1302 382 1303 386
rect 1307 382 1308 386
rect 1302 381 1308 382
rect 1870 384 1876 385
rect 1870 380 1871 384
rect 1875 380 1876 384
rect 2231 383 2232 387
rect 2236 386 2237 387
rect 2376 386 2378 393
rect 2533 392 2539 394
rect 2538 391 2539 392
rect 2543 391 2544 395
rect 2682 395 2688 396
rect 2682 394 2683 395
rect 2669 392 2683 394
rect 2538 390 2544 391
rect 2682 391 2683 392
rect 2687 391 2688 395
rect 2850 395 2856 396
rect 2850 394 2851 395
rect 2821 392 2851 394
rect 2682 390 2688 391
rect 2850 391 2851 392
rect 2855 391 2856 395
rect 3026 395 3032 396
rect 3026 394 3027 395
rect 2989 392 3027 394
rect 2850 390 2856 391
rect 3026 391 3027 392
rect 3031 391 3032 395
rect 3026 390 3032 391
rect 3034 395 3040 396
rect 3034 391 3035 395
rect 3039 394 3040 395
rect 3390 395 3396 396
rect 3390 394 3391 395
rect 3039 392 3129 394
rect 3365 392 3391 394
rect 3039 391 3040 392
rect 3034 390 3040 391
rect 3390 391 3391 392
rect 3395 391 3396 395
rect 3496 392 3513 394
rect 3390 390 3396 391
rect 3494 391 3500 392
rect 3494 387 3495 391
rect 3499 387 3500 391
rect 3494 386 3500 387
rect 2236 384 2378 386
rect 3590 384 3596 385
rect 2236 383 2237 384
rect 2231 382 2237 383
rect 1870 379 1876 380
rect 3590 380 3591 384
rect 3595 380 3596 384
rect 3590 379 3596 380
rect 223 375 229 376
rect 223 371 224 375
rect 228 374 229 375
rect 298 375 304 376
rect 298 374 299 375
rect 228 372 299 374
rect 228 371 229 372
rect 223 370 229 371
rect 298 371 299 372
rect 303 371 304 375
rect 298 370 304 371
rect 335 375 341 376
rect 335 371 336 375
rect 340 374 341 375
rect 402 375 408 376
rect 402 374 403 375
rect 340 372 403 374
rect 340 371 341 372
rect 335 370 341 371
rect 402 371 403 372
rect 407 371 408 375
rect 402 370 408 371
rect 446 375 453 376
rect 446 371 447 375
rect 452 371 453 375
rect 446 370 453 371
rect 559 375 565 376
rect 559 371 560 375
rect 564 374 565 375
rect 647 375 653 376
rect 647 374 648 375
rect 564 372 648 374
rect 564 371 565 372
rect 559 370 565 371
rect 647 371 648 372
rect 652 371 653 375
rect 647 370 653 371
rect 663 375 669 376
rect 663 371 664 375
rect 668 374 669 375
rect 730 375 736 376
rect 730 374 731 375
rect 668 372 731 374
rect 668 371 669 372
rect 663 370 669 371
rect 730 371 731 372
rect 735 371 736 375
rect 730 370 736 371
rect 751 375 757 376
rect 751 371 752 375
rect 756 374 757 375
rect 759 375 765 376
rect 759 374 760 375
rect 756 372 760 374
rect 756 371 757 372
rect 751 370 757 371
rect 759 371 760 372
rect 764 371 765 375
rect 759 370 765 371
rect 847 375 853 376
rect 847 371 848 375
rect 852 374 853 375
rect 914 375 920 376
rect 914 374 915 375
rect 852 372 915 374
rect 852 371 853 372
rect 847 370 853 371
rect 914 371 915 372
rect 919 371 920 375
rect 914 370 920 371
rect 935 375 941 376
rect 935 371 936 375
rect 940 374 941 375
rect 1002 375 1008 376
rect 1002 374 1003 375
rect 940 372 1003 374
rect 940 371 941 372
rect 935 370 941 371
rect 1002 371 1003 372
rect 1007 371 1008 375
rect 1002 370 1008 371
rect 1023 375 1029 376
rect 1023 371 1024 375
rect 1028 374 1029 375
rect 1090 375 1096 376
rect 1090 374 1091 375
rect 1028 372 1091 374
rect 1028 371 1029 372
rect 1023 370 1029 371
rect 1090 371 1091 372
rect 1095 371 1096 375
rect 1090 370 1096 371
rect 1111 375 1117 376
rect 1111 371 1112 375
rect 1116 374 1117 375
rect 1170 375 1176 376
rect 1170 374 1171 375
rect 1116 372 1171 374
rect 1116 371 1117 372
rect 1111 370 1117 371
rect 1170 371 1171 372
rect 1175 371 1176 375
rect 1170 370 1176 371
rect 1178 375 1184 376
rect 1178 371 1179 375
rect 1183 374 1184 375
rect 1199 375 1205 376
rect 1199 374 1200 375
rect 1183 372 1200 374
rect 1183 371 1184 372
rect 1178 370 1184 371
rect 1199 371 1200 372
rect 1204 371 1205 375
rect 1199 370 1205 371
rect 1266 375 1272 376
rect 1266 371 1267 375
rect 1271 374 1272 375
rect 1295 375 1301 376
rect 1295 374 1296 375
rect 1271 372 1296 374
rect 1271 371 1272 372
rect 1266 370 1272 371
rect 1295 371 1296 372
rect 1300 371 1301 375
rect 1295 370 1301 371
rect 1982 366 1988 367
rect 1982 362 1983 366
rect 1987 362 1988 366
rect 1982 361 1988 362
rect 2070 366 2076 367
rect 2070 362 2071 366
rect 2075 362 2076 366
rect 2070 361 2076 362
rect 2166 366 2172 367
rect 2166 362 2167 366
rect 2171 362 2172 366
rect 2166 361 2172 362
rect 2262 366 2268 367
rect 2262 362 2263 366
rect 2267 362 2268 366
rect 2262 361 2268 362
rect 2366 366 2372 367
rect 2366 362 2367 366
rect 2371 362 2372 366
rect 2366 361 2372 362
rect 2478 366 2484 367
rect 2478 362 2479 366
rect 2483 362 2484 366
rect 2478 361 2484 362
rect 2614 366 2620 367
rect 2614 362 2615 366
rect 2619 362 2620 366
rect 2614 361 2620 362
rect 2766 366 2772 367
rect 2766 362 2767 366
rect 2771 362 2772 366
rect 2766 361 2772 362
rect 2934 366 2940 367
rect 2934 362 2935 366
rect 2939 362 2940 366
rect 2934 361 2940 362
rect 3118 366 3124 367
rect 3118 362 3119 366
rect 3123 362 3124 366
rect 3118 361 3124 362
rect 3310 366 3316 367
rect 3310 362 3311 366
rect 3315 362 3316 366
rect 3310 361 3316 362
rect 3502 366 3508 367
rect 3502 362 3503 366
rect 3507 362 3508 366
rect 3502 361 3508 362
rect 1238 359 1244 360
rect 1238 358 1239 359
rect 956 356 1239 358
rect 127 351 133 352
rect 127 347 128 351
rect 132 350 133 351
rect 135 351 141 352
rect 135 350 136 351
rect 132 348 136 350
rect 132 347 133 348
rect 127 346 133 347
rect 135 347 136 348
rect 140 347 141 351
rect 135 346 141 347
rect 194 351 200 352
rect 194 347 195 351
rect 199 350 200 351
rect 255 351 261 352
rect 255 350 256 351
rect 199 348 256 350
rect 199 347 200 348
rect 194 346 200 347
rect 255 347 256 348
rect 260 347 261 351
rect 255 346 261 347
rect 314 351 320 352
rect 314 347 315 351
rect 319 350 320 351
rect 391 351 397 352
rect 391 350 392 351
rect 319 348 392 350
rect 319 347 320 348
rect 314 346 320 347
rect 391 347 392 348
rect 396 347 397 351
rect 391 346 397 347
rect 527 351 533 352
rect 527 347 528 351
rect 532 350 533 351
rect 535 351 541 352
rect 535 350 536 351
rect 532 348 536 350
rect 532 347 533 348
rect 527 346 533 347
rect 535 347 536 348
rect 540 347 541 351
rect 535 346 541 347
rect 586 351 592 352
rect 586 347 587 351
rect 591 350 592 351
rect 663 351 669 352
rect 663 350 664 351
rect 591 348 664 350
rect 591 347 592 348
rect 586 346 592 347
rect 663 347 664 348
rect 668 347 669 351
rect 663 346 669 347
rect 722 351 728 352
rect 722 347 723 351
rect 727 350 728 351
rect 783 351 789 352
rect 783 350 784 351
rect 727 348 784 350
rect 727 347 728 348
rect 722 346 728 347
rect 783 347 784 348
rect 788 347 789 351
rect 783 346 789 347
rect 903 351 909 352
rect 903 347 904 351
rect 908 350 909 351
rect 956 350 958 356
rect 1238 355 1239 356
rect 1243 355 1244 359
rect 1446 359 1452 360
rect 1446 358 1447 359
rect 1238 354 1244 355
rect 1304 356 1447 358
rect 908 348 958 350
rect 962 351 968 352
rect 908 347 909 348
rect 903 346 909 347
rect 962 347 963 351
rect 967 350 968 351
rect 1015 351 1021 352
rect 1015 350 1016 351
rect 967 348 1016 350
rect 967 347 968 348
rect 962 346 968 347
rect 1015 347 1016 348
rect 1020 347 1021 351
rect 1015 346 1021 347
rect 1074 351 1080 352
rect 1074 347 1075 351
rect 1079 350 1080 351
rect 1119 351 1125 352
rect 1119 350 1120 351
rect 1079 348 1120 350
rect 1079 347 1080 348
rect 1074 346 1080 347
rect 1119 347 1120 348
rect 1124 347 1125 351
rect 1119 346 1125 347
rect 1223 351 1229 352
rect 1223 347 1224 351
rect 1228 350 1229 351
rect 1304 350 1306 356
rect 1446 355 1447 356
rect 1451 355 1452 359
rect 1446 354 1452 355
rect 1975 355 1981 356
rect 1228 348 1306 350
rect 1310 351 1316 352
rect 1228 347 1229 348
rect 1223 346 1229 347
rect 1310 347 1311 351
rect 1315 350 1316 351
rect 1327 351 1333 352
rect 1327 350 1328 351
rect 1315 348 1328 350
rect 1315 347 1316 348
rect 1310 346 1316 347
rect 1327 347 1328 348
rect 1332 347 1333 351
rect 1327 346 1333 347
rect 1386 351 1392 352
rect 1386 347 1387 351
rect 1391 350 1392 351
rect 1431 351 1437 352
rect 1431 350 1432 351
rect 1391 348 1432 350
rect 1391 347 1392 348
rect 1386 346 1392 347
rect 1431 347 1432 348
rect 1436 347 1437 351
rect 1975 351 1976 355
rect 1980 354 1981 355
rect 1990 355 1996 356
rect 1990 354 1991 355
rect 1980 352 1991 354
rect 1980 351 1981 352
rect 1975 350 1981 351
rect 1990 351 1991 352
rect 1995 351 1996 355
rect 1990 350 1996 351
rect 2042 355 2048 356
rect 2042 351 2043 355
rect 2047 354 2048 355
rect 2063 355 2069 356
rect 2063 354 2064 355
rect 2047 352 2064 354
rect 2047 351 2048 352
rect 2042 350 2048 351
rect 2063 351 2064 352
rect 2068 351 2069 355
rect 2063 350 2069 351
rect 2130 355 2136 356
rect 2130 351 2131 355
rect 2135 354 2136 355
rect 2159 355 2165 356
rect 2159 354 2160 355
rect 2135 352 2160 354
rect 2135 351 2136 352
rect 2130 350 2136 351
rect 2159 351 2160 352
rect 2164 351 2165 355
rect 2159 350 2165 351
rect 2226 355 2232 356
rect 2226 351 2227 355
rect 2231 354 2232 355
rect 2255 355 2261 356
rect 2255 354 2256 355
rect 2231 352 2256 354
rect 2231 351 2232 352
rect 2226 350 2232 351
rect 2255 351 2256 352
rect 2260 351 2261 355
rect 2255 350 2261 351
rect 2327 355 2333 356
rect 2327 351 2328 355
rect 2332 354 2333 355
rect 2359 355 2365 356
rect 2359 354 2360 355
rect 2332 352 2360 354
rect 2332 351 2333 352
rect 2327 350 2333 351
rect 2359 351 2360 352
rect 2364 351 2365 355
rect 2359 350 2365 351
rect 2471 355 2477 356
rect 2471 351 2472 355
rect 2476 354 2477 355
rect 2486 355 2492 356
rect 2486 354 2487 355
rect 2476 352 2487 354
rect 2476 351 2477 352
rect 2471 350 2477 351
rect 2486 351 2487 352
rect 2491 351 2492 355
rect 2486 350 2492 351
rect 2538 355 2544 356
rect 2538 351 2539 355
rect 2543 354 2544 355
rect 2607 355 2613 356
rect 2607 354 2608 355
rect 2543 352 2608 354
rect 2543 351 2544 352
rect 2538 350 2544 351
rect 2607 351 2608 352
rect 2612 351 2613 355
rect 2607 350 2613 351
rect 2682 355 2688 356
rect 2682 351 2683 355
rect 2687 354 2688 355
rect 2759 355 2765 356
rect 2759 354 2760 355
rect 2687 352 2760 354
rect 2687 351 2688 352
rect 2682 350 2688 351
rect 2759 351 2760 352
rect 2764 351 2765 355
rect 2759 350 2765 351
rect 2850 355 2856 356
rect 2850 351 2851 355
rect 2855 354 2856 355
rect 2927 355 2933 356
rect 2927 354 2928 355
rect 2855 352 2928 354
rect 2855 351 2856 352
rect 2850 350 2856 351
rect 2927 351 2928 352
rect 2932 351 2933 355
rect 2927 350 2933 351
rect 3026 355 3032 356
rect 3026 351 3027 355
rect 3031 354 3032 355
rect 3111 355 3117 356
rect 3111 354 3112 355
rect 3031 352 3112 354
rect 3031 351 3032 352
rect 3026 350 3032 351
rect 3111 351 3112 352
rect 3116 351 3117 355
rect 3111 350 3117 351
rect 3303 355 3309 356
rect 3303 351 3304 355
rect 3308 354 3309 355
rect 3398 355 3404 356
rect 3398 354 3399 355
rect 3308 352 3399 354
rect 3308 351 3309 352
rect 3303 350 3309 351
rect 3398 351 3399 352
rect 3403 351 3404 355
rect 3398 350 3404 351
rect 3487 355 3493 356
rect 3487 351 3488 355
rect 3492 354 3493 355
rect 3495 355 3501 356
rect 3495 354 3496 355
rect 3492 352 3496 354
rect 3492 351 3493 352
rect 3487 350 3493 351
rect 3495 351 3496 352
rect 3500 351 3501 355
rect 3495 350 3501 351
rect 1431 346 1437 347
rect 142 342 148 343
rect 142 338 143 342
rect 147 338 148 342
rect 142 337 148 338
rect 262 342 268 343
rect 262 338 263 342
rect 267 338 268 342
rect 262 337 268 338
rect 398 342 404 343
rect 398 338 399 342
rect 403 338 404 342
rect 398 337 404 338
rect 534 342 540 343
rect 534 338 535 342
rect 539 338 540 342
rect 534 337 540 338
rect 670 342 676 343
rect 670 338 671 342
rect 675 338 676 342
rect 670 337 676 338
rect 790 342 796 343
rect 790 338 791 342
rect 795 338 796 342
rect 790 337 796 338
rect 910 342 916 343
rect 910 338 911 342
rect 915 338 916 342
rect 910 337 916 338
rect 1022 342 1028 343
rect 1022 338 1023 342
rect 1027 338 1028 342
rect 1022 337 1028 338
rect 1126 342 1132 343
rect 1126 338 1127 342
rect 1131 338 1132 342
rect 1126 337 1132 338
rect 1230 342 1236 343
rect 1230 338 1231 342
rect 1235 338 1236 342
rect 1230 337 1236 338
rect 1334 342 1340 343
rect 1334 338 1335 342
rect 1339 338 1340 342
rect 1334 337 1340 338
rect 1438 342 1444 343
rect 1438 338 1439 342
rect 1443 338 1444 342
rect 1438 337 1444 338
rect 2207 339 2213 340
rect 2207 335 2208 339
rect 2212 338 2213 339
rect 2231 339 2237 340
rect 2231 338 2232 339
rect 2212 336 2232 338
rect 2212 335 2213 336
rect 2207 334 2213 335
rect 2231 335 2232 336
rect 2236 335 2237 339
rect 2231 334 2237 335
rect 2274 339 2280 340
rect 2274 335 2275 339
rect 2279 338 2280 339
rect 2287 339 2293 340
rect 2287 338 2288 339
rect 2279 336 2288 338
rect 2279 335 2280 336
rect 2274 334 2280 335
rect 2287 335 2288 336
rect 2292 335 2293 339
rect 2287 334 2293 335
rect 2346 339 2352 340
rect 2346 335 2347 339
rect 2351 338 2352 339
rect 2375 339 2381 340
rect 2375 338 2376 339
rect 2351 336 2376 338
rect 2351 335 2352 336
rect 2346 334 2352 335
rect 2375 335 2376 336
rect 2380 335 2381 339
rect 2375 334 2381 335
rect 2434 339 2440 340
rect 2434 335 2435 339
rect 2439 338 2440 339
rect 2471 339 2477 340
rect 2471 338 2472 339
rect 2439 336 2472 338
rect 2439 335 2440 336
rect 2434 334 2440 335
rect 2471 335 2472 336
rect 2476 335 2477 339
rect 2471 334 2477 335
rect 2530 339 2536 340
rect 2530 335 2531 339
rect 2535 338 2536 339
rect 2583 339 2589 340
rect 2583 338 2584 339
rect 2535 336 2584 338
rect 2535 335 2536 336
rect 2530 334 2536 335
rect 2583 335 2584 336
rect 2588 335 2589 339
rect 2583 334 2589 335
rect 2642 339 2648 340
rect 2642 335 2643 339
rect 2647 338 2648 339
rect 2711 339 2717 340
rect 2711 338 2712 339
rect 2647 336 2712 338
rect 2647 335 2648 336
rect 2642 334 2648 335
rect 2711 335 2712 336
rect 2716 335 2717 339
rect 2711 334 2717 335
rect 2839 339 2845 340
rect 2839 335 2840 339
rect 2844 338 2845 339
rect 2906 339 2912 340
rect 2906 338 2907 339
rect 2844 336 2907 338
rect 2844 335 2845 336
rect 2839 334 2845 335
rect 2906 335 2907 336
rect 2911 335 2912 339
rect 2906 334 2912 335
rect 2975 339 2981 340
rect 2975 335 2976 339
rect 2980 338 2981 339
rect 3034 339 3040 340
rect 3034 338 3035 339
rect 2980 336 3035 338
rect 2980 335 2981 336
rect 2975 334 2981 335
rect 3034 335 3035 336
rect 3039 335 3040 339
rect 3034 334 3040 335
rect 3102 339 3108 340
rect 3102 335 3103 339
rect 3107 338 3108 339
rect 3111 339 3117 340
rect 3111 338 3112 339
rect 3107 336 3112 338
rect 3107 335 3108 336
rect 3102 334 3108 335
rect 3111 335 3112 336
rect 3116 335 3117 339
rect 3111 334 3117 335
rect 3170 339 3176 340
rect 3170 335 3171 339
rect 3175 338 3176 339
rect 3247 339 3253 340
rect 3247 338 3248 339
rect 3175 336 3248 338
rect 3175 335 3176 336
rect 3170 334 3176 335
rect 3247 335 3248 336
rect 3252 335 3253 339
rect 3247 334 3253 335
rect 3370 339 3376 340
rect 3370 335 3371 339
rect 3375 338 3376 339
rect 3383 339 3389 340
rect 3383 338 3384 339
rect 3375 336 3384 338
rect 3375 335 3376 336
rect 3370 334 3376 335
rect 3383 335 3384 336
rect 3388 335 3389 339
rect 3383 334 3389 335
rect 3494 339 3500 340
rect 3494 335 3495 339
rect 3499 338 3500 339
rect 3503 339 3509 340
rect 3503 338 3504 339
rect 3499 336 3504 338
rect 3499 335 3500 336
rect 3494 334 3500 335
rect 3503 335 3504 336
rect 3508 335 3509 339
rect 3503 334 3509 335
rect 2214 330 2220 331
rect 2214 326 2215 330
rect 2219 326 2220 330
rect 2214 325 2220 326
rect 2294 330 2300 331
rect 2294 326 2295 330
rect 2299 326 2300 330
rect 2294 325 2300 326
rect 2382 330 2388 331
rect 2382 326 2383 330
rect 2387 326 2388 330
rect 2382 325 2388 326
rect 2478 330 2484 331
rect 2478 326 2479 330
rect 2483 326 2484 330
rect 2478 325 2484 326
rect 2590 330 2596 331
rect 2590 326 2591 330
rect 2595 326 2596 330
rect 2590 325 2596 326
rect 2718 330 2724 331
rect 2718 326 2719 330
rect 2723 326 2724 330
rect 2718 325 2724 326
rect 2846 330 2852 331
rect 2846 326 2847 330
rect 2851 326 2852 330
rect 2846 325 2852 326
rect 2982 330 2988 331
rect 2982 326 2983 330
rect 2987 326 2988 330
rect 2982 325 2988 326
rect 3118 330 3124 331
rect 3118 326 3119 330
rect 3123 326 3124 330
rect 3118 325 3124 326
rect 3254 330 3260 331
rect 3254 326 3255 330
rect 3259 326 3260 330
rect 3254 325 3260 326
rect 3390 330 3396 331
rect 3390 326 3391 330
rect 3395 326 3396 330
rect 3390 325 3396 326
rect 3510 330 3516 331
rect 3510 326 3511 330
rect 3515 326 3516 330
rect 3510 325 3516 326
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 110 319 116 320
rect 1830 324 1836 325
rect 1830 320 1831 324
rect 1835 320 1836 324
rect 1830 319 1836 320
rect 194 315 200 316
rect 194 311 195 315
rect 199 311 200 315
rect 194 310 200 311
rect 314 315 320 316
rect 314 311 315 315
rect 319 311 320 315
rect 314 310 320 311
rect 446 315 452 316
rect 446 311 447 315
rect 451 311 452 315
rect 446 310 452 311
rect 586 315 592 316
rect 586 311 587 315
rect 591 311 592 315
rect 586 310 592 311
rect 722 315 728 316
rect 722 311 723 315
rect 727 311 728 315
rect 722 310 728 311
rect 838 315 844 316
rect 838 311 839 315
rect 843 311 844 315
rect 838 310 844 311
rect 962 315 968 316
rect 962 311 963 315
rect 967 311 968 315
rect 962 310 968 311
rect 1074 315 1080 316
rect 1074 311 1075 315
rect 1079 311 1080 315
rect 1074 310 1080 311
rect 1178 315 1184 316
rect 1178 311 1179 315
rect 1183 311 1184 315
rect 1178 310 1184 311
rect 1238 315 1244 316
rect 1238 311 1239 315
rect 1243 311 1244 315
rect 1238 310 1244 311
rect 1386 315 1392 316
rect 1386 311 1387 315
rect 1391 311 1392 315
rect 1386 310 1392 311
rect 1446 315 1452 316
rect 1446 311 1447 315
rect 1451 311 1452 315
rect 1446 310 1452 311
rect 1870 312 1876 313
rect 1870 308 1871 312
rect 1875 308 1876 312
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 1830 307 1836 308
rect 1870 307 1876 308
rect 3590 312 3596 313
rect 3590 308 3591 312
rect 3595 308 3596 312
rect 3590 307 3596 308
rect 110 302 116 303
rect 134 304 140 305
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 254 304 260 305
rect 254 300 255 304
rect 259 300 260 304
rect 254 299 260 300
rect 390 304 396 305
rect 390 300 391 304
rect 395 300 396 304
rect 390 299 396 300
rect 526 304 532 305
rect 526 300 527 304
rect 531 300 532 304
rect 526 299 532 300
rect 662 304 668 305
rect 662 300 663 304
rect 667 300 668 304
rect 662 299 668 300
rect 782 304 788 305
rect 782 300 783 304
rect 787 300 788 304
rect 782 299 788 300
rect 902 304 908 305
rect 902 300 903 304
rect 907 300 908 304
rect 902 299 908 300
rect 1014 304 1020 305
rect 1014 300 1015 304
rect 1019 300 1020 304
rect 1014 299 1020 300
rect 1118 304 1124 305
rect 1118 300 1119 304
rect 1123 300 1124 304
rect 1118 299 1124 300
rect 1222 304 1228 305
rect 1222 300 1223 304
rect 1227 300 1228 304
rect 1222 299 1228 300
rect 1326 304 1332 305
rect 1326 300 1327 304
rect 1331 300 1332 304
rect 1326 299 1332 300
rect 1430 304 1436 305
rect 1430 300 1431 304
rect 1435 300 1436 304
rect 1830 303 1831 307
rect 1835 303 1836 307
rect 1830 302 1836 303
rect 2274 303 2280 304
rect 2274 302 2275 303
rect 2269 300 2275 302
rect 1430 299 1436 300
rect 2274 299 2275 300
rect 2279 299 2280 303
rect 2274 298 2280 299
rect 2346 303 2352 304
rect 2346 299 2347 303
rect 2351 299 2352 303
rect 2346 298 2352 299
rect 2434 303 2440 304
rect 2434 299 2435 303
rect 2439 299 2440 303
rect 2434 298 2440 299
rect 2530 303 2536 304
rect 2530 299 2531 303
rect 2535 299 2536 303
rect 2530 298 2536 299
rect 2642 303 2648 304
rect 2642 299 2643 303
rect 2647 299 2648 303
rect 2642 298 2648 299
rect 2898 303 2904 304
rect 2898 299 2899 303
rect 2903 299 2904 303
rect 2898 298 2904 299
rect 2906 303 2912 304
rect 2906 299 2907 303
rect 2911 302 2912 303
rect 3170 303 3176 304
rect 2911 300 2993 302
rect 2911 299 2912 300
rect 2906 298 2912 299
rect 3170 299 3171 303
rect 3175 299 3176 303
rect 3370 303 3376 304
rect 3370 302 3371 303
rect 3309 300 3371 302
rect 3170 298 3176 299
rect 3370 299 3371 300
rect 3375 299 3376 303
rect 3370 298 3376 299
rect 3398 303 3404 304
rect 3398 299 3399 303
rect 3403 299 3404 303
rect 3398 298 3404 299
rect 1870 295 1876 296
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 3590 295 3596 296
rect 1870 290 1876 291
rect 2206 292 2212 293
rect 2206 288 2207 292
rect 2211 288 2212 292
rect 2206 287 2212 288
rect 2286 292 2292 293
rect 2286 288 2287 292
rect 2291 288 2292 292
rect 2286 287 2292 288
rect 2374 292 2380 293
rect 2374 288 2375 292
rect 2379 288 2380 292
rect 2374 287 2380 288
rect 2470 292 2476 293
rect 2470 288 2471 292
rect 2475 288 2476 292
rect 2470 287 2476 288
rect 2582 292 2588 293
rect 2582 288 2583 292
rect 2587 288 2588 292
rect 2582 287 2588 288
rect 2710 292 2716 293
rect 2710 288 2711 292
rect 2715 288 2716 292
rect 2710 287 2716 288
rect 2838 292 2844 293
rect 2838 288 2839 292
rect 2843 288 2844 292
rect 2838 287 2844 288
rect 2974 292 2980 293
rect 2974 288 2975 292
rect 2979 288 2980 292
rect 2974 287 2980 288
rect 3110 292 3116 293
rect 3110 288 3111 292
rect 3115 288 3116 292
rect 3110 287 3116 288
rect 3246 292 3252 293
rect 3246 288 3247 292
rect 3251 288 3252 292
rect 3246 287 3252 288
rect 3382 292 3388 293
rect 3382 288 3383 292
rect 3387 288 3388 292
rect 3382 287 3388 288
rect 3502 292 3508 293
rect 3502 288 3503 292
rect 3507 288 3508 292
rect 3590 291 3591 295
rect 3595 291 3596 295
rect 3590 290 3596 291
rect 3502 287 3508 288
rect 2550 275 2556 276
rect 2550 271 2551 275
rect 2555 274 2556 275
rect 2727 275 2733 276
rect 2727 274 2728 275
rect 2555 272 2728 274
rect 2555 271 2556 272
rect 2550 270 2556 271
rect 2727 271 2728 272
rect 2732 271 2733 275
rect 2727 270 2733 271
rect 3518 275 3525 276
rect 3518 271 3519 275
rect 3524 271 3525 275
rect 3518 270 3525 271
rect 134 252 140 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 246 252 252 253
rect 246 248 247 252
rect 251 248 252 252
rect 246 247 252 248
rect 390 252 396 253
rect 390 248 391 252
rect 395 248 396 252
rect 390 247 396 248
rect 542 252 548 253
rect 542 248 543 252
rect 547 248 548 252
rect 542 247 548 248
rect 694 252 700 253
rect 694 248 695 252
rect 699 248 700 252
rect 694 247 700 248
rect 846 252 852 253
rect 846 248 847 252
rect 851 248 852 252
rect 846 247 852 248
rect 990 252 996 253
rect 990 248 991 252
rect 995 248 996 252
rect 990 247 996 248
rect 1118 252 1124 253
rect 1118 248 1119 252
rect 1123 248 1124 252
rect 1118 247 1124 248
rect 1238 252 1244 253
rect 1238 248 1239 252
rect 1243 248 1244 252
rect 1238 247 1244 248
rect 1358 252 1364 253
rect 1358 248 1359 252
rect 1363 248 1364 252
rect 1358 247 1364 248
rect 1478 252 1484 253
rect 1478 248 1479 252
rect 1483 248 1484 252
rect 1478 247 1484 248
rect 1598 252 1604 253
rect 1598 248 1599 252
rect 1603 248 1604 252
rect 1598 247 1604 248
rect 1830 249 1836 250
rect 110 244 116 245
rect 1830 245 1831 249
rect 1835 245 1836 249
rect 1830 244 1836 245
rect 1990 244 1996 245
rect 127 243 133 244
rect 127 239 128 243
rect 132 242 133 243
rect 202 243 208 244
rect 132 240 153 242
rect 132 239 133 240
rect 127 238 133 239
rect 202 239 203 243
rect 207 242 208 243
rect 314 243 320 244
rect 207 240 265 242
rect 207 239 208 240
rect 202 238 208 239
rect 314 239 315 243
rect 319 242 320 243
rect 610 243 616 244
rect 610 242 611 243
rect 319 240 409 242
rect 605 240 611 242
rect 319 239 320 240
rect 314 238 320 239
rect 610 239 611 240
rect 615 239 616 243
rect 610 238 616 239
rect 647 243 653 244
rect 647 239 648 243
rect 652 242 653 243
rect 762 243 768 244
rect 652 240 713 242
rect 652 239 653 240
rect 647 238 653 239
rect 762 239 763 243
rect 767 242 768 243
rect 1062 243 1068 244
rect 1062 242 1063 243
rect 767 240 865 242
rect 1053 240 1063 242
rect 767 239 768 240
rect 762 238 768 239
rect 1062 239 1063 240
rect 1067 239 1068 243
rect 1186 243 1192 244
rect 1186 242 1187 243
rect 1181 240 1187 242
rect 1062 238 1068 239
rect 1186 239 1187 240
rect 1191 239 1192 243
rect 1310 243 1316 244
rect 1310 242 1311 243
rect 1301 240 1311 242
rect 1186 238 1192 239
rect 1310 239 1311 240
rect 1315 239 1316 243
rect 1426 243 1432 244
rect 1426 242 1427 243
rect 1421 240 1427 242
rect 1310 238 1316 239
rect 1426 239 1427 240
rect 1431 239 1432 243
rect 1546 243 1552 244
rect 1546 242 1547 243
rect 1541 240 1547 242
rect 1426 238 1432 239
rect 1546 239 1547 240
rect 1551 239 1552 243
rect 1870 241 1876 242
rect 1546 238 1552 239
rect 1050 235 1056 236
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 1050 231 1051 235
rect 1055 234 1056 235
rect 1616 234 1618 241
rect 1870 237 1871 241
rect 1875 237 1876 241
rect 1990 240 1991 244
rect 1995 240 1996 244
rect 1990 239 1996 240
rect 2118 244 2124 245
rect 2118 240 2119 244
rect 2123 240 2124 244
rect 2118 239 2124 240
rect 2254 244 2260 245
rect 2254 240 2255 244
rect 2259 240 2260 244
rect 2254 239 2260 240
rect 2390 244 2396 245
rect 2390 240 2391 244
rect 2395 240 2396 244
rect 2390 239 2396 240
rect 2534 244 2540 245
rect 2534 240 2535 244
rect 2539 240 2540 244
rect 2534 239 2540 240
rect 2678 244 2684 245
rect 2678 240 2679 244
rect 2683 240 2684 244
rect 2678 239 2684 240
rect 2814 244 2820 245
rect 2814 240 2815 244
rect 2819 240 2820 244
rect 2814 239 2820 240
rect 2950 244 2956 245
rect 2950 240 2951 244
rect 2955 240 2956 244
rect 2950 239 2956 240
rect 3094 244 3100 245
rect 3094 240 3095 244
rect 3099 240 3100 244
rect 3094 239 3100 240
rect 3238 244 3244 245
rect 3238 240 3239 244
rect 3243 240 3244 244
rect 3238 239 3244 240
rect 3382 244 3388 245
rect 3382 240 3383 244
rect 3387 240 3388 244
rect 3382 239 3388 240
rect 3502 244 3508 245
rect 3502 240 3503 244
rect 3507 240 3508 244
rect 3502 239 3508 240
rect 3590 241 3596 242
rect 1870 236 1876 237
rect 3590 237 3591 241
rect 3595 237 3596 241
rect 3590 236 3596 237
rect 2062 235 2068 236
rect 2062 234 2063 235
rect 1055 232 1618 234
rect 1830 232 1836 233
rect 2053 232 2063 234
rect 1055 231 1056 232
rect 1050 230 1056 231
rect 110 227 116 228
rect 1830 228 1831 232
rect 1835 228 1836 232
rect 2062 231 2063 232
rect 2067 231 2068 235
rect 2186 235 2192 236
rect 2186 234 2187 235
rect 2181 232 2187 234
rect 2062 230 2068 231
rect 2186 231 2187 232
rect 2191 231 2192 235
rect 2334 235 2340 236
rect 2186 230 2192 231
rect 1830 227 1836 228
rect 2050 227 2056 228
rect 1870 224 1876 225
rect 1870 220 1871 224
rect 1875 220 1876 224
rect 2050 223 2051 227
rect 2055 226 2056 227
rect 2272 226 2274 233
rect 2334 231 2335 235
rect 2339 234 2340 235
rect 2458 235 2464 236
rect 2339 232 2409 234
rect 2339 231 2340 232
rect 2334 230 2340 231
rect 2458 231 2459 235
rect 2463 234 2464 235
rect 2623 235 2629 236
rect 2463 232 2553 234
rect 2463 231 2464 232
rect 2458 230 2464 231
rect 2623 231 2624 235
rect 2628 234 2629 235
rect 2746 235 2752 236
rect 2628 232 2697 234
rect 2628 231 2629 232
rect 2623 230 2629 231
rect 2746 231 2747 235
rect 2751 234 2752 235
rect 2882 235 2888 236
rect 2751 232 2833 234
rect 2751 231 2752 232
rect 2746 230 2752 231
rect 2882 231 2883 235
rect 2887 234 2888 235
rect 3194 235 3200 236
rect 2887 232 2969 234
rect 2887 231 2888 232
rect 2882 230 2888 231
rect 3102 231 3108 232
rect 3102 227 3103 231
rect 3107 230 3108 231
rect 3112 230 3114 233
rect 3194 231 3195 235
rect 3199 234 3200 235
rect 3306 235 3312 236
rect 3199 232 3257 234
rect 3199 231 3200 232
rect 3194 230 3200 231
rect 3306 231 3307 235
rect 3311 234 3312 235
rect 3311 232 3401 234
rect 3504 232 3521 234
rect 3311 231 3312 232
rect 3306 230 3312 231
rect 3502 231 3508 232
rect 3107 228 3114 230
rect 3107 227 3108 228
rect 3102 226 3108 227
rect 3502 227 3503 231
rect 3507 227 3508 231
rect 3502 226 3508 227
rect 2055 224 2274 226
rect 3590 224 3596 225
rect 2055 223 2056 224
rect 2050 222 2056 223
rect 1870 219 1876 220
rect 3590 220 3591 224
rect 3595 220 3596 224
rect 3590 219 3596 220
rect 142 214 148 215
rect 142 210 143 214
rect 147 210 148 214
rect 142 209 148 210
rect 254 214 260 215
rect 254 210 255 214
rect 259 210 260 214
rect 254 209 260 210
rect 398 214 404 215
rect 398 210 399 214
rect 403 210 404 214
rect 398 209 404 210
rect 550 214 556 215
rect 550 210 551 214
rect 555 210 556 214
rect 550 209 556 210
rect 702 214 708 215
rect 702 210 703 214
rect 707 210 708 214
rect 702 209 708 210
rect 854 214 860 215
rect 854 210 855 214
rect 859 210 860 214
rect 854 209 860 210
rect 998 214 1004 215
rect 998 210 999 214
rect 1003 210 1004 214
rect 998 209 1004 210
rect 1126 214 1132 215
rect 1126 210 1127 214
rect 1131 210 1132 214
rect 1126 209 1132 210
rect 1246 214 1252 215
rect 1246 210 1247 214
rect 1251 210 1252 214
rect 1246 209 1252 210
rect 1366 214 1372 215
rect 1366 210 1367 214
rect 1371 210 1372 214
rect 1366 209 1372 210
rect 1486 214 1492 215
rect 1486 210 1487 214
rect 1491 210 1492 214
rect 1486 209 1492 210
rect 1606 214 1612 215
rect 1606 210 1607 214
rect 1611 210 1612 214
rect 1606 209 1612 210
rect 1998 206 2004 207
rect 135 203 141 204
rect 135 199 136 203
rect 140 202 141 203
rect 202 203 208 204
rect 202 202 203 203
rect 140 200 203 202
rect 140 199 141 200
rect 135 198 141 199
rect 202 199 203 200
rect 207 199 208 203
rect 202 198 208 199
rect 247 203 253 204
rect 247 199 248 203
rect 252 202 253 203
rect 314 203 320 204
rect 314 202 315 203
rect 252 200 315 202
rect 252 199 253 200
rect 247 198 253 199
rect 314 199 315 200
rect 319 199 320 203
rect 314 198 320 199
rect 354 203 360 204
rect 354 199 355 203
rect 359 202 360 203
rect 391 203 397 204
rect 391 202 392 203
rect 359 200 392 202
rect 359 199 360 200
rect 354 198 360 199
rect 391 199 392 200
rect 396 199 397 203
rect 391 198 397 199
rect 543 203 549 204
rect 543 199 544 203
rect 548 202 549 203
rect 647 203 653 204
rect 647 202 648 203
rect 548 200 648 202
rect 548 199 549 200
rect 543 198 549 199
rect 647 199 648 200
rect 652 199 653 203
rect 647 198 653 199
rect 695 203 701 204
rect 695 199 696 203
rect 700 202 701 203
rect 762 203 768 204
rect 762 202 763 203
rect 700 200 763 202
rect 700 199 701 200
rect 695 198 701 199
rect 762 199 763 200
rect 767 199 768 203
rect 762 198 768 199
rect 838 203 844 204
rect 838 199 839 203
rect 843 202 844 203
rect 847 203 853 204
rect 847 202 848 203
rect 843 200 848 202
rect 843 199 844 200
rect 838 198 844 199
rect 847 199 848 200
rect 852 199 853 203
rect 847 198 853 199
rect 991 203 997 204
rect 991 199 992 203
rect 996 202 997 203
rect 1050 203 1056 204
rect 1050 202 1051 203
rect 996 200 1051 202
rect 996 199 997 200
rect 991 198 997 199
rect 1050 199 1051 200
rect 1055 199 1056 203
rect 1050 198 1056 199
rect 1062 203 1068 204
rect 1062 199 1063 203
rect 1067 202 1068 203
rect 1119 203 1125 204
rect 1119 202 1120 203
rect 1067 200 1120 202
rect 1067 199 1068 200
rect 1062 198 1068 199
rect 1119 199 1120 200
rect 1124 199 1125 203
rect 1119 198 1125 199
rect 1186 203 1192 204
rect 1186 199 1187 203
rect 1191 202 1192 203
rect 1239 203 1245 204
rect 1239 202 1240 203
rect 1191 200 1240 202
rect 1191 199 1192 200
rect 1186 198 1192 199
rect 1239 199 1240 200
rect 1244 199 1245 203
rect 1239 198 1245 199
rect 1358 203 1365 204
rect 1358 199 1359 203
rect 1364 199 1365 203
rect 1358 198 1365 199
rect 1426 203 1432 204
rect 1426 199 1427 203
rect 1431 202 1432 203
rect 1479 203 1485 204
rect 1479 202 1480 203
rect 1431 200 1480 202
rect 1431 199 1432 200
rect 1426 198 1432 199
rect 1479 199 1480 200
rect 1484 199 1485 203
rect 1479 198 1485 199
rect 1546 203 1552 204
rect 1546 199 1547 203
rect 1551 202 1552 203
rect 1599 203 1605 204
rect 1599 202 1600 203
rect 1551 200 1600 202
rect 1551 199 1552 200
rect 1546 198 1552 199
rect 1599 199 1600 200
rect 1604 199 1605 203
rect 1998 202 1999 206
rect 2003 202 2004 206
rect 1998 201 2004 202
rect 2126 206 2132 207
rect 2126 202 2127 206
rect 2131 202 2132 206
rect 2126 201 2132 202
rect 2262 206 2268 207
rect 2262 202 2263 206
rect 2267 202 2268 206
rect 2262 201 2268 202
rect 2398 206 2404 207
rect 2398 202 2399 206
rect 2403 202 2404 206
rect 2398 201 2404 202
rect 2542 206 2548 207
rect 2542 202 2543 206
rect 2547 202 2548 206
rect 2542 201 2548 202
rect 2686 206 2692 207
rect 2686 202 2687 206
rect 2691 202 2692 206
rect 2686 201 2692 202
rect 2822 206 2828 207
rect 2822 202 2823 206
rect 2827 202 2828 206
rect 2822 201 2828 202
rect 2958 206 2964 207
rect 2958 202 2959 206
rect 2963 202 2964 206
rect 2958 201 2964 202
rect 3102 206 3108 207
rect 3102 202 3103 206
rect 3107 202 3108 206
rect 3102 201 3108 202
rect 3246 206 3252 207
rect 3246 202 3247 206
rect 3251 202 3252 206
rect 3246 201 3252 202
rect 3390 206 3396 207
rect 3390 202 3391 206
rect 3395 202 3396 206
rect 3390 201 3396 202
rect 3510 206 3516 207
rect 3510 202 3511 206
rect 3515 202 3516 206
rect 3510 201 3516 202
rect 1599 198 1605 199
rect 1991 195 1997 196
rect 1991 191 1992 195
rect 1996 194 1997 195
rect 2050 195 2056 196
rect 2050 194 2051 195
rect 1996 192 2051 194
rect 1996 191 1997 192
rect 1991 190 1997 191
rect 2050 191 2051 192
rect 2055 191 2056 195
rect 2050 190 2056 191
rect 2062 195 2068 196
rect 2062 191 2063 195
rect 2067 194 2068 195
rect 2119 195 2125 196
rect 2119 194 2120 195
rect 2067 192 2120 194
rect 2067 191 2068 192
rect 2062 190 2068 191
rect 2119 191 2120 192
rect 2124 191 2125 195
rect 2119 190 2125 191
rect 2255 195 2261 196
rect 2255 191 2256 195
rect 2260 194 2261 195
rect 2334 195 2340 196
rect 2334 194 2335 195
rect 2260 192 2335 194
rect 2260 191 2261 192
rect 2255 190 2261 191
rect 2334 191 2335 192
rect 2339 191 2340 195
rect 2334 190 2340 191
rect 2391 195 2397 196
rect 2391 191 2392 195
rect 2396 194 2397 195
rect 2458 195 2464 196
rect 2458 194 2459 195
rect 2396 192 2459 194
rect 2396 191 2397 192
rect 2391 190 2397 191
rect 2458 191 2459 192
rect 2463 191 2464 195
rect 2458 190 2464 191
rect 2535 195 2541 196
rect 2535 191 2536 195
rect 2540 194 2541 195
rect 2550 195 2556 196
rect 2550 194 2551 195
rect 2540 192 2551 194
rect 2540 191 2541 192
rect 2535 190 2541 191
rect 2550 191 2551 192
rect 2555 191 2556 195
rect 2550 190 2556 191
rect 2679 195 2685 196
rect 2679 191 2680 195
rect 2684 194 2685 195
rect 2746 195 2752 196
rect 2746 194 2747 195
rect 2684 192 2747 194
rect 2684 191 2685 192
rect 2679 190 2685 191
rect 2746 191 2747 192
rect 2751 191 2752 195
rect 2746 190 2752 191
rect 2815 195 2821 196
rect 2815 191 2816 195
rect 2820 194 2821 195
rect 2882 195 2888 196
rect 2882 194 2883 195
rect 2820 192 2883 194
rect 2820 191 2821 192
rect 2815 190 2821 191
rect 2882 191 2883 192
rect 2887 191 2888 195
rect 2882 190 2888 191
rect 2898 195 2904 196
rect 2898 191 2899 195
rect 2903 194 2904 195
rect 2951 195 2957 196
rect 2951 194 2952 195
rect 2903 192 2952 194
rect 2903 191 2904 192
rect 2898 190 2904 191
rect 2951 191 2952 192
rect 2956 191 2957 195
rect 2951 190 2957 191
rect 3095 195 3101 196
rect 3095 191 3096 195
rect 3100 194 3101 195
rect 3194 195 3200 196
rect 3194 194 3195 195
rect 3100 192 3195 194
rect 3100 191 3101 192
rect 3095 190 3101 191
rect 3194 191 3195 192
rect 3199 191 3200 195
rect 3194 190 3200 191
rect 3239 195 3245 196
rect 3239 191 3240 195
rect 3244 194 3245 195
rect 3306 195 3312 196
rect 3306 194 3307 195
rect 3244 192 3307 194
rect 3244 191 3245 192
rect 3239 190 3245 191
rect 3306 191 3307 192
rect 3311 191 3312 195
rect 3306 190 3312 191
rect 3382 195 3389 196
rect 3382 191 3383 195
rect 3388 191 3389 195
rect 3382 190 3389 191
rect 3503 195 3509 196
rect 3503 191 3504 195
rect 3508 194 3509 195
rect 3518 195 3524 196
rect 3518 194 3519 195
rect 3508 192 3519 194
rect 3508 191 3509 192
rect 3503 190 3509 191
rect 3518 191 3519 192
rect 3523 191 3524 195
rect 3518 190 3524 191
rect 2494 179 2500 180
rect 2494 178 2495 179
rect 2180 176 2495 178
rect 1895 171 1901 172
rect 1895 167 1896 171
rect 1900 170 1901 171
rect 1962 171 1968 172
rect 1962 170 1963 171
rect 1900 168 1963 170
rect 1900 167 1901 168
rect 1895 166 1901 167
rect 1962 167 1963 168
rect 1967 167 1968 171
rect 1962 166 1968 167
rect 1975 171 1981 172
rect 1975 167 1976 171
rect 1980 170 1981 171
rect 2042 171 2048 172
rect 2042 170 2043 171
rect 1980 168 2043 170
rect 1980 167 1981 168
rect 1975 166 1981 167
rect 2042 167 2043 168
rect 2047 167 2048 171
rect 2042 166 2048 167
rect 2079 171 2085 172
rect 2079 167 2080 171
rect 2084 170 2085 171
rect 2180 170 2182 176
rect 2494 175 2495 176
rect 2499 175 2500 179
rect 2494 174 2500 175
rect 2084 168 2182 170
rect 2186 171 2192 172
rect 2084 167 2085 168
rect 2079 166 2085 167
rect 2186 167 2187 171
rect 2191 170 2192 171
rect 2207 171 2213 172
rect 2207 170 2208 171
rect 2191 168 2208 170
rect 2191 167 2192 168
rect 2186 166 2192 167
rect 2207 167 2208 168
rect 2212 167 2213 171
rect 2207 166 2213 167
rect 2318 171 2324 172
rect 2318 167 2319 171
rect 2323 170 2324 171
rect 2343 171 2349 172
rect 2343 170 2344 171
rect 2323 168 2344 170
rect 2323 167 2324 168
rect 2318 166 2324 167
rect 2343 167 2344 168
rect 2348 167 2349 171
rect 2343 166 2349 167
rect 2478 171 2485 172
rect 2478 167 2479 171
rect 2484 167 2485 171
rect 2478 166 2485 167
rect 2615 171 2621 172
rect 2615 167 2616 171
rect 2620 170 2621 171
rect 2623 171 2629 172
rect 2623 170 2624 171
rect 2620 168 2624 170
rect 2620 167 2621 168
rect 2615 166 2621 167
rect 2623 167 2624 168
rect 2628 167 2629 171
rect 2623 166 2629 167
rect 2674 171 2680 172
rect 2674 167 2675 171
rect 2679 170 2680 171
rect 2735 171 2741 172
rect 2735 170 2736 171
rect 2679 168 2736 170
rect 2679 167 2680 168
rect 2674 166 2680 167
rect 2735 167 2736 168
rect 2740 167 2741 171
rect 2735 166 2741 167
rect 2794 171 2800 172
rect 2794 167 2795 171
rect 2799 170 2800 171
rect 2847 171 2853 172
rect 2847 170 2848 171
rect 2799 168 2848 170
rect 2799 167 2800 168
rect 2794 166 2800 167
rect 2847 167 2848 168
rect 2852 167 2853 171
rect 2847 166 2853 167
rect 2906 171 2912 172
rect 2906 167 2907 171
rect 2911 170 2912 171
rect 2951 171 2957 172
rect 2951 170 2952 171
rect 2911 168 2952 170
rect 2911 167 2912 168
rect 2906 166 2912 167
rect 2951 167 2952 168
rect 2956 167 2957 171
rect 2951 166 2957 167
rect 3010 171 3016 172
rect 3010 167 3011 171
rect 3015 170 3016 171
rect 3055 171 3061 172
rect 3055 170 3056 171
rect 3015 168 3056 170
rect 3015 167 3016 168
rect 3010 166 3016 167
rect 3055 167 3056 168
rect 3060 167 3061 171
rect 3055 166 3061 167
rect 3114 171 3120 172
rect 3114 167 3115 171
rect 3119 170 3120 171
rect 3151 171 3157 172
rect 3151 170 3152 171
rect 3119 168 3152 170
rect 3119 167 3120 168
rect 3114 166 3120 167
rect 3151 167 3152 168
rect 3156 167 3157 171
rect 3151 166 3157 167
rect 3210 171 3216 172
rect 3210 167 3211 171
rect 3215 170 3216 171
rect 3239 171 3245 172
rect 3239 170 3240 171
rect 3215 168 3240 170
rect 3215 167 3216 168
rect 3210 166 3216 167
rect 3239 167 3240 168
rect 3244 167 3245 171
rect 3239 166 3245 167
rect 3298 171 3304 172
rect 3298 167 3299 171
rect 3303 170 3304 171
rect 3335 171 3341 172
rect 3335 170 3336 171
rect 3303 168 3336 170
rect 3303 167 3304 168
rect 3298 166 3304 167
rect 3335 167 3336 168
rect 3340 167 3341 171
rect 3335 166 3341 167
rect 3423 171 3429 172
rect 3423 167 3424 171
rect 3428 170 3429 171
rect 3490 171 3496 172
rect 3490 170 3491 171
rect 3428 168 3491 170
rect 3428 167 3429 168
rect 3423 166 3429 167
rect 3490 167 3491 168
rect 3495 167 3496 171
rect 3490 166 3496 167
rect 3502 171 3509 172
rect 3502 167 3503 171
rect 3508 167 3509 171
rect 3502 166 3509 167
rect 390 163 396 164
rect 390 162 391 163
rect 188 160 391 162
rect 135 155 141 156
rect 135 151 136 155
rect 140 154 141 155
rect 188 154 190 160
rect 390 159 391 160
rect 395 159 396 163
rect 790 163 796 164
rect 790 162 791 163
rect 390 158 396 159
rect 537 160 791 162
rect 537 156 539 160
rect 790 159 791 160
rect 795 159 796 163
rect 1110 163 1116 164
rect 1110 162 1111 163
rect 790 158 796 159
rect 908 160 1111 162
rect 140 152 190 154
rect 194 155 200 156
rect 140 151 141 152
rect 135 150 141 151
rect 194 151 195 155
rect 199 154 200 155
rect 215 155 221 156
rect 215 154 216 155
rect 199 152 216 154
rect 199 151 200 152
rect 194 150 200 151
rect 215 151 216 152
rect 220 151 221 155
rect 215 150 221 151
rect 274 155 280 156
rect 274 151 275 155
rect 279 154 280 155
rect 295 155 301 156
rect 295 154 296 155
rect 279 152 296 154
rect 279 151 280 152
rect 274 150 280 151
rect 295 151 296 152
rect 300 151 301 155
rect 295 150 301 151
rect 375 155 381 156
rect 375 151 376 155
rect 380 154 381 155
rect 442 155 448 156
rect 442 154 443 155
rect 380 152 443 154
rect 380 151 381 152
rect 375 150 381 151
rect 442 151 443 152
rect 447 151 448 155
rect 442 150 448 151
rect 455 155 461 156
rect 455 151 456 155
rect 460 154 461 155
rect 522 155 528 156
rect 522 154 523 155
rect 460 152 523 154
rect 460 151 461 152
rect 455 150 461 151
rect 522 151 523 152
rect 527 151 528 155
rect 522 150 528 151
rect 535 155 541 156
rect 535 151 536 155
rect 540 151 541 155
rect 535 150 541 151
rect 610 155 621 156
rect 610 151 611 155
rect 615 151 616 155
rect 620 151 621 155
rect 610 150 621 151
rect 674 155 680 156
rect 674 151 675 155
rect 679 154 680 155
rect 695 155 701 156
rect 695 154 696 155
rect 679 152 696 154
rect 679 151 680 152
rect 674 150 680 151
rect 695 151 696 152
rect 700 151 701 155
rect 695 150 701 151
rect 754 155 760 156
rect 754 151 755 155
rect 759 154 760 155
rect 775 155 781 156
rect 775 154 776 155
rect 759 152 776 154
rect 759 151 760 152
rect 754 150 760 151
rect 775 151 776 152
rect 780 151 781 155
rect 775 150 781 151
rect 855 155 861 156
rect 855 151 856 155
rect 860 154 861 155
rect 908 154 910 160
rect 1110 159 1111 160
rect 1115 159 1116 163
rect 1110 158 1116 159
rect 1902 162 1908 163
rect 1902 158 1903 162
rect 1907 158 1908 162
rect 1902 157 1908 158
rect 1982 162 1988 163
rect 1982 158 1983 162
rect 1987 158 1988 162
rect 1982 157 1988 158
rect 2086 162 2092 163
rect 2086 158 2087 162
rect 2091 158 2092 162
rect 2086 157 2092 158
rect 2214 162 2220 163
rect 2214 158 2215 162
rect 2219 158 2220 162
rect 2214 157 2220 158
rect 2350 162 2356 163
rect 2350 158 2351 162
rect 2355 158 2356 162
rect 2350 157 2356 158
rect 2486 162 2492 163
rect 2486 158 2487 162
rect 2491 158 2492 162
rect 2486 157 2492 158
rect 2622 162 2628 163
rect 2622 158 2623 162
rect 2627 158 2628 162
rect 2622 157 2628 158
rect 2742 162 2748 163
rect 2742 158 2743 162
rect 2747 158 2748 162
rect 2742 157 2748 158
rect 2854 162 2860 163
rect 2854 158 2855 162
rect 2859 158 2860 162
rect 2854 157 2860 158
rect 2958 162 2964 163
rect 2958 158 2959 162
rect 2963 158 2964 162
rect 2958 157 2964 158
rect 3062 162 3068 163
rect 3062 158 3063 162
rect 3067 158 3068 162
rect 3062 157 3068 158
rect 3158 162 3164 163
rect 3158 158 3159 162
rect 3163 158 3164 162
rect 3158 157 3164 158
rect 3246 162 3252 163
rect 3246 158 3247 162
rect 3251 158 3252 162
rect 3246 157 3252 158
rect 3342 162 3348 163
rect 3342 158 3343 162
rect 3347 158 3348 162
rect 3342 157 3348 158
rect 3430 162 3436 163
rect 3430 158 3431 162
rect 3435 158 3436 162
rect 3430 157 3436 158
rect 3510 162 3516 163
rect 3510 158 3511 162
rect 3515 158 3516 162
rect 3510 157 3516 158
rect 860 152 910 154
rect 914 155 920 156
rect 860 151 861 152
rect 855 150 861 151
rect 914 151 915 155
rect 919 154 920 155
rect 935 155 941 156
rect 935 154 936 155
rect 919 152 936 154
rect 919 151 920 152
rect 914 150 920 151
rect 935 151 936 152
rect 940 151 941 155
rect 935 150 941 151
rect 1006 155 1012 156
rect 1006 151 1007 155
rect 1011 154 1012 155
rect 1015 155 1021 156
rect 1015 154 1016 155
rect 1011 152 1016 154
rect 1011 151 1012 152
rect 1006 150 1012 151
rect 1015 151 1016 152
rect 1020 151 1021 155
rect 1015 150 1021 151
rect 1095 155 1101 156
rect 1095 151 1096 155
rect 1100 154 1101 155
rect 1162 155 1168 156
rect 1162 154 1163 155
rect 1100 152 1163 154
rect 1100 151 1101 152
rect 1095 150 1101 151
rect 1162 151 1163 152
rect 1167 151 1168 155
rect 1162 150 1168 151
rect 1175 155 1181 156
rect 1175 151 1176 155
rect 1180 154 1181 155
rect 1247 155 1253 156
rect 1247 154 1248 155
rect 1180 152 1248 154
rect 1180 151 1181 152
rect 1175 150 1181 151
rect 1247 151 1248 152
rect 1252 151 1253 155
rect 1247 150 1253 151
rect 1255 155 1261 156
rect 1255 151 1256 155
rect 1260 154 1261 155
rect 1322 155 1328 156
rect 1322 154 1323 155
rect 1260 152 1323 154
rect 1260 151 1261 152
rect 1255 150 1261 151
rect 1322 151 1323 152
rect 1327 151 1328 155
rect 1322 150 1328 151
rect 1335 155 1341 156
rect 1335 151 1336 155
rect 1340 154 1341 155
rect 1402 155 1408 156
rect 1402 154 1403 155
rect 1340 152 1403 154
rect 1340 151 1341 152
rect 1335 150 1341 151
rect 1402 151 1403 152
rect 1407 151 1408 155
rect 1402 150 1408 151
rect 1415 155 1421 156
rect 1415 151 1416 155
rect 1420 154 1421 155
rect 1487 155 1493 156
rect 1487 154 1488 155
rect 1420 152 1488 154
rect 1420 151 1421 152
rect 1415 150 1421 151
rect 1487 151 1488 152
rect 1492 151 1493 155
rect 1487 150 1493 151
rect 1503 155 1509 156
rect 1503 151 1504 155
rect 1508 154 1509 155
rect 1570 155 1576 156
rect 1570 154 1571 155
rect 1508 152 1571 154
rect 1508 151 1509 152
rect 1503 150 1509 151
rect 1570 151 1571 152
rect 1575 151 1576 155
rect 1570 150 1576 151
rect 1583 155 1589 156
rect 1583 151 1584 155
rect 1588 154 1589 155
rect 1650 155 1656 156
rect 1650 154 1651 155
rect 1588 152 1651 154
rect 1588 151 1589 152
rect 1583 150 1589 151
rect 1650 151 1651 152
rect 1655 151 1656 155
rect 1650 150 1656 151
rect 1663 155 1669 156
rect 1663 151 1664 155
rect 1668 154 1669 155
rect 1730 155 1736 156
rect 1730 154 1731 155
rect 1668 152 1731 154
rect 1668 151 1669 152
rect 1663 150 1669 151
rect 1730 151 1731 152
rect 1735 151 1736 155
rect 1730 150 1736 151
rect 1743 155 1749 156
rect 1743 151 1744 155
rect 1748 154 1749 155
rect 1802 155 1808 156
rect 1802 154 1803 155
rect 1748 152 1803 154
rect 1748 151 1749 152
rect 1743 150 1749 151
rect 1802 151 1803 152
rect 1807 151 1808 155
rect 1802 150 1808 151
rect 142 146 148 147
rect 142 142 143 146
rect 147 142 148 146
rect 142 141 148 142
rect 222 146 228 147
rect 222 142 223 146
rect 227 142 228 146
rect 222 141 228 142
rect 302 146 308 147
rect 302 142 303 146
rect 307 142 308 146
rect 302 141 308 142
rect 382 146 388 147
rect 382 142 383 146
rect 387 142 388 146
rect 382 141 388 142
rect 462 146 468 147
rect 462 142 463 146
rect 467 142 468 146
rect 462 141 468 142
rect 542 146 548 147
rect 542 142 543 146
rect 547 142 548 146
rect 542 141 548 142
rect 622 146 628 147
rect 622 142 623 146
rect 627 142 628 146
rect 622 141 628 142
rect 702 146 708 147
rect 702 142 703 146
rect 707 142 708 146
rect 702 141 708 142
rect 782 146 788 147
rect 782 142 783 146
rect 787 142 788 146
rect 782 141 788 142
rect 862 146 868 147
rect 862 142 863 146
rect 867 142 868 146
rect 862 141 868 142
rect 942 146 948 147
rect 942 142 943 146
rect 947 142 948 146
rect 942 141 948 142
rect 1022 146 1028 147
rect 1022 142 1023 146
rect 1027 142 1028 146
rect 1022 141 1028 142
rect 1102 146 1108 147
rect 1102 142 1103 146
rect 1107 142 1108 146
rect 1102 141 1108 142
rect 1182 146 1188 147
rect 1182 142 1183 146
rect 1187 142 1188 146
rect 1182 141 1188 142
rect 1262 146 1268 147
rect 1262 142 1263 146
rect 1267 142 1268 146
rect 1262 141 1268 142
rect 1342 146 1348 147
rect 1342 142 1343 146
rect 1347 142 1348 146
rect 1342 141 1348 142
rect 1422 146 1428 147
rect 1422 142 1423 146
rect 1427 142 1428 146
rect 1422 141 1428 142
rect 1510 146 1516 147
rect 1510 142 1511 146
rect 1515 142 1516 146
rect 1510 141 1516 142
rect 1590 146 1596 147
rect 1590 142 1591 146
rect 1595 142 1596 146
rect 1590 141 1596 142
rect 1670 146 1676 147
rect 1670 142 1671 146
rect 1675 142 1676 146
rect 1670 141 1676 142
rect 1750 146 1756 147
rect 1750 142 1751 146
rect 1755 142 1756 146
rect 1750 141 1756 142
rect 1870 144 1876 145
rect 1870 140 1871 144
rect 1875 140 1876 144
rect 1870 139 1876 140
rect 3590 144 3596 145
rect 3590 140 3591 144
rect 3595 140 3596 144
rect 3590 139 3596 140
rect 1802 135 1808 136
rect 1802 131 1803 135
rect 1807 134 1808 135
rect 1962 135 1968 136
rect 1807 132 1913 134
rect 1807 131 1808 132
rect 1802 130 1808 131
rect 1962 131 1963 135
rect 1967 134 1968 135
rect 2042 135 2048 136
rect 1967 132 1993 134
rect 1967 131 1968 132
rect 1962 130 1968 131
rect 2042 131 2043 135
rect 2047 134 2048 135
rect 2318 135 2324 136
rect 2318 134 2319 135
rect 2047 132 2097 134
rect 2269 132 2319 134
rect 2047 131 2048 132
rect 2042 130 2048 131
rect 2318 131 2319 132
rect 2323 131 2324 135
rect 2478 135 2484 136
rect 2478 134 2479 135
rect 2405 132 2479 134
rect 2318 130 2324 131
rect 2478 131 2479 132
rect 2483 131 2484 135
rect 2478 130 2484 131
rect 2494 135 2500 136
rect 2494 131 2495 135
rect 2499 131 2500 135
rect 2494 130 2500 131
rect 2674 135 2680 136
rect 2674 131 2675 135
rect 2679 131 2680 135
rect 2674 130 2680 131
rect 2794 135 2800 136
rect 2794 131 2795 135
rect 2799 131 2800 135
rect 2794 130 2800 131
rect 2906 135 2912 136
rect 2906 131 2907 135
rect 2911 131 2912 135
rect 2906 130 2912 131
rect 3010 135 3016 136
rect 3010 131 3011 135
rect 3015 131 3016 135
rect 3010 130 3016 131
rect 3114 135 3120 136
rect 3114 131 3115 135
rect 3119 131 3120 135
rect 3114 130 3120 131
rect 3210 135 3216 136
rect 3210 131 3211 135
rect 3215 131 3216 135
rect 3210 130 3216 131
rect 3298 135 3304 136
rect 3298 131 3299 135
rect 3303 131 3304 135
rect 3298 130 3304 131
rect 3382 135 3388 136
rect 3382 131 3383 135
rect 3387 131 3388 135
rect 3382 130 3388 131
rect 3490 135 3496 136
rect 3490 131 3491 135
rect 3495 134 3496 135
rect 3495 132 3521 134
rect 3495 131 3496 132
rect 3490 130 3496 131
rect 110 128 116 129
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 1830 128 1836 129
rect 1830 124 1831 128
rect 1835 124 1836 128
rect 1830 123 1836 124
rect 1870 127 1876 128
rect 1870 123 1871 127
rect 1875 123 1876 127
rect 3590 127 3596 128
rect 1870 122 1876 123
rect 1894 124 1900 125
rect 1894 120 1895 124
rect 1899 120 1900 124
rect 194 119 200 120
rect 194 115 195 119
rect 199 115 200 119
rect 194 114 200 115
rect 274 119 280 120
rect 274 115 275 119
rect 279 115 280 119
rect 274 114 280 115
rect 354 119 360 120
rect 354 115 355 119
rect 359 115 360 119
rect 354 114 360 115
rect 390 119 396 120
rect 390 115 391 119
rect 395 115 396 119
rect 390 114 396 115
rect 442 119 448 120
rect 442 115 443 119
rect 447 118 448 119
rect 522 119 528 120
rect 447 116 473 118
rect 447 115 448 116
rect 442 114 448 115
rect 522 115 523 119
rect 527 118 528 119
rect 674 119 680 120
rect 527 116 553 118
rect 527 115 528 116
rect 522 114 528 115
rect 674 115 675 119
rect 679 115 680 119
rect 674 114 680 115
rect 754 119 760 120
rect 754 115 755 119
rect 759 115 760 119
rect 754 114 760 115
rect 790 119 796 120
rect 790 115 791 119
rect 795 115 796 119
rect 790 114 796 115
rect 914 119 920 120
rect 914 115 915 119
rect 919 115 920 119
rect 1006 119 1012 120
rect 1006 118 1007 119
rect 997 116 1007 118
rect 914 114 920 115
rect 1006 115 1007 116
rect 1011 115 1012 119
rect 1006 114 1012 115
rect 1074 119 1080 120
rect 1074 115 1075 119
rect 1079 115 1080 119
rect 1074 114 1080 115
rect 1110 119 1116 120
rect 1110 115 1111 119
rect 1115 115 1116 119
rect 1110 114 1116 115
rect 1162 119 1168 120
rect 1162 115 1163 119
rect 1167 118 1168 119
rect 1247 119 1253 120
rect 1167 116 1193 118
rect 1167 115 1168 116
rect 1162 114 1168 115
rect 1247 115 1248 119
rect 1252 118 1253 119
rect 1322 119 1328 120
rect 1252 116 1273 118
rect 1252 115 1253 116
rect 1247 114 1253 115
rect 1322 115 1323 119
rect 1327 118 1328 119
rect 1402 119 1408 120
rect 1327 116 1353 118
rect 1327 115 1328 116
rect 1322 114 1328 115
rect 1402 115 1403 119
rect 1407 118 1408 119
rect 1487 119 1493 120
rect 1407 116 1433 118
rect 1407 115 1408 116
rect 1402 114 1408 115
rect 1487 115 1488 119
rect 1492 118 1493 119
rect 1570 119 1576 120
rect 1492 116 1521 118
rect 1492 115 1493 116
rect 1487 114 1493 115
rect 1570 115 1571 119
rect 1575 118 1576 119
rect 1650 119 1656 120
rect 1575 116 1601 118
rect 1575 115 1576 116
rect 1570 114 1576 115
rect 1650 115 1651 119
rect 1655 118 1656 119
rect 1730 119 1736 120
rect 1894 119 1900 120
rect 1974 124 1980 125
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 2078 124 2084 125
rect 2078 120 2079 124
rect 2083 120 2084 124
rect 2078 119 2084 120
rect 2206 124 2212 125
rect 2206 120 2207 124
rect 2211 120 2212 124
rect 2206 119 2212 120
rect 2342 124 2348 125
rect 2342 120 2343 124
rect 2347 120 2348 124
rect 2342 119 2348 120
rect 2478 124 2484 125
rect 2478 120 2479 124
rect 2483 120 2484 124
rect 2478 119 2484 120
rect 2614 124 2620 125
rect 2614 120 2615 124
rect 2619 120 2620 124
rect 2614 119 2620 120
rect 2734 124 2740 125
rect 2734 120 2735 124
rect 2739 120 2740 124
rect 2734 119 2740 120
rect 2846 124 2852 125
rect 2846 120 2847 124
rect 2851 120 2852 124
rect 2846 119 2852 120
rect 2950 124 2956 125
rect 2950 120 2951 124
rect 2955 120 2956 124
rect 2950 119 2956 120
rect 3054 124 3060 125
rect 3054 120 3055 124
rect 3059 120 3060 124
rect 3054 119 3060 120
rect 3150 124 3156 125
rect 3150 120 3151 124
rect 3155 120 3156 124
rect 3150 119 3156 120
rect 3238 124 3244 125
rect 3238 120 3239 124
rect 3243 120 3244 124
rect 3238 119 3244 120
rect 3334 124 3340 125
rect 3334 120 3335 124
rect 3339 120 3340 124
rect 3334 119 3340 120
rect 3422 124 3428 125
rect 3422 120 3423 124
rect 3427 120 3428 124
rect 3422 119 3428 120
rect 3502 124 3508 125
rect 3502 120 3503 124
rect 3507 120 3508 124
rect 3590 123 3591 127
rect 3595 123 3596 127
rect 3590 122 3596 123
rect 3502 119 3508 120
rect 1655 116 1681 118
rect 1655 115 1656 116
rect 1650 114 1656 115
rect 1730 115 1731 119
rect 1735 118 1736 119
rect 1735 116 1761 118
rect 1735 115 1736 116
rect 1730 114 1736 115
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 1830 111 1836 112
rect 110 106 116 107
rect 134 108 140 109
rect 134 104 135 108
rect 139 104 140 108
rect 134 103 140 104
rect 214 108 220 109
rect 214 104 215 108
rect 219 104 220 108
rect 214 103 220 104
rect 294 108 300 109
rect 294 104 295 108
rect 299 104 300 108
rect 294 103 300 104
rect 374 108 380 109
rect 374 104 375 108
rect 379 104 380 108
rect 374 103 380 104
rect 454 108 460 109
rect 454 104 455 108
rect 459 104 460 108
rect 454 103 460 104
rect 534 108 540 109
rect 534 104 535 108
rect 539 104 540 108
rect 534 103 540 104
rect 614 108 620 109
rect 614 104 615 108
rect 619 104 620 108
rect 614 103 620 104
rect 694 108 700 109
rect 694 104 695 108
rect 699 104 700 108
rect 694 103 700 104
rect 774 108 780 109
rect 774 104 775 108
rect 779 104 780 108
rect 774 103 780 104
rect 854 108 860 109
rect 854 104 855 108
rect 859 104 860 108
rect 854 103 860 104
rect 934 108 940 109
rect 934 104 935 108
rect 939 104 940 108
rect 934 103 940 104
rect 1014 108 1020 109
rect 1014 104 1015 108
rect 1019 104 1020 108
rect 1014 103 1020 104
rect 1094 108 1100 109
rect 1094 104 1095 108
rect 1099 104 1100 108
rect 1094 103 1100 104
rect 1174 108 1180 109
rect 1174 104 1175 108
rect 1179 104 1180 108
rect 1174 103 1180 104
rect 1254 108 1260 109
rect 1254 104 1255 108
rect 1259 104 1260 108
rect 1254 103 1260 104
rect 1334 108 1340 109
rect 1334 104 1335 108
rect 1339 104 1340 108
rect 1334 103 1340 104
rect 1414 108 1420 109
rect 1414 104 1415 108
rect 1419 104 1420 108
rect 1414 103 1420 104
rect 1502 108 1508 109
rect 1502 104 1503 108
rect 1507 104 1508 108
rect 1502 103 1508 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1662 108 1668 109
rect 1662 104 1663 108
rect 1667 104 1668 108
rect 1662 103 1668 104
rect 1742 108 1748 109
rect 1742 104 1743 108
rect 1747 104 1748 108
rect 1830 107 1831 111
rect 1835 107 1836 111
rect 1830 106 1836 107
rect 1742 103 1748 104
<< m3c >>
rect 111 3641 115 3645
rect 135 3644 139 3648
rect 215 3644 219 3648
rect 295 3644 299 3648
rect 1831 3641 1835 3645
rect 135 3631 139 3635
rect 203 3635 207 3639
rect 283 3635 287 3639
rect 111 3624 115 3628
rect 1831 3624 1835 3628
rect 143 3606 147 3610
rect 223 3606 227 3610
rect 303 3606 307 3610
rect 203 3595 207 3599
rect 283 3595 287 3599
rect 2071 3591 2075 3595
rect 2115 3591 2119 3595
rect 2203 3591 2207 3595
rect 2307 3591 2311 3595
rect 2419 3591 2423 3595
rect 2531 3591 2535 3595
rect 2827 3599 2831 3603
rect 2755 3591 2759 3595
rect 2867 3591 2871 3595
rect 2971 3591 2975 3595
rect 3067 3591 3071 3595
rect 3163 3591 3167 3595
rect 3259 3591 3263 3595
rect 3355 3591 3359 3595
rect 135 3583 136 3587
rect 136 3583 139 3587
rect 195 3583 199 3587
rect 275 3583 279 3587
rect 395 3583 399 3587
rect 523 3583 527 3587
rect 659 3583 663 3587
rect 887 3583 891 3587
rect 931 3583 935 3587
rect 1051 3583 1055 3587
rect 1163 3583 1167 3587
rect 1275 3583 1279 3587
rect 1379 3583 1383 3587
rect 1475 3583 1479 3587
rect 1579 3583 1583 3587
rect 2063 3582 2067 3586
rect 2151 3582 2155 3586
rect 2255 3582 2259 3586
rect 2367 3582 2371 3586
rect 2479 3582 2483 3586
rect 2591 3582 2595 3586
rect 2703 3582 2707 3586
rect 2815 3582 2819 3586
rect 2919 3582 2923 3586
rect 3015 3582 3019 3586
rect 3111 3582 3115 3586
rect 3207 3582 3211 3586
rect 3303 3582 3307 3586
rect 3399 3582 3403 3586
rect 143 3574 147 3578
rect 223 3574 227 3578
rect 343 3574 347 3578
rect 471 3574 475 3578
rect 607 3574 611 3578
rect 743 3574 747 3578
rect 879 3574 883 3578
rect 999 3574 1003 3578
rect 1111 3574 1115 3578
rect 1223 3574 1227 3578
rect 1327 3574 1331 3578
rect 1423 3574 1427 3578
rect 1527 3574 1531 3578
rect 1631 3574 1635 3578
rect 1871 3564 1875 3568
rect 3591 3564 3595 3568
rect 111 3556 115 3560
rect 1831 3556 1835 3560
rect 2115 3555 2119 3559
rect 2203 3555 2207 3559
rect 2307 3555 2311 3559
rect 2419 3555 2423 3559
rect 2531 3555 2535 3559
rect 2755 3555 2759 3559
rect 2867 3555 2871 3559
rect 2971 3555 2975 3559
rect 3067 3555 3071 3559
rect 3163 3555 3167 3559
rect 3259 3555 3263 3559
rect 3355 3555 3359 3559
rect 195 3547 199 3551
rect 275 3547 279 3551
rect 395 3547 399 3551
rect 523 3547 527 3551
rect 659 3547 663 3551
rect 767 3547 771 3551
rect 931 3547 935 3551
rect 1051 3547 1055 3551
rect 1163 3547 1167 3551
rect 1275 3547 1279 3551
rect 1379 3547 1383 3551
rect 1475 3547 1479 3551
rect 1579 3547 1583 3551
rect 1871 3547 1875 3551
rect 2055 3544 2059 3548
rect 111 3539 115 3543
rect 2143 3544 2147 3548
rect 2247 3544 2251 3548
rect 2359 3544 2363 3548
rect 2471 3544 2475 3548
rect 2583 3544 2587 3548
rect 2695 3544 2699 3548
rect 2807 3544 2811 3548
rect 2911 3544 2915 3548
rect 3007 3544 3011 3548
rect 3103 3544 3107 3548
rect 3199 3544 3203 3548
rect 3295 3544 3299 3548
rect 3391 3544 3395 3548
rect 3591 3547 3595 3551
rect 135 3536 139 3540
rect 215 3536 219 3540
rect 335 3536 339 3540
rect 463 3536 467 3540
rect 599 3536 603 3540
rect 735 3536 739 3540
rect 871 3536 875 3540
rect 991 3536 995 3540
rect 1103 3536 1107 3540
rect 1215 3536 1219 3540
rect 1319 3536 1323 3540
rect 1415 3536 1419 3540
rect 1519 3536 1523 3540
rect 1623 3536 1627 3540
rect 1831 3539 1835 3543
rect 2383 3527 2387 3531
rect 3135 3527 3139 3531
rect 1583 3519 1587 3523
rect 1871 3497 1875 3501
rect 2087 3500 2091 3504
rect 2167 3500 2171 3504
rect 2263 3500 2267 3504
rect 2367 3500 2371 3504
rect 2487 3500 2491 3504
rect 2615 3500 2619 3504
rect 2743 3500 2747 3504
rect 2871 3500 2875 3504
rect 2991 3500 2995 3504
rect 3119 3500 3123 3504
rect 3247 3500 3251 3504
rect 3375 3500 3379 3504
rect 111 3489 115 3493
rect 191 3492 195 3496
rect 327 3492 331 3496
rect 471 3492 475 3496
rect 623 3492 627 3496
rect 775 3492 779 3496
rect 919 3492 923 3496
rect 1055 3492 1059 3496
rect 1183 3492 1187 3496
rect 1311 3492 1315 3496
rect 1439 3492 1443 3496
rect 3591 3497 3595 3501
rect 1567 3492 1571 3496
rect 1831 3489 1835 3493
rect 2071 3491 2075 3495
rect 2155 3491 2159 3495
rect 2235 3491 2239 3495
rect 2435 3491 2439 3495
rect 2559 3491 2563 3495
rect 2687 3491 2691 3495
rect 2827 3491 2831 3495
rect 2939 3491 2943 3495
rect 3319 3491 3323 3495
rect 259 3483 263 3487
rect 395 3483 399 3487
rect 539 3483 543 3487
rect 691 3483 695 3487
rect 887 3483 891 3487
rect 987 3483 991 3487
rect 1127 3483 1131 3487
rect 1379 3483 1383 3487
rect 1871 3480 1875 3484
rect 3435 3483 3439 3487
rect 3591 3480 3595 3484
rect 111 3472 115 3476
rect 1831 3472 1835 3476
rect 2095 3462 2099 3466
rect 2175 3462 2179 3466
rect 2271 3462 2275 3466
rect 2375 3462 2379 3466
rect 2495 3462 2499 3466
rect 2623 3462 2627 3466
rect 2751 3462 2755 3466
rect 2879 3462 2883 3466
rect 2999 3462 3003 3466
rect 3127 3462 3131 3466
rect 3255 3462 3259 3466
rect 3383 3462 3387 3466
rect 199 3454 203 3458
rect 335 3454 339 3458
rect 479 3454 483 3458
rect 631 3454 635 3458
rect 783 3454 787 3458
rect 927 3454 931 3458
rect 1063 3454 1067 3458
rect 1191 3454 1195 3458
rect 1319 3454 1323 3458
rect 1447 3454 1451 3458
rect 1575 3454 1579 3458
rect 2155 3451 2159 3455
rect 2235 3451 2239 3455
rect 2251 3451 2255 3455
rect 2383 3451 2387 3455
rect 2435 3451 2439 3455
rect 2559 3451 2563 3455
rect 2687 3451 2691 3455
rect 2939 3451 2943 3455
rect 2991 3451 2992 3455
rect 2992 3451 2995 3455
rect 3135 3451 3139 3455
rect 3319 3451 3323 3455
rect 259 3443 263 3447
rect 395 3443 399 3447
rect 539 3443 543 3447
rect 691 3443 695 3447
rect 767 3443 771 3447
rect 987 3443 991 3447
rect 1127 3443 1131 3447
rect 1171 3443 1175 3447
rect 1379 3443 1383 3447
rect 1583 3443 1587 3447
rect 287 3431 288 3435
rect 288 3431 291 3435
rect 347 3431 351 3435
rect 507 3431 511 3435
rect 675 3431 679 3435
rect 1011 3431 1015 3435
rect 1351 3431 1355 3435
rect 1467 3431 1471 3435
rect 1611 3431 1615 3435
rect 2155 3431 2159 3435
rect 2163 3431 2167 3435
rect 2295 3431 2296 3435
rect 2296 3431 2299 3435
rect 2423 3431 2427 3435
rect 2603 3431 2607 3435
rect 2739 3431 2743 3435
rect 3031 3431 3035 3435
rect 3135 3431 3139 3435
rect 3435 3431 3439 3435
rect 151 3422 155 3426
rect 295 3422 299 3426
rect 455 3422 459 3426
rect 623 3422 627 3426
rect 791 3422 795 3426
rect 959 3422 963 3426
rect 1119 3422 1123 3426
rect 1271 3422 1275 3426
rect 1415 3422 1419 3426
rect 1559 3422 1563 3426
rect 1711 3422 1715 3426
rect 2111 3422 2115 3426
rect 2199 3422 2203 3426
rect 2303 3422 2307 3426
rect 2415 3422 2419 3426
rect 2543 3422 2547 3426
rect 2679 3422 2683 3426
rect 2815 3422 2819 3426
rect 2959 3422 2963 3426
rect 3111 3422 3115 3426
rect 3263 3422 3267 3426
rect 3423 3422 3427 3426
rect 111 3404 115 3408
rect 1831 3404 1835 3408
rect 1871 3404 1875 3408
rect 3591 3404 3595 3408
rect 287 3395 291 3399
rect 347 3395 351 3399
rect 507 3395 511 3399
rect 675 3395 679 3399
rect 1011 3395 1015 3399
rect 1171 3395 1175 3399
rect 1351 3395 1355 3399
rect 1467 3395 1471 3399
rect 1611 3395 1615 3399
rect 1735 3395 1739 3399
rect 2163 3395 2167 3399
rect 2251 3395 2255 3399
rect 2295 3399 2299 3403
rect 2575 3395 2579 3399
rect 2603 3395 2607 3399
rect 2739 3395 2743 3399
rect 2991 3395 2995 3399
rect 3031 3395 3035 3399
rect 3303 3395 3307 3399
rect 111 3387 115 3391
rect 143 3384 147 3388
rect 287 3384 291 3388
rect 447 3384 451 3388
rect 615 3384 619 3388
rect 783 3384 787 3388
rect 951 3384 955 3388
rect 1111 3384 1115 3388
rect 1263 3384 1267 3388
rect 1407 3384 1411 3388
rect 1551 3384 1555 3388
rect 1703 3384 1707 3388
rect 1831 3387 1835 3391
rect 1871 3387 1875 3391
rect 2103 3384 2107 3388
rect 2191 3384 2195 3388
rect 2295 3384 2299 3388
rect 2407 3384 2411 3388
rect 2535 3384 2539 3388
rect 2671 3384 2675 3388
rect 2807 3384 2811 3388
rect 2951 3384 2955 3388
rect 3103 3384 3107 3388
rect 3255 3384 3259 3388
rect 3415 3384 3419 3388
rect 3591 3387 3595 3391
rect 679 3367 683 3371
rect 2155 3367 2159 3371
rect 111 3337 115 3341
rect 207 3340 211 3344
rect 335 3340 339 3344
rect 471 3340 475 3344
rect 623 3340 627 3344
rect 783 3340 787 3344
rect 943 3340 947 3344
rect 1103 3340 1107 3344
rect 1263 3340 1267 3344
rect 1423 3340 1427 3344
rect 1583 3340 1587 3344
rect 1743 3340 1747 3344
rect 1831 3337 1835 3341
rect 279 3331 283 3335
rect 411 3331 415 3335
rect 707 3331 711 3335
rect 111 3320 115 3324
rect 395 3323 399 3327
rect 1011 3331 1015 3335
rect 1171 3331 1175 3335
rect 1651 3331 1655 3335
rect 1871 3333 1875 3337
rect 2127 3336 2131 3340
rect 2223 3336 2227 3340
rect 2335 3336 2339 3340
rect 2455 3336 2459 3340
rect 2583 3336 2587 3340
rect 2719 3336 2723 3340
rect 2863 3336 2867 3340
rect 3007 3336 3011 3340
rect 3159 3336 3163 3340
rect 3311 3336 3315 3340
rect 3471 3336 3475 3340
rect 3591 3333 3595 3337
rect 2195 3327 2199 3331
rect 2291 3327 2295 3331
rect 2403 3327 2407 3331
rect 2423 3327 2427 3331
rect 2651 3327 2655 3331
rect 2799 3327 2803 3331
rect 3135 3327 3139 3331
rect 3395 3327 3399 3331
rect 1831 3320 1835 3324
rect 1871 3316 1875 3320
rect 3531 3319 3535 3323
rect 3591 3316 3595 3320
rect 215 3302 219 3306
rect 343 3302 347 3306
rect 479 3302 483 3306
rect 631 3302 635 3306
rect 791 3302 795 3306
rect 951 3302 955 3306
rect 1111 3302 1115 3306
rect 1271 3302 1275 3306
rect 1431 3302 1435 3306
rect 1591 3302 1595 3306
rect 1751 3302 1755 3306
rect 2135 3298 2139 3302
rect 2231 3298 2235 3302
rect 2343 3298 2347 3302
rect 2463 3298 2467 3302
rect 2591 3298 2595 3302
rect 2727 3298 2731 3302
rect 2871 3298 2875 3302
rect 3015 3298 3019 3302
rect 3167 3298 3171 3302
rect 3319 3298 3323 3302
rect 3479 3298 3483 3302
rect 223 3291 227 3295
rect 279 3291 283 3295
rect 411 3291 415 3295
rect 707 3291 711 3295
rect 1011 3291 1015 3295
rect 1171 3291 1175 3295
rect 1263 3291 1264 3295
rect 1264 3291 1267 3295
rect 1651 3291 1655 3295
rect 1735 3291 1739 3295
rect 2143 3287 2147 3291
rect 2195 3287 2199 3291
rect 2291 3287 2295 3291
rect 2403 3287 2407 3291
rect 2575 3287 2579 3291
rect 2651 3287 2655 3291
rect 2799 3287 2803 3291
rect 3007 3287 3008 3291
rect 3008 3287 3011 3291
rect 3303 3287 3307 3291
rect 3395 3287 3399 3291
rect 395 3275 399 3279
rect 403 3275 407 3279
rect 507 3275 511 3279
rect 755 3275 759 3279
rect 991 3275 995 3279
rect 1035 3275 1039 3279
rect 1171 3275 1175 3279
rect 1563 3275 1567 3279
rect 1691 3275 1695 3279
rect 351 3266 355 3270
rect 455 3266 459 3270
rect 575 3266 579 3270
rect 703 3266 707 3270
rect 839 3266 843 3270
rect 983 3266 987 3270
rect 1119 3266 1123 3270
rect 1255 3266 1259 3270
rect 1383 3266 1387 3270
rect 1511 3266 1515 3270
rect 1639 3266 1643 3270
rect 1751 3266 1755 3270
rect 2423 3271 2427 3275
rect 2255 3263 2259 3267
rect 2331 3263 2335 3267
rect 2611 3263 2615 3267
rect 2747 3263 2751 3267
rect 3023 3263 3027 3267
rect 3187 3263 3191 3267
rect 3267 3263 3271 3267
rect 3435 3263 3439 3267
rect 3531 3263 3535 3267
rect 2135 3254 2139 3258
rect 2279 3254 2283 3258
rect 2415 3254 2419 3258
rect 2551 3254 2555 3258
rect 2687 3254 2691 3258
rect 2823 3254 2827 3258
rect 2959 3254 2963 3258
rect 3095 3254 3099 3258
rect 3231 3254 3235 3258
rect 3375 3254 3379 3258
rect 3511 3254 3515 3258
rect 111 3248 115 3252
rect 1831 3248 1835 3252
rect 403 3239 407 3243
rect 507 3239 511 3243
rect 755 3239 759 3243
rect 1035 3239 1039 3243
rect 1171 3239 1175 3243
rect 1263 3239 1267 3243
rect 1563 3239 1567 3243
rect 1691 3239 1695 3243
rect 1871 3236 1875 3240
rect 111 3231 115 3235
rect 3591 3236 3595 3240
rect 343 3228 347 3232
rect 447 3228 451 3232
rect 567 3228 571 3232
rect 695 3228 699 3232
rect 831 3228 835 3232
rect 975 3228 979 3232
rect 1111 3228 1115 3232
rect 1247 3228 1251 3232
rect 1375 3228 1379 3232
rect 1503 3228 1507 3232
rect 1631 3228 1635 3232
rect 1743 3228 1747 3232
rect 1831 3231 1835 3235
rect 2143 3227 2147 3231
rect 2331 3227 2335 3231
rect 2423 3227 2427 3231
rect 2611 3227 2615 3231
rect 2747 3227 2751 3231
rect 3007 3227 3011 3231
rect 3023 3227 3027 3231
rect 3187 3227 3191 3231
rect 3427 3227 3431 3231
rect 3435 3227 3439 3231
rect 1871 3219 1875 3223
rect 2127 3216 2131 3220
rect 503 3211 507 3215
rect 2271 3216 2275 3220
rect 2407 3216 2411 3220
rect 2543 3216 2547 3220
rect 2679 3216 2683 3220
rect 2815 3216 2819 3220
rect 2951 3216 2955 3220
rect 3087 3216 3091 3220
rect 3223 3216 3227 3220
rect 3367 3216 3371 3220
rect 3503 3216 3507 3220
rect 3591 3219 3595 3223
rect 1759 3211 1760 3215
rect 1760 3211 1763 3215
rect 2551 3199 2555 3203
rect 111 3181 115 3185
rect 487 3184 491 3188
rect 575 3184 579 3188
rect 663 3184 667 3188
rect 767 3184 771 3188
rect 887 3184 891 3188
rect 1023 3184 1027 3188
rect 1191 3184 1195 3188
rect 1375 3184 1379 3188
rect 1567 3184 1571 3188
rect 1743 3184 1747 3188
rect 1831 3181 1835 3185
rect 555 3175 559 3179
rect 643 3175 647 3179
rect 731 3175 735 3179
rect 835 3175 839 3179
rect 843 3175 847 3179
rect 991 3175 995 3179
rect 1107 3175 1111 3179
rect 1479 3175 1483 3179
rect 1487 3175 1491 3179
rect 1819 3175 1823 3179
rect 111 3164 115 3168
rect 1831 3164 1835 3168
rect 1871 3165 1875 3169
rect 1895 3168 1899 3172
rect 1991 3168 1995 3172
rect 2119 3168 2123 3172
rect 2247 3168 2251 3172
rect 2383 3168 2387 3172
rect 2511 3168 2515 3172
rect 2639 3168 2643 3172
rect 2767 3168 2771 3172
rect 2895 3168 2899 3172
rect 3031 3168 3035 3172
rect 3175 3168 3179 3172
rect 3327 3168 3331 3172
rect 3487 3168 3491 3172
rect 3591 3165 3595 3169
rect 1963 3159 1967 3163
rect 2063 3159 2067 3163
rect 495 3146 499 3150
rect 583 3146 587 3150
rect 671 3146 675 3150
rect 775 3146 779 3150
rect 895 3146 899 3150
rect 1031 3146 1035 3150
rect 1199 3146 1203 3150
rect 1383 3146 1387 3150
rect 1575 3146 1579 3150
rect 1751 3146 1755 3150
rect 1871 3148 1875 3152
rect 2179 3151 2183 3155
rect 2255 3155 2259 3159
rect 2351 3159 2355 3163
rect 2583 3159 2587 3163
rect 2711 3159 2715 3163
rect 2839 3159 2843 3163
rect 2971 3159 2975 3163
rect 3099 3159 3103 3163
rect 3259 3159 3263 3163
rect 3267 3159 3271 3163
rect 3239 3151 3243 3155
rect 3591 3148 3595 3152
rect 503 3135 507 3139
rect 555 3135 559 3139
rect 643 3135 647 3139
rect 731 3135 735 3139
rect 835 3135 839 3139
rect 1107 3135 1111 3139
rect 1207 3135 1211 3139
rect 1391 3135 1395 3139
rect 1479 3135 1483 3139
rect 1759 3135 1763 3139
rect 1903 3130 1907 3134
rect 1999 3130 2003 3134
rect 2127 3130 2131 3134
rect 2255 3130 2259 3134
rect 2391 3130 2395 3134
rect 2519 3130 2523 3134
rect 2647 3130 2651 3134
rect 2775 3130 2779 3134
rect 2903 3130 2907 3134
rect 3039 3130 3043 3134
rect 3183 3130 3187 3134
rect 3335 3130 3339 3134
rect 3495 3130 3499 3134
rect 635 3119 639 3123
rect 643 3119 647 3123
rect 723 3119 727 3123
rect 811 3119 815 3123
rect 927 3119 928 3123
rect 928 3119 931 3123
rect 1067 3119 1071 3123
rect 1075 3119 1079 3123
rect 1163 3119 1167 3123
rect 1251 3119 1255 3123
rect 1339 3119 1343 3123
rect 1819 3119 1823 3123
rect 1963 3119 1967 3123
rect 2063 3119 2067 3123
rect 2351 3119 2355 3123
rect 2415 3119 2419 3123
rect 2551 3119 2555 3123
rect 2583 3119 2587 3123
rect 2711 3119 2715 3123
rect 2839 3119 2843 3123
rect 2971 3119 2975 3123
rect 3099 3119 3103 3123
rect 3259 3119 3263 3123
rect 3427 3119 3431 3123
rect 591 3110 595 3114
rect 671 3110 675 3114
rect 759 3110 763 3114
rect 847 3110 851 3114
rect 935 3110 939 3114
rect 1023 3110 1027 3114
rect 1111 3110 1115 3114
rect 1199 3110 1203 3114
rect 1287 3110 1291 3114
rect 1375 3110 1379 3114
rect 111 3092 115 3096
rect 1831 3092 1835 3096
rect 1911 3091 1915 3095
rect 1955 3091 1959 3095
rect 2179 3091 2183 3095
rect 2347 3091 2351 3095
rect 2459 3091 2463 3095
rect 2707 3091 2711 3095
rect 3239 3091 3243 3095
rect 3283 3091 3287 3095
rect 643 3083 647 3087
rect 723 3083 727 3087
rect 811 3083 815 3087
rect 927 3083 931 3087
rect 987 3083 991 3087
rect 1075 3083 1079 3087
rect 1163 3083 1167 3087
rect 1251 3083 1255 3087
rect 1339 3083 1343 3087
rect 1391 3083 1395 3087
rect 1903 3082 1907 3086
rect 2015 3082 2019 3086
rect 2191 3082 2195 3086
rect 2407 3082 2411 3086
rect 2655 3082 2659 3086
rect 2935 3082 2939 3086
rect 3231 3082 3235 3086
rect 3511 3082 3515 3086
rect 111 3075 115 3079
rect 583 3072 587 3076
rect 663 3072 667 3076
rect 751 3072 755 3076
rect 839 3072 843 3076
rect 927 3072 931 3076
rect 1015 3072 1019 3076
rect 1103 3072 1107 3076
rect 1191 3072 1195 3076
rect 1279 3072 1283 3076
rect 1367 3072 1371 3076
rect 1831 3075 1835 3079
rect 1871 3064 1875 3068
rect 3591 3064 3595 3068
rect 1955 3055 1959 3059
rect 2039 3055 2043 3059
rect 2199 3055 2203 3059
rect 2459 3055 2463 3059
rect 2707 3055 2711 3059
rect 2943 3055 2947 3059
rect 3283 3055 3287 3059
rect 1871 3047 1875 3051
rect 1895 3044 1899 3048
rect 2007 3044 2011 3048
rect 2183 3044 2187 3048
rect 2399 3044 2403 3048
rect 2647 3044 2651 3048
rect 2927 3044 2931 3048
rect 3223 3044 3227 3048
rect 3503 3044 3507 3048
rect 3591 3047 3595 3051
rect 111 3021 115 3025
rect 543 3024 547 3028
rect 623 3024 627 3028
rect 711 3024 715 3028
rect 807 3024 811 3028
rect 903 3024 907 3028
rect 999 3024 1003 3028
rect 1087 3024 1091 3028
rect 1183 3024 1187 3028
rect 1279 3024 1283 3028
rect 1375 3024 1379 3028
rect 1471 3024 1475 3028
rect 3519 3027 3520 3031
rect 3520 3027 3523 3031
rect 1831 3021 1835 3025
rect 611 3015 615 3019
rect 695 3015 699 3019
rect 111 3004 115 3008
rect 603 3007 607 3011
rect 779 3015 783 3019
rect 875 3015 879 3019
rect 971 3015 975 3019
rect 1067 3015 1071 3019
rect 1155 3015 1159 3019
rect 1255 3015 1259 3019
rect 1347 3015 1351 3019
rect 1443 3015 1447 3019
rect 1831 3004 1835 3008
rect 551 2986 555 2990
rect 631 2986 635 2990
rect 719 2986 723 2990
rect 815 2986 819 2990
rect 911 2986 915 2990
rect 1007 2986 1011 2990
rect 1095 2986 1099 2990
rect 1191 2986 1195 2990
rect 1287 2986 1291 2990
rect 1383 2986 1387 2990
rect 1479 2986 1483 2990
rect 1871 2989 1875 2993
rect 1895 2992 1899 2996
rect 2047 2992 2051 2996
rect 2223 2992 2227 2996
rect 2391 2992 2395 2996
rect 2543 2992 2547 2996
rect 2687 2992 2691 2996
rect 2815 2992 2819 2996
rect 2927 2992 2931 2996
rect 3039 2992 3043 2996
rect 3143 2992 3147 2996
rect 3239 2992 3243 2996
rect 3335 2992 3339 2996
rect 3423 2992 3427 2996
rect 3503 2992 3507 2996
rect 3591 2989 3595 2993
rect 603 2975 607 2979
rect 611 2975 615 2979
rect 779 2975 783 2979
rect 875 2975 879 2979
rect 971 2975 975 2979
rect 987 2975 991 2979
rect 1155 2975 1159 2979
rect 1255 2975 1259 2979
rect 1347 2975 1351 2979
rect 1443 2975 1447 2979
rect 1599 2975 1603 2979
rect 1895 2979 1899 2983
rect 1963 2983 1967 2987
rect 2347 2983 2351 2987
rect 2355 2983 2359 2987
rect 2611 2983 2615 2987
rect 2759 2983 2763 2987
rect 2911 2983 2915 2987
rect 2919 2983 2923 2987
rect 3107 2983 3111 2987
rect 3211 2983 3215 2987
rect 3403 2983 3407 2987
rect 3423 2979 3427 2983
rect 3491 2983 3495 2987
rect 1871 2972 1875 2976
rect 3591 2972 3595 2976
rect 531 2963 535 2967
rect 655 2963 659 2967
rect 695 2963 699 2967
rect 739 2963 743 2967
rect 859 2963 863 2967
rect 1103 2963 1107 2967
rect 1139 2963 1143 2967
rect 1299 2963 1303 2967
rect 1467 2963 1471 2967
rect 1799 2963 1803 2967
rect 3395 2963 3399 2967
rect 3491 2963 3495 2967
rect 471 2954 475 2958
rect 575 2954 579 2958
rect 687 2954 691 2958
rect 807 2954 811 2958
rect 943 2954 947 2958
rect 1087 2954 1091 2958
rect 1247 2954 1251 2958
rect 1415 2954 1419 2958
rect 1591 2954 1595 2958
rect 1751 2954 1755 2958
rect 1903 2954 1907 2958
rect 2055 2954 2059 2958
rect 2231 2954 2235 2958
rect 2399 2954 2403 2958
rect 2551 2954 2555 2958
rect 2695 2954 2699 2958
rect 2823 2954 2827 2958
rect 2935 2954 2939 2958
rect 3047 2954 3051 2958
rect 3151 2954 3155 2958
rect 3247 2954 3251 2958
rect 3343 2954 3347 2958
rect 3431 2954 3435 2958
rect 3511 2954 3515 2958
rect 1963 2943 1967 2947
rect 2039 2943 2043 2947
rect 2355 2943 2359 2947
rect 2495 2943 2499 2947
rect 2567 2943 2571 2947
rect 2611 2943 2615 2947
rect 2759 2943 2763 2947
rect 3107 2943 3111 2947
rect 3211 2943 3215 2947
rect 111 2936 115 2940
rect 1831 2936 1835 2940
rect 3395 2943 3399 2947
rect 3403 2943 3407 2947
rect 3519 2943 3523 2947
rect 523 2927 527 2931
rect 531 2927 535 2931
rect 739 2927 743 2931
rect 859 2927 863 2931
rect 951 2927 955 2931
rect 1139 2927 1143 2931
rect 1299 2927 1303 2931
rect 1467 2927 1471 2931
rect 1599 2927 1603 2931
rect 1895 2931 1896 2935
rect 1896 2931 1899 2935
rect 2095 2931 2099 2935
rect 2139 2931 2143 2935
rect 2347 2931 2351 2935
rect 2715 2931 2719 2935
rect 2723 2931 2727 2935
rect 2911 2931 2915 2935
rect 3099 2931 3103 2935
rect 3203 2931 3207 2935
rect 3363 2935 3367 2939
rect 3423 2931 3427 2935
rect 111 2919 115 2923
rect 463 2916 467 2920
rect 567 2916 571 2920
rect 679 2916 683 2920
rect 799 2916 803 2920
rect 935 2916 939 2920
rect 1079 2916 1083 2920
rect 1239 2916 1243 2920
rect 1407 2916 1411 2920
rect 1583 2916 1587 2920
rect 1743 2916 1747 2920
rect 1831 2919 1835 2923
rect 1903 2922 1907 2926
rect 2087 2922 2091 2926
rect 2295 2922 2299 2926
rect 2487 2922 2491 2926
rect 2671 2922 2675 2926
rect 2839 2922 2843 2926
rect 2999 2922 3003 2926
rect 3151 2922 3155 2926
rect 3303 2922 3307 2926
rect 3455 2922 3459 2926
rect 1871 2904 1875 2908
rect 3591 2904 3595 2908
rect 1759 2899 1760 2903
rect 1760 2899 1763 2903
rect 1799 2895 1803 2899
rect 2139 2895 2143 2899
rect 2347 2895 2351 2899
rect 2495 2895 2499 2899
rect 2723 2895 2727 2899
rect 2879 2895 2883 2899
rect 3099 2895 3103 2899
rect 3203 2895 3207 2899
rect 3311 2895 3315 2899
rect 3363 2895 3367 2899
rect 1871 2887 1875 2891
rect 1895 2884 1899 2888
rect 2079 2884 2083 2888
rect 2287 2884 2291 2888
rect 2479 2884 2483 2888
rect 2663 2884 2667 2888
rect 2831 2884 2835 2888
rect 2991 2884 2995 2888
rect 3143 2884 3147 2888
rect 3295 2884 3299 2888
rect 3447 2884 3451 2888
rect 3591 2887 3595 2891
rect 111 2869 115 2873
rect 311 2872 315 2876
rect 431 2872 435 2876
rect 551 2872 555 2876
rect 679 2872 683 2876
rect 815 2872 819 2876
rect 951 2872 955 2876
rect 1087 2872 1091 2876
rect 1223 2872 1227 2876
rect 1359 2872 1363 2876
rect 1495 2872 1499 2876
rect 1631 2872 1635 2876
rect 1743 2872 1747 2876
rect 1831 2869 1835 2873
rect 379 2863 383 2867
rect 431 2859 435 2863
rect 755 2863 759 2867
rect 763 2863 767 2867
rect 1027 2863 1031 2867
rect 1163 2863 1167 2867
rect 1299 2863 1303 2867
rect 1307 2863 1311 2867
rect 1563 2863 1567 2867
rect 1699 2863 1703 2867
rect 111 2852 115 2856
rect 1555 2855 1559 2859
rect 1831 2852 1835 2856
rect 319 2834 323 2838
rect 439 2834 443 2838
rect 559 2834 563 2838
rect 687 2834 691 2838
rect 823 2834 827 2838
rect 959 2834 963 2838
rect 1095 2834 1099 2838
rect 1231 2834 1235 2838
rect 1367 2834 1371 2838
rect 1503 2834 1507 2838
rect 1639 2834 1643 2838
rect 1751 2834 1755 2838
rect 1871 2829 1875 2833
rect 2135 2832 2139 2836
rect 2263 2832 2267 2836
rect 2391 2832 2395 2836
rect 2519 2832 2523 2836
rect 2647 2832 2651 2836
rect 2767 2832 2771 2836
rect 2887 2832 2891 2836
rect 3007 2832 3011 2836
rect 3135 2832 3139 2836
rect 3591 2829 3595 2833
rect 327 2823 331 2827
rect 379 2823 383 2827
rect 523 2823 527 2827
rect 755 2823 759 2827
rect 967 2823 971 2827
rect 1027 2823 1031 2827
rect 1163 2823 1167 2827
rect 1299 2823 1303 2827
rect 1563 2823 1567 2827
rect 1699 2823 1703 2827
rect 1759 2823 1763 2827
rect 2095 2823 2099 2827
rect 2203 2823 2207 2827
rect 2715 2823 2719 2827
rect 2955 2823 2959 2827
rect 3079 2823 3083 2827
rect 3087 2823 3091 2827
rect 211 2811 215 2815
rect 219 2811 223 2815
rect 431 2811 435 2815
rect 499 2811 503 2815
rect 659 2811 663 2815
rect 1019 2811 1023 2815
rect 1203 2811 1207 2815
rect 1267 2811 1271 2815
rect 1555 2811 1559 2815
rect 1587 2811 1591 2815
rect 1871 2812 1875 2816
rect 2827 2815 2831 2819
rect 3591 2812 3595 2816
rect 167 2802 171 2806
rect 303 2802 307 2806
rect 447 2802 451 2806
rect 607 2802 611 2806
rect 783 2802 787 2806
rect 959 2802 963 2806
rect 1143 2802 1147 2806
rect 1335 2802 1339 2806
rect 1535 2802 1539 2806
rect 1735 2802 1739 2806
rect 2143 2794 2147 2798
rect 2271 2794 2275 2798
rect 2399 2794 2403 2798
rect 2527 2794 2531 2798
rect 2655 2794 2659 2798
rect 2775 2794 2779 2798
rect 2895 2794 2899 2798
rect 3015 2794 3019 2798
rect 3143 2794 3147 2798
rect 111 2784 115 2788
rect 1831 2784 1835 2788
rect 2203 2783 2207 2787
rect 2559 2783 2563 2787
rect 2663 2783 2667 2787
rect 2715 2783 2719 2787
rect 2879 2783 2883 2787
rect 2955 2783 2959 2787
rect 3079 2783 3083 2787
rect 219 2775 223 2779
rect 355 2775 359 2779
rect 499 2775 503 2779
rect 659 2775 663 2779
rect 967 2775 971 2779
rect 1019 2775 1023 2779
rect 1203 2775 1207 2779
rect 1587 2775 1591 2779
rect 111 2767 115 2771
rect 159 2764 163 2768
rect 295 2764 299 2768
rect 439 2764 443 2768
rect 599 2764 603 2768
rect 775 2764 779 2768
rect 951 2764 955 2768
rect 1135 2764 1139 2768
rect 1327 2764 1331 2768
rect 1527 2764 1531 2768
rect 1727 2764 1731 2768
rect 1831 2767 1835 2771
rect 2283 2763 2287 2767
rect 2363 2763 2367 2767
rect 2443 2763 2447 2767
rect 2543 2763 2544 2767
rect 2544 2763 2547 2767
rect 2647 2763 2651 2767
rect 2691 2763 2695 2767
rect 2827 2763 2831 2767
rect 2867 2763 2871 2767
rect 2955 2763 2959 2767
rect 2231 2754 2235 2758
rect 2311 2754 2315 2758
rect 2391 2754 2395 2758
rect 2471 2754 2475 2758
rect 2551 2754 2555 2758
rect 2639 2754 2643 2758
rect 2727 2754 2731 2758
rect 2815 2754 2819 2758
rect 2903 2754 2907 2758
rect 2991 2754 2995 2758
rect 211 2747 215 2751
rect 1703 2747 1707 2751
rect 1871 2736 1875 2740
rect 3591 2736 3595 2740
rect 2283 2727 2287 2731
rect 2363 2727 2367 2731
rect 2443 2727 2447 2731
rect 2543 2727 2547 2731
rect 2559 2727 2563 2731
rect 2691 2727 2695 2731
rect 2779 2727 2783 2731
rect 2867 2727 2871 2731
rect 2955 2727 2959 2731
rect 2999 2727 3003 2731
rect 111 2713 115 2717
rect 135 2716 139 2720
rect 247 2716 251 2720
rect 391 2716 395 2720
rect 551 2716 555 2720
rect 711 2716 715 2720
rect 879 2716 883 2720
rect 1039 2716 1043 2720
rect 1199 2716 1203 2720
rect 1359 2716 1363 2720
rect 1519 2716 1523 2720
rect 1687 2716 1691 2720
rect 1871 2719 1875 2723
rect 1831 2713 1835 2717
rect 2223 2716 2227 2720
rect 2303 2716 2307 2720
rect 2383 2716 2387 2720
rect 2463 2716 2467 2720
rect 2543 2716 2547 2720
rect 2631 2716 2635 2720
rect 2719 2716 2723 2720
rect 2807 2716 2811 2720
rect 2895 2716 2899 2720
rect 2983 2716 2987 2720
rect 3591 2719 3595 2723
rect 135 2703 139 2707
rect 203 2707 207 2711
rect 479 2707 483 2711
rect 111 2696 115 2700
rect 651 2699 655 2703
rect 963 2707 967 2711
rect 1111 2707 1115 2711
rect 1267 2707 1271 2711
rect 1359 2703 1363 2707
rect 1427 2707 1431 2711
rect 1587 2707 1591 2711
rect 1831 2696 1835 2700
rect 143 2678 147 2682
rect 255 2678 259 2682
rect 399 2678 403 2682
rect 559 2678 563 2682
rect 719 2678 723 2682
rect 887 2678 891 2682
rect 1047 2678 1051 2682
rect 1207 2678 1211 2682
rect 1367 2678 1371 2682
rect 1527 2678 1531 2682
rect 1695 2678 1699 2682
rect 203 2667 207 2671
rect 263 2667 267 2671
rect 355 2667 359 2671
rect 479 2667 483 2671
rect 895 2667 899 2671
rect 963 2667 967 2671
rect 1111 2667 1115 2671
rect 1427 2667 1431 2671
rect 1587 2667 1591 2671
rect 1703 2667 1707 2671
rect 1871 2669 1875 2673
rect 2239 2672 2243 2676
rect 2319 2672 2323 2676
rect 2399 2672 2403 2676
rect 2479 2672 2483 2676
rect 2559 2672 2563 2676
rect 2639 2672 2643 2676
rect 2719 2672 2723 2676
rect 2799 2672 2803 2676
rect 2879 2672 2883 2676
rect 2959 2672 2963 2676
rect 3591 2669 3595 2673
rect 2387 2663 2391 2667
rect 2467 2663 2471 2667
rect 2547 2663 2551 2667
rect 135 2655 136 2659
rect 136 2655 139 2659
rect 195 2655 199 2659
rect 307 2655 311 2659
rect 451 2655 455 2659
rect 603 2655 607 2659
rect 939 2655 943 2659
rect 1135 2655 1139 2659
rect 1187 2655 1191 2659
rect 1359 2655 1363 2659
rect 1443 2655 1447 2659
rect 2639 2659 2643 2663
rect 2707 2663 2711 2667
rect 2867 2663 2871 2667
rect 2947 2663 2951 2667
rect 1871 2652 1875 2656
rect 2787 2655 2791 2659
rect 3591 2652 3595 2656
rect 143 2646 147 2650
rect 255 2646 259 2650
rect 399 2646 403 2650
rect 551 2646 555 2650
rect 711 2646 715 2650
rect 879 2646 883 2650
rect 1047 2646 1051 2650
rect 1215 2646 1219 2650
rect 1391 2646 1395 2650
rect 1567 2646 1571 2650
rect 2247 2634 2251 2638
rect 2327 2634 2331 2638
rect 2407 2634 2411 2638
rect 2487 2634 2491 2638
rect 2567 2634 2571 2638
rect 2647 2634 2651 2638
rect 2727 2634 2731 2638
rect 111 2628 115 2632
rect 1831 2628 1835 2632
rect 195 2619 199 2623
rect 307 2619 311 2623
rect 451 2619 455 2623
rect 603 2619 607 2623
rect 895 2619 899 2623
rect 939 2619 943 2623
rect 1135 2619 1139 2623
rect 1443 2619 1447 2623
rect 2387 2623 2391 2627
rect 2467 2623 2471 2627
rect 2547 2623 2551 2627
rect 2599 2623 2603 2627
rect 2707 2623 2711 2627
rect 2787 2631 2791 2635
rect 2807 2634 2811 2638
rect 2887 2634 2891 2638
rect 2967 2634 2971 2638
rect 2779 2623 2783 2627
rect 2867 2623 2871 2627
rect 2947 2623 2951 2627
rect 111 2611 115 2615
rect 135 2608 139 2612
rect 247 2608 251 2612
rect 391 2608 395 2612
rect 543 2608 547 2612
rect 703 2608 707 2612
rect 871 2608 875 2612
rect 1039 2608 1043 2612
rect 1207 2608 1211 2612
rect 1383 2608 1387 2612
rect 1559 2608 1563 2612
rect 1831 2611 1835 2615
rect 2475 2611 2479 2615
rect 2255 2603 2259 2607
rect 2335 2603 2339 2607
rect 2415 2603 2419 2607
rect 2495 2603 2499 2607
rect 2583 2603 2584 2607
rect 2584 2603 2587 2607
rect 2639 2603 2643 2607
rect 2735 2603 2739 2607
rect 2815 2603 2819 2607
rect 2895 2603 2899 2607
rect 2975 2603 2979 2607
rect 643 2591 647 2595
rect 1543 2591 1547 2595
rect 2191 2594 2195 2598
rect 2271 2594 2275 2598
rect 2351 2594 2355 2598
rect 2431 2594 2435 2598
rect 2511 2594 2515 2598
rect 2591 2594 2595 2598
rect 2671 2594 2675 2598
rect 2751 2594 2755 2598
rect 2831 2594 2835 2598
rect 2911 2594 2915 2598
rect 2991 2594 2995 2598
rect 1871 2576 1875 2580
rect 3591 2576 3595 2580
rect 2255 2567 2259 2571
rect 2335 2567 2339 2571
rect 2415 2567 2419 2571
rect 2495 2567 2499 2571
rect 2583 2567 2587 2571
rect 2599 2567 2603 2571
rect 2735 2567 2739 2571
rect 2815 2567 2819 2571
rect 2895 2567 2899 2571
rect 2975 2567 2979 2571
rect 111 2557 115 2561
rect 159 2560 163 2564
rect 279 2560 283 2564
rect 415 2560 419 2564
rect 559 2560 563 2564
rect 703 2560 707 2564
rect 847 2560 851 2564
rect 983 2560 987 2564
rect 1119 2560 1123 2564
rect 1255 2560 1259 2564
rect 1391 2560 1395 2564
rect 1527 2560 1531 2564
rect 1831 2557 1835 2561
rect 1871 2559 1875 2563
rect 2183 2556 2187 2560
rect 227 2551 231 2555
rect 347 2551 351 2555
rect 483 2551 487 2555
rect 635 2551 639 2555
rect 667 2551 671 2555
rect 915 2551 919 2555
rect 1051 2551 1055 2555
rect 1187 2551 1191 2555
rect 1331 2551 1335 2555
rect 2263 2556 2267 2560
rect 2343 2556 2347 2560
rect 2423 2556 2427 2560
rect 2503 2556 2507 2560
rect 2583 2556 2587 2560
rect 2663 2556 2667 2560
rect 2743 2556 2747 2560
rect 2823 2556 2827 2560
rect 2903 2556 2907 2560
rect 2983 2556 2987 2560
rect 3591 2559 3595 2563
rect 1479 2551 1483 2555
rect 111 2540 115 2544
rect 1315 2543 1319 2547
rect 1831 2540 1835 2544
rect 2607 2539 2611 2543
rect 167 2522 171 2526
rect 287 2522 291 2526
rect 423 2522 427 2526
rect 567 2522 571 2526
rect 711 2522 715 2526
rect 855 2522 859 2526
rect 991 2522 995 2526
rect 1127 2522 1131 2526
rect 1263 2522 1267 2526
rect 1399 2522 1403 2526
rect 1535 2522 1539 2526
rect 175 2511 179 2515
rect 227 2511 231 2515
rect 347 2511 351 2515
rect 483 2511 487 2515
rect 635 2511 639 2515
rect 887 2511 891 2515
rect 915 2511 919 2515
rect 1051 2511 1055 2515
rect 1331 2511 1335 2515
rect 1479 2511 1483 2515
rect 1543 2511 1547 2515
rect 1871 2501 1875 2505
rect 2119 2504 2123 2508
rect 2207 2504 2211 2508
rect 2303 2504 2307 2508
rect 2399 2504 2403 2508
rect 2495 2504 2499 2508
rect 2591 2504 2595 2508
rect 2687 2504 2691 2508
rect 2783 2504 2787 2508
rect 2879 2504 2883 2508
rect 2975 2504 2979 2508
rect 3079 2504 3083 2508
rect 3591 2501 3595 2505
rect 355 2495 359 2499
rect 387 2495 391 2499
rect 467 2495 471 2499
rect 555 2495 559 2499
rect 651 2495 655 2499
rect 755 2495 759 2499
rect 999 2495 1003 2499
rect 1271 2495 1275 2499
rect 1315 2495 1319 2499
rect 1379 2495 1383 2499
rect 2187 2495 2191 2499
rect 2275 2495 2279 2499
rect 2371 2495 2375 2499
rect 2467 2495 2471 2499
rect 2475 2495 2479 2499
rect 2659 2495 2663 2499
rect 2755 2495 2759 2499
rect 2851 2495 2855 2499
rect 2947 2495 2951 2499
rect 3043 2495 3047 2499
rect 3051 2495 3055 2499
rect 335 2486 339 2490
rect 415 2486 419 2490
rect 503 2486 507 2490
rect 599 2486 603 2490
rect 703 2486 707 2490
rect 815 2486 819 2490
rect 935 2486 939 2490
rect 1063 2486 1067 2490
rect 1191 2486 1195 2490
rect 1327 2486 1331 2490
rect 1471 2486 1475 2490
rect 1871 2484 1875 2488
rect 3591 2484 3595 2488
rect 111 2468 115 2472
rect 1831 2468 1835 2472
rect 2127 2466 2131 2470
rect 2215 2466 2219 2470
rect 2311 2466 2315 2470
rect 2407 2466 2411 2470
rect 2503 2466 2507 2470
rect 2599 2466 2603 2470
rect 2695 2466 2699 2470
rect 2791 2466 2795 2470
rect 2887 2466 2891 2470
rect 2983 2466 2987 2470
rect 3087 2466 3091 2470
rect 387 2459 391 2463
rect 467 2459 471 2463
rect 555 2459 559 2463
rect 651 2459 655 2463
rect 755 2459 759 2463
rect 887 2459 891 2463
rect 999 2459 1003 2463
rect 1379 2459 1383 2463
rect 1519 2459 1523 2463
rect 111 2451 115 2455
rect 327 2448 331 2452
rect 407 2448 411 2452
rect 495 2448 499 2452
rect 591 2448 595 2452
rect 695 2448 699 2452
rect 807 2448 811 2452
rect 927 2448 931 2452
rect 1055 2448 1059 2452
rect 1183 2448 1187 2452
rect 1319 2448 1323 2452
rect 1463 2448 1467 2452
rect 1831 2451 1835 2455
rect 2179 2455 2183 2459
rect 2187 2455 2191 2459
rect 2275 2455 2279 2459
rect 2371 2455 2375 2459
rect 2467 2455 2471 2459
rect 2607 2455 2611 2459
rect 2659 2455 2663 2459
rect 2755 2455 2759 2459
rect 2851 2455 2855 2459
rect 2947 2455 2951 2459
rect 3043 2455 3047 2459
rect 1947 2439 1951 2443
rect 1955 2439 1959 2443
rect 2043 2439 2047 2443
rect 2163 2439 2167 2443
rect 2299 2439 2303 2443
rect 2443 2439 2447 2443
rect 2703 2439 2707 2443
rect 2723 2439 2727 2443
rect 2859 2439 2863 2443
rect 2995 2439 2999 2443
rect 3131 2439 3135 2443
rect 799 2431 803 2435
rect 1903 2430 1907 2434
rect 1991 2430 1995 2434
rect 2111 2430 2115 2434
rect 2247 2430 2251 2434
rect 2391 2430 2395 2434
rect 2535 2430 2539 2434
rect 2671 2430 2675 2434
rect 2807 2430 2811 2434
rect 2943 2430 2947 2434
rect 3079 2430 3083 2434
rect 3215 2430 3219 2434
rect 1871 2412 1875 2416
rect 3591 2412 3595 2416
rect 1955 2403 1959 2407
rect 2043 2403 2047 2407
rect 2163 2403 2167 2407
rect 2299 2403 2303 2407
rect 2443 2403 2447 2407
rect 2543 2403 2547 2407
rect 2723 2403 2727 2407
rect 2859 2403 2863 2407
rect 2995 2403 2999 2407
rect 3131 2403 3135 2407
rect 111 2393 115 2397
rect 383 2396 387 2400
rect 463 2396 467 2400
rect 543 2396 547 2400
rect 623 2396 627 2400
rect 703 2396 707 2400
rect 783 2396 787 2400
rect 863 2396 867 2400
rect 943 2396 947 2400
rect 1023 2396 1027 2400
rect 1103 2396 1107 2400
rect 1183 2396 1187 2400
rect 1263 2396 1267 2400
rect 1351 2396 1355 2400
rect 1439 2396 1443 2400
rect 1527 2396 1531 2400
rect 1831 2393 1835 2397
rect 1871 2395 1875 2399
rect 1895 2392 1899 2396
rect 451 2387 455 2391
rect 531 2387 535 2391
rect 611 2387 615 2391
rect 691 2387 695 2391
rect 771 2387 775 2391
rect 863 2383 867 2387
rect 931 2387 935 2391
rect 1011 2387 1015 2391
rect 1091 2387 1095 2391
rect 1171 2387 1175 2391
rect 1251 2387 1255 2391
rect 1271 2383 1275 2387
rect 1419 2387 1423 2391
rect 1427 2387 1431 2391
rect 1983 2392 1987 2396
rect 2103 2392 2107 2396
rect 2239 2392 2243 2396
rect 2383 2392 2387 2396
rect 2527 2392 2531 2396
rect 2663 2392 2667 2396
rect 2799 2392 2803 2396
rect 2935 2392 2939 2396
rect 3071 2392 3075 2396
rect 3207 2392 3211 2396
rect 3591 2395 3595 2399
rect 1507 2387 1511 2391
rect 111 2376 115 2380
rect 1831 2376 1835 2380
rect 3139 2375 3143 2379
rect 391 2358 395 2362
rect 471 2358 475 2362
rect 551 2358 555 2362
rect 631 2358 635 2362
rect 711 2358 715 2362
rect 791 2358 795 2362
rect 871 2358 875 2362
rect 951 2358 955 2362
rect 1031 2358 1035 2362
rect 1111 2358 1115 2362
rect 1191 2358 1195 2362
rect 1271 2358 1275 2362
rect 1359 2358 1363 2362
rect 1447 2358 1451 2362
rect 1535 2358 1539 2362
rect 451 2347 455 2351
rect 531 2347 535 2351
rect 611 2347 615 2351
rect 691 2347 695 2351
rect 771 2347 775 2351
rect 863 2347 864 2351
rect 864 2347 867 2351
rect 931 2347 935 2351
rect 1011 2347 1015 2351
rect 1091 2347 1095 2351
rect 1171 2347 1175 2351
rect 1251 2347 1255 2351
rect 1427 2347 1431 2351
rect 1507 2347 1511 2351
rect 1519 2347 1523 2351
rect 799 2339 803 2343
rect 1419 2335 1423 2339
rect 1459 2335 1463 2339
rect 1559 2335 1560 2339
rect 1560 2335 1563 2339
rect 1619 2335 1623 2339
rect 1871 2337 1875 2341
rect 1895 2340 1899 2344
rect 2015 2340 2019 2344
rect 2175 2340 2179 2344
rect 2343 2340 2347 2344
rect 2511 2340 2515 2344
rect 2671 2340 2675 2344
rect 2823 2340 2827 2344
rect 2959 2340 2963 2344
rect 3079 2340 3083 2344
rect 3191 2340 3195 2344
rect 3303 2340 3307 2344
rect 3415 2340 3419 2344
rect 3503 2340 3507 2344
rect 3591 2337 3595 2341
rect 1963 2331 1967 2335
rect 1407 2326 1411 2330
rect 1487 2326 1491 2330
rect 1567 2326 1571 2330
rect 2099 2331 2103 2335
rect 2243 2331 2247 2335
rect 2435 2331 2439 2335
rect 2459 2331 2463 2335
rect 2755 2331 2759 2335
rect 2891 2331 2895 2335
rect 3031 2331 3035 2335
rect 3147 2331 3151 2335
rect 3263 2331 3267 2335
rect 3371 2331 3375 2335
rect 3483 2331 3487 2335
rect 1647 2326 1651 2330
rect 1871 2320 1875 2324
rect 3591 2320 3595 2324
rect 111 2308 115 2312
rect 1831 2308 1835 2312
rect 1459 2299 1463 2303
rect 1559 2299 1563 2303
rect 1619 2299 1623 2303
rect 1903 2302 1907 2306
rect 2023 2302 2027 2306
rect 2183 2302 2187 2306
rect 2351 2302 2355 2306
rect 2519 2302 2523 2306
rect 2679 2302 2683 2306
rect 2831 2302 2835 2306
rect 2967 2302 2971 2306
rect 3087 2302 3091 2306
rect 3199 2302 3203 2306
rect 3311 2302 3315 2306
rect 3423 2302 3427 2306
rect 3511 2302 3515 2306
rect 111 2291 115 2295
rect 1399 2288 1403 2292
rect 1479 2288 1483 2292
rect 1559 2288 1563 2292
rect 1639 2288 1643 2292
rect 1831 2291 1835 2295
rect 1911 2291 1915 2295
rect 1963 2291 1967 2295
rect 2099 2291 2103 2295
rect 2243 2291 2247 2295
rect 2435 2291 2439 2295
rect 2687 2291 2691 2295
rect 2755 2291 2759 2295
rect 2891 2291 2895 2295
rect 3031 2291 3035 2295
rect 3147 2291 3151 2295
rect 3263 2291 3267 2295
rect 3371 2291 3375 2295
rect 3483 2291 3487 2295
rect 1963 2279 1967 2283
rect 2375 2279 2379 2283
rect 2479 2279 2483 2283
rect 2627 2279 2631 2283
rect 1579 2271 1583 2275
rect 1903 2270 1907 2274
rect 2031 2270 2035 2274
rect 2183 2270 2187 2274
rect 2367 2270 2371 2274
rect 2575 2270 2579 2274
rect 2791 2270 2795 2274
rect 3023 2270 3027 2274
rect 3075 2279 3079 2283
rect 3343 2283 3347 2287
rect 3255 2270 3259 2274
rect 3495 2270 3499 2274
rect 1871 2252 1875 2256
rect 3591 2252 3595 2256
rect 1911 2243 1915 2247
rect 1963 2243 1967 2247
rect 2627 2243 2631 2247
rect 3075 2243 3079 2247
rect 3335 2243 3339 2247
rect 3343 2243 3347 2247
rect 111 2233 115 2237
rect 135 2236 139 2240
rect 215 2236 219 2240
rect 295 2236 299 2240
rect 383 2236 387 2240
rect 519 2236 523 2240
rect 671 2236 675 2240
rect 831 2236 835 2240
rect 999 2236 1003 2240
rect 1159 2236 1163 2240
rect 1311 2236 1315 2240
rect 1455 2236 1459 2240
rect 1607 2236 1611 2240
rect 1743 2236 1747 2240
rect 1831 2233 1835 2237
rect 1871 2235 1875 2239
rect 1895 2232 1899 2236
rect 203 2227 207 2231
rect 283 2227 287 2231
rect 363 2227 367 2231
rect 459 2227 463 2231
rect 587 2227 591 2231
rect 755 2227 759 2231
rect 923 2227 927 2231
rect 999 2223 1003 2227
rect 1235 2227 1239 2231
rect 1379 2227 1383 2231
rect 1531 2227 1535 2231
rect 1683 2227 1687 2231
rect 2023 2232 2027 2236
rect 2175 2232 2179 2236
rect 2359 2232 2363 2236
rect 2567 2232 2571 2236
rect 2783 2232 2787 2236
rect 3015 2232 3019 2236
rect 3247 2232 3251 2236
rect 3487 2232 3491 2236
rect 3591 2235 3595 2239
rect 1691 2227 1695 2231
rect 111 2216 115 2220
rect 1831 2216 1835 2220
rect 2375 2215 2379 2219
rect 143 2198 147 2202
rect 223 2198 227 2202
rect 303 2198 307 2202
rect 391 2198 395 2202
rect 527 2198 531 2202
rect 679 2198 683 2202
rect 839 2198 843 2202
rect 1007 2198 1011 2202
rect 1167 2198 1171 2202
rect 1319 2198 1323 2202
rect 1463 2198 1467 2202
rect 1615 2198 1619 2202
rect 1751 2198 1755 2202
rect 203 2187 207 2191
rect 283 2187 287 2191
rect 363 2187 367 2191
rect 459 2187 463 2191
rect 587 2187 591 2191
rect 755 2187 759 2191
rect 923 2187 927 2191
rect 1175 2187 1179 2191
rect 1235 2187 1239 2191
rect 1379 2187 1383 2191
rect 1531 2187 1535 2191
rect 1683 2187 1687 2191
rect 199 2171 203 2175
rect 283 2171 287 2175
rect 363 2171 367 2175
rect 647 2171 651 2175
rect 691 2171 695 2175
rect 999 2171 1003 2175
rect 1207 2171 1211 2175
rect 1251 2171 1255 2175
rect 1443 2171 1447 2175
rect 1635 2171 1639 2175
rect 191 2162 195 2166
rect 311 2162 315 2166
rect 463 2162 467 2166
rect 639 2162 643 2166
rect 823 2162 827 2166
rect 1015 2162 1019 2166
rect 1199 2162 1203 2166
rect 1391 2162 1395 2166
rect 1583 2162 1587 2166
rect 1751 2162 1755 2166
rect 1871 2165 1875 2169
rect 2199 2168 2203 2172
rect 2295 2168 2299 2172
rect 2399 2168 2403 2172
rect 2519 2168 2523 2172
rect 2639 2168 2643 2172
rect 2759 2168 2763 2172
rect 2879 2168 2883 2172
rect 2991 2168 2995 2172
rect 3095 2168 3099 2172
rect 3199 2168 3203 2172
rect 3303 2168 3307 2172
rect 3407 2168 3411 2172
rect 3503 2168 3507 2172
rect 3591 2165 3595 2169
rect 2267 2159 2271 2163
rect 2363 2159 2367 2163
rect 2479 2159 2483 2163
rect 2487 2159 2491 2163
rect 2587 2159 2591 2163
rect 2707 2159 2711 2163
rect 2947 2159 2951 2163
rect 3059 2159 3063 2163
rect 3175 2159 3179 2163
rect 3267 2159 3271 2163
rect 3475 2159 3479 2163
rect 3503 2155 3507 2159
rect 111 2144 115 2148
rect 1831 2144 1835 2148
rect 1871 2148 1875 2152
rect 3591 2148 3595 2152
rect 363 2135 367 2139
rect 471 2135 475 2139
rect 691 2135 695 2139
rect 875 2135 879 2139
rect 1023 2135 1027 2139
rect 1251 2135 1255 2139
rect 1443 2135 1447 2139
rect 1635 2135 1639 2139
rect 111 2127 115 2131
rect 183 2124 187 2128
rect 303 2124 307 2128
rect 455 2124 459 2128
rect 631 2124 635 2128
rect 815 2124 819 2128
rect 1007 2124 1011 2128
rect 1191 2124 1195 2128
rect 1383 2124 1387 2128
rect 1575 2124 1579 2128
rect 1743 2124 1747 2128
rect 1831 2127 1835 2131
rect 2207 2130 2211 2134
rect 2303 2130 2307 2134
rect 2407 2130 2411 2134
rect 2527 2130 2531 2134
rect 2647 2130 2651 2134
rect 2767 2130 2771 2134
rect 2887 2130 2891 2134
rect 2999 2130 3003 2134
rect 3103 2130 3107 2134
rect 3207 2130 3211 2134
rect 3311 2130 3315 2134
rect 3415 2130 3419 2134
rect 3511 2130 3515 2134
rect 2215 2119 2219 2123
rect 2267 2119 2271 2123
rect 2363 2119 2367 2123
rect 2587 2119 2591 2123
rect 2707 2119 2711 2123
rect 2759 2119 2760 2123
rect 2760 2119 2763 2123
rect 2947 2119 2951 2123
rect 3059 2119 3063 2123
rect 3175 2119 3179 2123
rect 3267 2119 3271 2123
rect 3319 2119 3323 2123
rect 3335 2119 3339 2123
rect 3475 2119 3479 2123
rect 1759 2107 1760 2111
rect 1760 2107 1763 2111
rect 2455 2103 2459 2107
rect 2227 2095 2231 2099
rect 2323 2095 2327 2099
rect 2427 2095 2431 2099
rect 2539 2095 2543 2099
rect 2659 2095 2663 2099
rect 2899 2095 2903 2099
rect 3019 2095 3023 2099
rect 3423 2103 3427 2107
rect 3243 2095 3247 2099
rect 3431 2095 3435 2099
rect 3503 2095 3504 2099
rect 3504 2095 3507 2099
rect 2175 2086 2179 2090
rect 2271 2086 2275 2090
rect 2375 2086 2379 2090
rect 2487 2086 2491 2090
rect 2607 2086 2611 2090
rect 2727 2086 2731 2090
rect 2847 2086 2851 2090
rect 2967 2086 2971 2090
rect 3079 2086 3083 2090
rect 3191 2086 3195 2090
rect 3303 2086 3307 2090
rect 3415 2086 3419 2090
rect 3511 2086 3515 2090
rect 111 2073 115 2077
rect 215 2076 219 2080
rect 359 2076 363 2080
rect 519 2076 523 2080
rect 703 2076 707 2080
rect 895 2076 899 2080
rect 1103 2076 1107 2080
rect 1311 2076 1315 2080
rect 1527 2076 1531 2080
rect 1743 2076 1747 2080
rect 1831 2073 1835 2077
rect 283 2067 287 2071
rect 291 2067 295 2071
rect 587 2067 591 2071
rect 771 2067 775 2071
rect 1215 2067 1219 2071
rect 111 2056 115 2060
rect 1595 2067 1599 2071
rect 1603 2067 1607 2071
rect 1871 2068 1875 2072
rect 3591 2068 3595 2072
rect 1831 2056 1835 2060
rect 2227 2059 2231 2063
rect 2323 2059 2327 2063
rect 2427 2059 2431 2063
rect 2539 2059 2543 2063
rect 2659 2059 2663 2063
rect 2759 2059 2763 2063
rect 2899 2059 2903 2063
rect 3019 2059 3023 2063
rect 3243 2059 3247 2063
rect 3319 2059 3323 2063
rect 3423 2059 3427 2063
rect 1871 2051 1875 2055
rect 2167 2048 2171 2052
rect 2263 2048 2267 2052
rect 2367 2048 2371 2052
rect 2479 2048 2483 2052
rect 2599 2048 2603 2052
rect 2719 2048 2723 2052
rect 2839 2048 2843 2052
rect 2959 2048 2963 2052
rect 3071 2048 3075 2052
rect 3183 2048 3187 2052
rect 3295 2048 3299 2052
rect 3407 2048 3411 2052
rect 3503 2048 3507 2052
rect 3591 2051 3595 2055
rect 223 2038 227 2042
rect 367 2038 371 2042
rect 527 2038 531 2042
rect 711 2038 715 2042
rect 903 2038 907 2042
rect 1111 2038 1115 2042
rect 1319 2038 1323 2042
rect 1535 2038 1539 2042
rect 1751 2038 1755 2042
rect 291 2027 295 2031
rect 391 2027 395 2031
rect 587 2027 591 2031
rect 771 2027 775 2031
rect 875 2027 879 2031
rect 1075 2027 1079 2031
rect 1215 2027 1219 2031
rect 1603 2027 1607 2031
rect 1759 2027 1763 2031
rect 3031 2031 3035 2035
rect 3519 2031 3520 2035
rect 3520 2031 3523 2035
rect 151 2015 155 2019
rect 195 2015 199 2019
rect 315 2015 319 2019
rect 547 2015 551 2019
rect 659 2015 663 2019
rect 867 2015 871 2019
rect 875 2015 879 2019
rect 979 2015 983 2019
rect 1163 2015 1167 2019
rect 1259 2015 1263 2019
rect 1347 2015 1351 2019
rect 1443 2015 1447 2019
rect 1595 2015 1599 2019
rect 1635 2015 1639 2019
rect 1723 2015 1727 2019
rect 143 2006 147 2010
rect 263 2006 267 2010
rect 383 2006 387 2010
rect 495 2006 499 2010
rect 607 2006 611 2010
rect 719 2006 723 2010
rect 823 2006 827 2010
rect 927 2006 931 2010
rect 1023 2006 1027 2010
rect 1111 2006 1115 2010
rect 1207 2006 1211 2010
rect 1295 2006 1299 2010
rect 1391 2006 1395 2010
rect 1487 2006 1491 2010
rect 1583 2006 1587 2010
rect 1671 2006 1675 2010
rect 1751 2006 1755 2010
rect 1871 1997 1875 2001
rect 2071 2000 2075 2004
rect 2207 2000 2211 2004
rect 2359 2000 2363 2004
rect 2519 2000 2523 2004
rect 2679 2000 2683 2004
rect 2847 2000 2851 2004
rect 3015 2000 3019 2004
rect 3183 2000 3187 2004
rect 3351 2000 3355 2004
rect 3503 2000 3507 2004
rect 3591 1997 3595 2001
rect 111 1988 115 1992
rect 1831 1988 1835 1992
rect 2147 1991 2151 1995
rect 2275 1991 2279 1995
rect 2447 1991 2451 1995
rect 2455 1991 2459 1995
rect 2599 1991 2603 1995
rect 2747 1991 2751 1995
rect 2915 1991 2919 1995
rect 3275 1991 3279 1995
rect 3431 1991 3435 1995
rect 195 1979 199 1983
rect 315 1979 319 1983
rect 391 1979 395 1983
rect 547 1979 551 1983
rect 659 1979 663 1983
rect 771 1979 775 1983
rect 875 1979 879 1983
rect 979 1979 983 1983
rect 1075 1979 1079 1983
rect 1163 1979 1167 1983
rect 1259 1979 1263 1983
rect 1347 1979 1351 1983
rect 1443 1979 1447 1983
rect 1635 1979 1639 1983
rect 1723 1979 1727 1983
rect 1871 1980 1875 1984
rect 3263 1983 3267 1987
rect 3591 1980 3595 1984
rect 111 1971 115 1975
rect 135 1968 139 1972
rect 255 1968 259 1972
rect 375 1968 379 1972
rect 487 1968 491 1972
rect 599 1968 603 1972
rect 711 1968 715 1972
rect 815 1968 819 1972
rect 919 1968 923 1972
rect 1015 1968 1019 1972
rect 1103 1968 1107 1972
rect 1199 1968 1203 1972
rect 1287 1968 1291 1972
rect 1383 1968 1387 1972
rect 1479 1968 1483 1972
rect 1575 1968 1579 1972
rect 1663 1968 1667 1972
rect 1743 1968 1747 1972
rect 1831 1971 1835 1975
rect 2079 1962 2083 1966
rect 2215 1962 2219 1966
rect 2367 1962 2371 1966
rect 2527 1962 2531 1966
rect 2687 1962 2691 1966
rect 2855 1962 2859 1966
rect 3023 1962 3027 1966
rect 3191 1962 3195 1966
rect 3359 1962 3363 1966
rect 3511 1962 3515 1966
rect 1231 1951 1235 1955
rect 1759 1951 1760 1955
rect 1760 1951 1763 1955
rect 2059 1951 2063 1955
rect 2147 1951 2151 1955
rect 2275 1951 2279 1955
rect 2447 1951 2451 1955
rect 2747 1951 2751 1955
rect 2915 1951 2919 1955
rect 3031 1951 3035 1955
rect 3263 1951 3267 1955
rect 3275 1951 3279 1955
rect 3519 1951 3523 1955
rect 1811 1939 1815 1943
rect 2067 1939 2071 1943
rect 2195 1939 2199 1943
rect 2351 1939 2355 1943
rect 2383 1939 2387 1943
rect 2427 1939 2431 1943
rect 2539 1939 2543 1943
rect 2651 1939 2655 1943
rect 2771 1939 2775 1943
rect 1903 1930 1907 1934
rect 2007 1930 2011 1934
rect 2135 1930 2139 1934
rect 2255 1930 2259 1934
rect 2375 1930 2379 1934
rect 2487 1930 2491 1934
rect 2599 1930 2603 1934
rect 2719 1930 2723 1934
rect 2839 1930 2843 1934
rect 111 1913 115 1917
rect 167 1916 171 1920
rect 327 1916 331 1920
rect 487 1916 491 1920
rect 647 1916 651 1920
rect 799 1916 803 1920
rect 943 1916 947 1920
rect 1079 1916 1083 1920
rect 1215 1916 1219 1920
rect 1351 1916 1355 1920
rect 1487 1916 1491 1920
rect 1623 1916 1627 1920
rect 1743 1916 1747 1920
rect 1831 1913 1835 1917
rect 1871 1912 1875 1916
rect 151 1907 155 1911
rect 235 1907 239 1911
rect 555 1907 559 1911
rect 563 1907 567 1911
rect 715 1907 719 1911
rect 867 1907 871 1911
rect 1011 1907 1015 1911
rect 1291 1907 1295 1911
rect 1419 1907 1423 1911
rect 1555 1907 1559 1911
rect 3591 1912 3595 1916
rect 111 1896 115 1900
rect 1343 1899 1347 1903
rect 1811 1907 1815 1911
rect 2059 1903 2063 1907
rect 2067 1903 2071 1907
rect 2195 1903 2199 1907
rect 2427 1903 2431 1907
rect 2539 1903 2543 1907
rect 2651 1903 2655 1907
rect 2771 1903 2775 1907
rect 1831 1896 1835 1900
rect 1871 1895 1875 1899
rect 1895 1892 1899 1896
rect 1999 1892 2003 1896
rect 2127 1892 2131 1896
rect 2247 1892 2251 1896
rect 2367 1892 2371 1896
rect 2479 1892 2483 1896
rect 2591 1892 2595 1896
rect 2711 1892 2715 1896
rect 2831 1892 2835 1896
rect 3591 1895 3595 1899
rect 175 1878 179 1882
rect 335 1878 339 1882
rect 495 1878 499 1882
rect 655 1878 659 1882
rect 807 1878 811 1882
rect 951 1878 955 1882
rect 1087 1878 1091 1882
rect 1223 1878 1227 1882
rect 1359 1878 1363 1882
rect 1495 1878 1499 1882
rect 1631 1878 1635 1882
rect 1751 1878 1755 1882
rect 1911 1875 1912 1879
rect 1912 1875 1915 1879
rect 2535 1875 2539 1879
rect 235 1867 239 1871
rect 327 1867 328 1871
rect 328 1867 331 1871
rect 563 1867 567 1871
rect 715 1867 719 1871
rect 771 1867 775 1871
rect 1011 1867 1015 1871
rect 1079 1867 1080 1871
rect 1080 1867 1083 1871
rect 1231 1867 1235 1871
rect 1291 1867 1295 1871
rect 1419 1867 1423 1871
rect 1555 1867 1559 1871
rect 1759 1867 1763 1871
rect 183 1855 187 1859
rect 211 1855 215 1859
rect 431 1855 435 1859
rect 555 1855 559 1859
rect 839 1855 843 1859
rect 1199 1855 1200 1859
rect 1200 1855 1203 1859
rect 1343 1855 1344 1859
rect 1344 1855 1347 1859
rect 1403 1855 1407 1859
rect 1539 1855 1543 1859
rect 1683 1855 1687 1859
rect 159 1846 163 1850
rect 303 1846 307 1850
rect 447 1846 451 1850
rect 599 1846 603 1850
rect 751 1846 755 1850
rect 903 1846 907 1850
rect 1055 1846 1059 1850
rect 1207 1846 1211 1850
rect 1351 1846 1355 1850
rect 1487 1846 1491 1850
rect 1631 1846 1635 1850
rect 1751 1846 1755 1850
rect 1871 1845 1875 1849
rect 1895 1848 1899 1852
rect 1991 1848 1995 1852
rect 2119 1848 2123 1852
rect 2247 1848 2251 1852
rect 2383 1848 2387 1852
rect 2519 1848 2523 1852
rect 2655 1848 2659 1852
rect 2807 1848 2811 1852
rect 2975 1848 2979 1852
rect 3151 1848 3155 1852
rect 3335 1848 3339 1852
rect 3503 1848 3507 1852
rect 3591 1845 3595 1849
rect 1963 1839 1967 1843
rect 1971 1839 1975 1843
rect 2191 1839 2195 1843
rect 2343 1839 2347 1843
rect 2351 1839 2355 1843
rect 2595 1839 2599 1843
rect 2731 1839 2735 1843
rect 2899 1839 2903 1843
rect 3051 1839 3055 1843
rect 3251 1839 3255 1843
rect 3259 1839 3263 1843
rect 3503 1835 3507 1839
rect 111 1828 115 1832
rect 1831 1828 1835 1832
rect 1871 1828 1875 1832
rect 3591 1828 3595 1832
rect 211 1819 215 1823
rect 327 1819 331 1823
rect 455 1819 459 1823
rect 839 1819 843 1823
rect 1079 1819 1083 1823
rect 1403 1819 1407 1823
rect 1539 1819 1543 1823
rect 1683 1819 1687 1823
rect 111 1811 115 1815
rect 151 1808 155 1812
rect 295 1808 299 1812
rect 439 1808 443 1812
rect 591 1808 595 1812
rect 743 1808 747 1812
rect 895 1808 899 1812
rect 1047 1808 1051 1812
rect 1199 1808 1203 1812
rect 1343 1808 1347 1812
rect 1479 1808 1483 1812
rect 1623 1808 1627 1812
rect 1743 1808 1747 1812
rect 1831 1811 1835 1815
rect 1903 1810 1907 1814
rect 1999 1810 2003 1814
rect 2127 1810 2131 1814
rect 2255 1810 2259 1814
rect 2391 1810 2395 1814
rect 2527 1810 2531 1814
rect 2663 1810 2667 1814
rect 2815 1810 2819 1814
rect 2983 1810 2987 1814
rect 3159 1810 3163 1814
rect 3343 1810 3347 1814
rect 3511 1810 3515 1814
rect 1911 1799 1915 1803
rect 1963 1799 1967 1803
rect 2191 1799 2195 1803
rect 2343 1799 2347 1803
rect 2535 1799 2539 1803
rect 2595 1799 2599 1803
rect 2731 1799 2735 1803
rect 2899 1799 2903 1803
rect 3051 1799 3055 1803
rect 3251 1799 3255 1803
rect 3527 1799 3531 1803
rect 767 1791 771 1795
rect 1971 1783 1975 1787
rect 1955 1775 1959 1779
rect 2083 1775 2087 1779
rect 2243 1775 2247 1779
rect 2411 1775 2415 1779
rect 2695 1775 2699 1779
rect 2739 1775 2743 1779
rect 2891 1775 2895 1779
rect 3035 1775 3039 1779
rect 3171 1775 3175 1779
rect 3307 1775 3311 1779
rect 3503 1775 3504 1779
rect 3504 1775 3507 1779
rect 1903 1766 1907 1770
rect 2031 1766 2035 1770
rect 2191 1766 2195 1770
rect 2359 1766 2363 1770
rect 2527 1766 2531 1770
rect 2687 1766 2691 1770
rect 2839 1766 2843 1770
rect 2983 1766 2987 1770
rect 3119 1766 3123 1770
rect 3255 1766 3259 1770
rect 3391 1766 3395 1770
rect 3511 1766 3515 1770
rect 111 1757 115 1761
rect 247 1760 251 1764
rect 423 1760 427 1764
rect 591 1760 595 1764
rect 751 1760 755 1764
rect 895 1760 899 1764
rect 1023 1760 1027 1764
rect 1143 1760 1147 1764
rect 1263 1760 1267 1764
rect 1391 1760 1395 1764
rect 1831 1757 1835 1761
rect 343 1751 347 1755
rect 431 1747 435 1751
rect 583 1751 587 1755
rect 679 1751 683 1755
rect 967 1751 971 1755
rect 1091 1751 1095 1755
rect 1211 1751 1215 1755
rect 1335 1751 1339 1755
rect 1343 1751 1347 1755
rect 1871 1748 1875 1752
rect 3591 1748 3595 1752
rect 111 1740 115 1744
rect 1831 1740 1835 1744
rect 1955 1739 1959 1743
rect 2083 1739 2087 1743
rect 2243 1739 2247 1743
rect 2411 1739 2415 1743
rect 2739 1739 2743 1743
rect 2891 1739 2895 1743
rect 3035 1739 3039 1743
rect 3171 1739 3175 1743
rect 3307 1739 3311 1743
rect 1871 1731 1875 1735
rect 1895 1728 1899 1732
rect 2023 1728 2027 1732
rect 2183 1728 2187 1732
rect 2351 1728 2355 1732
rect 2519 1728 2523 1732
rect 2679 1728 2683 1732
rect 2831 1728 2835 1732
rect 2975 1728 2979 1732
rect 3111 1728 3115 1732
rect 3247 1728 3251 1732
rect 3383 1728 3387 1732
rect 3503 1728 3507 1732
rect 3591 1731 3595 1735
rect 255 1722 259 1726
rect 431 1722 435 1726
rect 599 1722 603 1726
rect 759 1722 763 1726
rect 903 1722 907 1726
rect 1031 1722 1035 1726
rect 1151 1722 1155 1726
rect 1271 1722 1275 1726
rect 1399 1722 1403 1726
rect 343 1711 347 1715
rect 679 1711 683 1715
rect 767 1711 771 1715
rect 911 1711 915 1715
rect 967 1711 971 1715
rect 1091 1711 1095 1715
rect 1235 1711 1239 1715
rect 1335 1711 1339 1715
rect 2419 1711 2423 1715
rect 3399 1711 3400 1715
rect 3400 1711 3403 1715
rect 3519 1711 3520 1715
rect 3520 1711 3523 1715
rect 455 1703 459 1707
rect 175 1695 179 1699
rect 243 1695 247 1699
rect 363 1695 367 1699
rect 583 1695 584 1699
rect 584 1695 587 1699
rect 643 1695 647 1699
rect 795 1695 799 1699
rect 947 1695 951 1699
rect 1243 1695 1247 1699
rect 1379 1695 1383 1699
rect 1635 1695 1639 1699
rect 1727 1695 1731 1699
rect 191 1686 195 1690
rect 311 1686 315 1690
rect 447 1686 451 1690
rect 591 1686 595 1690
rect 743 1686 747 1690
rect 895 1686 899 1690
rect 1039 1686 1043 1690
rect 1183 1686 1187 1690
rect 1319 1686 1323 1690
rect 1447 1686 1451 1690
rect 1575 1686 1579 1690
rect 1711 1686 1715 1690
rect 1871 1677 1875 1681
rect 1895 1680 1899 1684
rect 1991 1680 1995 1684
rect 2135 1680 2139 1684
rect 2295 1680 2299 1684
rect 2471 1680 2475 1684
rect 2647 1680 2651 1684
rect 2815 1680 2819 1684
rect 2967 1680 2971 1684
rect 3111 1680 3115 1684
rect 3247 1680 3251 1684
rect 3383 1680 3387 1684
rect 3503 1680 3507 1684
rect 3591 1677 3595 1681
rect 111 1668 115 1672
rect 1831 1668 1835 1672
rect 1963 1671 1967 1675
rect 2071 1671 2075 1675
rect 2223 1671 2227 1675
rect 2391 1671 2395 1675
rect 2567 1671 2571 1675
rect 2575 1671 2579 1675
rect 2891 1671 2895 1675
rect 3047 1671 3051 1675
rect 3179 1671 3183 1675
rect 3187 1671 3191 1675
rect 3323 1671 3327 1675
rect 243 1659 247 1663
rect 363 1659 367 1663
rect 455 1659 459 1663
rect 643 1659 647 1663
rect 795 1659 799 1663
rect 947 1659 951 1663
rect 1235 1659 1239 1663
rect 1243 1659 1247 1663
rect 1379 1659 1383 1663
rect 1635 1659 1639 1663
rect 1871 1660 1875 1664
rect 3591 1660 3595 1664
rect 111 1651 115 1655
rect 183 1648 187 1652
rect 303 1648 307 1652
rect 439 1648 443 1652
rect 583 1648 587 1652
rect 735 1648 739 1652
rect 887 1648 891 1652
rect 1031 1648 1035 1652
rect 1175 1648 1179 1652
rect 1311 1648 1315 1652
rect 1439 1648 1443 1652
rect 1567 1648 1571 1652
rect 1703 1648 1707 1652
rect 1831 1651 1835 1655
rect 1903 1642 1907 1646
rect 1999 1642 2003 1646
rect 2143 1642 2147 1646
rect 2303 1642 2307 1646
rect 2479 1642 2483 1646
rect 2655 1642 2659 1646
rect 2823 1642 2827 1646
rect 2975 1642 2979 1646
rect 3119 1642 3123 1646
rect 3255 1642 3259 1646
rect 3391 1642 3395 1646
rect 3511 1642 3515 1646
rect 919 1631 923 1635
rect 1911 1631 1915 1635
rect 1963 1631 1967 1635
rect 2071 1631 2075 1635
rect 2223 1631 2227 1635
rect 2391 1631 2395 1635
rect 2567 1631 2571 1635
rect 2831 1631 2835 1635
rect 2891 1631 2895 1635
rect 3047 1631 3051 1635
rect 3323 1631 3327 1635
rect 3399 1631 3403 1635
rect 3519 1631 3523 1635
rect 2575 1623 2579 1627
rect 2027 1615 2031 1619
rect 2199 1615 2203 1619
rect 2283 1615 2287 1619
rect 2419 1615 2423 1619
rect 3063 1623 3067 1627
rect 2691 1615 2695 1619
rect 2867 1615 2871 1619
rect 3375 1623 3379 1627
rect 3179 1615 3183 1619
rect 3291 1615 3295 1619
rect 3487 1615 3491 1619
rect 1975 1606 1979 1610
rect 2095 1606 2099 1610
rect 2231 1606 2235 1610
rect 2367 1606 2371 1610
rect 2503 1606 2507 1610
rect 2639 1606 2643 1610
rect 2775 1606 2779 1610
rect 2911 1606 2915 1610
rect 3055 1606 3059 1610
rect 3207 1606 3211 1610
rect 3367 1606 3371 1610
rect 3511 1606 3515 1610
rect 111 1593 115 1597
rect 167 1596 171 1600
rect 351 1596 355 1600
rect 543 1596 547 1600
rect 727 1596 731 1600
rect 903 1596 907 1600
rect 1071 1596 1075 1600
rect 1223 1596 1227 1600
rect 1359 1596 1363 1600
rect 1495 1596 1499 1600
rect 1623 1596 1627 1600
rect 1743 1596 1747 1600
rect 1831 1593 1835 1597
rect 175 1583 179 1587
rect 235 1587 239 1591
rect 419 1587 423 1591
rect 611 1587 615 1591
rect 795 1587 799 1591
rect 1155 1587 1159 1591
rect 1291 1587 1295 1591
rect 1427 1587 1431 1591
rect 1567 1587 1571 1591
rect 1691 1587 1695 1591
rect 1727 1587 1731 1591
rect 1871 1588 1875 1592
rect 3591 1588 3595 1592
rect 111 1576 115 1580
rect 1831 1576 1835 1580
rect 2027 1579 2031 1583
rect 2199 1579 2203 1583
rect 2283 1579 2287 1583
rect 2419 1579 2423 1583
rect 2691 1579 2695 1583
rect 2867 1579 2871 1583
rect 2935 1579 2939 1583
rect 3063 1579 3067 1583
rect 3291 1579 3295 1583
rect 3375 1579 3379 1583
rect 3527 1579 3531 1583
rect 1871 1571 1875 1575
rect 1967 1568 1971 1572
rect 2087 1568 2091 1572
rect 2223 1568 2227 1572
rect 2359 1568 2363 1572
rect 2495 1568 2499 1572
rect 2631 1568 2635 1572
rect 2767 1568 2771 1572
rect 2903 1568 2907 1572
rect 3047 1568 3051 1572
rect 3199 1568 3203 1572
rect 3359 1568 3363 1572
rect 3503 1568 3507 1572
rect 3591 1571 3595 1575
rect 175 1558 179 1562
rect 359 1558 363 1562
rect 551 1558 555 1562
rect 735 1558 739 1562
rect 911 1558 915 1562
rect 1079 1558 1083 1562
rect 1231 1558 1235 1562
rect 1367 1558 1371 1562
rect 1503 1558 1507 1562
rect 1631 1558 1635 1562
rect 1751 1558 1755 1562
rect 235 1547 239 1551
rect 299 1547 303 1551
rect 611 1547 615 1551
rect 795 1547 799 1551
rect 919 1547 923 1551
rect 1155 1547 1159 1551
rect 1291 1547 1295 1551
rect 1427 1547 1431 1551
rect 1567 1547 1571 1551
rect 1691 1547 1695 1551
rect 2419 1551 2423 1555
rect 1479 1539 1483 1543
rect 195 1531 199 1535
rect 419 1531 423 1535
rect 435 1531 439 1535
rect 579 1531 583 1535
rect 723 1531 727 1535
rect 959 1531 963 1535
rect 1003 1531 1007 1535
rect 1131 1531 1135 1535
rect 1259 1531 1263 1535
rect 1387 1531 1391 1535
rect 143 1522 147 1526
rect 247 1522 251 1526
rect 383 1522 387 1526
rect 527 1522 531 1526
rect 671 1522 675 1526
rect 815 1522 819 1526
rect 951 1522 955 1526
rect 1079 1522 1083 1526
rect 1207 1522 1211 1526
rect 1335 1522 1339 1526
rect 1471 1522 1475 1526
rect 1871 1517 1875 1521
rect 2087 1520 2091 1524
rect 2167 1520 2171 1524
rect 2255 1520 2259 1524
rect 2343 1520 2347 1524
rect 2439 1520 2443 1524
rect 2535 1520 2539 1524
rect 2647 1520 2651 1524
rect 2783 1520 2787 1524
rect 2943 1520 2947 1524
rect 3119 1520 3123 1524
rect 3303 1520 3307 1524
rect 3495 1520 3499 1524
rect 3591 1517 3595 1521
rect 2155 1511 2159 1515
rect 2235 1511 2239 1515
rect 2323 1511 2327 1515
rect 2411 1511 2415 1515
rect 2507 1511 2511 1515
rect 111 1504 115 1508
rect 1831 1504 1835 1508
rect 2515 1507 2519 1511
rect 2723 1511 2727 1515
rect 2851 1511 2855 1515
rect 3039 1511 3043 1515
rect 3195 1511 3199 1515
rect 3203 1511 3207 1515
rect 1871 1500 1875 1504
rect 195 1495 199 1499
rect 299 1495 303 1499
rect 435 1495 439 1499
rect 579 1495 583 1499
rect 723 1495 727 1499
rect 1003 1495 1007 1499
rect 1131 1495 1135 1499
rect 1259 1495 1263 1499
rect 1387 1495 1391 1499
rect 3591 1500 3595 1504
rect 1479 1495 1483 1499
rect 111 1487 115 1491
rect 135 1484 139 1488
rect 239 1484 243 1488
rect 375 1484 379 1488
rect 519 1484 523 1488
rect 663 1484 667 1488
rect 807 1484 811 1488
rect 943 1484 947 1488
rect 1071 1484 1075 1488
rect 1199 1484 1203 1488
rect 1327 1484 1331 1488
rect 1463 1484 1467 1488
rect 1831 1487 1835 1491
rect 2095 1482 2099 1486
rect 2175 1482 2179 1486
rect 2263 1482 2267 1486
rect 2351 1482 2355 1486
rect 2447 1482 2451 1486
rect 2543 1482 2547 1486
rect 2655 1482 2659 1486
rect 2791 1482 2795 1486
rect 2951 1482 2955 1486
rect 3127 1482 3131 1486
rect 3311 1482 3315 1486
rect 3503 1482 3507 1486
rect 615 1467 619 1471
rect 2103 1471 2107 1475
rect 2155 1471 2159 1475
rect 2235 1471 2239 1475
rect 2323 1471 2327 1475
rect 2411 1471 2415 1475
rect 2507 1471 2511 1475
rect 2663 1471 2667 1475
rect 2723 1471 2727 1475
rect 2935 1471 2939 1475
rect 3039 1471 3043 1475
rect 3195 1471 3199 1475
rect 2271 1455 2275 1459
rect 2315 1455 2319 1459
rect 2395 1455 2399 1459
rect 2475 1455 2479 1459
rect 2667 1455 2671 1459
rect 2843 1455 2847 1459
rect 2851 1455 2855 1459
rect 3071 1455 3072 1459
rect 3072 1455 3075 1459
rect 3191 1455 3195 1459
rect 2263 1446 2267 1450
rect 2343 1446 2347 1450
rect 2423 1446 2427 1450
rect 2503 1446 2507 1450
rect 2607 1446 2611 1450
rect 2735 1446 2739 1450
rect 2895 1446 2899 1450
rect 3079 1446 3083 1450
rect 3279 1446 3283 1450
rect 3479 1446 3483 1450
rect 111 1433 115 1437
rect 135 1436 139 1440
rect 231 1436 235 1440
rect 359 1436 363 1440
rect 479 1436 483 1440
rect 599 1436 603 1440
rect 719 1436 723 1440
rect 831 1436 835 1440
rect 935 1436 939 1440
rect 1039 1436 1043 1440
rect 1143 1436 1147 1440
rect 1255 1436 1259 1440
rect 1831 1433 1835 1437
rect 203 1427 207 1431
rect 299 1427 303 1431
rect 427 1427 431 1431
rect 547 1427 551 1431
rect 787 1427 791 1431
rect 899 1427 903 1431
rect 1003 1427 1007 1431
rect 1107 1427 1111 1431
rect 1211 1427 1215 1431
rect 1219 1427 1223 1431
rect 1871 1428 1875 1432
rect 3591 1428 3595 1432
rect 111 1416 115 1420
rect 1831 1416 1835 1420
rect 2315 1419 2319 1423
rect 2395 1419 2399 1423
rect 2475 1419 2479 1423
rect 2667 1419 2671 1423
rect 3071 1419 3075 1423
rect 3191 1419 3195 1423
rect 3287 1419 3291 1423
rect 1871 1411 1875 1415
rect 2255 1408 2259 1412
rect 2335 1408 2339 1412
rect 2415 1408 2419 1412
rect 2495 1408 2499 1412
rect 2599 1408 2603 1412
rect 2727 1408 2731 1412
rect 2887 1408 2891 1412
rect 3071 1408 3075 1412
rect 3271 1408 3275 1412
rect 3471 1408 3475 1412
rect 3591 1411 3595 1415
rect 143 1398 147 1402
rect 203 1395 207 1399
rect 239 1398 243 1402
rect 367 1398 371 1402
rect 487 1398 491 1402
rect 607 1398 611 1402
rect 727 1398 731 1402
rect 839 1398 843 1402
rect 943 1398 947 1402
rect 1047 1398 1051 1402
rect 1151 1398 1155 1402
rect 1263 1398 1267 1402
rect 195 1387 199 1391
rect 427 1387 431 1391
rect 547 1387 551 1391
rect 615 1387 619 1391
rect 787 1387 791 1391
rect 899 1387 903 1391
rect 1003 1387 1007 1391
rect 1107 1387 1111 1391
rect 1211 1387 1215 1391
rect 2607 1391 2611 1395
rect 3415 1391 3419 1395
rect 1175 1379 1179 1383
rect 299 1359 303 1363
rect 339 1359 343 1363
rect 143 1350 147 1354
rect 287 1350 291 1354
rect 431 1350 435 1354
rect 583 1350 587 1354
rect 635 1359 639 1363
rect 787 1359 791 1363
rect 931 1359 935 1363
rect 1075 1359 1079 1363
rect 1551 1359 1555 1363
rect 1871 1361 1875 1365
rect 2263 1364 2267 1368
rect 2343 1364 2347 1368
rect 2423 1364 2427 1368
rect 2503 1364 2507 1368
rect 2591 1364 2595 1368
rect 2695 1364 2699 1368
rect 2807 1364 2811 1368
rect 2919 1364 2923 1368
rect 3039 1364 3043 1368
rect 3159 1364 3163 1368
rect 3279 1364 3283 1368
rect 3399 1364 3403 1368
rect 3503 1364 3507 1368
rect 3591 1361 3595 1365
rect 2331 1355 2335 1359
rect 663 1351 667 1355
rect 735 1350 739 1354
rect 879 1350 883 1354
rect 1023 1350 1027 1354
rect 1167 1350 1171 1354
rect 1319 1350 1323 1354
rect 1471 1350 1475 1354
rect 2415 1355 2419 1359
rect 1623 1350 1627 1354
rect 2423 1351 2427 1355
rect 2583 1355 2587 1359
rect 2659 1355 2663 1359
rect 2763 1355 2767 1359
rect 2771 1355 2775 1359
rect 2987 1355 2991 1359
rect 3039 1351 3043 1355
rect 3227 1355 3231 1359
rect 3235 1355 3239 1359
rect 3347 1355 3351 1359
rect 3487 1355 3491 1359
rect 1871 1344 1875 1348
rect 3591 1344 3595 1348
rect 111 1332 115 1336
rect 1831 1332 1835 1336
rect 2323 1335 2327 1339
rect 2771 1335 2775 1339
rect 195 1323 199 1327
rect 339 1323 343 1327
rect 635 1323 639 1327
rect 787 1323 791 1327
rect 931 1323 935 1327
rect 1075 1323 1079 1327
rect 1175 1323 1179 1327
rect 1343 1323 1347 1327
rect 1551 1323 1555 1327
rect 2271 1326 2275 1330
rect 2351 1326 2355 1330
rect 2431 1326 2435 1330
rect 2511 1326 2515 1330
rect 2599 1326 2603 1330
rect 2703 1326 2707 1330
rect 2815 1326 2819 1330
rect 2927 1326 2931 1330
rect 3047 1326 3051 1330
rect 3167 1326 3171 1330
rect 3287 1326 3291 1330
rect 3407 1326 3411 1330
rect 3511 1326 3515 1330
rect 111 1315 115 1319
rect 135 1312 139 1316
rect 279 1312 283 1316
rect 423 1312 427 1316
rect 575 1312 579 1316
rect 727 1312 731 1316
rect 871 1312 875 1316
rect 1015 1312 1019 1316
rect 1159 1312 1163 1316
rect 1311 1312 1315 1316
rect 1463 1312 1467 1316
rect 1615 1312 1619 1316
rect 1831 1315 1835 1319
rect 2323 1315 2327 1319
rect 2331 1315 2335 1319
rect 2415 1307 2419 1311
rect 2607 1315 2611 1319
rect 2659 1315 2663 1319
rect 2763 1315 2767 1319
rect 2839 1315 2843 1319
rect 2987 1315 2991 1319
rect 3235 1315 3239 1319
rect 3347 1315 3351 1319
rect 3415 1315 3419 1319
rect 3519 1315 3523 1319
rect 439 1295 440 1299
rect 440 1295 443 1299
rect 2671 1299 2675 1303
rect 2279 1291 2283 1295
rect 2359 1291 2363 1295
rect 2423 1291 2427 1295
rect 2655 1291 2656 1295
rect 2656 1291 2659 1295
rect 2851 1291 2855 1295
rect 2999 1291 3003 1295
rect 3039 1291 3043 1295
rect 3227 1291 3231 1295
rect 3267 1291 3271 1295
rect 2215 1282 2219 1286
rect 2295 1282 2299 1286
rect 2375 1282 2379 1286
rect 2455 1282 2459 1286
rect 2551 1282 2555 1286
rect 2663 1282 2667 1286
rect 2791 1282 2795 1286
rect 2927 1282 2931 1286
rect 3071 1282 3075 1286
rect 3215 1282 3219 1286
rect 3367 1282 3371 1286
rect 3511 1282 3515 1286
rect 111 1261 115 1265
rect 135 1264 139 1268
rect 263 1264 267 1268
rect 423 1264 427 1268
rect 591 1264 595 1268
rect 759 1264 763 1268
rect 927 1264 931 1268
rect 1079 1264 1083 1268
rect 1223 1264 1227 1268
rect 1351 1264 1355 1268
rect 1479 1264 1483 1268
rect 1607 1264 1611 1268
rect 1735 1264 1739 1268
rect 1831 1261 1835 1265
rect 1871 1264 1875 1268
rect 3591 1264 3595 1268
rect 499 1255 503 1259
rect 507 1255 511 1259
rect 663 1255 667 1259
rect 827 1255 831 1259
rect 1159 1255 1163 1259
rect 1291 1255 1295 1259
rect 1551 1255 1555 1259
rect 111 1244 115 1248
rect 1283 1247 1287 1251
rect 1539 1247 1543 1251
rect 2279 1255 2283 1259
rect 2359 1255 2363 1259
rect 2655 1255 2659 1259
rect 2671 1255 2675 1259
rect 2851 1255 2855 1259
rect 2999 1255 3003 1259
rect 3267 1255 3271 1259
rect 3519 1255 3523 1259
rect 1831 1244 1835 1248
rect 1871 1247 1875 1251
rect 2207 1244 2211 1248
rect 2287 1244 2291 1248
rect 2367 1244 2371 1248
rect 2447 1244 2451 1248
rect 2543 1244 2547 1248
rect 2655 1244 2659 1248
rect 2783 1244 2787 1248
rect 2919 1244 2923 1248
rect 3063 1244 3067 1248
rect 3207 1244 3211 1248
rect 3359 1244 3363 1248
rect 3503 1244 3507 1248
rect 3591 1247 3595 1251
rect 143 1226 147 1230
rect 271 1226 275 1230
rect 431 1226 435 1230
rect 599 1226 603 1230
rect 767 1226 771 1230
rect 935 1226 939 1230
rect 1087 1226 1091 1230
rect 1231 1226 1235 1230
rect 1359 1226 1363 1230
rect 1487 1226 1491 1230
rect 1615 1226 1619 1230
rect 1743 1226 1747 1230
rect 2127 1227 2131 1231
rect 2663 1227 2667 1231
rect 3367 1227 3371 1231
rect 195 1215 199 1219
rect 439 1215 443 1219
rect 499 1215 503 1219
rect 827 1215 831 1219
rect 899 1215 903 1219
rect 1095 1215 1099 1219
rect 1159 1215 1163 1219
rect 1343 1215 1347 1219
rect 1539 1215 1543 1219
rect 1551 1215 1555 1219
rect 1759 1215 1763 1219
rect 423 1195 427 1199
rect 507 1195 511 1199
rect 539 1195 543 1199
rect 855 1195 859 1199
rect 1303 1203 1307 1207
rect 1059 1195 1063 1199
rect 1283 1195 1287 1199
rect 1571 1203 1575 1207
rect 1467 1195 1471 1199
rect 1587 1195 1591 1199
rect 1707 1195 1711 1199
rect 1871 1193 1875 1197
rect 2111 1196 2115 1200
rect 2207 1196 2211 1200
rect 2303 1196 2307 1200
rect 2407 1196 2411 1200
rect 2527 1196 2531 1200
rect 2647 1196 2651 1200
rect 2775 1196 2779 1200
rect 2911 1196 2915 1200
rect 3055 1196 3059 1200
rect 3199 1196 3203 1200
rect 3343 1196 3347 1200
rect 3495 1196 3499 1200
rect 3591 1193 3595 1197
rect 143 1186 147 1190
rect 311 1186 315 1190
rect 487 1186 491 1190
rect 671 1186 675 1190
rect 847 1186 851 1190
rect 1007 1186 1011 1190
rect 1159 1186 1163 1190
rect 1295 1186 1299 1190
rect 1415 1186 1419 1190
rect 1535 1186 1539 1190
rect 1655 1186 1659 1190
rect 1751 1186 1755 1190
rect 2179 1187 2183 1191
rect 2275 1187 2279 1191
rect 2371 1187 2375 1191
rect 2475 1187 2479 1191
rect 2483 1187 2487 1191
rect 2719 1187 2723 1191
rect 2851 1187 2855 1191
rect 2991 1187 2995 1191
rect 2999 1187 3003 1191
rect 3275 1187 3279 1191
rect 3283 1187 3287 1191
rect 1871 1176 1875 1180
rect 3591 1176 3595 1180
rect 111 1168 115 1172
rect 1831 1168 1835 1172
rect 195 1159 199 1163
rect 539 1159 543 1163
rect 679 1159 683 1163
rect 899 1159 903 1163
rect 1059 1159 1063 1163
rect 1211 1159 1215 1163
rect 1303 1159 1307 1163
rect 1467 1159 1471 1163
rect 1587 1159 1591 1163
rect 1707 1159 1711 1163
rect 1759 1159 1763 1163
rect 2119 1158 2123 1162
rect 2215 1158 2219 1162
rect 2311 1158 2315 1162
rect 2415 1158 2419 1162
rect 2535 1158 2539 1162
rect 2655 1158 2659 1162
rect 2783 1158 2787 1162
rect 2919 1158 2923 1162
rect 3063 1158 3067 1162
rect 3207 1158 3211 1162
rect 3351 1158 3355 1162
rect 3503 1158 3507 1162
rect 111 1151 115 1155
rect 135 1148 139 1152
rect 303 1148 307 1152
rect 479 1148 483 1152
rect 663 1148 667 1152
rect 839 1148 843 1152
rect 999 1148 1003 1152
rect 1151 1148 1155 1152
rect 1287 1148 1291 1152
rect 1407 1148 1411 1152
rect 1527 1148 1531 1152
rect 1647 1148 1651 1152
rect 1743 1148 1747 1152
rect 1831 1151 1835 1155
rect 2127 1147 2131 1151
rect 2179 1147 2183 1151
rect 2275 1147 2279 1151
rect 2371 1147 2375 1151
rect 2475 1147 2479 1151
rect 2663 1147 2667 1151
rect 2719 1147 2723 1151
rect 2851 1147 2855 1151
rect 2991 1147 2995 1151
rect 3283 1147 3287 1151
rect 3367 1147 3371 1151
rect 3519 1147 3523 1151
rect 263 1131 267 1135
rect 2483 1127 2487 1131
rect 2583 1127 2587 1131
rect 2627 1127 2631 1131
rect 2827 1127 2831 1131
rect 3255 1127 3259 1131
rect 3275 1127 3279 1131
rect 1903 1118 1907 1122
rect 2127 1118 2131 1122
rect 2359 1118 2363 1122
rect 2575 1118 2579 1122
rect 2775 1118 2779 1122
rect 2967 1118 2971 1122
rect 3159 1118 3163 1122
rect 3343 1118 3347 1122
rect 3511 1118 3515 1122
rect 111 1101 115 1105
rect 135 1104 139 1108
rect 247 1104 251 1108
rect 383 1104 387 1108
rect 519 1104 523 1108
rect 647 1104 651 1108
rect 775 1104 779 1108
rect 895 1104 899 1108
rect 1015 1104 1019 1108
rect 1135 1104 1139 1108
rect 1255 1104 1259 1108
rect 1375 1104 1379 1108
rect 1503 1104 1507 1108
rect 1631 1104 1635 1108
rect 1743 1104 1747 1108
rect 1831 1101 1835 1105
rect 1871 1100 1875 1104
rect 315 1095 319 1099
rect 459 1095 463 1099
rect 111 1084 115 1088
rect 719 1095 723 1099
rect 855 1095 859 1099
rect 963 1095 967 1099
rect 1083 1095 1087 1099
rect 1323 1095 1327 1099
rect 1443 1095 1447 1099
rect 1195 1087 1199 1091
rect 1571 1095 1575 1099
rect 3591 1100 3595 1104
rect 1699 1095 1703 1099
rect 2215 1091 2219 1095
rect 2627 1091 2631 1095
rect 2827 1091 2831 1095
rect 3019 1091 3023 1095
rect 3211 1091 3215 1095
rect 3255 1091 3259 1095
rect 3519 1091 3523 1095
rect 1831 1084 1835 1088
rect 1871 1083 1875 1087
rect 1895 1080 1899 1084
rect 2119 1080 2123 1084
rect 2351 1080 2355 1084
rect 2567 1080 2571 1084
rect 2767 1080 2771 1084
rect 2959 1080 2963 1084
rect 3151 1080 3155 1084
rect 3335 1080 3339 1084
rect 3503 1080 3507 1084
rect 3591 1083 3595 1087
rect 143 1066 147 1070
rect 255 1066 259 1070
rect 391 1066 395 1070
rect 527 1066 531 1070
rect 655 1066 659 1070
rect 783 1066 787 1070
rect 903 1066 907 1070
rect 1023 1066 1027 1070
rect 1143 1066 1147 1070
rect 1263 1066 1267 1070
rect 1383 1066 1387 1070
rect 1511 1066 1515 1070
rect 1639 1066 1643 1070
rect 1751 1066 1755 1070
rect 151 1055 155 1059
rect 263 1055 267 1059
rect 315 1055 319 1059
rect 459 1055 463 1059
rect 627 1055 631 1059
rect 719 1055 723 1059
rect 963 1055 967 1059
rect 1083 1055 1087 1059
rect 1195 1055 1199 1059
rect 1211 1055 1215 1059
rect 1323 1055 1327 1059
rect 1443 1055 1447 1059
rect 1699 1055 1703 1059
rect 299 1031 303 1035
rect 679 1039 683 1043
rect 535 1031 539 1035
rect 687 1031 691 1035
rect 819 1031 823 1035
rect 935 1031 936 1035
rect 936 1031 939 1035
rect 995 1031 999 1035
rect 1083 1031 1087 1035
rect 1179 1031 1183 1035
rect 1871 1033 1875 1037
rect 1895 1036 1899 1040
rect 2015 1036 2019 1040
rect 2167 1036 2171 1040
rect 2327 1036 2331 1040
rect 2487 1036 2491 1040
rect 2639 1036 2643 1040
rect 2791 1036 2795 1040
rect 2935 1036 2939 1040
rect 3079 1036 3083 1040
rect 3223 1036 3227 1040
rect 3375 1036 3379 1040
rect 3503 1036 3507 1040
rect 3591 1033 3595 1037
rect 143 1022 147 1026
rect 239 1022 243 1026
rect 359 1022 363 1026
rect 471 1022 475 1026
rect 575 1022 579 1026
rect 671 1022 675 1026
rect 767 1022 771 1026
rect 855 1022 859 1026
rect 943 1022 947 1026
rect 1031 1022 1035 1026
rect 1127 1022 1131 1026
rect 1963 1027 1967 1031
rect 2083 1027 2087 1031
rect 2415 1027 2419 1031
rect 2707 1027 2711 1031
rect 2859 1027 2863 1031
rect 3003 1027 3007 1031
rect 3307 1027 3311 1031
rect 1223 1022 1227 1026
rect 1871 1016 1875 1020
rect 3591 1016 3595 1020
rect 111 1004 115 1008
rect 1831 1004 1835 1008
rect 151 995 155 999
rect 299 995 303 999
rect 535 995 539 999
rect 627 995 631 999
rect 679 995 683 999
rect 819 995 823 999
rect 935 995 939 999
rect 995 995 999 999
rect 1083 995 1087 999
rect 1179 995 1183 999
rect 1903 998 1907 1002
rect 2023 998 2027 1002
rect 2175 998 2179 1002
rect 2335 998 2339 1002
rect 2495 998 2499 1002
rect 2647 998 2651 1002
rect 2799 998 2803 1002
rect 2943 998 2947 1002
rect 3087 998 3091 1002
rect 3231 998 3235 1002
rect 3383 998 3387 1002
rect 3511 998 3515 1002
rect 111 987 115 991
rect 135 984 139 988
rect 231 984 235 988
rect 351 984 355 988
rect 463 984 467 988
rect 567 984 571 988
rect 663 984 667 988
rect 759 984 763 988
rect 847 984 851 988
rect 935 984 939 988
rect 1023 984 1027 988
rect 1119 984 1123 988
rect 1215 984 1219 988
rect 1831 987 1835 991
rect 1963 987 1967 991
rect 2083 987 2087 991
rect 2207 987 2211 991
rect 2215 987 2219 991
rect 2415 987 2419 991
rect 2707 987 2711 991
rect 2859 987 2863 991
rect 3003 987 3007 991
rect 3019 987 3023 991
rect 3211 987 3215 991
rect 3307 987 3311 991
rect 3519 987 3523 991
rect 1955 971 1959 975
rect 2035 971 2039 975
rect 2131 971 2135 975
rect 2407 971 2411 975
rect 2683 971 2687 975
rect 2843 971 2847 975
rect 3211 971 3215 975
rect 1903 962 1907 966
rect 1983 962 1987 966
rect 2079 962 2083 966
rect 2199 962 2203 966
rect 2335 962 2339 966
rect 2479 962 2483 966
rect 2631 962 2635 966
rect 2791 962 2795 966
rect 2967 962 2971 966
rect 3151 962 3155 966
rect 3343 962 3347 966
rect 3511 962 3515 966
rect 1871 944 1875 948
rect 3591 944 3595 948
rect 1955 935 1959 939
rect 2035 935 2039 939
rect 2131 935 2135 939
rect 2207 935 2211 939
rect 2407 935 2411 939
rect 2683 935 2687 939
rect 2843 935 2847 939
rect 3203 935 3207 939
rect 3211 935 3215 939
rect 3519 935 3523 939
rect 111 925 115 929
rect 135 928 139 932
rect 263 928 267 932
rect 415 928 419 932
rect 559 928 563 932
rect 703 928 707 932
rect 839 928 843 932
rect 975 928 979 932
rect 1103 928 1107 932
rect 1223 928 1227 932
rect 1335 928 1339 932
rect 1439 928 1443 932
rect 1543 928 1547 932
rect 1655 928 1659 932
rect 1743 928 1747 932
rect 1831 925 1835 929
rect 1871 927 1875 931
rect 1895 924 1899 928
rect 339 919 343 923
rect 495 919 499 923
rect 635 919 639 923
rect 687 919 691 923
rect 779 919 783 923
rect 1043 919 1047 923
rect 1171 919 1175 923
rect 1403 919 1407 923
rect 1507 919 1511 923
rect 1611 919 1615 923
rect 1975 924 1979 928
rect 2071 924 2075 928
rect 2191 924 2195 928
rect 2327 924 2331 928
rect 2471 924 2475 928
rect 2623 924 2627 928
rect 2783 924 2787 928
rect 2959 924 2963 928
rect 3143 924 3147 928
rect 3335 924 3339 928
rect 3503 924 3507 928
rect 3591 927 3595 931
rect 1723 919 1727 923
rect 1743 915 1747 919
rect 111 908 115 912
rect 1831 908 1835 912
rect 2311 907 2315 911
rect 2879 907 2883 911
rect 143 890 147 894
rect 271 890 275 894
rect 423 890 427 894
rect 567 890 571 894
rect 711 890 715 894
rect 847 890 851 894
rect 983 890 987 894
rect 1111 890 1115 894
rect 1231 890 1235 894
rect 1343 890 1347 894
rect 1447 890 1451 894
rect 1551 890 1555 894
rect 1663 890 1667 894
rect 1751 890 1755 894
rect 151 879 155 883
rect 339 879 343 883
rect 495 879 499 883
rect 779 879 783 883
rect 839 879 840 883
rect 840 879 843 883
rect 1043 879 1047 883
rect 1171 879 1175 883
rect 1391 879 1395 883
rect 1403 879 1407 883
rect 1507 879 1511 883
rect 1611 879 1615 883
rect 1723 879 1727 883
rect 203 863 207 867
rect 259 863 263 867
rect 367 863 371 867
rect 435 863 439 867
rect 635 863 639 867
rect 1011 863 1015 867
rect 1155 863 1159 867
rect 1647 871 1651 875
rect 1519 863 1523 867
rect 1563 863 1567 867
rect 1743 863 1744 867
rect 1744 863 1747 867
rect 1871 865 1875 869
rect 1919 868 1923 872
rect 2095 868 2099 872
rect 2271 868 2275 872
rect 2455 868 2459 872
rect 2655 868 2659 872
rect 2863 868 2867 872
rect 3079 868 3083 872
rect 3303 868 3307 872
rect 3503 868 3507 872
rect 3591 865 3595 869
rect 143 854 147 858
rect 247 854 251 858
rect 383 854 387 858
rect 519 854 523 858
rect 663 854 667 858
rect 815 854 819 858
rect 959 854 963 858
rect 1103 854 1107 858
rect 1247 854 1251 858
rect 1383 854 1387 858
rect 1511 854 1515 858
rect 1639 854 1643 858
rect 1987 859 1991 863
rect 2723 859 2727 863
rect 2931 859 2935 863
rect 3195 859 3199 863
rect 1751 854 1755 858
rect 1871 848 1875 852
rect 3591 848 3595 852
rect 111 836 115 840
rect 1831 836 1835 840
rect 151 827 155 831
rect 203 827 207 831
rect 435 827 439 831
rect 527 827 531 831
rect 839 827 843 831
rect 1011 827 1015 831
rect 1155 827 1159 831
rect 1391 827 1395 831
rect 1563 827 1567 831
rect 1647 827 1651 831
rect 1927 830 1931 834
rect 2103 830 2107 834
rect 2279 830 2283 834
rect 2463 830 2467 834
rect 2663 830 2667 834
rect 2871 830 2875 834
rect 3087 830 3091 834
rect 3311 830 3315 834
rect 3511 830 3515 834
rect 111 819 115 823
rect 135 816 139 820
rect 239 816 243 820
rect 375 816 379 820
rect 511 816 515 820
rect 655 816 659 820
rect 807 816 811 820
rect 951 816 955 820
rect 1095 816 1099 820
rect 1239 816 1243 820
rect 1375 816 1379 820
rect 1503 816 1507 820
rect 1631 816 1635 820
rect 1743 816 1747 820
rect 1831 819 1835 823
rect 1987 819 1991 823
rect 2311 819 2315 823
rect 2723 819 2727 823
rect 2879 819 2883 823
rect 3195 819 3199 823
rect 3203 819 3207 823
rect 3519 819 3523 823
rect 1955 807 1959 811
rect 2067 807 2071 811
rect 2219 807 2223 811
rect 2379 807 2383 811
rect 2931 807 2935 811
rect 2979 807 2983 811
rect 3011 807 3015 811
rect 3155 807 3159 811
rect 3299 807 3303 811
rect 1159 799 1163 803
rect 1903 798 1907 802
rect 2015 798 2019 802
rect 2167 798 2171 802
rect 2327 798 2331 802
rect 2487 798 2491 802
rect 2647 798 2651 802
rect 2807 798 2811 802
rect 2959 798 2963 802
rect 3103 798 3107 802
rect 3247 798 3251 802
rect 3391 798 3395 802
rect 3511 798 3515 802
rect 1871 780 1875 784
rect 3591 780 3595 784
rect 1955 771 1959 775
rect 2067 771 2071 775
rect 2219 771 2223 775
rect 2379 771 2383 775
rect 2699 771 2703 775
rect 2871 771 2875 775
rect 3011 771 3015 775
rect 3155 771 3159 775
rect 3299 771 3303 775
rect 3519 771 3523 775
rect 111 757 115 761
rect 135 760 139 764
rect 215 760 219 764
rect 303 760 307 764
rect 415 760 419 764
rect 543 760 547 764
rect 687 760 691 764
rect 839 760 843 764
rect 991 760 995 764
rect 1143 760 1147 764
rect 1295 760 1299 764
rect 1447 760 1451 764
rect 1607 760 1611 764
rect 1871 763 1875 767
rect 1831 757 1835 761
rect 1895 760 1899 764
rect 2007 760 2011 764
rect 2159 760 2163 764
rect 2319 760 2323 764
rect 2479 760 2483 764
rect 2639 760 2643 764
rect 2799 760 2803 764
rect 2951 760 2955 764
rect 3095 760 3099 764
rect 3239 760 3243 764
rect 3383 760 3387 764
rect 3503 760 3507 764
rect 3591 763 3595 767
rect 203 751 207 755
rect 283 751 287 755
rect 371 751 375 755
rect 487 751 491 755
rect 611 751 615 755
rect 655 751 659 755
rect 907 751 911 755
rect 915 751 919 755
rect 1059 751 1063 755
rect 1379 751 1383 755
rect 1519 751 1523 755
rect 1531 751 1535 755
rect 111 740 115 744
rect 1831 740 1835 744
rect 2419 743 2423 747
rect 3375 743 3379 747
rect 143 722 147 726
rect 223 722 227 726
rect 311 722 315 726
rect 423 722 427 726
rect 551 722 555 726
rect 695 722 699 726
rect 847 722 851 726
rect 999 722 1003 726
rect 1151 722 1155 726
rect 1303 722 1307 726
rect 1455 722 1459 726
rect 1615 722 1619 726
rect 151 711 155 715
rect 203 711 207 715
rect 283 711 287 715
rect 431 711 435 715
rect 487 711 491 715
rect 611 711 615 715
rect 915 711 919 715
rect 1059 711 1063 715
rect 1159 711 1163 715
rect 1311 711 1315 715
rect 1379 711 1383 715
rect 1607 711 1608 715
rect 1608 711 1611 715
rect 1871 713 1875 717
rect 1967 716 1971 720
rect 2063 716 2067 720
rect 2175 716 2179 720
rect 2303 716 2307 720
rect 2447 716 2451 720
rect 2599 716 2603 720
rect 2751 716 2755 720
rect 2903 716 2907 720
rect 3055 716 3059 720
rect 3207 716 3211 720
rect 3359 716 3363 720
rect 3503 716 3507 720
rect 3591 713 3595 717
rect 2035 707 2039 711
rect 2131 707 2135 711
rect 2247 707 2251 711
rect 2383 707 2387 711
rect 2607 703 2611 707
rect 2819 707 2823 711
rect 1871 696 1875 700
rect 2979 707 2983 711
rect 3275 707 3279 711
rect 3267 699 3271 703
rect 275 691 279 695
rect 283 691 287 695
rect 371 691 375 695
rect 603 691 607 695
rect 739 691 743 695
rect 855 691 859 695
rect 907 691 911 695
rect 1095 691 1099 695
rect 1139 691 1143 695
rect 1267 691 1271 695
rect 1387 691 1391 695
rect 1507 691 1511 695
rect 3591 696 3595 700
rect 231 682 235 686
rect 319 682 323 686
rect 423 682 427 686
rect 543 682 547 686
rect 679 682 683 686
rect 815 682 819 686
rect 951 682 955 686
rect 1087 682 1091 686
rect 1215 682 1219 686
rect 1335 682 1339 686
rect 1455 682 1459 686
rect 1583 682 1587 686
rect 1975 678 1979 682
rect 2071 678 2075 682
rect 2183 678 2187 682
rect 2311 678 2315 682
rect 2455 678 2459 682
rect 2607 678 2611 682
rect 2759 678 2763 682
rect 2911 678 2915 682
rect 3063 678 3067 682
rect 3215 678 3219 682
rect 3367 678 3371 682
rect 3511 678 3515 682
rect 111 664 115 668
rect 1831 664 1835 668
rect 1983 667 1987 671
rect 2035 667 2039 671
rect 2131 667 2135 671
rect 2247 667 2251 671
rect 2383 667 2387 671
rect 2699 667 2703 671
rect 2871 667 2875 671
rect 3127 667 3131 671
rect 3275 667 3279 671
rect 3375 671 3379 675
rect 3519 667 3523 671
rect 283 655 287 659
rect 371 655 375 659
rect 431 655 435 659
rect 551 655 555 659
rect 603 655 607 659
rect 739 655 743 659
rect 1139 655 1143 659
rect 1267 655 1271 659
rect 1387 655 1391 659
rect 1507 655 1511 659
rect 1607 655 1611 659
rect 2191 655 2195 659
rect 2227 655 2231 659
rect 2323 655 2327 659
rect 2427 655 2431 659
rect 2539 655 2543 659
rect 2819 655 2823 659
rect 2983 655 2984 659
rect 2984 655 2987 659
rect 3267 655 3271 659
rect 3299 655 3303 659
rect 3527 655 3531 659
rect 111 647 115 651
rect 223 644 227 648
rect 311 644 315 648
rect 415 644 419 648
rect 535 644 539 648
rect 671 644 675 648
rect 807 644 811 648
rect 943 644 947 648
rect 1079 644 1083 648
rect 1207 644 1211 648
rect 1327 644 1331 648
rect 1447 644 1451 648
rect 1575 644 1579 648
rect 1831 647 1835 651
rect 2175 646 2179 650
rect 2271 646 2275 650
rect 2375 646 2379 650
rect 2487 646 2491 650
rect 2607 646 2611 650
rect 2735 646 2739 650
rect 2863 646 2867 650
rect 2991 646 2995 650
rect 3119 646 3123 650
rect 3247 646 3251 650
rect 3375 646 3379 650
rect 3511 646 3515 650
rect 1871 628 1875 632
rect 3591 628 3595 632
rect 2227 619 2231 623
rect 2323 619 2327 623
rect 2427 619 2431 623
rect 2539 619 2543 623
rect 2787 619 2791 623
rect 2983 619 2987 623
rect 3043 619 3047 623
rect 3127 619 3131 623
rect 3299 619 3303 623
rect 3427 619 3431 623
rect 3519 619 3523 623
rect 1871 611 1875 615
rect 2167 608 2171 612
rect 2263 608 2267 612
rect 2367 608 2371 612
rect 2479 608 2483 612
rect 2599 608 2603 612
rect 2727 608 2731 612
rect 2855 608 2859 612
rect 2983 608 2987 612
rect 3111 608 3115 612
rect 3239 608 3243 612
rect 3367 608 3371 612
rect 3503 608 3507 612
rect 3591 611 3595 615
rect 111 589 115 593
rect 447 592 451 596
rect 527 592 531 596
rect 607 592 611 596
rect 687 592 691 596
rect 775 592 779 596
rect 871 592 875 596
rect 959 592 963 596
rect 1047 592 1051 596
rect 1143 592 1147 596
rect 1239 592 1243 596
rect 1335 592 1339 596
rect 1431 592 1435 596
rect 1831 589 1835 593
rect 2539 591 2543 595
rect 515 583 519 587
rect 595 583 599 587
rect 675 583 679 587
rect 755 583 759 587
rect 855 583 859 587
rect 863 583 867 587
rect 939 583 943 587
rect 1115 583 1119 587
rect 1211 583 1215 587
rect 1307 583 1311 587
rect 1403 583 1407 587
rect 1411 583 1415 587
rect 111 572 115 576
rect 1831 572 1835 576
rect 1871 561 1875 565
rect 2263 564 2267 568
rect 2343 564 2347 568
rect 2423 564 2427 568
rect 2503 564 2507 568
rect 2591 564 2595 568
rect 2695 564 2699 568
rect 2815 564 2819 568
rect 2959 564 2963 568
rect 3111 564 3115 568
rect 3279 564 3283 568
rect 3447 564 3451 568
rect 3591 561 3595 565
rect 455 554 459 558
rect 535 554 539 558
rect 615 554 619 558
rect 695 554 699 558
rect 783 554 787 558
rect 879 554 883 558
rect 967 554 971 558
rect 1055 554 1059 558
rect 1151 554 1155 558
rect 1247 554 1251 558
rect 1343 554 1347 558
rect 1439 554 1443 558
rect 2331 555 2335 559
rect 2411 555 2415 559
rect 2491 555 2495 559
rect 2571 555 2575 559
rect 2659 555 2663 559
rect 515 543 519 547
rect 595 543 599 547
rect 675 543 679 547
rect 755 543 759 547
rect 939 543 943 547
rect 599 535 603 539
rect 1115 543 1119 547
rect 1211 543 1215 547
rect 1307 543 1311 547
rect 1403 543 1407 547
rect 1871 544 1875 548
rect 2563 547 2567 551
rect 2895 555 2899 559
rect 2755 547 2759 551
rect 3027 555 3031 559
rect 3527 555 3531 559
rect 3591 544 3595 548
rect 1287 535 1291 539
rect 291 519 295 523
rect 387 519 391 523
rect 475 519 479 523
rect 563 519 567 523
rect 863 527 867 531
rect 2271 526 2275 530
rect 2351 526 2355 530
rect 2431 526 2435 530
rect 2511 526 2515 530
rect 2599 526 2603 530
rect 2703 526 2707 530
rect 2823 526 2827 530
rect 2967 526 2971 530
rect 3119 526 3123 530
rect 3287 526 3291 530
rect 3455 526 3459 530
rect 723 519 727 523
rect 855 519 859 523
rect 891 519 895 523
rect 979 519 983 523
rect 1067 519 1071 523
rect 1183 519 1184 523
rect 1184 519 1187 523
rect 1271 519 1272 523
rect 1272 519 1275 523
rect 335 510 339 514
rect 423 510 427 514
rect 511 510 515 514
rect 591 510 595 514
rect 671 510 675 514
rect 751 510 755 514
rect 839 510 843 514
rect 927 510 931 514
rect 1015 510 1019 514
rect 1103 510 1107 514
rect 1191 510 1195 514
rect 2283 515 2287 519
rect 2331 515 2335 519
rect 2411 515 2415 519
rect 2491 515 2495 519
rect 2571 515 2575 519
rect 2659 515 2663 519
rect 2787 515 2791 519
rect 2895 515 2899 519
rect 3043 515 3047 519
rect 3327 515 3331 519
rect 3427 515 3431 519
rect 1279 510 1283 514
rect 111 492 115 496
rect 1831 492 1835 496
rect 2251 495 2255 499
rect 2443 495 2447 499
rect 2563 495 2567 499
rect 2643 495 2647 499
rect 2755 495 2759 499
rect 3027 503 3031 507
rect 2843 495 2847 499
rect 3031 495 3032 499
rect 3032 495 3035 499
rect 3091 495 3095 499
rect 3227 495 3231 499
rect 3391 495 3395 499
rect 387 483 391 487
rect 475 483 479 487
rect 563 483 567 487
rect 599 483 603 487
rect 723 483 727 487
rect 891 483 895 487
rect 979 483 983 487
rect 1067 483 1071 487
rect 1183 483 1187 487
rect 1271 483 1275 487
rect 1287 483 1291 487
rect 2191 486 2195 490
rect 2287 486 2291 490
rect 2383 486 2387 490
rect 2487 486 2491 490
rect 2583 486 2587 490
rect 2687 486 2691 490
rect 2791 486 2795 490
rect 2911 486 2915 490
rect 3039 486 3043 490
rect 3175 486 3179 490
rect 3319 486 3323 490
rect 3471 486 3475 490
rect 111 475 115 479
rect 327 472 331 476
rect 415 472 419 476
rect 503 472 507 476
rect 583 472 587 476
rect 663 472 667 476
rect 743 472 747 476
rect 831 472 835 476
rect 919 472 923 476
rect 1007 472 1011 476
rect 1095 472 1099 476
rect 1183 472 1187 476
rect 1271 472 1275 476
rect 1831 475 1835 479
rect 1871 468 1875 472
rect 3591 468 3595 472
rect 2251 459 2255 463
rect 2443 459 2447 463
rect 2643 459 2647 463
rect 2843 459 2847 463
rect 3031 459 3035 463
rect 3091 459 3095 463
rect 3227 459 3231 463
rect 3327 459 3331 463
rect 1871 451 1875 455
rect 2183 448 2187 452
rect 2279 448 2283 452
rect 2375 448 2379 452
rect 2479 448 2483 452
rect 2575 448 2579 452
rect 2679 448 2683 452
rect 2783 448 2787 452
rect 2903 448 2907 452
rect 3031 448 3035 452
rect 3167 448 3171 452
rect 3311 448 3315 452
rect 3463 448 3467 452
rect 3591 451 3595 455
rect 1991 431 1995 435
rect 2487 431 2491 435
rect 111 417 115 421
rect 223 420 227 424
rect 335 420 339 424
rect 447 420 451 424
rect 559 420 563 424
rect 663 420 667 424
rect 759 420 763 424
rect 847 420 851 424
rect 935 420 939 424
rect 1023 420 1027 424
rect 1111 420 1115 424
rect 1199 420 1203 424
rect 1295 420 1299 424
rect 1831 417 1835 421
rect 291 411 295 415
rect 299 411 303 415
rect 403 411 407 415
rect 731 411 735 415
rect 855 407 859 411
rect 915 411 919 415
rect 1003 411 1007 415
rect 1091 411 1095 415
rect 1267 411 1271 415
rect 111 400 115 404
rect 1171 403 1175 407
rect 1831 400 1835 404
rect 1871 397 1875 401
rect 1975 400 1979 404
rect 2063 400 2067 404
rect 2159 400 2163 404
rect 2255 400 2259 404
rect 2359 400 2363 404
rect 2471 400 2475 404
rect 2607 400 2611 404
rect 2759 400 2763 404
rect 2927 400 2931 404
rect 3111 400 3115 404
rect 3303 400 3307 404
rect 3495 400 3499 404
rect 3591 397 3595 401
rect 2043 391 2047 395
rect 2131 391 2135 395
rect 2227 391 2231 395
rect 231 382 235 386
rect 343 382 347 386
rect 455 382 459 386
rect 567 382 571 386
rect 671 382 675 386
rect 767 382 771 386
rect 855 382 859 386
rect 943 382 947 386
rect 1031 382 1035 386
rect 1119 382 1123 386
rect 1207 382 1211 386
rect 1303 382 1307 386
rect 1871 380 1875 384
rect 2539 391 2543 395
rect 2683 391 2687 395
rect 2851 391 2855 395
rect 3027 391 3031 395
rect 3035 391 3039 395
rect 3391 391 3395 395
rect 3495 387 3499 391
rect 3591 380 3595 384
rect 299 371 303 375
rect 403 371 407 375
rect 447 371 448 375
rect 448 371 451 375
rect 731 371 735 375
rect 915 371 919 375
rect 1003 371 1007 375
rect 1091 371 1095 375
rect 1171 371 1175 375
rect 1179 371 1183 375
rect 1267 371 1271 375
rect 1983 362 1987 366
rect 2071 362 2075 366
rect 2167 362 2171 366
rect 2263 362 2267 366
rect 2367 362 2371 366
rect 2479 362 2483 366
rect 2615 362 2619 366
rect 2767 362 2771 366
rect 2935 362 2939 366
rect 3119 362 3123 366
rect 3311 362 3315 366
rect 3503 362 3507 366
rect 195 347 199 351
rect 315 347 319 351
rect 587 347 591 351
rect 723 347 727 351
rect 1239 355 1243 359
rect 963 347 967 351
rect 1075 347 1079 351
rect 1447 355 1451 359
rect 1311 347 1315 351
rect 1387 347 1391 351
rect 1991 351 1995 355
rect 2043 351 2047 355
rect 2131 351 2135 355
rect 2227 351 2231 355
rect 2487 351 2491 355
rect 2539 351 2543 355
rect 2683 351 2687 355
rect 2851 351 2855 355
rect 3027 351 3031 355
rect 3399 351 3403 355
rect 143 338 147 342
rect 263 338 267 342
rect 399 338 403 342
rect 535 338 539 342
rect 671 338 675 342
rect 791 338 795 342
rect 911 338 915 342
rect 1023 338 1027 342
rect 1127 338 1131 342
rect 1231 338 1235 342
rect 1335 338 1339 342
rect 1439 338 1443 342
rect 2275 335 2279 339
rect 2347 335 2351 339
rect 2435 335 2439 339
rect 2531 335 2535 339
rect 2643 335 2647 339
rect 2907 335 2911 339
rect 3035 335 3039 339
rect 3103 335 3107 339
rect 3171 335 3175 339
rect 3371 335 3375 339
rect 3495 335 3499 339
rect 2215 326 2219 330
rect 2295 326 2299 330
rect 2383 326 2387 330
rect 2479 326 2483 330
rect 2591 326 2595 330
rect 2719 326 2723 330
rect 2847 326 2851 330
rect 2983 326 2987 330
rect 3119 326 3123 330
rect 3255 326 3259 330
rect 3391 326 3395 330
rect 3511 326 3515 330
rect 111 320 115 324
rect 1831 320 1835 324
rect 195 311 199 315
rect 315 311 319 315
rect 447 311 451 315
rect 587 311 591 315
rect 723 311 727 315
rect 839 311 843 315
rect 963 311 967 315
rect 1075 311 1079 315
rect 1179 311 1183 315
rect 1239 311 1243 315
rect 1387 311 1391 315
rect 1447 311 1451 315
rect 1871 308 1875 312
rect 111 303 115 307
rect 3591 308 3595 312
rect 135 300 139 304
rect 255 300 259 304
rect 391 300 395 304
rect 527 300 531 304
rect 663 300 667 304
rect 783 300 787 304
rect 903 300 907 304
rect 1015 300 1019 304
rect 1119 300 1123 304
rect 1223 300 1227 304
rect 1327 300 1331 304
rect 1431 300 1435 304
rect 1831 303 1835 307
rect 2275 299 2279 303
rect 2347 299 2351 303
rect 2435 299 2439 303
rect 2531 299 2535 303
rect 2643 299 2647 303
rect 2899 299 2903 303
rect 2907 299 2911 303
rect 3171 299 3175 303
rect 3371 299 3375 303
rect 3399 299 3403 303
rect 1871 291 1875 295
rect 2207 288 2211 292
rect 2287 288 2291 292
rect 2375 288 2379 292
rect 2471 288 2475 292
rect 2583 288 2587 292
rect 2711 288 2715 292
rect 2839 288 2843 292
rect 2975 288 2979 292
rect 3111 288 3115 292
rect 3247 288 3251 292
rect 3383 288 3387 292
rect 3503 288 3507 292
rect 3591 291 3595 295
rect 2551 271 2555 275
rect 3519 271 3520 275
rect 3520 271 3523 275
rect 111 245 115 249
rect 135 248 139 252
rect 247 248 251 252
rect 391 248 395 252
rect 543 248 547 252
rect 695 248 699 252
rect 847 248 851 252
rect 991 248 995 252
rect 1119 248 1123 252
rect 1239 248 1243 252
rect 1359 248 1363 252
rect 1479 248 1483 252
rect 1599 248 1603 252
rect 1831 245 1835 249
rect 203 239 207 243
rect 315 239 319 243
rect 611 239 615 243
rect 763 239 767 243
rect 1063 239 1067 243
rect 1187 239 1191 243
rect 1311 239 1315 243
rect 1427 239 1431 243
rect 1547 239 1551 243
rect 111 228 115 232
rect 1051 231 1055 235
rect 1871 237 1875 241
rect 1991 240 1995 244
rect 2119 240 2123 244
rect 2255 240 2259 244
rect 2391 240 2395 244
rect 2535 240 2539 244
rect 2679 240 2683 244
rect 2815 240 2819 244
rect 2951 240 2955 244
rect 3095 240 3099 244
rect 3239 240 3243 244
rect 3383 240 3387 244
rect 3503 240 3507 244
rect 3591 237 3595 241
rect 1831 228 1835 232
rect 2063 231 2067 235
rect 2187 231 2191 235
rect 1871 220 1875 224
rect 2051 223 2055 227
rect 2335 231 2339 235
rect 2459 231 2463 235
rect 2747 231 2751 235
rect 2883 231 2887 235
rect 3103 227 3107 231
rect 3195 231 3199 235
rect 3307 231 3311 235
rect 3503 227 3507 231
rect 3591 220 3595 224
rect 143 210 147 214
rect 255 210 259 214
rect 399 210 403 214
rect 551 210 555 214
rect 703 210 707 214
rect 855 210 859 214
rect 999 210 1003 214
rect 1127 210 1131 214
rect 1247 210 1251 214
rect 1367 210 1371 214
rect 1487 210 1491 214
rect 1607 210 1611 214
rect 203 199 207 203
rect 315 199 319 203
rect 355 199 359 203
rect 763 199 767 203
rect 839 199 843 203
rect 1051 199 1055 203
rect 1063 199 1067 203
rect 1187 199 1191 203
rect 1359 199 1360 203
rect 1360 199 1363 203
rect 1427 199 1431 203
rect 1547 199 1551 203
rect 1999 202 2003 206
rect 2127 202 2131 206
rect 2263 202 2267 206
rect 2399 202 2403 206
rect 2543 202 2547 206
rect 2687 202 2691 206
rect 2823 202 2827 206
rect 2959 202 2963 206
rect 3103 202 3107 206
rect 3247 202 3251 206
rect 3391 202 3395 206
rect 3511 202 3515 206
rect 2051 191 2055 195
rect 2063 191 2067 195
rect 2335 191 2339 195
rect 2459 191 2463 195
rect 2551 191 2555 195
rect 2747 191 2751 195
rect 2883 191 2887 195
rect 2899 191 2903 195
rect 3195 191 3199 195
rect 3307 191 3311 195
rect 3383 191 3384 195
rect 3384 191 3387 195
rect 3519 191 3523 195
rect 1963 167 1967 171
rect 2043 167 2047 171
rect 2495 175 2499 179
rect 2187 167 2191 171
rect 2319 167 2323 171
rect 2479 167 2480 171
rect 2480 167 2483 171
rect 2675 167 2679 171
rect 2795 167 2799 171
rect 2907 167 2911 171
rect 3011 167 3015 171
rect 3115 167 3119 171
rect 3211 167 3215 171
rect 3299 167 3303 171
rect 3491 167 3495 171
rect 3503 167 3504 171
rect 3504 167 3507 171
rect 391 159 395 163
rect 791 159 795 163
rect 195 151 199 155
rect 275 151 279 155
rect 443 151 447 155
rect 523 151 527 155
rect 611 151 615 155
rect 675 151 679 155
rect 755 151 759 155
rect 1111 159 1115 163
rect 1903 158 1907 162
rect 1983 158 1987 162
rect 2087 158 2091 162
rect 2215 158 2219 162
rect 2351 158 2355 162
rect 2487 158 2491 162
rect 2623 158 2627 162
rect 2743 158 2747 162
rect 2855 158 2859 162
rect 2959 158 2963 162
rect 3063 158 3067 162
rect 3159 158 3163 162
rect 3247 158 3251 162
rect 3343 158 3347 162
rect 3431 158 3435 162
rect 3511 158 3515 162
rect 915 151 919 155
rect 1007 151 1011 155
rect 1163 151 1167 155
rect 1323 151 1327 155
rect 1403 151 1407 155
rect 1571 151 1575 155
rect 1651 151 1655 155
rect 1731 151 1735 155
rect 1803 151 1807 155
rect 143 142 147 146
rect 223 142 227 146
rect 303 142 307 146
rect 383 142 387 146
rect 463 142 467 146
rect 543 142 547 146
rect 623 142 627 146
rect 703 142 707 146
rect 783 142 787 146
rect 863 142 867 146
rect 943 142 947 146
rect 1023 142 1027 146
rect 1103 142 1107 146
rect 1183 142 1187 146
rect 1263 142 1267 146
rect 1343 142 1347 146
rect 1423 142 1427 146
rect 1511 142 1515 146
rect 1591 142 1595 146
rect 1671 142 1675 146
rect 1751 142 1755 146
rect 1871 140 1875 144
rect 3591 140 3595 144
rect 1803 131 1807 135
rect 1963 131 1967 135
rect 2043 131 2047 135
rect 2319 131 2323 135
rect 2479 131 2483 135
rect 2495 131 2499 135
rect 2675 131 2679 135
rect 2795 131 2799 135
rect 2907 131 2911 135
rect 3011 131 3015 135
rect 3115 131 3119 135
rect 3211 131 3215 135
rect 3299 131 3303 135
rect 3383 131 3387 135
rect 3491 131 3495 135
rect 111 124 115 128
rect 1831 124 1835 128
rect 1871 123 1875 127
rect 1895 120 1899 124
rect 195 115 199 119
rect 275 115 279 119
rect 355 115 359 119
rect 391 115 395 119
rect 443 115 447 119
rect 523 115 527 119
rect 675 115 679 119
rect 755 115 759 119
rect 791 115 795 119
rect 915 115 919 119
rect 1007 115 1011 119
rect 1075 115 1079 119
rect 1111 115 1115 119
rect 1163 115 1167 119
rect 1323 115 1327 119
rect 1403 115 1407 119
rect 1571 115 1575 119
rect 1651 115 1655 119
rect 1975 120 1979 124
rect 2079 120 2083 124
rect 2207 120 2211 124
rect 2343 120 2347 124
rect 2479 120 2483 124
rect 2615 120 2619 124
rect 2735 120 2739 124
rect 2847 120 2851 124
rect 2951 120 2955 124
rect 3055 120 3059 124
rect 3151 120 3155 124
rect 3239 120 3243 124
rect 3335 120 3339 124
rect 3423 120 3427 124
rect 3503 120 3507 124
rect 3591 123 3595 127
rect 1731 115 1735 119
rect 111 107 115 111
rect 135 104 139 108
rect 215 104 219 108
rect 295 104 299 108
rect 375 104 379 108
rect 455 104 459 108
rect 535 104 539 108
rect 615 104 619 108
rect 695 104 699 108
rect 775 104 779 108
rect 855 104 859 108
rect 935 104 939 108
rect 1015 104 1019 108
rect 1095 104 1099 108
rect 1175 104 1179 108
rect 1255 104 1259 108
rect 1335 104 1339 108
rect 1415 104 1419 108
rect 1503 104 1507 108
rect 1583 104 1587 108
rect 1663 104 1667 108
rect 1743 104 1747 108
rect 1831 107 1835 111
<< m3 >>
rect 111 3670 115 3671
rect 111 3665 115 3666
rect 135 3670 139 3671
rect 135 3665 139 3666
rect 215 3670 219 3671
rect 215 3665 219 3666
rect 295 3670 299 3671
rect 295 3665 299 3666
rect 1831 3670 1835 3671
rect 1831 3665 1835 3666
rect 112 3646 114 3665
rect 136 3649 138 3665
rect 216 3649 218 3665
rect 296 3649 298 3665
rect 134 3648 140 3649
rect 110 3645 116 3646
rect 110 3641 111 3645
rect 115 3641 116 3645
rect 134 3644 135 3648
rect 139 3644 140 3648
rect 134 3643 140 3644
rect 214 3648 220 3649
rect 214 3644 215 3648
rect 219 3644 220 3648
rect 214 3643 220 3644
rect 294 3648 300 3649
rect 294 3644 295 3648
rect 299 3644 300 3648
rect 1832 3646 1834 3665
rect 294 3643 300 3644
rect 1830 3645 1836 3646
rect 110 3640 116 3641
rect 1830 3641 1831 3645
rect 1835 3641 1836 3645
rect 1830 3640 1836 3641
rect 202 3639 208 3640
rect 134 3635 140 3636
rect 134 3631 135 3635
rect 139 3631 140 3635
rect 202 3635 203 3639
rect 207 3635 208 3639
rect 202 3634 208 3635
rect 282 3639 288 3640
rect 282 3635 283 3639
rect 287 3635 288 3639
rect 282 3634 288 3635
rect 134 3630 140 3631
rect 110 3628 116 3629
rect 110 3624 111 3628
rect 115 3624 116 3628
rect 110 3623 116 3624
rect 112 3595 114 3623
rect 111 3594 115 3595
rect 111 3589 115 3590
rect 112 3561 114 3589
rect 136 3588 138 3630
rect 142 3610 148 3611
rect 142 3606 143 3610
rect 147 3606 148 3610
rect 142 3605 148 3606
rect 144 3595 146 3605
rect 204 3600 206 3634
rect 222 3610 228 3611
rect 222 3606 223 3610
rect 227 3606 228 3610
rect 222 3605 228 3606
rect 202 3599 208 3600
rect 202 3595 203 3599
rect 207 3595 208 3599
rect 224 3595 226 3605
rect 284 3600 286 3634
rect 1830 3628 1836 3629
rect 1830 3624 1831 3628
rect 1835 3624 1836 3628
rect 1830 3623 1836 3624
rect 302 3610 308 3611
rect 302 3606 303 3610
rect 307 3606 308 3610
rect 302 3605 308 3606
rect 282 3599 288 3600
rect 282 3595 283 3599
rect 287 3595 288 3599
rect 304 3595 306 3605
rect 1832 3595 1834 3623
rect 2826 3603 2832 3604
rect 1871 3602 1875 3603
rect 1871 3597 1875 3598
rect 2063 3602 2067 3603
rect 2063 3597 2067 3598
rect 2151 3602 2155 3603
rect 2151 3597 2155 3598
rect 2255 3602 2259 3603
rect 2255 3597 2259 3598
rect 2367 3602 2371 3603
rect 2367 3597 2371 3598
rect 2479 3602 2483 3603
rect 2479 3597 2483 3598
rect 2591 3602 2595 3603
rect 2591 3597 2595 3598
rect 2703 3602 2707 3603
rect 2703 3597 2707 3598
rect 2815 3602 2819 3603
rect 2826 3599 2827 3603
rect 2831 3599 2832 3603
rect 2826 3598 2832 3599
rect 2919 3602 2923 3603
rect 2815 3597 2819 3598
rect 143 3594 147 3595
rect 202 3594 208 3595
rect 223 3594 227 3595
rect 282 3594 288 3595
rect 303 3594 307 3595
rect 143 3589 147 3590
rect 223 3589 227 3590
rect 303 3589 307 3590
rect 343 3594 347 3595
rect 343 3589 347 3590
rect 471 3594 475 3595
rect 471 3589 475 3590
rect 607 3594 611 3595
rect 607 3589 611 3590
rect 743 3594 747 3595
rect 743 3589 747 3590
rect 879 3594 883 3595
rect 879 3589 883 3590
rect 999 3594 1003 3595
rect 999 3589 1003 3590
rect 1111 3594 1115 3595
rect 1111 3589 1115 3590
rect 1223 3594 1227 3595
rect 1223 3589 1227 3590
rect 1327 3594 1331 3595
rect 1327 3589 1331 3590
rect 1423 3594 1427 3595
rect 1423 3589 1427 3590
rect 1527 3594 1531 3595
rect 1527 3589 1531 3590
rect 1631 3594 1635 3595
rect 1631 3589 1635 3590
rect 1831 3594 1835 3595
rect 1831 3589 1835 3590
rect 134 3587 140 3588
rect 134 3583 135 3587
rect 139 3583 140 3587
rect 134 3582 140 3583
rect 144 3579 146 3589
rect 194 3587 200 3588
rect 194 3583 195 3587
rect 199 3583 200 3587
rect 194 3582 200 3583
rect 142 3578 148 3579
rect 142 3574 143 3578
rect 147 3574 148 3578
rect 142 3573 148 3574
rect 110 3560 116 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 196 3552 198 3582
rect 224 3579 226 3589
rect 274 3587 280 3588
rect 274 3583 275 3587
rect 279 3583 280 3587
rect 274 3582 280 3583
rect 222 3578 228 3579
rect 222 3574 223 3578
rect 227 3574 228 3578
rect 222 3573 228 3574
rect 276 3552 278 3582
rect 344 3579 346 3589
rect 394 3587 400 3588
rect 394 3583 395 3587
rect 399 3583 400 3587
rect 394 3582 400 3583
rect 342 3578 348 3579
rect 342 3574 343 3578
rect 347 3574 348 3578
rect 342 3573 348 3574
rect 396 3552 398 3582
rect 472 3579 474 3589
rect 522 3587 528 3588
rect 522 3583 523 3587
rect 527 3583 528 3587
rect 522 3582 528 3583
rect 470 3578 476 3579
rect 470 3574 471 3578
rect 475 3574 476 3578
rect 470 3573 476 3574
rect 524 3552 526 3582
rect 608 3579 610 3589
rect 658 3587 664 3588
rect 658 3583 659 3587
rect 663 3583 664 3587
rect 658 3582 664 3583
rect 606 3578 612 3579
rect 606 3574 607 3578
rect 611 3574 612 3578
rect 606 3573 612 3574
rect 660 3552 662 3582
rect 744 3579 746 3589
rect 880 3579 882 3589
rect 886 3587 892 3588
rect 886 3583 887 3587
rect 891 3583 892 3587
rect 886 3582 892 3583
rect 930 3587 936 3588
rect 930 3583 931 3587
rect 935 3583 936 3587
rect 930 3582 936 3583
rect 742 3578 748 3579
rect 742 3574 743 3578
rect 747 3574 748 3578
rect 742 3573 748 3574
rect 878 3578 884 3579
rect 878 3574 879 3578
rect 883 3574 884 3578
rect 878 3573 884 3574
rect 194 3551 200 3552
rect 194 3547 195 3551
rect 199 3547 200 3551
rect 194 3546 200 3547
rect 274 3551 280 3552
rect 274 3547 275 3551
rect 279 3547 280 3551
rect 274 3546 280 3547
rect 394 3551 400 3552
rect 394 3547 395 3551
rect 399 3547 400 3551
rect 394 3546 400 3547
rect 522 3551 528 3552
rect 522 3547 523 3551
rect 527 3547 528 3551
rect 522 3546 528 3547
rect 658 3551 664 3552
rect 658 3547 659 3551
rect 663 3547 664 3551
rect 658 3546 664 3547
rect 766 3551 772 3552
rect 766 3547 767 3551
rect 771 3547 772 3551
rect 766 3546 772 3547
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 110 3538 116 3539
rect 134 3540 140 3541
rect 112 3519 114 3538
rect 134 3536 135 3540
rect 139 3536 140 3540
rect 134 3535 140 3536
rect 214 3540 220 3541
rect 214 3536 215 3540
rect 219 3536 220 3540
rect 214 3535 220 3536
rect 334 3540 340 3541
rect 334 3536 335 3540
rect 339 3536 340 3540
rect 334 3535 340 3536
rect 462 3540 468 3541
rect 462 3536 463 3540
rect 467 3536 468 3540
rect 462 3535 468 3536
rect 598 3540 604 3541
rect 598 3536 599 3540
rect 603 3536 604 3540
rect 598 3535 604 3536
rect 734 3540 740 3541
rect 734 3536 735 3540
rect 739 3536 740 3540
rect 734 3535 740 3536
rect 136 3519 138 3535
rect 216 3519 218 3535
rect 336 3519 338 3535
rect 464 3519 466 3535
rect 600 3519 602 3535
rect 736 3519 738 3535
rect 111 3518 115 3519
rect 111 3513 115 3514
rect 135 3518 139 3519
rect 135 3513 139 3514
rect 191 3518 195 3519
rect 191 3513 195 3514
rect 215 3518 219 3519
rect 215 3513 219 3514
rect 327 3518 331 3519
rect 327 3513 331 3514
rect 335 3518 339 3519
rect 335 3513 339 3514
rect 463 3518 467 3519
rect 463 3513 467 3514
rect 471 3518 475 3519
rect 471 3513 475 3514
rect 599 3518 603 3519
rect 599 3513 603 3514
rect 623 3518 627 3519
rect 623 3513 627 3514
rect 735 3518 739 3519
rect 735 3513 739 3514
rect 112 3494 114 3513
rect 192 3497 194 3513
rect 328 3497 330 3513
rect 472 3497 474 3513
rect 624 3497 626 3513
rect 190 3496 196 3497
rect 110 3493 116 3494
rect 110 3489 111 3493
rect 115 3489 116 3493
rect 190 3492 191 3496
rect 195 3492 196 3496
rect 190 3491 196 3492
rect 326 3496 332 3497
rect 326 3492 327 3496
rect 331 3492 332 3496
rect 326 3491 332 3492
rect 470 3496 476 3497
rect 470 3492 471 3496
rect 475 3492 476 3496
rect 470 3491 476 3492
rect 622 3496 628 3497
rect 622 3492 623 3496
rect 627 3492 628 3496
rect 622 3491 628 3492
rect 110 3488 116 3489
rect 258 3487 264 3488
rect 258 3483 259 3487
rect 263 3483 264 3487
rect 258 3482 264 3483
rect 394 3487 400 3488
rect 394 3483 395 3487
rect 399 3483 400 3487
rect 394 3482 400 3483
rect 538 3487 544 3488
rect 538 3483 539 3487
rect 543 3483 544 3487
rect 538 3482 544 3483
rect 690 3487 696 3488
rect 690 3483 691 3487
rect 695 3483 696 3487
rect 690 3482 696 3483
rect 110 3476 116 3477
rect 110 3472 111 3476
rect 115 3472 116 3476
rect 110 3471 116 3472
rect 112 3443 114 3471
rect 198 3458 204 3459
rect 198 3454 199 3458
rect 203 3454 204 3458
rect 198 3453 204 3454
rect 200 3443 202 3453
rect 260 3448 262 3482
rect 334 3458 340 3459
rect 334 3454 335 3458
rect 339 3454 340 3458
rect 334 3453 340 3454
rect 258 3447 264 3448
rect 258 3443 259 3447
rect 263 3443 264 3447
rect 336 3443 338 3453
rect 396 3448 398 3482
rect 478 3458 484 3459
rect 478 3454 479 3458
rect 483 3454 484 3458
rect 478 3453 484 3454
rect 394 3447 400 3448
rect 394 3443 395 3447
rect 399 3443 400 3447
rect 480 3443 482 3453
rect 540 3448 542 3482
rect 630 3458 636 3459
rect 630 3454 631 3458
rect 635 3454 636 3458
rect 630 3453 636 3454
rect 538 3447 544 3448
rect 538 3443 539 3447
rect 543 3443 544 3447
rect 632 3443 634 3453
rect 692 3448 694 3482
rect 768 3448 770 3546
rect 870 3540 876 3541
rect 870 3536 871 3540
rect 875 3536 876 3540
rect 870 3535 876 3536
rect 872 3519 874 3535
rect 775 3518 779 3519
rect 775 3513 779 3514
rect 871 3518 875 3519
rect 871 3513 875 3514
rect 776 3497 778 3513
rect 774 3496 780 3497
rect 774 3492 775 3496
rect 779 3492 780 3496
rect 774 3491 780 3492
rect 888 3488 890 3582
rect 932 3552 934 3582
rect 1000 3579 1002 3589
rect 1050 3587 1056 3588
rect 1050 3583 1051 3587
rect 1055 3583 1056 3587
rect 1050 3582 1056 3583
rect 998 3578 1004 3579
rect 998 3574 999 3578
rect 1003 3574 1004 3578
rect 998 3573 1004 3574
rect 1052 3552 1054 3582
rect 1112 3579 1114 3589
rect 1162 3587 1168 3588
rect 1162 3583 1163 3587
rect 1167 3583 1168 3587
rect 1162 3582 1168 3583
rect 1110 3578 1116 3579
rect 1110 3574 1111 3578
rect 1115 3574 1116 3578
rect 1110 3573 1116 3574
rect 1164 3552 1166 3582
rect 1224 3579 1226 3589
rect 1274 3587 1280 3588
rect 1274 3583 1275 3587
rect 1279 3583 1280 3587
rect 1274 3582 1280 3583
rect 1222 3578 1228 3579
rect 1222 3574 1223 3578
rect 1227 3574 1228 3578
rect 1222 3573 1228 3574
rect 1276 3552 1278 3582
rect 1328 3579 1330 3589
rect 1378 3587 1384 3588
rect 1378 3583 1379 3587
rect 1383 3583 1384 3587
rect 1378 3582 1384 3583
rect 1326 3578 1332 3579
rect 1326 3574 1327 3578
rect 1331 3574 1332 3578
rect 1326 3573 1332 3574
rect 1380 3552 1382 3582
rect 1424 3579 1426 3589
rect 1474 3587 1480 3588
rect 1474 3583 1475 3587
rect 1479 3583 1480 3587
rect 1474 3582 1480 3583
rect 1422 3578 1428 3579
rect 1422 3574 1423 3578
rect 1427 3574 1428 3578
rect 1422 3573 1428 3574
rect 1476 3552 1478 3582
rect 1528 3579 1530 3589
rect 1578 3587 1584 3588
rect 1578 3583 1579 3587
rect 1583 3583 1584 3587
rect 1578 3582 1584 3583
rect 1526 3578 1532 3579
rect 1526 3574 1527 3578
rect 1531 3574 1532 3578
rect 1526 3573 1532 3574
rect 1580 3552 1582 3582
rect 1632 3579 1634 3589
rect 1630 3578 1636 3579
rect 1630 3574 1631 3578
rect 1635 3574 1636 3578
rect 1630 3573 1636 3574
rect 1832 3561 1834 3589
rect 1872 3569 1874 3597
rect 2064 3587 2066 3597
rect 2070 3595 2076 3596
rect 2070 3591 2071 3595
rect 2075 3591 2076 3595
rect 2070 3590 2076 3591
rect 2114 3595 2120 3596
rect 2114 3591 2115 3595
rect 2119 3591 2120 3595
rect 2114 3590 2120 3591
rect 2062 3586 2068 3587
rect 2062 3582 2063 3586
rect 2067 3582 2068 3586
rect 2062 3581 2068 3582
rect 1870 3568 1876 3569
rect 1870 3564 1871 3568
rect 1875 3564 1876 3568
rect 1870 3563 1876 3564
rect 1830 3560 1836 3561
rect 1830 3556 1831 3560
rect 1835 3556 1836 3560
rect 1830 3555 1836 3556
rect 930 3551 936 3552
rect 930 3547 931 3551
rect 935 3547 936 3551
rect 930 3546 936 3547
rect 1050 3551 1056 3552
rect 1050 3547 1051 3551
rect 1055 3547 1056 3551
rect 1050 3546 1056 3547
rect 1162 3551 1168 3552
rect 1162 3547 1163 3551
rect 1167 3547 1168 3551
rect 1162 3546 1168 3547
rect 1274 3551 1280 3552
rect 1274 3547 1275 3551
rect 1279 3547 1280 3551
rect 1274 3546 1280 3547
rect 1378 3551 1384 3552
rect 1378 3547 1379 3551
rect 1383 3547 1384 3551
rect 1378 3546 1384 3547
rect 1474 3551 1480 3552
rect 1474 3547 1475 3551
rect 1479 3547 1480 3551
rect 1474 3546 1480 3547
rect 1578 3551 1584 3552
rect 1578 3547 1579 3551
rect 1583 3547 1584 3551
rect 1578 3546 1584 3547
rect 1870 3551 1876 3552
rect 1870 3547 1871 3551
rect 1875 3547 1876 3551
rect 1870 3546 1876 3547
rect 2054 3548 2060 3549
rect 1830 3543 1836 3544
rect 990 3540 996 3541
rect 990 3536 991 3540
rect 995 3536 996 3540
rect 990 3535 996 3536
rect 1102 3540 1108 3541
rect 1102 3536 1103 3540
rect 1107 3536 1108 3540
rect 1102 3535 1108 3536
rect 1214 3540 1220 3541
rect 1214 3536 1215 3540
rect 1219 3536 1220 3540
rect 1214 3535 1220 3536
rect 1318 3540 1324 3541
rect 1318 3536 1319 3540
rect 1323 3536 1324 3540
rect 1318 3535 1324 3536
rect 1414 3540 1420 3541
rect 1414 3536 1415 3540
rect 1419 3536 1420 3540
rect 1414 3535 1420 3536
rect 1518 3540 1524 3541
rect 1518 3536 1519 3540
rect 1523 3536 1524 3540
rect 1518 3535 1524 3536
rect 1622 3540 1628 3541
rect 1622 3536 1623 3540
rect 1627 3536 1628 3540
rect 1830 3539 1831 3543
rect 1835 3539 1836 3543
rect 1830 3538 1836 3539
rect 1622 3535 1628 3536
rect 992 3519 994 3535
rect 1104 3519 1106 3535
rect 1216 3519 1218 3535
rect 1320 3519 1322 3535
rect 1416 3519 1418 3535
rect 1520 3519 1522 3535
rect 1582 3523 1588 3524
rect 1582 3519 1583 3523
rect 1587 3519 1588 3523
rect 1624 3519 1626 3535
rect 1832 3519 1834 3538
rect 1872 3527 1874 3546
rect 2054 3544 2055 3548
rect 2059 3544 2060 3548
rect 2054 3543 2060 3544
rect 2056 3527 2058 3543
rect 1871 3526 1875 3527
rect 1871 3521 1875 3522
rect 2055 3526 2059 3527
rect 2055 3521 2059 3522
rect 919 3518 923 3519
rect 919 3513 923 3514
rect 991 3518 995 3519
rect 991 3513 995 3514
rect 1055 3518 1059 3519
rect 1055 3513 1059 3514
rect 1103 3518 1107 3519
rect 1103 3513 1107 3514
rect 1183 3518 1187 3519
rect 1183 3513 1187 3514
rect 1215 3518 1219 3519
rect 1215 3513 1219 3514
rect 1311 3518 1315 3519
rect 1311 3513 1315 3514
rect 1319 3518 1323 3519
rect 1319 3513 1323 3514
rect 1415 3518 1419 3519
rect 1415 3513 1419 3514
rect 1439 3518 1443 3519
rect 1439 3513 1443 3514
rect 1519 3518 1523 3519
rect 1519 3513 1523 3514
rect 1567 3518 1571 3519
rect 1582 3518 1588 3519
rect 1623 3518 1627 3519
rect 1567 3513 1571 3514
rect 920 3497 922 3513
rect 1056 3497 1058 3513
rect 1184 3497 1186 3513
rect 1312 3497 1314 3513
rect 1440 3497 1442 3513
rect 1568 3497 1570 3513
rect 918 3496 924 3497
rect 918 3492 919 3496
rect 923 3492 924 3496
rect 918 3491 924 3492
rect 1054 3496 1060 3497
rect 1054 3492 1055 3496
rect 1059 3492 1060 3496
rect 1054 3491 1060 3492
rect 1182 3496 1188 3497
rect 1182 3492 1183 3496
rect 1187 3492 1188 3496
rect 1182 3491 1188 3492
rect 1310 3496 1316 3497
rect 1310 3492 1311 3496
rect 1315 3492 1316 3496
rect 1310 3491 1316 3492
rect 1438 3496 1444 3497
rect 1438 3492 1439 3496
rect 1443 3492 1444 3496
rect 1438 3491 1444 3492
rect 1566 3496 1572 3497
rect 1566 3492 1567 3496
rect 1571 3492 1572 3496
rect 1566 3491 1572 3492
rect 886 3487 892 3488
rect 886 3483 887 3487
rect 891 3483 892 3487
rect 886 3482 892 3483
rect 986 3487 992 3488
rect 986 3483 987 3487
rect 991 3483 992 3487
rect 986 3482 992 3483
rect 1126 3487 1132 3488
rect 1126 3483 1127 3487
rect 1131 3483 1132 3487
rect 1126 3482 1132 3483
rect 1378 3487 1384 3488
rect 1378 3483 1379 3487
rect 1383 3483 1384 3487
rect 1378 3482 1384 3483
rect 782 3458 788 3459
rect 782 3454 783 3458
rect 787 3454 788 3458
rect 782 3453 788 3454
rect 926 3458 932 3459
rect 926 3454 927 3458
rect 931 3454 932 3458
rect 926 3453 932 3454
rect 690 3447 696 3448
rect 690 3443 691 3447
rect 695 3443 696 3447
rect 111 3442 115 3443
rect 111 3437 115 3438
rect 151 3442 155 3443
rect 151 3437 155 3438
rect 199 3442 203 3443
rect 258 3442 264 3443
rect 295 3442 299 3443
rect 199 3437 203 3438
rect 295 3437 299 3438
rect 335 3442 339 3443
rect 394 3442 400 3443
rect 455 3442 459 3443
rect 335 3437 339 3438
rect 455 3437 459 3438
rect 479 3442 483 3443
rect 538 3442 544 3443
rect 623 3442 627 3443
rect 479 3437 483 3438
rect 623 3437 627 3438
rect 631 3442 635 3443
rect 690 3442 696 3443
rect 766 3447 772 3448
rect 766 3443 767 3447
rect 771 3443 772 3447
rect 784 3443 786 3453
rect 928 3443 930 3453
rect 988 3448 990 3482
rect 1062 3458 1068 3459
rect 1062 3454 1063 3458
rect 1067 3454 1068 3458
rect 1062 3453 1068 3454
rect 986 3447 992 3448
rect 986 3443 987 3447
rect 991 3443 992 3447
rect 1064 3443 1066 3453
rect 1128 3448 1130 3482
rect 1190 3458 1196 3459
rect 1190 3454 1191 3458
rect 1195 3454 1196 3458
rect 1190 3453 1196 3454
rect 1318 3458 1324 3459
rect 1318 3454 1319 3458
rect 1323 3454 1324 3458
rect 1318 3453 1324 3454
rect 1126 3447 1132 3448
rect 1126 3443 1127 3447
rect 1131 3443 1132 3447
rect 766 3442 772 3443
rect 783 3442 787 3443
rect 631 3437 635 3438
rect 783 3437 787 3438
rect 791 3442 795 3443
rect 791 3437 795 3438
rect 927 3442 931 3443
rect 927 3437 931 3438
rect 959 3442 963 3443
rect 986 3442 992 3443
rect 1063 3442 1067 3443
rect 959 3437 963 3438
rect 1063 3437 1067 3438
rect 1119 3442 1123 3443
rect 1126 3442 1132 3443
rect 1170 3447 1176 3448
rect 1170 3443 1171 3447
rect 1175 3443 1176 3447
rect 1192 3443 1194 3453
rect 1320 3443 1322 3453
rect 1380 3448 1382 3482
rect 1446 3458 1452 3459
rect 1446 3454 1447 3458
rect 1451 3454 1452 3458
rect 1446 3453 1452 3454
rect 1574 3458 1580 3459
rect 1574 3454 1575 3458
rect 1579 3454 1580 3458
rect 1574 3453 1580 3454
rect 1378 3447 1384 3448
rect 1378 3443 1379 3447
rect 1383 3443 1384 3447
rect 1448 3443 1450 3453
rect 1576 3443 1578 3453
rect 1584 3448 1586 3518
rect 1623 3513 1627 3514
rect 1831 3518 1835 3519
rect 1831 3513 1835 3514
rect 1832 3494 1834 3513
rect 1872 3502 1874 3521
rect 1870 3501 1876 3502
rect 1870 3497 1871 3501
rect 1875 3497 1876 3501
rect 1870 3496 1876 3497
rect 2072 3496 2074 3590
rect 2116 3560 2118 3590
rect 2152 3587 2154 3597
rect 2202 3595 2208 3596
rect 2202 3591 2203 3595
rect 2207 3591 2208 3595
rect 2202 3590 2208 3591
rect 2150 3586 2156 3587
rect 2150 3582 2151 3586
rect 2155 3582 2156 3586
rect 2150 3581 2156 3582
rect 2204 3560 2206 3590
rect 2256 3587 2258 3597
rect 2306 3595 2312 3596
rect 2306 3591 2307 3595
rect 2311 3591 2312 3595
rect 2306 3590 2312 3591
rect 2254 3586 2260 3587
rect 2254 3582 2255 3586
rect 2259 3582 2260 3586
rect 2254 3581 2260 3582
rect 2308 3560 2310 3590
rect 2368 3587 2370 3597
rect 2418 3595 2424 3596
rect 2418 3591 2419 3595
rect 2423 3591 2424 3595
rect 2418 3590 2424 3591
rect 2366 3586 2372 3587
rect 2366 3582 2367 3586
rect 2371 3582 2372 3586
rect 2366 3581 2372 3582
rect 2420 3560 2422 3590
rect 2480 3587 2482 3597
rect 2530 3595 2536 3596
rect 2530 3591 2531 3595
rect 2535 3591 2536 3595
rect 2530 3590 2536 3591
rect 2478 3586 2484 3587
rect 2478 3582 2479 3586
rect 2483 3582 2484 3586
rect 2478 3581 2484 3582
rect 2532 3560 2534 3590
rect 2592 3587 2594 3597
rect 2704 3587 2706 3597
rect 2754 3595 2760 3596
rect 2754 3591 2755 3595
rect 2759 3591 2760 3595
rect 2754 3590 2760 3591
rect 2590 3586 2596 3587
rect 2590 3582 2591 3586
rect 2595 3582 2596 3586
rect 2590 3581 2596 3582
rect 2702 3586 2708 3587
rect 2702 3582 2703 3586
rect 2707 3582 2708 3586
rect 2702 3581 2708 3582
rect 2756 3560 2758 3590
rect 2816 3587 2818 3597
rect 2814 3586 2820 3587
rect 2814 3582 2815 3586
rect 2819 3582 2820 3586
rect 2814 3581 2820 3582
rect 2114 3559 2120 3560
rect 2114 3555 2115 3559
rect 2119 3555 2120 3559
rect 2114 3554 2120 3555
rect 2202 3559 2208 3560
rect 2202 3555 2203 3559
rect 2207 3555 2208 3559
rect 2202 3554 2208 3555
rect 2306 3559 2312 3560
rect 2306 3555 2307 3559
rect 2311 3555 2312 3559
rect 2306 3554 2312 3555
rect 2418 3559 2424 3560
rect 2418 3555 2419 3559
rect 2423 3555 2424 3559
rect 2418 3554 2424 3555
rect 2530 3559 2536 3560
rect 2530 3555 2531 3559
rect 2535 3555 2536 3559
rect 2530 3554 2536 3555
rect 2754 3559 2760 3560
rect 2754 3555 2755 3559
rect 2759 3555 2760 3559
rect 2754 3554 2760 3555
rect 2142 3548 2148 3549
rect 2142 3544 2143 3548
rect 2147 3544 2148 3548
rect 2142 3543 2148 3544
rect 2246 3548 2252 3549
rect 2246 3544 2247 3548
rect 2251 3544 2252 3548
rect 2246 3543 2252 3544
rect 2358 3548 2364 3549
rect 2358 3544 2359 3548
rect 2363 3544 2364 3548
rect 2358 3543 2364 3544
rect 2470 3548 2476 3549
rect 2470 3544 2471 3548
rect 2475 3544 2476 3548
rect 2470 3543 2476 3544
rect 2582 3548 2588 3549
rect 2582 3544 2583 3548
rect 2587 3544 2588 3548
rect 2582 3543 2588 3544
rect 2694 3548 2700 3549
rect 2694 3544 2695 3548
rect 2699 3544 2700 3548
rect 2694 3543 2700 3544
rect 2806 3548 2812 3549
rect 2806 3544 2807 3548
rect 2811 3544 2812 3548
rect 2806 3543 2812 3544
rect 2144 3527 2146 3543
rect 2248 3527 2250 3543
rect 2360 3527 2362 3543
rect 2382 3531 2388 3532
rect 2382 3527 2383 3531
rect 2387 3527 2388 3531
rect 2472 3527 2474 3543
rect 2584 3527 2586 3543
rect 2696 3527 2698 3543
rect 2808 3527 2810 3543
rect 2087 3526 2091 3527
rect 2087 3521 2091 3522
rect 2143 3526 2147 3527
rect 2143 3521 2147 3522
rect 2167 3526 2171 3527
rect 2167 3521 2171 3522
rect 2247 3526 2251 3527
rect 2247 3521 2251 3522
rect 2263 3526 2267 3527
rect 2263 3521 2267 3522
rect 2359 3526 2363 3527
rect 2359 3521 2363 3522
rect 2367 3526 2371 3527
rect 2382 3526 2388 3527
rect 2471 3526 2475 3527
rect 2367 3521 2371 3522
rect 2088 3505 2090 3521
rect 2168 3505 2170 3521
rect 2264 3505 2266 3521
rect 2368 3505 2370 3521
rect 2086 3504 2092 3505
rect 2086 3500 2087 3504
rect 2091 3500 2092 3504
rect 2086 3499 2092 3500
rect 2166 3504 2172 3505
rect 2166 3500 2167 3504
rect 2171 3500 2172 3504
rect 2166 3499 2172 3500
rect 2262 3504 2268 3505
rect 2262 3500 2263 3504
rect 2267 3500 2268 3504
rect 2262 3499 2268 3500
rect 2366 3504 2372 3505
rect 2366 3500 2367 3504
rect 2371 3500 2372 3504
rect 2366 3499 2372 3500
rect 2070 3495 2076 3496
rect 1830 3493 1836 3494
rect 1830 3489 1831 3493
rect 1835 3489 1836 3493
rect 2070 3491 2071 3495
rect 2075 3491 2076 3495
rect 2070 3490 2076 3491
rect 2154 3495 2160 3496
rect 2154 3491 2155 3495
rect 2159 3491 2160 3495
rect 2154 3490 2160 3491
rect 2234 3495 2240 3496
rect 2234 3491 2235 3495
rect 2239 3491 2240 3495
rect 2234 3490 2240 3491
rect 1830 3488 1836 3489
rect 1870 3484 1876 3485
rect 1870 3480 1871 3484
rect 1875 3480 1876 3484
rect 1870 3479 1876 3480
rect 1830 3476 1836 3477
rect 1830 3472 1831 3476
rect 1835 3472 1836 3476
rect 1830 3471 1836 3472
rect 1582 3447 1588 3448
rect 1582 3443 1583 3447
rect 1587 3443 1588 3447
rect 1832 3443 1834 3471
rect 1872 3443 1874 3479
rect 2094 3466 2100 3467
rect 2094 3462 2095 3466
rect 2099 3462 2100 3466
rect 2094 3461 2100 3462
rect 2096 3443 2098 3461
rect 2156 3456 2158 3490
rect 2174 3466 2180 3467
rect 2174 3462 2175 3466
rect 2179 3462 2180 3466
rect 2174 3461 2180 3462
rect 2154 3455 2160 3456
rect 2154 3451 2155 3455
rect 2159 3451 2160 3455
rect 2154 3450 2160 3451
rect 2176 3443 2178 3461
rect 2236 3456 2238 3490
rect 2270 3466 2276 3467
rect 2270 3462 2271 3466
rect 2275 3462 2276 3466
rect 2270 3461 2276 3462
rect 2374 3466 2380 3467
rect 2374 3462 2375 3466
rect 2379 3462 2380 3466
rect 2374 3461 2380 3462
rect 2234 3455 2240 3456
rect 2234 3451 2235 3455
rect 2239 3451 2240 3455
rect 2234 3450 2240 3451
rect 2250 3455 2256 3456
rect 2250 3451 2251 3455
rect 2255 3451 2256 3455
rect 2250 3450 2256 3451
rect 1170 3442 1176 3443
rect 1191 3442 1195 3443
rect 1119 3437 1123 3438
rect 112 3409 114 3437
rect 152 3427 154 3437
rect 286 3435 292 3436
rect 286 3431 287 3435
rect 291 3431 292 3435
rect 286 3430 292 3431
rect 150 3426 156 3427
rect 150 3422 151 3426
rect 155 3422 156 3426
rect 150 3421 156 3422
rect 110 3408 116 3409
rect 110 3404 111 3408
rect 115 3404 116 3408
rect 110 3403 116 3404
rect 288 3400 290 3430
rect 296 3427 298 3437
rect 346 3435 352 3436
rect 346 3431 347 3435
rect 351 3431 352 3435
rect 346 3430 352 3431
rect 294 3426 300 3427
rect 294 3422 295 3426
rect 299 3422 300 3426
rect 294 3421 300 3422
rect 348 3400 350 3430
rect 456 3427 458 3437
rect 506 3435 512 3436
rect 506 3431 507 3435
rect 511 3431 512 3435
rect 506 3430 512 3431
rect 454 3426 460 3427
rect 454 3422 455 3426
rect 459 3422 460 3426
rect 454 3421 460 3422
rect 508 3400 510 3430
rect 624 3427 626 3437
rect 674 3435 680 3436
rect 674 3431 675 3435
rect 679 3431 680 3435
rect 674 3430 680 3431
rect 622 3426 628 3427
rect 622 3422 623 3426
rect 627 3422 628 3426
rect 622 3421 628 3422
rect 676 3400 678 3430
rect 792 3427 794 3437
rect 960 3427 962 3437
rect 1010 3435 1016 3436
rect 1010 3431 1011 3435
rect 1015 3431 1016 3435
rect 1010 3430 1016 3431
rect 790 3426 796 3427
rect 790 3422 791 3426
rect 795 3422 796 3426
rect 790 3421 796 3422
rect 958 3426 964 3427
rect 958 3422 959 3426
rect 963 3422 964 3426
rect 958 3421 964 3422
rect 1012 3400 1014 3430
rect 1120 3427 1122 3437
rect 1118 3426 1124 3427
rect 1118 3422 1119 3426
rect 1123 3422 1124 3426
rect 1118 3421 1124 3422
rect 1172 3400 1174 3442
rect 1191 3437 1195 3438
rect 1271 3442 1275 3443
rect 1271 3437 1275 3438
rect 1319 3442 1323 3443
rect 1378 3442 1384 3443
rect 1415 3442 1419 3443
rect 1319 3437 1323 3438
rect 1415 3437 1419 3438
rect 1447 3442 1451 3443
rect 1447 3437 1451 3438
rect 1559 3442 1563 3443
rect 1559 3437 1563 3438
rect 1575 3442 1579 3443
rect 1582 3442 1588 3443
rect 1711 3442 1715 3443
rect 1575 3437 1579 3438
rect 1711 3437 1715 3438
rect 1831 3442 1835 3443
rect 1831 3437 1835 3438
rect 1871 3442 1875 3443
rect 1871 3437 1875 3438
rect 2095 3442 2099 3443
rect 2095 3437 2099 3438
rect 2111 3442 2115 3443
rect 2111 3437 2115 3438
rect 2175 3442 2179 3443
rect 2175 3437 2179 3438
rect 2199 3442 2203 3443
rect 2199 3437 2203 3438
rect 1272 3427 1274 3437
rect 1350 3435 1356 3436
rect 1350 3431 1351 3435
rect 1355 3431 1356 3435
rect 1350 3430 1356 3431
rect 1270 3426 1276 3427
rect 1270 3422 1271 3426
rect 1275 3422 1276 3426
rect 1270 3421 1276 3422
rect 1352 3400 1354 3430
rect 1416 3427 1418 3437
rect 1466 3435 1472 3436
rect 1466 3431 1467 3435
rect 1471 3431 1472 3435
rect 1466 3430 1472 3431
rect 1414 3426 1420 3427
rect 1414 3422 1415 3426
rect 1419 3422 1420 3426
rect 1414 3421 1420 3422
rect 1468 3400 1470 3430
rect 1560 3427 1562 3437
rect 1610 3435 1616 3436
rect 1610 3431 1611 3435
rect 1615 3431 1616 3435
rect 1610 3430 1616 3431
rect 1558 3426 1564 3427
rect 1558 3422 1559 3426
rect 1563 3422 1564 3426
rect 1558 3421 1564 3422
rect 1612 3400 1614 3430
rect 1712 3427 1714 3437
rect 1710 3426 1716 3427
rect 1710 3422 1711 3426
rect 1715 3422 1716 3426
rect 1710 3421 1716 3422
rect 1832 3409 1834 3437
rect 1872 3409 1874 3437
rect 2112 3427 2114 3437
rect 2154 3435 2160 3436
rect 2154 3431 2155 3435
rect 2159 3431 2160 3435
rect 2154 3430 2160 3431
rect 2162 3435 2168 3436
rect 2162 3431 2163 3435
rect 2167 3431 2168 3435
rect 2162 3430 2168 3431
rect 2110 3426 2116 3427
rect 2110 3422 2111 3426
rect 2115 3422 2116 3426
rect 2110 3421 2116 3422
rect 1830 3408 1836 3409
rect 1830 3404 1831 3408
rect 1835 3404 1836 3408
rect 1830 3403 1836 3404
rect 1870 3408 1876 3409
rect 1870 3404 1871 3408
rect 1875 3404 1876 3408
rect 1870 3403 1876 3404
rect 286 3399 292 3400
rect 286 3395 287 3399
rect 291 3395 292 3399
rect 286 3394 292 3395
rect 346 3399 352 3400
rect 346 3395 347 3399
rect 351 3395 352 3399
rect 346 3394 352 3395
rect 506 3399 512 3400
rect 506 3395 507 3399
rect 511 3395 512 3399
rect 506 3394 512 3395
rect 674 3399 680 3400
rect 674 3395 675 3399
rect 679 3395 680 3399
rect 674 3394 680 3395
rect 1010 3399 1016 3400
rect 1010 3395 1011 3399
rect 1015 3395 1016 3399
rect 1010 3394 1016 3395
rect 1170 3399 1176 3400
rect 1170 3395 1171 3399
rect 1175 3395 1176 3399
rect 1170 3394 1176 3395
rect 1350 3399 1356 3400
rect 1350 3395 1351 3399
rect 1355 3395 1356 3399
rect 1350 3394 1356 3395
rect 1466 3399 1472 3400
rect 1466 3395 1467 3399
rect 1471 3395 1472 3399
rect 1466 3394 1472 3395
rect 1610 3399 1616 3400
rect 1610 3395 1611 3399
rect 1615 3395 1616 3399
rect 1610 3394 1616 3395
rect 1734 3399 1740 3400
rect 1734 3395 1735 3399
rect 1739 3395 1740 3399
rect 1734 3394 1740 3395
rect 110 3391 116 3392
rect 110 3387 111 3391
rect 115 3387 116 3391
rect 110 3386 116 3387
rect 142 3388 148 3389
rect 112 3367 114 3386
rect 142 3384 143 3388
rect 147 3384 148 3388
rect 142 3383 148 3384
rect 286 3388 292 3389
rect 286 3384 287 3388
rect 291 3384 292 3388
rect 286 3383 292 3384
rect 446 3388 452 3389
rect 446 3384 447 3388
rect 451 3384 452 3388
rect 446 3383 452 3384
rect 614 3388 620 3389
rect 614 3384 615 3388
rect 619 3384 620 3388
rect 614 3383 620 3384
rect 782 3388 788 3389
rect 782 3384 783 3388
rect 787 3384 788 3388
rect 782 3383 788 3384
rect 950 3388 956 3389
rect 950 3384 951 3388
rect 955 3384 956 3388
rect 950 3383 956 3384
rect 1110 3388 1116 3389
rect 1110 3384 1111 3388
rect 1115 3384 1116 3388
rect 1110 3383 1116 3384
rect 1262 3388 1268 3389
rect 1262 3384 1263 3388
rect 1267 3384 1268 3388
rect 1262 3383 1268 3384
rect 1406 3388 1412 3389
rect 1406 3384 1407 3388
rect 1411 3384 1412 3388
rect 1406 3383 1412 3384
rect 1550 3388 1556 3389
rect 1550 3384 1551 3388
rect 1555 3384 1556 3388
rect 1550 3383 1556 3384
rect 1702 3388 1708 3389
rect 1702 3384 1703 3388
rect 1707 3384 1708 3388
rect 1702 3383 1708 3384
rect 144 3367 146 3383
rect 288 3367 290 3383
rect 448 3367 450 3383
rect 616 3367 618 3383
rect 678 3371 684 3372
rect 678 3367 679 3371
rect 683 3367 684 3371
rect 784 3367 786 3383
rect 952 3367 954 3383
rect 1112 3367 1114 3383
rect 1264 3367 1266 3383
rect 1408 3367 1410 3383
rect 1552 3367 1554 3383
rect 1704 3367 1706 3383
rect 111 3366 115 3367
rect 111 3361 115 3362
rect 143 3366 147 3367
rect 143 3361 147 3362
rect 207 3366 211 3367
rect 207 3361 211 3362
rect 287 3366 291 3367
rect 287 3361 291 3362
rect 335 3366 339 3367
rect 335 3361 339 3362
rect 447 3366 451 3367
rect 447 3361 451 3362
rect 471 3366 475 3367
rect 471 3361 475 3362
rect 615 3366 619 3367
rect 615 3361 619 3362
rect 623 3366 627 3367
rect 678 3366 684 3367
rect 783 3366 787 3367
rect 623 3361 627 3362
rect 112 3342 114 3361
rect 208 3345 210 3361
rect 336 3345 338 3361
rect 472 3345 474 3361
rect 624 3345 626 3361
rect 206 3344 212 3345
rect 110 3341 116 3342
rect 110 3337 111 3341
rect 115 3337 116 3341
rect 206 3340 207 3344
rect 211 3340 212 3344
rect 206 3339 212 3340
rect 334 3344 340 3345
rect 334 3340 335 3344
rect 339 3340 340 3344
rect 334 3339 340 3340
rect 470 3344 476 3345
rect 470 3340 471 3344
rect 475 3340 476 3344
rect 470 3339 476 3340
rect 622 3344 628 3345
rect 622 3340 623 3344
rect 627 3340 628 3344
rect 622 3339 628 3340
rect 110 3336 116 3337
rect 278 3335 284 3336
rect 278 3331 279 3335
rect 283 3331 284 3335
rect 278 3330 284 3331
rect 410 3335 416 3336
rect 410 3331 411 3335
rect 415 3331 416 3335
rect 410 3330 416 3331
rect 110 3324 116 3325
rect 110 3320 111 3324
rect 115 3320 116 3324
rect 110 3319 116 3320
rect 112 3287 114 3319
rect 214 3306 220 3307
rect 214 3302 215 3306
rect 219 3302 220 3306
rect 214 3301 220 3302
rect 216 3287 218 3301
rect 223 3300 227 3301
rect 280 3296 282 3330
rect 394 3327 400 3328
rect 394 3323 395 3327
rect 399 3323 400 3327
rect 394 3322 400 3323
rect 342 3306 348 3307
rect 342 3302 343 3306
rect 347 3302 348 3306
rect 342 3301 348 3302
rect 222 3295 228 3296
rect 222 3291 223 3295
rect 227 3291 228 3295
rect 222 3290 228 3291
rect 278 3295 284 3296
rect 278 3291 279 3295
rect 283 3291 284 3295
rect 278 3290 284 3291
rect 344 3287 346 3301
rect 111 3286 115 3287
rect 111 3281 115 3282
rect 215 3286 219 3287
rect 215 3281 219 3282
rect 343 3286 347 3287
rect 343 3281 347 3282
rect 351 3286 355 3287
rect 351 3281 355 3282
rect 112 3253 114 3281
rect 352 3271 354 3281
rect 396 3280 398 3322
rect 412 3296 414 3330
rect 478 3306 484 3307
rect 478 3302 479 3306
rect 483 3302 484 3306
rect 478 3301 484 3302
rect 630 3306 636 3307
rect 630 3302 631 3306
rect 635 3302 636 3306
rect 630 3301 636 3302
rect 680 3301 682 3366
rect 783 3361 787 3362
rect 943 3366 947 3367
rect 943 3361 947 3362
rect 951 3366 955 3367
rect 951 3361 955 3362
rect 1103 3366 1107 3367
rect 1103 3361 1107 3362
rect 1111 3366 1115 3367
rect 1111 3361 1115 3362
rect 1263 3366 1267 3367
rect 1263 3361 1267 3362
rect 1407 3366 1411 3367
rect 1407 3361 1411 3362
rect 1423 3366 1427 3367
rect 1423 3361 1427 3362
rect 1551 3366 1555 3367
rect 1551 3361 1555 3362
rect 1583 3366 1587 3367
rect 1583 3361 1587 3362
rect 1703 3366 1707 3367
rect 1703 3361 1707 3362
rect 784 3345 786 3361
rect 944 3345 946 3361
rect 1104 3345 1106 3361
rect 1264 3345 1266 3361
rect 1424 3345 1426 3361
rect 1584 3345 1586 3361
rect 782 3344 788 3345
rect 782 3340 783 3344
rect 787 3340 788 3344
rect 782 3339 788 3340
rect 942 3344 948 3345
rect 942 3340 943 3344
rect 947 3340 948 3344
rect 942 3339 948 3340
rect 1102 3344 1108 3345
rect 1102 3340 1103 3344
rect 1107 3340 1108 3344
rect 1102 3339 1108 3340
rect 1262 3344 1268 3345
rect 1262 3340 1263 3344
rect 1267 3340 1268 3344
rect 1262 3339 1268 3340
rect 1422 3344 1428 3345
rect 1422 3340 1423 3344
rect 1427 3340 1428 3344
rect 1422 3339 1428 3340
rect 1582 3344 1588 3345
rect 1582 3340 1583 3344
rect 1587 3340 1588 3344
rect 1582 3339 1588 3340
rect 706 3335 712 3336
rect 706 3331 707 3335
rect 711 3331 712 3335
rect 706 3330 712 3331
rect 1010 3335 1016 3336
rect 1010 3331 1011 3335
rect 1015 3331 1016 3335
rect 1010 3330 1016 3331
rect 1170 3335 1176 3336
rect 1170 3331 1171 3335
rect 1175 3331 1176 3335
rect 1170 3330 1176 3331
rect 1650 3335 1656 3336
rect 1650 3331 1651 3335
rect 1655 3331 1656 3335
rect 1650 3330 1656 3331
rect 410 3295 416 3296
rect 410 3291 411 3295
rect 415 3291 416 3295
rect 410 3290 416 3291
rect 480 3287 482 3301
rect 632 3287 634 3301
rect 679 3300 683 3301
rect 708 3296 710 3330
rect 790 3306 796 3307
rect 790 3302 791 3306
rect 795 3302 796 3306
rect 790 3301 796 3302
rect 950 3306 956 3307
rect 950 3302 951 3306
rect 955 3302 956 3306
rect 950 3301 956 3302
rect 679 3295 683 3296
rect 706 3295 712 3296
rect 706 3291 707 3295
rect 711 3291 712 3295
rect 706 3290 712 3291
rect 792 3287 794 3301
rect 952 3287 954 3301
rect 1012 3296 1014 3330
rect 1110 3306 1116 3307
rect 1110 3302 1111 3306
rect 1115 3302 1116 3306
rect 1110 3301 1116 3302
rect 1010 3295 1016 3296
rect 1010 3291 1011 3295
rect 1015 3291 1016 3295
rect 1010 3290 1016 3291
rect 1112 3287 1114 3301
rect 1172 3296 1174 3330
rect 1270 3306 1276 3307
rect 1270 3302 1271 3306
rect 1275 3302 1276 3306
rect 1270 3301 1276 3302
rect 1430 3306 1436 3307
rect 1430 3302 1431 3306
rect 1435 3302 1436 3306
rect 1430 3301 1436 3302
rect 1590 3306 1596 3307
rect 1590 3302 1591 3306
rect 1595 3302 1596 3306
rect 1590 3301 1596 3302
rect 1170 3295 1176 3296
rect 1170 3291 1171 3295
rect 1175 3291 1176 3295
rect 1170 3290 1176 3291
rect 1262 3295 1268 3296
rect 1262 3291 1263 3295
rect 1267 3291 1268 3295
rect 1262 3290 1268 3291
rect 455 3286 459 3287
rect 455 3281 459 3282
rect 479 3286 483 3287
rect 479 3281 483 3282
rect 575 3286 579 3287
rect 575 3281 579 3282
rect 631 3286 635 3287
rect 631 3281 635 3282
rect 703 3286 707 3287
rect 703 3281 707 3282
rect 791 3286 795 3287
rect 791 3281 795 3282
rect 839 3286 843 3287
rect 839 3281 843 3282
rect 951 3286 955 3287
rect 951 3281 955 3282
rect 983 3286 987 3287
rect 983 3281 987 3282
rect 1111 3286 1115 3287
rect 1111 3281 1115 3282
rect 1119 3286 1123 3287
rect 1119 3281 1123 3282
rect 1255 3286 1259 3287
rect 1255 3281 1259 3282
rect 394 3279 400 3280
rect 394 3275 395 3279
rect 399 3275 400 3279
rect 394 3274 400 3275
rect 402 3279 408 3280
rect 402 3275 403 3279
rect 407 3275 408 3279
rect 402 3274 408 3275
rect 350 3270 356 3271
rect 350 3266 351 3270
rect 355 3266 356 3270
rect 350 3265 356 3266
rect 110 3252 116 3253
rect 110 3248 111 3252
rect 115 3248 116 3252
rect 110 3247 116 3248
rect 404 3244 406 3274
rect 456 3271 458 3281
rect 506 3279 512 3280
rect 506 3275 507 3279
rect 511 3275 512 3279
rect 506 3274 512 3275
rect 454 3270 460 3271
rect 454 3266 455 3270
rect 459 3266 460 3270
rect 454 3265 460 3266
rect 508 3244 510 3274
rect 576 3271 578 3281
rect 704 3271 706 3281
rect 754 3279 760 3280
rect 754 3275 755 3279
rect 759 3275 760 3279
rect 754 3274 760 3275
rect 574 3270 580 3271
rect 574 3266 575 3270
rect 579 3266 580 3270
rect 574 3265 580 3266
rect 702 3270 708 3271
rect 702 3266 703 3270
rect 707 3266 708 3270
rect 702 3265 708 3266
rect 756 3244 758 3274
rect 840 3271 842 3281
rect 984 3271 986 3281
rect 990 3279 996 3280
rect 990 3275 991 3279
rect 995 3275 996 3279
rect 990 3274 996 3275
rect 1034 3279 1040 3280
rect 1034 3275 1035 3279
rect 1039 3275 1040 3279
rect 1034 3274 1040 3275
rect 838 3270 844 3271
rect 838 3266 839 3270
rect 843 3266 844 3270
rect 838 3265 844 3266
rect 982 3270 988 3271
rect 982 3266 983 3270
rect 987 3266 988 3270
rect 982 3265 988 3266
rect 402 3243 408 3244
rect 402 3239 403 3243
rect 407 3239 408 3243
rect 402 3238 408 3239
rect 506 3243 512 3244
rect 506 3239 507 3243
rect 511 3239 512 3243
rect 506 3238 512 3239
rect 754 3243 760 3244
rect 754 3239 755 3243
rect 759 3239 760 3243
rect 754 3238 760 3239
rect 110 3235 116 3236
rect 110 3231 111 3235
rect 115 3231 116 3235
rect 110 3230 116 3231
rect 342 3232 348 3233
rect 112 3211 114 3230
rect 342 3228 343 3232
rect 347 3228 348 3232
rect 342 3227 348 3228
rect 446 3232 452 3233
rect 446 3228 447 3232
rect 451 3228 452 3232
rect 446 3227 452 3228
rect 566 3232 572 3233
rect 566 3228 567 3232
rect 571 3228 572 3232
rect 566 3227 572 3228
rect 694 3232 700 3233
rect 694 3228 695 3232
rect 699 3228 700 3232
rect 694 3227 700 3228
rect 830 3232 836 3233
rect 830 3228 831 3232
rect 835 3228 836 3232
rect 830 3227 836 3228
rect 974 3232 980 3233
rect 974 3228 975 3232
rect 979 3228 980 3232
rect 974 3227 980 3228
rect 344 3211 346 3227
rect 448 3211 450 3227
rect 502 3215 508 3216
rect 502 3211 503 3215
rect 507 3211 508 3215
rect 568 3211 570 3227
rect 696 3211 698 3227
rect 832 3211 834 3227
rect 976 3211 978 3227
rect 111 3210 115 3211
rect 111 3205 115 3206
rect 343 3210 347 3211
rect 343 3205 347 3206
rect 447 3210 451 3211
rect 447 3205 451 3206
rect 487 3210 491 3211
rect 502 3210 508 3211
rect 567 3210 571 3211
rect 487 3205 491 3206
rect 112 3186 114 3205
rect 488 3189 490 3205
rect 486 3188 492 3189
rect 110 3185 116 3186
rect 110 3181 111 3185
rect 115 3181 116 3185
rect 486 3184 487 3188
rect 491 3184 492 3188
rect 486 3183 492 3184
rect 110 3180 116 3181
rect 110 3168 116 3169
rect 110 3164 111 3168
rect 115 3164 116 3168
rect 110 3163 116 3164
rect 112 3131 114 3163
rect 494 3150 500 3151
rect 494 3146 495 3150
rect 499 3146 500 3150
rect 494 3145 500 3146
rect 496 3131 498 3145
rect 504 3140 506 3210
rect 567 3205 571 3206
rect 575 3210 579 3211
rect 575 3205 579 3206
rect 663 3210 667 3211
rect 663 3205 667 3206
rect 695 3210 699 3211
rect 695 3205 699 3206
rect 767 3210 771 3211
rect 767 3205 771 3206
rect 831 3210 835 3211
rect 831 3205 835 3206
rect 887 3210 891 3211
rect 887 3205 891 3206
rect 975 3210 979 3211
rect 975 3205 979 3206
rect 576 3189 578 3205
rect 664 3189 666 3205
rect 768 3189 770 3205
rect 888 3189 890 3205
rect 574 3188 580 3189
rect 574 3184 575 3188
rect 579 3184 580 3188
rect 574 3183 580 3184
rect 662 3188 668 3189
rect 662 3184 663 3188
rect 667 3184 668 3188
rect 662 3183 668 3184
rect 766 3188 772 3189
rect 766 3184 767 3188
rect 771 3184 772 3188
rect 766 3183 772 3184
rect 886 3188 892 3189
rect 886 3184 887 3188
rect 891 3184 892 3188
rect 886 3183 892 3184
rect 992 3180 994 3274
rect 1036 3244 1038 3274
rect 1120 3271 1122 3281
rect 1170 3279 1176 3280
rect 1170 3275 1171 3279
rect 1175 3275 1176 3279
rect 1170 3274 1176 3275
rect 1118 3270 1124 3271
rect 1118 3266 1119 3270
rect 1123 3266 1124 3270
rect 1118 3265 1124 3266
rect 1172 3244 1174 3274
rect 1256 3271 1258 3281
rect 1254 3270 1260 3271
rect 1254 3266 1255 3270
rect 1259 3266 1260 3270
rect 1254 3265 1260 3266
rect 1264 3244 1266 3290
rect 1272 3287 1274 3301
rect 1432 3287 1434 3301
rect 1592 3287 1594 3301
rect 1652 3296 1654 3330
rect 1736 3296 1738 3394
rect 1830 3391 1836 3392
rect 1830 3387 1831 3391
rect 1835 3387 1836 3391
rect 1830 3386 1836 3387
rect 1870 3391 1876 3392
rect 1870 3387 1871 3391
rect 1875 3387 1876 3391
rect 1870 3386 1876 3387
rect 2102 3388 2108 3389
rect 1832 3367 1834 3386
rect 1743 3366 1747 3367
rect 1743 3361 1747 3362
rect 1831 3366 1835 3367
rect 1872 3363 1874 3386
rect 2102 3384 2103 3388
rect 2107 3384 2108 3388
rect 2102 3383 2108 3384
rect 2104 3363 2106 3383
rect 2156 3372 2158 3430
rect 2164 3400 2166 3430
rect 2200 3427 2202 3437
rect 2198 3426 2204 3427
rect 2198 3422 2199 3426
rect 2203 3422 2204 3426
rect 2198 3421 2204 3422
rect 2252 3400 2254 3450
rect 2272 3443 2274 3461
rect 2376 3443 2378 3461
rect 2384 3456 2386 3526
rect 2471 3521 2475 3522
rect 2487 3526 2491 3527
rect 2487 3521 2491 3522
rect 2583 3526 2587 3527
rect 2583 3521 2587 3522
rect 2615 3526 2619 3527
rect 2615 3521 2619 3522
rect 2695 3526 2699 3527
rect 2695 3521 2699 3522
rect 2743 3526 2747 3527
rect 2743 3521 2747 3522
rect 2807 3526 2811 3527
rect 2807 3521 2811 3522
rect 2488 3505 2490 3521
rect 2616 3505 2618 3521
rect 2744 3505 2746 3521
rect 2486 3504 2492 3505
rect 2486 3500 2487 3504
rect 2491 3500 2492 3504
rect 2486 3499 2492 3500
rect 2614 3504 2620 3505
rect 2614 3500 2615 3504
rect 2619 3500 2620 3504
rect 2614 3499 2620 3500
rect 2742 3504 2748 3505
rect 2742 3500 2743 3504
rect 2747 3500 2748 3504
rect 2742 3499 2748 3500
rect 2828 3496 2830 3598
rect 2919 3597 2923 3598
rect 3015 3602 3019 3603
rect 3015 3597 3019 3598
rect 3111 3602 3115 3603
rect 3111 3597 3115 3598
rect 3207 3602 3211 3603
rect 3207 3597 3211 3598
rect 3303 3602 3307 3603
rect 3303 3597 3307 3598
rect 3399 3602 3403 3603
rect 3399 3597 3403 3598
rect 3591 3602 3595 3603
rect 3591 3597 3595 3598
rect 2866 3595 2872 3596
rect 2866 3591 2867 3595
rect 2871 3591 2872 3595
rect 2866 3590 2872 3591
rect 2868 3560 2870 3590
rect 2920 3587 2922 3597
rect 2970 3595 2976 3596
rect 2970 3591 2971 3595
rect 2975 3591 2976 3595
rect 2970 3590 2976 3591
rect 2918 3586 2924 3587
rect 2918 3582 2919 3586
rect 2923 3582 2924 3586
rect 2918 3581 2924 3582
rect 2972 3560 2974 3590
rect 3016 3587 3018 3597
rect 3066 3595 3072 3596
rect 3066 3591 3067 3595
rect 3071 3591 3072 3595
rect 3066 3590 3072 3591
rect 3014 3586 3020 3587
rect 3014 3582 3015 3586
rect 3019 3582 3020 3586
rect 3014 3581 3020 3582
rect 3068 3560 3070 3590
rect 3112 3587 3114 3597
rect 3162 3595 3168 3596
rect 3162 3591 3163 3595
rect 3167 3591 3168 3595
rect 3162 3590 3168 3591
rect 3110 3586 3116 3587
rect 3110 3582 3111 3586
rect 3115 3582 3116 3586
rect 3110 3581 3116 3582
rect 3164 3560 3166 3590
rect 3208 3587 3210 3597
rect 3258 3595 3264 3596
rect 3258 3591 3259 3595
rect 3263 3591 3264 3595
rect 3258 3590 3264 3591
rect 3206 3586 3212 3587
rect 3206 3582 3207 3586
rect 3211 3582 3212 3586
rect 3206 3581 3212 3582
rect 3260 3560 3262 3590
rect 3304 3587 3306 3597
rect 3354 3595 3360 3596
rect 3354 3591 3355 3595
rect 3359 3591 3360 3595
rect 3354 3590 3360 3591
rect 3302 3586 3308 3587
rect 3302 3582 3303 3586
rect 3307 3582 3308 3586
rect 3302 3581 3308 3582
rect 3356 3560 3358 3590
rect 3400 3587 3402 3597
rect 3398 3586 3404 3587
rect 3398 3582 3399 3586
rect 3403 3582 3404 3586
rect 3398 3581 3404 3582
rect 3592 3569 3594 3597
rect 3590 3568 3596 3569
rect 3590 3564 3591 3568
rect 3595 3564 3596 3568
rect 3590 3563 3596 3564
rect 2866 3559 2872 3560
rect 2866 3555 2867 3559
rect 2871 3555 2872 3559
rect 2866 3554 2872 3555
rect 2970 3559 2976 3560
rect 2970 3555 2971 3559
rect 2975 3555 2976 3559
rect 2970 3554 2976 3555
rect 3066 3559 3072 3560
rect 3066 3555 3067 3559
rect 3071 3555 3072 3559
rect 3066 3554 3072 3555
rect 3162 3559 3168 3560
rect 3162 3555 3163 3559
rect 3167 3555 3168 3559
rect 3162 3554 3168 3555
rect 3258 3559 3264 3560
rect 3258 3555 3259 3559
rect 3263 3555 3264 3559
rect 3258 3554 3264 3555
rect 3354 3559 3360 3560
rect 3354 3555 3355 3559
rect 3359 3555 3360 3559
rect 3354 3554 3360 3555
rect 3590 3551 3596 3552
rect 2910 3548 2916 3549
rect 2910 3544 2911 3548
rect 2915 3544 2916 3548
rect 2910 3543 2916 3544
rect 3006 3548 3012 3549
rect 3006 3544 3007 3548
rect 3011 3544 3012 3548
rect 3006 3543 3012 3544
rect 3102 3548 3108 3549
rect 3102 3544 3103 3548
rect 3107 3544 3108 3548
rect 3102 3543 3108 3544
rect 3198 3548 3204 3549
rect 3198 3544 3199 3548
rect 3203 3544 3204 3548
rect 3198 3543 3204 3544
rect 3294 3548 3300 3549
rect 3294 3544 3295 3548
rect 3299 3544 3300 3548
rect 3294 3543 3300 3544
rect 3390 3548 3396 3549
rect 3390 3544 3391 3548
rect 3395 3544 3396 3548
rect 3590 3547 3591 3551
rect 3595 3547 3596 3551
rect 3590 3546 3596 3547
rect 3390 3543 3396 3544
rect 2912 3527 2914 3543
rect 3008 3527 3010 3543
rect 3104 3527 3106 3543
rect 3134 3531 3140 3532
rect 3134 3527 3135 3531
rect 3139 3527 3140 3531
rect 3200 3527 3202 3543
rect 3296 3527 3298 3543
rect 3392 3527 3394 3543
rect 3592 3527 3594 3546
rect 2871 3526 2875 3527
rect 2871 3521 2875 3522
rect 2911 3526 2915 3527
rect 2911 3521 2915 3522
rect 2991 3526 2995 3527
rect 2991 3521 2995 3522
rect 3007 3526 3011 3527
rect 3007 3521 3011 3522
rect 3103 3526 3107 3527
rect 3103 3521 3107 3522
rect 3119 3526 3123 3527
rect 3134 3526 3140 3527
rect 3199 3526 3203 3527
rect 3119 3521 3123 3522
rect 2872 3505 2874 3521
rect 2992 3505 2994 3521
rect 3120 3505 3122 3521
rect 2870 3504 2876 3505
rect 2870 3500 2871 3504
rect 2875 3500 2876 3504
rect 2870 3499 2876 3500
rect 2990 3504 2996 3505
rect 2990 3500 2991 3504
rect 2995 3500 2996 3504
rect 2990 3499 2996 3500
rect 3118 3504 3124 3505
rect 3118 3500 3119 3504
rect 3123 3500 3124 3504
rect 3118 3499 3124 3500
rect 2434 3495 2440 3496
rect 2434 3491 2435 3495
rect 2439 3491 2440 3495
rect 2434 3490 2440 3491
rect 2558 3495 2564 3496
rect 2558 3491 2559 3495
rect 2563 3491 2564 3495
rect 2558 3490 2564 3491
rect 2686 3495 2692 3496
rect 2686 3491 2687 3495
rect 2691 3491 2692 3495
rect 2686 3490 2692 3491
rect 2826 3495 2832 3496
rect 2826 3491 2827 3495
rect 2831 3491 2832 3495
rect 2826 3490 2832 3491
rect 2938 3495 2944 3496
rect 2938 3491 2939 3495
rect 2943 3491 2944 3495
rect 2938 3490 2944 3491
rect 2436 3456 2438 3490
rect 2494 3466 2500 3467
rect 2494 3462 2495 3466
rect 2499 3462 2500 3466
rect 2494 3461 2500 3462
rect 2382 3455 2388 3456
rect 2382 3451 2383 3455
rect 2387 3451 2388 3455
rect 2382 3450 2388 3451
rect 2434 3455 2440 3456
rect 2434 3451 2435 3455
rect 2439 3451 2440 3455
rect 2434 3450 2440 3451
rect 2496 3443 2498 3461
rect 2560 3456 2562 3490
rect 2622 3466 2628 3467
rect 2622 3462 2623 3466
rect 2627 3462 2628 3466
rect 2622 3461 2628 3462
rect 2558 3455 2564 3456
rect 2558 3451 2559 3455
rect 2563 3451 2564 3455
rect 2558 3450 2564 3451
rect 2624 3443 2626 3461
rect 2688 3456 2690 3490
rect 2750 3466 2756 3467
rect 2750 3462 2751 3466
rect 2755 3462 2756 3466
rect 2750 3461 2756 3462
rect 2878 3466 2884 3467
rect 2878 3462 2879 3466
rect 2883 3462 2884 3466
rect 2878 3461 2884 3462
rect 2686 3455 2692 3456
rect 2686 3451 2687 3455
rect 2691 3451 2692 3455
rect 2686 3450 2692 3451
rect 2752 3443 2754 3461
rect 2880 3443 2882 3461
rect 2940 3456 2942 3490
rect 2998 3466 3004 3467
rect 2998 3462 2999 3466
rect 3003 3462 3004 3466
rect 2998 3461 3004 3462
rect 3126 3466 3132 3467
rect 3126 3462 3127 3466
rect 3131 3462 3132 3466
rect 3126 3461 3132 3462
rect 2938 3455 2944 3456
rect 2938 3451 2939 3455
rect 2943 3451 2944 3455
rect 2938 3450 2944 3451
rect 2990 3455 2996 3456
rect 2990 3451 2991 3455
rect 2995 3451 2996 3455
rect 2990 3450 2996 3451
rect 2271 3442 2275 3443
rect 2271 3437 2275 3438
rect 2303 3442 2307 3443
rect 2303 3437 2307 3438
rect 2375 3442 2379 3443
rect 2375 3437 2379 3438
rect 2415 3442 2419 3443
rect 2415 3437 2419 3438
rect 2495 3442 2499 3443
rect 2495 3437 2499 3438
rect 2543 3442 2547 3443
rect 2543 3437 2547 3438
rect 2623 3442 2627 3443
rect 2623 3437 2627 3438
rect 2679 3442 2683 3443
rect 2679 3437 2683 3438
rect 2751 3442 2755 3443
rect 2751 3437 2755 3438
rect 2815 3442 2819 3443
rect 2815 3437 2819 3438
rect 2879 3442 2883 3443
rect 2879 3437 2883 3438
rect 2959 3442 2963 3443
rect 2959 3437 2963 3438
rect 2294 3435 2300 3436
rect 2294 3431 2295 3435
rect 2299 3431 2300 3435
rect 2294 3430 2300 3431
rect 2296 3404 2298 3430
rect 2304 3427 2306 3437
rect 2416 3427 2418 3437
rect 2422 3435 2428 3436
rect 2422 3431 2423 3435
rect 2427 3431 2428 3435
rect 2422 3430 2428 3431
rect 2302 3426 2308 3427
rect 2302 3422 2303 3426
rect 2307 3422 2308 3426
rect 2302 3421 2308 3422
rect 2414 3426 2420 3427
rect 2414 3422 2415 3426
rect 2419 3422 2420 3426
rect 2414 3421 2420 3422
rect 2294 3403 2300 3404
rect 2162 3399 2168 3400
rect 2162 3395 2163 3399
rect 2167 3395 2168 3399
rect 2162 3394 2168 3395
rect 2250 3399 2256 3400
rect 2250 3395 2251 3399
rect 2255 3395 2256 3399
rect 2294 3399 2295 3403
rect 2299 3399 2300 3403
rect 2294 3398 2300 3399
rect 2250 3394 2256 3395
rect 2190 3388 2196 3389
rect 2190 3384 2191 3388
rect 2195 3384 2196 3388
rect 2190 3383 2196 3384
rect 2294 3388 2300 3389
rect 2294 3384 2295 3388
rect 2299 3384 2300 3388
rect 2294 3383 2300 3384
rect 2406 3388 2412 3389
rect 2406 3384 2407 3388
rect 2411 3384 2412 3388
rect 2406 3383 2412 3384
rect 2154 3371 2160 3372
rect 2154 3367 2155 3371
rect 2159 3367 2160 3371
rect 2154 3366 2160 3367
rect 2192 3363 2194 3383
rect 2296 3363 2298 3383
rect 2408 3363 2410 3383
rect 1831 3361 1835 3362
rect 1871 3362 1875 3363
rect 1744 3345 1746 3361
rect 1742 3344 1748 3345
rect 1742 3340 1743 3344
rect 1747 3340 1748 3344
rect 1832 3342 1834 3361
rect 1871 3357 1875 3358
rect 2103 3362 2107 3363
rect 2103 3357 2107 3358
rect 2127 3362 2131 3363
rect 2127 3357 2131 3358
rect 2191 3362 2195 3363
rect 2191 3357 2195 3358
rect 2223 3362 2227 3363
rect 2223 3357 2227 3358
rect 2295 3362 2299 3363
rect 2295 3357 2299 3358
rect 2335 3362 2339 3363
rect 2335 3357 2339 3358
rect 2407 3362 2411 3363
rect 2407 3357 2411 3358
rect 1742 3339 1748 3340
rect 1830 3341 1836 3342
rect 1830 3337 1831 3341
rect 1835 3337 1836 3341
rect 1872 3338 1874 3357
rect 2128 3341 2130 3357
rect 2224 3341 2226 3357
rect 2336 3341 2338 3357
rect 2126 3340 2132 3341
rect 1830 3336 1836 3337
rect 1870 3337 1876 3338
rect 1870 3333 1871 3337
rect 1875 3333 1876 3337
rect 2126 3336 2127 3340
rect 2131 3336 2132 3340
rect 2126 3335 2132 3336
rect 2222 3340 2228 3341
rect 2222 3336 2223 3340
rect 2227 3336 2228 3340
rect 2222 3335 2228 3336
rect 2334 3340 2340 3341
rect 2334 3336 2335 3340
rect 2339 3336 2340 3340
rect 2334 3335 2340 3336
rect 1870 3332 1876 3333
rect 2424 3332 2426 3430
rect 2544 3427 2546 3437
rect 2602 3435 2608 3436
rect 2602 3431 2603 3435
rect 2607 3431 2608 3435
rect 2602 3430 2608 3431
rect 2542 3426 2548 3427
rect 2542 3422 2543 3426
rect 2547 3422 2548 3426
rect 2542 3421 2548 3422
rect 2604 3400 2606 3430
rect 2680 3427 2682 3437
rect 2738 3435 2744 3436
rect 2738 3431 2739 3435
rect 2743 3431 2744 3435
rect 2738 3430 2744 3431
rect 2678 3426 2684 3427
rect 2678 3422 2679 3426
rect 2683 3422 2684 3426
rect 2678 3421 2684 3422
rect 2740 3400 2742 3430
rect 2816 3427 2818 3437
rect 2960 3427 2962 3437
rect 2814 3426 2820 3427
rect 2814 3422 2815 3426
rect 2819 3422 2820 3426
rect 2814 3421 2820 3422
rect 2958 3426 2964 3427
rect 2958 3422 2959 3426
rect 2963 3422 2964 3426
rect 2958 3421 2964 3422
rect 2992 3400 2994 3450
rect 3000 3443 3002 3461
rect 3128 3443 3130 3461
rect 3136 3456 3138 3526
rect 3199 3521 3203 3522
rect 3247 3526 3251 3527
rect 3247 3521 3251 3522
rect 3295 3526 3299 3527
rect 3295 3521 3299 3522
rect 3375 3526 3379 3527
rect 3375 3521 3379 3522
rect 3391 3526 3395 3527
rect 3391 3521 3395 3522
rect 3591 3526 3595 3527
rect 3591 3521 3595 3522
rect 3248 3505 3250 3521
rect 3376 3505 3378 3521
rect 3246 3504 3252 3505
rect 3246 3500 3247 3504
rect 3251 3500 3252 3504
rect 3246 3499 3252 3500
rect 3374 3504 3380 3505
rect 3374 3500 3375 3504
rect 3379 3500 3380 3504
rect 3592 3502 3594 3521
rect 3374 3499 3380 3500
rect 3590 3501 3596 3502
rect 3590 3497 3591 3501
rect 3595 3497 3596 3501
rect 3590 3496 3596 3497
rect 3318 3495 3324 3496
rect 3318 3491 3319 3495
rect 3323 3491 3324 3495
rect 3318 3490 3324 3491
rect 3254 3466 3260 3467
rect 3254 3462 3255 3466
rect 3259 3462 3260 3466
rect 3254 3461 3260 3462
rect 3134 3455 3140 3456
rect 3134 3451 3135 3455
rect 3139 3451 3140 3455
rect 3134 3450 3140 3451
rect 3256 3443 3258 3461
rect 3320 3456 3322 3490
rect 3434 3487 3440 3488
rect 3434 3483 3435 3487
rect 3439 3483 3440 3487
rect 3434 3482 3440 3483
rect 3590 3484 3596 3485
rect 3382 3466 3388 3467
rect 3382 3462 3383 3466
rect 3387 3462 3388 3466
rect 3382 3461 3388 3462
rect 3318 3455 3324 3456
rect 3318 3451 3319 3455
rect 3323 3451 3324 3455
rect 3318 3450 3324 3451
rect 3384 3443 3386 3461
rect 2999 3442 3003 3443
rect 2999 3437 3003 3438
rect 3111 3442 3115 3443
rect 3111 3437 3115 3438
rect 3127 3442 3131 3443
rect 3127 3437 3131 3438
rect 3255 3442 3259 3443
rect 3255 3437 3259 3438
rect 3263 3442 3267 3443
rect 3263 3437 3267 3438
rect 3383 3442 3387 3443
rect 3383 3437 3387 3438
rect 3423 3442 3427 3443
rect 3423 3437 3427 3438
rect 3030 3435 3036 3436
rect 3030 3431 3031 3435
rect 3035 3431 3036 3435
rect 3030 3430 3036 3431
rect 3032 3400 3034 3430
rect 3112 3427 3114 3437
rect 3134 3435 3140 3436
rect 3134 3431 3135 3435
rect 3139 3431 3140 3435
rect 3134 3430 3140 3431
rect 3110 3426 3116 3427
rect 3110 3422 3111 3426
rect 3115 3422 3116 3426
rect 3110 3421 3116 3422
rect 2574 3399 2580 3400
rect 2574 3395 2575 3399
rect 2579 3395 2580 3399
rect 2574 3394 2580 3395
rect 2602 3399 2608 3400
rect 2602 3395 2603 3399
rect 2607 3395 2608 3399
rect 2602 3394 2608 3395
rect 2738 3399 2744 3400
rect 2738 3395 2739 3399
rect 2743 3395 2744 3399
rect 2738 3394 2744 3395
rect 2990 3399 2996 3400
rect 2990 3395 2991 3399
rect 2995 3395 2996 3399
rect 2990 3394 2996 3395
rect 3030 3399 3036 3400
rect 3030 3395 3031 3399
rect 3035 3395 3036 3399
rect 3030 3394 3036 3395
rect 2534 3388 2540 3389
rect 2534 3384 2535 3388
rect 2539 3384 2540 3388
rect 2534 3383 2540 3384
rect 2536 3363 2538 3383
rect 2455 3362 2459 3363
rect 2455 3357 2459 3358
rect 2535 3362 2539 3363
rect 2535 3357 2539 3358
rect 2456 3341 2458 3357
rect 2454 3340 2460 3341
rect 2454 3336 2455 3340
rect 2459 3336 2460 3340
rect 2454 3335 2460 3336
rect 2194 3331 2200 3332
rect 2194 3327 2195 3331
rect 2199 3327 2200 3331
rect 2194 3326 2200 3327
rect 2290 3331 2296 3332
rect 2290 3327 2291 3331
rect 2295 3327 2296 3331
rect 2290 3326 2296 3327
rect 2402 3331 2408 3332
rect 2402 3327 2403 3331
rect 2407 3327 2408 3331
rect 2402 3326 2408 3327
rect 2422 3331 2428 3332
rect 2422 3327 2423 3331
rect 2427 3327 2428 3331
rect 2422 3326 2428 3327
rect 1830 3324 1836 3325
rect 1830 3320 1831 3324
rect 1835 3320 1836 3324
rect 1830 3319 1836 3320
rect 1870 3320 1876 3321
rect 1750 3306 1756 3307
rect 1750 3302 1751 3306
rect 1755 3302 1756 3306
rect 1750 3301 1756 3302
rect 1650 3295 1656 3296
rect 1650 3291 1651 3295
rect 1655 3291 1656 3295
rect 1650 3290 1656 3291
rect 1734 3295 1740 3296
rect 1734 3291 1735 3295
rect 1739 3291 1740 3295
rect 1734 3290 1740 3291
rect 1752 3287 1754 3301
rect 1832 3287 1834 3319
rect 1870 3316 1871 3320
rect 1875 3316 1876 3320
rect 1870 3315 1876 3316
rect 1271 3286 1275 3287
rect 1271 3281 1275 3282
rect 1383 3286 1387 3287
rect 1383 3281 1387 3282
rect 1431 3286 1435 3287
rect 1431 3281 1435 3282
rect 1511 3286 1515 3287
rect 1511 3281 1515 3282
rect 1591 3286 1595 3287
rect 1591 3281 1595 3282
rect 1639 3286 1643 3287
rect 1639 3281 1643 3282
rect 1751 3286 1755 3287
rect 1751 3281 1755 3282
rect 1831 3286 1835 3287
rect 1831 3281 1835 3282
rect 1384 3271 1386 3281
rect 1512 3271 1514 3281
rect 1562 3279 1568 3280
rect 1562 3275 1563 3279
rect 1567 3275 1568 3279
rect 1562 3274 1568 3275
rect 1382 3270 1388 3271
rect 1382 3266 1383 3270
rect 1387 3266 1388 3270
rect 1382 3265 1388 3266
rect 1510 3270 1516 3271
rect 1510 3266 1511 3270
rect 1515 3266 1516 3270
rect 1510 3265 1516 3266
rect 1564 3244 1566 3274
rect 1640 3271 1642 3281
rect 1690 3279 1696 3280
rect 1690 3275 1691 3279
rect 1695 3275 1696 3279
rect 1690 3274 1696 3275
rect 1638 3270 1644 3271
rect 1638 3266 1639 3270
rect 1643 3266 1644 3270
rect 1638 3265 1644 3266
rect 1692 3244 1694 3274
rect 1752 3271 1754 3281
rect 1750 3270 1756 3271
rect 1750 3266 1751 3270
rect 1755 3266 1756 3270
rect 1750 3265 1756 3266
rect 1832 3253 1834 3281
rect 1872 3275 1874 3315
rect 2134 3302 2140 3303
rect 2134 3298 2135 3302
rect 2139 3298 2140 3302
rect 2134 3297 2140 3298
rect 2136 3275 2138 3297
rect 2196 3292 2198 3326
rect 2230 3302 2236 3303
rect 2230 3298 2231 3302
rect 2235 3298 2236 3302
rect 2230 3297 2236 3298
rect 2142 3291 2148 3292
rect 2142 3287 2143 3291
rect 2147 3287 2148 3291
rect 2142 3286 2148 3287
rect 2194 3291 2200 3292
rect 2194 3287 2195 3291
rect 2199 3287 2200 3291
rect 2194 3286 2200 3287
rect 1871 3274 1875 3275
rect 1871 3269 1875 3270
rect 2135 3274 2139 3275
rect 2135 3269 2139 3270
rect 1830 3252 1836 3253
rect 1830 3248 1831 3252
rect 1835 3248 1836 3252
rect 1830 3247 1836 3248
rect 1034 3243 1040 3244
rect 1034 3239 1035 3243
rect 1039 3239 1040 3243
rect 1034 3238 1040 3239
rect 1170 3243 1176 3244
rect 1170 3239 1171 3243
rect 1175 3239 1176 3243
rect 1170 3238 1176 3239
rect 1262 3243 1268 3244
rect 1262 3239 1263 3243
rect 1267 3239 1268 3243
rect 1262 3238 1268 3239
rect 1562 3243 1568 3244
rect 1562 3239 1563 3243
rect 1567 3239 1568 3243
rect 1562 3238 1568 3239
rect 1690 3243 1696 3244
rect 1690 3239 1691 3243
rect 1695 3239 1696 3243
rect 1872 3241 1874 3269
rect 2136 3259 2138 3269
rect 2134 3258 2140 3259
rect 2134 3254 2135 3258
rect 2139 3254 2140 3258
rect 2134 3253 2140 3254
rect 1690 3238 1696 3239
rect 1870 3240 1876 3241
rect 1870 3236 1871 3240
rect 1875 3236 1876 3240
rect 1830 3235 1836 3236
rect 1870 3235 1876 3236
rect 1110 3232 1116 3233
rect 1110 3228 1111 3232
rect 1115 3228 1116 3232
rect 1110 3227 1116 3228
rect 1246 3232 1252 3233
rect 1246 3228 1247 3232
rect 1251 3228 1252 3232
rect 1246 3227 1252 3228
rect 1374 3232 1380 3233
rect 1374 3228 1375 3232
rect 1379 3228 1380 3232
rect 1374 3227 1380 3228
rect 1502 3232 1508 3233
rect 1502 3228 1503 3232
rect 1507 3228 1508 3232
rect 1502 3227 1508 3228
rect 1630 3232 1636 3233
rect 1630 3228 1631 3232
rect 1635 3228 1636 3232
rect 1630 3227 1636 3228
rect 1742 3232 1748 3233
rect 1742 3228 1743 3232
rect 1747 3228 1748 3232
rect 1830 3231 1831 3235
rect 1835 3231 1836 3235
rect 2144 3232 2146 3286
rect 2232 3275 2234 3297
rect 2292 3292 2294 3326
rect 2342 3302 2348 3303
rect 2342 3298 2343 3302
rect 2347 3298 2348 3302
rect 2342 3297 2348 3298
rect 2290 3291 2296 3292
rect 2290 3287 2291 3291
rect 2295 3287 2296 3291
rect 2290 3286 2296 3287
rect 2344 3275 2346 3297
rect 2404 3292 2406 3326
rect 2462 3302 2468 3303
rect 2462 3298 2463 3302
rect 2467 3298 2468 3302
rect 2462 3297 2468 3298
rect 2402 3291 2408 3292
rect 2402 3287 2403 3291
rect 2407 3287 2408 3291
rect 2402 3286 2408 3287
rect 2422 3275 2428 3276
rect 2464 3275 2466 3297
rect 2576 3292 2578 3394
rect 2670 3388 2676 3389
rect 2670 3384 2671 3388
rect 2675 3384 2676 3388
rect 2670 3383 2676 3384
rect 2806 3388 2812 3389
rect 2806 3384 2807 3388
rect 2811 3384 2812 3388
rect 2806 3383 2812 3384
rect 2950 3388 2956 3389
rect 2950 3384 2951 3388
rect 2955 3384 2956 3388
rect 2950 3383 2956 3384
rect 3102 3388 3108 3389
rect 3102 3384 3103 3388
rect 3107 3384 3108 3388
rect 3102 3383 3108 3384
rect 2672 3363 2674 3383
rect 2808 3363 2810 3383
rect 2952 3363 2954 3383
rect 3104 3363 3106 3383
rect 2583 3362 2587 3363
rect 2583 3357 2587 3358
rect 2671 3362 2675 3363
rect 2671 3357 2675 3358
rect 2719 3362 2723 3363
rect 2719 3357 2723 3358
rect 2807 3362 2811 3363
rect 2807 3357 2811 3358
rect 2863 3362 2867 3363
rect 2863 3357 2867 3358
rect 2951 3362 2955 3363
rect 2951 3357 2955 3358
rect 3007 3362 3011 3363
rect 3007 3357 3011 3358
rect 3103 3362 3107 3363
rect 3103 3357 3107 3358
rect 2584 3341 2586 3357
rect 2720 3341 2722 3357
rect 2864 3341 2866 3357
rect 3008 3341 3010 3357
rect 2582 3340 2588 3341
rect 2582 3336 2583 3340
rect 2587 3336 2588 3340
rect 2582 3335 2588 3336
rect 2718 3340 2724 3341
rect 2718 3336 2719 3340
rect 2723 3336 2724 3340
rect 2718 3335 2724 3336
rect 2862 3340 2868 3341
rect 2862 3336 2863 3340
rect 2867 3336 2868 3340
rect 2862 3335 2868 3336
rect 3006 3340 3012 3341
rect 3006 3336 3007 3340
rect 3011 3336 3012 3340
rect 3006 3335 3012 3336
rect 3136 3332 3138 3430
rect 3264 3427 3266 3437
rect 3424 3427 3426 3437
rect 3436 3436 3438 3482
rect 3590 3480 3591 3484
rect 3595 3480 3596 3484
rect 3590 3479 3596 3480
rect 3592 3443 3594 3479
rect 3591 3442 3595 3443
rect 3591 3437 3595 3438
rect 3434 3435 3440 3436
rect 3434 3431 3435 3435
rect 3439 3431 3440 3435
rect 3434 3430 3440 3431
rect 3262 3426 3268 3427
rect 3262 3422 3263 3426
rect 3267 3422 3268 3426
rect 3262 3421 3268 3422
rect 3422 3426 3428 3427
rect 3422 3422 3423 3426
rect 3427 3422 3428 3426
rect 3422 3421 3428 3422
rect 3592 3409 3594 3437
rect 3590 3408 3596 3409
rect 3590 3404 3591 3408
rect 3595 3404 3596 3408
rect 3590 3403 3596 3404
rect 3302 3399 3308 3400
rect 3302 3395 3303 3399
rect 3307 3395 3308 3399
rect 3302 3394 3308 3395
rect 3254 3388 3260 3389
rect 3254 3384 3255 3388
rect 3259 3384 3260 3388
rect 3254 3383 3260 3384
rect 3256 3363 3258 3383
rect 3159 3362 3163 3363
rect 3159 3357 3163 3358
rect 3255 3362 3259 3363
rect 3255 3357 3259 3358
rect 3160 3341 3162 3357
rect 3158 3340 3164 3341
rect 3158 3336 3159 3340
rect 3163 3336 3164 3340
rect 3158 3335 3164 3336
rect 2650 3331 2656 3332
rect 2650 3327 2651 3331
rect 2655 3327 2656 3331
rect 2650 3326 2656 3327
rect 2798 3331 2804 3332
rect 2798 3327 2799 3331
rect 2803 3327 2804 3331
rect 2798 3326 2804 3327
rect 3134 3331 3140 3332
rect 3134 3327 3135 3331
rect 3139 3327 3140 3331
rect 3134 3326 3140 3327
rect 2590 3302 2596 3303
rect 2590 3298 2591 3302
rect 2595 3298 2596 3302
rect 2590 3297 2596 3298
rect 2574 3291 2580 3292
rect 2574 3287 2575 3291
rect 2579 3287 2580 3291
rect 2574 3286 2580 3287
rect 2592 3275 2594 3297
rect 2652 3292 2654 3326
rect 2726 3302 2732 3303
rect 2726 3298 2727 3302
rect 2731 3298 2732 3302
rect 2726 3297 2732 3298
rect 2650 3291 2656 3292
rect 2650 3287 2651 3291
rect 2655 3287 2656 3291
rect 2650 3286 2656 3287
rect 2728 3275 2730 3297
rect 2800 3292 2802 3326
rect 2870 3302 2876 3303
rect 2870 3298 2871 3302
rect 2875 3298 2876 3302
rect 2870 3297 2876 3298
rect 3014 3302 3020 3303
rect 3014 3298 3015 3302
rect 3019 3298 3020 3302
rect 3014 3297 3020 3298
rect 3166 3302 3172 3303
rect 3166 3298 3167 3302
rect 3171 3298 3172 3302
rect 3166 3297 3172 3298
rect 2798 3291 2804 3292
rect 2798 3287 2799 3291
rect 2803 3287 2804 3291
rect 2798 3286 2804 3287
rect 2872 3275 2874 3297
rect 3006 3291 3012 3292
rect 3006 3287 3007 3291
rect 3011 3287 3012 3291
rect 3006 3286 3012 3287
rect 2231 3274 2235 3275
rect 2231 3269 2235 3270
rect 2279 3274 2283 3275
rect 2279 3269 2283 3270
rect 2343 3274 2347 3275
rect 2343 3269 2347 3270
rect 2415 3274 2419 3275
rect 2422 3271 2423 3275
rect 2427 3271 2428 3275
rect 2422 3270 2428 3271
rect 2463 3274 2467 3275
rect 2415 3269 2419 3270
rect 2254 3267 2260 3268
rect 2254 3263 2255 3267
rect 2259 3263 2260 3267
rect 2254 3262 2260 3263
rect 1830 3230 1836 3231
rect 2142 3231 2148 3232
rect 1742 3227 1748 3228
rect 1112 3211 1114 3227
rect 1248 3211 1250 3227
rect 1376 3211 1378 3227
rect 1504 3211 1506 3227
rect 1632 3211 1634 3227
rect 1744 3211 1746 3227
rect 1758 3215 1764 3216
rect 1758 3211 1759 3215
rect 1763 3211 1764 3215
rect 1832 3211 1834 3230
rect 2142 3227 2143 3231
rect 2147 3227 2148 3231
rect 2142 3226 2148 3227
rect 1870 3223 1876 3224
rect 1870 3219 1871 3223
rect 1875 3219 1876 3223
rect 1870 3218 1876 3219
rect 2126 3220 2132 3221
rect 1023 3210 1027 3211
rect 1023 3205 1027 3206
rect 1111 3210 1115 3211
rect 1111 3205 1115 3206
rect 1191 3210 1195 3211
rect 1191 3205 1195 3206
rect 1247 3210 1251 3211
rect 1247 3205 1251 3206
rect 1375 3210 1379 3211
rect 1375 3205 1379 3206
rect 1503 3210 1507 3211
rect 1503 3205 1507 3206
rect 1567 3210 1571 3211
rect 1567 3205 1571 3206
rect 1631 3210 1635 3211
rect 1631 3205 1635 3206
rect 1743 3210 1747 3211
rect 1758 3210 1764 3211
rect 1831 3210 1835 3211
rect 1743 3205 1747 3206
rect 1024 3189 1026 3205
rect 1192 3189 1194 3205
rect 1376 3189 1378 3205
rect 1568 3189 1570 3205
rect 1744 3189 1746 3205
rect 1022 3188 1028 3189
rect 1022 3184 1023 3188
rect 1027 3184 1028 3188
rect 1022 3183 1028 3184
rect 1190 3188 1196 3189
rect 1190 3184 1191 3188
rect 1195 3184 1196 3188
rect 1190 3183 1196 3184
rect 1374 3188 1380 3189
rect 1374 3184 1375 3188
rect 1379 3184 1380 3188
rect 1374 3183 1380 3184
rect 1566 3188 1572 3189
rect 1566 3184 1567 3188
rect 1571 3184 1572 3188
rect 1566 3183 1572 3184
rect 1742 3188 1748 3189
rect 1742 3184 1743 3188
rect 1747 3184 1748 3188
rect 1742 3183 1748 3184
rect 554 3179 560 3180
rect 554 3175 555 3179
rect 559 3175 560 3179
rect 554 3174 560 3175
rect 642 3179 648 3180
rect 642 3175 643 3179
rect 647 3175 648 3179
rect 642 3174 648 3175
rect 730 3179 736 3180
rect 730 3175 731 3179
rect 735 3175 736 3179
rect 730 3174 736 3175
rect 834 3179 840 3180
rect 834 3175 835 3179
rect 839 3175 840 3179
rect 834 3174 840 3175
rect 842 3179 848 3180
rect 842 3175 843 3179
rect 847 3175 848 3179
rect 842 3174 848 3175
rect 990 3179 996 3180
rect 990 3175 991 3179
rect 995 3175 996 3179
rect 990 3174 996 3175
rect 1106 3179 1112 3180
rect 1106 3175 1107 3179
rect 1111 3175 1112 3179
rect 1106 3174 1112 3175
rect 1478 3179 1484 3180
rect 1478 3175 1479 3179
rect 1483 3175 1484 3179
rect 1478 3174 1484 3175
rect 1486 3179 1492 3180
rect 1486 3175 1487 3179
rect 1491 3175 1492 3179
rect 1486 3174 1492 3175
rect 556 3140 558 3174
rect 582 3150 588 3151
rect 582 3146 583 3150
rect 587 3146 588 3150
rect 582 3145 588 3146
rect 635 3148 639 3149
rect 502 3139 508 3140
rect 502 3135 503 3139
rect 507 3135 508 3139
rect 502 3134 508 3135
rect 554 3139 560 3140
rect 554 3135 555 3139
rect 559 3135 560 3139
rect 554 3134 560 3135
rect 584 3131 586 3145
rect 635 3143 639 3144
rect 111 3130 115 3131
rect 111 3125 115 3126
rect 495 3130 499 3131
rect 495 3125 499 3126
rect 583 3130 587 3131
rect 583 3125 587 3126
rect 591 3130 595 3131
rect 591 3125 595 3126
rect 112 3097 114 3125
rect 592 3115 594 3125
rect 636 3124 638 3143
rect 644 3140 646 3174
rect 670 3150 676 3151
rect 670 3146 671 3150
rect 675 3146 676 3150
rect 670 3145 676 3146
rect 642 3139 648 3140
rect 642 3135 643 3139
rect 647 3135 648 3139
rect 642 3134 648 3135
rect 672 3131 674 3145
rect 732 3140 734 3174
rect 774 3150 780 3151
rect 774 3146 775 3150
rect 779 3146 780 3150
rect 774 3145 780 3146
rect 730 3139 736 3140
rect 730 3135 731 3139
rect 735 3135 736 3139
rect 730 3134 736 3135
rect 776 3131 778 3145
rect 836 3140 838 3174
rect 844 3149 846 3174
rect 894 3150 900 3151
rect 843 3148 847 3149
rect 894 3146 895 3150
rect 899 3146 900 3150
rect 894 3145 900 3146
rect 1030 3150 1036 3151
rect 1030 3146 1031 3150
rect 1035 3146 1036 3150
rect 1030 3145 1036 3146
rect 843 3143 847 3144
rect 834 3139 840 3140
rect 834 3135 835 3139
rect 839 3135 840 3139
rect 834 3134 840 3135
rect 896 3131 898 3145
rect 1032 3131 1034 3145
rect 1108 3140 1110 3174
rect 1198 3150 1204 3151
rect 1198 3146 1199 3150
rect 1203 3146 1204 3150
rect 1382 3150 1388 3151
rect 1198 3145 1204 3146
rect 1207 3148 1211 3149
rect 1106 3139 1112 3140
rect 1106 3135 1107 3139
rect 1111 3135 1112 3139
rect 1106 3134 1112 3135
rect 1200 3131 1202 3145
rect 1382 3146 1383 3150
rect 1387 3146 1388 3150
rect 1382 3145 1388 3146
rect 1207 3143 1211 3144
rect 1208 3140 1210 3143
rect 1206 3139 1212 3140
rect 1206 3135 1207 3139
rect 1211 3135 1212 3139
rect 1206 3134 1212 3135
rect 1384 3131 1386 3145
rect 1480 3140 1482 3174
rect 1488 3149 1490 3174
rect 1574 3150 1580 3151
rect 1487 3148 1491 3149
rect 1574 3146 1575 3150
rect 1579 3146 1580 3150
rect 1574 3145 1580 3146
rect 1750 3150 1756 3151
rect 1750 3146 1751 3150
rect 1755 3146 1756 3150
rect 1750 3145 1756 3146
rect 1487 3143 1491 3144
rect 1390 3139 1396 3140
rect 1390 3135 1391 3139
rect 1395 3135 1396 3139
rect 1390 3134 1396 3135
rect 1478 3139 1484 3140
rect 1478 3135 1479 3139
rect 1483 3135 1484 3139
rect 1478 3134 1484 3135
rect 671 3130 675 3131
rect 671 3125 675 3126
rect 759 3130 763 3131
rect 759 3125 763 3126
rect 775 3130 779 3131
rect 775 3125 779 3126
rect 847 3130 851 3131
rect 847 3125 851 3126
rect 895 3130 899 3131
rect 895 3125 899 3126
rect 935 3130 939 3131
rect 935 3125 939 3126
rect 1023 3130 1027 3131
rect 1023 3125 1027 3126
rect 1031 3130 1035 3131
rect 1031 3125 1035 3126
rect 1111 3130 1115 3131
rect 1111 3125 1115 3126
rect 1199 3130 1203 3131
rect 1199 3125 1203 3126
rect 1287 3130 1291 3131
rect 1287 3125 1291 3126
rect 1375 3130 1379 3131
rect 1375 3125 1379 3126
rect 1383 3130 1387 3131
rect 1383 3125 1387 3126
rect 634 3123 640 3124
rect 634 3119 635 3123
rect 639 3119 640 3123
rect 634 3118 640 3119
rect 642 3123 648 3124
rect 642 3119 643 3123
rect 647 3119 648 3123
rect 642 3118 648 3119
rect 590 3114 596 3115
rect 590 3110 591 3114
rect 595 3110 596 3114
rect 590 3109 596 3110
rect 110 3096 116 3097
rect 110 3092 111 3096
rect 115 3092 116 3096
rect 110 3091 116 3092
rect 644 3088 646 3118
rect 672 3115 674 3125
rect 722 3123 728 3124
rect 722 3119 723 3123
rect 727 3119 728 3123
rect 722 3118 728 3119
rect 670 3114 676 3115
rect 670 3110 671 3114
rect 675 3110 676 3114
rect 670 3109 676 3110
rect 724 3088 726 3118
rect 760 3115 762 3125
rect 810 3123 816 3124
rect 810 3119 811 3123
rect 815 3119 816 3123
rect 810 3118 816 3119
rect 758 3114 764 3115
rect 758 3110 759 3114
rect 763 3110 764 3114
rect 758 3109 764 3110
rect 812 3088 814 3118
rect 848 3115 850 3125
rect 926 3123 932 3124
rect 926 3119 927 3123
rect 931 3119 932 3123
rect 926 3118 932 3119
rect 846 3114 852 3115
rect 846 3110 847 3114
rect 851 3110 852 3114
rect 846 3109 852 3110
rect 928 3088 930 3118
rect 936 3115 938 3125
rect 1024 3115 1026 3125
rect 1066 3123 1072 3124
rect 1066 3119 1067 3123
rect 1071 3119 1072 3123
rect 1066 3118 1072 3119
rect 1074 3123 1080 3124
rect 1074 3119 1075 3123
rect 1079 3119 1080 3123
rect 1074 3118 1080 3119
rect 934 3114 940 3115
rect 934 3110 935 3114
rect 939 3110 940 3114
rect 934 3109 940 3110
rect 1022 3114 1028 3115
rect 1022 3110 1023 3114
rect 1027 3110 1028 3114
rect 1022 3109 1028 3110
rect 642 3087 648 3088
rect 642 3083 643 3087
rect 647 3083 648 3087
rect 642 3082 648 3083
rect 722 3087 728 3088
rect 722 3083 723 3087
rect 727 3083 728 3087
rect 722 3082 728 3083
rect 810 3087 816 3088
rect 810 3083 811 3087
rect 815 3083 816 3087
rect 810 3082 816 3083
rect 926 3087 932 3088
rect 926 3083 927 3087
rect 931 3083 932 3087
rect 926 3082 932 3083
rect 986 3087 992 3088
rect 986 3083 987 3087
rect 991 3083 992 3087
rect 986 3082 992 3083
rect 110 3079 116 3080
rect 110 3075 111 3079
rect 115 3075 116 3079
rect 110 3074 116 3075
rect 582 3076 588 3077
rect 112 3051 114 3074
rect 582 3072 583 3076
rect 587 3072 588 3076
rect 582 3071 588 3072
rect 662 3076 668 3077
rect 662 3072 663 3076
rect 667 3072 668 3076
rect 662 3071 668 3072
rect 750 3076 756 3077
rect 750 3072 751 3076
rect 755 3072 756 3076
rect 750 3071 756 3072
rect 838 3076 844 3077
rect 838 3072 839 3076
rect 843 3072 844 3076
rect 838 3071 844 3072
rect 926 3076 932 3077
rect 926 3072 927 3076
rect 931 3072 932 3076
rect 926 3071 932 3072
rect 584 3051 586 3071
rect 664 3051 666 3071
rect 752 3051 754 3071
rect 840 3051 842 3071
rect 928 3051 930 3071
rect 111 3050 115 3051
rect 111 3045 115 3046
rect 543 3050 547 3051
rect 543 3045 547 3046
rect 583 3050 587 3051
rect 583 3045 587 3046
rect 623 3050 627 3051
rect 623 3045 627 3046
rect 663 3050 667 3051
rect 663 3045 667 3046
rect 711 3050 715 3051
rect 711 3045 715 3046
rect 751 3050 755 3051
rect 751 3045 755 3046
rect 807 3050 811 3051
rect 807 3045 811 3046
rect 839 3050 843 3051
rect 839 3045 843 3046
rect 903 3050 907 3051
rect 903 3045 907 3046
rect 927 3050 931 3051
rect 927 3045 931 3046
rect 112 3026 114 3045
rect 544 3029 546 3045
rect 624 3029 626 3045
rect 712 3029 714 3045
rect 808 3029 810 3045
rect 904 3029 906 3045
rect 542 3028 548 3029
rect 110 3025 116 3026
rect 110 3021 111 3025
rect 115 3021 116 3025
rect 542 3024 543 3028
rect 547 3024 548 3028
rect 542 3023 548 3024
rect 622 3028 628 3029
rect 622 3024 623 3028
rect 627 3024 628 3028
rect 622 3023 628 3024
rect 710 3028 716 3029
rect 710 3024 711 3028
rect 715 3024 716 3028
rect 710 3023 716 3024
rect 806 3028 812 3029
rect 806 3024 807 3028
rect 811 3024 812 3028
rect 806 3023 812 3024
rect 902 3028 908 3029
rect 902 3024 903 3028
rect 907 3024 908 3028
rect 902 3023 908 3024
rect 110 3020 116 3021
rect 610 3019 616 3020
rect 610 3015 611 3019
rect 615 3015 616 3019
rect 610 3014 616 3015
rect 694 3019 700 3020
rect 694 3015 695 3019
rect 699 3015 700 3019
rect 694 3014 700 3015
rect 778 3019 784 3020
rect 778 3015 779 3019
rect 783 3015 784 3019
rect 778 3014 784 3015
rect 874 3019 880 3020
rect 874 3015 875 3019
rect 879 3015 880 3019
rect 874 3014 880 3015
rect 970 3019 976 3020
rect 970 3015 971 3019
rect 975 3015 976 3019
rect 970 3014 976 3015
rect 602 3011 608 3012
rect 110 3008 116 3009
rect 110 3004 111 3008
rect 115 3004 116 3008
rect 602 3007 603 3011
rect 607 3007 608 3011
rect 602 3006 608 3007
rect 110 3003 116 3004
rect 112 2975 114 3003
rect 550 2990 556 2991
rect 550 2986 551 2990
rect 555 2986 556 2990
rect 550 2985 556 2986
rect 552 2975 554 2985
rect 604 2980 606 3006
rect 612 2980 614 3014
rect 630 2990 636 2991
rect 630 2986 631 2990
rect 635 2986 636 2990
rect 630 2985 636 2986
rect 602 2979 608 2980
rect 602 2975 603 2979
rect 607 2975 608 2979
rect 111 2974 115 2975
rect 111 2969 115 2970
rect 471 2974 475 2975
rect 471 2969 475 2970
rect 551 2974 555 2975
rect 551 2969 555 2970
rect 575 2974 579 2975
rect 602 2974 608 2975
rect 610 2979 616 2980
rect 610 2975 611 2979
rect 615 2975 616 2979
rect 632 2975 634 2985
rect 610 2974 616 2975
rect 631 2974 635 2975
rect 575 2969 579 2970
rect 631 2969 635 2970
rect 687 2974 691 2975
rect 687 2969 691 2970
rect 112 2941 114 2969
rect 472 2959 474 2969
rect 530 2967 536 2968
rect 530 2963 531 2967
rect 535 2963 536 2967
rect 530 2962 536 2963
rect 470 2958 476 2959
rect 470 2954 471 2958
rect 475 2954 476 2958
rect 470 2953 476 2954
rect 110 2940 116 2941
rect 110 2936 111 2940
rect 115 2936 116 2940
rect 110 2935 116 2936
rect 532 2932 534 2962
rect 576 2959 578 2969
rect 654 2967 660 2968
rect 654 2963 655 2967
rect 659 2963 660 2967
rect 654 2962 660 2963
rect 574 2958 580 2959
rect 574 2954 575 2958
rect 579 2954 580 2958
rect 574 2953 580 2954
rect 656 2949 658 2962
rect 688 2959 690 2969
rect 696 2968 698 3014
rect 718 2990 724 2991
rect 718 2986 719 2990
rect 723 2986 724 2990
rect 718 2985 724 2986
rect 720 2975 722 2985
rect 780 2980 782 3014
rect 814 2990 820 2991
rect 814 2986 815 2990
rect 819 2986 820 2990
rect 814 2985 820 2986
rect 778 2979 784 2980
rect 778 2975 779 2979
rect 783 2975 784 2979
rect 816 2975 818 2985
rect 876 2980 878 3014
rect 910 2990 916 2991
rect 910 2986 911 2990
rect 915 2986 916 2990
rect 910 2985 916 2986
rect 874 2979 880 2980
rect 874 2975 875 2979
rect 879 2975 880 2979
rect 912 2975 914 2985
rect 972 2980 974 3014
rect 988 2980 990 3082
rect 1014 3076 1020 3077
rect 1014 3072 1015 3076
rect 1019 3072 1020 3076
rect 1014 3071 1020 3072
rect 1016 3051 1018 3071
rect 999 3050 1003 3051
rect 999 3045 1003 3046
rect 1015 3050 1019 3051
rect 1015 3045 1019 3046
rect 1000 3029 1002 3045
rect 998 3028 1004 3029
rect 998 3024 999 3028
rect 1003 3024 1004 3028
rect 998 3023 1004 3024
rect 1068 3020 1070 3118
rect 1076 3088 1078 3118
rect 1112 3115 1114 3125
rect 1162 3123 1168 3124
rect 1162 3119 1163 3123
rect 1167 3119 1168 3123
rect 1162 3118 1168 3119
rect 1110 3114 1116 3115
rect 1110 3110 1111 3114
rect 1115 3110 1116 3114
rect 1110 3109 1116 3110
rect 1164 3088 1166 3118
rect 1200 3115 1202 3125
rect 1250 3123 1256 3124
rect 1250 3119 1251 3123
rect 1255 3119 1256 3123
rect 1250 3118 1256 3119
rect 1198 3114 1204 3115
rect 1198 3110 1199 3114
rect 1203 3110 1204 3114
rect 1198 3109 1204 3110
rect 1252 3088 1254 3118
rect 1288 3115 1290 3125
rect 1338 3123 1344 3124
rect 1338 3119 1339 3123
rect 1343 3119 1344 3123
rect 1338 3118 1344 3119
rect 1286 3114 1292 3115
rect 1286 3110 1287 3114
rect 1291 3110 1292 3114
rect 1286 3109 1292 3110
rect 1340 3088 1342 3118
rect 1376 3115 1378 3125
rect 1374 3114 1380 3115
rect 1374 3110 1375 3114
rect 1379 3110 1380 3114
rect 1374 3109 1380 3110
rect 1392 3088 1394 3134
rect 1576 3131 1578 3145
rect 1752 3131 1754 3145
rect 1760 3140 1762 3210
rect 1831 3205 1835 3206
rect 1832 3186 1834 3205
rect 1872 3195 1874 3218
rect 2126 3216 2127 3220
rect 2131 3216 2132 3220
rect 2126 3215 2132 3216
rect 2128 3195 2130 3215
rect 1871 3194 1875 3195
rect 1871 3189 1875 3190
rect 1895 3194 1899 3195
rect 1895 3189 1899 3190
rect 1991 3194 1995 3195
rect 1991 3189 1995 3190
rect 2119 3194 2123 3195
rect 2119 3189 2123 3190
rect 2127 3194 2131 3195
rect 2127 3189 2131 3190
rect 2247 3194 2251 3195
rect 2247 3189 2251 3190
rect 1830 3185 1836 3186
rect 1830 3181 1831 3185
rect 1835 3181 1836 3185
rect 1830 3180 1836 3181
rect 1818 3179 1824 3180
rect 1818 3175 1819 3179
rect 1823 3175 1824 3179
rect 1818 3174 1824 3175
rect 1758 3139 1764 3140
rect 1758 3135 1759 3139
rect 1763 3135 1764 3139
rect 1758 3134 1764 3135
rect 1575 3130 1579 3131
rect 1575 3125 1579 3126
rect 1751 3130 1755 3131
rect 1751 3125 1755 3126
rect 1820 3124 1822 3174
rect 1872 3170 1874 3189
rect 1896 3173 1898 3189
rect 1992 3173 1994 3189
rect 2120 3173 2122 3189
rect 2248 3173 2250 3189
rect 1894 3172 1900 3173
rect 1870 3169 1876 3170
rect 1830 3168 1836 3169
rect 1830 3164 1831 3168
rect 1835 3164 1836 3168
rect 1870 3165 1871 3169
rect 1875 3165 1876 3169
rect 1894 3168 1895 3172
rect 1899 3168 1900 3172
rect 1894 3167 1900 3168
rect 1990 3172 1996 3173
rect 1990 3168 1991 3172
rect 1995 3168 1996 3172
rect 1990 3167 1996 3168
rect 2118 3172 2124 3173
rect 2118 3168 2119 3172
rect 2123 3168 2124 3172
rect 2118 3167 2124 3168
rect 2246 3172 2252 3173
rect 2246 3168 2247 3172
rect 2251 3168 2252 3172
rect 2246 3167 2252 3168
rect 1870 3164 1876 3165
rect 1830 3163 1836 3164
rect 1962 3163 1968 3164
rect 1832 3131 1834 3163
rect 1962 3159 1963 3163
rect 1967 3159 1968 3163
rect 1962 3158 1968 3159
rect 2062 3163 2068 3164
rect 2062 3159 2063 3163
rect 2067 3159 2068 3163
rect 2256 3160 2258 3262
rect 2280 3259 2282 3269
rect 2330 3267 2336 3268
rect 2330 3263 2331 3267
rect 2335 3263 2336 3267
rect 2330 3262 2336 3263
rect 2278 3258 2284 3259
rect 2278 3254 2279 3258
rect 2283 3254 2284 3258
rect 2278 3253 2284 3254
rect 2332 3232 2334 3262
rect 2416 3259 2418 3269
rect 2414 3258 2420 3259
rect 2414 3254 2415 3258
rect 2419 3254 2420 3258
rect 2414 3253 2420 3254
rect 2424 3232 2426 3270
rect 2463 3269 2467 3270
rect 2551 3274 2555 3275
rect 2551 3269 2555 3270
rect 2591 3274 2595 3275
rect 2591 3269 2595 3270
rect 2687 3274 2691 3275
rect 2687 3269 2691 3270
rect 2727 3274 2731 3275
rect 2727 3269 2731 3270
rect 2823 3274 2827 3275
rect 2823 3269 2827 3270
rect 2871 3274 2875 3275
rect 2871 3269 2875 3270
rect 2959 3274 2963 3275
rect 2959 3269 2963 3270
rect 2552 3259 2554 3269
rect 2610 3267 2616 3268
rect 2610 3263 2611 3267
rect 2615 3263 2616 3267
rect 2610 3262 2616 3263
rect 2550 3258 2556 3259
rect 2550 3254 2551 3258
rect 2555 3254 2556 3258
rect 2550 3253 2556 3254
rect 2612 3232 2614 3262
rect 2688 3259 2690 3269
rect 2746 3267 2752 3268
rect 2746 3263 2747 3267
rect 2751 3263 2752 3267
rect 2746 3262 2752 3263
rect 2686 3258 2692 3259
rect 2686 3254 2687 3258
rect 2691 3254 2692 3258
rect 2686 3253 2692 3254
rect 2748 3232 2750 3262
rect 2824 3259 2826 3269
rect 2960 3259 2962 3269
rect 2822 3258 2828 3259
rect 2822 3254 2823 3258
rect 2827 3254 2828 3258
rect 2822 3253 2828 3254
rect 2958 3258 2964 3259
rect 2958 3254 2959 3258
rect 2963 3254 2964 3258
rect 2958 3253 2964 3254
rect 3008 3232 3010 3286
rect 3016 3275 3018 3297
rect 3168 3275 3170 3297
rect 3304 3292 3306 3394
rect 3590 3391 3596 3392
rect 3414 3388 3420 3389
rect 3414 3384 3415 3388
rect 3419 3384 3420 3388
rect 3590 3387 3591 3391
rect 3595 3387 3596 3391
rect 3590 3386 3596 3387
rect 3414 3383 3420 3384
rect 3416 3363 3418 3383
rect 3592 3363 3594 3386
rect 3311 3362 3315 3363
rect 3311 3357 3315 3358
rect 3415 3362 3419 3363
rect 3415 3357 3419 3358
rect 3471 3362 3475 3363
rect 3471 3357 3475 3358
rect 3591 3362 3595 3363
rect 3591 3357 3595 3358
rect 3312 3341 3314 3357
rect 3472 3341 3474 3357
rect 3310 3340 3316 3341
rect 3310 3336 3311 3340
rect 3315 3336 3316 3340
rect 3310 3335 3316 3336
rect 3470 3340 3476 3341
rect 3470 3336 3471 3340
rect 3475 3336 3476 3340
rect 3592 3338 3594 3357
rect 3470 3335 3476 3336
rect 3590 3337 3596 3338
rect 3590 3333 3591 3337
rect 3595 3333 3596 3337
rect 3590 3332 3596 3333
rect 3394 3331 3400 3332
rect 3394 3327 3395 3331
rect 3399 3327 3400 3331
rect 3394 3326 3400 3327
rect 3318 3302 3324 3303
rect 3318 3298 3319 3302
rect 3323 3298 3324 3302
rect 3318 3297 3324 3298
rect 3302 3291 3308 3292
rect 3302 3287 3303 3291
rect 3307 3287 3308 3291
rect 3302 3286 3308 3287
rect 3320 3275 3322 3297
rect 3396 3292 3398 3326
rect 3530 3323 3536 3324
rect 3530 3319 3531 3323
rect 3535 3319 3536 3323
rect 3530 3318 3536 3319
rect 3590 3320 3596 3321
rect 3478 3302 3484 3303
rect 3478 3298 3479 3302
rect 3483 3298 3484 3302
rect 3478 3297 3484 3298
rect 3394 3291 3400 3292
rect 3394 3287 3395 3291
rect 3399 3287 3400 3291
rect 3394 3286 3400 3287
rect 3480 3275 3482 3297
rect 3015 3274 3019 3275
rect 3015 3269 3019 3270
rect 3095 3274 3099 3275
rect 3095 3269 3099 3270
rect 3167 3274 3171 3275
rect 3167 3269 3171 3270
rect 3231 3274 3235 3275
rect 3231 3269 3235 3270
rect 3319 3274 3323 3275
rect 3319 3269 3323 3270
rect 3375 3274 3379 3275
rect 3375 3269 3379 3270
rect 3479 3274 3483 3275
rect 3479 3269 3483 3270
rect 3511 3274 3515 3275
rect 3511 3269 3515 3270
rect 3022 3267 3028 3268
rect 3022 3263 3023 3267
rect 3027 3263 3028 3267
rect 3022 3262 3028 3263
rect 3024 3232 3026 3262
rect 3096 3259 3098 3269
rect 3186 3267 3192 3268
rect 3186 3263 3187 3267
rect 3191 3263 3192 3267
rect 3186 3262 3192 3263
rect 3094 3258 3100 3259
rect 3094 3254 3095 3258
rect 3099 3254 3100 3258
rect 3094 3253 3100 3254
rect 3188 3232 3190 3262
rect 3232 3259 3234 3269
rect 3266 3267 3272 3268
rect 3266 3263 3267 3267
rect 3271 3263 3272 3267
rect 3266 3262 3272 3263
rect 3230 3258 3236 3259
rect 3230 3254 3231 3258
rect 3235 3254 3236 3258
rect 3230 3253 3236 3254
rect 2330 3231 2336 3232
rect 2330 3227 2331 3231
rect 2335 3227 2336 3231
rect 2330 3226 2336 3227
rect 2422 3231 2428 3232
rect 2422 3227 2423 3231
rect 2427 3227 2428 3231
rect 2422 3226 2428 3227
rect 2610 3231 2616 3232
rect 2610 3227 2611 3231
rect 2615 3227 2616 3231
rect 2610 3226 2616 3227
rect 2746 3231 2752 3232
rect 2746 3227 2747 3231
rect 2751 3227 2752 3231
rect 2746 3226 2752 3227
rect 3006 3231 3012 3232
rect 3006 3227 3007 3231
rect 3011 3227 3012 3231
rect 3006 3226 3012 3227
rect 3022 3231 3028 3232
rect 3022 3227 3023 3231
rect 3027 3227 3028 3231
rect 3022 3226 3028 3227
rect 3186 3231 3192 3232
rect 3186 3227 3187 3231
rect 3191 3227 3192 3231
rect 3186 3226 3192 3227
rect 2270 3220 2276 3221
rect 2270 3216 2271 3220
rect 2275 3216 2276 3220
rect 2270 3215 2276 3216
rect 2406 3220 2412 3221
rect 2406 3216 2407 3220
rect 2411 3216 2412 3220
rect 2406 3215 2412 3216
rect 2542 3220 2548 3221
rect 2542 3216 2543 3220
rect 2547 3216 2548 3220
rect 2542 3215 2548 3216
rect 2678 3220 2684 3221
rect 2678 3216 2679 3220
rect 2683 3216 2684 3220
rect 2678 3215 2684 3216
rect 2814 3220 2820 3221
rect 2814 3216 2815 3220
rect 2819 3216 2820 3220
rect 2814 3215 2820 3216
rect 2950 3220 2956 3221
rect 2950 3216 2951 3220
rect 2955 3216 2956 3220
rect 2950 3215 2956 3216
rect 3086 3220 3092 3221
rect 3086 3216 3087 3220
rect 3091 3216 3092 3220
rect 3086 3215 3092 3216
rect 3222 3220 3228 3221
rect 3222 3216 3223 3220
rect 3227 3216 3228 3220
rect 3222 3215 3228 3216
rect 2272 3195 2274 3215
rect 2408 3195 2410 3215
rect 2544 3195 2546 3215
rect 2550 3203 2556 3204
rect 2550 3199 2551 3203
rect 2555 3199 2556 3203
rect 2550 3198 2556 3199
rect 2271 3194 2275 3195
rect 2271 3189 2275 3190
rect 2383 3194 2387 3195
rect 2383 3189 2387 3190
rect 2407 3194 2411 3195
rect 2407 3189 2411 3190
rect 2511 3194 2515 3195
rect 2511 3189 2515 3190
rect 2543 3194 2547 3195
rect 2543 3189 2547 3190
rect 2384 3173 2386 3189
rect 2512 3173 2514 3189
rect 2382 3172 2388 3173
rect 2382 3168 2383 3172
rect 2387 3168 2388 3172
rect 2382 3167 2388 3168
rect 2510 3172 2516 3173
rect 2510 3168 2511 3172
rect 2515 3168 2516 3172
rect 2510 3167 2516 3168
rect 2350 3163 2356 3164
rect 2062 3158 2068 3159
rect 2254 3159 2260 3160
rect 1870 3152 1876 3153
rect 1870 3148 1871 3152
rect 1875 3148 1876 3152
rect 1870 3147 1876 3148
rect 1831 3130 1835 3131
rect 1831 3125 1835 3126
rect 1818 3123 1824 3124
rect 1818 3119 1819 3123
rect 1823 3119 1824 3123
rect 1818 3118 1824 3119
rect 1832 3097 1834 3125
rect 1872 3103 1874 3147
rect 1902 3134 1908 3135
rect 1902 3130 1903 3134
rect 1907 3130 1908 3134
rect 1902 3129 1908 3130
rect 1904 3103 1906 3129
rect 1964 3124 1966 3158
rect 1998 3134 2004 3135
rect 1998 3130 1999 3134
rect 2003 3130 2004 3134
rect 1998 3129 2004 3130
rect 1962 3123 1968 3124
rect 1962 3119 1963 3123
rect 1967 3119 1968 3123
rect 1962 3118 1968 3119
rect 2000 3103 2002 3129
rect 2064 3124 2066 3158
rect 2178 3155 2184 3156
rect 2178 3151 2179 3155
rect 2183 3151 2184 3155
rect 2254 3155 2255 3159
rect 2259 3155 2260 3159
rect 2350 3159 2351 3163
rect 2355 3159 2356 3163
rect 2350 3158 2356 3159
rect 2254 3154 2260 3155
rect 2178 3150 2184 3151
rect 2126 3134 2132 3135
rect 2126 3130 2127 3134
rect 2131 3130 2132 3134
rect 2126 3129 2132 3130
rect 2062 3123 2068 3124
rect 2062 3119 2063 3123
rect 2067 3119 2068 3123
rect 2062 3118 2068 3119
rect 2128 3103 2130 3129
rect 1871 3102 1875 3103
rect 1871 3097 1875 3098
rect 1903 3102 1907 3103
rect 1903 3097 1907 3098
rect 1999 3102 2003 3103
rect 1999 3097 2003 3098
rect 2015 3102 2019 3103
rect 2015 3097 2019 3098
rect 2127 3102 2131 3103
rect 2127 3097 2131 3098
rect 1830 3096 1836 3097
rect 1830 3092 1831 3096
rect 1835 3092 1836 3096
rect 1830 3091 1836 3092
rect 1074 3087 1080 3088
rect 1074 3083 1075 3087
rect 1079 3083 1080 3087
rect 1074 3082 1080 3083
rect 1162 3087 1168 3088
rect 1162 3083 1163 3087
rect 1167 3083 1168 3087
rect 1162 3082 1168 3083
rect 1250 3087 1256 3088
rect 1250 3083 1251 3087
rect 1255 3083 1256 3087
rect 1250 3082 1256 3083
rect 1338 3087 1344 3088
rect 1338 3083 1339 3087
rect 1343 3083 1344 3087
rect 1338 3082 1344 3083
rect 1390 3087 1396 3088
rect 1390 3083 1391 3087
rect 1395 3083 1396 3087
rect 1390 3082 1396 3083
rect 1830 3079 1836 3080
rect 1102 3076 1108 3077
rect 1102 3072 1103 3076
rect 1107 3072 1108 3076
rect 1102 3071 1108 3072
rect 1190 3076 1196 3077
rect 1190 3072 1191 3076
rect 1195 3072 1196 3076
rect 1190 3071 1196 3072
rect 1278 3076 1284 3077
rect 1278 3072 1279 3076
rect 1283 3072 1284 3076
rect 1278 3071 1284 3072
rect 1366 3076 1372 3077
rect 1366 3072 1367 3076
rect 1371 3072 1372 3076
rect 1830 3075 1831 3079
rect 1835 3075 1836 3079
rect 1830 3074 1836 3075
rect 1366 3071 1372 3072
rect 1104 3051 1106 3071
rect 1192 3051 1194 3071
rect 1280 3051 1282 3071
rect 1368 3051 1370 3071
rect 1832 3051 1834 3074
rect 1872 3069 1874 3097
rect 1904 3087 1906 3097
rect 1910 3095 1916 3096
rect 1910 3090 1911 3095
rect 1915 3090 1916 3095
rect 1954 3095 1960 3096
rect 1954 3091 1955 3095
rect 1959 3091 1960 3095
rect 1954 3090 1960 3091
rect 1911 3087 1915 3088
rect 1902 3086 1908 3087
rect 1902 3082 1903 3086
rect 1907 3082 1908 3086
rect 1902 3081 1908 3082
rect 1870 3068 1876 3069
rect 1870 3064 1871 3068
rect 1875 3064 1876 3068
rect 1870 3063 1876 3064
rect 1956 3060 1958 3090
rect 2016 3087 2018 3097
rect 2180 3096 2182 3150
rect 2254 3134 2260 3135
rect 2254 3130 2255 3134
rect 2259 3130 2260 3134
rect 2254 3129 2260 3130
rect 2256 3103 2258 3129
rect 2352 3124 2354 3158
rect 2390 3134 2396 3135
rect 2390 3130 2391 3134
rect 2395 3130 2396 3134
rect 2390 3129 2396 3130
rect 2518 3134 2524 3135
rect 2518 3130 2519 3134
rect 2523 3130 2524 3134
rect 2518 3129 2524 3130
rect 2350 3123 2356 3124
rect 2350 3119 2351 3123
rect 2355 3119 2356 3123
rect 2350 3118 2356 3119
rect 2392 3103 2394 3129
rect 2414 3123 2420 3124
rect 2414 3119 2415 3123
rect 2419 3119 2420 3123
rect 2414 3118 2420 3119
rect 2191 3102 2195 3103
rect 2191 3097 2195 3098
rect 2255 3102 2259 3103
rect 2255 3097 2259 3098
rect 2391 3102 2395 3103
rect 2391 3097 2395 3098
rect 2407 3102 2411 3103
rect 2407 3097 2411 3098
rect 2178 3095 2184 3096
rect 2178 3091 2179 3095
rect 2183 3091 2184 3095
rect 2178 3090 2184 3091
rect 2192 3087 2194 3097
rect 2346 3095 2352 3096
rect 2199 3092 2203 3093
rect 2346 3091 2347 3095
rect 2351 3091 2352 3095
rect 2346 3090 2352 3091
rect 2199 3087 2203 3088
rect 2014 3086 2020 3087
rect 2014 3082 2015 3086
rect 2019 3082 2020 3086
rect 2014 3081 2020 3082
rect 2190 3086 2196 3087
rect 2190 3082 2191 3086
rect 2195 3082 2196 3086
rect 2190 3081 2196 3082
rect 2200 3060 2202 3087
rect 1954 3059 1960 3060
rect 1954 3055 1955 3059
rect 1959 3055 1960 3059
rect 1954 3054 1960 3055
rect 2038 3059 2044 3060
rect 2038 3055 2039 3059
rect 2043 3055 2044 3059
rect 2038 3054 2044 3055
rect 2198 3059 2204 3060
rect 2198 3055 2199 3059
rect 2203 3055 2204 3059
rect 2198 3054 2204 3055
rect 1870 3051 1876 3052
rect 1087 3050 1091 3051
rect 1087 3045 1091 3046
rect 1103 3050 1107 3051
rect 1103 3045 1107 3046
rect 1183 3050 1187 3051
rect 1183 3045 1187 3046
rect 1191 3050 1195 3051
rect 1191 3045 1195 3046
rect 1279 3050 1283 3051
rect 1279 3045 1283 3046
rect 1367 3050 1371 3051
rect 1367 3045 1371 3046
rect 1375 3050 1379 3051
rect 1375 3045 1379 3046
rect 1471 3050 1475 3051
rect 1471 3045 1475 3046
rect 1831 3050 1835 3051
rect 1870 3047 1871 3051
rect 1875 3047 1876 3051
rect 1870 3046 1876 3047
rect 1894 3048 1900 3049
rect 1831 3045 1835 3046
rect 1088 3029 1090 3045
rect 1184 3029 1186 3045
rect 1280 3029 1282 3045
rect 1376 3029 1378 3045
rect 1472 3029 1474 3045
rect 1086 3028 1092 3029
rect 1086 3024 1087 3028
rect 1091 3024 1092 3028
rect 1086 3023 1092 3024
rect 1182 3028 1188 3029
rect 1182 3024 1183 3028
rect 1187 3024 1188 3028
rect 1182 3023 1188 3024
rect 1278 3028 1284 3029
rect 1278 3024 1279 3028
rect 1283 3024 1284 3028
rect 1278 3023 1284 3024
rect 1374 3028 1380 3029
rect 1374 3024 1375 3028
rect 1379 3024 1380 3028
rect 1374 3023 1380 3024
rect 1470 3028 1476 3029
rect 1470 3024 1471 3028
rect 1475 3024 1476 3028
rect 1832 3026 1834 3045
rect 1470 3023 1476 3024
rect 1830 3025 1836 3026
rect 1830 3021 1831 3025
rect 1835 3021 1836 3025
rect 1830 3020 1836 3021
rect 1066 3019 1072 3020
rect 1066 3015 1067 3019
rect 1071 3015 1072 3019
rect 1066 3014 1072 3015
rect 1154 3019 1160 3020
rect 1154 3015 1155 3019
rect 1159 3015 1160 3019
rect 1154 3014 1160 3015
rect 1254 3019 1260 3020
rect 1254 3015 1255 3019
rect 1259 3015 1260 3019
rect 1254 3014 1260 3015
rect 1346 3019 1352 3020
rect 1346 3015 1347 3019
rect 1351 3015 1352 3019
rect 1346 3014 1352 3015
rect 1442 3019 1448 3020
rect 1872 3019 1874 3046
rect 1894 3044 1895 3048
rect 1899 3044 1900 3048
rect 1894 3043 1900 3044
rect 2006 3048 2012 3049
rect 2006 3044 2007 3048
rect 2011 3044 2012 3048
rect 2006 3043 2012 3044
rect 1896 3019 1898 3043
rect 2008 3019 2010 3043
rect 1442 3015 1443 3019
rect 1447 3015 1448 3019
rect 1442 3014 1448 3015
rect 1871 3018 1875 3019
rect 1006 2990 1012 2991
rect 1006 2986 1007 2990
rect 1011 2986 1012 2990
rect 1006 2985 1012 2986
rect 1094 2990 1100 2991
rect 1094 2986 1095 2990
rect 1099 2986 1100 2990
rect 1094 2985 1100 2986
rect 970 2979 976 2980
rect 970 2975 971 2979
rect 975 2975 976 2979
rect 719 2974 723 2975
rect 778 2974 784 2975
rect 807 2974 811 2975
rect 719 2969 723 2970
rect 807 2969 811 2970
rect 815 2974 819 2975
rect 874 2974 880 2975
rect 911 2974 915 2975
rect 815 2969 819 2970
rect 911 2969 915 2970
rect 943 2974 947 2975
rect 970 2974 976 2975
rect 986 2979 992 2980
rect 986 2975 987 2979
rect 991 2975 992 2979
rect 1008 2975 1010 2985
rect 1096 2975 1098 2985
rect 1156 2980 1158 3014
rect 1190 2990 1196 2991
rect 1190 2986 1191 2990
rect 1195 2986 1196 2990
rect 1190 2985 1196 2986
rect 1154 2979 1160 2980
rect 1154 2975 1155 2979
rect 1159 2975 1160 2979
rect 1192 2975 1194 2985
rect 1256 2980 1258 3014
rect 1286 2990 1292 2991
rect 1286 2986 1287 2990
rect 1291 2986 1292 2990
rect 1286 2985 1292 2986
rect 1254 2979 1260 2980
rect 1254 2975 1255 2979
rect 1259 2975 1260 2979
rect 1288 2975 1290 2985
rect 1348 2980 1350 3014
rect 1382 2990 1388 2991
rect 1382 2986 1383 2990
rect 1387 2986 1388 2990
rect 1382 2985 1388 2986
rect 1346 2979 1352 2980
rect 1346 2975 1347 2979
rect 1351 2975 1352 2979
rect 1384 2975 1386 2985
rect 1444 2980 1446 3014
rect 1871 3013 1875 3014
rect 1895 3018 1899 3019
rect 1895 3013 1899 3014
rect 2007 3018 2011 3019
rect 2007 3013 2011 3014
rect 1830 3008 1836 3009
rect 1830 3004 1831 3008
rect 1835 3004 1836 3008
rect 1830 3003 1836 3004
rect 1478 2990 1484 2991
rect 1478 2986 1479 2990
rect 1483 2986 1484 2990
rect 1478 2985 1484 2986
rect 1442 2979 1448 2980
rect 1442 2975 1443 2979
rect 1447 2975 1448 2979
rect 1480 2975 1482 2985
rect 1598 2979 1604 2980
rect 1598 2975 1599 2979
rect 1603 2975 1604 2979
rect 1832 2975 1834 3003
rect 1872 2994 1874 3013
rect 1896 2997 1898 3013
rect 1894 2996 1900 2997
rect 1870 2993 1876 2994
rect 1870 2989 1871 2993
rect 1875 2989 1876 2993
rect 1894 2992 1895 2996
rect 1899 2992 1900 2996
rect 1894 2991 1900 2992
rect 1870 2988 1876 2989
rect 1962 2987 1968 2988
rect 1894 2983 1900 2984
rect 1894 2979 1895 2983
rect 1899 2979 1900 2983
rect 1962 2983 1963 2987
rect 1967 2983 1968 2987
rect 1962 2982 1968 2983
rect 1894 2978 1900 2979
rect 1870 2976 1876 2977
rect 986 2974 992 2975
rect 1007 2974 1011 2975
rect 943 2969 947 2970
rect 1007 2969 1011 2970
rect 1087 2974 1091 2975
rect 1087 2969 1091 2970
rect 1095 2974 1099 2975
rect 1154 2974 1160 2975
rect 1191 2974 1195 2975
rect 1095 2969 1099 2970
rect 1191 2969 1195 2970
rect 1247 2974 1251 2975
rect 1254 2974 1260 2975
rect 1287 2974 1291 2975
rect 1346 2974 1352 2975
rect 1383 2974 1387 2975
rect 1247 2969 1251 2970
rect 1287 2969 1291 2970
rect 1383 2969 1387 2970
rect 1415 2974 1419 2975
rect 1442 2974 1448 2975
rect 1479 2974 1483 2975
rect 1415 2969 1419 2970
rect 1479 2969 1483 2970
rect 1591 2974 1595 2975
rect 1598 2974 1604 2975
rect 1751 2974 1755 2975
rect 1591 2969 1595 2970
rect 694 2967 700 2968
rect 694 2963 695 2967
rect 699 2963 700 2967
rect 694 2962 700 2963
rect 738 2967 744 2968
rect 738 2963 739 2967
rect 743 2963 744 2967
rect 738 2962 744 2963
rect 686 2958 692 2959
rect 686 2954 687 2958
rect 691 2954 692 2958
rect 686 2953 692 2954
rect 655 2948 659 2949
rect 655 2943 659 2944
rect 740 2932 742 2962
rect 808 2959 810 2969
rect 858 2967 864 2968
rect 858 2963 859 2967
rect 863 2963 864 2967
rect 858 2962 864 2963
rect 806 2958 812 2959
rect 806 2954 807 2958
rect 811 2954 812 2958
rect 806 2953 812 2954
rect 860 2932 862 2962
rect 944 2959 946 2969
rect 1088 2959 1090 2969
rect 1102 2967 1108 2968
rect 1102 2963 1103 2967
rect 1107 2963 1108 2967
rect 1102 2962 1108 2963
rect 1138 2967 1144 2968
rect 1138 2963 1139 2967
rect 1143 2963 1144 2967
rect 1138 2962 1144 2963
rect 942 2958 948 2959
rect 942 2954 943 2958
rect 947 2954 948 2958
rect 942 2953 948 2954
rect 1086 2958 1092 2959
rect 1086 2954 1087 2958
rect 1091 2954 1092 2958
rect 1086 2953 1092 2954
rect 1104 2949 1106 2962
rect 951 2948 955 2949
rect 951 2943 955 2944
rect 1103 2948 1107 2949
rect 1103 2943 1107 2944
rect 952 2932 954 2943
rect 1140 2932 1142 2962
rect 1248 2959 1250 2969
rect 1298 2967 1304 2968
rect 1298 2963 1299 2967
rect 1303 2963 1304 2967
rect 1298 2962 1304 2963
rect 1246 2958 1252 2959
rect 1246 2954 1247 2958
rect 1251 2954 1252 2958
rect 1246 2953 1252 2954
rect 1300 2932 1302 2962
rect 1416 2959 1418 2969
rect 1466 2967 1472 2968
rect 1466 2963 1467 2967
rect 1471 2963 1472 2967
rect 1466 2962 1472 2963
rect 1414 2958 1420 2959
rect 1414 2954 1415 2958
rect 1419 2954 1420 2958
rect 1414 2953 1420 2954
rect 1307 2948 1311 2949
rect 1307 2943 1311 2944
rect 522 2931 528 2932
rect 522 2927 523 2931
rect 527 2927 528 2931
rect 522 2926 528 2927
rect 530 2931 536 2932
rect 530 2927 531 2931
rect 535 2927 536 2931
rect 530 2926 536 2927
rect 738 2931 744 2932
rect 738 2927 739 2931
rect 743 2927 744 2931
rect 738 2926 744 2927
rect 858 2931 864 2932
rect 858 2927 859 2931
rect 863 2927 864 2931
rect 858 2926 864 2927
rect 950 2931 956 2932
rect 950 2927 951 2931
rect 955 2927 956 2931
rect 950 2926 956 2927
rect 1138 2931 1144 2932
rect 1138 2927 1139 2931
rect 1143 2927 1144 2931
rect 1138 2926 1144 2927
rect 1298 2931 1304 2932
rect 1298 2927 1299 2931
rect 1303 2927 1304 2931
rect 1298 2926 1304 2927
rect 110 2923 116 2924
rect 110 2919 111 2923
rect 115 2919 116 2923
rect 110 2918 116 2919
rect 462 2920 468 2921
rect 112 2899 114 2918
rect 462 2916 463 2920
rect 467 2916 468 2920
rect 462 2915 468 2916
rect 464 2899 466 2915
rect 111 2898 115 2899
rect 111 2893 115 2894
rect 311 2898 315 2899
rect 311 2893 315 2894
rect 431 2898 435 2899
rect 431 2893 435 2894
rect 463 2898 467 2899
rect 463 2893 467 2894
rect 112 2874 114 2893
rect 312 2877 314 2893
rect 432 2877 434 2893
rect 310 2876 316 2877
rect 110 2873 116 2874
rect 110 2869 111 2873
rect 115 2869 116 2873
rect 310 2872 311 2876
rect 315 2872 316 2876
rect 310 2871 316 2872
rect 430 2876 436 2877
rect 430 2872 431 2876
rect 435 2872 436 2876
rect 430 2871 436 2872
rect 110 2868 116 2869
rect 378 2867 384 2868
rect 378 2863 379 2867
rect 383 2863 384 2867
rect 378 2862 384 2863
rect 430 2863 436 2864
rect 110 2856 116 2857
rect 110 2852 111 2856
rect 115 2852 116 2856
rect 110 2851 116 2852
rect 112 2823 114 2851
rect 318 2838 324 2839
rect 318 2834 319 2838
rect 323 2834 324 2838
rect 318 2833 324 2834
rect 327 2836 331 2837
rect 320 2823 322 2833
rect 327 2831 331 2832
rect 328 2828 330 2831
rect 380 2828 382 2862
rect 430 2859 431 2863
rect 435 2859 436 2863
rect 430 2858 436 2859
rect 326 2827 332 2828
rect 326 2823 327 2827
rect 331 2823 332 2827
rect 111 2822 115 2823
rect 111 2817 115 2818
rect 167 2822 171 2823
rect 167 2817 171 2818
rect 303 2822 307 2823
rect 303 2817 307 2818
rect 319 2822 323 2823
rect 326 2822 332 2823
rect 378 2827 384 2828
rect 378 2823 379 2827
rect 383 2823 384 2827
rect 378 2822 384 2823
rect 319 2817 323 2818
rect 112 2789 114 2817
rect 168 2807 170 2817
rect 210 2815 216 2816
rect 210 2811 211 2815
rect 215 2811 216 2815
rect 210 2810 216 2811
rect 218 2815 224 2816
rect 218 2811 219 2815
rect 223 2811 224 2815
rect 218 2810 224 2811
rect 166 2806 172 2807
rect 166 2802 167 2806
rect 171 2802 172 2806
rect 166 2801 172 2802
rect 110 2788 116 2789
rect 110 2784 111 2788
rect 115 2784 116 2788
rect 110 2783 116 2784
rect 110 2771 116 2772
rect 110 2767 111 2771
rect 115 2767 116 2771
rect 110 2766 116 2767
rect 158 2768 164 2769
rect 112 2743 114 2766
rect 158 2764 159 2768
rect 163 2764 164 2768
rect 158 2763 164 2764
rect 160 2743 162 2763
rect 212 2752 214 2810
rect 220 2780 222 2810
rect 304 2807 306 2817
rect 432 2816 434 2858
rect 438 2838 444 2839
rect 438 2834 439 2838
rect 443 2834 444 2838
rect 438 2833 444 2834
rect 440 2823 442 2833
rect 524 2828 526 2926
rect 566 2920 572 2921
rect 566 2916 567 2920
rect 571 2916 572 2920
rect 566 2915 572 2916
rect 678 2920 684 2921
rect 678 2916 679 2920
rect 683 2916 684 2920
rect 678 2915 684 2916
rect 798 2920 804 2921
rect 798 2916 799 2920
rect 803 2916 804 2920
rect 798 2915 804 2916
rect 934 2920 940 2921
rect 934 2916 935 2920
rect 939 2916 940 2920
rect 934 2915 940 2916
rect 1078 2920 1084 2921
rect 1078 2916 1079 2920
rect 1083 2916 1084 2920
rect 1078 2915 1084 2916
rect 1238 2920 1244 2921
rect 1238 2916 1239 2920
rect 1243 2916 1244 2920
rect 1238 2915 1244 2916
rect 568 2899 570 2915
rect 680 2899 682 2915
rect 800 2899 802 2915
rect 936 2899 938 2915
rect 1080 2899 1082 2915
rect 1240 2899 1242 2915
rect 551 2898 555 2899
rect 551 2893 555 2894
rect 567 2898 571 2899
rect 567 2893 571 2894
rect 679 2898 683 2899
rect 679 2893 683 2894
rect 799 2898 803 2899
rect 799 2893 803 2894
rect 815 2898 819 2899
rect 815 2893 819 2894
rect 935 2898 939 2899
rect 935 2893 939 2894
rect 951 2898 955 2899
rect 951 2893 955 2894
rect 1079 2898 1083 2899
rect 1079 2893 1083 2894
rect 1087 2898 1091 2899
rect 1087 2893 1091 2894
rect 1223 2898 1227 2899
rect 1223 2893 1227 2894
rect 1239 2898 1243 2899
rect 1239 2893 1243 2894
rect 552 2877 554 2893
rect 680 2877 682 2893
rect 816 2877 818 2893
rect 952 2877 954 2893
rect 1088 2877 1090 2893
rect 1224 2877 1226 2893
rect 550 2876 556 2877
rect 550 2872 551 2876
rect 555 2872 556 2876
rect 550 2871 556 2872
rect 678 2876 684 2877
rect 678 2872 679 2876
rect 683 2872 684 2876
rect 678 2871 684 2872
rect 814 2876 820 2877
rect 814 2872 815 2876
rect 819 2872 820 2876
rect 814 2871 820 2872
rect 950 2876 956 2877
rect 950 2872 951 2876
rect 955 2872 956 2876
rect 950 2871 956 2872
rect 1086 2876 1092 2877
rect 1086 2872 1087 2876
rect 1091 2872 1092 2876
rect 1086 2871 1092 2872
rect 1222 2876 1228 2877
rect 1222 2872 1223 2876
rect 1227 2872 1228 2876
rect 1222 2871 1228 2872
rect 1308 2868 1310 2943
rect 1468 2932 1470 2962
rect 1592 2959 1594 2969
rect 1590 2958 1596 2959
rect 1590 2954 1591 2958
rect 1595 2954 1596 2958
rect 1590 2953 1596 2954
rect 1600 2932 1602 2974
rect 1751 2969 1755 2970
rect 1831 2974 1835 2975
rect 1870 2972 1871 2976
rect 1875 2972 1876 2976
rect 1870 2971 1876 2972
rect 1831 2969 1835 2970
rect 1752 2959 1754 2969
rect 1798 2967 1804 2968
rect 1798 2963 1799 2967
rect 1803 2963 1804 2967
rect 1798 2962 1804 2963
rect 1750 2958 1756 2959
rect 1750 2954 1751 2958
rect 1755 2954 1756 2958
rect 1750 2953 1756 2954
rect 1466 2931 1472 2932
rect 1466 2927 1467 2931
rect 1471 2927 1472 2931
rect 1466 2926 1472 2927
rect 1598 2931 1604 2932
rect 1598 2927 1599 2931
rect 1603 2927 1604 2931
rect 1598 2926 1604 2927
rect 1406 2920 1412 2921
rect 1406 2916 1407 2920
rect 1411 2916 1412 2920
rect 1406 2915 1412 2916
rect 1582 2920 1588 2921
rect 1582 2916 1583 2920
rect 1587 2916 1588 2920
rect 1582 2915 1588 2916
rect 1742 2920 1748 2921
rect 1742 2916 1743 2920
rect 1747 2916 1748 2920
rect 1742 2915 1748 2916
rect 1408 2899 1410 2915
rect 1584 2899 1586 2915
rect 1744 2899 1746 2915
rect 1758 2903 1764 2904
rect 1758 2899 1759 2903
rect 1763 2899 1764 2903
rect 1800 2900 1802 2962
rect 1832 2941 1834 2969
rect 1872 2943 1874 2971
rect 1871 2942 1875 2943
rect 1830 2940 1836 2941
rect 1830 2936 1831 2940
rect 1835 2936 1836 2940
rect 1871 2937 1875 2938
rect 1830 2935 1836 2936
rect 1830 2923 1836 2924
rect 1830 2919 1831 2923
rect 1835 2919 1836 2923
rect 1830 2918 1836 2919
rect 1359 2898 1363 2899
rect 1359 2893 1363 2894
rect 1407 2898 1411 2899
rect 1407 2893 1411 2894
rect 1495 2898 1499 2899
rect 1495 2893 1499 2894
rect 1583 2898 1587 2899
rect 1583 2893 1587 2894
rect 1631 2898 1635 2899
rect 1631 2893 1635 2894
rect 1743 2898 1747 2899
rect 1758 2898 1764 2899
rect 1798 2899 1804 2900
rect 1832 2899 1834 2918
rect 1872 2909 1874 2937
rect 1896 2936 1898 2978
rect 1902 2958 1908 2959
rect 1902 2954 1903 2958
rect 1907 2954 1908 2958
rect 1902 2953 1908 2954
rect 1904 2943 1906 2953
rect 1964 2948 1966 2982
rect 2040 2948 2042 3054
rect 2182 3048 2188 3049
rect 2182 3044 2183 3048
rect 2187 3044 2188 3048
rect 2182 3043 2188 3044
rect 2184 3019 2186 3043
rect 2047 3018 2051 3019
rect 2047 3013 2051 3014
rect 2183 3018 2187 3019
rect 2183 3013 2187 3014
rect 2223 3018 2227 3019
rect 2223 3013 2227 3014
rect 2048 2997 2050 3013
rect 2224 2997 2226 3013
rect 2046 2996 2052 2997
rect 2046 2992 2047 2996
rect 2051 2992 2052 2996
rect 2046 2991 2052 2992
rect 2222 2996 2228 2997
rect 2222 2992 2223 2996
rect 2227 2992 2228 2996
rect 2222 2991 2228 2992
rect 2348 2988 2350 3090
rect 2408 3087 2410 3097
rect 2416 3093 2418 3118
rect 2520 3103 2522 3129
rect 2552 3124 2554 3198
rect 2680 3195 2682 3215
rect 2816 3195 2818 3215
rect 2952 3195 2954 3215
rect 3088 3195 3090 3215
rect 3224 3195 3226 3215
rect 2639 3194 2643 3195
rect 2639 3189 2643 3190
rect 2679 3194 2683 3195
rect 2679 3189 2683 3190
rect 2767 3194 2771 3195
rect 2767 3189 2771 3190
rect 2815 3194 2819 3195
rect 2815 3189 2819 3190
rect 2895 3194 2899 3195
rect 2895 3189 2899 3190
rect 2951 3194 2955 3195
rect 2951 3189 2955 3190
rect 3031 3194 3035 3195
rect 3031 3189 3035 3190
rect 3087 3194 3091 3195
rect 3087 3189 3091 3190
rect 3175 3194 3179 3195
rect 3175 3189 3179 3190
rect 3223 3194 3227 3195
rect 3223 3189 3227 3190
rect 2640 3173 2642 3189
rect 2768 3173 2770 3189
rect 2896 3173 2898 3189
rect 3032 3173 3034 3189
rect 3176 3173 3178 3189
rect 2638 3172 2644 3173
rect 2638 3168 2639 3172
rect 2643 3168 2644 3172
rect 2638 3167 2644 3168
rect 2766 3172 2772 3173
rect 2766 3168 2767 3172
rect 2771 3168 2772 3172
rect 2766 3167 2772 3168
rect 2894 3172 2900 3173
rect 2894 3168 2895 3172
rect 2899 3168 2900 3172
rect 2894 3167 2900 3168
rect 3030 3172 3036 3173
rect 3030 3168 3031 3172
rect 3035 3168 3036 3172
rect 3030 3167 3036 3168
rect 3174 3172 3180 3173
rect 3174 3168 3175 3172
rect 3179 3168 3180 3172
rect 3174 3167 3180 3168
rect 3268 3164 3270 3262
rect 3376 3259 3378 3269
rect 3434 3267 3440 3268
rect 3434 3263 3435 3267
rect 3439 3263 3440 3267
rect 3434 3262 3440 3263
rect 3374 3258 3380 3259
rect 3374 3254 3375 3258
rect 3379 3254 3380 3258
rect 3374 3253 3380 3254
rect 3436 3232 3438 3262
rect 3512 3259 3514 3269
rect 3532 3268 3534 3318
rect 3590 3316 3591 3320
rect 3595 3316 3596 3320
rect 3590 3315 3596 3316
rect 3592 3275 3594 3315
rect 3591 3274 3595 3275
rect 3591 3269 3595 3270
rect 3530 3267 3536 3268
rect 3530 3263 3531 3267
rect 3535 3263 3536 3267
rect 3530 3262 3536 3263
rect 3510 3258 3516 3259
rect 3510 3254 3511 3258
rect 3515 3254 3516 3258
rect 3510 3253 3516 3254
rect 3592 3241 3594 3269
rect 3590 3240 3596 3241
rect 3590 3236 3591 3240
rect 3595 3236 3596 3240
rect 3590 3235 3596 3236
rect 3426 3231 3432 3232
rect 3426 3227 3427 3231
rect 3431 3227 3432 3231
rect 3426 3226 3432 3227
rect 3434 3231 3440 3232
rect 3434 3227 3435 3231
rect 3439 3227 3440 3231
rect 3434 3226 3440 3227
rect 3366 3220 3372 3221
rect 3366 3216 3367 3220
rect 3371 3216 3372 3220
rect 3366 3215 3372 3216
rect 3368 3195 3370 3215
rect 3327 3194 3331 3195
rect 3327 3189 3331 3190
rect 3367 3194 3371 3195
rect 3367 3189 3371 3190
rect 3328 3173 3330 3189
rect 3326 3172 3332 3173
rect 3326 3168 3327 3172
rect 3331 3168 3332 3172
rect 3326 3167 3332 3168
rect 2582 3163 2588 3164
rect 2582 3159 2583 3163
rect 2587 3159 2588 3163
rect 2582 3158 2588 3159
rect 2710 3163 2716 3164
rect 2710 3159 2711 3163
rect 2715 3159 2716 3163
rect 2710 3158 2716 3159
rect 2838 3163 2844 3164
rect 2838 3159 2839 3163
rect 2843 3159 2844 3163
rect 2838 3158 2844 3159
rect 2970 3163 2976 3164
rect 2970 3159 2971 3163
rect 2975 3159 2976 3163
rect 2970 3158 2976 3159
rect 3098 3163 3104 3164
rect 3098 3159 3099 3163
rect 3103 3159 3104 3163
rect 3098 3158 3104 3159
rect 3258 3163 3264 3164
rect 3258 3159 3259 3163
rect 3263 3159 3264 3163
rect 3258 3158 3264 3159
rect 3266 3163 3272 3164
rect 3266 3159 3267 3163
rect 3271 3159 3272 3163
rect 3266 3158 3272 3159
rect 2584 3124 2586 3158
rect 2646 3134 2652 3135
rect 2646 3130 2647 3134
rect 2651 3130 2652 3134
rect 2646 3129 2652 3130
rect 2550 3123 2556 3124
rect 2550 3119 2551 3123
rect 2555 3119 2556 3123
rect 2550 3118 2556 3119
rect 2582 3123 2588 3124
rect 2582 3119 2583 3123
rect 2587 3119 2588 3123
rect 2582 3118 2588 3119
rect 2648 3103 2650 3129
rect 2712 3124 2714 3158
rect 2774 3134 2780 3135
rect 2774 3130 2775 3134
rect 2779 3130 2780 3134
rect 2774 3129 2780 3130
rect 2710 3123 2716 3124
rect 2710 3119 2711 3123
rect 2715 3119 2716 3123
rect 2710 3118 2716 3119
rect 2776 3103 2778 3129
rect 2840 3124 2842 3158
rect 2902 3134 2908 3135
rect 2902 3130 2903 3134
rect 2907 3130 2908 3134
rect 2902 3129 2908 3130
rect 2838 3123 2844 3124
rect 2838 3119 2839 3123
rect 2843 3119 2844 3123
rect 2838 3118 2844 3119
rect 2904 3103 2906 3129
rect 2972 3124 2974 3158
rect 3038 3134 3044 3135
rect 3038 3130 3039 3134
rect 3043 3130 3044 3134
rect 3038 3129 3044 3130
rect 2970 3123 2976 3124
rect 2970 3119 2971 3123
rect 2975 3119 2976 3123
rect 2970 3118 2976 3119
rect 3040 3103 3042 3129
rect 3100 3124 3102 3158
rect 3238 3155 3244 3156
rect 3238 3151 3239 3155
rect 3243 3151 3244 3155
rect 3238 3150 3244 3151
rect 3182 3134 3188 3135
rect 3182 3130 3183 3134
rect 3187 3130 3188 3134
rect 3182 3129 3188 3130
rect 3098 3123 3104 3124
rect 3098 3119 3099 3123
rect 3103 3119 3104 3123
rect 3098 3118 3104 3119
rect 3184 3103 3186 3129
rect 2519 3102 2523 3103
rect 2519 3097 2523 3098
rect 2647 3102 2651 3103
rect 2647 3097 2651 3098
rect 2655 3102 2659 3103
rect 2655 3097 2659 3098
rect 2775 3102 2779 3103
rect 2775 3097 2779 3098
rect 2903 3102 2907 3103
rect 2903 3097 2907 3098
rect 2935 3102 2939 3103
rect 2935 3097 2939 3098
rect 3039 3102 3043 3103
rect 3039 3097 3043 3098
rect 3183 3102 3187 3103
rect 3183 3097 3187 3098
rect 3231 3102 3235 3103
rect 3231 3097 3235 3098
rect 2458 3095 2464 3096
rect 2415 3092 2419 3093
rect 2458 3091 2459 3095
rect 2463 3091 2464 3095
rect 2458 3090 2464 3091
rect 2415 3087 2419 3088
rect 2406 3086 2412 3087
rect 2406 3082 2407 3086
rect 2411 3082 2412 3086
rect 2406 3081 2412 3082
rect 2460 3060 2462 3090
rect 2656 3087 2658 3097
rect 2706 3095 2712 3096
rect 2706 3091 2707 3095
rect 2711 3091 2712 3095
rect 2706 3090 2712 3091
rect 2654 3086 2660 3087
rect 2654 3082 2655 3086
rect 2659 3082 2660 3086
rect 2654 3081 2660 3082
rect 2708 3060 2710 3090
rect 2936 3087 2938 3097
rect 2943 3092 2947 3093
rect 2943 3087 2947 3088
rect 3232 3087 3234 3097
rect 3240 3096 3242 3150
rect 3260 3124 3262 3158
rect 3334 3134 3340 3135
rect 3334 3130 3335 3134
rect 3339 3130 3340 3134
rect 3334 3129 3340 3130
rect 3258 3123 3264 3124
rect 3258 3119 3259 3123
rect 3263 3119 3264 3123
rect 3258 3118 3264 3119
rect 3336 3103 3338 3129
rect 3428 3124 3430 3226
rect 3590 3223 3596 3224
rect 3502 3220 3508 3221
rect 3502 3216 3503 3220
rect 3507 3216 3508 3220
rect 3590 3219 3591 3223
rect 3595 3219 3596 3223
rect 3590 3218 3596 3219
rect 3502 3215 3508 3216
rect 3504 3195 3506 3215
rect 3592 3195 3594 3218
rect 3487 3194 3491 3195
rect 3487 3189 3491 3190
rect 3503 3194 3507 3195
rect 3503 3189 3507 3190
rect 3591 3194 3595 3195
rect 3591 3189 3595 3190
rect 3488 3173 3490 3189
rect 3486 3172 3492 3173
rect 3486 3168 3487 3172
rect 3491 3168 3492 3172
rect 3592 3170 3594 3189
rect 3486 3167 3492 3168
rect 3590 3169 3596 3170
rect 3590 3165 3591 3169
rect 3595 3165 3596 3169
rect 3590 3164 3596 3165
rect 3590 3152 3596 3153
rect 3590 3148 3591 3152
rect 3595 3148 3596 3152
rect 3590 3147 3596 3148
rect 3494 3134 3500 3135
rect 3494 3130 3495 3134
rect 3499 3130 3500 3134
rect 3494 3129 3500 3130
rect 3426 3123 3432 3124
rect 3426 3119 3427 3123
rect 3431 3119 3432 3123
rect 3426 3118 3432 3119
rect 3496 3103 3498 3129
rect 3592 3103 3594 3147
rect 3335 3102 3339 3103
rect 3335 3097 3339 3098
rect 3495 3102 3499 3103
rect 3495 3097 3499 3098
rect 3511 3102 3515 3103
rect 3511 3097 3515 3098
rect 3591 3102 3595 3103
rect 3591 3097 3595 3098
rect 3238 3095 3244 3096
rect 3238 3091 3239 3095
rect 3243 3091 3244 3095
rect 3238 3090 3244 3091
rect 3282 3095 3288 3096
rect 3282 3091 3283 3095
rect 3287 3091 3288 3095
rect 3282 3090 3288 3091
rect 2934 3086 2940 3087
rect 2934 3082 2935 3086
rect 2939 3082 2940 3086
rect 2934 3081 2940 3082
rect 2944 3060 2946 3087
rect 3230 3086 3236 3087
rect 3230 3082 3231 3086
rect 3235 3082 3236 3086
rect 3230 3081 3236 3082
rect 3284 3060 3286 3090
rect 3512 3087 3514 3097
rect 3510 3086 3516 3087
rect 3510 3082 3511 3086
rect 3515 3082 3516 3086
rect 3510 3081 3516 3082
rect 3592 3069 3594 3097
rect 3590 3068 3596 3069
rect 3590 3064 3591 3068
rect 3595 3064 3596 3068
rect 3590 3063 3596 3064
rect 2458 3059 2464 3060
rect 2458 3055 2459 3059
rect 2463 3055 2464 3059
rect 2458 3054 2464 3055
rect 2706 3059 2712 3060
rect 2706 3055 2707 3059
rect 2711 3055 2712 3059
rect 2706 3054 2712 3055
rect 2942 3059 2948 3060
rect 2942 3055 2943 3059
rect 2947 3055 2948 3059
rect 2942 3054 2948 3055
rect 3282 3059 3288 3060
rect 3282 3055 3283 3059
rect 3287 3055 3288 3059
rect 3282 3054 3288 3055
rect 3590 3051 3596 3052
rect 2398 3048 2404 3049
rect 2398 3044 2399 3048
rect 2403 3044 2404 3048
rect 2398 3043 2404 3044
rect 2646 3048 2652 3049
rect 2646 3044 2647 3048
rect 2651 3044 2652 3048
rect 2646 3043 2652 3044
rect 2926 3048 2932 3049
rect 2926 3044 2927 3048
rect 2931 3044 2932 3048
rect 2926 3043 2932 3044
rect 3222 3048 3228 3049
rect 3222 3044 3223 3048
rect 3227 3044 3228 3048
rect 3222 3043 3228 3044
rect 3502 3048 3508 3049
rect 3502 3044 3503 3048
rect 3507 3044 3508 3048
rect 3590 3047 3591 3051
rect 3595 3047 3596 3051
rect 3590 3046 3596 3047
rect 3502 3043 3508 3044
rect 2400 3019 2402 3043
rect 2648 3019 2650 3043
rect 2928 3019 2930 3043
rect 3224 3019 3226 3043
rect 3504 3019 3506 3043
rect 3518 3031 3524 3032
rect 3518 3027 3519 3031
rect 3523 3027 3524 3031
rect 3518 3026 3524 3027
rect 2391 3018 2395 3019
rect 2391 3013 2395 3014
rect 2399 3018 2403 3019
rect 2399 3013 2403 3014
rect 2543 3018 2547 3019
rect 2543 3013 2547 3014
rect 2647 3018 2651 3019
rect 2647 3013 2651 3014
rect 2687 3018 2691 3019
rect 2687 3013 2691 3014
rect 2815 3018 2819 3019
rect 2815 3013 2819 3014
rect 2927 3018 2931 3019
rect 2927 3013 2931 3014
rect 3039 3018 3043 3019
rect 3039 3013 3043 3014
rect 3143 3018 3147 3019
rect 3143 3013 3147 3014
rect 3223 3018 3227 3019
rect 3223 3013 3227 3014
rect 3239 3018 3243 3019
rect 3239 3013 3243 3014
rect 3335 3018 3339 3019
rect 3335 3013 3339 3014
rect 3423 3018 3427 3019
rect 3423 3013 3427 3014
rect 3503 3018 3507 3019
rect 3503 3013 3507 3014
rect 2392 2997 2394 3013
rect 2544 2997 2546 3013
rect 2688 2997 2690 3013
rect 2816 2997 2818 3013
rect 2928 2997 2930 3013
rect 3040 2997 3042 3013
rect 3144 2997 3146 3013
rect 3240 2997 3242 3013
rect 3336 2997 3338 3013
rect 3424 2997 3426 3013
rect 3504 2997 3506 3013
rect 2390 2996 2396 2997
rect 2390 2992 2391 2996
rect 2395 2992 2396 2996
rect 2390 2991 2396 2992
rect 2542 2996 2548 2997
rect 2542 2992 2543 2996
rect 2547 2992 2548 2996
rect 2542 2991 2548 2992
rect 2686 2996 2692 2997
rect 2686 2992 2687 2996
rect 2691 2992 2692 2996
rect 2686 2991 2692 2992
rect 2814 2996 2820 2997
rect 2814 2992 2815 2996
rect 2819 2992 2820 2996
rect 2814 2991 2820 2992
rect 2926 2996 2932 2997
rect 2926 2992 2927 2996
rect 2931 2992 2932 2996
rect 2926 2991 2932 2992
rect 3038 2996 3044 2997
rect 3038 2992 3039 2996
rect 3043 2992 3044 2996
rect 3038 2991 3044 2992
rect 3142 2996 3148 2997
rect 3142 2992 3143 2996
rect 3147 2992 3148 2996
rect 3142 2991 3148 2992
rect 3238 2996 3244 2997
rect 3238 2992 3239 2996
rect 3243 2992 3244 2996
rect 3238 2991 3244 2992
rect 3334 2996 3340 2997
rect 3334 2992 3335 2996
rect 3339 2992 3340 2996
rect 3334 2991 3340 2992
rect 3422 2996 3428 2997
rect 3422 2992 3423 2996
rect 3427 2992 3428 2996
rect 3422 2991 3428 2992
rect 3502 2996 3508 2997
rect 3502 2992 3503 2996
rect 3507 2992 3508 2996
rect 3502 2991 3508 2992
rect 2346 2987 2352 2988
rect 2346 2983 2347 2987
rect 2351 2983 2352 2987
rect 2346 2982 2352 2983
rect 2354 2987 2360 2988
rect 2354 2983 2355 2987
rect 2359 2983 2360 2987
rect 2354 2982 2360 2983
rect 2610 2987 2616 2988
rect 2610 2983 2611 2987
rect 2615 2983 2616 2987
rect 2610 2982 2616 2983
rect 2758 2987 2764 2988
rect 2758 2983 2759 2987
rect 2763 2983 2764 2987
rect 2758 2982 2764 2983
rect 2910 2987 2916 2988
rect 2910 2983 2911 2987
rect 2915 2983 2916 2987
rect 2910 2982 2916 2983
rect 2918 2987 2924 2988
rect 2918 2983 2919 2987
rect 2923 2983 2924 2987
rect 2918 2982 2924 2983
rect 3106 2987 3112 2988
rect 3106 2983 3107 2987
rect 3111 2983 3112 2987
rect 3106 2982 3112 2983
rect 3210 2987 3216 2988
rect 3210 2983 3211 2987
rect 3215 2983 3216 2987
rect 3210 2982 3216 2983
rect 3402 2987 3408 2988
rect 3402 2983 3403 2987
rect 3407 2983 3408 2987
rect 3490 2987 3496 2988
rect 3402 2982 3408 2983
rect 3422 2983 3428 2984
rect 2054 2958 2060 2959
rect 2054 2954 2055 2958
rect 2059 2954 2060 2958
rect 2054 2953 2060 2954
rect 2230 2958 2236 2959
rect 2230 2954 2231 2958
rect 2235 2954 2236 2958
rect 2230 2953 2236 2954
rect 1962 2947 1968 2948
rect 1962 2943 1963 2947
rect 1967 2943 1968 2947
rect 1903 2942 1907 2943
rect 1962 2942 1968 2943
rect 2038 2947 2044 2948
rect 2038 2943 2039 2947
rect 2043 2943 2044 2947
rect 2056 2943 2058 2953
rect 2232 2943 2234 2953
rect 2356 2948 2358 2982
rect 2398 2958 2404 2959
rect 2398 2954 2399 2958
rect 2403 2954 2404 2958
rect 2398 2953 2404 2954
rect 2550 2958 2556 2959
rect 2550 2954 2551 2958
rect 2555 2954 2556 2958
rect 2550 2953 2556 2954
rect 2567 2956 2571 2957
rect 2354 2947 2360 2948
rect 2354 2943 2355 2947
rect 2359 2943 2360 2947
rect 2400 2943 2402 2953
rect 2494 2947 2500 2948
rect 2494 2943 2495 2947
rect 2499 2943 2500 2947
rect 2552 2943 2554 2953
rect 2567 2951 2571 2952
rect 2568 2948 2570 2951
rect 2612 2948 2614 2982
rect 2694 2958 2700 2959
rect 2694 2954 2695 2958
rect 2699 2954 2700 2958
rect 2694 2953 2700 2954
rect 2566 2947 2572 2948
rect 2566 2943 2567 2947
rect 2571 2943 2572 2947
rect 2038 2942 2044 2943
rect 2055 2942 2059 2943
rect 1903 2937 1907 2938
rect 2055 2937 2059 2938
rect 2087 2942 2091 2943
rect 2087 2937 2091 2938
rect 2231 2942 2235 2943
rect 2231 2937 2235 2938
rect 2295 2942 2299 2943
rect 2354 2942 2360 2943
rect 2399 2942 2403 2943
rect 2295 2937 2299 2938
rect 2399 2937 2403 2938
rect 2487 2942 2491 2943
rect 2494 2942 2500 2943
rect 2551 2942 2555 2943
rect 2566 2942 2572 2943
rect 2610 2947 2616 2948
rect 2610 2943 2611 2947
rect 2615 2943 2616 2947
rect 2696 2943 2698 2953
rect 2760 2948 2762 2982
rect 2822 2958 2828 2959
rect 2822 2954 2823 2958
rect 2827 2954 2828 2958
rect 2822 2953 2828 2954
rect 2758 2947 2764 2948
rect 2758 2943 2759 2947
rect 2763 2943 2764 2947
rect 2824 2943 2826 2953
rect 2610 2942 2616 2943
rect 2671 2942 2675 2943
rect 2487 2937 2491 2938
rect 1894 2935 1900 2936
rect 1894 2931 1895 2935
rect 1899 2931 1900 2935
rect 1894 2930 1900 2931
rect 1904 2927 1906 2937
rect 2088 2927 2090 2937
rect 2094 2935 2100 2936
rect 2094 2931 2095 2935
rect 2099 2931 2100 2935
rect 2094 2930 2100 2931
rect 2138 2935 2144 2936
rect 2138 2931 2139 2935
rect 2143 2931 2144 2935
rect 2138 2930 2144 2931
rect 1902 2926 1908 2927
rect 1902 2922 1903 2926
rect 1907 2922 1908 2926
rect 1902 2921 1908 2922
rect 2086 2926 2092 2927
rect 2086 2922 2087 2926
rect 2091 2922 2092 2926
rect 2086 2921 2092 2922
rect 1870 2908 1876 2909
rect 1870 2904 1871 2908
rect 1875 2904 1876 2908
rect 1870 2903 1876 2904
rect 1743 2893 1747 2894
rect 1360 2877 1362 2893
rect 1496 2877 1498 2893
rect 1632 2877 1634 2893
rect 1744 2877 1746 2893
rect 1358 2876 1364 2877
rect 1358 2872 1359 2876
rect 1363 2872 1364 2876
rect 1358 2871 1364 2872
rect 1494 2876 1500 2877
rect 1494 2872 1495 2876
rect 1499 2872 1500 2876
rect 1494 2871 1500 2872
rect 1630 2876 1636 2877
rect 1630 2872 1631 2876
rect 1635 2872 1636 2876
rect 1630 2871 1636 2872
rect 1742 2876 1748 2877
rect 1742 2872 1743 2876
rect 1747 2872 1748 2876
rect 1742 2871 1748 2872
rect 754 2867 760 2868
rect 754 2863 755 2867
rect 759 2863 760 2867
rect 754 2862 760 2863
rect 762 2867 768 2868
rect 762 2863 763 2867
rect 767 2863 768 2867
rect 762 2862 768 2863
rect 1026 2867 1032 2868
rect 1026 2863 1027 2867
rect 1031 2863 1032 2867
rect 1026 2862 1032 2863
rect 1162 2867 1168 2868
rect 1162 2863 1163 2867
rect 1167 2863 1168 2867
rect 1162 2862 1168 2863
rect 1298 2867 1304 2868
rect 1298 2863 1299 2867
rect 1303 2863 1304 2867
rect 1298 2862 1304 2863
rect 1306 2867 1312 2868
rect 1306 2863 1307 2867
rect 1311 2863 1312 2867
rect 1306 2862 1312 2863
rect 1562 2867 1568 2868
rect 1562 2863 1563 2867
rect 1567 2863 1568 2867
rect 1562 2862 1568 2863
rect 1698 2867 1704 2868
rect 1698 2863 1699 2867
rect 1703 2863 1704 2867
rect 1698 2862 1704 2863
rect 558 2838 564 2839
rect 558 2834 559 2838
rect 563 2834 564 2838
rect 558 2833 564 2834
rect 686 2838 692 2839
rect 686 2834 687 2838
rect 691 2834 692 2838
rect 686 2833 692 2834
rect 522 2827 528 2828
rect 522 2823 523 2827
rect 527 2823 528 2827
rect 560 2823 562 2833
rect 688 2823 690 2833
rect 756 2828 758 2862
rect 764 2837 766 2862
rect 822 2838 828 2839
rect 763 2836 767 2837
rect 822 2834 823 2838
rect 827 2834 828 2838
rect 822 2833 828 2834
rect 958 2838 964 2839
rect 958 2834 959 2838
rect 963 2834 964 2838
rect 958 2833 964 2834
rect 763 2831 767 2832
rect 754 2827 760 2828
rect 754 2823 755 2827
rect 759 2823 760 2827
rect 824 2823 826 2833
rect 960 2823 962 2833
rect 1028 2828 1030 2862
rect 1094 2838 1100 2839
rect 1094 2834 1095 2838
rect 1099 2834 1100 2838
rect 1094 2833 1100 2834
rect 966 2827 972 2828
rect 966 2823 967 2827
rect 971 2823 972 2827
rect 439 2822 443 2823
rect 439 2817 443 2818
rect 447 2822 451 2823
rect 522 2822 528 2823
rect 559 2822 563 2823
rect 447 2817 451 2818
rect 559 2817 563 2818
rect 607 2822 611 2823
rect 607 2817 611 2818
rect 687 2822 691 2823
rect 754 2822 760 2823
rect 783 2822 787 2823
rect 687 2817 691 2818
rect 783 2817 787 2818
rect 823 2822 827 2823
rect 823 2817 827 2818
rect 959 2822 963 2823
rect 966 2822 972 2823
rect 1026 2827 1032 2828
rect 1026 2823 1027 2827
rect 1031 2823 1032 2827
rect 1096 2823 1098 2833
rect 1164 2828 1166 2862
rect 1230 2838 1236 2839
rect 1230 2834 1231 2838
rect 1235 2834 1236 2838
rect 1230 2833 1236 2834
rect 1162 2827 1168 2828
rect 1162 2823 1163 2827
rect 1167 2823 1168 2827
rect 1232 2823 1234 2833
rect 1300 2828 1302 2862
rect 1554 2859 1560 2860
rect 1554 2855 1555 2859
rect 1559 2855 1560 2859
rect 1554 2854 1560 2855
rect 1366 2838 1372 2839
rect 1366 2834 1367 2838
rect 1371 2834 1372 2838
rect 1366 2833 1372 2834
rect 1502 2838 1508 2839
rect 1502 2834 1503 2838
rect 1507 2834 1508 2838
rect 1502 2833 1508 2834
rect 1298 2827 1304 2828
rect 1298 2823 1299 2827
rect 1303 2823 1304 2827
rect 1368 2823 1370 2833
rect 1504 2823 1506 2833
rect 1026 2822 1032 2823
rect 1095 2822 1099 2823
rect 959 2817 963 2818
rect 430 2815 436 2816
rect 430 2811 431 2815
rect 435 2811 436 2815
rect 430 2810 436 2811
rect 448 2807 450 2817
rect 498 2815 504 2816
rect 498 2811 499 2815
rect 503 2811 504 2815
rect 498 2810 504 2811
rect 302 2806 308 2807
rect 302 2802 303 2806
rect 307 2802 308 2806
rect 302 2801 308 2802
rect 446 2806 452 2807
rect 446 2802 447 2806
rect 451 2802 452 2806
rect 446 2801 452 2802
rect 500 2780 502 2810
rect 608 2807 610 2817
rect 658 2815 664 2816
rect 658 2811 659 2815
rect 663 2811 664 2815
rect 658 2810 664 2811
rect 606 2806 612 2807
rect 606 2802 607 2806
rect 611 2802 612 2806
rect 606 2801 612 2802
rect 660 2780 662 2810
rect 784 2807 786 2817
rect 960 2807 962 2817
rect 782 2806 788 2807
rect 782 2802 783 2806
rect 787 2802 788 2806
rect 782 2801 788 2802
rect 958 2806 964 2807
rect 958 2802 959 2806
rect 963 2802 964 2806
rect 958 2801 964 2802
rect 968 2780 970 2822
rect 1095 2817 1099 2818
rect 1143 2822 1147 2823
rect 1162 2822 1168 2823
rect 1231 2822 1235 2823
rect 1298 2822 1304 2823
rect 1335 2822 1339 2823
rect 1143 2817 1147 2818
rect 1231 2817 1235 2818
rect 1335 2817 1339 2818
rect 1367 2822 1371 2823
rect 1367 2817 1371 2818
rect 1503 2822 1507 2823
rect 1503 2817 1507 2818
rect 1535 2822 1539 2823
rect 1535 2817 1539 2818
rect 1018 2815 1024 2816
rect 1018 2811 1019 2815
rect 1023 2811 1024 2815
rect 1018 2810 1024 2811
rect 1020 2780 1022 2810
rect 1144 2807 1146 2817
rect 1202 2815 1208 2816
rect 1202 2811 1203 2815
rect 1207 2811 1208 2815
rect 1202 2810 1208 2811
rect 1266 2815 1272 2816
rect 1266 2811 1267 2815
rect 1271 2811 1272 2815
rect 1266 2810 1272 2811
rect 1142 2806 1148 2807
rect 1142 2802 1143 2806
rect 1147 2802 1148 2806
rect 1142 2801 1148 2802
rect 1204 2780 1206 2810
rect 218 2779 224 2780
rect 218 2775 219 2779
rect 223 2775 224 2779
rect 218 2774 224 2775
rect 354 2779 360 2780
rect 354 2775 355 2779
rect 359 2775 360 2779
rect 354 2774 360 2775
rect 498 2779 504 2780
rect 498 2775 499 2779
rect 503 2775 504 2779
rect 498 2774 504 2775
rect 658 2779 664 2780
rect 658 2775 659 2779
rect 663 2775 664 2779
rect 658 2774 664 2775
rect 966 2779 972 2780
rect 966 2775 967 2779
rect 971 2775 972 2779
rect 966 2774 972 2775
rect 1018 2779 1024 2780
rect 1018 2775 1019 2779
rect 1023 2775 1024 2779
rect 1018 2774 1024 2775
rect 1202 2779 1208 2780
rect 1202 2775 1203 2779
rect 1207 2775 1208 2779
rect 1202 2774 1208 2775
rect 294 2768 300 2769
rect 294 2764 295 2768
rect 299 2764 300 2768
rect 294 2763 300 2764
rect 210 2751 216 2752
rect 210 2747 211 2751
rect 215 2747 216 2751
rect 210 2746 216 2747
rect 296 2743 298 2763
rect 111 2742 115 2743
rect 111 2737 115 2738
rect 135 2742 139 2743
rect 135 2737 139 2738
rect 159 2742 163 2743
rect 159 2737 163 2738
rect 247 2742 251 2743
rect 247 2737 251 2738
rect 295 2742 299 2743
rect 295 2737 299 2738
rect 112 2718 114 2737
rect 136 2721 138 2737
rect 248 2721 250 2737
rect 134 2720 140 2721
rect 110 2717 116 2718
rect 110 2713 111 2717
rect 115 2713 116 2717
rect 134 2716 135 2720
rect 139 2716 140 2720
rect 134 2715 140 2716
rect 246 2720 252 2721
rect 246 2716 247 2720
rect 251 2716 252 2720
rect 246 2715 252 2716
rect 110 2712 116 2713
rect 202 2711 208 2712
rect 134 2707 140 2708
rect 134 2703 135 2707
rect 139 2703 140 2707
rect 202 2707 203 2711
rect 207 2707 208 2711
rect 202 2706 208 2707
rect 134 2702 140 2703
rect 110 2700 116 2701
rect 110 2696 111 2700
rect 115 2696 116 2700
rect 110 2695 116 2696
rect 112 2667 114 2695
rect 111 2666 115 2667
rect 111 2661 115 2662
rect 112 2633 114 2661
rect 136 2660 138 2702
rect 142 2682 148 2683
rect 142 2678 143 2682
rect 147 2678 148 2682
rect 142 2677 148 2678
rect 144 2667 146 2677
rect 204 2672 206 2706
rect 254 2682 260 2683
rect 254 2678 255 2682
rect 259 2678 260 2682
rect 254 2677 260 2678
rect 202 2671 208 2672
rect 202 2667 203 2671
rect 207 2667 208 2671
rect 256 2667 258 2677
rect 263 2676 267 2677
rect 356 2672 358 2774
rect 438 2768 444 2769
rect 438 2764 439 2768
rect 443 2764 444 2768
rect 438 2763 444 2764
rect 598 2768 604 2769
rect 598 2764 599 2768
rect 603 2764 604 2768
rect 598 2763 604 2764
rect 774 2768 780 2769
rect 774 2764 775 2768
rect 779 2764 780 2768
rect 774 2763 780 2764
rect 950 2768 956 2769
rect 950 2764 951 2768
rect 955 2764 956 2768
rect 950 2763 956 2764
rect 1134 2768 1140 2769
rect 1134 2764 1135 2768
rect 1139 2764 1140 2768
rect 1134 2763 1140 2764
rect 440 2743 442 2763
rect 600 2743 602 2763
rect 776 2743 778 2763
rect 952 2743 954 2763
rect 1136 2743 1138 2763
rect 391 2742 395 2743
rect 391 2737 395 2738
rect 439 2742 443 2743
rect 439 2737 443 2738
rect 551 2742 555 2743
rect 551 2737 555 2738
rect 599 2742 603 2743
rect 599 2737 603 2738
rect 711 2742 715 2743
rect 711 2737 715 2738
rect 775 2742 779 2743
rect 775 2737 779 2738
rect 879 2742 883 2743
rect 879 2737 883 2738
rect 951 2742 955 2743
rect 951 2737 955 2738
rect 1039 2742 1043 2743
rect 1039 2737 1043 2738
rect 1135 2742 1139 2743
rect 1135 2737 1139 2738
rect 1199 2742 1203 2743
rect 1199 2737 1203 2738
rect 392 2721 394 2737
rect 552 2721 554 2737
rect 712 2721 714 2737
rect 880 2721 882 2737
rect 1040 2721 1042 2737
rect 1200 2721 1202 2737
rect 390 2720 396 2721
rect 390 2716 391 2720
rect 395 2716 396 2720
rect 390 2715 396 2716
rect 550 2720 556 2721
rect 550 2716 551 2720
rect 555 2716 556 2720
rect 550 2715 556 2716
rect 710 2720 716 2721
rect 710 2716 711 2720
rect 715 2716 716 2720
rect 710 2715 716 2716
rect 878 2720 884 2721
rect 878 2716 879 2720
rect 883 2716 884 2720
rect 878 2715 884 2716
rect 1038 2720 1044 2721
rect 1038 2716 1039 2720
rect 1043 2716 1044 2720
rect 1038 2715 1044 2716
rect 1198 2720 1204 2721
rect 1198 2716 1199 2720
rect 1203 2716 1204 2720
rect 1198 2715 1204 2716
rect 1268 2712 1270 2810
rect 1336 2807 1338 2817
rect 1536 2807 1538 2817
rect 1556 2816 1558 2854
rect 1564 2828 1566 2862
rect 1638 2838 1644 2839
rect 1638 2834 1639 2838
rect 1643 2834 1644 2838
rect 1638 2833 1644 2834
rect 1562 2827 1568 2828
rect 1562 2823 1563 2827
rect 1567 2823 1568 2827
rect 1640 2823 1642 2833
rect 1700 2828 1702 2862
rect 1750 2838 1756 2839
rect 1750 2834 1751 2838
rect 1755 2834 1756 2838
rect 1750 2833 1756 2834
rect 1698 2827 1704 2828
rect 1698 2823 1699 2827
rect 1703 2823 1704 2827
rect 1752 2823 1754 2833
rect 1760 2828 1762 2898
rect 1798 2895 1799 2899
rect 1803 2895 1804 2899
rect 1798 2894 1804 2895
rect 1831 2898 1835 2899
rect 1831 2893 1835 2894
rect 1832 2874 1834 2893
rect 1870 2891 1876 2892
rect 1870 2887 1871 2891
rect 1875 2887 1876 2891
rect 1870 2886 1876 2887
rect 1894 2888 1900 2889
rect 1830 2873 1836 2874
rect 1830 2869 1831 2873
rect 1835 2869 1836 2873
rect 1830 2868 1836 2869
rect 1872 2859 1874 2886
rect 1894 2884 1895 2888
rect 1899 2884 1900 2888
rect 1894 2883 1900 2884
rect 2078 2888 2084 2889
rect 2078 2884 2079 2888
rect 2083 2884 2084 2888
rect 2078 2883 2084 2884
rect 1896 2859 1898 2883
rect 2080 2859 2082 2883
rect 1871 2858 1875 2859
rect 1830 2856 1836 2857
rect 1830 2852 1831 2856
rect 1835 2852 1836 2856
rect 1871 2853 1875 2854
rect 1895 2858 1899 2859
rect 1895 2853 1899 2854
rect 2079 2858 2083 2859
rect 2079 2853 2083 2854
rect 1830 2851 1836 2852
rect 1758 2827 1764 2828
rect 1758 2823 1759 2827
rect 1763 2823 1764 2827
rect 1832 2823 1834 2851
rect 1872 2834 1874 2853
rect 1870 2833 1876 2834
rect 1870 2829 1871 2833
rect 1875 2829 1876 2833
rect 1870 2828 1876 2829
rect 2096 2828 2098 2930
rect 2140 2900 2142 2930
rect 2296 2927 2298 2937
rect 2346 2935 2352 2936
rect 2346 2931 2347 2935
rect 2351 2931 2352 2935
rect 2346 2930 2352 2931
rect 2294 2926 2300 2927
rect 2294 2922 2295 2926
rect 2299 2922 2300 2926
rect 2294 2921 2300 2922
rect 2348 2900 2350 2930
rect 2488 2927 2490 2937
rect 2486 2926 2492 2927
rect 2486 2922 2487 2926
rect 2491 2922 2492 2926
rect 2486 2921 2492 2922
rect 2496 2900 2498 2942
rect 2551 2937 2555 2938
rect 2671 2937 2675 2938
rect 2695 2942 2699 2943
rect 2758 2942 2764 2943
rect 2823 2942 2827 2943
rect 2695 2937 2699 2938
rect 2823 2937 2827 2938
rect 2839 2942 2843 2943
rect 2839 2937 2843 2938
rect 2672 2927 2674 2937
rect 2714 2935 2720 2936
rect 2714 2930 2715 2935
rect 2719 2930 2720 2935
rect 2722 2935 2728 2936
rect 2722 2931 2723 2935
rect 2727 2931 2728 2935
rect 2722 2930 2728 2931
rect 2715 2927 2719 2928
rect 2670 2926 2676 2927
rect 2670 2922 2671 2926
rect 2675 2922 2676 2926
rect 2670 2921 2676 2922
rect 2724 2900 2726 2930
rect 2840 2927 2842 2937
rect 2912 2936 2914 2982
rect 2920 2957 2922 2982
rect 2934 2958 2940 2959
rect 2919 2956 2923 2957
rect 2934 2954 2935 2958
rect 2939 2954 2940 2958
rect 2934 2953 2940 2954
rect 3046 2958 3052 2959
rect 3046 2954 3047 2958
rect 3051 2954 3052 2958
rect 3046 2953 3052 2954
rect 2919 2951 2923 2952
rect 2936 2943 2938 2953
rect 3048 2943 3050 2953
rect 3108 2948 3110 2982
rect 3150 2958 3156 2959
rect 3150 2954 3151 2958
rect 3155 2954 3156 2958
rect 3150 2953 3156 2954
rect 3106 2947 3112 2948
rect 3106 2943 3107 2947
rect 3111 2943 3112 2947
rect 3152 2943 3154 2953
rect 3212 2948 3214 2982
rect 3394 2967 3400 2968
rect 3394 2963 3395 2967
rect 3399 2963 3400 2967
rect 3394 2962 3400 2963
rect 3246 2958 3252 2959
rect 3246 2954 3247 2958
rect 3251 2954 3252 2958
rect 3246 2953 3252 2954
rect 3342 2958 3348 2959
rect 3342 2954 3343 2958
rect 3347 2954 3348 2958
rect 3342 2953 3348 2954
rect 3210 2947 3216 2948
rect 3210 2943 3211 2947
rect 3215 2943 3216 2947
rect 3248 2943 3250 2953
rect 3344 2943 3346 2953
rect 3396 2948 3398 2962
rect 3404 2948 3406 2982
rect 3422 2979 3423 2983
rect 3427 2979 3428 2983
rect 3490 2983 3491 2987
rect 3495 2983 3496 2987
rect 3490 2982 3496 2983
rect 3422 2978 3428 2979
rect 3394 2947 3400 2948
rect 3394 2943 3395 2947
rect 3399 2943 3400 2947
rect 2935 2942 2939 2943
rect 2935 2937 2939 2938
rect 2999 2942 3003 2943
rect 2999 2937 3003 2938
rect 3047 2942 3051 2943
rect 3106 2942 3112 2943
rect 3151 2942 3155 2943
rect 3210 2942 3216 2943
rect 3247 2942 3251 2943
rect 3047 2937 3051 2938
rect 3151 2937 3155 2938
rect 3247 2937 3251 2938
rect 3303 2942 3307 2943
rect 3303 2937 3307 2938
rect 3343 2942 3347 2943
rect 3394 2942 3400 2943
rect 3402 2947 3408 2948
rect 3402 2943 3403 2947
rect 3407 2943 3408 2947
rect 3402 2942 3408 2943
rect 3343 2937 3347 2938
rect 3362 2939 3368 2940
rect 2910 2935 2916 2936
rect 2910 2931 2911 2935
rect 2915 2931 2916 2935
rect 2910 2930 2916 2931
rect 3000 2927 3002 2937
rect 3098 2935 3104 2936
rect 3098 2931 3099 2935
rect 3103 2931 3104 2935
rect 3098 2930 3104 2931
rect 2838 2926 2844 2927
rect 2838 2922 2839 2926
rect 2843 2922 2844 2926
rect 2838 2921 2844 2922
rect 2998 2926 3004 2927
rect 2998 2922 2999 2926
rect 3003 2922 3004 2926
rect 2998 2921 3004 2922
rect 3100 2900 3102 2930
rect 3152 2927 3154 2937
rect 3202 2935 3208 2936
rect 3202 2931 3203 2935
rect 3207 2931 3208 2935
rect 3202 2930 3208 2931
rect 3150 2926 3156 2927
rect 3150 2922 3151 2926
rect 3155 2922 3156 2926
rect 3150 2921 3156 2922
rect 3204 2900 3206 2930
rect 3304 2927 3306 2937
rect 3362 2935 3363 2939
rect 3367 2935 3368 2939
rect 3424 2936 3426 2978
rect 3492 2968 3494 2982
rect 3490 2967 3496 2968
rect 3490 2963 3491 2967
rect 3495 2963 3496 2967
rect 3490 2962 3496 2963
rect 3430 2958 3436 2959
rect 3430 2954 3431 2958
rect 3435 2954 3436 2958
rect 3430 2953 3436 2954
rect 3510 2958 3516 2959
rect 3510 2954 3511 2958
rect 3515 2954 3516 2958
rect 3510 2953 3516 2954
rect 3432 2943 3434 2953
rect 3512 2943 3514 2953
rect 3520 2948 3522 3026
rect 3592 3019 3594 3046
rect 3591 3018 3595 3019
rect 3591 3013 3595 3014
rect 3592 2994 3594 3013
rect 3590 2993 3596 2994
rect 3590 2989 3591 2993
rect 3595 2989 3596 2993
rect 3590 2988 3596 2989
rect 3590 2976 3596 2977
rect 3590 2972 3591 2976
rect 3595 2972 3596 2976
rect 3590 2971 3596 2972
rect 3518 2947 3524 2948
rect 3518 2943 3519 2947
rect 3523 2943 3524 2947
rect 3592 2943 3594 2971
rect 3431 2942 3435 2943
rect 3431 2937 3435 2938
rect 3455 2942 3459 2943
rect 3455 2937 3459 2938
rect 3511 2942 3515 2943
rect 3518 2942 3524 2943
rect 3591 2942 3595 2943
rect 3511 2937 3515 2938
rect 3591 2937 3595 2938
rect 3362 2934 3368 2935
rect 3422 2935 3428 2936
rect 3311 2932 3315 2933
rect 3311 2927 3315 2928
rect 3302 2926 3308 2927
rect 3302 2922 3303 2926
rect 3307 2922 3308 2926
rect 3302 2921 3308 2922
rect 3312 2900 3314 2927
rect 3364 2900 3366 2934
rect 3422 2931 3423 2935
rect 3427 2931 3428 2935
rect 3422 2930 3428 2931
rect 3456 2927 3458 2937
rect 3454 2926 3460 2927
rect 3454 2922 3455 2926
rect 3459 2922 3460 2926
rect 3454 2921 3460 2922
rect 3592 2909 3594 2937
rect 3590 2908 3596 2909
rect 3590 2904 3591 2908
rect 3595 2904 3596 2908
rect 3590 2903 3596 2904
rect 2138 2899 2144 2900
rect 2138 2895 2139 2899
rect 2143 2895 2144 2899
rect 2138 2894 2144 2895
rect 2346 2899 2352 2900
rect 2346 2895 2347 2899
rect 2351 2895 2352 2899
rect 2346 2894 2352 2895
rect 2494 2899 2500 2900
rect 2494 2895 2495 2899
rect 2499 2895 2500 2899
rect 2494 2894 2500 2895
rect 2722 2899 2728 2900
rect 2722 2895 2723 2899
rect 2727 2895 2728 2899
rect 2722 2894 2728 2895
rect 2878 2899 2884 2900
rect 2878 2895 2879 2899
rect 2883 2895 2884 2899
rect 2878 2894 2884 2895
rect 3098 2899 3104 2900
rect 3098 2895 3099 2899
rect 3103 2895 3104 2899
rect 3098 2894 3104 2895
rect 3202 2899 3208 2900
rect 3202 2895 3203 2899
rect 3207 2895 3208 2899
rect 3202 2894 3208 2895
rect 3310 2899 3316 2900
rect 3310 2895 3311 2899
rect 3315 2895 3316 2899
rect 3310 2894 3316 2895
rect 3362 2899 3368 2900
rect 3362 2895 3363 2899
rect 3367 2895 3368 2899
rect 3362 2894 3368 2895
rect 2286 2888 2292 2889
rect 2286 2884 2287 2888
rect 2291 2884 2292 2888
rect 2286 2883 2292 2884
rect 2478 2888 2484 2889
rect 2478 2884 2479 2888
rect 2483 2884 2484 2888
rect 2478 2883 2484 2884
rect 2662 2888 2668 2889
rect 2662 2884 2663 2888
rect 2667 2884 2668 2888
rect 2662 2883 2668 2884
rect 2830 2888 2836 2889
rect 2830 2884 2831 2888
rect 2835 2884 2836 2888
rect 2830 2883 2836 2884
rect 2288 2859 2290 2883
rect 2480 2859 2482 2883
rect 2664 2859 2666 2883
rect 2832 2859 2834 2883
rect 2135 2858 2139 2859
rect 2135 2853 2139 2854
rect 2263 2858 2267 2859
rect 2263 2853 2267 2854
rect 2287 2858 2291 2859
rect 2287 2853 2291 2854
rect 2391 2858 2395 2859
rect 2391 2853 2395 2854
rect 2479 2858 2483 2859
rect 2479 2853 2483 2854
rect 2519 2858 2523 2859
rect 2519 2853 2523 2854
rect 2647 2858 2651 2859
rect 2647 2853 2651 2854
rect 2663 2858 2667 2859
rect 2663 2853 2667 2854
rect 2767 2858 2771 2859
rect 2767 2853 2771 2854
rect 2831 2858 2835 2859
rect 2831 2853 2835 2854
rect 2136 2837 2138 2853
rect 2264 2837 2266 2853
rect 2392 2837 2394 2853
rect 2520 2837 2522 2853
rect 2648 2837 2650 2853
rect 2768 2837 2770 2853
rect 2134 2836 2140 2837
rect 2134 2832 2135 2836
rect 2139 2832 2140 2836
rect 2134 2831 2140 2832
rect 2262 2836 2268 2837
rect 2262 2832 2263 2836
rect 2267 2832 2268 2836
rect 2262 2831 2268 2832
rect 2390 2836 2396 2837
rect 2390 2832 2391 2836
rect 2395 2832 2396 2836
rect 2390 2831 2396 2832
rect 2518 2836 2524 2837
rect 2518 2832 2519 2836
rect 2523 2832 2524 2836
rect 2518 2831 2524 2832
rect 2646 2836 2652 2837
rect 2646 2832 2647 2836
rect 2651 2832 2652 2836
rect 2646 2831 2652 2832
rect 2766 2836 2772 2837
rect 2766 2832 2767 2836
rect 2771 2832 2772 2836
rect 2766 2831 2772 2832
rect 2094 2827 2100 2828
rect 2094 2823 2095 2827
rect 2099 2823 2100 2827
rect 1562 2822 1568 2823
rect 1639 2822 1643 2823
rect 1698 2822 1704 2823
rect 1735 2822 1739 2823
rect 1639 2817 1643 2818
rect 1735 2817 1739 2818
rect 1751 2822 1755 2823
rect 1758 2822 1764 2823
rect 1831 2822 1835 2823
rect 2094 2822 2100 2823
rect 2202 2827 2208 2828
rect 2202 2823 2203 2827
rect 2207 2823 2208 2827
rect 2202 2822 2208 2823
rect 2714 2827 2720 2828
rect 2714 2823 2715 2827
rect 2719 2823 2720 2827
rect 2714 2822 2720 2823
rect 1751 2817 1755 2818
rect 1831 2817 1835 2818
rect 1554 2815 1560 2816
rect 1554 2811 1555 2815
rect 1559 2811 1560 2815
rect 1554 2810 1560 2811
rect 1586 2815 1592 2816
rect 1586 2811 1587 2815
rect 1591 2811 1592 2815
rect 1586 2810 1592 2811
rect 1334 2806 1340 2807
rect 1334 2802 1335 2806
rect 1339 2802 1340 2806
rect 1334 2801 1340 2802
rect 1534 2806 1540 2807
rect 1534 2802 1535 2806
rect 1539 2802 1540 2806
rect 1534 2801 1540 2802
rect 1588 2780 1590 2810
rect 1736 2807 1738 2817
rect 1734 2806 1740 2807
rect 1734 2802 1735 2806
rect 1739 2802 1740 2806
rect 1734 2801 1740 2802
rect 1832 2789 1834 2817
rect 1870 2816 1876 2817
rect 1870 2812 1871 2816
rect 1875 2812 1876 2816
rect 1870 2811 1876 2812
rect 1830 2788 1836 2789
rect 1830 2784 1831 2788
rect 1835 2784 1836 2788
rect 1830 2783 1836 2784
rect 1586 2779 1592 2780
rect 1586 2775 1587 2779
rect 1591 2775 1592 2779
rect 1872 2775 1874 2811
rect 2142 2798 2148 2799
rect 2142 2794 2143 2798
rect 2147 2794 2148 2798
rect 2142 2793 2148 2794
rect 2144 2775 2146 2793
rect 2204 2788 2206 2822
rect 2663 2804 2667 2805
rect 2663 2799 2667 2800
rect 2270 2798 2276 2799
rect 2270 2794 2271 2798
rect 2275 2794 2276 2798
rect 2270 2793 2276 2794
rect 2398 2798 2404 2799
rect 2398 2794 2399 2798
rect 2403 2794 2404 2798
rect 2398 2793 2404 2794
rect 2526 2798 2532 2799
rect 2526 2794 2527 2798
rect 2531 2794 2532 2798
rect 2526 2793 2532 2794
rect 2654 2798 2660 2799
rect 2654 2794 2655 2798
rect 2659 2794 2660 2798
rect 2654 2793 2660 2794
rect 2202 2787 2208 2788
rect 2202 2783 2203 2787
rect 2207 2783 2208 2787
rect 2202 2782 2208 2783
rect 2272 2775 2274 2793
rect 2400 2775 2402 2793
rect 2528 2775 2530 2793
rect 2558 2787 2564 2788
rect 2558 2783 2559 2787
rect 2563 2783 2564 2787
rect 2558 2782 2564 2783
rect 1586 2774 1592 2775
rect 1871 2774 1875 2775
rect 1830 2771 1836 2772
rect 1326 2768 1332 2769
rect 1326 2764 1327 2768
rect 1331 2764 1332 2768
rect 1326 2763 1332 2764
rect 1526 2768 1532 2769
rect 1526 2764 1527 2768
rect 1531 2764 1532 2768
rect 1526 2763 1532 2764
rect 1726 2768 1732 2769
rect 1726 2764 1727 2768
rect 1731 2764 1732 2768
rect 1830 2767 1831 2771
rect 1835 2767 1836 2771
rect 1871 2769 1875 2770
rect 2143 2774 2147 2775
rect 2143 2769 2147 2770
rect 2231 2774 2235 2775
rect 2231 2769 2235 2770
rect 2271 2774 2275 2775
rect 2271 2769 2275 2770
rect 2311 2774 2315 2775
rect 2311 2769 2315 2770
rect 2391 2774 2395 2775
rect 2391 2769 2395 2770
rect 2399 2774 2403 2775
rect 2399 2769 2403 2770
rect 2471 2774 2475 2775
rect 2471 2769 2475 2770
rect 2527 2774 2531 2775
rect 2527 2769 2531 2770
rect 2551 2774 2555 2775
rect 2551 2769 2555 2770
rect 1830 2766 1836 2767
rect 1726 2763 1732 2764
rect 1328 2743 1330 2763
rect 1528 2743 1530 2763
rect 1702 2751 1708 2752
rect 1702 2747 1703 2751
rect 1707 2747 1708 2751
rect 1702 2746 1708 2747
rect 1327 2742 1331 2743
rect 1327 2737 1331 2738
rect 1359 2742 1363 2743
rect 1359 2737 1363 2738
rect 1519 2742 1523 2743
rect 1519 2737 1523 2738
rect 1527 2742 1531 2743
rect 1527 2737 1531 2738
rect 1687 2742 1691 2743
rect 1687 2737 1691 2738
rect 1360 2721 1362 2737
rect 1520 2721 1522 2737
rect 1688 2721 1690 2737
rect 1358 2720 1364 2721
rect 1358 2716 1359 2720
rect 1363 2716 1364 2720
rect 1358 2715 1364 2716
rect 1518 2720 1524 2721
rect 1518 2716 1519 2720
rect 1523 2716 1524 2720
rect 1518 2715 1524 2716
rect 1686 2720 1692 2721
rect 1686 2716 1687 2720
rect 1691 2716 1692 2720
rect 1686 2715 1692 2716
rect 478 2711 484 2712
rect 478 2707 479 2711
rect 483 2707 484 2711
rect 478 2706 484 2707
rect 962 2711 968 2712
rect 962 2707 963 2711
rect 967 2707 968 2711
rect 962 2706 968 2707
rect 1110 2711 1116 2712
rect 1110 2707 1111 2711
rect 1115 2707 1116 2711
rect 1110 2706 1116 2707
rect 1266 2711 1272 2712
rect 1266 2707 1267 2711
rect 1271 2707 1272 2711
rect 1426 2711 1432 2712
rect 1266 2706 1272 2707
rect 1358 2707 1364 2708
rect 398 2682 404 2683
rect 398 2678 399 2682
rect 403 2678 404 2682
rect 398 2677 404 2678
rect 262 2671 268 2672
rect 262 2667 263 2671
rect 267 2667 268 2671
rect 143 2666 147 2667
rect 202 2666 208 2667
rect 255 2666 259 2667
rect 262 2666 268 2667
rect 354 2671 360 2672
rect 354 2667 355 2671
rect 359 2667 360 2671
rect 400 2667 402 2677
rect 480 2672 482 2706
rect 650 2703 656 2704
rect 650 2699 651 2703
rect 655 2699 656 2703
rect 650 2698 656 2699
rect 558 2682 564 2683
rect 558 2678 559 2682
rect 563 2678 564 2682
rect 558 2677 564 2678
rect 652 2677 654 2698
rect 718 2682 724 2683
rect 718 2678 719 2682
rect 723 2678 724 2682
rect 718 2677 724 2678
rect 886 2682 892 2683
rect 886 2678 887 2682
rect 891 2678 892 2682
rect 886 2677 892 2678
rect 478 2671 484 2672
rect 478 2667 479 2671
rect 483 2667 484 2671
rect 560 2667 562 2677
rect 651 2676 655 2677
rect 651 2671 655 2672
rect 720 2667 722 2677
rect 888 2667 890 2677
rect 964 2672 966 2706
rect 1046 2682 1052 2683
rect 1046 2678 1047 2682
rect 1051 2678 1052 2682
rect 1046 2677 1052 2678
rect 894 2671 900 2672
rect 894 2667 895 2671
rect 899 2667 900 2671
rect 354 2666 360 2667
rect 399 2666 403 2667
rect 478 2666 484 2667
rect 551 2666 555 2667
rect 143 2661 147 2662
rect 255 2661 259 2662
rect 399 2661 403 2662
rect 551 2661 555 2662
rect 559 2666 563 2667
rect 559 2661 563 2662
rect 711 2666 715 2667
rect 711 2661 715 2662
rect 719 2666 723 2667
rect 719 2661 723 2662
rect 879 2666 883 2667
rect 879 2661 883 2662
rect 887 2666 891 2667
rect 894 2666 900 2667
rect 962 2671 968 2672
rect 962 2667 963 2671
rect 967 2667 968 2671
rect 1048 2667 1050 2677
rect 1112 2672 1114 2706
rect 1358 2703 1359 2707
rect 1363 2703 1364 2707
rect 1426 2707 1427 2711
rect 1431 2707 1432 2711
rect 1426 2706 1432 2707
rect 1586 2711 1592 2712
rect 1586 2707 1587 2711
rect 1591 2707 1592 2711
rect 1586 2706 1592 2707
rect 1358 2702 1364 2703
rect 1206 2682 1212 2683
rect 1206 2678 1207 2682
rect 1211 2678 1212 2682
rect 1206 2677 1212 2678
rect 1110 2671 1116 2672
rect 1110 2667 1111 2671
rect 1115 2667 1116 2671
rect 1208 2667 1210 2677
rect 962 2666 968 2667
rect 1047 2666 1051 2667
rect 1110 2666 1116 2667
rect 1207 2666 1211 2667
rect 887 2661 891 2662
rect 134 2659 140 2660
rect 134 2655 135 2659
rect 139 2655 140 2659
rect 134 2654 140 2655
rect 144 2651 146 2661
rect 194 2659 200 2660
rect 194 2655 195 2659
rect 199 2655 200 2659
rect 194 2654 200 2655
rect 142 2650 148 2651
rect 142 2646 143 2650
rect 147 2646 148 2650
rect 142 2645 148 2646
rect 110 2632 116 2633
rect 110 2628 111 2632
rect 115 2628 116 2632
rect 110 2627 116 2628
rect 196 2624 198 2654
rect 256 2651 258 2661
rect 306 2659 312 2660
rect 306 2655 307 2659
rect 311 2655 312 2659
rect 306 2654 312 2655
rect 254 2650 260 2651
rect 254 2646 255 2650
rect 259 2646 260 2650
rect 254 2645 260 2646
rect 308 2624 310 2654
rect 400 2651 402 2661
rect 450 2659 456 2660
rect 450 2655 451 2659
rect 455 2655 456 2659
rect 450 2654 456 2655
rect 398 2650 404 2651
rect 398 2646 399 2650
rect 403 2646 404 2650
rect 398 2645 404 2646
rect 452 2624 454 2654
rect 552 2651 554 2661
rect 602 2659 608 2660
rect 602 2655 603 2659
rect 607 2655 608 2659
rect 602 2654 608 2655
rect 550 2650 556 2651
rect 550 2646 551 2650
rect 555 2646 556 2650
rect 550 2645 556 2646
rect 604 2624 606 2654
rect 712 2651 714 2661
rect 880 2651 882 2661
rect 710 2650 716 2651
rect 710 2646 711 2650
rect 715 2646 716 2650
rect 710 2645 716 2646
rect 878 2650 884 2651
rect 878 2646 879 2650
rect 883 2646 884 2650
rect 878 2645 884 2646
rect 896 2624 898 2666
rect 1047 2661 1051 2662
rect 1207 2661 1211 2662
rect 1215 2666 1219 2667
rect 1215 2661 1219 2662
rect 938 2659 944 2660
rect 938 2655 939 2659
rect 943 2655 944 2659
rect 938 2654 944 2655
rect 940 2624 942 2654
rect 1048 2651 1050 2661
rect 1134 2659 1140 2660
rect 1134 2655 1135 2659
rect 1139 2655 1140 2659
rect 1134 2654 1140 2655
rect 1186 2659 1192 2660
rect 1186 2655 1187 2659
rect 1191 2655 1192 2659
rect 1186 2654 1192 2655
rect 1046 2650 1052 2651
rect 1046 2646 1047 2650
rect 1051 2646 1052 2650
rect 1046 2645 1052 2646
rect 1136 2624 1138 2654
rect 194 2623 200 2624
rect 194 2619 195 2623
rect 199 2619 200 2623
rect 194 2618 200 2619
rect 306 2623 312 2624
rect 306 2619 307 2623
rect 311 2619 312 2623
rect 306 2618 312 2619
rect 450 2623 456 2624
rect 450 2619 451 2623
rect 455 2619 456 2623
rect 450 2618 456 2619
rect 602 2623 608 2624
rect 602 2619 603 2623
rect 607 2619 608 2623
rect 602 2618 608 2619
rect 894 2623 900 2624
rect 894 2619 895 2623
rect 899 2619 900 2623
rect 894 2618 900 2619
rect 938 2623 944 2624
rect 938 2619 939 2623
rect 943 2619 944 2623
rect 938 2618 944 2619
rect 1134 2623 1140 2624
rect 1134 2619 1135 2623
rect 1139 2619 1140 2623
rect 1134 2618 1140 2619
rect 110 2615 116 2616
rect 110 2611 111 2615
rect 115 2611 116 2615
rect 110 2610 116 2611
rect 134 2612 140 2613
rect 112 2587 114 2610
rect 134 2608 135 2612
rect 139 2608 140 2612
rect 134 2607 140 2608
rect 246 2612 252 2613
rect 246 2608 247 2612
rect 251 2608 252 2612
rect 246 2607 252 2608
rect 390 2612 396 2613
rect 390 2608 391 2612
rect 395 2608 396 2612
rect 390 2607 396 2608
rect 542 2612 548 2613
rect 542 2608 543 2612
rect 547 2608 548 2612
rect 542 2607 548 2608
rect 702 2612 708 2613
rect 702 2608 703 2612
rect 707 2608 708 2612
rect 702 2607 708 2608
rect 870 2612 876 2613
rect 870 2608 871 2612
rect 875 2608 876 2612
rect 870 2607 876 2608
rect 1038 2612 1044 2613
rect 1038 2608 1039 2612
rect 1043 2608 1044 2612
rect 1038 2607 1044 2608
rect 136 2587 138 2607
rect 248 2587 250 2607
rect 392 2587 394 2607
rect 544 2587 546 2607
rect 642 2595 648 2596
rect 642 2591 643 2595
rect 647 2591 648 2595
rect 642 2590 648 2591
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 135 2586 139 2587
rect 135 2581 139 2582
rect 159 2586 163 2587
rect 159 2581 163 2582
rect 247 2586 251 2587
rect 247 2581 251 2582
rect 279 2586 283 2587
rect 279 2581 283 2582
rect 391 2586 395 2587
rect 391 2581 395 2582
rect 415 2586 419 2587
rect 415 2581 419 2582
rect 543 2586 547 2587
rect 543 2581 547 2582
rect 559 2586 563 2587
rect 559 2581 563 2582
rect 112 2562 114 2581
rect 160 2565 162 2581
rect 280 2565 282 2581
rect 416 2565 418 2581
rect 560 2565 562 2581
rect 158 2564 164 2565
rect 110 2561 116 2562
rect 110 2557 111 2561
rect 115 2557 116 2561
rect 158 2560 159 2564
rect 163 2560 164 2564
rect 158 2559 164 2560
rect 278 2564 284 2565
rect 278 2560 279 2564
rect 283 2560 284 2564
rect 278 2559 284 2560
rect 414 2564 420 2565
rect 414 2560 415 2564
rect 419 2560 420 2564
rect 414 2559 420 2560
rect 558 2564 564 2565
rect 558 2560 559 2564
rect 563 2560 564 2564
rect 558 2559 564 2560
rect 644 2557 646 2590
rect 704 2587 706 2607
rect 872 2587 874 2607
rect 1040 2587 1042 2607
rect 703 2586 707 2587
rect 703 2581 707 2582
rect 847 2586 851 2587
rect 847 2581 851 2582
rect 871 2586 875 2587
rect 871 2581 875 2582
rect 983 2586 987 2587
rect 983 2581 987 2582
rect 1039 2586 1043 2587
rect 1039 2581 1043 2582
rect 1119 2586 1123 2587
rect 1119 2581 1123 2582
rect 704 2565 706 2581
rect 848 2565 850 2581
rect 984 2565 986 2581
rect 1120 2565 1122 2581
rect 702 2564 708 2565
rect 702 2560 703 2564
rect 707 2560 708 2564
rect 702 2559 708 2560
rect 846 2564 852 2565
rect 846 2560 847 2564
rect 851 2560 852 2564
rect 846 2559 852 2560
rect 982 2564 988 2565
rect 982 2560 983 2564
rect 987 2560 988 2564
rect 982 2559 988 2560
rect 1118 2564 1124 2565
rect 1118 2560 1119 2564
rect 1123 2560 1124 2564
rect 1118 2559 1124 2560
rect 110 2556 116 2557
rect 175 2556 179 2557
rect 643 2556 647 2557
rect 1188 2556 1190 2654
rect 1216 2651 1218 2661
rect 1360 2660 1362 2702
rect 1366 2682 1372 2683
rect 1366 2678 1367 2682
rect 1371 2678 1372 2682
rect 1366 2677 1372 2678
rect 1368 2667 1370 2677
rect 1428 2672 1430 2706
rect 1526 2682 1532 2683
rect 1526 2678 1527 2682
rect 1531 2678 1532 2682
rect 1526 2677 1532 2678
rect 1426 2671 1432 2672
rect 1426 2667 1427 2671
rect 1431 2667 1432 2671
rect 1528 2667 1530 2677
rect 1588 2672 1590 2706
rect 1694 2682 1700 2683
rect 1694 2678 1695 2682
rect 1699 2678 1700 2682
rect 1694 2677 1700 2678
rect 1586 2671 1592 2672
rect 1586 2667 1587 2671
rect 1591 2667 1592 2671
rect 1696 2667 1698 2677
rect 1704 2672 1706 2746
rect 1728 2743 1730 2763
rect 1832 2743 1834 2766
rect 1727 2742 1731 2743
rect 1727 2737 1731 2738
rect 1831 2742 1835 2743
rect 1872 2741 1874 2769
rect 2232 2759 2234 2769
rect 2282 2767 2288 2768
rect 2282 2763 2283 2767
rect 2287 2763 2288 2767
rect 2282 2762 2288 2763
rect 2230 2758 2236 2759
rect 2230 2754 2231 2758
rect 2235 2754 2236 2758
rect 2230 2753 2236 2754
rect 1831 2737 1835 2738
rect 1870 2740 1876 2741
rect 1832 2718 1834 2737
rect 1870 2736 1871 2740
rect 1875 2736 1876 2740
rect 1870 2735 1876 2736
rect 2284 2732 2286 2762
rect 2312 2759 2314 2769
rect 2362 2767 2368 2768
rect 2362 2763 2363 2767
rect 2367 2763 2368 2767
rect 2362 2762 2368 2763
rect 2310 2758 2316 2759
rect 2310 2754 2311 2758
rect 2315 2754 2316 2758
rect 2310 2753 2316 2754
rect 2364 2732 2366 2762
rect 2392 2759 2394 2769
rect 2442 2767 2448 2768
rect 2442 2763 2443 2767
rect 2447 2763 2448 2767
rect 2442 2762 2448 2763
rect 2390 2758 2396 2759
rect 2390 2754 2391 2758
rect 2395 2754 2396 2758
rect 2390 2753 2396 2754
rect 2444 2732 2446 2762
rect 2472 2759 2474 2769
rect 2542 2767 2548 2768
rect 2542 2763 2543 2767
rect 2547 2763 2548 2767
rect 2542 2762 2548 2763
rect 2470 2758 2476 2759
rect 2470 2754 2471 2758
rect 2475 2754 2476 2758
rect 2470 2753 2476 2754
rect 2544 2732 2546 2762
rect 2552 2759 2554 2769
rect 2550 2758 2556 2759
rect 2550 2754 2551 2758
rect 2555 2754 2556 2758
rect 2550 2753 2556 2754
rect 2560 2732 2562 2782
rect 2656 2775 2658 2793
rect 2664 2788 2666 2799
rect 2716 2788 2718 2822
rect 2826 2819 2832 2820
rect 2826 2815 2827 2819
rect 2831 2815 2832 2819
rect 2826 2814 2832 2815
rect 2774 2798 2780 2799
rect 2774 2794 2775 2798
rect 2779 2794 2780 2798
rect 2774 2793 2780 2794
rect 2662 2787 2668 2788
rect 2662 2783 2663 2787
rect 2667 2783 2668 2787
rect 2662 2782 2668 2783
rect 2714 2787 2720 2788
rect 2714 2783 2715 2787
rect 2719 2783 2720 2787
rect 2714 2782 2720 2783
rect 2776 2775 2778 2793
rect 2639 2774 2643 2775
rect 2639 2769 2643 2770
rect 2655 2774 2659 2775
rect 2655 2769 2659 2770
rect 2727 2774 2731 2775
rect 2727 2769 2731 2770
rect 2775 2774 2779 2775
rect 2775 2769 2779 2770
rect 2815 2774 2819 2775
rect 2815 2769 2819 2770
rect 2640 2759 2642 2769
rect 2646 2767 2652 2768
rect 2646 2762 2647 2767
rect 2651 2762 2652 2767
rect 2690 2767 2696 2768
rect 2690 2763 2691 2767
rect 2695 2763 2696 2767
rect 2690 2762 2696 2763
rect 2647 2759 2651 2760
rect 2638 2758 2644 2759
rect 2638 2754 2639 2758
rect 2643 2754 2644 2758
rect 2638 2753 2644 2754
rect 2692 2732 2694 2762
rect 2728 2759 2730 2769
rect 2816 2759 2818 2769
rect 2828 2768 2830 2814
rect 2880 2788 2882 2894
rect 3590 2891 3596 2892
rect 2990 2888 2996 2889
rect 2990 2884 2991 2888
rect 2995 2884 2996 2888
rect 2990 2883 2996 2884
rect 3142 2888 3148 2889
rect 3142 2884 3143 2888
rect 3147 2884 3148 2888
rect 3142 2883 3148 2884
rect 3294 2888 3300 2889
rect 3294 2884 3295 2888
rect 3299 2884 3300 2888
rect 3294 2883 3300 2884
rect 3446 2888 3452 2889
rect 3446 2884 3447 2888
rect 3451 2884 3452 2888
rect 3590 2887 3591 2891
rect 3595 2887 3596 2891
rect 3590 2886 3596 2887
rect 3446 2883 3452 2884
rect 2992 2859 2994 2883
rect 3144 2859 3146 2883
rect 3296 2859 3298 2883
rect 3448 2859 3450 2883
rect 3592 2859 3594 2886
rect 2887 2858 2891 2859
rect 2887 2853 2891 2854
rect 2991 2858 2995 2859
rect 2991 2853 2995 2854
rect 3007 2858 3011 2859
rect 3007 2853 3011 2854
rect 3135 2858 3139 2859
rect 3135 2853 3139 2854
rect 3143 2858 3147 2859
rect 3143 2853 3147 2854
rect 3295 2858 3299 2859
rect 3295 2853 3299 2854
rect 3447 2858 3451 2859
rect 3447 2853 3451 2854
rect 3591 2858 3595 2859
rect 3591 2853 3595 2854
rect 2888 2837 2890 2853
rect 3008 2837 3010 2853
rect 3136 2837 3138 2853
rect 2886 2836 2892 2837
rect 2886 2832 2887 2836
rect 2891 2832 2892 2836
rect 2886 2831 2892 2832
rect 3006 2836 3012 2837
rect 3006 2832 3007 2836
rect 3011 2832 3012 2836
rect 3006 2831 3012 2832
rect 3134 2836 3140 2837
rect 3134 2832 3135 2836
rect 3139 2832 3140 2836
rect 3592 2834 3594 2853
rect 3134 2831 3140 2832
rect 3590 2833 3596 2834
rect 3590 2829 3591 2833
rect 3595 2829 3596 2833
rect 3590 2828 3596 2829
rect 2954 2827 2960 2828
rect 2954 2823 2955 2827
rect 2959 2823 2960 2827
rect 2954 2822 2960 2823
rect 3078 2827 3084 2828
rect 3078 2823 3079 2827
rect 3083 2823 3084 2827
rect 3078 2822 3084 2823
rect 3086 2827 3092 2828
rect 3086 2823 3087 2827
rect 3091 2823 3092 2827
rect 3086 2822 3092 2823
rect 2894 2798 2900 2799
rect 2894 2794 2895 2798
rect 2899 2794 2900 2798
rect 2894 2793 2900 2794
rect 2878 2787 2884 2788
rect 2878 2783 2879 2787
rect 2883 2783 2884 2787
rect 2878 2782 2884 2783
rect 2896 2775 2898 2793
rect 2956 2788 2958 2822
rect 3014 2798 3020 2799
rect 3014 2794 3015 2798
rect 3019 2794 3020 2798
rect 3014 2793 3020 2794
rect 2954 2787 2960 2788
rect 2954 2783 2955 2787
rect 2959 2783 2960 2787
rect 2954 2782 2960 2783
rect 3016 2775 3018 2793
rect 3080 2788 3082 2822
rect 3088 2805 3090 2822
rect 3590 2816 3596 2817
rect 3590 2812 3591 2816
rect 3595 2812 3596 2816
rect 3590 2811 3596 2812
rect 3087 2804 3091 2805
rect 3087 2799 3091 2800
rect 3142 2798 3148 2799
rect 3142 2794 3143 2798
rect 3147 2794 3148 2798
rect 3142 2793 3148 2794
rect 3078 2787 3084 2788
rect 3078 2783 3079 2787
rect 3083 2783 3084 2787
rect 3078 2782 3084 2783
rect 3144 2775 3146 2793
rect 3592 2775 3594 2811
rect 2895 2774 2899 2775
rect 2895 2769 2899 2770
rect 2903 2774 2907 2775
rect 2903 2769 2907 2770
rect 2991 2774 2995 2775
rect 2991 2769 2995 2770
rect 3015 2774 3019 2775
rect 3015 2769 3019 2770
rect 3143 2774 3147 2775
rect 3143 2769 3147 2770
rect 3591 2774 3595 2775
rect 3591 2769 3595 2770
rect 2826 2767 2832 2768
rect 2826 2763 2827 2767
rect 2831 2763 2832 2767
rect 2826 2762 2832 2763
rect 2866 2767 2872 2768
rect 2866 2763 2867 2767
rect 2871 2763 2872 2767
rect 2866 2762 2872 2763
rect 2726 2758 2732 2759
rect 2726 2754 2727 2758
rect 2731 2754 2732 2758
rect 2726 2753 2732 2754
rect 2814 2758 2820 2759
rect 2814 2754 2815 2758
rect 2819 2754 2820 2758
rect 2814 2753 2820 2754
rect 2868 2732 2870 2762
rect 2904 2759 2906 2769
rect 2954 2767 2960 2768
rect 2954 2763 2955 2767
rect 2959 2763 2960 2767
rect 2954 2762 2960 2763
rect 2902 2758 2908 2759
rect 2902 2754 2903 2758
rect 2907 2754 2908 2758
rect 2902 2753 2908 2754
rect 2956 2732 2958 2762
rect 2992 2759 2994 2769
rect 2999 2764 3003 2765
rect 2999 2759 3003 2760
rect 2990 2758 2996 2759
rect 2990 2754 2991 2758
rect 2995 2754 2996 2758
rect 2990 2753 2996 2754
rect 3000 2732 3002 2759
rect 3592 2741 3594 2769
rect 3590 2740 3596 2741
rect 3590 2736 3591 2740
rect 3595 2736 3596 2740
rect 3590 2735 3596 2736
rect 2282 2731 2288 2732
rect 2282 2727 2283 2731
rect 2287 2727 2288 2731
rect 2282 2726 2288 2727
rect 2362 2731 2368 2732
rect 2362 2727 2363 2731
rect 2367 2727 2368 2731
rect 2362 2726 2368 2727
rect 2442 2731 2448 2732
rect 2442 2727 2443 2731
rect 2447 2727 2448 2731
rect 2442 2726 2448 2727
rect 2542 2731 2548 2732
rect 2542 2727 2543 2731
rect 2547 2727 2548 2731
rect 2542 2726 2548 2727
rect 2558 2731 2564 2732
rect 2558 2727 2559 2731
rect 2563 2727 2564 2731
rect 2558 2726 2564 2727
rect 2690 2731 2696 2732
rect 2690 2727 2691 2731
rect 2695 2727 2696 2731
rect 2690 2726 2696 2727
rect 2778 2731 2784 2732
rect 2778 2727 2779 2731
rect 2783 2727 2784 2731
rect 2778 2726 2784 2727
rect 2866 2731 2872 2732
rect 2866 2727 2867 2731
rect 2871 2727 2872 2731
rect 2866 2726 2872 2727
rect 2954 2731 2960 2732
rect 2954 2727 2955 2731
rect 2959 2727 2960 2731
rect 2954 2726 2960 2727
rect 2998 2731 3004 2732
rect 2998 2727 2999 2731
rect 3003 2727 3004 2731
rect 2998 2726 3004 2727
rect 1870 2723 1876 2724
rect 1870 2719 1871 2723
rect 1875 2719 1876 2723
rect 1870 2718 1876 2719
rect 2222 2720 2228 2721
rect 1830 2717 1836 2718
rect 1830 2713 1831 2717
rect 1835 2713 1836 2717
rect 1830 2712 1836 2713
rect 1830 2700 1836 2701
rect 1830 2696 1831 2700
rect 1835 2696 1836 2700
rect 1872 2699 1874 2718
rect 2222 2716 2223 2720
rect 2227 2716 2228 2720
rect 2222 2715 2228 2716
rect 2302 2720 2308 2721
rect 2302 2716 2303 2720
rect 2307 2716 2308 2720
rect 2302 2715 2308 2716
rect 2382 2720 2388 2721
rect 2382 2716 2383 2720
rect 2387 2716 2388 2720
rect 2382 2715 2388 2716
rect 2462 2720 2468 2721
rect 2462 2716 2463 2720
rect 2467 2716 2468 2720
rect 2462 2715 2468 2716
rect 2542 2720 2548 2721
rect 2542 2716 2543 2720
rect 2547 2716 2548 2720
rect 2542 2715 2548 2716
rect 2630 2720 2636 2721
rect 2630 2716 2631 2720
rect 2635 2716 2636 2720
rect 2630 2715 2636 2716
rect 2718 2720 2724 2721
rect 2718 2716 2719 2720
rect 2723 2716 2724 2720
rect 2718 2715 2724 2716
rect 2224 2699 2226 2715
rect 2304 2699 2306 2715
rect 2384 2699 2386 2715
rect 2464 2699 2466 2715
rect 2544 2699 2546 2715
rect 2632 2699 2634 2715
rect 2720 2699 2722 2715
rect 1830 2695 1836 2696
rect 1871 2698 1875 2699
rect 1702 2671 1708 2672
rect 1702 2667 1703 2671
rect 1707 2667 1708 2671
rect 1832 2667 1834 2695
rect 1871 2693 1875 2694
rect 2223 2698 2227 2699
rect 2223 2693 2227 2694
rect 2239 2698 2243 2699
rect 2239 2693 2243 2694
rect 2303 2698 2307 2699
rect 2303 2693 2307 2694
rect 2319 2698 2323 2699
rect 2319 2693 2323 2694
rect 2383 2698 2387 2699
rect 2383 2693 2387 2694
rect 2399 2698 2403 2699
rect 2399 2693 2403 2694
rect 2463 2698 2467 2699
rect 2463 2693 2467 2694
rect 2479 2698 2483 2699
rect 2479 2693 2483 2694
rect 2543 2698 2547 2699
rect 2543 2693 2547 2694
rect 2559 2698 2563 2699
rect 2559 2693 2563 2694
rect 2631 2698 2635 2699
rect 2631 2693 2635 2694
rect 2639 2698 2643 2699
rect 2639 2693 2643 2694
rect 2719 2698 2723 2699
rect 2719 2693 2723 2694
rect 1872 2674 1874 2693
rect 2240 2677 2242 2693
rect 2320 2677 2322 2693
rect 2400 2677 2402 2693
rect 2480 2677 2482 2693
rect 2560 2677 2562 2693
rect 2640 2677 2642 2693
rect 2720 2677 2722 2693
rect 2238 2676 2244 2677
rect 1870 2673 1876 2674
rect 1870 2669 1871 2673
rect 1875 2669 1876 2673
rect 2238 2672 2239 2676
rect 2243 2672 2244 2676
rect 2238 2671 2244 2672
rect 2318 2676 2324 2677
rect 2318 2672 2319 2676
rect 2323 2672 2324 2676
rect 2318 2671 2324 2672
rect 2398 2676 2404 2677
rect 2398 2672 2399 2676
rect 2403 2672 2404 2676
rect 2398 2671 2404 2672
rect 2478 2676 2484 2677
rect 2478 2672 2479 2676
rect 2483 2672 2484 2676
rect 2478 2671 2484 2672
rect 2558 2676 2564 2677
rect 2558 2672 2559 2676
rect 2563 2672 2564 2676
rect 2558 2671 2564 2672
rect 2638 2676 2644 2677
rect 2638 2672 2639 2676
rect 2643 2672 2644 2676
rect 2638 2671 2644 2672
rect 2718 2676 2724 2677
rect 2718 2672 2719 2676
rect 2723 2672 2724 2676
rect 2718 2671 2724 2672
rect 1870 2668 1876 2669
rect 2386 2667 2392 2668
rect 1367 2666 1371 2667
rect 1367 2661 1371 2662
rect 1391 2666 1395 2667
rect 1426 2666 1432 2667
rect 1527 2666 1531 2667
rect 1391 2661 1395 2662
rect 1527 2661 1531 2662
rect 1567 2666 1571 2667
rect 1586 2666 1592 2667
rect 1695 2666 1699 2667
rect 1702 2666 1708 2667
rect 1831 2666 1835 2667
rect 1567 2661 1571 2662
rect 1695 2661 1699 2662
rect 2386 2663 2387 2667
rect 2391 2663 2392 2667
rect 2386 2662 2392 2663
rect 2466 2667 2472 2668
rect 2466 2663 2467 2667
rect 2471 2663 2472 2667
rect 2466 2662 2472 2663
rect 2546 2667 2552 2668
rect 2546 2663 2547 2667
rect 2551 2663 2552 2667
rect 2706 2667 2712 2668
rect 2546 2662 2552 2663
rect 2638 2663 2644 2664
rect 1831 2661 1835 2662
rect 1358 2659 1364 2660
rect 1358 2655 1359 2659
rect 1363 2655 1364 2659
rect 1358 2654 1364 2655
rect 1392 2651 1394 2661
rect 1442 2659 1448 2660
rect 1442 2655 1443 2659
rect 1447 2655 1448 2659
rect 1442 2654 1448 2655
rect 1214 2650 1220 2651
rect 1214 2646 1215 2650
rect 1219 2646 1220 2650
rect 1214 2645 1220 2646
rect 1390 2650 1396 2651
rect 1390 2646 1391 2650
rect 1395 2646 1396 2650
rect 1390 2645 1396 2646
rect 1444 2624 1446 2654
rect 1568 2651 1570 2661
rect 1566 2650 1572 2651
rect 1566 2646 1567 2650
rect 1571 2646 1572 2650
rect 1566 2645 1572 2646
rect 1832 2633 1834 2661
rect 1870 2656 1876 2657
rect 1870 2652 1871 2656
rect 1875 2652 1876 2656
rect 1870 2651 1876 2652
rect 1830 2632 1836 2633
rect 1830 2628 1831 2632
rect 1835 2628 1836 2632
rect 1830 2627 1836 2628
rect 1442 2623 1448 2624
rect 1442 2619 1443 2623
rect 1447 2619 1448 2623
rect 1442 2618 1448 2619
rect 1830 2615 1836 2616
rect 1872 2615 1874 2651
rect 2246 2638 2252 2639
rect 2246 2634 2247 2638
rect 2251 2634 2252 2638
rect 2246 2633 2252 2634
rect 2326 2638 2332 2639
rect 2326 2634 2327 2638
rect 2331 2634 2332 2638
rect 2326 2633 2332 2634
rect 2248 2615 2250 2633
rect 2328 2615 2330 2633
rect 2388 2628 2390 2662
rect 2406 2638 2412 2639
rect 2406 2634 2407 2638
rect 2411 2634 2412 2638
rect 2406 2633 2412 2634
rect 2386 2627 2392 2628
rect 2386 2623 2387 2627
rect 2391 2623 2392 2627
rect 2386 2622 2392 2623
rect 2408 2615 2410 2633
rect 2468 2628 2470 2662
rect 2486 2638 2492 2639
rect 2486 2634 2487 2638
rect 2491 2634 2492 2638
rect 2486 2633 2492 2634
rect 2466 2627 2472 2628
rect 2466 2623 2467 2627
rect 2471 2623 2472 2627
rect 2466 2622 2472 2623
rect 2474 2615 2480 2616
rect 2488 2615 2490 2633
rect 2548 2628 2550 2662
rect 2638 2659 2639 2663
rect 2643 2659 2644 2663
rect 2706 2663 2707 2667
rect 2711 2663 2712 2667
rect 2706 2662 2712 2663
rect 2638 2658 2644 2659
rect 2566 2638 2572 2639
rect 2566 2634 2567 2638
rect 2571 2634 2572 2638
rect 2566 2633 2572 2634
rect 2546 2627 2552 2628
rect 2546 2623 2547 2627
rect 2551 2623 2552 2627
rect 2546 2622 2552 2623
rect 2568 2615 2570 2633
rect 2598 2627 2604 2628
rect 2598 2623 2599 2627
rect 2603 2623 2604 2627
rect 2598 2622 2604 2623
rect 1206 2612 1212 2613
rect 1206 2608 1207 2612
rect 1211 2608 1212 2612
rect 1206 2607 1212 2608
rect 1382 2612 1388 2613
rect 1382 2608 1383 2612
rect 1387 2608 1388 2612
rect 1382 2607 1388 2608
rect 1558 2612 1564 2613
rect 1558 2608 1559 2612
rect 1563 2608 1564 2612
rect 1830 2611 1831 2615
rect 1835 2611 1836 2615
rect 1830 2610 1836 2611
rect 1871 2614 1875 2615
rect 1558 2607 1564 2608
rect 1208 2587 1210 2607
rect 1384 2587 1386 2607
rect 1542 2595 1548 2596
rect 1542 2591 1543 2595
rect 1547 2591 1548 2595
rect 1542 2590 1548 2591
rect 1207 2586 1211 2587
rect 1207 2581 1211 2582
rect 1255 2586 1259 2587
rect 1255 2581 1259 2582
rect 1383 2586 1387 2587
rect 1383 2581 1387 2582
rect 1391 2586 1395 2587
rect 1391 2581 1395 2582
rect 1527 2586 1531 2587
rect 1527 2581 1531 2582
rect 1256 2565 1258 2581
rect 1392 2565 1394 2581
rect 1528 2565 1530 2581
rect 1254 2564 1260 2565
rect 1254 2560 1255 2564
rect 1259 2560 1260 2564
rect 1254 2559 1260 2560
rect 1390 2564 1396 2565
rect 1390 2560 1391 2564
rect 1395 2560 1396 2564
rect 1390 2559 1396 2560
rect 1526 2564 1532 2565
rect 1526 2560 1527 2564
rect 1531 2560 1532 2564
rect 1526 2559 1532 2560
rect 175 2551 179 2552
rect 226 2555 232 2556
rect 226 2551 227 2555
rect 231 2551 232 2555
rect 110 2544 116 2545
rect 110 2540 111 2544
rect 115 2540 116 2544
rect 110 2539 116 2540
rect 112 2507 114 2539
rect 166 2526 172 2527
rect 166 2522 167 2526
rect 171 2522 172 2526
rect 166 2521 172 2522
rect 168 2507 170 2521
rect 176 2516 178 2551
rect 226 2550 232 2551
rect 346 2555 352 2556
rect 346 2551 347 2555
rect 351 2551 352 2555
rect 346 2550 352 2551
rect 482 2555 488 2556
rect 482 2551 483 2555
rect 487 2551 488 2555
rect 482 2550 488 2551
rect 634 2555 640 2556
rect 634 2551 635 2555
rect 639 2551 640 2555
rect 643 2551 647 2552
rect 666 2555 672 2556
rect 666 2551 667 2555
rect 671 2551 672 2555
rect 634 2550 640 2551
rect 666 2550 672 2551
rect 914 2555 920 2556
rect 914 2551 915 2555
rect 919 2551 920 2555
rect 914 2550 920 2551
rect 1050 2555 1056 2556
rect 1050 2551 1051 2555
rect 1055 2551 1056 2555
rect 1050 2550 1056 2551
rect 1186 2555 1192 2556
rect 1186 2551 1187 2555
rect 1191 2551 1192 2555
rect 1186 2550 1192 2551
rect 1330 2555 1336 2556
rect 1330 2551 1331 2555
rect 1335 2551 1336 2555
rect 1330 2550 1336 2551
rect 1478 2555 1484 2556
rect 1478 2551 1479 2555
rect 1483 2551 1484 2555
rect 1478 2550 1484 2551
rect 228 2516 230 2550
rect 286 2526 292 2527
rect 286 2522 287 2526
rect 291 2522 292 2526
rect 286 2521 292 2522
rect 174 2515 180 2516
rect 174 2511 175 2515
rect 179 2511 180 2515
rect 174 2510 180 2511
rect 226 2515 232 2516
rect 226 2511 227 2515
rect 231 2511 232 2515
rect 226 2510 232 2511
rect 288 2507 290 2521
rect 348 2516 350 2550
rect 422 2526 428 2527
rect 355 2524 359 2525
rect 422 2522 423 2526
rect 427 2522 428 2526
rect 422 2521 428 2522
rect 355 2519 359 2520
rect 346 2515 352 2516
rect 346 2511 347 2515
rect 351 2511 352 2515
rect 346 2510 352 2511
rect 111 2506 115 2507
rect 111 2501 115 2502
rect 167 2506 171 2507
rect 167 2501 171 2502
rect 287 2506 291 2507
rect 287 2501 291 2502
rect 335 2506 339 2507
rect 335 2501 339 2502
rect 112 2473 114 2501
rect 336 2491 338 2501
rect 356 2500 358 2519
rect 424 2507 426 2521
rect 484 2516 486 2550
rect 566 2526 572 2527
rect 566 2522 567 2526
rect 571 2522 572 2526
rect 566 2521 572 2522
rect 482 2515 488 2516
rect 482 2511 483 2515
rect 487 2511 488 2515
rect 482 2510 488 2511
rect 568 2507 570 2521
rect 636 2516 638 2550
rect 668 2525 670 2550
rect 710 2526 716 2527
rect 667 2524 671 2525
rect 710 2522 711 2526
rect 715 2522 716 2526
rect 710 2521 716 2522
rect 854 2526 860 2527
rect 854 2522 855 2526
rect 859 2522 860 2526
rect 854 2521 860 2522
rect 667 2519 671 2520
rect 634 2515 640 2516
rect 634 2511 635 2515
rect 639 2511 640 2515
rect 634 2510 640 2511
rect 712 2507 714 2521
rect 856 2507 858 2521
rect 916 2516 918 2550
rect 990 2526 996 2527
rect 990 2522 991 2526
rect 995 2522 996 2526
rect 990 2521 996 2522
rect 886 2515 892 2516
rect 886 2511 887 2515
rect 891 2511 892 2515
rect 886 2510 892 2511
rect 914 2515 920 2516
rect 914 2511 915 2515
rect 919 2511 920 2515
rect 914 2510 920 2511
rect 415 2506 419 2507
rect 415 2501 419 2502
rect 423 2506 427 2507
rect 423 2501 427 2502
rect 503 2506 507 2507
rect 503 2501 507 2502
rect 567 2506 571 2507
rect 567 2501 571 2502
rect 599 2506 603 2507
rect 599 2501 603 2502
rect 703 2506 707 2507
rect 703 2501 707 2502
rect 711 2506 715 2507
rect 711 2501 715 2502
rect 815 2506 819 2507
rect 815 2501 819 2502
rect 855 2506 859 2507
rect 855 2501 859 2502
rect 354 2499 360 2500
rect 354 2495 355 2499
rect 359 2495 360 2499
rect 354 2494 360 2495
rect 386 2499 392 2500
rect 386 2495 387 2499
rect 391 2495 392 2499
rect 386 2494 392 2495
rect 334 2490 340 2491
rect 334 2486 335 2490
rect 339 2486 340 2490
rect 334 2485 340 2486
rect 110 2472 116 2473
rect 110 2468 111 2472
rect 115 2468 116 2472
rect 110 2467 116 2468
rect 388 2464 390 2494
rect 416 2491 418 2501
rect 466 2499 472 2500
rect 466 2495 467 2499
rect 471 2495 472 2499
rect 466 2494 472 2495
rect 414 2490 420 2491
rect 414 2486 415 2490
rect 419 2486 420 2490
rect 414 2485 420 2486
rect 468 2464 470 2494
rect 504 2491 506 2501
rect 554 2499 560 2500
rect 554 2495 555 2499
rect 559 2495 560 2499
rect 554 2494 560 2495
rect 502 2490 508 2491
rect 502 2486 503 2490
rect 507 2486 508 2490
rect 502 2485 508 2486
rect 556 2464 558 2494
rect 600 2491 602 2501
rect 650 2499 656 2500
rect 650 2495 651 2499
rect 655 2495 656 2499
rect 650 2494 656 2495
rect 598 2490 604 2491
rect 598 2486 599 2490
rect 603 2486 604 2490
rect 598 2485 604 2486
rect 652 2464 654 2494
rect 704 2491 706 2501
rect 754 2499 760 2500
rect 754 2495 755 2499
rect 759 2495 760 2499
rect 754 2494 760 2495
rect 702 2490 708 2491
rect 702 2486 703 2490
rect 707 2486 708 2490
rect 702 2485 708 2486
rect 756 2464 758 2494
rect 816 2491 818 2501
rect 814 2490 820 2491
rect 814 2486 815 2490
rect 819 2486 820 2490
rect 814 2485 820 2486
rect 888 2464 890 2510
rect 992 2507 994 2521
rect 1052 2516 1054 2550
rect 1314 2547 1320 2548
rect 1314 2543 1315 2547
rect 1319 2543 1320 2547
rect 1314 2542 1320 2543
rect 1126 2526 1132 2527
rect 1126 2522 1127 2526
rect 1131 2522 1132 2526
rect 1126 2521 1132 2522
rect 1262 2526 1268 2527
rect 1262 2522 1263 2526
rect 1267 2522 1268 2526
rect 1262 2521 1268 2522
rect 1050 2515 1056 2516
rect 1050 2511 1051 2515
rect 1055 2511 1056 2515
rect 1050 2510 1056 2511
rect 1128 2507 1130 2521
rect 1264 2507 1266 2521
rect 935 2506 939 2507
rect 935 2501 939 2502
rect 991 2506 995 2507
rect 991 2501 995 2502
rect 1063 2506 1067 2507
rect 1063 2501 1067 2502
rect 1127 2506 1131 2507
rect 1127 2501 1131 2502
rect 1191 2506 1195 2507
rect 1191 2501 1195 2502
rect 1263 2506 1267 2507
rect 1263 2501 1267 2502
rect 936 2491 938 2501
rect 998 2499 1004 2500
rect 998 2495 999 2499
rect 1003 2495 1004 2499
rect 998 2494 1004 2495
rect 934 2490 940 2491
rect 934 2486 935 2490
rect 939 2486 940 2490
rect 934 2485 940 2486
rect 1000 2464 1002 2494
rect 1064 2491 1066 2501
rect 1192 2491 1194 2501
rect 1316 2500 1318 2542
rect 1332 2516 1334 2550
rect 1398 2526 1404 2527
rect 1398 2522 1399 2526
rect 1403 2522 1404 2526
rect 1398 2521 1404 2522
rect 1330 2515 1336 2516
rect 1330 2511 1331 2515
rect 1335 2511 1336 2515
rect 1330 2510 1336 2511
rect 1400 2507 1402 2521
rect 1480 2516 1482 2550
rect 1534 2526 1540 2527
rect 1534 2522 1535 2526
rect 1539 2522 1540 2526
rect 1534 2521 1540 2522
rect 1478 2515 1484 2516
rect 1478 2511 1479 2515
rect 1483 2511 1484 2515
rect 1478 2510 1484 2511
rect 1536 2507 1538 2521
rect 1544 2516 1546 2590
rect 1560 2587 1562 2607
rect 1832 2587 1834 2610
rect 1871 2609 1875 2610
rect 2191 2614 2195 2615
rect 2191 2609 2195 2610
rect 2247 2614 2251 2615
rect 2247 2609 2251 2610
rect 2271 2614 2275 2615
rect 2271 2609 2275 2610
rect 2327 2614 2331 2615
rect 2327 2609 2331 2610
rect 2351 2614 2355 2615
rect 2351 2609 2355 2610
rect 2407 2614 2411 2615
rect 2407 2609 2411 2610
rect 2431 2614 2435 2615
rect 2474 2611 2475 2615
rect 2479 2611 2480 2615
rect 2474 2610 2480 2611
rect 2487 2614 2491 2615
rect 2431 2609 2435 2610
rect 1559 2586 1563 2587
rect 1559 2581 1563 2582
rect 1831 2586 1835 2587
rect 1831 2581 1835 2582
rect 1872 2581 1874 2609
rect 2192 2599 2194 2609
rect 2254 2607 2260 2608
rect 2254 2603 2255 2607
rect 2259 2603 2260 2607
rect 2254 2602 2260 2603
rect 2190 2598 2196 2599
rect 2190 2594 2191 2598
rect 2195 2594 2196 2598
rect 2190 2593 2196 2594
rect 1832 2562 1834 2581
rect 1870 2580 1876 2581
rect 1870 2576 1871 2580
rect 1875 2576 1876 2580
rect 1870 2575 1876 2576
rect 2256 2572 2258 2602
rect 2272 2599 2274 2609
rect 2334 2607 2340 2608
rect 2334 2603 2335 2607
rect 2339 2603 2340 2607
rect 2334 2602 2340 2603
rect 2270 2598 2276 2599
rect 2270 2594 2271 2598
rect 2275 2594 2276 2598
rect 2270 2593 2276 2594
rect 2336 2572 2338 2602
rect 2352 2599 2354 2609
rect 2414 2607 2420 2608
rect 2414 2603 2415 2607
rect 2419 2603 2420 2607
rect 2414 2602 2420 2603
rect 2350 2598 2356 2599
rect 2350 2594 2351 2598
rect 2355 2594 2356 2598
rect 2350 2593 2356 2594
rect 2416 2572 2418 2602
rect 2432 2599 2434 2609
rect 2430 2598 2436 2599
rect 2430 2594 2431 2598
rect 2435 2594 2436 2598
rect 2430 2593 2436 2594
rect 2254 2571 2260 2572
rect 2254 2567 2255 2571
rect 2259 2567 2260 2571
rect 2254 2566 2260 2567
rect 2334 2571 2340 2572
rect 2334 2567 2335 2571
rect 2339 2567 2340 2571
rect 2334 2566 2340 2567
rect 2414 2571 2420 2572
rect 2414 2567 2415 2571
rect 2419 2567 2420 2571
rect 2414 2566 2420 2567
rect 1870 2563 1876 2564
rect 1830 2561 1836 2562
rect 1830 2557 1831 2561
rect 1835 2557 1836 2561
rect 1870 2559 1871 2563
rect 1875 2559 1876 2563
rect 1870 2558 1876 2559
rect 2182 2560 2188 2561
rect 1830 2556 1836 2557
rect 1830 2544 1836 2545
rect 1830 2540 1831 2544
rect 1835 2540 1836 2544
rect 1830 2539 1836 2540
rect 1542 2515 1548 2516
rect 1542 2511 1543 2515
rect 1547 2511 1548 2515
rect 1542 2510 1548 2511
rect 1832 2507 1834 2539
rect 1872 2531 1874 2558
rect 2182 2556 2183 2560
rect 2187 2556 2188 2560
rect 2182 2555 2188 2556
rect 2262 2560 2268 2561
rect 2262 2556 2263 2560
rect 2267 2556 2268 2560
rect 2262 2555 2268 2556
rect 2342 2560 2348 2561
rect 2342 2556 2343 2560
rect 2347 2556 2348 2560
rect 2342 2555 2348 2556
rect 2422 2560 2428 2561
rect 2422 2556 2423 2560
rect 2427 2556 2428 2560
rect 2422 2555 2428 2556
rect 2184 2531 2186 2555
rect 2264 2531 2266 2555
rect 2344 2531 2346 2555
rect 2424 2531 2426 2555
rect 1871 2530 1875 2531
rect 1871 2525 1875 2526
rect 2119 2530 2123 2531
rect 2119 2525 2123 2526
rect 2183 2530 2187 2531
rect 2183 2525 2187 2526
rect 2207 2530 2211 2531
rect 2207 2525 2211 2526
rect 2263 2530 2267 2531
rect 2263 2525 2267 2526
rect 2303 2530 2307 2531
rect 2303 2525 2307 2526
rect 2343 2530 2347 2531
rect 2343 2525 2347 2526
rect 2399 2530 2403 2531
rect 2399 2525 2403 2526
rect 2423 2530 2427 2531
rect 2423 2525 2427 2526
rect 1327 2506 1331 2507
rect 1327 2501 1331 2502
rect 1399 2506 1403 2507
rect 1399 2501 1403 2502
rect 1471 2506 1475 2507
rect 1471 2501 1475 2502
rect 1535 2506 1539 2507
rect 1535 2501 1539 2502
rect 1831 2506 1835 2507
rect 1872 2506 1874 2525
rect 2120 2509 2122 2525
rect 2208 2509 2210 2525
rect 2304 2509 2306 2525
rect 2400 2509 2402 2525
rect 2118 2508 2124 2509
rect 1831 2501 1835 2502
rect 1870 2505 1876 2506
rect 1870 2501 1871 2505
rect 1875 2501 1876 2505
rect 2118 2504 2119 2508
rect 2123 2504 2124 2508
rect 2118 2503 2124 2504
rect 2206 2508 2212 2509
rect 2206 2504 2207 2508
rect 2211 2504 2212 2508
rect 2206 2503 2212 2504
rect 2302 2508 2308 2509
rect 2302 2504 2303 2508
rect 2307 2504 2308 2508
rect 2302 2503 2308 2504
rect 2398 2508 2404 2509
rect 2398 2504 2399 2508
rect 2403 2504 2404 2508
rect 2398 2503 2404 2504
rect 1270 2499 1276 2500
rect 1270 2495 1271 2499
rect 1275 2495 1276 2499
rect 1270 2494 1276 2495
rect 1314 2499 1320 2500
rect 1314 2495 1315 2499
rect 1319 2495 1320 2499
rect 1314 2494 1320 2495
rect 1062 2490 1068 2491
rect 1062 2486 1063 2490
rect 1067 2486 1068 2490
rect 1062 2485 1068 2486
rect 1190 2490 1196 2491
rect 1190 2486 1191 2490
rect 1195 2486 1196 2490
rect 1190 2485 1196 2486
rect 386 2463 392 2464
rect 386 2459 387 2463
rect 391 2459 392 2463
rect 386 2458 392 2459
rect 466 2463 472 2464
rect 466 2459 467 2463
rect 471 2459 472 2463
rect 466 2458 472 2459
rect 554 2463 560 2464
rect 554 2459 555 2463
rect 559 2459 560 2463
rect 554 2458 560 2459
rect 650 2463 656 2464
rect 650 2459 651 2463
rect 655 2459 656 2463
rect 650 2458 656 2459
rect 754 2463 760 2464
rect 754 2459 755 2463
rect 759 2459 760 2463
rect 754 2458 760 2459
rect 886 2463 892 2464
rect 886 2459 887 2463
rect 891 2459 892 2463
rect 886 2458 892 2459
rect 998 2463 1004 2464
rect 998 2459 999 2463
rect 1003 2459 1004 2463
rect 998 2458 1004 2459
rect 110 2455 116 2456
rect 110 2451 111 2455
rect 115 2451 116 2455
rect 110 2450 116 2451
rect 326 2452 332 2453
rect 112 2423 114 2450
rect 326 2448 327 2452
rect 331 2448 332 2452
rect 326 2447 332 2448
rect 406 2452 412 2453
rect 406 2448 407 2452
rect 411 2448 412 2452
rect 406 2447 412 2448
rect 494 2452 500 2453
rect 494 2448 495 2452
rect 499 2448 500 2452
rect 494 2447 500 2448
rect 590 2452 596 2453
rect 590 2448 591 2452
rect 595 2448 596 2452
rect 590 2447 596 2448
rect 694 2452 700 2453
rect 694 2448 695 2452
rect 699 2448 700 2452
rect 694 2447 700 2448
rect 806 2452 812 2453
rect 806 2448 807 2452
rect 811 2448 812 2452
rect 806 2447 812 2448
rect 926 2452 932 2453
rect 926 2448 927 2452
rect 931 2448 932 2452
rect 926 2447 932 2448
rect 1054 2452 1060 2453
rect 1054 2448 1055 2452
rect 1059 2448 1060 2452
rect 1054 2447 1060 2448
rect 1182 2452 1188 2453
rect 1182 2448 1183 2452
rect 1187 2448 1188 2452
rect 1182 2447 1188 2448
rect 328 2423 330 2447
rect 408 2423 410 2447
rect 496 2423 498 2447
rect 592 2423 594 2447
rect 696 2423 698 2447
rect 798 2435 804 2436
rect 798 2431 799 2435
rect 803 2431 804 2435
rect 798 2430 804 2431
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 327 2422 331 2423
rect 327 2417 331 2418
rect 383 2422 387 2423
rect 383 2417 387 2418
rect 407 2422 411 2423
rect 407 2417 411 2418
rect 463 2422 467 2423
rect 463 2417 467 2418
rect 495 2422 499 2423
rect 495 2417 499 2418
rect 543 2422 547 2423
rect 543 2417 547 2418
rect 591 2422 595 2423
rect 591 2417 595 2418
rect 623 2422 627 2423
rect 623 2417 627 2418
rect 695 2422 699 2423
rect 695 2417 699 2418
rect 703 2422 707 2423
rect 703 2417 707 2418
rect 783 2422 787 2423
rect 783 2417 787 2418
rect 112 2398 114 2417
rect 384 2401 386 2417
rect 464 2401 466 2417
rect 544 2401 546 2417
rect 624 2401 626 2417
rect 704 2401 706 2417
rect 784 2401 786 2417
rect 382 2400 388 2401
rect 110 2397 116 2398
rect 110 2393 111 2397
rect 115 2393 116 2397
rect 382 2396 383 2400
rect 387 2396 388 2400
rect 382 2395 388 2396
rect 462 2400 468 2401
rect 462 2396 463 2400
rect 467 2396 468 2400
rect 462 2395 468 2396
rect 542 2400 548 2401
rect 542 2396 543 2400
rect 547 2396 548 2400
rect 542 2395 548 2396
rect 622 2400 628 2401
rect 622 2396 623 2400
rect 627 2396 628 2400
rect 622 2395 628 2396
rect 702 2400 708 2401
rect 702 2396 703 2400
rect 707 2396 708 2400
rect 702 2395 708 2396
rect 782 2400 788 2401
rect 782 2396 783 2400
rect 787 2396 788 2400
rect 782 2395 788 2396
rect 110 2392 116 2393
rect 450 2391 456 2392
rect 450 2387 451 2391
rect 455 2387 456 2391
rect 450 2386 456 2387
rect 530 2391 536 2392
rect 530 2387 531 2391
rect 535 2387 536 2391
rect 530 2386 536 2387
rect 610 2391 616 2392
rect 610 2387 611 2391
rect 615 2387 616 2391
rect 610 2386 616 2387
rect 690 2391 696 2392
rect 690 2387 691 2391
rect 695 2387 696 2391
rect 690 2386 696 2387
rect 770 2391 776 2392
rect 770 2387 771 2391
rect 775 2387 776 2391
rect 770 2386 776 2387
rect 110 2380 116 2381
rect 110 2376 111 2380
rect 115 2376 116 2380
rect 110 2375 116 2376
rect 112 2347 114 2375
rect 390 2362 396 2363
rect 390 2358 391 2362
rect 395 2358 396 2362
rect 390 2357 396 2358
rect 392 2347 394 2357
rect 452 2352 454 2386
rect 470 2362 476 2363
rect 470 2358 471 2362
rect 475 2358 476 2362
rect 470 2357 476 2358
rect 450 2351 456 2352
rect 450 2347 451 2351
rect 455 2347 456 2351
rect 472 2347 474 2357
rect 532 2352 534 2386
rect 550 2362 556 2363
rect 550 2358 551 2362
rect 555 2358 556 2362
rect 550 2357 556 2358
rect 530 2351 536 2352
rect 530 2347 531 2351
rect 535 2347 536 2351
rect 552 2347 554 2357
rect 612 2352 614 2386
rect 630 2362 636 2363
rect 630 2358 631 2362
rect 635 2358 636 2362
rect 630 2357 636 2358
rect 610 2351 616 2352
rect 610 2347 611 2351
rect 615 2347 616 2351
rect 632 2347 634 2357
rect 692 2352 694 2386
rect 710 2362 716 2363
rect 710 2358 711 2362
rect 715 2358 716 2362
rect 710 2357 716 2358
rect 690 2351 696 2352
rect 690 2347 691 2351
rect 695 2347 696 2351
rect 712 2347 714 2357
rect 772 2352 774 2386
rect 790 2362 796 2363
rect 790 2358 791 2362
rect 795 2358 796 2362
rect 790 2357 796 2358
rect 770 2351 776 2352
rect 770 2347 771 2351
rect 775 2347 776 2351
rect 792 2347 794 2357
rect 111 2346 115 2347
rect 111 2341 115 2342
rect 391 2346 395 2347
rect 450 2346 456 2347
rect 471 2346 475 2347
rect 530 2346 536 2347
rect 551 2346 555 2347
rect 610 2346 616 2347
rect 631 2346 635 2347
rect 690 2346 696 2347
rect 711 2346 715 2347
rect 770 2346 776 2347
rect 791 2346 795 2347
rect 391 2341 395 2342
rect 471 2341 475 2342
rect 551 2341 555 2342
rect 631 2341 635 2342
rect 711 2341 715 2342
rect 800 2344 802 2430
rect 808 2423 810 2447
rect 928 2423 930 2447
rect 1056 2423 1058 2447
rect 1184 2423 1186 2447
rect 807 2422 811 2423
rect 807 2417 811 2418
rect 863 2422 867 2423
rect 863 2417 867 2418
rect 927 2422 931 2423
rect 927 2417 931 2418
rect 943 2422 947 2423
rect 943 2417 947 2418
rect 1023 2422 1027 2423
rect 1023 2417 1027 2418
rect 1055 2422 1059 2423
rect 1055 2417 1059 2418
rect 1103 2422 1107 2423
rect 1103 2417 1107 2418
rect 1183 2422 1187 2423
rect 1183 2417 1187 2418
rect 1263 2422 1267 2423
rect 1263 2417 1267 2418
rect 864 2401 866 2417
rect 944 2401 946 2417
rect 1024 2401 1026 2417
rect 1104 2401 1106 2417
rect 1184 2401 1186 2417
rect 1264 2401 1266 2417
rect 862 2400 868 2401
rect 862 2396 863 2400
rect 867 2396 868 2400
rect 862 2395 868 2396
rect 942 2400 948 2401
rect 942 2396 943 2400
rect 947 2396 948 2400
rect 942 2395 948 2396
rect 1022 2400 1028 2401
rect 1022 2396 1023 2400
rect 1027 2396 1028 2400
rect 1022 2395 1028 2396
rect 1102 2400 1108 2401
rect 1102 2396 1103 2400
rect 1107 2396 1108 2400
rect 1102 2395 1108 2396
rect 1182 2400 1188 2401
rect 1182 2396 1183 2400
rect 1187 2396 1188 2400
rect 1182 2395 1188 2396
rect 1262 2400 1268 2401
rect 1262 2396 1263 2400
rect 1267 2396 1268 2400
rect 1262 2395 1268 2396
rect 930 2391 936 2392
rect 862 2387 868 2388
rect 862 2383 863 2387
rect 867 2383 868 2387
rect 930 2387 931 2391
rect 935 2387 936 2391
rect 930 2386 936 2387
rect 1010 2391 1016 2392
rect 1010 2387 1011 2391
rect 1015 2387 1016 2391
rect 1010 2386 1016 2387
rect 1090 2391 1096 2392
rect 1090 2387 1091 2391
rect 1095 2387 1096 2391
rect 1090 2386 1096 2387
rect 1170 2391 1176 2392
rect 1170 2387 1171 2391
rect 1175 2387 1176 2391
rect 1170 2386 1176 2387
rect 1250 2391 1256 2392
rect 1250 2387 1251 2391
rect 1255 2387 1256 2391
rect 1272 2388 1274 2494
rect 1328 2491 1330 2501
rect 1378 2499 1384 2500
rect 1378 2495 1379 2499
rect 1383 2495 1384 2499
rect 1378 2494 1384 2495
rect 1326 2490 1332 2491
rect 1326 2486 1327 2490
rect 1331 2486 1332 2490
rect 1326 2485 1332 2486
rect 1380 2464 1382 2494
rect 1472 2491 1474 2501
rect 1470 2490 1476 2491
rect 1470 2486 1471 2490
rect 1475 2486 1476 2490
rect 1470 2485 1476 2486
rect 1832 2473 1834 2501
rect 1870 2500 1876 2501
rect 2476 2500 2478 2610
rect 2487 2609 2491 2610
rect 2511 2614 2515 2615
rect 2511 2609 2515 2610
rect 2567 2614 2571 2615
rect 2567 2609 2571 2610
rect 2591 2614 2595 2615
rect 2591 2609 2595 2610
rect 2494 2607 2500 2608
rect 2494 2603 2495 2607
rect 2499 2603 2500 2607
rect 2494 2602 2500 2603
rect 2496 2572 2498 2602
rect 2512 2599 2514 2609
rect 2582 2607 2588 2608
rect 2582 2603 2583 2607
rect 2587 2603 2588 2607
rect 2582 2602 2588 2603
rect 2510 2598 2516 2599
rect 2510 2594 2511 2598
rect 2515 2594 2516 2598
rect 2510 2593 2516 2594
rect 2584 2572 2586 2602
rect 2592 2599 2594 2609
rect 2590 2598 2596 2599
rect 2590 2594 2591 2598
rect 2595 2594 2596 2598
rect 2590 2593 2596 2594
rect 2600 2572 2602 2622
rect 2640 2608 2642 2658
rect 2646 2638 2652 2639
rect 2646 2634 2647 2638
rect 2651 2634 2652 2638
rect 2646 2633 2652 2634
rect 2648 2615 2650 2633
rect 2708 2628 2710 2662
rect 2726 2638 2732 2639
rect 2726 2634 2727 2638
rect 2731 2634 2732 2638
rect 2726 2633 2732 2634
rect 2706 2627 2712 2628
rect 2706 2623 2707 2627
rect 2711 2623 2712 2627
rect 2706 2622 2712 2623
rect 2728 2615 2730 2633
rect 2780 2628 2782 2726
rect 3590 2723 3596 2724
rect 2806 2720 2812 2721
rect 2806 2716 2807 2720
rect 2811 2716 2812 2720
rect 2806 2715 2812 2716
rect 2894 2720 2900 2721
rect 2894 2716 2895 2720
rect 2899 2716 2900 2720
rect 2894 2715 2900 2716
rect 2982 2720 2988 2721
rect 2982 2716 2983 2720
rect 2987 2716 2988 2720
rect 3590 2719 3591 2723
rect 3595 2719 3596 2723
rect 3590 2718 3596 2719
rect 2982 2715 2988 2716
rect 2808 2699 2810 2715
rect 2896 2699 2898 2715
rect 2984 2699 2986 2715
rect 3592 2699 3594 2718
rect 2799 2698 2803 2699
rect 2799 2693 2803 2694
rect 2807 2698 2811 2699
rect 2807 2693 2811 2694
rect 2879 2698 2883 2699
rect 2879 2693 2883 2694
rect 2895 2698 2899 2699
rect 2895 2693 2899 2694
rect 2959 2698 2963 2699
rect 2959 2693 2963 2694
rect 2983 2698 2987 2699
rect 2983 2693 2987 2694
rect 3591 2698 3595 2699
rect 3591 2693 3595 2694
rect 2800 2677 2802 2693
rect 2880 2677 2882 2693
rect 2960 2677 2962 2693
rect 2798 2676 2804 2677
rect 2798 2672 2799 2676
rect 2803 2672 2804 2676
rect 2798 2671 2804 2672
rect 2878 2676 2884 2677
rect 2878 2672 2879 2676
rect 2883 2672 2884 2676
rect 2878 2671 2884 2672
rect 2958 2676 2964 2677
rect 2958 2672 2959 2676
rect 2963 2672 2964 2676
rect 3592 2674 3594 2693
rect 2958 2671 2964 2672
rect 3590 2673 3596 2674
rect 3590 2669 3591 2673
rect 3595 2669 3596 2673
rect 3590 2668 3596 2669
rect 2866 2667 2872 2668
rect 2866 2663 2867 2667
rect 2871 2663 2872 2667
rect 2866 2662 2872 2663
rect 2946 2667 2952 2668
rect 2946 2663 2947 2667
rect 2951 2663 2952 2667
rect 2946 2662 2952 2663
rect 2786 2659 2792 2660
rect 2786 2655 2787 2659
rect 2791 2655 2792 2659
rect 2786 2654 2792 2655
rect 2788 2636 2790 2654
rect 2806 2638 2812 2639
rect 2786 2635 2792 2636
rect 2786 2631 2787 2635
rect 2791 2631 2792 2635
rect 2806 2634 2807 2638
rect 2811 2634 2812 2638
rect 2806 2633 2812 2634
rect 2786 2630 2792 2631
rect 2778 2627 2784 2628
rect 2778 2623 2779 2627
rect 2783 2623 2784 2627
rect 2778 2622 2784 2623
rect 2808 2615 2810 2633
rect 2868 2628 2870 2662
rect 2886 2638 2892 2639
rect 2886 2634 2887 2638
rect 2891 2634 2892 2638
rect 2886 2633 2892 2634
rect 2866 2627 2872 2628
rect 2866 2623 2867 2627
rect 2871 2623 2872 2627
rect 2866 2622 2872 2623
rect 2888 2615 2890 2633
rect 2948 2628 2950 2662
rect 3590 2656 3596 2657
rect 3590 2652 3591 2656
rect 3595 2652 3596 2656
rect 3590 2651 3596 2652
rect 2966 2638 2972 2639
rect 2966 2634 2967 2638
rect 2971 2634 2972 2638
rect 2966 2633 2972 2634
rect 2946 2627 2952 2628
rect 2946 2623 2947 2627
rect 2951 2623 2952 2627
rect 2946 2622 2952 2623
rect 2968 2615 2970 2633
rect 3592 2615 3594 2651
rect 2647 2614 2651 2615
rect 2647 2609 2651 2610
rect 2671 2614 2675 2615
rect 2671 2609 2675 2610
rect 2727 2614 2731 2615
rect 2727 2609 2731 2610
rect 2751 2614 2755 2615
rect 2751 2609 2755 2610
rect 2807 2614 2811 2615
rect 2807 2609 2811 2610
rect 2831 2614 2835 2615
rect 2831 2609 2835 2610
rect 2887 2614 2891 2615
rect 2887 2609 2891 2610
rect 2911 2614 2915 2615
rect 2911 2609 2915 2610
rect 2967 2614 2971 2615
rect 2967 2609 2971 2610
rect 2991 2614 2995 2615
rect 2991 2609 2995 2610
rect 3591 2614 3595 2615
rect 3591 2609 3595 2610
rect 2638 2607 2644 2608
rect 2638 2603 2639 2607
rect 2643 2603 2644 2607
rect 2638 2602 2644 2603
rect 2672 2599 2674 2609
rect 2734 2607 2740 2608
rect 2734 2603 2735 2607
rect 2739 2603 2740 2607
rect 2734 2602 2740 2603
rect 2670 2598 2676 2599
rect 2670 2594 2671 2598
rect 2675 2594 2676 2598
rect 2670 2593 2676 2594
rect 2736 2572 2738 2602
rect 2752 2599 2754 2609
rect 2814 2607 2820 2608
rect 2814 2603 2815 2607
rect 2819 2603 2820 2607
rect 2814 2602 2820 2603
rect 2750 2598 2756 2599
rect 2750 2594 2751 2598
rect 2755 2594 2756 2598
rect 2750 2593 2756 2594
rect 2816 2572 2818 2602
rect 2832 2599 2834 2609
rect 2894 2607 2900 2608
rect 2894 2603 2895 2607
rect 2899 2603 2900 2607
rect 2894 2602 2900 2603
rect 2830 2598 2836 2599
rect 2830 2594 2831 2598
rect 2835 2594 2836 2598
rect 2830 2593 2836 2594
rect 2896 2572 2898 2602
rect 2912 2599 2914 2609
rect 2974 2607 2980 2608
rect 2974 2603 2975 2607
rect 2979 2603 2980 2607
rect 2974 2602 2980 2603
rect 2910 2598 2916 2599
rect 2910 2594 2911 2598
rect 2915 2594 2916 2598
rect 2910 2593 2916 2594
rect 2976 2572 2978 2602
rect 2992 2599 2994 2609
rect 2990 2598 2996 2599
rect 2990 2594 2991 2598
rect 2995 2594 2996 2598
rect 2990 2593 2996 2594
rect 3592 2581 3594 2609
rect 3590 2580 3596 2581
rect 3590 2576 3591 2580
rect 3595 2576 3596 2580
rect 3590 2575 3596 2576
rect 2494 2571 2500 2572
rect 2494 2567 2495 2571
rect 2499 2567 2500 2571
rect 2494 2566 2500 2567
rect 2582 2571 2588 2572
rect 2582 2567 2583 2571
rect 2587 2567 2588 2571
rect 2582 2566 2588 2567
rect 2598 2571 2604 2572
rect 2598 2567 2599 2571
rect 2603 2567 2604 2571
rect 2598 2566 2604 2567
rect 2734 2571 2740 2572
rect 2734 2567 2735 2571
rect 2739 2567 2740 2571
rect 2734 2566 2740 2567
rect 2814 2571 2820 2572
rect 2814 2567 2815 2571
rect 2819 2567 2820 2571
rect 2814 2566 2820 2567
rect 2894 2571 2900 2572
rect 2894 2567 2895 2571
rect 2899 2567 2900 2571
rect 2894 2566 2900 2567
rect 2974 2571 2980 2572
rect 2974 2567 2975 2571
rect 2979 2567 2980 2571
rect 2974 2566 2980 2567
rect 3590 2563 3596 2564
rect 2502 2560 2508 2561
rect 2502 2556 2503 2560
rect 2507 2556 2508 2560
rect 2502 2555 2508 2556
rect 2582 2560 2588 2561
rect 2582 2556 2583 2560
rect 2587 2556 2588 2560
rect 2582 2555 2588 2556
rect 2662 2560 2668 2561
rect 2662 2556 2663 2560
rect 2667 2556 2668 2560
rect 2662 2555 2668 2556
rect 2742 2560 2748 2561
rect 2742 2556 2743 2560
rect 2747 2556 2748 2560
rect 2742 2555 2748 2556
rect 2822 2560 2828 2561
rect 2822 2556 2823 2560
rect 2827 2556 2828 2560
rect 2822 2555 2828 2556
rect 2902 2560 2908 2561
rect 2902 2556 2903 2560
rect 2907 2556 2908 2560
rect 2902 2555 2908 2556
rect 2982 2560 2988 2561
rect 2982 2556 2983 2560
rect 2987 2556 2988 2560
rect 3590 2559 3591 2563
rect 3595 2559 3596 2563
rect 3590 2558 3596 2559
rect 2982 2555 2988 2556
rect 2504 2531 2506 2555
rect 2584 2531 2586 2555
rect 2606 2543 2612 2544
rect 2606 2539 2607 2543
rect 2611 2539 2612 2543
rect 2606 2538 2612 2539
rect 2495 2530 2499 2531
rect 2495 2525 2499 2526
rect 2503 2530 2507 2531
rect 2503 2525 2507 2526
rect 2583 2530 2587 2531
rect 2583 2525 2587 2526
rect 2591 2530 2595 2531
rect 2591 2525 2595 2526
rect 2496 2509 2498 2525
rect 2592 2509 2594 2525
rect 2494 2508 2500 2509
rect 2494 2504 2495 2508
rect 2499 2504 2500 2508
rect 2494 2503 2500 2504
rect 2590 2508 2596 2509
rect 2590 2504 2591 2508
rect 2595 2504 2596 2508
rect 2590 2503 2596 2504
rect 2186 2499 2192 2500
rect 2186 2495 2187 2499
rect 2191 2495 2192 2499
rect 2186 2494 2192 2495
rect 2274 2499 2280 2500
rect 2274 2495 2275 2499
rect 2279 2495 2280 2499
rect 2274 2494 2280 2495
rect 2370 2499 2376 2500
rect 2370 2495 2371 2499
rect 2375 2495 2376 2499
rect 2370 2494 2376 2495
rect 2466 2499 2472 2500
rect 2466 2495 2467 2499
rect 2471 2495 2472 2499
rect 2466 2494 2472 2495
rect 2474 2499 2480 2500
rect 2474 2495 2475 2499
rect 2479 2495 2480 2499
rect 2474 2494 2480 2495
rect 1870 2488 1876 2489
rect 1870 2484 1871 2488
rect 1875 2484 1876 2488
rect 1870 2483 1876 2484
rect 1830 2472 1836 2473
rect 1830 2468 1831 2472
rect 1835 2468 1836 2472
rect 1830 2467 1836 2468
rect 1378 2463 1384 2464
rect 1378 2459 1379 2463
rect 1383 2459 1384 2463
rect 1378 2458 1384 2459
rect 1518 2463 1524 2464
rect 1518 2459 1519 2463
rect 1523 2459 1524 2463
rect 1518 2458 1524 2459
rect 1318 2452 1324 2453
rect 1318 2448 1319 2452
rect 1323 2448 1324 2452
rect 1318 2447 1324 2448
rect 1462 2452 1468 2453
rect 1462 2448 1463 2452
rect 1467 2448 1468 2452
rect 1462 2447 1468 2448
rect 1320 2423 1322 2447
rect 1464 2423 1466 2447
rect 1319 2422 1323 2423
rect 1319 2417 1323 2418
rect 1351 2422 1355 2423
rect 1351 2417 1355 2418
rect 1439 2422 1443 2423
rect 1439 2417 1443 2418
rect 1463 2422 1467 2423
rect 1463 2417 1467 2418
rect 1352 2401 1354 2417
rect 1440 2401 1442 2417
rect 1350 2400 1356 2401
rect 1350 2396 1351 2400
rect 1355 2396 1356 2400
rect 1350 2395 1356 2396
rect 1438 2400 1444 2401
rect 1438 2396 1439 2400
rect 1443 2396 1444 2400
rect 1438 2395 1444 2396
rect 1418 2391 1424 2392
rect 1250 2386 1256 2387
rect 1270 2387 1276 2388
rect 862 2382 868 2383
rect 864 2352 866 2382
rect 870 2362 876 2363
rect 870 2358 871 2362
rect 875 2358 876 2362
rect 870 2357 876 2358
rect 862 2351 868 2352
rect 862 2347 863 2351
rect 867 2347 868 2351
rect 872 2347 874 2357
rect 932 2352 934 2386
rect 950 2362 956 2363
rect 950 2358 951 2362
rect 955 2358 956 2362
rect 950 2357 956 2358
rect 930 2351 936 2352
rect 930 2347 931 2351
rect 935 2347 936 2351
rect 952 2347 954 2357
rect 1012 2352 1014 2386
rect 1030 2362 1036 2363
rect 1030 2358 1031 2362
rect 1035 2358 1036 2362
rect 1030 2357 1036 2358
rect 1010 2351 1016 2352
rect 1010 2347 1011 2351
rect 1015 2347 1016 2351
rect 1032 2347 1034 2357
rect 1092 2352 1094 2386
rect 1110 2362 1116 2363
rect 1110 2358 1111 2362
rect 1115 2358 1116 2362
rect 1110 2357 1116 2358
rect 1090 2351 1096 2352
rect 1090 2347 1091 2351
rect 1095 2347 1096 2351
rect 1112 2347 1114 2357
rect 1172 2352 1174 2386
rect 1190 2362 1196 2363
rect 1190 2358 1191 2362
rect 1195 2358 1196 2362
rect 1190 2357 1196 2358
rect 1170 2351 1176 2352
rect 1170 2347 1171 2351
rect 1175 2347 1176 2351
rect 1192 2347 1194 2357
rect 1252 2352 1254 2386
rect 1270 2383 1271 2387
rect 1275 2383 1276 2387
rect 1418 2387 1419 2391
rect 1423 2387 1424 2391
rect 1418 2386 1424 2387
rect 1426 2391 1432 2392
rect 1426 2387 1427 2391
rect 1431 2387 1432 2391
rect 1426 2386 1432 2387
rect 1506 2391 1512 2392
rect 1506 2387 1507 2391
rect 1511 2387 1512 2391
rect 1506 2386 1512 2387
rect 1270 2382 1276 2383
rect 1270 2362 1276 2363
rect 1270 2358 1271 2362
rect 1275 2358 1276 2362
rect 1270 2357 1276 2358
rect 1358 2362 1364 2363
rect 1358 2358 1359 2362
rect 1363 2358 1364 2362
rect 1358 2357 1364 2358
rect 1250 2351 1256 2352
rect 1250 2347 1251 2351
rect 1255 2347 1256 2351
rect 1272 2347 1274 2357
rect 1360 2347 1362 2357
rect 862 2346 868 2347
rect 871 2346 875 2347
rect 930 2346 936 2347
rect 951 2346 955 2347
rect 1010 2346 1016 2347
rect 1031 2346 1035 2347
rect 1090 2346 1096 2347
rect 1111 2346 1115 2347
rect 1170 2346 1176 2347
rect 1191 2346 1195 2347
rect 1250 2346 1256 2347
rect 1271 2346 1275 2347
rect 791 2341 795 2342
rect 798 2343 804 2344
rect 112 2313 114 2341
rect 798 2339 799 2343
rect 803 2339 804 2343
rect 871 2341 875 2342
rect 951 2341 955 2342
rect 1031 2341 1035 2342
rect 1111 2341 1115 2342
rect 1191 2341 1195 2342
rect 1271 2341 1275 2342
rect 1359 2346 1363 2347
rect 1359 2341 1363 2342
rect 1407 2346 1411 2347
rect 1407 2341 1411 2342
rect 798 2338 804 2339
rect 1408 2331 1410 2341
rect 1420 2340 1422 2386
rect 1428 2352 1430 2386
rect 1446 2362 1452 2363
rect 1446 2358 1447 2362
rect 1451 2358 1452 2362
rect 1446 2357 1452 2358
rect 1426 2351 1432 2352
rect 1426 2347 1427 2351
rect 1431 2347 1432 2351
rect 1448 2347 1450 2357
rect 1508 2352 1510 2386
rect 1520 2352 1522 2458
rect 1830 2455 1836 2456
rect 1830 2451 1831 2455
rect 1835 2451 1836 2455
rect 1872 2451 1874 2483
rect 2126 2470 2132 2471
rect 2126 2466 2127 2470
rect 2131 2466 2132 2470
rect 2126 2465 2132 2466
rect 2128 2451 2130 2465
rect 2188 2460 2190 2494
rect 2214 2470 2220 2471
rect 2214 2466 2215 2470
rect 2219 2466 2220 2470
rect 2214 2465 2220 2466
rect 2178 2459 2184 2460
rect 2178 2455 2179 2459
rect 2183 2455 2184 2459
rect 2178 2454 2184 2455
rect 2186 2459 2192 2460
rect 2186 2455 2187 2459
rect 2191 2455 2192 2459
rect 2186 2454 2192 2455
rect 1830 2450 1836 2451
rect 1871 2450 1875 2451
rect 1832 2423 1834 2450
rect 1871 2445 1875 2446
rect 1903 2450 1907 2451
rect 1903 2445 1907 2446
rect 1991 2450 1995 2451
rect 1991 2445 1995 2446
rect 2111 2450 2115 2451
rect 2111 2445 2115 2446
rect 2127 2450 2131 2451
rect 2127 2445 2131 2446
rect 1527 2422 1531 2423
rect 1527 2417 1531 2418
rect 1831 2422 1835 2423
rect 1831 2417 1835 2418
rect 1872 2417 1874 2445
rect 1904 2435 1906 2445
rect 1946 2443 1952 2444
rect 1946 2439 1947 2443
rect 1951 2439 1952 2443
rect 1946 2438 1952 2439
rect 1954 2443 1960 2444
rect 1954 2439 1955 2443
rect 1959 2439 1960 2443
rect 1954 2438 1960 2439
rect 1902 2434 1908 2435
rect 1902 2430 1903 2434
rect 1907 2430 1908 2434
rect 1902 2429 1908 2430
rect 1528 2401 1530 2417
rect 1526 2400 1532 2401
rect 1526 2396 1527 2400
rect 1531 2396 1532 2400
rect 1832 2398 1834 2417
rect 1870 2416 1876 2417
rect 1870 2412 1871 2416
rect 1875 2412 1876 2416
rect 1948 2413 1950 2438
rect 1870 2411 1876 2412
rect 1947 2412 1951 2413
rect 1956 2408 1958 2438
rect 1992 2435 1994 2445
rect 2042 2443 2048 2444
rect 2042 2439 2043 2443
rect 2047 2439 2048 2443
rect 2042 2438 2048 2439
rect 1990 2434 1996 2435
rect 1990 2430 1991 2434
rect 1995 2430 1996 2434
rect 1990 2429 1996 2430
rect 2044 2408 2046 2438
rect 2112 2435 2114 2445
rect 2162 2443 2168 2444
rect 2162 2439 2163 2443
rect 2167 2439 2168 2443
rect 2162 2438 2168 2439
rect 2110 2434 2116 2435
rect 2110 2430 2111 2434
rect 2115 2430 2116 2434
rect 2110 2429 2116 2430
rect 2164 2408 2166 2438
rect 2180 2437 2182 2454
rect 2216 2451 2218 2465
rect 2276 2460 2278 2494
rect 2310 2470 2316 2471
rect 2310 2466 2311 2470
rect 2315 2466 2316 2470
rect 2310 2465 2316 2466
rect 2274 2459 2280 2460
rect 2274 2455 2275 2459
rect 2279 2455 2280 2459
rect 2274 2454 2280 2455
rect 2312 2451 2314 2465
rect 2372 2460 2374 2494
rect 2406 2470 2412 2471
rect 2406 2466 2407 2470
rect 2411 2466 2412 2470
rect 2406 2465 2412 2466
rect 2370 2459 2376 2460
rect 2370 2455 2371 2459
rect 2375 2455 2376 2459
rect 2370 2454 2376 2455
rect 2408 2451 2410 2465
rect 2468 2460 2470 2494
rect 2502 2470 2508 2471
rect 2502 2466 2503 2470
rect 2507 2466 2508 2470
rect 2502 2465 2508 2466
rect 2598 2470 2604 2471
rect 2598 2466 2599 2470
rect 2603 2466 2604 2470
rect 2598 2465 2604 2466
rect 2466 2459 2472 2460
rect 2466 2455 2467 2459
rect 2471 2455 2472 2459
rect 2466 2454 2472 2455
rect 2504 2451 2506 2465
rect 2600 2451 2602 2465
rect 2608 2460 2610 2538
rect 2664 2531 2666 2555
rect 2744 2531 2746 2555
rect 2824 2531 2826 2555
rect 2904 2531 2906 2555
rect 2984 2531 2986 2555
rect 3592 2531 3594 2558
rect 2663 2530 2667 2531
rect 2663 2525 2667 2526
rect 2687 2530 2691 2531
rect 2687 2525 2691 2526
rect 2743 2530 2747 2531
rect 2743 2525 2747 2526
rect 2783 2530 2787 2531
rect 2783 2525 2787 2526
rect 2823 2530 2827 2531
rect 2823 2525 2827 2526
rect 2879 2530 2883 2531
rect 2879 2525 2883 2526
rect 2903 2530 2907 2531
rect 2903 2525 2907 2526
rect 2975 2530 2979 2531
rect 2975 2525 2979 2526
rect 2983 2530 2987 2531
rect 2983 2525 2987 2526
rect 3079 2530 3083 2531
rect 3079 2525 3083 2526
rect 3591 2530 3595 2531
rect 3591 2525 3595 2526
rect 2688 2509 2690 2525
rect 2784 2509 2786 2525
rect 2880 2509 2882 2525
rect 2976 2509 2978 2525
rect 3080 2509 3082 2525
rect 2686 2508 2692 2509
rect 2686 2504 2687 2508
rect 2691 2504 2692 2508
rect 2686 2503 2692 2504
rect 2782 2508 2788 2509
rect 2782 2504 2783 2508
rect 2787 2504 2788 2508
rect 2782 2503 2788 2504
rect 2878 2508 2884 2509
rect 2878 2504 2879 2508
rect 2883 2504 2884 2508
rect 2878 2503 2884 2504
rect 2974 2508 2980 2509
rect 2974 2504 2975 2508
rect 2979 2504 2980 2508
rect 2974 2503 2980 2504
rect 3078 2508 3084 2509
rect 3078 2504 3079 2508
rect 3083 2504 3084 2508
rect 3592 2506 3594 2525
rect 3078 2503 3084 2504
rect 3590 2505 3596 2506
rect 3590 2501 3591 2505
rect 3595 2501 3596 2505
rect 3590 2500 3596 2501
rect 2658 2499 2664 2500
rect 2658 2495 2659 2499
rect 2663 2495 2664 2499
rect 2658 2494 2664 2495
rect 2754 2499 2760 2500
rect 2754 2495 2755 2499
rect 2759 2495 2760 2499
rect 2754 2494 2760 2495
rect 2850 2499 2856 2500
rect 2850 2495 2851 2499
rect 2855 2495 2856 2499
rect 2850 2494 2856 2495
rect 2946 2499 2952 2500
rect 2946 2495 2947 2499
rect 2951 2495 2952 2499
rect 2946 2494 2952 2495
rect 3042 2499 3048 2500
rect 3042 2495 3043 2499
rect 3047 2495 3048 2499
rect 3042 2494 3048 2495
rect 3050 2499 3056 2500
rect 3050 2495 3051 2499
rect 3055 2495 3056 2499
rect 3050 2494 3056 2495
rect 2660 2460 2662 2494
rect 2694 2470 2700 2471
rect 2694 2466 2695 2470
rect 2699 2466 2700 2470
rect 2694 2465 2700 2466
rect 2703 2468 2707 2469
rect 2606 2459 2612 2460
rect 2606 2455 2607 2459
rect 2611 2455 2612 2459
rect 2606 2454 2612 2455
rect 2658 2459 2664 2460
rect 2658 2455 2659 2459
rect 2663 2455 2664 2459
rect 2658 2454 2664 2455
rect 2696 2451 2698 2465
rect 2703 2463 2707 2464
rect 2215 2450 2219 2451
rect 2215 2445 2219 2446
rect 2247 2450 2251 2451
rect 2247 2445 2251 2446
rect 2311 2450 2315 2451
rect 2311 2445 2315 2446
rect 2391 2450 2395 2451
rect 2391 2445 2395 2446
rect 2407 2450 2411 2451
rect 2407 2445 2411 2446
rect 2503 2450 2507 2451
rect 2503 2445 2507 2446
rect 2535 2450 2539 2451
rect 2535 2445 2539 2446
rect 2599 2450 2603 2451
rect 2599 2445 2603 2446
rect 2671 2450 2675 2451
rect 2671 2445 2675 2446
rect 2695 2450 2699 2451
rect 2695 2445 2699 2446
rect 2179 2436 2183 2437
rect 2248 2435 2250 2445
rect 2298 2443 2304 2444
rect 2298 2439 2299 2443
rect 2303 2439 2304 2443
rect 2298 2438 2304 2439
rect 2179 2431 2183 2432
rect 2246 2434 2252 2435
rect 2246 2430 2247 2434
rect 2251 2430 2252 2434
rect 2246 2429 2252 2430
rect 2300 2408 2302 2438
rect 2392 2435 2394 2445
rect 2442 2443 2448 2444
rect 2442 2439 2443 2443
rect 2447 2439 2448 2443
rect 2442 2438 2448 2439
rect 2390 2434 2396 2435
rect 2390 2430 2391 2434
rect 2395 2430 2396 2434
rect 2390 2429 2396 2430
rect 2444 2408 2446 2438
rect 2536 2435 2538 2445
rect 2543 2436 2547 2437
rect 2534 2434 2540 2435
rect 2534 2430 2535 2434
rect 2539 2430 2540 2434
rect 2672 2435 2674 2445
rect 2704 2444 2706 2463
rect 2756 2460 2758 2494
rect 2790 2470 2796 2471
rect 2790 2466 2791 2470
rect 2795 2466 2796 2470
rect 2790 2465 2796 2466
rect 2754 2459 2760 2460
rect 2754 2455 2755 2459
rect 2759 2455 2760 2459
rect 2754 2454 2760 2455
rect 2792 2451 2794 2465
rect 2852 2460 2854 2494
rect 2886 2470 2892 2471
rect 2886 2466 2887 2470
rect 2891 2466 2892 2470
rect 2886 2465 2892 2466
rect 2850 2459 2856 2460
rect 2850 2455 2851 2459
rect 2855 2455 2856 2459
rect 2850 2454 2856 2455
rect 2888 2451 2890 2465
rect 2948 2460 2950 2494
rect 2982 2470 2988 2471
rect 2982 2466 2983 2470
rect 2987 2466 2988 2470
rect 2982 2465 2988 2466
rect 2946 2459 2952 2460
rect 2946 2455 2947 2459
rect 2951 2455 2952 2459
rect 2946 2454 2952 2455
rect 2984 2451 2986 2465
rect 3044 2460 3046 2494
rect 3052 2469 3054 2494
rect 3590 2488 3596 2489
rect 3590 2484 3591 2488
rect 3595 2484 3596 2488
rect 3590 2483 3596 2484
rect 3086 2470 3092 2471
rect 3051 2468 3055 2469
rect 3086 2466 3087 2470
rect 3091 2466 3092 2470
rect 3086 2465 3092 2466
rect 3051 2463 3055 2464
rect 3042 2459 3048 2460
rect 3042 2455 3043 2459
rect 3047 2455 3048 2459
rect 3042 2454 3048 2455
rect 3088 2451 3090 2465
rect 3592 2451 3594 2483
rect 2791 2450 2795 2451
rect 2791 2445 2795 2446
rect 2807 2450 2811 2451
rect 2807 2445 2811 2446
rect 2887 2450 2891 2451
rect 2887 2445 2891 2446
rect 2943 2450 2947 2451
rect 2943 2445 2947 2446
rect 2983 2450 2987 2451
rect 2983 2445 2987 2446
rect 3079 2450 3083 2451
rect 3079 2445 3083 2446
rect 3087 2450 3091 2451
rect 3087 2445 3091 2446
rect 3215 2450 3219 2451
rect 3215 2445 3219 2446
rect 3591 2450 3595 2451
rect 3591 2445 3595 2446
rect 2702 2443 2708 2444
rect 2702 2439 2703 2443
rect 2707 2439 2708 2443
rect 2702 2438 2708 2439
rect 2722 2443 2728 2444
rect 2722 2439 2723 2443
rect 2727 2439 2728 2443
rect 2722 2438 2728 2439
rect 2543 2431 2547 2432
rect 2670 2434 2676 2435
rect 2534 2429 2540 2430
rect 2459 2412 2463 2413
rect 2544 2408 2546 2431
rect 2670 2430 2671 2434
rect 2675 2430 2676 2434
rect 2670 2429 2676 2430
rect 2724 2408 2726 2438
rect 2808 2435 2810 2445
rect 2858 2443 2864 2444
rect 2858 2439 2859 2443
rect 2863 2439 2864 2443
rect 2858 2438 2864 2439
rect 2806 2434 2812 2435
rect 2806 2430 2807 2434
rect 2811 2430 2812 2434
rect 2806 2429 2812 2430
rect 2860 2408 2862 2438
rect 2944 2435 2946 2445
rect 2994 2443 3000 2444
rect 2994 2439 2995 2443
rect 2999 2439 3000 2443
rect 2994 2438 3000 2439
rect 2942 2434 2948 2435
rect 2942 2430 2943 2434
rect 2947 2430 2948 2434
rect 2942 2429 2948 2430
rect 2996 2408 2998 2438
rect 3080 2435 3082 2445
rect 3130 2443 3136 2444
rect 3130 2439 3131 2443
rect 3135 2439 3136 2443
rect 3130 2438 3136 2439
rect 3078 2434 3084 2435
rect 3078 2430 3079 2434
rect 3083 2430 3084 2434
rect 3078 2429 3084 2430
rect 3132 2408 3134 2438
rect 3216 2435 3218 2445
rect 3214 2434 3220 2435
rect 3214 2430 3215 2434
rect 3219 2430 3220 2434
rect 3214 2429 3220 2430
rect 3592 2417 3594 2445
rect 3590 2416 3596 2417
rect 3590 2412 3591 2416
rect 3595 2412 3596 2416
rect 3590 2411 3596 2412
rect 1947 2407 1951 2408
rect 1954 2407 1960 2408
rect 1954 2403 1955 2407
rect 1959 2403 1960 2407
rect 1954 2402 1960 2403
rect 2042 2407 2048 2408
rect 2042 2403 2043 2407
rect 2047 2403 2048 2407
rect 2042 2402 2048 2403
rect 2162 2407 2168 2408
rect 2162 2403 2163 2407
rect 2167 2403 2168 2407
rect 2162 2402 2168 2403
rect 2298 2407 2304 2408
rect 2298 2403 2299 2407
rect 2303 2403 2304 2407
rect 2298 2402 2304 2403
rect 2442 2407 2448 2408
rect 2459 2407 2463 2408
rect 2542 2407 2548 2408
rect 2442 2403 2443 2407
rect 2447 2403 2448 2407
rect 2442 2402 2448 2403
rect 1870 2399 1876 2400
rect 1526 2395 1532 2396
rect 1830 2397 1836 2398
rect 1830 2393 1831 2397
rect 1835 2393 1836 2397
rect 1870 2395 1871 2399
rect 1875 2395 1876 2399
rect 1870 2394 1876 2395
rect 1894 2396 1900 2397
rect 1830 2392 1836 2393
rect 1830 2380 1836 2381
rect 1830 2376 1831 2380
rect 1835 2376 1836 2380
rect 1830 2375 1836 2376
rect 1534 2362 1540 2363
rect 1534 2358 1535 2362
rect 1539 2358 1540 2362
rect 1534 2357 1540 2358
rect 1506 2351 1512 2352
rect 1506 2347 1507 2351
rect 1511 2347 1512 2351
rect 1426 2346 1432 2347
rect 1447 2346 1451 2347
rect 1447 2341 1451 2342
rect 1487 2346 1491 2347
rect 1506 2346 1512 2347
rect 1518 2351 1524 2352
rect 1518 2347 1519 2351
rect 1523 2347 1524 2351
rect 1536 2347 1538 2357
rect 1832 2347 1834 2375
rect 1872 2367 1874 2394
rect 1894 2392 1895 2396
rect 1899 2392 1900 2396
rect 1894 2391 1900 2392
rect 1982 2396 1988 2397
rect 1982 2392 1983 2396
rect 1987 2392 1988 2396
rect 1982 2391 1988 2392
rect 2102 2396 2108 2397
rect 2102 2392 2103 2396
rect 2107 2392 2108 2396
rect 2102 2391 2108 2392
rect 2238 2396 2244 2397
rect 2238 2392 2239 2396
rect 2243 2392 2244 2396
rect 2238 2391 2244 2392
rect 2382 2396 2388 2397
rect 2382 2392 2383 2396
rect 2387 2392 2388 2396
rect 2382 2391 2388 2392
rect 1896 2367 1898 2391
rect 1984 2367 1986 2391
rect 2104 2367 2106 2391
rect 2240 2367 2242 2391
rect 2384 2367 2386 2391
rect 1871 2366 1875 2367
rect 1871 2361 1875 2362
rect 1895 2366 1899 2367
rect 1895 2361 1899 2362
rect 1983 2366 1987 2367
rect 1983 2361 1987 2362
rect 2015 2366 2019 2367
rect 2015 2361 2019 2362
rect 2103 2366 2107 2367
rect 2103 2361 2107 2362
rect 2175 2366 2179 2367
rect 2175 2361 2179 2362
rect 2239 2366 2243 2367
rect 2239 2361 2243 2362
rect 2343 2366 2347 2367
rect 2343 2361 2347 2362
rect 2383 2366 2387 2367
rect 2383 2361 2387 2362
rect 1518 2346 1524 2347
rect 1535 2346 1539 2347
rect 1487 2341 1491 2342
rect 1535 2341 1539 2342
rect 1567 2346 1571 2347
rect 1567 2341 1571 2342
rect 1647 2346 1651 2347
rect 1647 2341 1651 2342
rect 1831 2346 1835 2347
rect 1872 2342 1874 2361
rect 1896 2345 1898 2361
rect 2016 2345 2018 2361
rect 2176 2345 2178 2361
rect 2344 2345 2346 2361
rect 1894 2344 1900 2345
rect 1831 2341 1835 2342
rect 1870 2341 1876 2342
rect 1418 2339 1424 2340
rect 1418 2335 1419 2339
rect 1423 2335 1424 2339
rect 1418 2334 1424 2335
rect 1458 2339 1464 2340
rect 1458 2335 1459 2339
rect 1463 2335 1464 2339
rect 1458 2334 1464 2335
rect 1406 2330 1412 2331
rect 1406 2326 1407 2330
rect 1411 2326 1412 2330
rect 1406 2325 1412 2326
rect 110 2312 116 2313
rect 110 2308 111 2312
rect 115 2308 116 2312
rect 110 2307 116 2308
rect 1460 2304 1462 2334
rect 1488 2331 1490 2341
rect 1558 2339 1564 2340
rect 1558 2335 1559 2339
rect 1563 2335 1564 2339
rect 1558 2334 1564 2335
rect 1486 2330 1492 2331
rect 1486 2326 1487 2330
rect 1491 2326 1492 2330
rect 1486 2325 1492 2326
rect 1560 2304 1562 2334
rect 1568 2331 1570 2341
rect 1618 2339 1624 2340
rect 1618 2335 1619 2339
rect 1623 2335 1624 2339
rect 1618 2334 1624 2335
rect 1566 2330 1572 2331
rect 1566 2326 1567 2330
rect 1571 2326 1572 2330
rect 1566 2325 1572 2326
rect 1620 2304 1622 2334
rect 1648 2331 1650 2341
rect 1646 2330 1652 2331
rect 1646 2326 1647 2330
rect 1651 2326 1652 2330
rect 1646 2325 1652 2326
rect 1832 2313 1834 2341
rect 1870 2337 1871 2341
rect 1875 2337 1876 2341
rect 1894 2340 1895 2344
rect 1899 2340 1900 2344
rect 1894 2339 1900 2340
rect 2014 2344 2020 2345
rect 2014 2340 2015 2344
rect 2019 2340 2020 2344
rect 2014 2339 2020 2340
rect 2174 2344 2180 2345
rect 2174 2340 2175 2344
rect 2179 2340 2180 2344
rect 2174 2339 2180 2340
rect 2342 2344 2348 2345
rect 2342 2340 2343 2344
rect 2347 2340 2348 2344
rect 2342 2339 2348 2340
rect 1870 2336 1876 2337
rect 2460 2336 2462 2407
rect 2542 2403 2543 2407
rect 2547 2403 2548 2407
rect 2542 2402 2548 2403
rect 2722 2407 2728 2408
rect 2722 2403 2723 2407
rect 2727 2403 2728 2407
rect 2722 2402 2728 2403
rect 2858 2407 2864 2408
rect 2858 2403 2859 2407
rect 2863 2403 2864 2407
rect 2858 2402 2864 2403
rect 2994 2407 3000 2408
rect 2994 2403 2995 2407
rect 2999 2403 3000 2407
rect 2994 2402 3000 2403
rect 3130 2407 3136 2408
rect 3130 2403 3131 2407
rect 3135 2403 3136 2407
rect 3130 2402 3136 2403
rect 3590 2399 3596 2400
rect 2526 2396 2532 2397
rect 2526 2392 2527 2396
rect 2531 2392 2532 2396
rect 2526 2391 2532 2392
rect 2662 2396 2668 2397
rect 2662 2392 2663 2396
rect 2667 2392 2668 2396
rect 2662 2391 2668 2392
rect 2798 2396 2804 2397
rect 2798 2392 2799 2396
rect 2803 2392 2804 2396
rect 2798 2391 2804 2392
rect 2934 2396 2940 2397
rect 2934 2392 2935 2396
rect 2939 2392 2940 2396
rect 2934 2391 2940 2392
rect 3070 2396 3076 2397
rect 3070 2392 3071 2396
rect 3075 2392 3076 2396
rect 3070 2391 3076 2392
rect 3206 2396 3212 2397
rect 3206 2392 3207 2396
rect 3211 2392 3212 2396
rect 3590 2395 3591 2399
rect 3595 2395 3596 2399
rect 3590 2394 3596 2395
rect 3206 2391 3212 2392
rect 2528 2367 2530 2391
rect 2664 2367 2666 2391
rect 2800 2367 2802 2391
rect 2936 2367 2938 2391
rect 3072 2367 3074 2391
rect 3138 2379 3144 2380
rect 3138 2375 3139 2379
rect 3143 2375 3144 2379
rect 3138 2374 3144 2375
rect 2511 2366 2515 2367
rect 2511 2361 2515 2362
rect 2527 2366 2531 2367
rect 2527 2361 2531 2362
rect 2663 2366 2667 2367
rect 2663 2361 2667 2362
rect 2671 2366 2675 2367
rect 2671 2361 2675 2362
rect 2799 2366 2803 2367
rect 2799 2361 2803 2362
rect 2823 2366 2827 2367
rect 2823 2361 2827 2362
rect 2935 2366 2939 2367
rect 2935 2361 2939 2362
rect 2959 2366 2963 2367
rect 2959 2361 2963 2362
rect 3071 2366 3075 2367
rect 3071 2361 3075 2362
rect 3079 2366 3083 2367
rect 3079 2361 3083 2362
rect 2512 2345 2514 2361
rect 2672 2345 2674 2361
rect 2824 2345 2826 2361
rect 2960 2345 2962 2361
rect 3080 2345 3082 2361
rect 2510 2344 2516 2345
rect 2510 2340 2511 2344
rect 2515 2340 2516 2344
rect 2510 2339 2516 2340
rect 2670 2344 2676 2345
rect 2670 2340 2671 2344
rect 2675 2340 2676 2344
rect 2670 2339 2676 2340
rect 2822 2344 2828 2345
rect 2822 2340 2823 2344
rect 2827 2340 2828 2344
rect 2822 2339 2828 2340
rect 2958 2344 2964 2345
rect 2958 2340 2959 2344
rect 2963 2340 2964 2344
rect 2958 2339 2964 2340
rect 3078 2344 3084 2345
rect 3078 2340 3079 2344
rect 3083 2340 3084 2344
rect 3078 2339 3084 2340
rect 1962 2335 1968 2336
rect 1962 2331 1963 2335
rect 1967 2331 1968 2335
rect 1962 2330 1968 2331
rect 2098 2335 2104 2336
rect 2098 2331 2099 2335
rect 2103 2331 2104 2335
rect 2098 2330 2104 2331
rect 2242 2335 2248 2336
rect 2242 2331 2243 2335
rect 2247 2331 2248 2335
rect 2242 2330 2248 2331
rect 2434 2335 2440 2336
rect 2434 2331 2435 2335
rect 2439 2331 2440 2335
rect 2434 2330 2440 2331
rect 2458 2335 2464 2336
rect 2458 2331 2459 2335
rect 2463 2331 2464 2335
rect 2458 2330 2464 2331
rect 2754 2335 2760 2336
rect 2754 2331 2755 2335
rect 2759 2331 2760 2335
rect 2754 2330 2760 2331
rect 2890 2335 2896 2336
rect 2890 2331 2891 2335
rect 2895 2331 2896 2335
rect 2890 2330 2896 2331
rect 3030 2335 3036 2336
rect 3030 2331 3031 2335
rect 3035 2331 3036 2335
rect 3030 2330 3036 2331
rect 1870 2324 1876 2325
rect 1870 2320 1871 2324
rect 1875 2320 1876 2324
rect 1870 2319 1876 2320
rect 1830 2312 1836 2313
rect 1830 2308 1831 2312
rect 1835 2308 1836 2312
rect 1830 2307 1836 2308
rect 1458 2303 1464 2304
rect 1458 2299 1459 2303
rect 1463 2299 1464 2303
rect 1458 2298 1464 2299
rect 1558 2303 1564 2304
rect 1558 2299 1559 2303
rect 1563 2299 1564 2303
rect 1558 2298 1564 2299
rect 1618 2303 1624 2304
rect 1618 2299 1619 2303
rect 1623 2299 1624 2303
rect 1618 2298 1624 2299
rect 110 2295 116 2296
rect 110 2291 111 2295
rect 115 2291 116 2295
rect 1830 2295 1836 2296
rect 110 2290 116 2291
rect 1398 2292 1404 2293
rect 112 2263 114 2290
rect 1398 2288 1399 2292
rect 1403 2288 1404 2292
rect 1398 2287 1404 2288
rect 1478 2292 1484 2293
rect 1478 2288 1479 2292
rect 1483 2288 1484 2292
rect 1478 2287 1484 2288
rect 1558 2292 1564 2293
rect 1558 2288 1559 2292
rect 1563 2288 1564 2292
rect 1558 2287 1564 2288
rect 1638 2292 1644 2293
rect 1638 2288 1639 2292
rect 1643 2288 1644 2292
rect 1830 2291 1831 2295
rect 1835 2291 1836 2295
rect 1872 2291 1874 2319
rect 1902 2306 1908 2307
rect 1902 2302 1903 2306
rect 1907 2302 1908 2306
rect 1902 2301 1908 2302
rect 1904 2291 1906 2301
rect 1964 2296 1966 2330
rect 2022 2306 2028 2307
rect 2022 2302 2023 2306
rect 2027 2302 2028 2306
rect 2022 2301 2028 2302
rect 1910 2295 1916 2296
rect 1910 2291 1911 2295
rect 1915 2291 1916 2295
rect 1830 2290 1836 2291
rect 1871 2290 1875 2291
rect 1638 2287 1644 2288
rect 1400 2263 1402 2287
rect 1480 2263 1482 2287
rect 1560 2263 1562 2287
rect 1578 2275 1584 2276
rect 1578 2271 1579 2275
rect 1583 2271 1584 2275
rect 1578 2270 1584 2271
rect 111 2262 115 2263
rect 111 2257 115 2258
rect 135 2262 139 2263
rect 135 2257 139 2258
rect 215 2262 219 2263
rect 215 2257 219 2258
rect 295 2262 299 2263
rect 295 2257 299 2258
rect 383 2262 387 2263
rect 383 2257 387 2258
rect 519 2262 523 2263
rect 519 2257 523 2258
rect 671 2262 675 2263
rect 671 2257 675 2258
rect 831 2262 835 2263
rect 831 2257 835 2258
rect 999 2262 1003 2263
rect 999 2257 1003 2258
rect 1159 2262 1163 2263
rect 1159 2257 1163 2258
rect 1311 2262 1315 2263
rect 1311 2257 1315 2258
rect 1399 2262 1403 2263
rect 1399 2257 1403 2258
rect 1455 2262 1459 2263
rect 1455 2257 1459 2258
rect 1479 2262 1483 2263
rect 1479 2257 1483 2258
rect 1559 2262 1563 2263
rect 1559 2257 1563 2258
rect 112 2238 114 2257
rect 136 2241 138 2257
rect 216 2241 218 2257
rect 296 2241 298 2257
rect 384 2241 386 2257
rect 520 2241 522 2257
rect 672 2241 674 2257
rect 832 2241 834 2257
rect 1000 2241 1002 2257
rect 1160 2241 1162 2257
rect 1175 2244 1179 2245
rect 134 2240 140 2241
rect 110 2237 116 2238
rect 110 2233 111 2237
rect 115 2233 116 2237
rect 134 2236 135 2240
rect 139 2236 140 2240
rect 134 2235 140 2236
rect 214 2240 220 2241
rect 214 2236 215 2240
rect 219 2236 220 2240
rect 214 2235 220 2236
rect 294 2240 300 2241
rect 294 2236 295 2240
rect 299 2236 300 2240
rect 294 2235 300 2236
rect 382 2240 388 2241
rect 382 2236 383 2240
rect 387 2236 388 2240
rect 382 2235 388 2236
rect 518 2240 524 2241
rect 518 2236 519 2240
rect 523 2236 524 2240
rect 518 2235 524 2236
rect 670 2240 676 2241
rect 670 2236 671 2240
rect 675 2236 676 2240
rect 670 2235 676 2236
rect 830 2240 836 2241
rect 830 2236 831 2240
rect 835 2236 836 2240
rect 830 2235 836 2236
rect 998 2240 1004 2241
rect 998 2236 999 2240
rect 1003 2236 1004 2240
rect 998 2235 1004 2236
rect 1158 2240 1164 2241
rect 1158 2236 1159 2240
rect 1163 2236 1164 2240
rect 1312 2241 1314 2257
rect 1456 2241 1458 2257
rect 1580 2245 1582 2270
rect 1640 2263 1642 2287
rect 1832 2263 1834 2290
rect 1871 2285 1875 2286
rect 1903 2290 1907 2291
rect 1910 2290 1916 2291
rect 1962 2295 1968 2296
rect 1962 2291 1963 2295
rect 1967 2291 1968 2295
rect 2024 2291 2026 2301
rect 2100 2296 2102 2330
rect 2182 2306 2188 2307
rect 2182 2302 2183 2306
rect 2187 2302 2188 2306
rect 2182 2301 2188 2302
rect 2098 2295 2104 2296
rect 2098 2291 2099 2295
rect 2103 2291 2104 2295
rect 2184 2291 2186 2301
rect 2244 2296 2246 2330
rect 2350 2306 2356 2307
rect 2350 2302 2351 2306
rect 2355 2302 2356 2306
rect 2350 2301 2356 2302
rect 2242 2295 2248 2296
rect 2242 2291 2243 2295
rect 2247 2291 2248 2295
rect 2352 2291 2354 2301
rect 2436 2296 2438 2330
rect 2518 2306 2524 2307
rect 2518 2302 2519 2306
rect 2523 2302 2524 2306
rect 2518 2301 2524 2302
rect 2678 2306 2684 2307
rect 2678 2302 2679 2306
rect 2683 2302 2684 2306
rect 2678 2301 2684 2302
rect 2434 2295 2440 2296
rect 2434 2291 2435 2295
rect 2439 2291 2440 2295
rect 2520 2291 2522 2301
rect 2680 2291 2682 2301
rect 2687 2300 2691 2301
rect 2756 2296 2758 2330
rect 2830 2306 2836 2307
rect 2830 2302 2831 2306
rect 2835 2302 2836 2306
rect 2830 2301 2836 2302
rect 2686 2295 2692 2296
rect 2686 2291 2687 2295
rect 2691 2291 2692 2295
rect 1962 2290 1968 2291
rect 2023 2290 2027 2291
rect 1903 2285 1907 2286
rect 1607 2262 1611 2263
rect 1607 2257 1611 2258
rect 1639 2262 1643 2263
rect 1639 2257 1643 2258
rect 1743 2262 1747 2263
rect 1743 2257 1747 2258
rect 1831 2262 1835 2263
rect 1831 2257 1835 2258
rect 1872 2257 1874 2285
rect 1904 2275 1906 2285
rect 1902 2274 1908 2275
rect 1902 2270 1903 2274
rect 1907 2270 1908 2274
rect 1902 2269 1908 2270
rect 1579 2244 1583 2245
rect 1175 2239 1179 2240
rect 1310 2240 1316 2241
rect 1158 2235 1164 2236
rect 110 2232 116 2233
rect 202 2231 208 2232
rect 202 2227 203 2231
rect 207 2227 208 2231
rect 202 2226 208 2227
rect 282 2231 288 2232
rect 282 2227 283 2231
rect 287 2227 288 2231
rect 282 2226 288 2227
rect 362 2231 368 2232
rect 362 2227 363 2231
rect 367 2227 368 2231
rect 362 2226 368 2227
rect 458 2231 464 2232
rect 458 2227 459 2231
rect 463 2227 464 2231
rect 458 2226 464 2227
rect 586 2231 592 2232
rect 586 2227 587 2231
rect 591 2227 592 2231
rect 586 2226 592 2227
rect 754 2231 760 2232
rect 754 2227 755 2231
rect 759 2227 760 2231
rect 754 2226 760 2227
rect 922 2231 928 2232
rect 922 2227 923 2231
rect 927 2227 928 2231
rect 922 2226 928 2227
rect 998 2227 1004 2228
rect 110 2220 116 2221
rect 110 2216 111 2220
rect 115 2216 116 2220
rect 110 2215 116 2216
rect 112 2183 114 2215
rect 142 2202 148 2203
rect 142 2198 143 2202
rect 147 2198 148 2202
rect 142 2197 148 2198
rect 144 2183 146 2197
rect 204 2192 206 2226
rect 222 2202 228 2203
rect 222 2198 223 2202
rect 227 2198 228 2202
rect 222 2197 228 2198
rect 202 2191 208 2192
rect 202 2187 203 2191
rect 207 2187 208 2191
rect 202 2186 208 2187
rect 224 2183 226 2197
rect 284 2192 286 2226
rect 302 2202 308 2203
rect 302 2198 303 2202
rect 307 2198 308 2202
rect 302 2197 308 2198
rect 282 2191 288 2192
rect 282 2187 283 2191
rect 287 2187 288 2191
rect 282 2186 288 2187
rect 304 2183 306 2197
rect 364 2192 366 2226
rect 390 2202 396 2203
rect 390 2198 391 2202
rect 395 2198 396 2202
rect 390 2197 396 2198
rect 362 2191 368 2192
rect 362 2187 363 2191
rect 367 2187 368 2191
rect 362 2186 368 2187
rect 392 2183 394 2197
rect 460 2192 462 2226
rect 526 2202 532 2203
rect 526 2198 527 2202
rect 531 2198 532 2202
rect 526 2197 532 2198
rect 458 2191 464 2192
rect 458 2187 459 2191
rect 463 2187 464 2191
rect 458 2186 464 2187
rect 528 2183 530 2197
rect 588 2192 590 2226
rect 678 2202 684 2203
rect 678 2198 679 2202
rect 683 2198 684 2202
rect 678 2197 684 2198
rect 586 2191 592 2192
rect 586 2187 587 2191
rect 591 2187 592 2191
rect 586 2186 592 2187
rect 680 2183 682 2197
rect 756 2192 758 2226
rect 838 2202 844 2203
rect 838 2198 839 2202
rect 843 2198 844 2202
rect 838 2197 844 2198
rect 754 2191 760 2192
rect 754 2187 755 2191
rect 759 2187 760 2191
rect 754 2186 760 2187
rect 840 2183 842 2197
rect 924 2192 926 2226
rect 998 2223 999 2227
rect 1003 2223 1004 2227
rect 998 2222 1004 2223
rect 922 2191 928 2192
rect 922 2187 923 2191
rect 927 2187 928 2191
rect 922 2186 928 2187
rect 111 2182 115 2183
rect 111 2177 115 2178
rect 143 2182 147 2183
rect 143 2177 147 2178
rect 191 2182 195 2183
rect 191 2177 195 2178
rect 223 2182 227 2183
rect 223 2177 227 2178
rect 303 2182 307 2183
rect 303 2177 307 2178
rect 311 2182 315 2183
rect 311 2177 315 2178
rect 391 2182 395 2183
rect 391 2177 395 2178
rect 463 2182 467 2183
rect 463 2177 467 2178
rect 527 2182 531 2183
rect 527 2177 531 2178
rect 639 2182 643 2183
rect 639 2177 643 2178
rect 679 2182 683 2183
rect 679 2177 683 2178
rect 823 2182 827 2183
rect 823 2177 827 2178
rect 839 2182 843 2183
rect 839 2177 843 2178
rect 112 2149 114 2177
rect 192 2167 194 2177
rect 198 2175 204 2176
rect 198 2170 199 2175
rect 203 2170 204 2175
rect 282 2175 288 2176
rect 282 2171 283 2175
rect 287 2171 288 2175
rect 282 2170 288 2171
rect 199 2167 203 2168
rect 190 2166 196 2167
rect 190 2162 191 2166
rect 195 2162 196 2166
rect 190 2161 196 2162
rect 110 2148 116 2149
rect 110 2144 111 2148
rect 115 2144 116 2148
rect 110 2143 116 2144
rect 110 2131 116 2132
rect 110 2127 111 2131
rect 115 2127 116 2131
rect 110 2126 116 2127
rect 182 2128 188 2129
rect 112 2103 114 2126
rect 182 2124 183 2128
rect 187 2124 188 2128
rect 182 2123 188 2124
rect 184 2103 186 2123
rect 111 2102 115 2103
rect 111 2097 115 2098
rect 183 2102 187 2103
rect 183 2097 187 2098
rect 215 2102 219 2103
rect 215 2097 219 2098
rect 112 2078 114 2097
rect 216 2081 218 2097
rect 214 2080 220 2081
rect 110 2077 116 2078
rect 110 2073 111 2077
rect 115 2073 116 2077
rect 214 2076 215 2080
rect 219 2076 220 2080
rect 214 2075 220 2076
rect 110 2072 116 2073
rect 284 2072 286 2170
rect 312 2167 314 2177
rect 362 2175 368 2176
rect 362 2171 363 2175
rect 367 2171 368 2175
rect 362 2170 368 2171
rect 310 2166 316 2167
rect 310 2162 311 2166
rect 315 2162 316 2166
rect 310 2161 316 2162
rect 364 2140 366 2170
rect 464 2167 466 2177
rect 471 2172 475 2173
rect 471 2167 475 2168
rect 640 2167 642 2177
rect 646 2175 652 2176
rect 646 2170 647 2175
rect 651 2170 652 2175
rect 690 2175 696 2176
rect 690 2171 691 2175
rect 695 2171 696 2175
rect 690 2170 696 2171
rect 647 2167 651 2168
rect 462 2166 468 2167
rect 462 2162 463 2166
rect 467 2162 468 2166
rect 462 2161 468 2162
rect 472 2140 474 2167
rect 638 2166 644 2167
rect 638 2162 639 2166
rect 643 2162 644 2166
rect 638 2161 644 2162
rect 692 2140 694 2170
rect 824 2167 826 2177
rect 1000 2176 1002 2222
rect 1006 2202 1012 2203
rect 1006 2198 1007 2202
rect 1011 2198 1012 2202
rect 1006 2197 1012 2198
rect 1166 2202 1172 2203
rect 1166 2198 1167 2202
rect 1171 2198 1172 2202
rect 1166 2197 1172 2198
rect 1008 2183 1010 2197
rect 1168 2183 1170 2197
rect 1176 2192 1178 2239
rect 1310 2236 1311 2240
rect 1315 2236 1316 2240
rect 1310 2235 1316 2236
rect 1454 2240 1460 2241
rect 1454 2236 1455 2240
rect 1459 2236 1460 2240
rect 1608 2241 1610 2257
rect 1744 2241 1746 2257
rect 1579 2239 1583 2240
rect 1606 2240 1612 2241
rect 1454 2235 1460 2236
rect 1606 2236 1607 2240
rect 1611 2236 1612 2240
rect 1606 2235 1612 2236
rect 1742 2240 1748 2241
rect 1742 2236 1743 2240
rect 1747 2236 1748 2240
rect 1832 2238 1834 2257
rect 1870 2256 1876 2257
rect 1870 2252 1871 2256
rect 1875 2252 1876 2256
rect 1870 2251 1876 2252
rect 1912 2248 1914 2290
rect 2023 2285 2027 2286
rect 2031 2290 2035 2291
rect 2098 2290 2104 2291
rect 2183 2290 2187 2291
rect 2242 2290 2248 2291
rect 2351 2290 2355 2291
rect 2031 2285 2035 2286
rect 2183 2285 2187 2286
rect 2351 2285 2355 2286
rect 2367 2290 2371 2291
rect 2434 2290 2440 2291
rect 2519 2290 2523 2291
rect 2367 2285 2371 2286
rect 2519 2285 2523 2286
rect 2575 2290 2579 2291
rect 2575 2285 2579 2286
rect 2679 2290 2683 2291
rect 2686 2290 2692 2291
rect 2754 2295 2760 2296
rect 2754 2291 2755 2295
rect 2759 2291 2760 2295
rect 2832 2291 2834 2301
rect 2892 2296 2894 2330
rect 2966 2306 2972 2307
rect 2966 2302 2967 2306
rect 2971 2302 2972 2306
rect 2966 2301 2972 2302
rect 2890 2295 2896 2296
rect 2890 2291 2891 2295
rect 2895 2291 2896 2295
rect 2968 2291 2970 2301
rect 3032 2296 3034 2330
rect 3086 2306 3092 2307
rect 3086 2302 3087 2306
rect 3091 2302 3092 2306
rect 3086 2301 3092 2302
rect 3140 2301 3142 2374
rect 3208 2367 3210 2391
rect 3592 2367 3594 2394
rect 3191 2366 3195 2367
rect 3191 2361 3195 2362
rect 3207 2366 3211 2367
rect 3207 2361 3211 2362
rect 3303 2366 3307 2367
rect 3303 2361 3307 2362
rect 3415 2366 3419 2367
rect 3415 2361 3419 2362
rect 3503 2366 3507 2367
rect 3503 2361 3507 2362
rect 3591 2366 3595 2367
rect 3591 2361 3595 2362
rect 3192 2345 3194 2361
rect 3304 2345 3306 2361
rect 3416 2345 3418 2361
rect 3504 2345 3506 2361
rect 3190 2344 3196 2345
rect 3190 2340 3191 2344
rect 3195 2340 3196 2344
rect 3190 2339 3196 2340
rect 3302 2344 3308 2345
rect 3302 2340 3303 2344
rect 3307 2340 3308 2344
rect 3302 2339 3308 2340
rect 3414 2344 3420 2345
rect 3414 2340 3415 2344
rect 3419 2340 3420 2344
rect 3414 2339 3420 2340
rect 3502 2344 3508 2345
rect 3502 2340 3503 2344
rect 3507 2340 3508 2344
rect 3592 2342 3594 2361
rect 3502 2339 3508 2340
rect 3590 2341 3596 2342
rect 3590 2337 3591 2341
rect 3595 2337 3596 2341
rect 3590 2336 3596 2337
rect 3146 2335 3152 2336
rect 3146 2331 3147 2335
rect 3151 2331 3152 2335
rect 3146 2330 3152 2331
rect 3262 2335 3268 2336
rect 3262 2331 3263 2335
rect 3267 2331 3268 2335
rect 3262 2330 3268 2331
rect 3370 2335 3376 2336
rect 3370 2331 3371 2335
rect 3375 2331 3376 2335
rect 3370 2330 3376 2331
rect 3482 2335 3488 2336
rect 3482 2331 3483 2335
rect 3487 2331 3488 2335
rect 3482 2330 3488 2331
rect 3030 2295 3036 2296
rect 3030 2291 3031 2295
rect 3035 2291 3036 2295
rect 3088 2291 3090 2301
rect 3139 2300 3143 2301
rect 3148 2296 3150 2330
rect 3198 2306 3204 2307
rect 3198 2302 3199 2306
rect 3203 2302 3204 2306
rect 3198 2301 3204 2302
rect 3139 2295 3143 2296
rect 3146 2295 3152 2296
rect 3146 2291 3147 2295
rect 3151 2291 3152 2295
rect 3200 2291 3202 2301
rect 3264 2296 3266 2330
rect 3310 2306 3316 2307
rect 3310 2302 3311 2306
rect 3315 2302 3316 2306
rect 3310 2301 3316 2302
rect 3262 2295 3268 2296
rect 3262 2291 3263 2295
rect 3267 2291 3268 2295
rect 3312 2291 3314 2301
rect 3372 2296 3374 2330
rect 3422 2306 3428 2307
rect 3422 2302 3423 2306
rect 3427 2302 3428 2306
rect 3422 2301 3428 2302
rect 3370 2295 3376 2296
rect 3370 2291 3371 2295
rect 3375 2291 3376 2295
rect 3424 2291 3426 2301
rect 3484 2296 3486 2330
rect 3590 2324 3596 2325
rect 3590 2320 3591 2324
rect 3595 2320 3596 2324
rect 3590 2319 3596 2320
rect 3510 2306 3516 2307
rect 3510 2302 3511 2306
rect 3515 2302 3516 2306
rect 3510 2301 3516 2302
rect 3482 2295 3488 2296
rect 3482 2291 3483 2295
rect 3487 2291 3488 2295
rect 3512 2291 3514 2301
rect 3592 2291 3594 2319
rect 2754 2290 2760 2291
rect 2791 2290 2795 2291
rect 2679 2285 2683 2286
rect 2791 2285 2795 2286
rect 2831 2290 2835 2291
rect 2890 2290 2896 2291
rect 2967 2290 2971 2291
rect 2831 2285 2835 2286
rect 2967 2285 2971 2286
rect 3023 2290 3027 2291
rect 3030 2290 3036 2291
rect 3087 2290 3091 2291
rect 3146 2290 3152 2291
rect 3199 2290 3203 2291
rect 3023 2285 3027 2286
rect 3087 2285 3091 2286
rect 3199 2285 3203 2286
rect 3255 2290 3259 2291
rect 3262 2290 3268 2291
rect 3311 2290 3315 2291
rect 3370 2290 3376 2291
rect 3423 2290 3427 2291
rect 3482 2290 3488 2291
rect 3495 2290 3499 2291
rect 3255 2285 3259 2286
rect 3311 2285 3315 2286
rect 3342 2287 3348 2288
rect 1962 2283 1968 2284
rect 1962 2279 1963 2283
rect 1967 2279 1968 2283
rect 1962 2278 1968 2279
rect 1964 2248 1966 2278
rect 2032 2275 2034 2285
rect 2184 2275 2186 2285
rect 2368 2275 2370 2285
rect 2374 2283 2380 2284
rect 2374 2279 2375 2283
rect 2379 2279 2380 2283
rect 2374 2278 2380 2279
rect 2478 2283 2484 2284
rect 2478 2279 2479 2283
rect 2483 2279 2484 2283
rect 2478 2278 2484 2279
rect 2030 2274 2036 2275
rect 2030 2270 2031 2274
rect 2035 2270 2036 2274
rect 2030 2269 2036 2270
rect 2182 2274 2188 2275
rect 2182 2270 2183 2274
rect 2187 2270 2188 2274
rect 2182 2269 2188 2270
rect 2366 2274 2372 2275
rect 2366 2270 2367 2274
rect 2371 2270 2372 2274
rect 2366 2269 2372 2270
rect 1910 2247 1916 2248
rect 1910 2243 1911 2247
rect 1915 2243 1916 2247
rect 1910 2242 1916 2243
rect 1962 2247 1968 2248
rect 1962 2243 1963 2247
rect 1967 2243 1968 2247
rect 1962 2242 1968 2243
rect 1870 2239 1876 2240
rect 1742 2235 1748 2236
rect 1830 2237 1836 2238
rect 1830 2233 1831 2237
rect 1835 2233 1836 2237
rect 1870 2235 1871 2239
rect 1875 2235 1876 2239
rect 1870 2234 1876 2235
rect 1894 2236 1900 2237
rect 1830 2232 1836 2233
rect 1234 2231 1240 2232
rect 1234 2227 1235 2231
rect 1239 2227 1240 2231
rect 1234 2226 1240 2227
rect 1378 2231 1384 2232
rect 1378 2227 1379 2231
rect 1383 2227 1384 2231
rect 1378 2226 1384 2227
rect 1530 2231 1536 2232
rect 1530 2227 1531 2231
rect 1535 2227 1536 2231
rect 1530 2226 1536 2227
rect 1682 2231 1688 2232
rect 1682 2227 1683 2231
rect 1687 2227 1688 2231
rect 1682 2226 1688 2227
rect 1690 2231 1696 2232
rect 1690 2227 1691 2231
rect 1695 2227 1696 2231
rect 1690 2226 1696 2227
rect 1207 2196 1211 2197
rect 1236 2192 1238 2226
rect 1318 2202 1324 2203
rect 1318 2198 1319 2202
rect 1323 2198 1324 2202
rect 1318 2197 1324 2198
rect 1174 2191 1180 2192
rect 1207 2191 1211 2192
rect 1234 2191 1240 2192
rect 1174 2187 1175 2191
rect 1179 2187 1180 2191
rect 1174 2186 1180 2187
rect 1007 2182 1011 2183
rect 1007 2177 1011 2178
rect 1015 2182 1019 2183
rect 1015 2177 1019 2178
rect 1167 2182 1171 2183
rect 1167 2177 1171 2178
rect 1199 2182 1203 2183
rect 1199 2177 1203 2178
rect 998 2175 1004 2176
rect 998 2171 999 2175
rect 1003 2171 1004 2175
rect 998 2170 1004 2171
rect 1016 2167 1018 2177
rect 1023 2172 1027 2173
rect 1023 2167 1027 2168
rect 1200 2167 1202 2177
rect 1208 2176 1210 2191
rect 1234 2187 1235 2191
rect 1239 2187 1240 2191
rect 1234 2186 1240 2187
rect 1320 2183 1322 2197
rect 1380 2192 1382 2226
rect 1462 2202 1468 2203
rect 1462 2198 1463 2202
rect 1467 2198 1468 2202
rect 1462 2197 1468 2198
rect 1378 2191 1384 2192
rect 1378 2187 1379 2191
rect 1383 2187 1384 2191
rect 1378 2186 1384 2187
rect 1464 2183 1466 2197
rect 1532 2192 1534 2226
rect 1614 2202 1620 2203
rect 1614 2198 1615 2202
rect 1619 2198 1620 2202
rect 1614 2197 1620 2198
rect 1530 2191 1536 2192
rect 1530 2187 1531 2191
rect 1535 2187 1536 2191
rect 1530 2186 1536 2187
rect 1616 2183 1618 2197
rect 1684 2192 1686 2226
rect 1692 2197 1694 2226
rect 1830 2220 1836 2221
rect 1830 2216 1831 2220
rect 1835 2216 1836 2220
rect 1830 2215 1836 2216
rect 1750 2202 1756 2203
rect 1750 2198 1751 2202
rect 1755 2198 1756 2202
rect 1750 2197 1756 2198
rect 1691 2196 1695 2197
rect 1682 2191 1688 2192
rect 1691 2191 1695 2192
rect 1682 2187 1683 2191
rect 1687 2187 1688 2191
rect 1682 2186 1688 2187
rect 1752 2183 1754 2197
rect 1832 2183 1834 2215
rect 1872 2195 1874 2234
rect 1894 2232 1895 2236
rect 1899 2232 1900 2236
rect 1894 2231 1900 2232
rect 2022 2236 2028 2237
rect 2022 2232 2023 2236
rect 2027 2232 2028 2236
rect 2022 2231 2028 2232
rect 2174 2236 2180 2237
rect 2174 2232 2175 2236
rect 2179 2232 2180 2236
rect 2174 2231 2180 2232
rect 2358 2236 2364 2237
rect 2358 2232 2359 2236
rect 2363 2232 2364 2236
rect 2358 2231 2364 2232
rect 1896 2195 1898 2231
rect 2024 2195 2026 2231
rect 2176 2195 2178 2231
rect 2360 2195 2362 2231
rect 2376 2220 2378 2278
rect 2374 2219 2380 2220
rect 2374 2215 2375 2219
rect 2379 2215 2380 2219
rect 2374 2214 2380 2215
rect 1871 2194 1875 2195
rect 1871 2189 1875 2190
rect 1895 2194 1899 2195
rect 1895 2189 1899 2190
rect 2023 2194 2027 2195
rect 2023 2189 2027 2190
rect 2175 2194 2179 2195
rect 2175 2189 2179 2190
rect 2199 2194 2203 2195
rect 2199 2189 2203 2190
rect 2295 2194 2299 2195
rect 2295 2189 2299 2190
rect 2359 2194 2363 2195
rect 2359 2189 2363 2190
rect 2399 2194 2403 2195
rect 2399 2189 2403 2190
rect 1319 2182 1323 2183
rect 1319 2177 1323 2178
rect 1391 2182 1395 2183
rect 1391 2177 1395 2178
rect 1463 2182 1467 2183
rect 1463 2177 1467 2178
rect 1583 2182 1587 2183
rect 1583 2177 1587 2178
rect 1615 2182 1619 2183
rect 1615 2177 1619 2178
rect 1751 2182 1755 2183
rect 1751 2177 1755 2178
rect 1831 2182 1835 2183
rect 1831 2177 1835 2178
rect 1206 2175 1212 2176
rect 1206 2171 1207 2175
rect 1211 2171 1212 2175
rect 1206 2170 1212 2171
rect 1250 2175 1256 2176
rect 1250 2171 1251 2175
rect 1255 2171 1256 2175
rect 1250 2170 1256 2171
rect 822 2166 828 2167
rect 822 2162 823 2166
rect 827 2162 828 2166
rect 822 2161 828 2162
rect 1014 2166 1020 2167
rect 1014 2162 1015 2166
rect 1019 2162 1020 2166
rect 1014 2161 1020 2162
rect 1024 2140 1026 2167
rect 1198 2166 1204 2167
rect 1198 2162 1199 2166
rect 1203 2162 1204 2166
rect 1198 2161 1204 2162
rect 1252 2140 1254 2170
rect 1392 2167 1394 2177
rect 1442 2175 1448 2176
rect 1442 2171 1443 2175
rect 1447 2171 1448 2175
rect 1442 2170 1448 2171
rect 1390 2166 1396 2167
rect 1390 2162 1391 2166
rect 1395 2162 1396 2166
rect 1390 2161 1396 2162
rect 1444 2140 1446 2170
rect 1584 2167 1586 2177
rect 1634 2175 1640 2176
rect 1634 2171 1635 2175
rect 1639 2171 1640 2175
rect 1634 2170 1640 2171
rect 1582 2166 1588 2167
rect 1582 2162 1583 2166
rect 1587 2162 1588 2166
rect 1582 2161 1588 2162
rect 1636 2140 1638 2170
rect 1752 2167 1754 2177
rect 1750 2166 1756 2167
rect 1750 2162 1751 2166
rect 1755 2162 1756 2166
rect 1750 2161 1756 2162
rect 1832 2149 1834 2177
rect 1872 2170 1874 2189
rect 2200 2173 2202 2189
rect 2296 2173 2298 2189
rect 2400 2173 2402 2189
rect 2198 2172 2204 2173
rect 1870 2169 1876 2170
rect 1870 2165 1871 2169
rect 1875 2165 1876 2169
rect 2198 2168 2199 2172
rect 2203 2168 2204 2172
rect 2198 2167 2204 2168
rect 2294 2172 2300 2173
rect 2294 2168 2295 2172
rect 2299 2168 2300 2172
rect 2294 2167 2300 2168
rect 2398 2172 2404 2173
rect 2398 2168 2399 2172
rect 2403 2168 2404 2172
rect 2398 2167 2404 2168
rect 1870 2164 1876 2165
rect 2480 2164 2482 2278
rect 2576 2275 2578 2285
rect 2626 2283 2632 2284
rect 2626 2279 2627 2283
rect 2631 2279 2632 2283
rect 2626 2278 2632 2279
rect 2574 2274 2580 2275
rect 2574 2270 2575 2274
rect 2579 2270 2580 2274
rect 2574 2269 2580 2270
rect 2628 2248 2630 2278
rect 2792 2275 2794 2285
rect 3024 2275 3026 2285
rect 3074 2283 3080 2284
rect 3074 2279 3075 2283
rect 3079 2279 3080 2283
rect 3074 2278 3080 2279
rect 2790 2274 2796 2275
rect 2790 2270 2791 2274
rect 2795 2270 2796 2274
rect 2790 2269 2796 2270
rect 3022 2274 3028 2275
rect 3022 2270 3023 2274
rect 3027 2270 3028 2274
rect 3022 2269 3028 2270
rect 3076 2248 3078 2278
rect 3256 2275 3258 2285
rect 3342 2283 3343 2287
rect 3347 2283 3348 2287
rect 3423 2285 3427 2286
rect 3495 2285 3499 2286
rect 3511 2290 3515 2291
rect 3511 2285 3515 2286
rect 3591 2290 3595 2291
rect 3591 2285 3595 2286
rect 3342 2282 3348 2283
rect 3254 2274 3260 2275
rect 3254 2270 3255 2274
rect 3259 2270 3260 2274
rect 3254 2269 3260 2270
rect 3344 2248 3346 2282
rect 3496 2275 3498 2285
rect 3494 2274 3500 2275
rect 3494 2270 3495 2274
rect 3499 2270 3500 2274
rect 3494 2269 3500 2270
rect 3592 2257 3594 2285
rect 3590 2256 3596 2257
rect 3590 2252 3591 2256
rect 3595 2252 3596 2256
rect 3590 2251 3596 2252
rect 2626 2247 2632 2248
rect 2626 2243 2627 2247
rect 2631 2243 2632 2247
rect 2626 2242 2632 2243
rect 3074 2247 3080 2248
rect 3074 2243 3075 2247
rect 3079 2243 3080 2247
rect 3074 2242 3080 2243
rect 3334 2247 3340 2248
rect 3334 2243 3335 2247
rect 3339 2243 3340 2247
rect 3334 2242 3340 2243
rect 3342 2247 3348 2248
rect 3342 2243 3343 2247
rect 3347 2243 3348 2247
rect 3342 2242 3348 2243
rect 2566 2236 2572 2237
rect 2566 2232 2567 2236
rect 2571 2232 2572 2236
rect 2566 2231 2572 2232
rect 2782 2236 2788 2237
rect 2782 2232 2783 2236
rect 2787 2232 2788 2236
rect 2782 2231 2788 2232
rect 3014 2236 3020 2237
rect 3014 2232 3015 2236
rect 3019 2232 3020 2236
rect 3014 2231 3020 2232
rect 3246 2236 3252 2237
rect 3246 2232 3247 2236
rect 3251 2232 3252 2236
rect 3246 2231 3252 2232
rect 2568 2195 2570 2231
rect 2784 2195 2786 2231
rect 3016 2195 3018 2231
rect 3248 2195 3250 2231
rect 2519 2194 2523 2195
rect 2519 2189 2523 2190
rect 2567 2194 2571 2195
rect 2567 2189 2571 2190
rect 2639 2194 2643 2195
rect 2639 2189 2643 2190
rect 2759 2194 2763 2195
rect 2759 2189 2763 2190
rect 2783 2194 2787 2195
rect 2783 2189 2787 2190
rect 2879 2194 2883 2195
rect 2879 2189 2883 2190
rect 2991 2194 2995 2195
rect 2991 2189 2995 2190
rect 3015 2194 3019 2195
rect 3015 2189 3019 2190
rect 3095 2194 3099 2195
rect 3095 2189 3099 2190
rect 3199 2194 3203 2195
rect 3199 2189 3203 2190
rect 3247 2194 3251 2195
rect 3247 2189 3251 2190
rect 3303 2194 3307 2195
rect 3303 2189 3307 2190
rect 2520 2173 2522 2189
rect 2640 2173 2642 2189
rect 2760 2173 2762 2189
rect 2880 2173 2882 2189
rect 2992 2173 2994 2189
rect 3096 2173 3098 2189
rect 3200 2173 3202 2189
rect 3304 2173 3306 2189
rect 2518 2172 2524 2173
rect 2518 2168 2519 2172
rect 2523 2168 2524 2172
rect 2518 2167 2524 2168
rect 2638 2172 2644 2173
rect 2638 2168 2639 2172
rect 2643 2168 2644 2172
rect 2638 2167 2644 2168
rect 2758 2172 2764 2173
rect 2758 2168 2759 2172
rect 2763 2168 2764 2172
rect 2758 2167 2764 2168
rect 2878 2172 2884 2173
rect 2878 2168 2879 2172
rect 2883 2168 2884 2172
rect 2878 2167 2884 2168
rect 2990 2172 2996 2173
rect 2990 2168 2991 2172
rect 2995 2168 2996 2172
rect 2990 2167 2996 2168
rect 3094 2172 3100 2173
rect 3094 2168 3095 2172
rect 3099 2168 3100 2172
rect 3094 2167 3100 2168
rect 3198 2172 3204 2173
rect 3198 2168 3199 2172
rect 3203 2168 3204 2172
rect 3198 2167 3204 2168
rect 3302 2172 3308 2173
rect 3302 2168 3303 2172
rect 3307 2168 3308 2172
rect 3302 2167 3308 2168
rect 2266 2163 2272 2164
rect 2266 2159 2267 2163
rect 2271 2159 2272 2163
rect 2266 2158 2272 2159
rect 2362 2163 2368 2164
rect 2362 2159 2363 2163
rect 2367 2159 2368 2163
rect 2362 2158 2368 2159
rect 2478 2163 2484 2164
rect 2478 2159 2479 2163
rect 2483 2159 2484 2163
rect 2478 2158 2484 2159
rect 2486 2163 2492 2164
rect 2486 2159 2487 2163
rect 2491 2159 2492 2163
rect 2486 2158 2492 2159
rect 2586 2163 2592 2164
rect 2586 2159 2587 2163
rect 2591 2159 2592 2163
rect 2586 2158 2592 2159
rect 2706 2163 2712 2164
rect 2706 2159 2707 2163
rect 2711 2159 2712 2163
rect 2706 2158 2712 2159
rect 2946 2163 2952 2164
rect 2946 2159 2947 2163
rect 2951 2159 2952 2163
rect 2946 2158 2952 2159
rect 3058 2163 3064 2164
rect 3058 2159 3059 2163
rect 3063 2159 3064 2163
rect 3058 2158 3064 2159
rect 3174 2163 3180 2164
rect 3174 2159 3175 2163
rect 3179 2159 3180 2163
rect 3174 2158 3180 2159
rect 3266 2163 3272 2164
rect 3266 2159 3267 2163
rect 3271 2159 3272 2163
rect 3266 2158 3272 2159
rect 1870 2152 1876 2153
rect 1830 2148 1836 2149
rect 1830 2144 1831 2148
rect 1835 2144 1836 2148
rect 1870 2148 1871 2152
rect 1875 2148 1876 2152
rect 1870 2147 1876 2148
rect 1830 2143 1836 2144
rect 362 2139 368 2140
rect 362 2135 363 2139
rect 367 2135 368 2139
rect 362 2134 368 2135
rect 470 2139 476 2140
rect 470 2135 471 2139
rect 475 2135 476 2139
rect 470 2134 476 2135
rect 690 2139 696 2140
rect 690 2135 691 2139
rect 695 2135 696 2139
rect 690 2134 696 2135
rect 874 2139 880 2140
rect 874 2135 875 2139
rect 879 2135 880 2139
rect 874 2134 880 2135
rect 1022 2139 1028 2140
rect 1022 2135 1023 2139
rect 1027 2135 1028 2139
rect 1022 2134 1028 2135
rect 1250 2139 1256 2140
rect 1250 2135 1251 2139
rect 1255 2135 1256 2139
rect 1250 2134 1256 2135
rect 1442 2139 1448 2140
rect 1442 2135 1443 2139
rect 1447 2135 1448 2139
rect 1442 2134 1448 2135
rect 1634 2139 1640 2140
rect 1634 2135 1635 2139
rect 1639 2135 1640 2139
rect 1634 2134 1640 2135
rect 302 2128 308 2129
rect 302 2124 303 2128
rect 307 2124 308 2128
rect 302 2123 308 2124
rect 454 2128 460 2129
rect 454 2124 455 2128
rect 459 2124 460 2128
rect 454 2123 460 2124
rect 630 2128 636 2129
rect 630 2124 631 2128
rect 635 2124 636 2128
rect 630 2123 636 2124
rect 814 2128 820 2129
rect 814 2124 815 2128
rect 819 2124 820 2128
rect 814 2123 820 2124
rect 304 2103 306 2123
rect 456 2103 458 2123
rect 632 2103 634 2123
rect 816 2103 818 2123
rect 303 2102 307 2103
rect 303 2097 307 2098
rect 359 2102 363 2103
rect 359 2097 363 2098
rect 455 2102 459 2103
rect 455 2097 459 2098
rect 519 2102 523 2103
rect 519 2097 523 2098
rect 631 2102 635 2103
rect 631 2097 635 2098
rect 703 2102 707 2103
rect 703 2097 707 2098
rect 815 2102 819 2103
rect 815 2097 819 2098
rect 360 2081 362 2097
rect 520 2081 522 2097
rect 704 2081 706 2097
rect 358 2080 364 2081
rect 358 2076 359 2080
rect 363 2076 364 2080
rect 358 2075 364 2076
rect 518 2080 524 2081
rect 518 2076 519 2080
rect 523 2076 524 2080
rect 518 2075 524 2076
rect 702 2080 708 2081
rect 702 2076 703 2080
rect 707 2076 708 2080
rect 702 2075 708 2076
rect 282 2071 288 2072
rect 282 2067 283 2071
rect 287 2067 288 2071
rect 282 2066 288 2067
rect 290 2071 296 2072
rect 290 2067 291 2071
rect 295 2067 296 2071
rect 290 2066 296 2067
rect 586 2071 592 2072
rect 586 2067 587 2071
rect 591 2067 592 2071
rect 586 2066 592 2067
rect 770 2071 776 2072
rect 770 2067 771 2071
rect 775 2067 776 2071
rect 770 2066 776 2067
rect 110 2060 116 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 112 2027 114 2055
rect 222 2042 228 2043
rect 222 2038 223 2042
rect 227 2038 228 2042
rect 222 2037 228 2038
rect 224 2027 226 2037
rect 292 2032 294 2066
rect 366 2042 372 2043
rect 366 2038 367 2042
rect 371 2038 372 2042
rect 366 2037 372 2038
rect 526 2042 532 2043
rect 526 2038 527 2042
rect 531 2038 532 2042
rect 526 2037 532 2038
rect 290 2031 296 2032
rect 290 2027 291 2031
rect 295 2027 296 2031
rect 368 2027 370 2037
rect 390 2031 396 2032
rect 390 2027 391 2031
rect 395 2027 396 2031
rect 528 2027 530 2037
rect 588 2032 590 2066
rect 710 2042 716 2043
rect 710 2038 711 2042
rect 715 2038 716 2042
rect 710 2037 716 2038
rect 586 2031 592 2032
rect 586 2027 587 2031
rect 591 2027 592 2031
rect 712 2027 714 2037
rect 772 2032 774 2066
rect 876 2032 878 2134
rect 1830 2131 1836 2132
rect 1006 2128 1012 2129
rect 1006 2124 1007 2128
rect 1011 2124 1012 2128
rect 1006 2123 1012 2124
rect 1190 2128 1196 2129
rect 1190 2124 1191 2128
rect 1195 2124 1196 2128
rect 1190 2123 1196 2124
rect 1382 2128 1388 2129
rect 1382 2124 1383 2128
rect 1387 2124 1388 2128
rect 1382 2123 1388 2124
rect 1574 2128 1580 2129
rect 1574 2124 1575 2128
rect 1579 2124 1580 2128
rect 1574 2123 1580 2124
rect 1742 2128 1748 2129
rect 1742 2124 1743 2128
rect 1747 2124 1748 2128
rect 1830 2127 1831 2131
rect 1835 2127 1836 2131
rect 1830 2126 1836 2127
rect 1742 2123 1748 2124
rect 1008 2103 1010 2123
rect 1192 2103 1194 2123
rect 1384 2103 1386 2123
rect 1576 2103 1578 2123
rect 1744 2103 1746 2123
rect 1758 2111 1764 2112
rect 1758 2107 1759 2111
rect 1763 2107 1764 2111
rect 1758 2106 1764 2107
rect 895 2102 899 2103
rect 895 2097 899 2098
rect 1007 2102 1011 2103
rect 1007 2097 1011 2098
rect 1103 2102 1107 2103
rect 1103 2097 1107 2098
rect 1191 2102 1195 2103
rect 1191 2097 1195 2098
rect 1311 2102 1315 2103
rect 1311 2097 1315 2098
rect 1383 2102 1387 2103
rect 1383 2097 1387 2098
rect 1527 2102 1531 2103
rect 1527 2097 1531 2098
rect 1575 2102 1579 2103
rect 1575 2097 1579 2098
rect 1743 2102 1747 2103
rect 1743 2097 1747 2098
rect 896 2081 898 2097
rect 1104 2081 1106 2097
rect 1312 2081 1314 2097
rect 1528 2081 1530 2097
rect 1744 2081 1746 2097
rect 894 2080 900 2081
rect 894 2076 895 2080
rect 899 2076 900 2080
rect 894 2075 900 2076
rect 1102 2080 1108 2081
rect 1102 2076 1103 2080
rect 1107 2076 1108 2080
rect 1102 2075 1108 2076
rect 1310 2080 1316 2081
rect 1310 2076 1311 2080
rect 1315 2076 1316 2080
rect 1310 2075 1316 2076
rect 1526 2080 1532 2081
rect 1526 2076 1527 2080
rect 1531 2076 1532 2080
rect 1526 2075 1532 2076
rect 1742 2080 1748 2081
rect 1742 2076 1743 2080
rect 1747 2076 1748 2080
rect 1742 2075 1748 2076
rect 1214 2071 1220 2072
rect 1214 2067 1215 2071
rect 1219 2067 1220 2071
rect 1214 2066 1220 2067
rect 1594 2071 1600 2072
rect 1594 2067 1595 2071
rect 1599 2067 1600 2071
rect 1594 2066 1600 2067
rect 1602 2071 1608 2072
rect 1602 2067 1603 2071
rect 1607 2067 1608 2071
rect 1602 2066 1608 2067
rect 902 2042 908 2043
rect 902 2038 903 2042
rect 907 2038 908 2042
rect 902 2037 908 2038
rect 1110 2042 1116 2043
rect 1110 2038 1111 2042
rect 1115 2038 1116 2042
rect 1110 2037 1116 2038
rect 770 2031 776 2032
rect 770 2027 771 2031
rect 775 2027 776 2031
rect 874 2031 880 2032
rect 874 2027 875 2031
rect 879 2027 880 2031
rect 904 2027 906 2037
rect 1074 2031 1080 2032
rect 1074 2027 1075 2031
rect 1079 2027 1080 2031
rect 1112 2027 1114 2037
rect 1216 2032 1218 2066
rect 1318 2042 1324 2043
rect 1318 2038 1319 2042
rect 1323 2038 1324 2042
rect 1318 2037 1324 2038
rect 1534 2042 1540 2043
rect 1534 2038 1535 2042
rect 1539 2038 1540 2042
rect 1534 2037 1540 2038
rect 1214 2031 1220 2032
rect 1214 2027 1215 2031
rect 1219 2027 1220 2031
rect 1320 2027 1322 2037
rect 1536 2027 1538 2037
rect 111 2026 115 2027
rect 111 2021 115 2022
rect 143 2026 147 2027
rect 143 2021 147 2022
rect 223 2026 227 2027
rect 223 2021 227 2022
rect 263 2026 267 2027
rect 290 2026 296 2027
rect 367 2026 371 2027
rect 263 2021 267 2022
rect 367 2021 371 2022
rect 383 2026 387 2027
rect 390 2026 396 2027
rect 495 2026 499 2027
rect 383 2021 387 2022
rect 112 1993 114 2021
rect 144 2011 146 2021
rect 150 2019 156 2020
rect 150 2015 151 2019
rect 155 2015 156 2019
rect 150 2014 156 2015
rect 194 2019 200 2020
rect 194 2015 195 2019
rect 199 2015 200 2019
rect 194 2014 200 2015
rect 142 2010 148 2011
rect 142 2006 143 2010
rect 147 2006 148 2010
rect 142 2005 148 2006
rect 110 1992 116 1993
rect 110 1988 111 1992
rect 115 1988 116 1992
rect 110 1987 116 1988
rect 110 1975 116 1976
rect 110 1971 111 1975
rect 115 1971 116 1975
rect 110 1970 116 1971
rect 134 1972 140 1973
rect 112 1943 114 1970
rect 134 1968 135 1972
rect 139 1968 140 1972
rect 134 1967 140 1968
rect 136 1943 138 1967
rect 111 1942 115 1943
rect 111 1937 115 1938
rect 135 1942 139 1943
rect 135 1937 139 1938
rect 112 1918 114 1937
rect 110 1917 116 1918
rect 110 1913 111 1917
rect 115 1913 116 1917
rect 110 1912 116 1913
rect 152 1912 154 2014
rect 196 1984 198 2014
rect 264 2011 266 2021
rect 314 2019 320 2020
rect 314 2015 315 2019
rect 319 2015 320 2019
rect 314 2014 320 2015
rect 262 2010 268 2011
rect 262 2006 263 2010
rect 267 2006 268 2010
rect 262 2005 268 2006
rect 316 1984 318 2014
rect 384 2011 386 2021
rect 382 2010 388 2011
rect 382 2006 383 2010
rect 387 2006 388 2010
rect 382 2005 388 2006
rect 392 1984 394 2026
rect 495 2021 499 2022
rect 527 2026 531 2027
rect 586 2026 592 2027
rect 607 2026 611 2027
rect 527 2021 531 2022
rect 607 2021 611 2022
rect 711 2026 715 2027
rect 711 2021 715 2022
rect 719 2026 723 2027
rect 770 2026 776 2027
rect 823 2026 827 2027
rect 874 2026 880 2027
rect 903 2026 907 2027
rect 719 2021 723 2022
rect 823 2021 827 2022
rect 903 2021 907 2022
rect 927 2026 931 2027
rect 927 2021 931 2022
rect 1023 2026 1027 2027
rect 1074 2026 1080 2027
rect 1111 2026 1115 2027
rect 1023 2021 1027 2022
rect 496 2011 498 2021
rect 546 2019 552 2020
rect 546 2015 547 2019
rect 551 2015 552 2019
rect 546 2014 552 2015
rect 494 2010 500 2011
rect 494 2006 495 2010
rect 499 2006 500 2010
rect 494 2005 500 2006
rect 548 1984 550 2014
rect 608 2011 610 2021
rect 658 2019 664 2020
rect 658 2015 659 2019
rect 663 2015 664 2019
rect 658 2014 664 2015
rect 606 2010 612 2011
rect 606 2006 607 2010
rect 611 2006 612 2010
rect 606 2005 612 2006
rect 660 1984 662 2014
rect 720 2011 722 2021
rect 824 2011 826 2021
rect 866 2019 872 2020
rect 866 2015 867 2019
rect 871 2015 872 2019
rect 866 2014 872 2015
rect 874 2019 880 2020
rect 874 2015 875 2019
rect 879 2015 880 2019
rect 874 2014 880 2015
rect 718 2010 724 2011
rect 718 2006 719 2010
rect 723 2006 724 2010
rect 718 2005 724 2006
rect 822 2010 828 2011
rect 822 2006 823 2010
rect 827 2006 828 2010
rect 822 2005 828 2006
rect 194 1983 200 1984
rect 194 1979 195 1983
rect 199 1979 200 1983
rect 194 1978 200 1979
rect 314 1983 320 1984
rect 314 1979 315 1983
rect 319 1979 320 1983
rect 314 1978 320 1979
rect 390 1983 396 1984
rect 390 1979 391 1983
rect 395 1979 396 1983
rect 390 1978 396 1979
rect 546 1983 552 1984
rect 546 1979 547 1983
rect 551 1979 552 1983
rect 546 1978 552 1979
rect 658 1983 664 1984
rect 658 1979 659 1983
rect 663 1979 664 1983
rect 658 1978 664 1979
rect 770 1983 776 1984
rect 770 1979 771 1983
rect 775 1979 776 1983
rect 770 1978 776 1979
rect 254 1972 260 1973
rect 254 1968 255 1972
rect 259 1968 260 1972
rect 254 1967 260 1968
rect 374 1972 380 1973
rect 374 1968 375 1972
rect 379 1968 380 1972
rect 374 1967 380 1968
rect 486 1972 492 1973
rect 486 1968 487 1972
rect 491 1968 492 1972
rect 486 1967 492 1968
rect 598 1972 604 1973
rect 598 1968 599 1972
rect 603 1968 604 1972
rect 598 1967 604 1968
rect 710 1972 716 1973
rect 710 1968 711 1972
rect 715 1968 716 1972
rect 710 1967 716 1968
rect 256 1943 258 1967
rect 376 1943 378 1967
rect 488 1943 490 1967
rect 600 1943 602 1967
rect 712 1943 714 1967
rect 167 1942 171 1943
rect 167 1937 171 1938
rect 255 1942 259 1943
rect 255 1937 259 1938
rect 327 1942 331 1943
rect 327 1937 331 1938
rect 375 1942 379 1943
rect 375 1937 379 1938
rect 487 1942 491 1943
rect 487 1937 491 1938
rect 599 1942 603 1943
rect 599 1937 603 1938
rect 647 1942 651 1943
rect 647 1937 651 1938
rect 711 1942 715 1943
rect 711 1937 715 1938
rect 168 1921 170 1937
rect 328 1921 330 1937
rect 488 1921 490 1937
rect 648 1921 650 1937
rect 166 1920 172 1921
rect 166 1916 167 1920
rect 171 1916 172 1920
rect 166 1915 172 1916
rect 326 1920 332 1921
rect 326 1916 327 1920
rect 331 1916 332 1920
rect 326 1915 332 1916
rect 486 1920 492 1921
rect 486 1916 487 1920
rect 491 1916 492 1920
rect 486 1915 492 1916
rect 646 1920 652 1921
rect 646 1916 647 1920
rect 651 1916 652 1920
rect 646 1915 652 1916
rect 150 1911 156 1912
rect 150 1907 151 1911
rect 155 1907 156 1911
rect 150 1906 156 1907
rect 234 1911 240 1912
rect 234 1907 235 1911
rect 239 1907 240 1911
rect 234 1906 240 1907
rect 554 1911 560 1912
rect 554 1907 555 1911
rect 559 1907 560 1911
rect 554 1906 560 1907
rect 562 1911 568 1912
rect 562 1907 563 1911
rect 567 1907 568 1911
rect 562 1906 568 1907
rect 714 1911 720 1912
rect 714 1907 715 1911
rect 719 1907 720 1911
rect 714 1906 720 1907
rect 110 1900 116 1901
rect 110 1896 111 1900
rect 115 1896 116 1900
rect 110 1895 116 1896
rect 112 1867 114 1895
rect 174 1882 180 1883
rect 174 1878 175 1882
rect 179 1878 180 1882
rect 174 1877 180 1878
rect 176 1867 178 1877
rect 236 1872 238 1906
rect 334 1882 340 1883
rect 334 1878 335 1882
rect 339 1878 340 1882
rect 334 1877 340 1878
rect 494 1882 500 1883
rect 494 1878 495 1882
rect 499 1878 500 1882
rect 494 1877 500 1878
rect 234 1871 240 1872
rect 234 1867 235 1871
rect 239 1867 240 1871
rect 326 1871 332 1872
rect 326 1867 327 1871
rect 331 1867 332 1871
rect 336 1867 338 1877
rect 496 1867 498 1877
rect 111 1866 115 1867
rect 111 1861 115 1862
rect 159 1866 163 1867
rect 159 1861 163 1862
rect 175 1866 179 1867
rect 234 1866 240 1867
rect 303 1866 307 1867
rect 326 1866 332 1867
rect 335 1866 339 1867
rect 175 1861 179 1862
rect 303 1861 307 1862
rect 112 1833 114 1861
rect 160 1851 162 1861
rect 182 1859 188 1860
rect 182 1855 183 1859
rect 187 1855 188 1859
rect 182 1854 188 1855
rect 210 1859 216 1860
rect 210 1855 211 1859
rect 215 1855 216 1859
rect 210 1854 216 1855
rect 158 1850 164 1851
rect 158 1846 159 1850
rect 163 1846 164 1850
rect 158 1845 164 1846
rect 184 1845 186 1854
rect 183 1844 187 1845
rect 183 1839 187 1840
rect 110 1832 116 1833
rect 110 1828 111 1832
rect 115 1828 116 1832
rect 110 1827 116 1828
rect 212 1824 214 1854
rect 304 1851 306 1861
rect 302 1850 308 1851
rect 302 1846 303 1850
rect 307 1846 308 1850
rect 302 1845 308 1846
rect 328 1824 330 1866
rect 335 1861 339 1862
rect 447 1866 451 1867
rect 447 1861 451 1862
rect 495 1866 499 1867
rect 495 1861 499 1862
rect 430 1859 436 1860
rect 430 1855 431 1859
rect 435 1855 436 1859
rect 430 1854 436 1855
rect 210 1823 216 1824
rect 210 1819 211 1823
rect 215 1819 216 1823
rect 210 1818 216 1819
rect 326 1823 332 1824
rect 326 1819 327 1823
rect 331 1819 332 1823
rect 326 1818 332 1819
rect 110 1815 116 1816
rect 110 1811 111 1815
rect 115 1811 116 1815
rect 110 1810 116 1811
rect 150 1812 156 1813
rect 112 1787 114 1810
rect 150 1808 151 1812
rect 155 1808 156 1812
rect 150 1807 156 1808
rect 294 1812 300 1813
rect 294 1808 295 1812
rect 299 1808 300 1812
rect 294 1807 300 1808
rect 152 1787 154 1807
rect 296 1787 298 1807
rect 111 1786 115 1787
rect 111 1781 115 1782
rect 151 1786 155 1787
rect 151 1781 155 1782
rect 247 1786 251 1787
rect 247 1781 251 1782
rect 295 1786 299 1787
rect 295 1781 299 1782
rect 423 1786 427 1787
rect 423 1781 427 1782
rect 112 1762 114 1781
rect 248 1765 250 1781
rect 424 1765 426 1781
rect 246 1764 252 1765
rect 110 1761 116 1762
rect 110 1757 111 1761
rect 115 1757 116 1761
rect 246 1760 247 1764
rect 251 1760 252 1764
rect 246 1759 252 1760
rect 422 1764 428 1765
rect 422 1760 423 1764
rect 427 1760 428 1764
rect 422 1759 428 1760
rect 110 1756 116 1757
rect 342 1755 348 1756
rect 342 1751 343 1755
rect 347 1751 348 1755
rect 432 1752 434 1854
rect 448 1851 450 1861
rect 556 1860 558 1906
rect 564 1872 566 1906
rect 654 1882 660 1883
rect 654 1878 655 1882
rect 659 1878 660 1882
rect 654 1877 660 1878
rect 562 1871 568 1872
rect 562 1867 563 1871
rect 567 1867 568 1871
rect 656 1867 658 1877
rect 716 1872 718 1906
rect 772 1872 774 1978
rect 814 1972 820 1973
rect 814 1968 815 1972
rect 819 1968 820 1972
rect 814 1967 820 1968
rect 816 1943 818 1967
rect 799 1942 803 1943
rect 799 1937 803 1938
rect 815 1942 819 1943
rect 815 1937 819 1938
rect 800 1921 802 1937
rect 798 1920 804 1921
rect 798 1916 799 1920
rect 803 1916 804 1920
rect 798 1915 804 1916
rect 868 1912 870 2014
rect 876 1984 878 2014
rect 928 2011 930 2021
rect 978 2019 984 2020
rect 978 2015 979 2019
rect 983 2015 984 2019
rect 978 2014 984 2015
rect 926 2010 932 2011
rect 926 2006 927 2010
rect 931 2006 932 2010
rect 926 2005 932 2006
rect 980 1984 982 2014
rect 1024 2011 1026 2021
rect 1022 2010 1028 2011
rect 1022 2006 1023 2010
rect 1027 2006 1028 2010
rect 1022 2005 1028 2006
rect 1076 1984 1078 2026
rect 1111 2021 1115 2022
rect 1207 2026 1211 2027
rect 1214 2026 1220 2027
rect 1295 2026 1299 2027
rect 1207 2021 1211 2022
rect 1295 2021 1299 2022
rect 1319 2026 1323 2027
rect 1319 2021 1323 2022
rect 1391 2026 1395 2027
rect 1391 2021 1395 2022
rect 1487 2026 1491 2027
rect 1487 2021 1491 2022
rect 1535 2026 1539 2027
rect 1535 2021 1539 2022
rect 1583 2026 1587 2027
rect 1583 2021 1587 2022
rect 1112 2011 1114 2021
rect 1162 2019 1168 2020
rect 1162 2015 1163 2019
rect 1167 2015 1168 2019
rect 1162 2014 1168 2015
rect 1110 2010 1116 2011
rect 1110 2006 1111 2010
rect 1115 2006 1116 2010
rect 1110 2005 1116 2006
rect 1164 1984 1166 2014
rect 1208 2011 1210 2021
rect 1258 2019 1264 2020
rect 1258 2015 1259 2019
rect 1263 2015 1264 2019
rect 1258 2014 1264 2015
rect 1206 2010 1212 2011
rect 1206 2006 1207 2010
rect 1211 2006 1212 2010
rect 1206 2005 1212 2006
rect 1260 1984 1262 2014
rect 1296 2011 1298 2021
rect 1346 2019 1352 2020
rect 1346 2015 1347 2019
rect 1351 2015 1352 2019
rect 1346 2014 1352 2015
rect 1294 2010 1300 2011
rect 1294 2006 1295 2010
rect 1299 2006 1300 2010
rect 1294 2005 1300 2006
rect 1348 1984 1350 2014
rect 1392 2011 1394 2021
rect 1442 2019 1448 2020
rect 1442 2015 1443 2019
rect 1447 2015 1448 2019
rect 1442 2014 1448 2015
rect 1390 2010 1396 2011
rect 1390 2006 1391 2010
rect 1395 2006 1396 2010
rect 1390 2005 1396 2006
rect 1444 1984 1446 2014
rect 1488 2011 1490 2021
rect 1584 2011 1586 2021
rect 1596 2020 1598 2066
rect 1604 2032 1606 2066
rect 1750 2042 1756 2043
rect 1750 2038 1751 2042
rect 1755 2038 1756 2042
rect 1750 2037 1756 2038
rect 1602 2031 1608 2032
rect 1602 2027 1603 2031
rect 1607 2027 1608 2031
rect 1752 2027 1754 2037
rect 1760 2032 1762 2106
rect 1832 2103 1834 2126
rect 1872 2107 1874 2147
rect 2206 2134 2212 2135
rect 2206 2130 2207 2134
rect 2211 2130 2212 2134
rect 2206 2129 2212 2130
rect 2215 2132 2219 2133
rect 2208 2107 2210 2129
rect 2215 2127 2219 2128
rect 2216 2124 2218 2127
rect 2268 2124 2270 2158
rect 2302 2134 2308 2135
rect 2302 2130 2303 2134
rect 2307 2130 2308 2134
rect 2302 2129 2308 2130
rect 2214 2123 2220 2124
rect 2214 2119 2215 2123
rect 2219 2119 2220 2123
rect 2214 2118 2220 2119
rect 2266 2123 2272 2124
rect 2266 2119 2267 2123
rect 2271 2119 2272 2123
rect 2266 2118 2272 2119
rect 2304 2107 2306 2129
rect 2364 2124 2366 2158
rect 2406 2134 2412 2135
rect 2406 2130 2407 2134
rect 2411 2130 2412 2134
rect 2488 2133 2490 2158
rect 2526 2134 2532 2135
rect 2406 2129 2412 2130
rect 2487 2132 2491 2133
rect 2362 2123 2368 2124
rect 2362 2119 2363 2123
rect 2367 2119 2368 2123
rect 2362 2118 2368 2119
rect 2408 2107 2410 2129
rect 2526 2130 2527 2134
rect 2531 2130 2532 2134
rect 2526 2129 2532 2130
rect 2487 2127 2491 2128
rect 2454 2107 2460 2108
rect 2528 2107 2530 2129
rect 2588 2124 2590 2158
rect 2646 2134 2652 2135
rect 2646 2130 2647 2134
rect 2651 2130 2652 2134
rect 2646 2129 2652 2130
rect 2586 2123 2592 2124
rect 2586 2119 2587 2123
rect 2591 2119 2592 2123
rect 2586 2118 2592 2119
rect 2648 2107 2650 2129
rect 2708 2124 2710 2158
rect 2766 2134 2772 2135
rect 2766 2130 2767 2134
rect 2771 2130 2772 2134
rect 2766 2129 2772 2130
rect 2886 2134 2892 2135
rect 2886 2130 2887 2134
rect 2891 2130 2892 2134
rect 2886 2129 2892 2130
rect 2706 2123 2712 2124
rect 2706 2119 2707 2123
rect 2711 2119 2712 2123
rect 2706 2118 2712 2119
rect 2758 2123 2764 2124
rect 2758 2119 2759 2123
rect 2763 2119 2764 2123
rect 2758 2118 2764 2119
rect 1871 2106 1875 2107
rect 1831 2102 1835 2103
rect 1871 2101 1875 2102
rect 2175 2106 2179 2107
rect 2175 2101 2179 2102
rect 2207 2106 2211 2107
rect 2207 2101 2211 2102
rect 2271 2106 2275 2107
rect 2271 2101 2275 2102
rect 2303 2106 2307 2107
rect 2303 2101 2307 2102
rect 2375 2106 2379 2107
rect 2375 2101 2379 2102
rect 2407 2106 2411 2107
rect 2454 2103 2455 2107
rect 2459 2103 2460 2107
rect 2454 2102 2460 2103
rect 2487 2106 2491 2107
rect 2407 2101 2411 2102
rect 1831 2097 1835 2098
rect 1832 2078 1834 2097
rect 1830 2077 1836 2078
rect 1830 2073 1831 2077
rect 1835 2073 1836 2077
rect 1872 2073 1874 2101
rect 2176 2091 2178 2101
rect 2226 2099 2232 2100
rect 2226 2095 2227 2099
rect 2231 2095 2232 2099
rect 2226 2094 2232 2095
rect 2174 2090 2180 2091
rect 2174 2086 2175 2090
rect 2179 2086 2180 2090
rect 2174 2085 2180 2086
rect 1830 2072 1836 2073
rect 1870 2072 1876 2073
rect 1870 2068 1871 2072
rect 1875 2068 1876 2072
rect 1870 2067 1876 2068
rect 2228 2064 2230 2094
rect 2272 2091 2274 2101
rect 2322 2099 2328 2100
rect 2322 2095 2323 2099
rect 2327 2095 2328 2099
rect 2322 2094 2328 2095
rect 2270 2090 2276 2091
rect 2270 2086 2271 2090
rect 2275 2086 2276 2090
rect 2270 2085 2276 2086
rect 2324 2064 2326 2094
rect 2376 2091 2378 2101
rect 2426 2099 2432 2100
rect 2426 2095 2427 2099
rect 2431 2095 2432 2099
rect 2426 2094 2432 2095
rect 2374 2090 2380 2091
rect 2374 2086 2375 2090
rect 2379 2086 2380 2090
rect 2374 2085 2380 2086
rect 2428 2064 2430 2094
rect 2226 2063 2232 2064
rect 1830 2060 1836 2061
rect 1830 2056 1831 2060
rect 1835 2056 1836 2060
rect 2226 2059 2227 2063
rect 2231 2059 2232 2063
rect 2226 2058 2232 2059
rect 2322 2063 2328 2064
rect 2322 2059 2323 2063
rect 2327 2059 2328 2063
rect 2322 2058 2328 2059
rect 2426 2063 2432 2064
rect 2426 2059 2427 2063
rect 2431 2059 2432 2063
rect 2426 2058 2432 2059
rect 1830 2055 1836 2056
rect 1870 2055 1876 2056
rect 1758 2031 1764 2032
rect 1758 2027 1759 2031
rect 1763 2027 1764 2031
rect 1832 2027 1834 2055
rect 1870 2051 1871 2055
rect 1875 2051 1876 2055
rect 1870 2050 1876 2051
rect 2166 2052 2172 2053
rect 1872 2027 1874 2050
rect 2166 2048 2167 2052
rect 2171 2048 2172 2052
rect 2166 2047 2172 2048
rect 2262 2052 2268 2053
rect 2262 2048 2263 2052
rect 2267 2048 2268 2052
rect 2262 2047 2268 2048
rect 2366 2052 2372 2053
rect 2366 2048 2367 2052
rect 2371 2048 2372 2052
rect 2366 2047 2372 2048
rect 2168 2027 2170 2047
rect 2264 2027 2266 2047
rect 2368 2027 2370 2047
rect 1602 2026 1608 2027
rect 1671 2026 1675 2027
rect 1671 2021 1675 2022
rect 1751 2026 1755 2027
rect 1758 2026 1764 2027
rect 1831 2026 1835 2027
rect 1751 2021 1755 2022
rect 1831 2021 1835 2022
rect 1871 2026 1875 2027
rect 1871 2021 1875 2022
rect 2071 2026 2075 2027
rect 2071 2021 2075 2022
rect 2167 2026 2171 2027
rect 2167 2021 2171 2022
rect 2207 2026 2211 2027
rect 2207 2021 2211 2022
rect 2263 2026 2267 2027
rect 2263 2021 2267 2022
rect 2359 2026 2363 2027
rect 2359 2021 2363 2022
rect 2367 2026 2371 2027
rect 2367 2021 2371 2022
rect 1594 2019 1600 2020
rect 1594 2015 1595 2019
rect 1599 2015 1600 2019
rect 1594 2014 1600 2015
rect 1634 2019 1640 2020
rect 1634 2015 1635 2019
rect 1639 2015 1640 2019
rect 1634 2014 1640 2015
rect 1486 2010 1492 2011
rect 1486 2006 1487 2010
rect 1491 2006 1492 2010
rect 1486 2005 1492 2006
rect 1582 2010 1588 2011
rect 1582 2006 1583 2010
rect 1587 2006 1588 2010
rect 1582 2005 1588 2006
rect 1636 1984 1638 2014
rect 1672 2011 1674 2021
rect 1722 2019 1728 2020
rect 1722 2015 1723 2019
rect 1727 2015 1728 2019
rect 1722 2014 1728 2015
rect 1670 2010 1676 2011
rect 1670 2006 1671 2010
rect 1675 2006 1676 2010
rect 1670 2005 1676 2006
rect 1724 1984 1726 2014
rect 1752 2011 1754 2021
rect 1750 2010 1756 2011
rect 1750 2006 1751 2010
rect 1755 2006 1756 2010
rect 1750 2005 1756 2006
rect 1832 1993 1834 2021
rect 1872 2002 1874 2021
rect 2072 2005 2074 2021
rect 2208 2005 2210 2021
rect 2360 2005 2362 2021
rect 2070 2004 2076 2005
rect 1870 2001 1876 2002
rect 1870 1997 1871 2001
rect 1875 1997 1876 2001
rect 2070 2000 2071 2004
rect 2075 2000 2076 2004
rect 2070 1999 2076 2000
rect 2206 2004 2212 2005
rect 2206 2000 2207 2004
rect 2211 2000 2212 2004
rect 2206 1999 2212 2000
rect 2358 2004 2364 2005
rect 2358 2000 2359 2004
rect 2363 2000 2364 2004
rect 2358 1999 2364 2000
rect 1870 1996 1876 1997
rect 2456 1996 2458 2102
rect 2487 2101 2491 2102
rect 2527 2106 2531 2107
rect 2527 2101 2531 2102
rect 2607 2106 2611 2107
rect 2607 2101 2611 2102
rect 2647 2106 2651 2107
rect 2647 2101 2651 2102
rect 2727 2106 2731 2107
rect 2727 2101 2731 2102
rect 2488 2091 2490 2101
rect 2538 2099 2544 2100
rect 2538 2095 2539 2099
rect 2543 2095 2544 2099
rect 2538 2094 2544 2095
rect 2486 2090 2492 2091
rect 2486 2086 2487 2090
rect 2491 2086 2492 2090
rect 2486 2085 2492 2086
rect 2540 2064 2542 2094
rect 2608 2091 2610 2101
rect 2658 2099 2664 2100
rect 2658 2095 2659 2099
rect 2663 2095 2664 2099
rect 2658 2094 2664 2095
rect 2606 2090 2612 2091
rect 2606 2086 2607 2090
rect 2611 2086 2612 2090
rect 2606 2085 2612 2086
rect 2660 2064 2662 2094
rect 2728 2091 2730 2101
rect 2726 2090 2732 2091
rect 2726 2086 2727 2090
rect 2731 2086 2732 2090
rect 2726 2085 2732 2086
rect 2760 2064 2762 2118
rect 2768 2107 2770 2129
rect 2888 2107 2890 2129
rect 2948 2124 2950 2158
rect 2998 2134 3004 2135
rect 2998 2130 2999 2134
rect 3003 2130 3004 2134
rect 2998 2129 3004 2130
rect 2946 2123 2952 2124
rect 2946 2119 2947 2123
rect 2951 2119 2952 2123
rect 2946 2118 2952 2119
rect 3000 2107 3002 2129
rect 3060 2124 3062 2158
rect 3102 2134 3108 2135
rect 3102 2130 3103 2134
rect 3107 2130 3108 2134
rect 3102 2129 3108 2130
rect 3058 2123 3064 2124
rect 3058 2119 3059 2123
rect 3063 2119 3064 2123
rect 3058 2118 3064 2119
rect 3104 2107 3106 2129
rect 3176 2124 3178 2158
rect 3206 2134 3212 2135
rect 3206 2130 3207 2134
rect 3211 2130 3212 2134
rect 3206 2129 3212 2130
rect 3174 2123 3180 2124
rect 3174 2119 3175 2123
rect 3179 2119 3180 2123
rect 3174 2118 3180 2119
rect 3208 2107 3210 2129
rect 3268 2124 3270 2158
rect 3310 2134 3316 2135
rect 3310 2130 3311 2134
rect 3315 2130 3316 2134
rect 3310 2129 3316 2130
rect 3266 2123 3272 2124
rect 3266 2119 3267 2123
rect 3271 2119 3272 2123
rect 3266 2118 3272 2119
rect 3312 2107 3314 2129
rect 3336 2124 3338 2242
rect 3590 2239 3596 2240
rect 3486 2236 3492 2237
rect 3486 2232 3487 2236
rect 3491 2232 3492 2236
rect 3590 2235 3591 2239
rect 3595 2235 3596 2239
rect 3590 2234 3596 2235
rect 3486 2231 3492 2232
rect 3488 2195 3490 2231
rect 3592 2195 3594 2234
rect 3407 2194 3411 2195
rect 3407 2189 3411 2190
rect 3487 2194 3491 2195
rect 3487 2189 3491 2190
rect 3503 2194 3507 2195
rect 3503 2189 3507 2190
rect 3591 2194 3595 2195
rect 3591 2189 3595 2190
rect 3408 2173 3410 2189
rect 3504 2173 3506 2189
rect 3406 2172 3412 2173
rect 3406 2168 3407 2172
rect 3411 2168 3412 2172
rect 3406 2167 3412 2168
rect 3502 2172 3508 2173
rect 3502 2168 3503 2172
rect 3507 2168 3508 2172
rect 3592 2170 3594 2189
rect 3502 2167 3508 2168
rect 3590 2169 3596 2170
rect 3590 2165 3591 2169
rect 3595 2165 3596 2169
rect 3590 2164 3596 2165
rect 3474 2163 3480 2164
rect 3474 2159 3475 2163
rect 3479 2159 3480 2163
rect 3474 2158 3480 2159
rect 3502 2159 3508 2160
rect 3414 2134 3420 2135
rect 3414 2130 3415 2134
rect 3419 2130 3420 2134
rect 3414 2129 3420 2130
rect 3318 2123 3324 2124
rect 3318 2119 3319 2123
rect 3323 2119 3324 2123
rect 3318 2118 3324 2119
rect 3334 2123 3340 2124
rect 3334 2119 3335 2123
rect 3339 2119 3340 2123
rect 3334 2118 3340 2119
rect 2767 2106 2771 2107
rect 2767 2101 2771 2102
rect 2847 2106 2851 2107
rect 2847 2101 2851 2102
rect 2887 2106 2891 2107
rect 2887 2101 2891 2102
rect 2967 2106 2971 2107
rect 2967 2101 2971 2102
rect 2999 2106 3003 2107
rect 2999 2101 3003 2102
rect 3079 2106 3083 2107
rect 3079 2101 3083 2102
rect 3103 2106 3107 2107
rect 3103 2101 3107 2102
rect 3191 2106 3195 2107
rect 3191 2101 3195 2102
rect 3207 2106 3211 2107
rect 3207 2101 3211 2102
rect 3303 2106 3307 2107
rect 3303 2101 3307 2102
rect 3311 2106 3315 2107
rect 3311 2101 3315 2102
rect 2848 2091 2850 2101
rect 2898 2099 2904 2100
rect 2898 2095 2899 2099
rect 2903 2095 2904 2099
rect 2898 2094 2904 2095
rect 2846 2090 2852 2091
rect 2846 2086 2847 2090
rect 2851 2086 2852 2090
rect 2846 2085 2852 2086
rect 2900 2064 2902 2094
rect 2968 2091 2970 2101
rect 3018 2099 3024 2100
rect 3018 2095 3019 2099
rect 3023 2095 3024 2099
rect 3018 2094 3024 2095
rect 2966 2090 2972 2091
rect 2966 2086 2967 2090
rect 2971 2086 2972 2090
rect 2966 2085 2972 2086
rect 3020 2064 3022 2094
rect 3080 2091 3082 2101
rect 3192 2091 3194 2101
rect 3242 2099 3248 2100
rect 3242 2095 3243 2099
rect 3247 2095 3248 2099
rect 3242 2094 3248 2095
rect 3078 2090 3084 2091
rect 3078 2086 3079 2090
rect 3083 2086 3084 2090
rect 3078 2085 3084 2086
rect 3190 2090 3196 2091
rect 3190 2086 3191 2090
rect 3195 2086 3196 2090
rect 3190 2085 3196 2086
rect 3244 2064 3246 2094
rect 3304 2091 3306 2101
rect 3302 2090 3308 2091
rect 3302 2086 3303 2090
rect 3307 2086 3308 2090
rect 3302 2085 3308 2086
rect 3320 2064 3322 2118
rect 3416 2107 3418 2129
rect 3476 2124 3478 2158
rect 3502 2155 3503 2159
rect 3507 2155 3508 2159
rect 3502 2154 3508 2155
rect 3474 2123 3480 2124
rect 3474 2119 3475 2123
rect 3479 2119 3480 2123
rect 3474 2118 3480 2119
rect 3422 2107 3428 2108
rect 3415 2106 3419 2107
rect 3422 2103 3423 2107
rect 3427 2103 3428 2107
rect 3422 2102 3428 2103
rect 3415 2101 3419 2102
rect 3416 2091 3418 2101
rect 3414 2090 3420 2091
rect 3414 2086 3415 2090
rect 3419 2086 3420 2090
rect 3414 2085 3420 2086
rect 3424 2064 3426 2102
rect 3504 2100 3506 2154
rect 3590 2152 3596 2153
rect 3590 2148 3591 2152
rect 3595 2148 3596 2152
rect 3590 2147 3596 2148
rect 3510 2134 3516 2135
rect 3510 2130 3511 2134
rect 3515 2130 3516 2134
rect 3510 2129 3516 2130
rect 3512 2107 3514 2129
rect 3592 2107 3594 2147
rect 3511 2106 3515 2107
rect 3511 2101 3515 2102
rect 3591 2106 3595 2107
rect 3591 2101 3595 2102
rect 3430 2099 3436 2100
rect 3430 2095 3431 2099
rect 3435 2095 3436 2099
rect 3430 2094 3436 2095
rect 3502 2099 3508 2100
rect 3502 2095 3503 2099
rect 3507 2095 3508 2099
rect 3502 2094 3508 2095
rect 2538 2063 2544 2064
rect 2538 2059 2539 2063
rect 2543 2059 2544 2063
rect 2538 2058 2544 2059
rect 2658 2063 2664 2064
rect 2658 2059 2659 2063
rect 2663 2059 2664 2063
rect 2658 2058 2664 2059
rect 2758 2063 2764 2064
rect 2758 2059 2759 2063
rect 2763 2059 2764 2063
rect 2758 2058 2764 2059
rect 2898 2063 2904 2064
rect 2898 2059 2899 2063
rect 2903 2059 2904 2063
rect 2898 2058 2904 2059
rect 3018 2063 3024 2064
rect 3018 2059 3019 2063
rect 3023 2059 3024 2063
rect 3018 2058 3024 2059
rect 3242 2063 3248 2064
rect 3242 2059 3243 2063
rect 3247 2059 3248 2063
rect 3242 2058 3248 2059
rect 3318 2063 3324 2064
rect 3318 2059 3319 2063
rect 3323 2059 3324 2063
rect 3318 2058 3324 2059
rect 3422 2063 3428 2064
rect 3422 2059 3423 2063
rect 3427 2059 3428 2063
rect 3422 2058 3428 2059
rect 2478 2052 2484 2053
rect 2478 2048 2479 2052
rect 2483 2048 2484 2052
rect 2478 2047 2484 2048
rect 2598 2052 2604 2053
rect 2598 2048 2599 2052
rect 2603 2048 2604 2052
rect 2598 2047 2604 2048
rect 2718 2052 2724 2053
rect 2718 2048 2719 2052
rect 2723 2048 2724 2052
rect 2718 2047 2724 2048
rect 2838 2052 2844 2053
rect 2838 2048 2839 2052
rect 2843 2048 2844 2052
rect 2838 2047 2844 2048
rect 2958 2052 2964 2053
rect 2958 2048 2959 2052
rect 2963 2048 2964 2052
rect 2958 2047 2964 2048
rect 3070 2052 3076 2053
rect 3070 2048 3071 2052
rect 3075 2048 3076 2052
rect 3070 2047 3076 2048
rect 3182 2052 3188 2053
rect 3182 2048 3183 2052
rect 3187 2048 3188 2052
rect 3182 2047 3188 2048
rect 3294 2052 3300 2053
rect 3294 2048 3295 2052
rect 3299 2048 3300 2052
rect 3294 2047 3300 2048
rect 3406 2052 3412 2053
rect 3406 2048 3407 2052
rect 3411 2048 3412 2052
rect 3406 2047 3412 2048
rect 2480 2027 2482 2047
rect 2600 2027 2602 2047
rect 2720 2027 2722 2047
rect 2840 2027 2842 2047
rect 2960 2027 2962 2047
rect 3030 2035 3036 2036
rect 3030 2031 3031 2035
rect 3035 2031 3036 2035
rect 3030 2030 3036 2031
rect 2479 2026 2483 2027
rect 2479 2021 2483 2022
rect 2519 2026 2523 2027
rect 2519 2021 2523 2022
rect 2599 2026 2603 2027
rect 2599 2021 2603 2022
rect 2679 2026 2683 2027
rect 2679 2021 2683 2022
rect 2719 2026 2723 2027
rect 2719 2021 2723 2022
rect 2839 2026 2843 2027
rect 2839 2021 2843 2022
rect 2847 2026 2851 2027
rect 2847 2021 2851 2022
rect 2959 2026 2963 2027
rect 2959 2021 2963 2022
rect 3015 2026 3019 2027
rect 3015 2021 3019 2022
rect 2520 2005 2522 2021
rect 2680 2005 2682 2021
rect 2848 2005 2850 2021
rect 3016 2005 3018 2021
rect 2518 2004 2524 2005
rect 2518 2000 2519 2004
rect 2523 2000 2524 2004
rect 2518 1999 2524 2000
rect 2678 2004 2684 2005
rect 2678 2000 2679 2004
rect 2683 2000 2684 2004
rect 2678 1999 2684 2000
rect 2846 2004 2852 2005
rect 2846 2000 2847 2004
rect 2851 2000 2852 2004
rect 2846 1999 2852 2000
rect 3014 2004 3020 2005
rect 3014 2000 3015 2004
rect 3019 2000 3020 2004
rect 3014 1999 3020 2000
rect 2146 1995 2152 1996
rect 1830 1992 1836 1993
rect 1830 1988 1831 1992
rect 1835 1988 1836 1992
rect 2146 1991 2147 1995
rect 2151 1991 2152 1995
rect 2146 1990 2152 1991
rect 2274 1995 2280 1996
rect 2274 1991 2275 1995
rect 2279 1991 2280 1995
rect 2274 1990 2280 1991
rect 2446 1995 2452 1996
rect 2446 1991 2447 1995
rect 2451 1991 2452 1995
rect 2446 1990 2452 1991
rect 2454 1995 2460 1996
rect 2454 1991 2455 1995
rect 2459 1991 2460 1995
rect 2454 1990 2460 1991
rect 2598 1995 2604 1996
rect 2598 1991 2599 1995
rect 2603 1991 2604 1995
rect 2598 1990 2604 1991
rect 2746 1995 2752 1996
rect 2746 1991 2747 1995
rect 2751 1991 2752 1995
rect 2746 1990 2752 1991
rect 2914 1995 2920 1996
rect 2914 1991 2915 1995
rect 2919 1991 2920 1995
rect 2914 1990 2920 1991
rect 1830 1987 1836 1988
rect 1870 1984 1876 1985
rect 874 1983 880 1984
rect 874 1979 875 1983
rect 879 1979 880 1983
rect 874 1978 880 1979
rect 978 1983 984 1984
rect 978 1979 979 1983
rect 983 1979 984 1983
rect 978 1978 984 1979
rect 1074 1983 1080 1984
rect 1074 1979 1075 1983
rect 1079 1979 1080 1983
rect 1074 1978 1080 1979
rect 1162 1983 1168 1984
rect 1162 1979 1163 1983
rect 1167 1979 1168 1983
rect 1162 1978 1168 1979
rect 1258 1983 1264 1984
rect 1258 1979 1259 1983
rect 1263 1979 1264 1983
rect 1258 1978 1264 1979
rect 1346 1983 1352 1984
rect 1346 1979 1347 1983
rect 1351 1979 1352 1983
rect 1346 1978 1352 1979
rect 1442 1983 1448 1984
rect 1442 1979 1443 1983
rect 1447 1979 1448 1983
rect 1442 1978 1448 1979
rect 1634 1983 1640 1984
rect 1634 1979 1635 1983
rect 1639 1979 1640 1983
rect 1634 1978 1640 1979
rect 1722 1983 1728 1984
rect 1722 1979 1723 1983
rect 1727 1979 1728 1983
rect 1870 1980 1871 1984
rect 1875 1980 1876 1984
rect 1870 1979 1876 1980
rect 1722 1978 1728 1979
rect 1830 1975 1836 1976
rect 918 1972 924 1973
rect 918 1968 919 1972
rect 923 1968 924 1972
rect 918 1967 924 1968
rect 1014 1972 1020 1973
rect 1014 1968 1015 1972
rect 1019 1968 1020 1972
rect 1014 1967 1020 1968
rect 1102 1972 1108 1973
rect 1102 1968 1103 1972
rect 1107 1968 1108 1972
rect 1102 1967 1108 1968
rect 1198 1972 1204 1973
rect 1198 1968 1199 1972
rect 1203 1968 1204 1972
rect 1198 1967 1204 1968
rect 1286 1972 1292 1973
rect 1286 1968 1287 1972
rect 1291 1968 1292 1972
rect 1286 1967 1292 1968
rect 1382 1972 1388 1973
rect 1382 1968 1383 1972
rect 1387 1968 1388 1972
rect 1382 1967 1388 1968
rect 1478 1972 1484 1973
rect 1478 1968 1479 1972
rect 1483 1968 1484 1972
rect 1478 1967 1484 1968
rect 1574 1972 1580 1973
rect 1574 1968 1575 1972
rect 1579 1968 1580 1972
rect 1574 1967 1580 1968
rect 1662 1972 1668 1973
rect 1662 1968 1663 1972
rect 1667 1968 1668 1972
rect 1662 1967 1668 1968
rect 1742 1972 1748 1973
rect 1742 1968 1743 1972
rect 1747 1968 1748 1972
rect 1830 1971 1831 1975
rect 1835 1971 1836 1975
rect 1830 1970 1836 1971
rect 1742 1967 1748 1968
rect 920 1943 922 1967
rect 1016 1943 1018 1967
rect 1104 1943 1106 1967
rect 1200 1943 1202 1967
rect 1230 1955 1236 1956
rect 1230 1951 1231 1955
rect 1235 1951 1236 1955
rect 1230 1950 1236 1951
rect 919 1942 923 1943
rect 919 1937 923 1938
rect 943 1942 947 1943
rect 943 1937 947 1938
rect 1015 1942 1019 1943
rect 1015 1937 1019 1938
rect 1079 1942 1083 1943
rect 1079 1937 1083 1938
rect 1103 1942 1107 1943
rect 1103 1937 1107 1938
rect 1199 1942 1203 1943
rect 1199 1937 1203 1938
rect 1215 1942 1219 1943
rect 1215 1937 1219 1938
rect 944 1921 946 1937
rect 1080 1921 1082 1937
rect 1216 1921 1218 1937
rect 942 1920 948 1921
rect 942 1916 943 1920
rect 947 1916 948 1920
rect 942 1915 948 1916
rect 1078 1920 1084 1921
rect 1078 1916 1079 1920
rect 1083 1916 1084 1920
rect 1078 1915 1084 1916
rect 1214 1920 1220 1921
rect 1214 1916 1215 1920
rect 1219 1916 1220 1920
rect 1214 1915 1220 1916
rect 866 1911 872 1912
rect 866 1907 867 1911
rect 871 1907 872 1911
rect 866 1906 872 1907
rect 1010 1911 1016 1912
rect 1010 1907 1011 1911
rect 1015 1907 1016 1911
rect 1010 1906 1016 1907
rect 806 1882 812 1883
rect 806 1878 807 1882
rect 811 1878 812 1882
rect 806 1877 812 1878
rect 950 1882 956 1883
rect 950 1878 951 1882
rect 955 1878 956 1882
rect 950 1877 956 1878
rect 714 1871 720 1872
rect 714 1867 715 1871
rect 719 1867 720 1871
rect 770 1871 776 1872
rect 770 1867 771 1871
rect 775 1867 776 1871
rect 808 1867 810 1877
rect 952 1867 954 1877
rect 1012 1872 1014 1906
rect 1086 1882 1092 1883
rect 1086 1878 1087 1882
rect 1091 1878 1092 1882
rect 1086 1877 1092 1878
rect 1222 1882 1228 1883
rect 1222 1878 1223 1882
rect 1227 1878 1228 1882
rect 1222 1877 1228 1878
rect 1010 1871 1016 1872
rect 1010 1867 1011 1871
rect 1015 1867 1016 1871
rect 1078 1871 1084 1872
rect 1078 1867 1079 1871
rect 1083 1867 1084 1871
rect 1088 1867 1090 1877
rect 1224 1867 1226 1877
rect 1232 1872 1234 1950
rect 1288 1943 1290 1967
rect 1384 1943 1386 1967
rect 1480 1943 1482 1967
rect 1576 1943 1578 1967
rect 1664 1943 1666 1967
rect 1744 1943 1746 1967
rect 1758 1955 1764 1956
rect 1758 1951 1759 1955
rect 1763 1951 1764 1955
rect 1758 1950 1764 1951
rect 1287 1942 1291 1943
rect 1287 1937 1291 1938
rect 1351 1942 1355 1943
rect 1351 1937 1355 1938
rect 1383 1942 1387 1943
rect 1383 1937 1387 1938
rect 1479 1942 1483 1943
rect 1479 1937 1483 1938
rect 1487 1942 1491 1943
rect 1487 1937 1491 1938
rect 1575 1942 1579 1943
rect 1575 1937 1579 1938
rect 1623 1942 1627 1943
rect 1623 1937 1627 1938
rect 1663 1942 1667 1943
rect 1663 1937 1667 1938
rect 1743 1942 1747 1943
rect 1743 1937 1747 1938
rect 1352 1921 1354 1937
rect 1488 1921 1490 1937
rect 1624 1921 1626 1937
rect 1744 1921 1746 1937
rect 1350 1920 1356 1921
rect 1350 1916 1351 1920
rect 1355 1916 1356 1920
rect 1350 1915 1356 1916
rect 1486 1920 1492 1921
rect 1486 1916 1487 1920
rect 1491 1916 1492 1920
rect 1486 1915 1492 1916
rect 1622 1920 1628 1921
rect 1622 1916 1623 1920
rect 1627 1916 1628 1920
rect 1622 1915 1628 1916
rect 1742 1920 1748 1921
rect 1742 1916 1743 1920
rect 1747 1916 1748 1920
rect 1742 1915 1748 1916
rect 1290 1911 1296 1912
rect 1290 1907 1291 1911
rect 1295 1907 1296 1911
rect 1290 1906 1296 1907
rect 1418 1911 1424 1912
rect 1418 1907 1419 1911
rect 1423 1907 1424 1911
rect 1418 1906 1424 1907
rect 1554 1911 1560 1912
rect 1554 1907 1555 1911
rect 1559 1907 1560 1911
rect 1554 1906 1560 1907
rect 1292 1872 1294 1906
rect 1342 1903 1348 1904
rect 1342 1899 1343 1903
rect 1347 1899 1348 1903
rect 1342 1898 1348 1899
rect 1230 1871 1236 1872
rect 1230 1867 1231 1871
rect 1235 1867 1236 1871
rect 562 1866 568 1867
rect 599 1866 603 1867
rect 599 1861 603 1862
rect 655 1866 659 1867
rect 714 1866 720 1867
rect 751 1866 755 1867
rect 770 1866 776 1867
rect 807 1866 811 1867
rect 655 1861 659 1862
rect 751 1861 755 1862
rect 807 1861 811 1862
rect 903 1866 907 1867
rect 903 1861 907 1862
rect 951 1866 955 1867
rect 1010 1866 1016 1867
rect 1055 1866 1059 1867
rect 1078 1866 1084 1867
rect 1087 1866 1091 1867
rect 951 1861 955 1862
rect 1055 1861 1059 1862
rect 554 1859 560 1860
rect 554 1855 555 1859
rect 559 1855 560 1859
rect 554 1854 560 1855
rect 600 1851 602 1861
rect 752 1851 754 1861
rect 838 1859 844 1860
rect 838 1855 839 1859
rect 843 1855 844 1859
rect 838 1854 844 1855
rect 446 1850 452 1851
rect 446 1846 447 1850
rect 451 1846 452 1850
rect 446 1845 452 1846
rect 598 1850 604 1851
rect 598 1846 599 1850
rect 603 1846 604 1850
rect 598 1845 604 1846
rect 750 1850 756 1851
rect 750 1846 751 1850
rect 755 1846 756 1850
rect 750 1845 756 1846
rect 455 1844 459 1845
rect 455 1839 459 1840
rect 456 1824 458 1839
rect 840 1824 842 1854
rect 904 1851 906 1861
rect 1056 1851 1058 1861
rect 902 1850 908 1851
rect 902 1846 903 1850
rect 907 1846 908 1850
rect 902 1845 908 1846
rect 1054 1850 1060 1851
rect 1054 1846 1055 1850
rect 1059 1846 1060 1850
rect 1054 1845 1060 1846
rect 1080 1824 1082 1866
rect 1087 1861 1091 1862
rect 1207 1866 1211 1867
rect 1207 1861 1211 1862
rect 1223 1866 1227 1867
rect 1230 1866 1236 1867
rect 1290 1871 1296 1872
rect 1290 1867 1291 1871
rect 1295 1867 1296 1871
rect 1290 1866 1296 1867
rect 1223 1861 1227 1862
rect 1198 1859 1204 1860
rect 1198 1855 1199 1859
rect 1203 1855 1204 1859
rect 1198 1854 1204 1855
rect 1200 1843 1202 1854
rect 1208 1851 1210 1861
rect 1344 1860 1346 1898
rect 1358 1882 1364 1883
rect 1358 1878 1359 1882
rect 1363 1878 1364 1882
rect 1358 1877 1364 1878
rect 1360 1867 1362 1877
rect 1420 1872 1422 1906
rect 1494 1882 1500 1883
rect 1494 1878 1495 1882
rect 1499 1878 1500 1882
rect 1494 1877 1500 1878
rect 1418 1871 1424 1872
rect 1418 1867 1419 1871
rect 1423 1867 1424 1871
rect 1496 1867 1498 1877
rect 1556 1872 1558 1906
rect 1630 1882 1636 1883
rect 1630 1878 1631 1882
rect 1635 1878 1636 1882
rect 1630 1877 1636 1878
rect 1750 1882 1756 1883
rect 1750 1878 1751 1882
rect 1755 1878 1756 1882
rect 1750 1877 1756 1878
rect 1554 1871 1560 1872
rect 1554 1867 1555 1871
rect 1559 1867 1560 1871
rect 1632 1867 1634 1877
rect 1752 1867 1754 1877
rect 1760 1872 1762 1950
rect 1810 1943 1816 1944
rect 1832 1943 1834 1970
rect 1872 1951 1874 1979
rect 2078 1966 2084 1967
rect 2078 1962 2079 1966
rect 2083 1962 2084 1966
rect 2078 1961 2084 1962
rect 2058 1955 2064 1956
rect 2058 1951 2059 1955
rect 2063 1951 2064 1955
rect 2080 1951 2082 1961
rect 2148 1956 2150 1990
rect 2214 1966 2220 1967
rect 2214 1962 2215 1966
rect 2219 1962 2220 1966
rect 2214 1961 2220 1962
rect 2146 1955 2152 1956
rect 2146 1951 2147 1955
rect 2151 1951 2152 1955
rect 2216 1951 2218 1961
rect 2276 1956 2278 1990
rect 2383 1972 2387 1973
rect 2383 1967 2387 1968
rect 2366 1966 2372 1967
rect 2366 1962 2367 1966
rect 2371 1962 2372 1966
rect 2366 1961 2372 1962
rect 2274 1955 2280 1956
rect 2274 1951 2275 1955
rect 2279 1951 2280 1955
rect 2368 1951 2370 1961
rect 1871 1950 1875 1951
rect 1871 1945 1875 1946
rect 1903 1950 1907 1951
rect 1903 1945 1907 1946
rect 2007 1950 2011 1951
rect 2058 1950 2064 1951
rect 2079 1950 2083 1951
rect 2007 1945 2011 1946
rect 1810 1939 1811 1943
rect 1815 1939 1816 1943
rect 1810 1938 1816 1939
rect 1831 1942 1835 1943
rect 1812 1912 1814 1938
rect 1831 1937 1835 1938
rect 1832 1918 1834 1937
rect 1830 1917 1836 1918
rect 1872 1917 1874 1945
rect 1904 1935 1906 1945
rect 2008 1935 2010 1945
rect 1902 1934 1908 1935
rect 1902 1930 1903 1934
rect 1907 1930 1908 1934
rect 1902 1929 1908 1930
rect 2006 1934 2012 1935
rect 2006 1930 2007 1934
rect 2011 1930 2012 1934
rect 2006 1929 2012 1930
rect 1830 1913 1831 1917
rect 1835 1913 1836 1917
rect 1830 1912 1836 1913
rect 1870 1916 1876 1917
rect 1870 1912 1871 1916
rect 1875 1912 1876 1916
rect 1810 1911 1816 1912
rect 1870 1911 1876 1912
rect 1810 1907 1811 1911
rect 1815 1907 1816 1911
rect 2060 1908 2062 1950
rect 2079 1945 2083 1946
rect 2135 1950 2139 1951
rect 2146 1950 2152 1951
rect 2215 1950 2219 1951
rect 2135 1945 2139 1946
rect 2215 1945 2219 1946
rect 2255 1950 2259 1951
rect 2274 1950 2280 1951
rect 2367 1950 2371 1951
rect 2255 1945 2259 1946
rect 2367 1945 2371 1946
rect 2375 1950 2379 1951
rect 2375 1945 2379 1946
rect 2066 1943 2072 1944
rect 2066 1939 2067 1943
rect 2071 1939 2072 1943
rect 2066 1938 2072 1939
rect 2068 1908 2070 1938
rect 2136 1935 2138 1945
rect 2194 1943 2200 1944
rect 2194 1939 2195 1943
rect 2199 1939 2200 1943
rect 2194 1938 2200 1939
rect 2134 1934 2140 1935
rect 2134 1930 2135 1934
rect 2139 1930 2140 1934
rect 2134 1929 2140 1930
rect 2196 1908 2198 1938
rect 2256 1935 2258 1945
rect 2350 1943 2356 1944
rect 2350 1939 2351 1943
rect 2355 1939 2356 1943
rect 2350 1938 2356 1939
rect 2254 1934 2260 1935
rect 2254 1930 2255 1934
rect 2259 1930 2260 1934
rect 2254 1929 2260 1930
rect 1810 1906 1816 1907
rect 2058 1907 2064 1908
rect 2058 1903 2059 1907
rect 2063 1903 2064 1907
rect 2058 1902 2064 1903
rect 2066 1907 2072 1908
rect 2066 1903 2067 1907
rect 2071 1903 2072 1907
rect 2066 1902 2072 1903
rect 2194 1907 2200 1908
rect 2194 1903 2195 1907
rect 2199 1903 2200 1907
rect 2194 1902 2200 1903
rect 1830 1900 1836 1901
rect 1830 1896 1831 1900
rect 1835 1896 1836 1900
rect 1830 1895 1836 1896
rect 1870 1899 1876 1900
rect 1870 1895 1871 1899
rect 1875 1895 1876 1899
rect 1758 1871 1764 1872
rect 1758 1867 1759 1871
rect 1763 1867 1764 1871
rect 1832 1867 1834 1895
rect 1870 1894 1876 1895
rect 1894 1896 1900 1897
rect 1872 1875 1874 1894
rect 1894 1892 1895 1896
rect 1899 1892 1900 1896
rect 1894 1891 1900 1892
rect 1998 1896 2004 1897
rect 1998 1892 1999 1896
rect 2003 1892 2004 1896
rect 1998 1891 2004 1892
rect 2126 1896 2132 1897
rect 2126 1892 2127 1896
rect 2131 1892 2132 1896
rect 2126 1891 2132 1892
rect 2246 1896 2252 1897
rect 2246 1892 2247 1896
rect 2251 1892 2252 1896
rect 2246 1891 2252 1892
rect 1896 1875 1898 1891
rect 1910 1879 1916 1880
rect 1910 1875 1911 1879
rect 1915 1875 1916 1879
rect 2000 1875 2002 1891
rect 2128 1875 2130 1891
rect 2248 1875 2250 1891
rect 1871 1874 1875 1875
rect 1871 1869 1875 1870
rect 1895 1874 1899 1875
rect 1910 1874 1916 1875
rect 1991 1874 1995 1875
rect 1895 1869 1899 1870
rect 1351 1866 1355 1867
rect 1351 1861 1355 1862
rect 1359 1866 1363 1867
rect 1418 1866 1424 1867
rect 1487 1866 1491 1867
rect 1359 1861 1363 1862
rect 1487 1861 1491 1862
rect 1495 1866 1499 1867
rect 1554 1866 1560 1867
rect 1631 1866 1635 1867
rect 1495 1861 1499 1862
rect 1631 1861 1635 1862
rect 1751 1866 1755 1867
rect 1758 1866 1764 1867
rect 1831 1866 1835 1867
rect 1751 1861 1755 1862
rect 1831 1861 1835 1862
rect 1342 1859 1348 1860
rect 1342 1855 1343 1859
rect 1347 1855 1348 1859
rect 1342 1854 1348 1855
rect 1352 1851 1354 1861
rect 1402 1859 1408 1860
rect 1402 1855 1403 1859
rect 1407 1855 1408 1859
rect 1402 1854 1408 1855
rect 1206 1850 1212 1851
rect 1206 1846 1207 1850
rect 1211 1846 1212 1850
rect 1206 1845 1212 1846
rect 1350 1850 1356 1851
rect 1350 1846 1351 1850
rect 1355 1846 1356 1850
rect 1350 1845 1356 1846
rect 1200 1841 1210 1843
rect 454 1823 460 1824
rect 454 1819 455 1823
rect 459 1819 460 1823
rect 454 1818 460 1819
rect 838 1823 844 1824
rect 838 1819 839 1823
rect 843 1819 844 1823
rect 838 1818 844 1819
rect 1078 1823 1084 1824
rect 1078 1819 1079 1823
rect 1083 1819 1084 1823
rect 1078 1818 1084 1819
rect 438 1812 444 1813
rect 438 1808 439 1812
rect 443 1808 444 1812
rect 438 1807 444 1808
rect 590 1812 596 1813
rect 590 1808 591 1812
rect 595 1808 596 1812
rect 590 1807 596 1808
rect 742 1812 748 1813
rect 742 1808 743 1812
rect 747 1808 748 1812
rect 742 1807 748 1808
rect 894 1812 900 1813
rect 894 1808 895 1812
rect 899 1808 900 1812
rect 894 1807 900 1808
rect 1046 1812 1052 1813
rect 1046 1808 1047 1812
rect 1051 1808 1052 1812
rect 1046 1807 1052 1808
rect 1198 1812 1204 1813
rect 1198 1808 1199 1812
rect 1203 1808 1204 1812
rect 1208 1811 1210 1841
rect 1404 1824 1406 1854
rect 1488 1851 1490 1861
rect 1538 1859 1544 1860
rect 1538 1855 1539 1859
rect 1543 1855 1544 1859
rect 1538 1854 1544 1855
rect 1486 1850 1492 1851
rect 1486 1846 1487 1850
rect 1491 1846 1492 1850
rect 1486 1845 1492 1846
rect 1540 1824 1542 1854
rect 1632 1851 1634 1861
rect 1682 1859 1688 1860
rect 1682 1855 1683 1859
rect 1687 1855 1688 1859
rect 1682 1854 1688 1855
rect 1630 1850 1636 1851
rect 1630 1846 1631 1850
rect 1635 1846 1636 1850
rect 1630 1845 1636 1846
rect 1684 1824 1686 1854
rect 1752 1851 1754 1861
rect 1750 1850 1756 1851
rect 1750 1846 1751 1850
rect 1755 1846 1756 1850
rect 1750 1845 1756 1846
rect 1832 1833 1834 1861
rect 1872 1850 1874 1869
rect 1896 1853 1898 1869
rect 1894 1852 1900 1853
rect 1870 1849 1876 1850
rect 1870 1845 1871 1849
rect 1875 1845 1876 1849
rect 1894 1848 1895 1852
rect 1899 1848 1900 1852
rect 1894 1847 1900 1848
rect 1870 1844 1876 1845
rect 1830 1832 1836 1833
rect 1830 1828 1831 1832
rect 1835 1828 1836 1832
rect 1830 1827 1836 1828
rect 1870 1832 1876 1833
rect 1870 1828 1871 1832
rect 1875 1828 1876 1832
rect 1870 1827 1876 1828
rect 1402 1823 1408 1824
rect 1402 1819 1403 1823
rect 1407 1819 1408 1823
rect 1402 1818 1408 1819
rect 1538 1823 1544 1824
rect 1538 1819 1539 1823
rect 1543 1819 1544 1823
rect 1538 1818 1544 1819
rect 1682 1823 1688 1824
rect 1682 1819 1683 1823
rect 1687 1819 1688 1823
rect 1682 1818 1688 1819
rect 1830 1815 1836 1816
rect 1342 1812 1348 1813
rect 1208 1809 1214 1811
rect 1198 1807 1204 1808
rect 440 1787 442 1807
rect 592 1787 594 1807
rect 744 1787 746 1807
rect 766 1795 772 1796
rect 766 1791 767 1795
rect 771 1791 772 1795
rect 766 1790 772 1791
rect 439 1786 443 1787
rect 439 1781 443 1782
rect 591 1786 595 1787
rect 591 1781 595 1782
rect 743 1786 747 1787
rect 743 1781 747 1782
rect 751 1786 755 1787
rect 751 1781 755 1782
rect 592 1765 594 1781
rect 752 1765 754 1781
rect 590 1764 596 1765
rect 590 1760 591 1764
rect 595 1760 596 1764
rect 590 1759 596 1760
rect 750 1764 756 1765
rect 750 1760 751 1764
rect 755 1760 756 1764
rect 750 1759 756 1760
rect 582 1755 588 1756
rect 342 1750 348 1751
rect 430 1751 436 1752
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 110 1739 116 1740
rect 112 1707 114 1739
rect 254 1726 260 1727
rect 254 1722 255 1726
rect 259 1722 260 1726
rect 254 1721 260 1722
rect 256 1707 258 1721
rect 344 1716 346 1750
rect 430 1747 431 1751
rect 435 1747 436 1751
rect 582 1751 583 1755
rect 587 1751 588 1755
rect 582 1750 588 1751
rect 678 1755 684 1756
rect 678 1751 679 1755
rect 683 1751 684 1755
rect 678 1750 684 1751
rect 430 1746 436 1747
rect 430 1726 436 1727
rect 430 1722 431 1726
rect 435 1722 436 1726
rect 430 1721 436 1722
rect 342 1715 348 1716
rect 342 1711 343 1715
rect 347 1711 348 1715
rect 342 1710 348 1711
rect 432 1707 434 1721
rect 454 1707 460 1708
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 191 1706 195 1707
rect 191 1701 195 1702
rect 255 1706 259 1707
rect 255 1701 259 1702
rect 311 1706 315 1707
rect 311 1701 315 1702
rect 431 1706 435 1707
rect 431 1701 435 1702
rect 447 1706 451 1707
rect 454 1703 455 1707
rect 459 1703 460 1707
rect 454 1702 460 1703
rect 447 1701 451 1702
rect 112 1673 114 1701
rect 174 1699 180 1700
rect 174 1695 175 1699
rect 179 1695 180 1699
rect 174 1694 180 1695
rect 110 1672 116 1673
rect 110 1668 111 1672
rect 115 1668 116 1672
rect 110 1667 116 1668
rect 110 1655 116 1656
rect 110 1651 111 1655
rect 115 1651 116 1655
rect 110 1650 116 1651
rect 112 1623 114 1650
rect 111 1622 115 1623
rect 111 1617 115 1618
rect 167 1622 171 1623
rect 167 1617 171 1618
rect 112 1598 114 1617
rect 168 1601 170 1617
rect 166 1600 172 1601
rect 110 1597 116 1598
rect 110 1593 111 1597
rect 115 1593 116 1597
rect 166 1596 167 1600
rect 171 1596 172 1600
rect 166 1595 172 1596
rect 110 1592 116 1593
rect 176 1588 178 1694
rect 192 1691 194 1701
rect 242 1699 248 1700
rect 242 1695 243 1699
rect 247 1695 248 1699
rect 242 1694 248 1695
rect 190 1690 196 1691
rect 190 1686 191 1690
rect 195 1686 196 1690
rect 190 1685 196 1686
rect 244 1664 246 1694
rect 312 1691 314 1701
rect 362 1699 368 1700
rect 362 1695 363 1699
rect 367 1695 368 1699
rect 362 1694 368 1695
rect 310 1690 316 1691
rect 310 1686 311 1690
rect 315 1686 316 1690
rect 310 1685 316 1686
rect 364 1664 366 1694
rect 448 1691 450 1701
rect 446 1690 452 1691
rect 446 1686 447 1690
rect 451 1686 452 1690
rect 446 1685 452 1686
rect 456 1664 458 1702
rect 584 1700 586 1750
rect 598 1726 604 1727
rect 598 1722 599 1726
rect 603 1722 604 1726
rect 598 1721 604 1722
rect 600 1707 602 1721
rect 680 1716 682 1750
rect 758 1726 764 1727
rect 758 1722 759 1726
rect 763 1722 764 1726
rect 758 1721 764 1722
rect 678 1715 684 1716
rect 678 1711 679 1715
rect 683 1711 684 1715
rect 678 1710 684 1711
rect 760 1707 762 1721
rect 768 1716 770 1790
rect 896 1787 898 1807
rect 1048 1787 1050 1807
rect 1200 1787 1202 1807
rect 895 1786 899 1787
rect 895 1781 899 1782
rect 1023 1786 1027 1787
rect 1023 1781 1027 1782
rect 1047 1786 1051 1787
rect 1047 1781 1051 1782
rect 1143 1786 1147 1787
rect 1143 1781 1147 1782
rect 1199 1786 1203 1787
rect 1199 1781 1203 1782
rect 896 1765 898 1781
rect 1024 1765 1026 1781
rect 1144 1765 1146 1781
rect 894 1764 900 1765
rect 894 1760 895 1764
rect 899 1760 900 1764
rect 894 1759 900 1760
rect 1022 1764 1028 1765
rect 1022 1760 1023 1764
rect 1027 1760 1028 1764
rect 1022 1759 1028 1760
rect 1142 1764 1148 1765
rect 1142 1760 1143 1764
rect 1147 1760 1148 1764
rect 1142 1759 1148 1760
rect 1212 1756 1214 1809
rect 1342 1808 1343 1812
rect 1347 1808 1348 1812
rect 1342 1807 1348 1808
rect 1478 1812 1484 1813
rect 1478 1808 1479 1812
rect 1483 1808 1484 1812
rect 1478 1807 1484 1808
rect 1622 1812 1628 1813
rect 1622 1808 1623 1812
rect 1627 1808 1628 1812
rect 1622 1807 1628 1808
rect 1742 1812 1748 1813
rect 1742 1808 1743 1812
rect 1747 1808 1748 1812
rect 1830 1811 1831 1815
rect 1835 1811 1836 1815
rect 1830 1810 1836 1811
rect 1742 1807 1748 1808
rect 1344 1787 1346 1807
rect 1480 1787 1482 1807
rect 1624 1787 1626 1807
rect 1744 1787 1746 1807
rect 1832 1787 1834 1810
rect 1872 1787 1874 1827
rect 1902 1814 1908 1815
rect 1902 1810 1903 1814
rect 1907 1810 1908 1814
rect 1902 1809 1908 1810
rect 1904 1787 1906 1809
rect 1912 1804 1914 1874
rect 1991 1869 1995 1870
rect 1999 1874 2003 1875
rect 1999 1869 2003 1870
rect 2119 1874 2123 1875
rect 2119 1869 2123 1870
rect 2127 1874 2131 1875
rect 2127 1869 2131 1870
rect 2247 1874 2251 1875
rect 2247 1869 2251 1870
rect 1992 1853 1994 1869
rect 2120 1853 2122 1869
rect 2248 1853 2250 1869
rect 1990 1852 1996 1853
rect 1990 1848 1991 1852
rect 1995 1848 1996 1852
rect 1990 1847 1996 1848
rect 2118 1852 2124 1853
rect 2118 1848 2119 1852
rect 2123 1848 2124 1852
rect 2118 1847 2124 1848
rect 2246 1852 2252 1853
rect 2246 1848 2247 1852
rect 2251 1848 2252 1852
rect 2246 1847 2252 1848
rect 2352 1844 2354 1938
rect 2376 1935 2378 1945
rect 2384 1944 2386 1967
rect 2448 1956 2450 1990
rect 2600 1973 2602 1990
rect 2599 1972 2603 1973
rect 2599 1967 2603 1968
rect 2526 1966 2532 1967
rect 2526 1962 2527 1966
rect 2531 1962 2532 1966
rect 2526 1961 2532 1962
rect 2686 1966 2692 1967
rect 2686 1962 2687 1966
rect 2691 1962 2692 1966
rect 2686 1961 2692 1962
rect 2446 1955 2452 1956
rect 2446 1951 2447 1955
rect 2451 1951 2452 1955
rect 2528 1951 2530 1961
rect 2688 1951 2690 1961
rect 2748 1956 2750 1990
rect 2854 1966 2860 1967
rect 2854 1962 2855 1966
rect 2859 1962 2860 1966
rect 2854 1961 2860 1962
rect 2746 1955 2752 1956
rect 2746 1951 2747 1955
rect 2751 1951 2752 1955
rect 2856 1951 2858 1961
rect 2916 1956 2918 1990
rect 3022 1966 3028 1967
rect 3022 1962 3023 1966
rect 3027 1962 3028 1966
rect 3022 1961 3028 1962
rect 2914 1955 2920 1956
rect 2914 1951 2915 1955
rect 2919 1951 2920 1955
rect 3024 1951 3026 1961
rect 3032 1956 3034 2030
rect 3072 2027 3074 2047
rect 3184 2027 3186 2047
rect 3296 2027 3298 2047
rect 3408 2027 3410 2047
rect 3071 2026 3075 2027
rect 3071 2021 3075 2022
rect 3183 2026 3187 2027
rect 3183 2021 3187 2022
rect 3295 2026 3299 2027
rect 3295 2021 3299 2022
rect 3351 2026 3355 2027
rect 3351 2021 3355 2022
rect 3407 2026 3411 2027
rect 3407 2021 3411 2022
rect 3184 2005 3186 2021
rect 3352 2005 3354 2021
rect 3182 2004 3188 2005
rect 3182 2000 3183 2004
rect 3187 2000 3188 2004
rect 3182 1999 3188 2000
rect 3350 2004 3356 2005
rect 3350 2000 3351 2004
rect 3355 2000 3356 2004
rect 3350 1999 3356 2000
rect 3432 1996 3434 2094
rect 3512 2091 3514 2101
rect 3510 2090 3516 2091
rect 3510 2086 3511 2090
rect 3515 2086 3516 2090
rect 3510 2085 3516 2086
rect 3592 2073 3594 2101
rect 3590 2072 3596 2073
rect 3590 2068 3591 2072
rect 3595 2068 3596 2072
rect 3590 2067 3596 2068
rect 3590 2055 3596 2056
rect 3502 2052 3508 2053
rect 3502 2048 3503 2052
rect 3507 2048 3508 2052
rect 3590 2051 3591 2055
rect 3595 2051 3596 2055
rect 3590 2050 3596 2051
rect 3502 2047 3508 2048
rect 3504 2027 3506 2047
rect 3518 2035 3524 2036
rect 3518 2031 3519 2035
rect 3523 2031 3524 2035
rect 3518 2030 3524 2031
rect 3503 2026 3507 2027
rect 3503 2021 3507 2022
rect 3504 2005 3506 2021
rect 3502 2004 3508 2005
rect 3502 2000 3503 2004
rect 3507 2000 3508 2004
rect 3502 1999 3508 2000
rect 3274 1995 3280 1996
rect 3274 1991 3275 1995
rect 3279 1991 3280 1995
rect 3274 1990 3280 1991
rect 3430 1995 3436 1996
rect 3430 1991 3431 1995
rect 3435 1991 3436 1995
rect 3430 1990 3436 1991
rect 3262 1987 3268 1988
rect 3262 1983 3263 1987
rect 3267 1983 3268 1987
rect 3262 1982 3268 1983
rect 3190 1966 3196 1967
rect 3190 1962 3191 1966
rect 3195 1962 3196 1966
rect 3190 1961 3196 1962
rect 3030 1955 3036 1956
rect 3030 1951 3031 1955
rect 3035 1951 3036 1955
rect 3192 1951 3194 1961
rect 3264 1956 3266 1982
rect 3276 1956 3278 1990
rect 3358 1966 3364 1967
rect 3358 1962 3359 1966
rect 3363 1962 3364 1966
rect 3358 1961 3364 1962
rect 3510 1966 3516 1967
rect 3510 1962 3511 1966
rect 3515 1962 3516 1966
rect 3510 1961 3516 1962
rect 3262 1955 3268 1956
rect 3262 1951 3263 1955
rect 3267 1951 3268 1955
rect 2446 1950 2452 1951
rect 2487 1950 2491 1951
rect 2487 1945 2491 1946
rect 2527 1950 2531 1951
rect 2527 1945 2531 1946
rect 2599 1950 2603 1951
rect 2599 1945 2603 1946
rect 2687 1950 2691 1951
rect 2687 1945 2691 1946
rect 2719 1950 2723 1951
rect 2746 1950 2752 1951
rect 2839 1950 2843 1951
rect 2719 1945 2723 1946
rect 2839 1945 2843 1946
rect 2855 1950 2859 1951
rect 2914 1950 2920 1951
rect 3023 1950 3027 1951
rect 3030 1950 3036 1951
rect 3191 1950 3195 1951
rect 3262 1950 3268 1951
rect 3274 1955 3280 1956
rect 3274 1951 3275 1955
rect 3279 1951 3280 1955
rect 3360 1951 3362 1961
rect 3512 1951 3514 1961
rect 3520 1956 3522 2030
rect 3592 2027 3594 2050
rect 3591 2026 3595 2027
rect 3591 2021 3595 2022
rect 3592 2002 3594 2021
rect 3590 2001 3596 2002
rect 3590 1997 3591 2001
rect 3595 1997 3596 2001
rect 3590 1996 3596 1997
rect 3590 1984 3596 1985
rect 3590 1980 3591 1984
rect 3595 1980 3596 1984
rect 3590 1979 3596 1980
rect 3518 1955 3524 1956
rect 3518 1951 3519 1955
rect 3523 1951 3524 1955
rect 3592 1951 3594 1979
rect 3274 1950 3280 1951
rect 3359 1950 3363 1951
rect 2855 1945 2859 1946
rect 3023 1945 3027 1946
rect 3191 1945 3195 1946
rect 3359 1945 3363 1946
rect 3511 1950 3515 1951
rect 3518 1950 3524 1951
rect 3591 1950 3595 1951
rect 3511 1945 3515 1946
rect 3591 1945 3595 1946
rect 2382 1943 2388 1944
rect 2382 1939 2383 1943
rect 2387 1939 2388 1943
rect 2382 1938 2388 1939
rect 2426 1943 2432 1944
rect 2426 1939 2427 1943
rect 2431 1939 2432 1943
rect 2426 1938 2432 1939
rect 2374 1934 2380 1935
rect 2374 1930 2375 1934
rect 2379 1930 2380 1934
rect 2374 1929 2380 1930
rect 2428 1908 2430 1938
rect 2488 1935 2490 1945
rect 2538 1943 2544 1944
rect 2538 1939 2539 1943
rect 2543 1939 2544 1943
rect 2538 1938 2544 1939
rect 2486 1934 2492 1935
rect 2486 1930 2487 1934
rect 2491 1930 2492 1934
rect 2486 1929 2492 1930
rect 2540 1908 2542 1938
rect 2600 1935 2602 1945
rect 2650 1943 2656 1944
rect 2650 1939 2651 1943
rect 2655 1939 2656 1943
rect 2650 1938 2656 1939
rect 2598 1934 2604 1935
rect 2598 1930 2599 1934
rect 2603 1930 2604 1934
rect 2598 1929 2604 1930
rect 2652 1908 2654 1938
rect 2720 1935 2722 1945
rect 2770 1943 2776 1944
rect 2770 1939 2771 1943
rect 2775 1939 2776 1943
rect 2770 1938 2776 1939
rect 2718 1934 2724 1935
rect 2718 1930 2719 1934
rect 2723 1930 2724 1934
rect 2718 1929 2724 1930
rect 2772 1908 2774 1938
rect 2840 1935 2842 1945
rect 2838 1934 2844 1935
rect 2838 1930 2839 1934
rect 2843 1930 2844 1934
rect 2838 1929 2844 1930
rect 3592 1917 3594 1945
rect 3590 1916 3596 1917
rect 3590 1912 3591 1916
rect 3595 1912 3596 1916
rect 3590 1911 3596 1912
rect 2426 1907 2432 1908
rect 2426 1903 2427 1907
rect 2431 1903 2432 1907
rect 2426 1902 2432 1903
rect 2538 1907 2544 1908
rect 2538 1903 2539 1907
rect 2543 1903 2544 1907
rect 2538 1902 2544 1903
rect 2650 1907 2656 1908
rect 2650 1903 2651 1907
rect 2655 1903 2656 1907
rect 2650 1902 2656 1903
rect 2770 1907 2776 1908
rect 2770 1903 2771 1907
rect 2775 1903 2776 1907
rect 2770 1902 2776 1903
rect 3590 1899 3596 1900
rect 2366 1896 2372 1897
rect 2366 1892 2367 1896
rect 2371 1892 2372 1896
rect 2366 1891 2372 1892
rect 2478 1896 2484 1897
rect 2478 1892 2479 1896
rect 2483 1892 2484 1896
rect 2478 1891 2484 1892
rect 2590 1896 2596 1897
rect 2590 1892 2591 1896
rect 2595 1892 2596 1896
rect 2590 1891 2596 1892
rect 2710 1896 2716 1897
rect 2710 1892 2711 1896
rect 2715 1892 2716 1896
rect 2710 1891 2716 1892
rect 2830 1896 2836 1897
rect 2830 1892 2831 1896
rect 2835 1892 2836 1896
rect 3590 1895 3591 1899
rect 3595 1895 3596 1899
rect 3590 1894 3596 1895
rect 2830 1891 2836 1892
rect 2368 1875 2370 1891
rect 2480 1875 2482 1891
rect 2534 1879 2540 1880
rect 2534 1875 2535 1879
rect 2539 1875 2540 1879
rect 2592 1875 2594 1891
rect 2712 1875 2714 1891
rect 2832 1875 2834 1891
rect 3592 1875 3594 1894
rect 2367 1874 2371 1875
rect 2367 1869 2371 1870
rect 2383 1874 2387 1875
rect 2383 1869 2387 1870
rect 2479 1874 2483 1875
rect 2479 1869 2483 1870
rect 2519 1874 2523 1875
rect 2534 1874 2540 1875
rect 2591 1874 2595 1875
rect 2519 1869 2523 1870
rect 2384 1853 2386 1869
rect 2520 1853 2522 1869
rect 2382 1852 2388 1853
rect 2382 1848 2383 1852
rect 2387 1848 2388 1852
rect 2382 1847 2388 1848
rect 2518 1852 2524 1853
rect 2518 1848 2519 1852
rect 2523 1848 2524 1852
rect 2518 1847 2524 1848
rect 1962 1843 1968 1844
rect 1962 1839 1963 1843
rect 1967 1839 1968 1843
rect 1962 1838 1968 1839
rect 1970 1843 1976 1844
rect 1970 1839 1971 1843
rect 1975 1839 1976 1843
rect 1970 1838 1976 1839
rect 2190 1843 2196 1844
rect 2190 1839 2191 1843
rect 2195 1839 2196 1843
rect 2190 1838 2196 1839
rect 2342 1843 2348 1844
rect 2342 1839 2343 1843
rect 2347 1839 2348 1843
rect 2342 1838 2348 1839
rect 2350 1843 2356 1844
rect 2350 1839 2351 1843
rect 2355 1839 2356 1843
rect 2350 1838 2356 1839
rect 1964 1804 1966 1838
rect 1910 1803 1916 1804
rect 1910 1799 1911 1803
rect 1915 1799 1916 1803
rect 1910 1798 1916 1799
rect 1962 1803 1968 1804
rect 1962 1799 1963 1803
rect 1967 1799 1968 1803
rect 1962 1798 1968 1799
rect 1972 1788 1974 1838
rect 1998 1814 2004 1815
rect 1998 1810 1999 1814
rect 2003 1810 2004 1814
rect 1998 1809 2004 1810
rect 2126 1814 2132 1815
rect 2126 1810 2127 1814
rect 2131 1810 2132 1814
rect 2126 1809 2132 1810
rect 1970 1787 1976 1788
rect 2000 1787 2002 1809
rect 2128 1787 2130 1809
rect 2192 1804 2194 1838
rect 2254 1814 2260 1815
rect 2254 1810 2255 1814
rect 2259 1810 2260 1814
rect 2254 1809 2260 1810
rect 2190 1803 2196 1804
rect 2190 1799 2191 1803
rect 2195 1799 2196 1803
rect 2190 1798 2196 1799
rect 2256 1787 2258 1809
rect 2344 1804 2346 1838
rect 2390 1814 2396 1815
rect 2390 1810 2391 1814
rect 2395 1810 2396 1814
rect 2390 1809 2396 1810
rect 2526 1814 2532 1815
rect 2526 1810 2527 1814
rect 2531 1810 2532 1814
rect 2526 1809 2532 1810
rect 2342 1803 2348 1804
rect 2342 1799 2343 1803
rect 2347 1799 2348 1803
rect 2342 1798 2348 1799
rect 2392 1787 2394 1809
rect 2528 1787 2530 1809
rect 2536 1804 2538 1874
rect 2591 1869 2595 1870
rect 2655 1874 2659 1875
rect 2655 1869 2659 1870
rect 2711 1874 2715 1875
rect 2711 1869 2715 1870
rect 2807 1874 2811 1875
rect 2807 1869 2811 1870
rect 2831 1874 2835 1875
rect 2831 1869 2835 1870
rect 2975 1874 2979 1875
rect 2975 1869 2979 1870
rect 3151 1874 3155 1875
rect 3151 1869 3155 1870
rect 3335 1874 3339 1875
rect 3335 1869 3339 1870
rect 3503 1874 3507 1875
rect 3503 1869 3507 1870
rect 3591 1874 3595 1875
rect 3591 1869 3595 1870
rect 2656 1853 2658 1869
rect 2808 1853 2810 1869
rect 2976 1853 2978 1869
rect 3152 1853 3154 1869
rect 3336 1853 3338 1869
rect 3504 1853 3506 1869
rect 2654 1852 2660 1853
rect 2654 1848 2655 1852
rect 2659 1848 2660 1852
rect 2654 1847 2660 1848
rect 2806 1852 2812 1853
rect 2806 1848 2807 1852
rect 2811 1848 2812 1852
rect 2806 1847 2812 1848
rect 2974 1852 2980 1853
rect 2974 1848 2975 1852
rect 2979 1848 2980 1852
rect 2974 1847 2980 1848
rect 3150 1852 3156 1853
rect 3150 1848 3151 1852
rect 3155 1848 3156 1852
rect 3150 1847 3156 1848
rect 3334 1852 3340 1853
rect 3334 1848 3335 1852
rect 3339 1848 3340 1852
rect 3334 1847 3340 1848
rect 3502 1852 3508 1853
rect 3502 1848 3503 1852
rect 3507 1848 3508 1852
rect 3592 1850 3594 1869
rect 3502 1847 3508 1848
rect 3590 1849 3596 1850
rect 3590 1845 3591 1849
rect 3595 1845 3596 1849
rect 3590 1844 3596 1845
rect 2594 1843 2600 1844
rect 2594 1839 2595 1843
rect 2599 1839 2600 1843
rect 2594 1838 2600 1839
rect 2730 1843 2736 1844
rect 2730 1839 2731 1843
rect 2735 1839 2736 1843
rect 2730 1838 2736 1839
rect 2898 1843 2904 1844
rect 2898 1839 2899 1843
rect 2903 1839 2904 1843
rect 2898 1838 2904 1839
rect 3050 1843 3056 1844
rect 3050 1839 3051 1843
rect 3055 1839 3056 1843
rect 3050 1838 3056 1839
rect 3250 1843 3256 1844
rect 3250 1839 3251 1843
rect 3255 1839 3256 1843
rect 3250 1838 3256 1839
rect 3258 1843 3264 1844
rect 3258 1839 3259 1843
rect 3263 1839 3264 1843
rect 3258 1838 3264 1839
rect 3502 1839 3508 1840
rect 2596 1804 2598 1838
rect 2662 1814 2668 1815
rect 2662 1810 2663 1814
rect 2667 1810 2668 1814
rect 2662 1809 2668 1810
rect 2534 1803 2540 1804
rect 2534 1799 2535 1803
rect 2539 1799 2540 1803
rect 2534 1798 2540 1799
rect 2594 1803 2600 1804
rect 2594 1799 2595 1803
rect 2599 1799 2600 1803
rect 2594 1798 2600 1799
rect 2664 1787 2666 1809
rect 2732 1804 2734 1838
rect 2814 1814 2820 1815
rect 2814 1810 2815 1814
rect 2819 1810 2820 1814
rect 2814 1809 2820 1810
rect 2730 1803 2736 1804
rect 2730 1799 2731 1803
rect 2735 1799 2736 1803
rect 2730 1798 2736 1799
rect 2695 1796 2699 1797
rect 2695 1791 2699 1792
rect 1263 1786 1267 1787
rect 1263 1781 1267 1782
rect 1343 1786 1347 1787
rect 1343 1781 1347 1782
rect 1391 1786 1395 1787
rect 1391 1781 1395 1782
rect 1479 1786 1483 1787
rect 1479 1781 1483 1782
rect 1623 1786 1627 1787
rect 1623 1781 1627 1782
rect 1743 1786 1747 1787
rect 1743 1781 1747 1782
rect 1831 1786 1835 1787
rect 1831 1781 1835 1782
rect 1871 1786 1875 1787
rect 1871 1781 1875 1782
rect 1903 1786 1907 1787
rect 1970 1783 1971 1787
rect 1975 1783 1976 1787
rect 1970 1782 1976 1783
rect 1999 1786 2003 1787
rect 1903 1781 1907 1782
rect 1999 1781 2003 1782
rect 2031 1786 2035 1787
rect 2031 1781 2035 1782
rect 2127 1786 2131 1787
rect 2127 1781 2131 1782
rect 2191 1786 2195 1787
rect 2191 1781 2195 1782
rect 2255 1786 2259 1787
rect 2255 1781 2259 1782
rect 2359 1786 2363 1787
rect 2359 1781 2363 1782
rect 2391 1786 2395 1787
rect 2391 1781 2395 1782
rect 2527 1786 2531 1787
rect 2527 1781 2531 1782
rect 2663 1786 2667 1787
rect 2663 1781 2667 1782
rect 2687 1786 2691 1787
rect 2687 1781 2691 1782
rect 1264 1765 1266 1781
rect 1392 1765 1394 1781
rect 1262 1764 1268 1765
rect 1262 1760 1263 1764
rect 1267 1760 1268 1764
rect 1262 1759 1268 1760
rect 1390 1764 1396 1765
rect 1390 1760 1391 1764
rect 1395 1760 1396 1764
rect 1832 1762 1834 1781
rect 1390 1759 1396 1760
rect 1830 1761 1836 1762
rect 1830 1757 1831 1761
rect 1835 1757 1836 1761
rect 1830 1756 1836 1757
rect 966 1755 972 1756
rect 966 1751 967 1755
rect 971 1751 972 1755
rect 966 1750 972 1751
rect 1090 1755 1096 1756
rect 1090 1751 1091 1755
rect 1095 1751 1096 1755
rect 1090 1750 1096 1751
rect 1210 1755 1216 1756
rect 1210 1751 1211 1755
rect 1215 1751 1216 1755
rect 1210 1750 1216 1751
rect 1334 1755 1340 1756
rect 1334 1751 1335 1755
rect 1339 1751 1340 1755
rect 1334 1750 1340 1751
rect 1342 1755 1348 1756
rect 1342 1751 1343 1755
rect 1347 1751 1348 1755
rect 1872 1753 1874 1781
rect 1904 1771 1906 1781
rect 1954 1779 1960 1780
rect 1954 1775 1955 1779
rect 1959 1775 1960 1779
rect 1954 1774 1960 1775
rect 1902 1770 1908 1771
rect 1902 1766 1903 1770
rect 1907 1766 1908 1770
rect 1902 1765 1908 1766
rect 1342 1750 1348 1751
rect 1870 1752 1876 1753
rect 902 1726 908 1727
rect 902 1722 903 1726
rect 907 1722 908 1726
rect 902 1721 908 1722
rect 911 1724 915 1725
rect 766 1715 772 1716
rect 766 1711 767 1715
rect 771 1711 772 1715
rect 766 1710 772 1711
rect 904 1707 906 1721
rect 911 1719 915 1720
rect 912 1716 914 1719
rect 968 1716 970 1750
rect 1030 1726 1036 1727
rect 1030 1722 1031 1726
rect 1035 1722 1036 1726
rect 1030 1721 1036 1722
rect 910 1715 916 1716
rect 910 1711 911 1715
rect 915 1711 916 1715
rect 910 1710 916 1711
rect 966 1715 972 1716
rect 966 1711 967 1715
rect 971 1711 972 1715
rect 966 1710 972 1711
rect 1032 1707 1034 1721
rect 1092 1716 1094 1750
rect 1150 1726 1156 1727
rect 1150 1722 1151 1726
rect 1155 1722 1156 1726
rect 1150 1721 1156 1722
rect 1270 1726 1276 1727
rect 1270 1722 1271 1726
rect 1275 1722 1276 1726
rect 1270 1721 1276 1722
rect 1090 1715 1096 1716
rect 1090 1711 1091 1715
rect 1095 1711 1096 1715
rect 1090 1710 1096 1711
rect 1152 1707 1154 1721
rect 1234 1715 1240 1716
rect 1234 1711 1235 1715
rect 1239 1711 1240 1715
rect 1234 1710 1240 1711
rect 591 1706 595 1707
rect 591 1701 595 1702
rect 599 1706 603 1707
rect 599 1701 603 1702
rect 743 1706 747 1707
rect 743 1701 747 1702
rect 759 1706 763 1707
rect 759 1701 763 1702
rect 895 1706 899 1707
rect 895 1701 899 1702
rect 903 1706 907 1707
rect 903 1701 907 1702
rect 1031 1706 1035 1707
rect 1031 1701 1035 1702
rect 1039 1706 1043 1707
rect 1039 1701 1043 1702
rect 1151 1706 1155 1707
rect 1151 1701 1155 1702
rect 1183 1706 1187 1707
rect 1183 1701 1187 1702
rect 582 1699 588 1700
rect 582 1695 583 1699
rect 587 1695 588 1699
rect 582 1694 588 1695
rect 592 1691 594 1701
rect 642 1699 648 1700
rect 642 1695 643 1699
rect 647 1695 648 1699
rect 642 1694 648 1695
rect 590 1690 596 1691
rect 590 1686 591 1690
rect 595 1686 596 1690
rect 590 1685 596 1686
rect 644 1664 646 1694
rect 744 1691 746 1701
rect 794 1699 800 1700
rect 794 1695 795 1699
rect 799 1695 800 1699
rect 794 1694 800 1695
rect 742 1690 748 1691
rect 742 1686 743 1690
rect 747 1686 748 1690
rect 742 1685 748 1686
rect 796 1664 798 1694
rect 896 1691 898 1701
rect 946 1699 952 1700
rect 946 1695 947 1699
rect 951 1695 952 1699
rect 946 1694 952 1695
rect 894 1690 900 1691
rect 894 1686 895 1690
rect 899 1686 900 1690
rect 894 1685 900 1686
rect 948 1664 950 1694
rect 1040 1691 1042 1701
rect 1184 1691 1186 1701
rect 1038 1690 1044 1691
rect 1038 1686 1039 1690
rect 1043 1686 1044 1690
rect 1038 1685 1044 1686
rect 1182 1690 1188 1691
rect 1182 1686 1183 1690
rect 1187 1686 1188 1690
rect 1182 1685 1188 1686
rect 1236 1664 1238 1710
rect 1272 1707 1274 1721
rect 1336 1716 1338 1750
rect 1344 1725 1346 1750
rect 1870 1748 1871 1752
rect 1875 1748 1876 1752
rect 1870 1747 1876 1748
rect 1830 1744 1836 1745
rect 1956 1744 1958 1774
rect 2032 1771 2034 1781
rect 2082 1779 2088 1780
rect 2082 1775 2083 1779
rect 2087 1775 2088 1779
rect 2082 1774 2088 1775
rect 2030 1770 2036 1771
rect 2030 1766 2031 1770
rect 2035 1766 2036 1770
rect 2030 1765 2036 1766
rect 2084 1744 2086 1774
rect 2192 1771 2194 1781
rect 2242 1779 2248 1780
rect 2242 1775 2243 1779
rect 2247 1775 2248 1779
rect 2242 1774 2248 1775
rect 2190 1770 2196 1771
rect 2190 1766 2191 1770
rect 2195 1766 2196 1770
rect 2190 1765 2196 1766
rect 2244 1744 2246 1774
rect 2360 1771 2362 1781
rect 2410 1779 2416 1780
rect 2410 1775 2411 1779
rect 2415 1775 2416 1779
rect 2410 1774 2416 1775
rect 2358 1770 2364 1771
rect 2358 1766 2359 1770
rect 2363 1766 2364 1770
rect 2358 1765 2364 1766
rect 2412 1744 2414 1774
rect 2528 1771 2530 1781
rect 2688 1771 2690 1781
rect 2696 1780 2698 1791
rect 2816 1787 2818 1809
rect 2900 1804 2902 1838
rect 2982 1814 2988 1815
rect 2982 1810 2983 1814
rect 2987 1810 2988 1814
rect 2982 1809 2988 1810
rect 2898 1803 2904 1804
rect 2898 1799 2899 1803
rect 2903 1799 2904 1803
rect 2898 1798 2904 1799
rect 2984 1787 2986 1809
rect 3052 1804 3054 1838
rect 3158 1814 3164 1815
rect 3158 1810 3159 1814
rect 3163 1810 3164 1814
rect 3158 1809 3164 1810
rect 3050 1803 3056 1804
rect 3050 1799 3051 1803
rect 3055 1799 3056 1803
rect 3050 1798 3056 1799
rect 3160 1787 3162 1809
rect 3252 1804 3254 1838
rect 3250 1803 3256 1804
rect 3250 1799 3251 1803
rect 3255 1799 3256 1803
rect 3250 1798 3256 1799
rect 3260 1797 3262 1838
rect 3502 1835 3503 1839
rect 3507 1835 3508 1839
rect 3502 1834 3508 1835
rect 3342 1814 3348 1815
rect 3342 1810 3343 1814
rect 3347 1810 3348 1814
rect 3342 1809 3348 1810
rect 3259 1796 3263 1797
rect 3259 1791 3263 1792
rect 3344 1787 3346 1809
rect 2815 1786 2819 1787
rect 2815 1781 2819 1782
rect 2839 1786 2843 1787
rect 2839 1781 2843 1782
rect 2983 1786 2987 1787
rect 2983 1781 2987 1782
rect 3119 1786 3123 1787
rect 3119 1781 3123 1782
rect 3159 1786 3163 1787
rect 3159 1781 3163 1782
rect 3255 1786 3259 1787
rect 3255 1781 3259 1782
rect 3343 1786 3347 1787
rect 3343 1781 3347 1782
rect 3391 1786 3395 1787
rect 3391 1781 3395 1782
rect 2694 1779 2700 1780
rect 2694 1775 2695 1779
rect 2699 1775 2700 1779
rect 2694 1774 2700 1775
rect 2738 1779 2744 1780
rect 2738 1775 2739 1779
rect 2743 1775 2744 1779
rect 2738 1774 2744 1775
rect 2526 1770 2532 1771
rect 2526 1766 2527 1770
rect 2531 1766 2532 1770
rect 2526 1765 2532 1766
rect 2686 1770 2692 1771
rect 2686 1766 2687 1770
rect 2691 1766 2692 1770
rect 2686 1765 2692 1766
rect 2740 1744 2742 1774
rect 2840 1771 2842 1781
rect 2890 1779 2896 1780
rect 2890 1775 2891 1779
rect 2895 1775 2896 1779
rect 2890 1774 2896 1775
rect 2838 1770 2844 1771
rect 2838 1766 2839 1770
rect 2843 1766 2844 1770
rect 2838 1765 2844 1766
rect 2892 1744 2894 1774
rect 2984 1771 2986 1781
rect 3034 1779 3040 1780
rect 3034 1775 3035 1779
rect 3039 1775 3040 1779
rect 3034 1774 3040 1775
rect 2982 1770 2988 1771
rect 2982 1766 2983 1770
rect 2987 1766 2988 1770
rect 2982 1765 2988 1766
rect 3036 1744 3038 1774
rect 3120 1771 3122 1781
rect 3170 1779 3176 1780
rect 3170 1775 3171 1779
rect 3175 1775 3176 1779
rect 3170 1774 3176 1775
rect 3118 1770 3124 1771
rect 3118 1766 3119 1770
rect 3123 1766 3124 1770
rect 3118 1765 3124 1766
rect 3172 1744 3174 1774
rect 3256 1771 3258 1781
rect 3306 1779 3312 1780
rect 3306 1775 3307 1779
rect 3311 1775 3312 1779
rect 3306 1774 3312 1775
rect 3254 1770 3260 1771
rect 3254 1766 3255 1770
rect 3259 1766 3260 1770
rect 3254 1765 3260 1766
rect 3308 1744 3310 1774
rect 3392 1771 3394 1781
rect 3504 1780 3506 1834
rect 3590 1832 3596 1833
rect 3590 1828 3591 1832
rect 3595 1828 3596 1832
rect 3590 1827 3596 1828
rect 3510 1814 3516 1815
rect 3510 1810 3511 1814
rect 3515 1810 3516 1814
rect 3510 1809 3516 1810
rect 3512 1787 3514 1809
rect 3526 1803 3532 1804
rect 3526 1799 3527 1803
rect 3531 1799 3532 1803
rect 3526 1798 3532 1799
rect 3511 1786 3515 1787
rect 3511 1781 3515 1782
rect 3502 1779 3508 1780
rect 3502 1775 3503 1779
rect 3507 1775 3508 1779
rect 3502 1774 3508 1775
rect 3512 1771 3514 1781
rect 3390 1770 3396 1771
rect 3390 1766 3391 1770
rect 3395 1766 3396 1770
rect 3390 1765 3396 1766
rect 3510 1770 3516 1771
rect 3510 1766 3511 1770
rect 3515 1766 3516 1770
rect 3510 1765 3516 1766
rect 1830 1740 1831 1744
rect 1835 1740 1836 1744
rect 1830 1739 1836 1740
rect 1954 1743 1960 1744
rect 1954 1739 1955 1743
rect 1959 1739 1960 1743
rect 1398 1726 1404 1727
rect 1343 1724 1347 1725
rect 1398 1722 1399 1726
rect 1403 1722 1404 1726
rect 1398 1721 1404 1722
rect 1343 1719 1347 1720
rect 1334 1715 1340 1716
rect 1334 1711 1335 1715
rect 1339 1711 1340 1715
rect 1334 1710 1340 1711
rect 1400 1707 1402 1721
rect 1832 1707 1834 1739
rect 1954 1738 1960 1739
rect 2082 1743 2088 1744
rect 2082 1739 2083 1743
rect 2087 1739 2088 1743
rect 2082 1738 2088 1739
rect 2242 1743 2248 1744
rect 2242 1739 2243 1743
rect 2247 1739 2248 1743
rect 2242 1738 2248 1739
rect 2410 1743 2416 1744
rect 2410 1739 2411 1743
rect 2415 1739 2416 1743
rect 2410 1738 2416 1739
rect 2738 1743 2744 1744
rect 2738 1739 2739 1743
rect 2743 1739 2744 1743
rect 2738 1738 2744 1739
rect 2890 1743 2896 1744
rect 2890 1739 2891 1743
rect 2895 1739 2896 1743
rect 2890 1738 2896 1739
rect 3034 1743 3040 1744
rect 3034 1739 3035 1743
rect 3039 1739 3040 1743
rect 3034 1738 3040 1739
rect 3170 1743 3176 1744
rect 3170 1739 3171 1743
rect 3175 1739 3176 1743
rect 3170 1738 3176 1739
rect 3306 1743 3312 1744
rect 3306 1739 3307 1743
rect 3311 1739 3312 1743
rect 3306 1738 3312 1739
rect 1870 1735 1876 1736
rect 1870 1731 1871 1735
rect 1875 1731 1876 1735
rect 1870 1730 1876 1731
rect 1894 1732 1900 1733
rect 1872 1707 1874 1730
rect 1894 1728 1895 1732
rect 1899 1728 1900 1732
rect 1894 1727 1900 1728
rect 2022 1732 2028 1733
rect 2022 1728 2023 1732
rect 2027 1728 2028 1732
rect 2022 1727 2028 1728
rect 2182 1732 2188 1733
rect 2182 1728 2183 1732
rect 2187 1728 2188 1732
rect 2182 1727 2188 1728
rect 2350 1732 2356 1733
rect 2350 1728 2351 1732
rect 2355 1728 2356 1732
rect 2350 1727 2356 1728
rect 2518 1732 2524 1733
rect 2518 1728 2519 1732
rect 2523 1728 2524 1732
rect 2518 1727 2524 1728
rect 2678 1732 2684 1733
rect 2678 1728 2679 1732
rect 2683 1728 2684 1732
rect 2678 1727 2684 1728
rect 2830 1732 2836 1733
rect 2830 1728 2831 1732
rect 2835 1728 2836 1732
rect 2830 1727 2836 1728
rect 2974 1732 2980 1733
rect 2974 1728 2975 1732
rect 2979 1728 2980 1732
rect 2974 1727 2980 1728
rect 3110 1732 3116 1733
rect 3110 1728 3111 1732
rect 3115 1728 3116 1732
rect 3110 1727 3116 1728
rect 3246 1732 3252 1733
rect 3246 1728 3247 1732
rect 3251 1728 3252 1732
rect 3246 1727 3252 1728
rect 3382 1732 3388 1733
rect 3382 1728 3383 1732
rect 3387 1728 3388 1732
rect 3382 1727 3388 1728
rect 3502 1732 3508 1733
rect 3502 1728 3503 1732
rect 3507 1728 3508 1732
rect 3502 1727 3508 1728
rect 1896 1707 1898 1727
rect 2024 1707 2026 1727
rect 2184 1707 2186 1727
rect 2352 1707 2354 1727
rect 2418 1715 2424 1716
rect 2418 1711 2419 1715
rect 2423 1711 2424 1715
rect 2418 1710 2424 1711
rect 1271 1706 1275 1707
rect 1271 1701 1275 1702
rect 1319 1706 1323 1707
rect 1319 1701 1323 1702
rect 1399 1706 1403 1707
rect 1399 1701 1403 1702
rect 1447 1706 1451 1707
rect 1447 1701 1451 1702
rect 1575 1706 1579 1707
rect 1575 1701 1579 1702
rect 1711 1706 1715 1707
rect 1711 1701 1715 1702
rect 1831 1706 1835 1707
rect 1831 1701 1835 1702
rect 1871 1706 1875 1707
rect 1871 1701 1875 1702
rect 1895 1706 1899 1707
rect 1895 1701 1899 1702
rect 1991 1706 1995 1707
rect 1991 1701 1995 1702
rect 2023 1706 2027 1707
rect 2023 1701 2027 1702
rect 2135 1706 2139 1707
rect 2135 1701 2139 1702
rect 2183 1706 2187 1707
rect 2183 1701 2187 1702
rect 2295 1706 2299 1707
rect 2295 1701 2299 1702
rect 2351 1706 2355 1707
rect 2351 1701 2355 1702
rect 1242 1699 1248 1700
rect 1242 1695 1243 1699
rect 1247 1695 1248 1699
rect 1242 1694 1248 1695
rect 1244 1664 1246 1694
rect 1320 1691 1322 1701
rect 1378 1699 1384 1700
rect 1378 1695 1379 1699
rect 1383 1695 1384 1699
rect 1378 1694 1384 1695
rect 1318 1690 1324 1691
rect 1318 1686 1319 1690
rect 1323 1686 1324 1690
rect 1318 1685 1324 1686
rect 1380 1664 1382 1694
rect 1448 1691 1450 1701
rect 1576 1691 1578 1701
rect 1634 1699 1640 1700
rect 1634 1695 1635 1699
rect 1639 1695 1640 1699
rect 1634 1694 1640 1695
rect 1446 1690 1452 1691
rect 1446 1686 1447 1690
rect 1451 1686 1452 1690
rect 1446 1685 1452 1686
rect 1574 1690 1580 1691
rect 1574 1686 1575 1690
rect 1579 1686 1580 1690
rect 1574 1685 1580 1686
rect 1636 1664 1638 1694
rect 1712 1691 1714 1701
rect 1726 1699 1732 1700
rect 1726 1695 1727 1699
rect 1731 1695 1732 1699
rect 1726 1694 1732 1695
rect 1710 1690 1716 1691
rect 1710 1686 1711 1690
rect 1715 1686 1716 1690
rect 1710 1685 1716 1686
rect 242 1663 248 1664
rect 242 1659 243 1663
rect 247 1659 248 1663
rect 242 1658 248 1659
rect 362 1663 368 1664
rect 362 1659 363 1663
rect 367 1659 368 1663
rect 362 1658 368 1659
rect 454 1663 460 1664
rect 454 1659 455 1663
rect 459 1659 460 1663
rect 454 1658 460 1659
rect 642 1663 648 1664
rect 642 1659 643 1663
rect 647 1659 648 1663
rect 642 1658 648 1659
rect 794 1663 800 1664
rect 794 1659 795 1663
rect 799 1659 800 1663
rect 794 1658 800 1659
rect 946 1663 952 1664
rect 946 1659 947 1663
rect 951 1659 952 1663
rect 946 1658 952 1659
rect 1234 1663 1240 1664
rect 1234 1659 1235 1663
rect 1239 1659 1240 1663
rect 1234 1658 1240 1659
rect 1242 1663 1248 1664
rect 1242 1659 1243 1663
rect 1247 1659 1248 1663
rect 1242 1658 1248 1659
rect 1378 1663 1384 1664
rect 1378 1659 1379 1663
rect 1383 1659 1384 1663
rect 1378 1658 1384 1659
rect 1634 1663 1640 1664
rect 1634 1659 1635 1663
rect 1639 1659 1640 1663
rect 1634 1658 1640 1659
rect 182 1652 188 1653
rect 182 1648 183 1652
rect 187 1648 188 1652
rect 182 1647 188 1648
rect 302 1652 308 1653
rect 302 1648 303 1652
rect 307 1648 308 1652
rect 302 1647 308 1648
rect 438 1652 444 1653
rect 438 1648 439 1652
rect 443 1648 444 1652
rect 438 1647 444 1648
rect 582 1652 588 1653
rect 582 1648 583 1652
rect 587 1648 588 1652
rect 582 1647 588 1648
rect 734 1652 740 1653
rect 734 1648 735 1652
rect 739 1648 740 1652
rect 734 1647 740 1648
rect 886 1652 892 1653
rect 886 1648 887 1652
rect 891 1648 892 1652
rect 886 1647 892 1648
rect 1030 1652 1036 1653
rect 1030 1648 1031 1652
rect 1035 1648 1036 1652
rect 1030 1647 1036 1648
rect 1174 1652 1180 1653
rect 1174 1648 1175 1652
rect 1179 1648 1180 1652
rect 1174 1647 1180 1648
rect 1310 1652 1316 1653
rect 1310 1648 1311 1652
rect 1315 1648 1316 1652
rect 1310 1647 1316 1648
rect 1438 1652 1444 1653
rect 1438 1648 1439 1652
rect 1443 1648 1444 1652
rect 1438 1647 1444 1648
rect 1566 1652 1572 1653
rect 1566 1648 1567 1652
rect 1571 1648 1572 1652
rect 1566 1647 1572 1648
rect 1702 1652 1708 1653
rect 1702 1648 1703 1652
rect 1707 1648 1708 1652
rect 1702 1647 1708 1648
rect 184 1623 186 1647
rect 304 1623 306 1647
rect 440 1623 442 1647
rect 584 1623 586 1647
rect 736 1623 738 1647
rect 888 1623 890 1647
rect 918 1635 924 1636
rect 918 1631 919 1635
rect 923 1631 924 1635
rect 918 1630 924 1631
rect 183 1622 187 1623
rect 183 1617 187 1618
rect 303 1622 307 1623
rect 303 1617 307 1618
rect 351 1622 355 1623
rect 351 1617 355 1618
rect 439 1622 443 1623
rect 439 1617 443 1618
rect 543 1622 547 1623
rect 543 1617 547 1618
rect 583 1622 587 1623
rect 583 1617 587 1618
rect 727 1622 731 1623
rect 727 1617 731 1618
rect 735 1622 739 1623
rect 735 1617 739 1618
rect 887 1622 891 1623
rect 887 1617 891 1618
rect 903 1622 907 1623
rect 903 1617 907 1618
rect 352 1601 354 1617
rect 544 1601 546 1617
rect 728 1601 730 1617
rect 904 1601 906 1617
rect 350 1600 356 1601
rect 350 1596 351 1600
rect 355 1596 356 1600
rect 350 1595 356 1596
rect 542 1600 548 1601
rect 542 1596 543 1600
rect 547 1596 548 1600
rect 542 1595 548 1596
rect 726 1600 732 1601
rect 726 1596 727 1600
rect 731 1596 732 1600
rect 726 1595 732 1596
rect 902 1600 908 1601
rect 902 1596 903 1600
rect 907 1596 908 1600
rect 902 1595 908 1596
rect 234 1591 240 1592
rect 174 1587 180 1588
rect 174 1583 175 1587
rect 179 1583 180 1587
rect 234 1587 235 1591
rect 239 1587 240 1591
rect 234 1586 240 1587
rect 418 1591 424 1592
rect 418 1587 419 1591
rect 423 1587 424 1591
rect 418 1586 424 1587
rect 610 1591 616 1592
rect 610 1587 611 1591
rect 615 1587 616 1591
rect 610 1586 616 1587
rect 794 1591 800 1592
rect 794 1587 795 1591
rect 799 1587 800 1591
rect 794 1586 800 1587
rect 174 1582 180 1583
rect 110 1580 116 1581
rect 110 1576 111 1580
rect 115 1576 116 1580
rect 110 1575 116 1576
rect 112 1543 114 1575
rect 174 1562 180 1563
rect 174 1558 175 1562
rect 179 1558 180 1562
rect 174 1557 180 1558
rect 176 1543 178 1557
rect 236 1552 238 1586
rect 358 1562 364 1563
rect 358 1558 359 1562
rect 363 1558 364 1562
rect 358 1557 364 1558
rect 234 1551 240 1552
rect 234 1547 235 1551
rect 239 1547 240 1551
rect 234 1546 240 1547
rect 298 1551 304 1552
rect 298 1547 299 1551
rect 303 1547 304 1551
rect 298 1546 304 1547
rect 111 1542 115 1543
rect 111 1537 115 1538
rect 143 1542 147 1543
rect 143 1537 147 1538
rect 175 1542 179 1543
rect 175 1537 179 1538
rect 247 1542 251 1543
rect 247 1537 251 1538
rect 112 1509 114 1537
rect 144 1527 146 1537
rect 194 1535 200 1536
rect 194 1531 195 1535
rect 199 1531 200 1535
rect 194 1530 200 1531
rect 142 1526 148 1527
rect 142 1522 143 1526
rect 147 1522 148 1526
rect 142 1521 148 1522
rect 110 1508 116 1509
rect 110 1504 111 1508
rect 115 1504 116 1508
rect 110 1503 116 1504
rect 196 1500 198 1530
rect 248 1527 250 1537
rect 246 1526 252 1527
rect 246 1522 247 1526
rect 251 1522 252 1526
rect 246 1521 252 1522
rect 300 1500 302 1546
rect 360 1543 362 1557
rect 359 1542 363 1543
rect 359 1537 363 1538
rect 383 1542 387 1543
rect 383 1537 387 1538
rect 384 1527 386 1537
rect 420 1536 422 1586
rect 550 1562 556 1563
rect 550 1558 551 1562
rect 555 1558 556 1562
rect 550 1557 556 1558
rect 552 1543 554 1557
rect 612 1552 614 1586
rect 734 1562 740 1563
rect 734 1558 735 1562
rect 739 1558 740 1562
rect 734 1557 740 1558
rect 610 1551 616 1552
rect 610 1547 611 1551
rect 615 1547 616 1551
rect 610 1546 616 1547
rect 736 1543 738 1557
rect 796 1552 798 1586
rect 910 1562 916 1563
rect 910 1558 911 1562
rect 915 1558 916 1562
rect 910 1557 916 1558
rect 794 1551 800 1552
rect 794 1547 795 1551
rect 799 1547 800 1551
rect 794 1546 800 1547
rect 912 1543 914 1557
rect 920 1552 922 1630
rect 1032 1623 1034 1647
rect 1176 1623 1178 1647
rect 1312 1623 1314 1647
rect 1440 1623 1442 1647
rect 1568 1623 1570 1647
rect 1704 1623 1706 1647
rect 1031 1622 1035 1623
rect 1031 1617 1035 1618
rect 1071 1622 1075 1623
rect 1071 1617 1075 1618
rect 1175 1622 1179 1623
rect 1175 1617 1179 1618
rect 1223 1622 1227 1623
rect 1223 1617 1227 1618
rect 1311 1622 1315 1623
rect 1311 1617 1315 1618
rect 1359 1622 1363 1623
rect 1359 1617 1363 1618
rect 1439 1622 1443 1623
rect 1439 1617 1443 1618
rect 1495 1622 1499 1623
rect 1495 1617 1499 1618
rect 1567 1622 1571 1623
rect 1567 1617 1571 1618
rect 1623 1622 1627 1623
rect 1623 1617 1627 1618
rect 1703 1622 1707 1623
rect 1703 1617 1707 1618
rect 1072 1601 1074 1617
rect 1224 1601 1226 1617
rect 1360 1601 1362 1617
rect 1496 1601 1498 1617
rect 1624 1601 1626 1617
rect 1070 1600 1076 1601
rect 1070 1596 1071 1600
rect 1075 1596 1076 1600
rect 1070 1595 1076 1596
rect 1222 1600 1228 1601
rect 1222 1596 1223 1600
rect 1227 1596 1228 1600
rect 1222 1595 1228 1596
rect 1358 1600 1364 1601
rect 1358 1596 1359 1600
rect 1363 1596 1364 1600
rect 1358 1595 1364 1596
rect 1494 1600 1500 1601
rect 1494 1596 1495 1600
rect 1499 1596 1500 1600
rect 1494 1595 1500 1596
rect 1622 1600 1628 1601
rect 1622 1596 1623 1600
rect 1627 1596 1628 1600
rect 1622 1595 1628 1596
rect 1728 1592 1730 1694
rect 1832 1673 1834 1701
rect 1872 1682 1874 1701
rect 1896 1685 1898 1701
rect 1911 1692 1915 1693
rect 1911 1687 1915 1688
rect 1894 1684 1900 1685
rect 1870 1681 1876 1682
rect 1870 1677 1871 1681
rect 1875 1677 1876 1681
rect 1894 1680 1895 1684
rect 1899 1680 1900 1684
rect 1894 1679 1900 1680
rect 1870 1676 1876 1677
rect 1830 1672 1836 1673
rect 1830 1668 1831 1672
rect 1835 1668 1836 1672
rect 1830 1667 1836 1668
rect 1870 1664 1876 1665
rect 1870 1660 1871 1664
rect 1875 1660 1876 1664
rect 1870 1659 1876 1660
rect 1830 1655 1836 1656
rect 1830 1651 1831 1655
rect 1835 1651 1836 1655
rect 1830 1650 1836 1651
rect 1832 1623 1834 1650
rect 1872 1627 1874 1659
rect 1902 1646 1908 1647
rect 1902 1642 1903 1646
rect 1907 1642 1908 1646
rect 1902 1641 1908 1642
rect 1904 1627 1906 1641
rect 1912 1636 1914 1687
rect 1992 1685 1994 1701
rect 2136 1685 2138 1701
rect 2296 1685 2298 1701
rect 2420 1693 2422 1710
rect 2520 1707 2522 1727
rect 2680 1707 2682 1727
rect 2832 1707 2834 1727
rect 2976 1707 2978 1727
rect 3112 1707 3114 1727
rect 3248 1707 3250 1727
rect 3384 1707 3386 1727
rect 3398 1715 3404 1716
rect 3398 1711 3399 1715
rect 3403 1711 3404 1715
rect 3398 1710 3404 1711
rect 2471 1706 2475 1707
rect 2471 1701 2475 1702
rect 2519 1706 2523 1707
rect 2519 1701 2523 1702
rect 2647 1706 2651 1707
rect 2647 1701 2651 1702
rect 2679 1706 2683 1707
rect 2679 1701 2683 1702
rect 2815 1706 2819 1707
rect 2815 1701 2819 1702
rect 2831 1706 2835 1707
rect 2831 1701 2835 1702
rect 2967 1706 2971 1707
rect 2967 1701 2971 1702
rect 2975 1706 2979 1707
rect 2975 1701 2979 1702
rect 3111 1706 3115 1707
rect 3111 1701 3115 1702
rect 3247 1706 3251 1707
rect 3247 1701 3251 1702
rect 3383 1706 3387 1707
rect 3383 1701 3387 1702
rect 2419 1692 2423 1693
rect 2419 1687 2423 1688
rect 2472 1685 2474 1701
rect 2648 1685 2650 1701
rect 2816 1685 2818 1701
rect 2968 1685 2970 1701
rect 3112 1685 3114 1701
rect 3248 1685 3250 1701
rect 3384 1685 3386 1701
rect 1990 1684 1996 1685
rect 1990 1680 1991 1684
rect 1995 1680 1996 1684
rect 1990 1679 1996 1680
rect 2134 1684 2140 1685
rect 2134 1680 2135 1684
rect 2139 1680 2140 1684
rect 2134 1679 2140 1680
rect 2294 1684 2300 1685
rect 2294 1680 2295 1684
rect 2299 1680 2300 1684
rect 2294 1679 2300 1680
rect 2470 1684 2476 1685
rect 2470 1680 2471 1684
rect 2475 1680 2476 1684
rect 2470 1679 2476 1680
rect 2646 1684 2652 1685
rect 2646 1680 2647 1684
rect 2651 1680 2652 1684
rect 2646 1679 2652 1680
rect 2814 1684 2820 1685
rect 2814 1680 2815 1684
rect 2819 1680 2820 1684
rect 2814 1679 2820 1680
rect 2966 1684 2972 1685
rect 2966 1680 2967 1684
rect 2971 1680 2972 1684
rect 2966 1679 2972 1680
rect 3110 1684 3116 1685
rect 3110 1680 3111 1684
rect 3115 1680 3116 1684
rect 3110 1679 3116 1680
rect 3246 1684 3252 1685
rect 3246 1680 3247 1684
rect 3251 1680 3252 1684
rect 3246 1679 3252 1680
rect 3382 1684 3388 1685
rect 3382 1680 3383 1684
rect 3387 1680 3388 1684
rect 3382 1679 3388 1680
rect 1962 1675 1968 1676
rect 1962 1671 1963 1675
rect 1967 1671 1968 1675
rect 1962 1670 1968 1671
rect 2070 1675 2076 1676
rect 2070 1671 2071 1675
rect 2075 1671 2076 1675
rect 2070 1670 2076 1671
rect 2222 1675 2228 1676
rect 2222 1671 2223 1675
rect 2227 1671 2228 1675
rect 2222 1670 2228 1671
rect 2390 1675 2396 1676
rect 2390 1671 2391 1675
rect 2395 1671 2396 1675
rect 2390 1670 2396 1671
rect 2566 1675 2572 1676
rect 2566 1671 2567 1675
rect 2571 1671 2572 1675
rect 2566 1670 2572 1671
rect 2574 1675 2580 1676
rect 2574 1671 2575 1675
rect 2579 1671 2580 1675
rect 2574 1670 2580 1671
rect 2890 1675 2896 1676
rect 2890 1671 2891 1675
rect 2895 1671 2896 1675
rect 2890 1670 2896 1671
rect 3046 1675 3052 1676
rect 3046 1671 3047 1675
rect 3051 1671 3052 1675
rect 3046 1670 3052 1671
rect 3178 1675 3184 1676
rect 3178 1671 3179 1675
rect 3183 1671 3184 1675
rect 3178 1670 3184 1671
rect 3186 1675 3192 1676
rect 3186 1671 3187 1675
rect 3191 1671 3192 1675
rect 3186 1670 3192 1671
rect 3322 1675 3328 1676
rect 3322 1671 3323 1675
rect 3327 1671 3328 1675
rect 3322 1670 3328 1671
rect 1964 1636 1966 1670
rect 1998 1646 2004 1647
rect 1998 1642 1999 1646
rect 2003 1642 2004 1646
rect 1998 1641 2004 1642
rect 1910 1635 1916 1636
rect 1910 1631 1911 1635
rect 1915 1631 1916 1635
rect 1910 1630 1916 1631
rect 1962 1635 1968 1636
rect 1962 1631 1963 1635
rect 1967 1631 1968 1635
rect 1962 1630 1968 1631
rect 2000 1627 2002 1641
rect 2072 1636 2074 1670
rect 2142 1646 2148 1647
rect 2142 1642 2143 1646
rect 2147 1642 2148 1646
rect 2142 1641 2148 1642
rect 2070 1635 2076 1636
rect 2070 1631 2071 1635
rect 2075 1631 2076 1635
rect 2070 1630 2076 1631
rect 2144 1627 2146 1641
rect 2224 1636 2226 1670
rect 2302 1646 2308 1647
rect 2302 1642 2303 1646
rect 2307 1642 2308 1646
rect 2302 1641 2308 1642
rect 2222 1635 2228 1636
rect 2222 1631 2223 1635
rect 2227 1631 2228 1635
rect 2222 1630 2228 1631
rect 2304 1627 2306 1641
rect 2392 1636 2394 1670
rect 2478 1646 2484 1647
rect 2478 1642 2479 1646
rect 2483 1642 2484 1646
rect 2478 1641 2484 1642
rect 2390 1635 2396 1636
rect 2390 1631 2391 1635
rect 2395 1631 2396 1635
rect 2390 1630 2396 1631
rect 2480 1627 2482 1641
rect 2568 1636 2570 1670
rect 2566 1635 2572 1636
rect 2566 1631 2567 1635
rect 2571 1631 2572 1635
rect 2566 1630 2572 1631
rect 2576 1628 2578 1670
rect 2654 1646 2660 1647
rect 2654 1642 2655 1646
rect 2659 1642 2660 1646
rect 2654 1641 2660 1642
rect 2822 1646 2828 1647
rect 2822 1642 2823 1646
rect 2827 1642 2828 1646
rect 2822 1641 2828 1642
rect 2831 1644 2835 1645
rect 2574 1627 2580 1628
rect 2656 1627 2658 1641
rect 2824 1627 2826 1641
rect 2831 1639 2835 1640
rect 2832 1636 2834 1639
rect 2892 1636 2894 1670
rect 2974 1646 2980 1647
rect 2974 1642 2975 1646
rect 2979 1642 2980 1646
rect 2974 1641 2980 1642
rect 2830 1635 2836 1636
rect 2830 1631 2831 1635
rect 2835 1631 2836 1635
rect 2830 1630 2836 1631
rect 2890 1635 2896 1636
rect 2890 1631 2891 1635
rect 2895 1631 2896 1635
rect 2890 1630 2896 1631
rect 2976 1627 2978 1641
rect 3048 1636 3050 1670
rect 3118 1646 3124 1647
rect 3118 1642 3119 1646
rect 3123 1642 3124 1646
rect 3118 1641 3124 1642
rect 3046 1635 3052 1636
rect 3046 1631 3047 1635
rect 3051 1631 3052 1635
rect 3046 1630 3052 1631
rect 3062 1627 3068 1628
rect 3120 1627 3122 1641
rect 1871 1626 1875 1627
rect 1743 1622 1747 1623
rect 1743 1617 1747 1618
rect 1831 1622 1835 1623
rect 1871 1621 1875 1622
rect 1903 1626 1907 1627
rect 1903 1621 1907 1622
rect 1975 1626 1979 1627
rect 1975 1621 1979 1622
rect 1999 1626 2003 1627
rect 1999 1621 2003 1622
rect 2095 1626 2099 1627
rect 2095 1621 2099 1622
rect 2143 1626 2147 1627
rect 2143 1621 2147 1622
rect 2231 1626 2235 1627
rect 2231 1621 2235 1622
rect 2303 1626 2307 1627
rect 2303 1621 2307 1622
rect 2367 1626 2371 1627
rect 2367 1621 2371 1622
rect 2479 1626 2483 1627
rect 2479 1621 2483 1622
rect 2503 1626 2507 1627
rect 2574 1623 2575 1627
rect 2579 1623 2580 1627
rect 2574 1622 2580 1623
rect 2639 1626 2643 1627
rect 2503 1621 2507 1622
rect 2639 1621 2643 1622
rect 2655 1626 2659 1627
rect 2655 1621 2659 1622
rect 2775 1626 2779 1627
rect 2775 1621 2779 1622
rect 2823 1626 2827 1627
rect 2823 1621 2827 1622
rect 2911 1626 2915 1627
rect 2911 1621 2915 1622
rect 2975 1626 2979 1627
rect 2975 1621 2979 1622
rect 3055 1626 3059 1627
rect 3062 1623 3063 1627
rect 3067 1623 3068 1627
rect 3062 1622 3068 1623
rect 3119 1626 3123 1627
rect 3055 1621 3059 1622
rect 1831 1617 1835 1618
rect 1744 1601 1746 1617
rect 1742 1600 1748 1601
rect 1742 1596 1743 1600
rect 1747 1596 1748 1600
rect 1832 1598 1834 1617
rect 1742 1595 1748 1596
rect 1830 1597 1836 1598
rect 1830 1593 1831 1597
rect 1835 1593 1836 1597
rect 1872 1593 1874 1621
rect 1976 1611 1978 1621
rect 2026 1619 2032 1620
rect 2026 1615 2027 1619
rect 2031 1615 2032 1619
rect 2026 1614 2032 1615
rect 1974 1610 1980 1611
rect 1974 1606 1975 1610
rect 1979 1606 1980 1610
rect 1974 1605 1980 1606
rect 1830 1592 1836 1593
rect 1870 1592 1876 1593
rect 1154 1591 1160 1592
rect 1154 1587 1155 1591
rect 1159 1587 1160 1591
rect 1154 1586 1160 1587
rect 1290 1591 1296 1592
rect 1290 1587 1291 1591
rect 1295 1587 1296 1591
rect 1290 1586 1296 1587
rect 1426 1591 1432 1592
rect 1426 1587 1427 1591
rect 1431 1587 1432 1591
rect 1426 1586 1432 1587
rect 1566 1591 1572 1592
rect 1566 1587 1567 1591
rect 1571 1587 1572 1591
rect 1566 1586 1572 1587
rect 1690 1591 1696 1592
rect 1690 1587 1691 1591
rect 1695 1587 1696 1591
rect 1690 1586 1696 1587
rect 1726 1591 1732 1592
rect 1726 1587 1727 1591
rect 1731 1587 1732 1591
rect 1870 1588 1871 1592
rect 1875 1588 1876 1592
rect 1870 1587 1876 1588
rect 1726 1586 1732 1587
rect 1078 1562 1084 1563
rect 1078 1558 1079 1562
rect 1083 1558 1084 1562
rect 1078 1557 1084 1558
rect 918 1551 924 1552
rect 918 1547 919 1551
rect 923 1547 924 1551
rect 918 1546 924 1547
rect 1080 1543 1082 1557
rect 1156 1552 1158 1586
rect 1230 1562 1236 1563
rect 1230 1558 1231 1562
rect 1235 1558 1236 1562
rect 1230 1557 1236 1558
rect 1154 1551 1160 1552
rect 1154 1547 1155 1551
rect 1159 1547 1160 1551
rect 1154 1546 1160 1547
rect 1232 1543 1234 1557
rect 1292 1552 1294 1586
rect 1366 1562 1372 1563
rect 1366 1558 1367 1562
rect 1371 1558 1372 1562
rect 1366 1557 1372 1558
rect 1290 1551 1296 1552
rect 1290 1547 1291 1551
rect 1295 1547 1296 1551
rect 1290 1546 1296 1547
rect 1368 1543 1370 1557
rect 1428 1552 1430 1586
rect 1502 1562 1508 1563
rect 1502 1558 1503 1562
rect 1507 1558 1508 1562
rect 1502 1557 1508 1558
rect 1426 1551 1432 1552
rect 1426 1547 1427 1551
rect 1431 1547 1432 1551
rect 1426 1546 1432 1547
rect 1478 1543 1484 1544
rect 1504 1543 1506 1557
rect 1568 1552 1570 1586
rect 1630 1562 1636 1563
rect 1630 1558 1631 1562
rect 1635 1558 1636 1562
rect 1630 1557 1636 1558
rect 1566 1551 1572 1552
rect 1566 1547 1567 1551
rect 1571 1547 1572 1551
rect 1566 1546 1572 1547
rect 1632 1543 1634 1557
rect 1692 1552 1694 1586
rect 2028 1584 2030 1614
rect 2096 1611 2098 1621
rect 2198 1619 2204 1620
rect 2198 1615 2199 1619
rect 2203 1615 2204 1619
rect 2198 1614 2204 1615
rect 2094 1610 2100 1611
rect 2094 1606 2095 1610
rect 2099 1606 2100 1610
rect 2094 1605 2100 1606
rect 2200 1584 2202 1614
rect 2232 1611 2234 1621
rect 2282 1619 2288 1620
rect 2282 1615 2283 1619
rect 2287 1615 2288 1619
rect 2282 1614 2288 1615
rect 2230 1610 2236 1611
rect 2230 1606 2231 1610
rect 2235 1606 2236 1610
rect 2230 1605 2236 1606
rect 2284 1584 2286 1614
rect 2368 1611 2370 1621
rect 2418 1619 2424 1620
rect 2418 1615 2419 1619
rect 2423 1615 2424 1619
rect 2418 1614 2424 1615
rect 2366 1610 2372 1611
rect 2366 1606 2367 1610
rect 2371 1606 2372 1610
rect 2366 1605 2372 1606
rect 2420 1584 2422 1614
rect 2504 1611 2506 1621
rect 2640 1611 2642 1621
rect 2690 1619 2696 1620
rect 2690 1615 2691 1619
rect 2695 1615 2696 1619
rect 2690 1614 2696 1615
rect 2502 1610 2508 1611
rect 2502 1606 2503 1610
rect 2507 1606 2508 1610
rect 2502 1605 2508 1606
rect 2638 1610 2644 1611
rect 2638 1606 2639 1610
rect 2643 1606 2644 1610
rect 2638 1605 2644 1606
rect 2692 1584 2694 1614
rect 2776 1611 2778 1621
rect 2866 1619 2872 1620
rect 2866 1615 2867 1619
rect 2871 1615 2872 1619
rect 2866 1614 2872 1615
rect 2774 1610 2780 1611
rect 2774 1606 2775 1610
rect 2779 1606 2780 1610
rect 2774 1605 2780 1606
rect 2868 1584 2870 1614
rect 2912 1611 2914 1621
rect 3056 1611 3058 1621
rect 2910 1610 2916 1611
rect 2910 1606 2911 1610
rect 2915 1606 2916 1610
rect 2910 1605 2916 1606
rect 3054 1610 3060 1611
rect 3054 1606 3055 1610
rect 3059 1606 3060 1610
rect 3054 1605 3060 1606
rect 3064 1584 3066 1622
rect 3119 1621 3123 1622
rect 3180 1620 3182 1670
rect 3188 1645 3190 1670
rect 3254 1646 3260 1647
rect 3187 1644 3191 1645
rect 3254 1642 3255 1646
rect 3259 1642 3260 1646
rect 3254 1641 3260 1642
rect 3187 1639 3191 1640
rect 3256 1627 3258 1641
rect 3324 1636 3326 1670
rect 3390 1646 3396 1647
rect 3390 1642 3391 1646
rect 3395 1642 3396 1646
rect 3390 1641 3396 1642
rect 3322 1635 3328 1636
rect 3322 1631 3323 1635
rect 3327 1631 3328 1635
rect 3322 1630 3328 1631
rect 3374 1627 3380 1628
rect 3392 1627 3394 1641
rect 3400 1636 3402 1710
rect 3504 1707 3506 1727
rect 3518 1715 3524 1716
rect 3518 1711 3519 1715
rect 3523 1711 3524 1715
rect 3518 1710 3524 1711
rect 3503 1706 3507 1707
rect 3503 1701 3507 1702
rect 3504 1685 3506 1701
rect 3502 1684 3508 1685
rect 3502 1680 3503 1684
rect 3507 1680 3508 1684
rect 3502 1679 3508 1680
rect 3510 1646 3516 1647
rect 3510 1642 3511 1646
rect 3515 1642 3516 1646
rect 3510 1641 3516 1642
rect 3398 1635 3404 1636
rect 3398 1631 3399 1635
rect 3403 1631 3404 1635
rect 3398 1630 3404 1631
rect 3512 1627 3514 1641
rect 3520 1636 3522 1710
rect 3518 1635 3524 1636
rect 3518 1631 3519 1635
rect 3523 1631 3524 1635
rect 3518 1630 3524 1631
rect 3207 1626 3211 1627
rect 3207 1621 3211 1622
rect 3255 1626 3259 1627
rect 3255 1621 3259 1622
rect 3367 1626 3371 1627
rect 3374 1623 3375 1627
rect 3379 1623 3380 1627
rect 3374 1622 3380 1623
rect 3391 1626 3395 1627
rect 3367 1621 3371 1622
rect 3178 1619 3184 1620
rect 3178 1615 3179 1619
rect 3183 1615 3184 1619
rect 3178 1614 3184 1615
rect 3208 1611 3210 1621
rect 3290 1619 3296 1620
rect 3290 1615 3291 1619
rect 3295 1615 3296 1619
rect 3290 1614 3296 1615
rect 3206 1610 3212 1611
rect 3206 1606 3207 1610
rect 3211 1606 3212 1610
rect 3206 1605 3212 1606
rect 3292 1584 3294 1614
rect 3368 1611 3370 1621
rect 3366 1610 3372 1611
rect 3366 1606 3367 1610
rect 3371 1606 3372 1610
rect 3366 1605 3372 1606
rect 3376 1584 3378 1622
rect 3391 1621 3395 1622
rect 3511 1626 3515 1627
rect 3511 1621 3515 1622
rect 3486 1619 3492 1620
rect 3486 1615 3487 1619
rect 3491 1615 3492 1619
rect 3486 1614 3492 1615
rect 2026 1583 2032 1584
rect 1830 1580 1836 1581
rect 1830 1576 1831 1580
rect 1835 1576 1836 1580
rect 2026 1579 2027 1583
rect 2031 1579 2032 1583
rect 2026 1578 2032 1579
rect 2198 1583 2204 1584
rect 2198 1579 2199 1583
rect 2203 1579 2204 1583
rect 2198 1578 2204 1579
rect 2282 1583 2288 1584
rect 2282 1579 2283 1583
rect 2287 1579 2288 1583
rect 2282 1578 2288 1579
rect 2418 1583 2424 1584
rect 2418 1579 2419 1583
rect 2423 1579 2424 1583
rect 2418 1578 2424 1579
rect 2690 1583 2696 1584
rect 2690 1579 2691 1583
rect 2695 1579 2696 1583
rect 2690 1578 2696 1579
rect 2866 1583 2872 1584
rect 2866 1579 2867 1583
rect 2871 1579 2872 1583
rect 2866 1578 2872 1579
rect 2934 1583 2940 1584
rect 2934 1579 2935 1583
rect 2939 1579 2940 1583
rect 2934 1578 2940 1579
rect 3062 1583 3068 1584
rect 3062 1579 3063 1583
rect 3067 1579 3068 1583
rect 3062 1578 3068 1579
rect 3290 1583 3296 1584
rect 3290 1579 3291 1583
rect 3295 1579 3296 1583
rect 3290 1578 3296 1579
rect 3374 1583 3380 1584
rect 3374 1579 3375 1583
rect 3379 1579 3380 1583
rect 3374 1578 3380 1579
rect 1830 1575 1836 1576
rect 1870 1575 1876 1576
rect 1750 1562 1756 1563
rect 1750 1558 1751 1562
rect 1755 1558 1756 1562
rect 1750 1557 1756 1558
rect 1690 1551 1696 1552
rect 1690 1547 1691 1551
rect 1695 1547 1696 1551
rect 1690 1546 1696 1547
rect 1752 1543 1754 1557
rect 1832 1543 1834 1575
rect 1870 1571 1871 1575
rect 1875 1571 1876 1575
rect 1870 1570 1876 1571
rect 1966 1572 1972 1573
rect 1872 1547 1874 1570
rect 1966 1568 1967 1572
rect 1971 1568 1972 1572
rect 1966 1567 1972 1568
rect 2086 1572 2092 1573
rect 2086 1568 2087 1572
rect 2091 1568 2092 1572
rect 2086 1567 2092 1568
rect 2222 1572 2228 1573
rect 2222 1568 2223 1572
rect 2227 1568 2228 1572
rect 2222 1567 2228 1568
rect 2358 1572 2364 1573
rect 2358 1568 2359 1572
rect 2363 1568 2364 1572
rect 2358 1567 2364 1568
rect 2494 1572 2500 1573
rect 2494 1568 2495 1572
rect 2499 1568 2500 1572
rect 2494 1567 2500 1568
rect 2630 1572 2636 1573
rect 2630 1568 2631 1572
rect 2635 1568 2636 1572
rect 2630 1567 2636 1568
rect 2766 1572 2772 1573
rect 2766 1568 2767 1572
rect 2771 1568 2772 1572
rect 2766 1567 2772 1568
rect 2902 1572 2908 1573
rect 2902 1568 2903 1572
rect 2907 1568 2908 1572
rect 2902 1567 2908 1568
rect 1968 1547 1970 1567
rect 2088 1547 2090 1567
rect 2224 1547 2226 1567
rect 2360 1547 2362 1567
rect 2418 1555 2424 1556
rect 2418 1551 2419 1555
rect 2423 1551 2424 1555
rect 2418 1550 2424 1551
rect 1871 1546 1875 1547
rect 527 1542 531 1543
rect 527 1537 531 1538
rect 551 1542 555 1543
rect 551 1537 555 1538
rect 671 1542 675 1543
rect 671 1537 675 1538
rect 735 1542 739 1543
rect 735 1537 739 1538
rect 815 1542 819 1543
rect 815 1537 819 1538
rect 911 1542 915 1543
rect 911 1537 915 1538
rect 951 1542 955 1543
rect 951 1537 955 1538
rect 1079 1542 1083 1543
rect 1079 1537 1083 1538
rect 1207 1542 1211 1543
rect 1207 1537 1211 1538
rect 1231 1542 1235 1543
rect 1231 1537 1235 1538
rect 1335 1542 1339 1543
rect 1335 1537 1339 1538
rect 1367 1542 1371 1543
rect 1367 1537 1371 1538
rect 1471 1542 1475 1543
rect 1478 1539 1479 1543
rect 1483 1539 1484 1543
rect 1478 1538 1484 1539
rect 1503 1542 1507 1543
rect 1471 1537 1475 1538
rect 418 1535 424 1536
rect 418 1531 419 1535
rect 423 1531 424 1535
rect 418 1530 424 1531
rect 434 1535 440 1536
rect 434 1531 435 1535
rect 439 1531 440 1535
rect 434 1530 440 1531
rect 382 1526 388 1527
rect 382 1522 383 1526
rect 387 1522 388 1526
rect 382 1521 388 1522
rect 436 1500 438 1530
rect 528 1527 530 1537
rect 578 1535 584 1536
rect 578 1531 579 1535
rect 583 1531 584 1535
rect 578 1530 584 1531
rect 526 1526 532 1527
rect 526 1522 527 1526
rect 531 1522 532 1526
rect 526 1521 532 1522
rect 580 1500 582 1530
rect 672 1527 674 1537
rect 722 1535 728 1536
rect 722 1531 723 1535
rect 727 1531 728 1535
rect 722 1530 728 1531
rect 670 1526 676 1527
rect 670 1522 671 1526
rect 675 1522 676 1526
rect 670 1521 676 1522
rect 724 1500 726 1530
rect 816 1527 818 1537
rect 952 1527 954 1537
rect 958 1535 964 1536
rect 958 1531 959 1535
rect 963 1531 964 1535
rect 958 1530 964 1531
rect 1002 1535 1008 1536
rect 1002 1531 1003 1535
rect 1007 1531 1008 1535
rect 1002 1530 1008 1531
rect 814 1526 820 1527
rect 814 1522 815 1526
rect 819 1522 820 1526
rect 814 1521 820 1522
rect 950 1526 956 1527
rect 950 1522 951 1526
rect 955 1522 956 1526
rect 950 1521 956 1522
rect 194 1499 200 1500
rect 194 1495 195 1499
rect 199 1495 200 1499
rect 194 1494 200 1495
rect 298 1499 304 1500
rect 298 1495 299 1499
rect 303 1495 304 1499
rect 298 1494 304 1495
rect 434 1499 440 1500
rect 434 1495 435 1499
rect 439 1495 440 1499
rect 434 1494 440 1495
rect 578 1499 584 1500
rect 578 1495 579 1499
rect 583 1495 584 1499
rect 578 1494 584 1495
rect 722 1499 728 1500
rect 722 1495 723 1499
rect 727 1495 728 1499
rect 722 1494 728 1495
rect 110 1491 116 1492
rect 110 1487 111 1491
rect 115 1487 116 1491
rect 110 1486 116 1487
rect 134 1488 140 1489
rect 112 1463 114 1486
rect 134 1484 135 1488
rect 139 1484 140 1488
rect 134 1483 140 1484
rect 238 1488 244 1489
rect 238 1484 239 1488
rect 243 1484 244 1488
rect 238 1483 244 1484
rect 374 1488 380 1489
rect 374 1484 375 1488
rect 379 1484 380 1488
rect 374 1483 380 1484
rect 518 1488 524 1489
rect 518 1484 519 1488
rect 523 1484 524 1488
rect 518 1483 524 1484
rect 662 1488 668 1489
rect 662 1484 663 1488
rect 667 1484 668 1488
rect 662 1483 668 1484
rect 806 1488 812 1489
rect 806 1484 807 1488
rect 811 1484 812 1488
rect 806 1483 812 1484
rect 942 1488 948 1489
rect 942 1484 943 1488
rect 947 1484 948 1488
rect 942 1483 948 1484
rect 136 1463 138 1483
rect 240 1463 242 1483
rect 376 1463 378 1483
rect 520 1463 522 1483
rect 614 1471 620 1472
rect 614 1467 615 1471
rect 619 1467 620 1471
rect 614 1466 620 1467
rect 111 1462 115 1463
rect 111 1457 115 1458
rect 135 1462 139 1463
rect 135 1457 139 1458
rect 231 1462 235 1463
rect 231 1457 235 1458
rect 239 1462 243 1463
rect 239 1457 243 1458
rect 359 1462 363 1463
rect 359 1457 363 1458
rect 375 1462 379 1463
rect 375 1457 379 1458
rect 479 1462 483 1463
rect 479 1457 483 1458
rect 519 1462 523 1463
rect 519 1457 523 1458
rect 599 1462 603 1463
rect 599 1457 603 1458
rect 112 1438 114 1457
rect 136 1441 138 1457
rect 232 1441 234 1457
rect 360 1441 362 1457
rect 480 1441 482 1457
rect 600 1441 602 1457
rect 134 1440 140 1441
rect 110 1437 116 1438
rect 110 1433 111 1437
rect 115 1433 116 1437
rect 134 1436 135 1440
rect 139 1436 140 1440
rect 134 1435 140 1436
rect 230 1440 236 1441
rect 230 1436 231 1440
rect 235 1436 236 1440
rect 230 1435 236 1436
rect 358 1440 364 1441
rect 358 1436 359 1440
rect 363 1436 364 1440
rect 358 1435 364 1436
rect 478 1440 484 1441
rect 478 1436 479 1440
rect 483 1436 484 1440
rect 478 1435 484 1436
rect 598 1440 604 1441
rect 598 1436 599 1440
rect 603 1436 604 1440
rect 598 1435 604 1436
rect 110 1432 116 1433
rect 202 1431 208 1432
rect 202 1427 203 1431
rect 207 1427 208 1431
rect 202 1426 208 1427
rect 298 1431 304 1432
rect 298 1427 299 1431
rect 303 1427 304 1431
rect 298 1426 304 1427
rect 426 1431 432 1432
rect 426 1427 427 1431
rect 431 1427 432 1431
rect 426 1426 432 1427
rect 546 1431 552 1432
rect 546 1427 547 1431
rect 551 1427 552 1431
rect 546 1426 552 1427
rect 110 1420 116 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 110 1415 116 1416
rect 112 1371 114 1415
rect 142 1402 148 1403
rect 142 1398 143 1402
rect 147 1398 148 1402
rect 204 1400 206 1426
rect 238 1402 244 1403
rect 142 1397 148 1398
rect 202 1399 208 1400
rect 144 1371 146 1397
rect 202 1395 203 1399
rect 207 1395 208 1399
rect 238 1398 239 1402
rect 243 1398 244 1402
rect 238 1397 244 1398
rect 202 1394 208 1395
rect 194 1391 200 1392
rect 194 1387 195 1391
rect 199 1387 200 1391
rect 194 1386 200 1387
rect 111 1370 115 1371
rect 111 1365 115 1366
rect 143 1370 147 1371
rect 143 1365 147 1366
rect 112 1337 114 1365
rect 144 1355 146 1365
rect 142 1354 148 1355
rect 142 1350 143 1354
rect 147 1350 148 1354
rect 142 1349 148 1350
rect 110 1336 116 1337
rect 110 1332 111 1336
rect 115 1332 116 1336
rect 110 1331 116 1332
rect 196 1328 198 1386
rect 240 1371 242 1397
rect 239 1370 243 1371
rect 239 1365 243 1366
rect 287 1370 291 1371
rect 287 1365 291 1366
rect 288 1355 290 1365
rect 300 1364 302 1426
rect 366 1402 372 1403
rect 366 1398 367 1402
rect 371 1398 372 1402
rect 366 1397 372 1398
rect 368 1371 370 1397
rect 428 1392 430 1426
rect 486 1402 492 1403
rect 486 1398 487 1402
rect 491 1398 492 1402
rect 486 1397 492 1398
rect 426 1391 432 1392
rect 426 1387 427 1391
rect 431 1387 432 1391
rect 426 1386 432 1387
rect 488 1371 490 1397
rect 548 1392 550 1426
rect 606 1402 612 1403
rect 606 1398 607 1402
rect 611 1398 612 1402
rect 606 1397 612 1398
rect 546 1391 552 1392
rect 546 1387 547 1391
rect 551 1387 552 1391
rect 546 1386 552 1387
rect 608 1371 610 1397
rect 616 1392 618 1466
rect 664 1463 666 1483
rect 808 1463 810 1483
rect 944 1463 946 1483
rect 960 1477 962 1530
rect 1004 1500 1006 1530
rect 1080 1527 1082 1537
rect 1130 1535 1136 1536
rect 1130 1531 1131 1535
rect 1135 1531 1136 1535
rect 1130 1530 1136 1531
rect 1078 1526 1084 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1132 1500 1134 1530
rect 1208 1527 1210 1537
rect 1258 1535 1264 1536
rect 1258 1531 1259 1535
rect 1263 1531 1264 1535
rect 1258 1530 1264 1531
rect 1206 1526 1212 1527
rect 1206 1522 1207 1526
rect 1211 1522 1212 1526
rect 1206 1521 1212 1522
rect 1260 1500 1262 1530
rect 1336 1527 1338 1537
rect 1386 1535 1392 1536
rect 1386 1531 1387 1535
rect 1391 1531 1392 1535
rect 1386 1530 1392 1531
rect 1334 1526 1340 1527
rect 1334 1522 1335 1526
rect 1339 1522 1340 1526
rect 1334 1521 1340 1522
rect 1388 1500 1390 1530
rect 1472 1527 1474 1537
rect 1470 1526 1476 1527
rect 1470 1522 1471 1526
rect 1475 1522 1476 1526
rect 1470 1521 1476 1522
rect 1480 1500 1482 1538
rect 1503 1537 1507 1538
rect 1631 1542 1635 1543
rect 1631 1537 1635 1538
rect 1751 1542 1755 1543
rect 1751 1537 1755 1538
rect 1831 1542 1835 1543
rect 1871 1541 1875 1542
rect 1967 1546 1971 1547
rect 1967 1541 1971 1542
rect 2087 1546 2091 1547
rect 2087 1541 2091 1542
rect 2167 1546 2171 1547
rect 2167 1541 2171 1542
rect 2223 1546 2227 1547
rect 2223 1541 2227 1542
rect 2255 1546 2259 1547
rect 2255 1541 2259 1542
rect 2343 1546 2347 1547
rect 2343 1541 2347 1542
rect 2359 1546 2363 1547
rect 2359 1541 2363 1542
rect 1831 1537 1835 1538
rect 1832 1509 1834 1537
rect 1872 1522 1874 1541
rect 2088 1525 2090 1541
rect 2103 1532 2107 1533
rect 2103 1527 2107 1528
rect 2086 1524 2092 1525
rect 1870 1521 1876 1522
rect 1870 1517 1871 1521
rect 1875 1517 1876 1521
rect 2086 1520 2087 1524
rect 2091 1520 2092 1524
rect 2086 1519 2092 1520
rect 1870 1516 1876 1517
rect 1830 1508 1836 1509
rect 1830 1504 1831 1508
rect 1835 1504 1836 1508
rect 1830 1503 1836 1504
rect 1870 1504 1876 1505
rect 1870 1500 1871 1504
rect 1875 1500 1876 1504
rect 1002 1499 1008 1500
rect 1002 1495 1003 1499
rect 1007 1495 1008 1499
rect 1002 1494 1008 1495
rect 1130 1499 1136 1500
rect 1130 1495 1131 1499
rect 1135 1495 1136 1499
rect 1130 1494 1136 1495
rect 1258 1499 1264 1500
rect 1258 1495 1259 1499
rect 1263 1495 1264 1499
rect 1258 1494 1264 1495
rect 1386 1499 1392 1500
rect 1386 1495 1387 1499
rect 1391 1495 1392 1499
rect 1386 1494 1392 1495
rect 1478 1499 1484 1500
rect 1870 1499 1876 1500
rect 1478 1495 1479 1499
rect 1483 1495 1484 1499
rect 1478 1494 1484 1495
rect 1830 1491 1836 1492
rect 1070 1488 1076 1489
rect 1070 1484 1071 1488
rect 1075 1484 1076 1488
rect 1070 1483 1076 1484
rect 1198 1488 1204 1489
rect 1198 1484 1199 1488
rect 1203 1484 1204 1488
rect 1198 1483 1204 1484
rect 1326 1488 1332 1489
rect 1326 1484 1327 1488
rect 1331 1484 1332 1488
rect 1326 1483 1332 1484
rect 1462 1488 1468 1489
rect 1462 1484 1463 1488
rect 1467 1484 1468 1488
rect 1830 1487 1831 1491
rect 1835 1487 1836 1491
rect 1830 1486 1836 1487
rect 1462 1483 1468 1484
rect 959 1476 963 1477
rect 959 1471 963 1472
rect 1072 1463 1074 1483
rect 1200 1463 1202 1483
rect 1219 1476 1223 1477
rect 1219 1471 1223 1472
rect 663 1462 667 1463
rect 663 1457 667 1458
rect 719 1462 723 1463
rect 719 1457 723 1458
rect 807 1462 811 1463
rect 807 1457 811 1458
rect 831 1462 835 1463
rect 831 1457 835 1458
rect 935 1462 939 1463
rect 935 1457 939 1458
rect 943 1462 947 1463
rect 943 1457 947 1458
rect 1039 1462 1043 1463
rect 1039 1457 1043 1458
rect 1071 1462 1075 1463
rect 1071 1457 1075 1458
rect 1143 1462 1147 1463
rect 1143 1457 1147 1458
rect 1199 1462 1203 1463
rect 1199 1457 1203 1458
rect 720 1441 722 1457
rect 832 1441 834 1457
rect 936 1441 938 1457
rect 1040 1441 1042 1457
rect 1144 1441 1146 1457
rect 718 1440 724 1441
rect 718 1436 719 1440
rect 723 1436 724 1440
rect 718 1435 724 1436
rect 830 1440 836 1441
rect 830 1436 831 1440
rect 835 1436 836 1440
rect 830 1435 836 1436
rect 934 1440 940 1441
rect 934 1436 935 1440
rect 939 1436 940 1440
rect 934 1435 940 1436
rect 1038 1440 1044 1441
rect 1038 1436 1039 1440
rect 1043 1436 1044 1440
rect 1038 1435 1044 1436
rect 1142 1440 1148 1441
rect 1142 1436 1143 1440
rect 1147 1436 1148 1440
rect 1142 1435 1148 1436
rect 1220 1432 1222 1471
rect 1328 1463 1330 1483
rect 1464 1463 1466 1483
rect 1832 1463 1834 1486
rect 1872 1467 1874 1499
rect 2094 1486 2100 1487
rect 2094 1482 2095 1486
rect 2099 1482 2100 1486
rect 2094 1481 2100 1482
rect 2096 1467 2098 1481
rect 2104 1476 2106 1527
rect 2168 1525 2170 1541
rect 2256 1525 2258 1541
rect 2344 1525 2346 1541
rect 2420 1533 2422 1550
rect 2496 1547 2498 1567
rect 2632 1547 2634 1567
rect 2768 1547 2770 1567
rect 2904 1547 2906 1567
rect 2439 1546 2443 1547
rect 2439 1541 2443 1542
rect 2495 1546 2499 1547
rect 2495 1541 2499 1542
rect 2535 1546 2539 1547
rect 2535 1541 2539 1542
rect 2631 1546 2635 1547
rect 2631 1541 2635 1542
rect 2647 1546 2651 1547
rect 2647 1541 2651 1542
rect 2767 1546 2771 1547
rect 2767 1541 2771 1542
rect 2783 1546 2787 1547
rect 2783 1541 2787 1542
rect 2903 1546 2907 1547
rect 2903 1541 2907 1542
rect 2419 1532 2423 1533
rect 2419 1527 2423 1528
rect 2440 1525 2442 1541
rect 2536 1525 2538 1541
rect 2648 1525 2650 1541
rect 2784 1525 2786 1541
rect 2166 1524 2172 1525
rect 2166 1520 2167 1524
rect 2171 1520 2172 1524
rect 2166 1519 2172 1520
rect 2254 1524 2260 1525
rect 2254 1520 2255 1524
rect 2259 1520 2260 1524
rect 2254 1519 2260 1520
rect 2342 1524 2348 1525
rect 2342 1520 2343 1524
rect 2347 1520 2348 1524
rect 2342 1519 2348 1520
rect 2438 1524 2444 1525
rect 2438 1520 2439 1524
rect 2443 1520 2444 1524
rect 2438 1519 2444 1520
rect 2534 1524 2540 1525
rect 2534 1520 2535 1524
rect 2539 1520 2540 1524
rect 2534 1519 2540 1520
rect 2646 1524 2652 1525
rect 2646 1520 2647 1524
rect 2651 1520 2652 1524
rect 2646 1519 2652 1520
rect 2782 1524 2788 1525
rect 2782 1520 2783 1524
rect 2787 1520 2788 1524
rect 2782 1519 2788 1520
rect 2154 1515 2160 1516
rect 2154 1511 2155 1515
rect 2159 1511 2160 1515
rect 2154 1510 2160 1511
rect 2234 1515 2240 1516
rect 2234 1511 2235 1515
rect 2239 1511 2240 1515
rect 2234 1510 2240 1511
rect 2322 1515 2328 1516
rect 2322 1511 2323 1515
rect 2327 1511 2328 1515
rect 2322 1510 2328 1511
rect 2410 1515 2416 1516
rect 2410 1511 2411 1515
rect 2415 1511 2416 1515
rect 2410 1510 2416 1511
rect 2506 1515 2512 1516
rect 2506 1511 2507 1515
rect 2511 1511 2512 1515
rect 2722 1515 2728 1516
rect 2506 1510 2512 1511
rect 2514 1511 2520 1512
rect 2156 1476 2158 1510
rect 2174 1486 2180 1487
rect 2174 1482 2175 1486
rect 2179 1482 2180 1486
rect 2174 1481 2180 1482
rect 2102 1475 2108 1476
rect 2102 1471 2103 1475
rect 2107 1471 2108 1475
rect 2102 1470 2108 1471
rect 2154 1475 2160 1476
rect 2154 1471 2155 1475
rect 2159 1471 2160 1475
rect 2154 1470 2160 1471
rect 2176 1467 2178 1481
rect 2236 1476 2238 1510
rect 2262 1486 2268 1487
rect 2262 1482 2263 1486
rect 2267 1482 2268 1486
rect 2262 1481 2268 1482
rect 2234 1475 2240 1476
rect 2234 1471 2235 1475
rect 2239 1471 2240 1475
rect 2234 1470 2240 1471
rect 2264 1467 2266 1481
rect 2271 1476 2275 1477
rect 2324 1476 2326 1510
rect 2350 1486 2356 1487
rect 2350 1482 2351 1486
rect 2355 1482 2356 1486
rect 2350 1481 2356 1482
rect 2271 1471 2275 1472
rect 2322 1475 2328 1476
rect 2322 1471 2323 1475
rect 2327 1471 2328 1475
rect 1871 1466 1875 1467
rect 1255 1462 1259 1463
rect 1255 1457 1259 1458
rect 1327 1462 1331 1463
rect 1327 1457 1331 1458
rect 1463 1462 1467 1463
rect 1463 1457 1467 1458
rect 1831 1462 1835 1463
rect 1871 1461 1875 1462
rect 2095 1466 2099 1467
rect 2095 1461 2099 1462
rect 2175 1466 2179 1467
rect 2175 1461 2179 1462
rect 2263 1466 2267 1467
rect 2263 1461 2267 1462
rect 1831 1457 1835 1458
rect 1256 1441 1258 1457
rect 1254 1440 1260 1441
rect 1254 1436 1255 1440
rect 1259 1436 1260 1440
rect 1832 1438 1834 1457
rect 1254 1435 1260 1436
rect 1830 1437 1836 1438
rect 1830 1433 1831 1437
rect 1835 1433 1836 1437
rect 1872 1433 1874 1461
rect 2264 1451 2266 1461
rect 2272 1460 2274 1471
rect 2322 1470 2328 1471
rect 2352 1467 2354 1481
rect 2412 1476 2414 1510
rect 2446 1486 2452 1487
rect 2446 1482 2447 1486
rect 2451 1482 2452 1486
rect 2446 1481 2452 1482
rect 2410 1475 2416 1476
rect 2410 1471 2411 1475
rect 2415 1471 2416 1475
rect 2410 1470 2416 1471
rect 2448 1467 2450 1481
rect 2508 1476 2510 1510
rect 2514 1507 2515 1511
rect 2519 1507 2520 1511
rect 2722 1511 2723 1515
rect 2727 1511 2728 1515
rect 2722 1510 2728 1511
rect 2850 1515 2856 1516
rect 2850 1511 2851 1515
rect 2855 1511 2856 1515
rect 2850 1510 2856 1511
rect 2514 1506 2520 1507
rect 2516 1477 2518 1506
rect 2542 1486 2548 1487
rect 2542 1482 2543 1486
rect 2547 1482 2548 1486
rect 2542 1481 2548 1482
rect 2654 1486 2660 1487
rect 2654 1482 2655 1486
rect 2659 1482 2660 1486
rect 2654 1481 2660 1482
rect 2663 1484 2667 1485
rect 2515 1476 2519 1477
rect 2506 1475 2512 1476
rect 2506 1471 2507 1475
rect 2511 1471 2512 1475
rect 2515 1471 2519 1472
rect 2506 1470 2512 1471
rect 2544 1467 2546 1481
rect 2656 1467 2658 1481
rect 2663 1479 2667 1480
rect 2664 1476 2666 1479
rect 2724 1476 2726 1510
rect 2790 1486 2796 1487
rect 2790 1482 2791 1486
rect 2795 1482 2796 1486
rect 2790 1481 2796 1482
rect 2662 1475 2668 1476
rect 2662 1471 2663 1475
rect 2667 1471 2668 1475
rect 2662 1470 2668 1471
rect 2722 1475 2728 1476
rect 2722 1471 2723 1475
rect 2727 1471 2728 1475
rect 2722 1470 2728 1471
rect 2792 1467 2794 1481
rect 2343 1466 2347 1467
rect 2343 1461 2347 1462
rect 2351 1466 2355 1467
rect 2351 1461 2355 1462
rect 2423 1466 2427 1467
rect 2423 1461 2427 1462
rect 2447 1466 2451 1467
rect 2447 1461 2451 1462
rect 2503 1466 2507 1467
rect 2503 1461 2507 1462
rect 2543 1466 2547 1467
rect 2543 1461 2547 1462
rect 2607 1466 2611 1467
rect 2607 1461 2611 1462
rect 2655 1466 2659 1467
rect 2655 1461 2659 1462
rect 2735 1466 2739 1467
rect 2735 1461 2739 1462
rect 2791 1466 2795 1467
rect 2791 1461 2795 1462
rect 2270 1459 2276 1460
rect 2270 1455 2271 1459
rect 2275 1455 2276 1459
rect 2270 1454 2276 1455
rect 2314 1459 2320 1460
rect 2314 1455 2315 1459
rect 2319 1455 2320 1459
rect 2314 1454 2320 1455
rect 2262 1450 2268 1451
rect 2262 1446 2263 1450
rect 2267 1446 2268 1450
rect 2262 1445 2268 1446
rect 1830 1432 1836 1433
rect 1870 1432 1876 1433
rect 786 1431 792 1432
rect 786 1427 787 1431
rect 791 1427 792 1431
rect 786 1426 792 1427
rect 898 1431 904 1432
rect 898 1427 899 1431
rect 903 1427 904 1431
rect 898 1426 904 1427
rect 1002 1431 1008 1432
rect 1002 1427 1003 1431
rect 1007 1427 1008 1431
rect 1002 1426 1008 1427
rect 1106 1431 1112 1432
rect 1106 1427 1107 1431
rect 1111 1427 1112 1431
rect 1106 1426 1112 1427
rect 1210 1431 1216 1432
rect 1210 1427 1211 1431
rect 1215 1427 1216 1431
rect 1210 1426 1216 1427
rect 1218 1431 1224 1432
rect 1218 1427 1219 1431
rect 1223 1427 1224 1431
rect 1870 1428 1871 1432
rect 1875 1428 1876 1432
rect 1870 1427 1876 1428
rect 1218 1426 1224 1427
rect 726 1402 732 1403
rect 726 1398 727 1402
rect 731 1398 732 1402
rect 726 1397 732 1398
rect 614 1391 620 1392
rect 614 1387 615 1391
rect 619 1387 620 1391
rect 614 1386 620 1387
rect 728 1371 730 1397
rect 788 1392 790 1426
rect 838 1402 844 1403
rect 838 1398 839 1402
rect 843 1398 844 1402
rect 838 1397 844 1398
rect 786 1391 792 1392
rect 786 1387 787 1391
rect 791 1387 792 1391
rect 786 1386 792 1387
rect 840 1371 842 1397
rect 900 1392 902 1426
rect 942 1402 948 1403
rect 942 1398 943 1402
rect 947 1398 948 1402
rect 942 1397 948 1398
rect 898 1391 904 1392
rect 898 1387 899 1391
rect 903 1387 904 1391
rect 898 1386 904 1387
rect 944 1371 946 1397
rect 1004 1392 1006 1426
rect 1046 1402 1052 1403
rect 1046 1398 1047 1402
rect 1051 1398 1052 1402
rect 1046 1397 1052 1398
rect 1002 1391 1008 1392
rect 1002 1387 1003 1391
rect 1007 1387 1008 1391
rect 1002 1386 1008 1387
rect 1048 1371 1050 1397
rect 1108 1392 1110 1426
rect 1150 1402 1156 1403
rect 1150 1398 1151 1402
rect 1155 1398 1156 1402
rect 1150 1397 1156 1398
rect 1106 1391 1112 1392
rect 1106 1387 1107 1391
rect 1111 1387 1112 1391
rect 1106 1386 1112 1387
rect 1152 1371 1154 1397
rect 1212 1392 1214 1426
rect 2316 1424 2318 1454
rect 2344 1451 2346 1461
rect 2394 1459 2400 1460
rect 2394 1455 2395 1459
rect 2399 1455 2400 1459
rect 2394 1454 2400 1455
rect 2342 1450 2348 1451
rect 2342 1446 2343 1450
rect 2347 1446 2348 1450
rect 2342 1445 2348 1446
rect 2396 1424 2398 1454
rect 2424 1451 2426 1461
rect 2474 1459 2480 1460
rect 2474 1455 2475 1459
rect 2479 1455 2480 1459
rect 2474 1454 2480 1455
rect 2422 1450 2428 1451
rect 2422 1446 2423 1450
rect 2427 1446 2428 1450
rect 2422 1445 2428 1446
rect 2476 1424 2478 1454
rect 2504 1451 2506 1461
rect 2608 1451 2610 1461
rect 2666 1459 2672 1460
rect 2666 1455 2667 1459
rect 2671 1455 2672 1459
rect 2666 1454 2672 1455
rect 2502 1450 2508 1451
rect 2502 1446 2503 1450
rect 2507 1446 2508 1450
rect 2502 1445 2508 1446
rect 2606 1450 2612 1451
rect 2606 1446 2607 1450
rect 2611 1446 2612 1450
rect 2606 1445 2612 1446
rect 2668 1424 2670 1454
rect 2736 1451 2738 1461
rect 2852 1460 2854 1510
rect 2936 1476 2938 1578
rect 3046 1572 3052 1573
rect 3046 1568 3047 1572
rect 3051 1568 3052 1572
rect 3046 1567 3052 1568
rect 3198 1572 3204 1573
rect 3198 1568 3199 1572
rect 3203 1568 3204 1572
rect 3198 1567 3204 1568
rect 3358 1572 3364 1573
rect 3358 1568 3359 1572
rect 3363 1568 3364 1572
rect 3358 1567 3364 1568
rect 3048 1547 3050 1567
rect 3200 1547 3202 1567
rect 3360 1547 3362 1567
rect 2943 1546 2947 1547
rect 2943 1541 2947 1542
rect 3047 1546 3051 1547
rect 3047 1541 3051 1542
rect 3119 1546 3123 1547
rect 3119 1541 3123 1542
rect 3199 1546 3203 1547
rect 3199 1541 3203 1542
rect 3303 1546 3307 1547
rect 3303 1541 3307 1542
rect 3359 1546 3363 1547
rect 3359 1541 3363 1542
rect 2944 1525 2946 1541
rect 3120 1525 3122 1541
rect 3304 1525 3306 1541
rect 2942 1524 2948 1525
rect 2942 1520 2943 1524
rect 2947 1520 2948 1524
rect 2942 1519 2948 1520
rect 3118 1524 3124 1525
rect 3118 1520 3119 1524
rect 3123 1520 3124 1524
rect 3118 1519 3124 1520
rect 3302 1524 3308 1525
rect 3302 1520 3303 1524
rect 3307 1520 3308 1524
rect 3302 1519 3308 1520
rect 3038 1515 3044 1516
rect 3038 1511 3039 1515
rect 3043 1511 3044 1515
rect 3038 1510 3044 1511
rect 3194 1515 3200 1516
rect 3194 1511 3195 1515
rect 3199 1511 3200 1515
rect 3194 1510 3200 1511
rect 3202 1515 3208 1516
rect 3202 1511 3203 1515
rect 3207 1511 3208 1515
rect 3202 1510 3208 1511
rect 2950 1486 2956 1487
rect 2950 1482 2951 1486
rect 2955 1482 2956 1486
rect 2950 1481 2956 1482
rect 2934 1475 2940 1476
rect 2934 1471 2935 1475
rect 2939 1471 2940 1475
rect 2934 1470 2940 1471
rect 2952 1467 2954 1481
rect 3040 1476 3042 1510
rect 3126 1486 3132 1487
rect 3126 1482 3127 1486
rect 3131 1482 3132 1486
rect 3126 1481 3132 1482
rect 3038 1475 3044 1476
rect 3038 1471 3039 1475
rect 3043 1471 3044 1475
rect 3038 1470 3044 1471
rect 3128 1467 3130 1481
rect 3196 1476 3198 1510
rect 3204 1485 3206 1510
rect 3310 1486 3316 1487
rect 3203 1484 3207 1485
rect 3310 1482 3311 1486
rect 3315 1482 3316 1486
rect 3310 1481 3316 1482
rect 3203 1479 3207 1480
rect 3194 1475 3200 1476
rect 3194 1471 3195 1475
rect 3199 1471 3200 1475
rect 3194 1470 3200 1471
rect 3312 1467 3314 1481
rect 2895 1466 2899 1467
rect 2895 1461 2899 1462
rect 2951 1466 2955 1467
rect 2951 1461 2955 1462
rect 3079 1466 3083 1467
rect 3079 1461 3083 1462
rect 3127 1466 3131 1467
rect 3127 1461 3131 1462
rect 3279 1466 3283 1467
rect 3279 1461 3283 1462
rect 3311 1466 3315 1467
rect 3311 1461 3315 1462
rect 3479 1466 3483 1467
rect 3479 1461 3483 1462
rect 2842 1459 2848 1460
rect 2842 1455 2843 1459
rect 2847 1455 2848 1459
rect 2842 1454 2848 1455
rect 2850 1459 2856 1460
rect 2850 1455 2851 1459
rect 2855 1455 2856 1459
rect 2850 1454 2856 1455
rect 2734 1450 2740 1451
rect 2734 1446 2735 1450
rect 2739 1446 2740 1450
rect 2734 1445 2740 1446
rect 2844 1437 2846 1454
rect 2896 1451 2898 1461
rect 3070 1459 3076 1460
rect 3070 1455 3071 1459
rect 3075 1455 3076 1459
rect 3070 1454 3076 1455
rect 2894 1450 2900 1451
rect 2894 1446 2895 1450
rect 2899 1446 2900 1450
rect 2894 1445 2900 1446
rect 2843 1436 2847 1437
rect 2843 1431 2847 1432
rect 3072 1424 3074 1454
rect 3080 1451 3082 1461
rect 3190 1459 3196 1460
rect 3190 1455 3191 1459
rect 3195 1455 3196 1459
rect 3190 1454 3196 1455
rect 3078 1450 3084 1451
rect 3078 1446 3079 1450
rect 3083 1446 3084 1450
rect 3078 1445 3084 1446
rect 3192 1424 3194 1454
rect 3280 1451 3282 1461
rect 3480 1451 3482 1461
rect 3278 1450 3284 1451
rect 3278 1446 3279 1450
rect 3283 1446 3284 1450
rect 3278 1445 3284 1446
rect 3478 1450 3484 1451
rect 3478 1446 3479 1450
rect 3483 1446 3484 1450
rect 3478 1445 3484 1446
rect 3287 1436 3291 1437
rect 3287 1431 3291 1432
rect 3288 1424 3290 1431
rect 2314 1423 2320 1424
rect 1830 1420 1836 1421
rect 1830 1416 1831 1420
rect 1835 1416 1836 1420
rect 2314 1419 2315 1423
rect 2319 1419 2320 1423
rect 2314 1418 2320 1419
rect 2394 1423 2400 1424
rect 2394 1419 2395 1423
rect 2399 1419 2400 1423
rect 2394 1418 2400 1419
rect 2474 1423 2480 1424
rect 2474 1419 2475 1423
rect 2479 1419 2480 1423
rect 2474 1418 2480 1419
rect 2666 1423 2672 1424
rect 2666 1419 2667 1423
rect 2671 1419 2672 1423
rect 2666 1418 2672 1419
rect 3070 1423 3076 1424
rect 3070 1419 3071 1423
rect 3075 1419 3076 1423
rect 3070 1418 3076 1419
rect 3190 1423 3196 1424
rect 3190 1419 3191 1423
rect 3195 1419 3196 1423
rect 3190 1418 3196 1419
rect 3286 1423 3292 1424
rect 3286 1419 3287 1423
rect 3291 1419 3292 1423
rect 3286 1418 3292 1419
rect 1830 1415 1836 1416
rect 1870 1415 1876 1416
rect 1262 1402 1268 1403
rect 1262 1398 1263 1402
rect 1267 1398 1268 1402
rect 1262 1397 1268 1398
rect 1210 1391 1216 1392
rect 1210 1387 1211 1391
rect 1215 1387 1216 1391
rect 1210 1386 1216 1387
rect 1174 1383 1180 1384
rect 1174 1379 1175 1383
rect 1179 1379 1180 1383
rect 1174 1378 1180 1379
rect 367 1370 371 1371
rect 367 1365 371 1366
rect 431 1370 435 1371
rect 431 1365 435 1366
rect 487 1370 491 1371
rect 487 1365 491 1366
rect 583 1370 587 1371
rect 583 1365 587 1366
rect 607 1370 611 1371
rect 607 1365 611 1366
rect 727 1370 731 1371
rect 727 1365 731 1366
rect 735 1370 739 1371
rect 735 1365 739 1366
rect 839 1370 843 1371
rect 839 1365 843 1366
rect 879 1370 883 1371
rect 879 1365 883 1366
rect 943 1370 947 1371
rect 943 1365 947 1366
rect 1023 1370 1027 1371
rect 1023 1365 1027 1366
rect 1047 1370 1051 1371
rect 1047 1365 1051 1366
rect 1151 1370 1155 1371
rect 1151 1365 1155 1366
rect 1167 1370 1171 1371
rect 1167 1365 1171 1366
rect 298 1363 304 1364
rect 298 1359 299 1363
rect 303 1359 304 1363
rect 298 1358 304 1359
rect 338 1363 344 1364
rect 338 1359 339 1363
rect 343 1359 344 1363
rect 338 1358 344 1359
rect 286 1354 292 1355
rect 286 1350 287 1354
rect 291 1350 292 1354
rect 286 1349 292 1350
rect 340 1328 342 1358
rect 432 1355 434 1365
rect 584 1355 586 1365
rect 634 1363 640 1364
rect 634 1359 635 1363
rect 639 1359 640 1363
rect 634 1358 640 1359
rect 430 1354 436 1355
rect 430 1350 431 1354
rect 435 1350 436 1354
rect 430 1349 436 1350
rect 582 1354 588 1355
rect 582 1350 583 1354
rect 587 1350 588 1354
rect 582 1349 588 1350
rect 636 1328 638 1358
rect 662 1355 668 1356
rect 736 1355 738 1365
rect 786 1363 792 1364
rect 786 1359 787 1363
rect 791 1359 792 1363
rect 786 1358 792 1359
rect 662 1351 663 1355
rect 667 1351 668 1355
rect 662 1350 668 1351
rect 734 1354 740 1355
rect 734 1350 735 1354
rect 739 1350 740 1354
rect 194 1327 200 1328
rect 194 1323 195 1327
rect 199 1323 200 1327
rect 194 1322 200 1323
rect 338 1327 344 1328
rect 338 1323 339 1327
rect 343 1323 344 1327
rect 338 1322 344 1323
rect 634 1327 640 1328
rect 634 1323 635 1327
rect 639 1323 640 1327
rect 634 1322 640 1323
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 110 1314 116 1315
rect 134 1316 140 1317
rect 112 1291 114 1314
rect 134 1312 135 1316
rect 139 1312 140 1316
rect 134 1311 140 1312
rect 278 1316 284 1317
rect 278 1312 279 1316
rect 283 1312 284 1316
rect 278 1311 284 1312
rect 422 1316 428 1317
rect 422 1312 423 1316
rect 427 1312 428 1316
rect 422 1311 428 1312
rect 574 1316 580 1317
rect 574 1312 575 1316
rect 579 1312 580 1316
rect 574 1311 580 1312
rect 136 1291 138 1311
rect 280 1291 282 1311
rect 424 1291 426 1311
rect 438 1299 444 1300
rect 438 1295 439 1299
rect 443 1295 444 1299
rect 438 1294 444 1295
rect 111 1290 115 1291
rect 111 1285 115 1286
rect 135 1290 139 1291
rect 135 1285 139 1286
rect 263 1290 267 1291
rect 263 1285 267 1286
rect 279 1290 283 1291
rect 279 1285 283 1286
rect 423 1290 427 1291
rect 423 1285 427 1286
rect 112 1266 114 1285
rect 136 1269 138 1285
rect 264 1269 266 1285
rect 424 1269 426 1285
rect 134 1268 140 1269
rect 110 1265 116 1266
rect 110 1261 111 1265
rect 115 1261 116 1265
rect 134 1264 135 1268
rect 139 1264 140 1268
rect 134 1263 140 1264
rect 262 1268 268 1269
rect 262 1264 263 1268
rect 267 1264 268 1268
rect 262 1263 268 1264
rect 422 1268 428 1269
rect 422 1264 423 1268
rect 427 1264 428 1268
rect 422 1263 428 1264
rect 110 1260 116 1261
rect 110 1248 116 1249
rect 110 1244 111 1248
rect 115 1244 116 1248
rect 110 1243 116 1244
rect 112 1207 114 1243
rect 142 1230 148 1231
rect 142 1226 143 1230
rect 147 1226 148 1230
rect 142 1225 148 1226
rect 270 1230 276 1231
rect 270 1226 271 1230
rect 275 1226 276 1230
rect 270 1225 276 1226
rect 430 1230 436 1231
rect 430 1226 431 1230
rect 435 1226 436 1230
rect 430 1225 436 1226
rect 144 1207 146 1225
rect 194 1219 200 1220
rect 194 1215 195 1219
rect 199 1215 200 1219
rect 194 1214 200 1215
rect 111 1206 115 1207
rect 111 1201 115 1202
rect 143 1206 147 1207
rect 143 1201 147 1202
rect 112 1173 114 1201
rect 144 1191 146 1201
rect 142 1190 148 1191
rect 142 1186 143 1190
rect 147 1186 148 1190
rect 142 1185 148 1186
rect 110 1172 116 1173
rect 110 1168 111 1172
rect 115 1168 116 1172
rect 110 1167 116 1168
rect 196 1164 198 1214
rect 272 1207 274 1225
rect 432 1207 434 1225
rect 440 1220 442 1294
rect 576 1291 578 1311
rect 575 1290 579 1291
rect 575 1285 579 1286
rect 591 1290 595 1291
rect 591 1285 595 1286
rect 592 1269 594 1285
rect 590 1268 596 1269
rect 590 1264 591 1268
rect 595 1264 596 1268
rect 590 1263 596 1264
rect 664 1260 666 1350
rect 734 1349 740 1350
rect 788 1328 790 1358
rect 880 1355 882 1365
rect 930 1363 936 1364
rect 930 1359 931 1363
rect 935 1359 936 1363
rect 930 1358 936 1359
rect 878 1354 884 1355
rect 878 1350 879 1354
rect 883 1350 884 1354
rect 878 1349 884 1350
rect 932 1328 934 1358
rect 1024 1355 1026 1365
rect 1074 1363 1080 1364
rect 1074 1359 1075 1363
rect 1079 1359 1080 1363
rect 1074 1358 1080 1359
rect 1022 1354 1028 1355
rect 1022 1350 1023 1354
rect 1027 1350 1028 1354
rect 1022 1349 1028 1350
rect 1076 1328 1078 1358
rect 1168 1355 1170 1365
rect 1166 1354 1172 1355
rect 1166 1350 1167 1354
rect 1171 1350 1172 1354
rect 1166 1349 1172 1350
rect 1176 1328 1178 1378
rect 1264 1371 1266 1397
rect 1832 1371 1834 1415
rect 1870 1411 1871 1415
rect 1875 1411 1876 1415
rect 1870 1410 1876 1411
rect 2254 1412 2260 1413
rect 1872 1391 1874 1410
rect 2254 1408 2255 1412
rect 2259 1408 2260 1412
rect 2254 1407 2260 1408
rect 2334 1412 2340 1413
rect 2334 1408 2335 1412
rect 2339 1408 2340 1412
rect 2334 1407 2340 1408
rect 2414 1412 2420 1413
rect 2414 1408 2415 1412
rect 2419 1408 2420 1412
rect 2414 1407 2420 1408
rect 2494 1412 2500 1413
rect 2494 1408 2495 1412
rect 2499 1408 2500 1412
rect 2494 1407 2500 1408
rect 2598 1412 2604 1413
rect 2598 1408 2599 1412
rect 2603 1408 2604 1412
rect 2598 1407 2604 1408
rect 2726 1412 2732 1413
rect 2726 1408 2727 1412
rect 2731 1408 2732 1412
rect 2726 1407 2732 1408
rect 2886 1412 2892 1413
rect 2886 1408 2887 1412
rect 2891 1408 2892 1412
rect 2886 1407 2892 1408
rect 3070 1412 3076 1413
rect 3070 1408 3071 1412
rect 3075 1408 3076 1412
rect 3070 1407 3076 1408
rect 3270 1412 3276 1413
rect 3270 1408 3271 1412
rect 3275 1408 3276 1412
rect 3270 1407 3276 1408
rect 3470 1412 3476 1413
rect 3470 1408 3471 1412
rect 3475 1408 3476 1412
rect 3470 1407 3476 1408
rect 2256 1391 2258 1407
rect 2336 1391 2338 1407
rect 2416 1391 2418 1407
rect 2496 1391 2498 1407
rect 2600 1391 2602 1407
rect 2606 1395 2612 1396
rect 2606 1391 2607 1395
rect 2611 1391 2612 1395
rect 2728 1391 2730 1407
rect 2888 1391 2890 1407
rect 3072 1391 3074 1407
rect 3272 1391 3274 1407
rect 3414 1395 3420 1396
rect 3414 1391 3415 1395
rect 3419 1391 3420 1395
rect 3472 1391 3474 1407
rect 1871 1390 1875 1391
rect 1871 1385 1875 1386
rect 2255 1390 2259 1391
rect 2255 1385 2259 1386
rect 2263 1390 2267 1391
rect 2263 1385 2267 1386
rect 2335 1390 2339 1391
rect 2335 1385 2339 1386
rect 2343 1390 2347 1391
rect 2343 1385 2347 1386
rect 2415 1390 2419 1391
rect 2415 1385 2419 1386
rect 2423 1390 2427 1391
rect 2423 1385 2427 1386
rect 2495 1390 2499 1391
rect 2495 1385 2499 1386
rect 2503 1390 2507 1391
rect 2503 1385 2507 1386
rect 2591 1390 2595 1391
rect 2591 1385 2595 1386
rect 2599 1390 2603 1391
rect 2606 1390 2612 1391
rect 2695 1390 2699 1391
rect 2599 1385 2603 1386
rect 1263 1370 1267 1371
rect 1263 1365 1267 1366
rect 1319 1370 1323 1371
rect 1319 1365 1323 1366
rect 1471 1370 1475 1371
rect 1471 1365 1475 1366
rect 1623 1370 1627 1371
rect 1623 1365 1627 1366
rect 1831 1370 1835 1371
rect 1872 1366 1874 1385
rect 2264 1369 2266 1385
rect 2344 1369 2346 1385
rect 2424 1369 2426 1385
rect 2504 1369 2506 1385
rect 2592 1369 2594 1385
rect 2262 1368 2268 1369
rect 1831 1365 1835 1366
rect 1870 1365 1876 1366
rect 1320 1355 1322 1365
rect 1472 1355 1474 1365
rect 1550 1363 1556 1364
rect 1550 1359 1551 1363
rect 1555 1359 1556 1363
rect 1550 1358 1556 1359
rect 1318 1354 1324 1355
rect 1318 1350 1319 1354
rect 1323 1350 1324 1354
rect 1318 1349 1324 1350
rect 1470 1354 1476 1355
rect 1470 1350 1471 1354
rect 1475 1350 1476 1354
rect 1470 1349 1476 1350
rect 1552 1328 1554 1358
rect 1624 1355 1626 1365
rect 1622 1354 1628 1355
rect 1622 1350 1623 1354
rect 1627 1350 1628 1354
rect 1622 1349 1628 1350
rect 1832 1337 1834 1365
rect 1870 1361 1871 1365
rect 1875 1361 1876 1365
rect 2262 1364 2263 1368
rect 2267 1364 2268 1368
rect 2262 1363 2268 1364
rect 2342 1368 2348 1369
rect 2342 1364 2343 1368
rect 2347 1364 2348 1368
rect 2342 1363 2348 1364
rect 2422 1368 2428 1369
rect 2422 1364 2423 1368
rect 2427 1364 2428 1368
rect 2422 1363 2428 1364
rect 2502 1368 2508 1369
rect 2502 1364 2503 1368
rect 2507 1364 2508 1368
rect 2502 1363 2508 1364
rect 2590 1368 2596 1369
rect 2590 1364 2591 1368
rect 2595 1364 2596 1368
rect 2590 1363 2596 1364
rect 1870 1360 1876 1361
rect 2330 1359 2336 1360
rect 2330 1355 2331 1359
rect 2335 1355 2336 1359
rect 2330 1354 2336 1355
rect 2414 1359 2420 1360
rect 2414 1355 2415 1359
rect 2419 1355 2420 1359
rect 2582 1359 2588 1360
rect 2414 1354 2420 1355
rect 2422 1355 2428 1356
rect 1870 1348 1876 1349
rect 1870 1344 1871 1348
rect 1875 1344 1876 1348
rect 1870 1343 1876 1344
rect 1830 1336 1836 1337
rect 1830 1332 1831 1336
rect 1835 1332 1836 1336
rect 1830 1331 1836 1332
rect 786 1327 792 1328
rect 786 1323 787 1327
rect 791 1323 792 1327
rect 786 1322 792 1323
rect 930 1327 936 1328
rect 930 1323 931 1327
rect 935 1323 936 1327
rect 930 1322 936 1323
rect 1074 1327 1080 1328
rect 1074 1323 1075 1327
rect 1079 1323 1080 1327
rect 1074 1322 1080 1323
rect 1174 1327 1180 1328
rect 1174 1323 1175 1327
rect 1179 1323 1180 1327
rect 1174 1322 1180 1323
rect 1342 1327 1348 1328
rect 1342 1323 1343 1327
rect 1347 1323 1348 1327
rect 1342 1322 1348 1323
rect 1550 1327 1556 1328
rect 1550 1323 1551 1327
rect 1555 1323 1556 1327
rect 1550 1322 1556 1323
rect 726 1316 732 1317
rect 726 1312 727 1316
rect 731 1312 732 1316
rect 726 1311 732 1312
rect 870 1316 876 1317
rect 870 1312 871 1316
rect 875 1312 876 1316
rect 870 1311 876 1312
rect 1014 1316 1020 1317
rect 1014 1312 1015 1316
rect 1019 1312 1020 1316
rect 1014 1311 1020 1312
rect 1158 1316 1164 1317
rect 1158 1312 1159 1316
rect 1163 1312 1164 1316
rect 1158 1311 1164 1312
rect 1310 1316 1316 1317
rect 1310 1312 1311 1316
rect 1315 1312 1316 1316
rect 1310 1311 1316 1312
rect 728 1291 730 1311
rect 872 1291 874 1311
rect 1016 1291 1018 1311
rect 1160 1291 1162 1311
rect 1312 1291 1314 1311
rect 727 1290 731 1291
rect 727 1285 731 1286
rect 759 1290 763 1291
rect 759 1285 763 1286
rect 871 1290 875 1291
rect 871 1285 875 1286
rect 927 1290 931 1291
rect 927 1285 931 1286
rect 1015 1290 1019 1291
rect 1015 1285 1019 1286
rect 1079 1290 1083 1291
rect 1079 1285 1083 1286
rect 1159 1290 1163 1291
rect 1159 1285 1163 1286
rect 1223 1290 1227 1291
rect 1223 1285 1227 1286
rect 1311 1290 1315 1291
rect 1311 1285 1315 1286
rect 760 1269 762 1285
rect 928 1269 930 1285
rect 1080 1269 1082 1285
rect 1224 1269 1226 1285
rect 758 1268 764 1269
rect 758 1264 759 1268
rect 763 1264 764 1268
rect 758 1263 764 1264
rect 926 1268 932 1269
rect 926 1264 927 1268
rect 931 1264 932 1268
rect 926 1263 932 1264
rect 1078 1268 1084 1269
rect 1078 1264 1079 1268
rect 1083 1264 1084 1268
rect 1078 1263 1084 1264
rect 1222 1268 1228 1269
rect 1222 1264 1223 1268
rect 1227 1264 1228 1268
rect 1222 1263 1228 1264
rect 498 1259 504 1260
rect 498 1255 499 1259
rect 503 1255 504 1259
rect 498 1254 504 1255
rect 506 1259 512 1260
rect 506 1255 507 1259
rect 511 1255 512 1259
rect 506 1254 512 1255
rect 662 1259 668 1260
rect 662 1255 663 1259
rect 667 1255 668 1259
rect 662 1254 668 1255
rect 826 1259 832 1260
rect 826 1255 827 1259
rect 831 1255 832 1259
rect 826 1254 832 1255
rect 1158 1259 1164 1260
rect 1158 1255 1159 1259
rect 1163 1255 1164 1259
rect 1158 1254 1164 1255
rect 1290 1259 1296 1260
rect 1290 1255 1291 1259
rect 1295 1255 1296 1259
rect 1290 1254 1296 1255
rect 500 1220 502 1254
rect 438 1219 444 1220
rect 438 1215 439 1219
rect 443 1215 444 1219
rect 438 1214 444 1215
rect 498 1219 504 1220
rect 498 1215 499 1219
rect 503 1215 504 1219
rect 498 1214 504 1215
rect 271 1206 275 1207
rect 271 1201 275 1202
rect 311 1206 315 1207
rect 311 1201 315 1202
rect 431 1206 435 1207
rect 431 1201 435 1202
rect 487 1206 491 1207
rect 487 1201 491 1202
rect 312 1191 314 1201
rect 422 1199 428 1200
rect 422 1194 423 1199
rect 427 1194 428 1199
rect 423 1191 427 1192
rect 488 1191 490 1201
rect 508 1200 510 1254
rect 598 1230 604 1231
rect 598 1226 599 1230
rect 603 1226 604 1230
rect 598 1225 604 1226
rect 766 1230 772 1231
rect 766 1226 767 1230
rect 771 1226 772 1230
rect 766 1225 772 1226
rect 600 1207 602 1225
rect 768 1207 770 1225
rect 828 1220 830 1254
rect 934 1230 940 1231
rect 934 1226 935 1230
rect 939 1226 940 1230
rect 934 1225 940 1226
rect 1086 1230 1092 1231
rect 1086 1226 1087 1230
rect 1091 1226 1092 1230
rect 1086 1225 1092 1226
rect 1095 1228 1099 1229
rect 826 1219 832 1220
rect 826 1215 827 1219
rect 831 1215 832 1219
rect 826 1214 832 1215
rect 898 1219 904 1220
rect 898 1215 899 1219
rect 903 1215 904 1219
rect 898 1214 904 1215
rect 599 1206 603 1207
rect 599 1201 603 1202
rect 671 1206 675 1207
rect 671 1201 675 1202
rect 767 1206 771 1207
rect 767 1201 771 1202
rect 847 1206 851 1207
rect 847 1201 851 1202
rect 506 1199 512 1200
rect 506 1195 507 1199
rect 511 1195 512 1199
rect 506 1194 512 1195
rect 538 1199 544 1200
rect 538 1195 539 1199
rect 543 1195 544 1199
rect 538 1194 544 1195
rect 310 1190 316 1191
rect 310 1186 311 1190
rect 315 1186 316 1190
rect 310 1185 316 1186
rect 486 1190 492 1191
rect 486 1186 487 1190
rect 491 1186 492 1190
rect 486 1185 492 1186
rect 540 1164 542 1194
rect 672 1191 674 1201
rect 679 1196 683 1197
rect 679 1191 683 1192
rect 848 1191 850 1201
rect 854 1199 860 1200
rect 854 1195 855 1199
rect 859 1195 860 1199
rect 854 1194 860 1195
rect 670 1190 676 1191
rect 670 1186 671 1190
rect 675 1186 676 1190
rect 670 1185 676 1186
rect 680 1164 682 1191
rect 846 1190 852 1191
rect 846 1186 847 1190
rect 851 1186 852 1190
rect 846 1185 852 1186
rect 194 1163 200 1164
rect 194 1159 195 1163
rect 199 1159 200 1163
rect 194 1158 200 1159
rect 538 1163 544 1164
rect 538 1159 539 1163
rect 543 1159 544 1163
rect 538 1158 544 1159
rect 678 1163 684 1164
rect 678 1159 679 1163
rect 683 1159 684 1163
rect 678 1158 684 1159
rect 110 1155 116 1156
rect 110 1151 111 1155
rect 115 1151 116 1155
rect 110 1150 116 1151
rect 134 1152 140 1153
rect 112 1131 114 1150
rect 134 1148 135 1152
rect 139 1148 140 1152
rect 134 1147 140 1148
rect 302 1152 308 1153
rect 302 1148 303 1152
rect 307 1148 308 1152
rect 302 1147 308 1148
rect 478 1152 484 1153
rect 478 1148 479 1152
rect 483 1148 484 1152
rect 478 1147 484 1148
rect 662 1152 668 1153
rect 662 1148 663 1152
rect 667 1148 668 1152
rect 662 1147 668 1148
rect 838 1152 844 1153
rect 838 1148 839 1152
rect 843 1148 844 1152
rect 838 1147 844 1148
rect 136 1131 138 1147
rect 262 1135 268 1136
rect 262 1131 263 1135
rect 267 1131 268 1135
rect 304 1131 306 1147
rect 480 1131 482 1147
rect 664 1131 666 1147
rect 840 1131 842 1147
rect 111 1130 115 1131
rect 111 1125 115 1126
rect 135 1130 139 1131
rect 135 1125 139 1126
rect 247 1130 251 1131
rect 262 1130 268 1131
rect 303 1130 307 1131
rect 247 1125 251 1126
rect 112 1106 114 1125
rect 136 1109 138 1125
rect 248 1109 250 1125
rect 134 1108 140 1109
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 134 1104 135 1108
rect 139 1104 140 1108
rect 134 1103 140 1104
rect 246 1108 252 1109
rect 246 1104 247 1108
rect 251 1104 252 1108
rect 246 1103 252 1104
rect 110 1100 116 1101
rect 110 1088 116 1089
rect 110 1084 111 1088
rect 115 1084 116 1088
rect 110 1083 116 1084
rect 112 1043 114 1083
rect 142 1070 148 1071
rect 142 1066 143 1070
rect 147 1066 148 1070
rect 142 1065 148 1066
rect 254 1070 260 1071
rect 254 1066 255 1070
rect 259 1066 260 1070
rect 254 1065 260 1066
rect 144 1043 146 1065
rect 150 1059 156 1060
rect 150 1055 151 1059
rect 155 1055 156 1059
rect 150 1054 156 1055
rect 111 1042 115 1043
rect 111 1037 115 1038
rect 143 1042 147 1043
rect 143 1037 147 1038
rect 112 1009 114 1037
rect 144 1027 146 1037
rect 142 1026 148 1027
rect 142 1022 143 1026
rect 147 1022 148 1026
rect 142 1021 148 1022
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 152 1000 154 1054
rect 256 1043 258 1065
rect 264 1060 266 1130
rect 303 1125 307 1126
rect 383 1130 387 1131
rect 383 1125 387 1126
rect 479 1130 483 1131
rect 479 1125 483 1126
rect 519 1130 523 1131
rect 519 1125 523 1126
rect 647 1130 651 1131
rect 647 1125 651 1126
rect 663 1130 667 1131
rect 663 1125 667 1126
rect 775 1130 779 1131
rect 775 1125 779 1126
rect 839 1130 843 1131
rect 839 1125 843 1126
rect 384 1109 386 1125
rect 520 1109 522 1125
rect 648 1109 650 1125
rect 776 1109 778 1125
rect 382 1108 388 1109
rect 382 1104 383 1108
rect 387 1104 388 1108
rect 382 1103 388 1104
rect 518 1108 524 1109
rect 518 1104 519 1108
rect 523 1104 524 1108
rect 518 1103 524 1104
rect 646 1108 652 1109
rect 646 1104 647 1108
rect 651 1104 652 1108
rect 646 1103 652 1104
rect 774 1108 780 1109
rect 774 1104 775 1108
rect 779 1104 780 1108
rect 774 1103 780 1104
rect 856 1100 858 1194
rect 900 1164 902 1214
rect 936 1207 938 1225
rect 1088 1207 1090 1225
rect 1095 1223 1099 1224
rect 1096 1220 1098 1223
rect 1160 1220 1162 1254
rect 1282 1251 1288 1252
rect 1282 1247 1283 1251
rect 1287 1247 1288 1251
rect 1282 1246 1288 1247
rect 1230 1230 1236 1231
rect 1230 1226 1231 1230
rect 1235 1226 1236 1230
rect 1230 1225 1236 1226
rect 1094 1219 1100 1220
rect 1094 1215 1095 1219
rect 1099 1215 1100 1219
rect 1094 1214 1100 1215
rect 1158 1219 1164 1220
rect 1158 1215 1159 1219
rect 1163 1215 1164 1219
rect 1158 1214 1164 1215
rect 1232 1207 1234 1225
rect 935 1206 939 1207
rect 935 1201 939 1202
rect 1007 1206 1011 1207
rect 1007 1201 1011 1202
rect 1087 1206 1091 1207
rect 1087 1201 1091 1202
rect 1159 1206 1163 1207
rect 1159 1201 1163 1202
rect 1231 1206 1235 1207
rect 1231 1201 1235 1202
rect 1008 1191 1010 1201
rect 1058 1199 1064 1200
rect 1058 1195 1059 1199
rect 1063 1195 1064 1199
rect 1058 1194 1064 1195
rect 1006 1190 1012 1191
rect 1006 1186 1007 1190
rect 1011 1186 1012 1190
rect 1006 1185 1012 1186
rect 1060 1164 1062 1194
rect 1160 1191 1162 1201
rect 1284 1200 1286 1246
rect 1292 1229 1294 1254
rect 1291 1228 1295 1229
rect 1291 1223 1295 1224
rect 1344 1220 1346 1322
rect 1830 1319 1836 1320
rect 1462 1316 1468 1317
rect 1462 1312 1463 1316
rect 1467 1312 1468 1316
rect 1462 1311 1468 1312
rect 1614 1316 1620 1317
rect 1614 1312 1615 1316
rect 1619 1312 1620 1316
rect 1830 1315 1831 1319
rect 1835 1315 1836 1319
rect 1830 1314 1836 1315
rect 1614 1311 1620 1312
rect 1464 1291 1466 1311
rect 1616 1291 1618 1311
rect 1832 1291 1834 1314
rect 1872 1303 1874 1343
rect 2322 1339 2328 1340
rect 2322 1335 2323 1339
rect 2327 1335 2328 1339
rect 2322 1334 2328 1335
rect 2270 1330 2276 1331
rect 2270 1326 2271 1330
rect 2275 1326 2276 1330
rect 2270 1325 2276 1326
rect 2272 1303 2274 1325
rect 2324 1320 2326 1334
rect 2332 1320 2334 1354
rect 2350 1330 2356 1331
rect 2350 1326 2351 1330
rect 2355 1326 2356 1330
rect 2350 1325 2356 1326
rect 2322 1319 2328 1320
rect 2322 1315 2323 1319
rect 2327 1315 2328 1319
rect 2322 1314 2328 1315
rect 2330 1319 2336 1320
rect 2330 1315 2331 1319
rect 2335 1315 2336 1319
rect 2330 1314 2336 1315
rect 2352 1303 2354 1325
rect 2416 1312 2418 1354
rect 2422 1351 2423 1355
rect 2427 1351 2428 1355
rect 2582 1355 2583 1359
rect 2587 1355 2588 1359
rect 2582 1354 2588 1355
rect 2422 1350 2428 1351
rect 2414 1311 2420 1312
rect 2414 1307 2415 1311
rect 2419 1307 2420 1311
rect 2414 1306 2420 1307
rect 1871 1302 1875 1303
rect 1871 1297 1875 1298
rect 2215 1302 2219 1303
rect 2215 1297 2219 1298
rect 2271 1302 2275 1303
rect 2271 1297 2275 1298
rect 2295 1302 2299 1303
rect 2295 1297 2299 1298
rect 2351 1302 2355 1303
rect 2351 1297 2355 1298
rect 2375 1302 2379 1303
rect 2375 1297 2379 1298
rect 1351 1290 1355 1291
rect 1351 1285 1355 1286
rect 1463 1290 1467 1291
rect 1463 1285 1467 1286
rect 1479 1290 1483 1291
rect 1479 1285 1483 1286
rect 1607 1290 1611 1291
rect 1607 1285 1611 1286
rect 1615 1290 1619 1291
rect 1615 1285 1619 1286
rect 1735 1290 1739 1291
rect 1735 1285 1739 1286
rect 1831 1290 1835 1291
rect 1831 1285 1835 1286
rect 1352 1269 1354 1285
rect 1480 1269 1482 1285
rect 1608 1269 1610 1285
rect 1736 1269 1738 1285
rect 1350 1268 1356 1269
rect 1350 1264 1351 1268
rect 1355 1264 1356 1268
rect 1350 1263 1356 1264
rect 1478 1268 1484 1269
rect 1478 1264 1479 1268
rect 1483 1264 1484 1268
rect 1478 1263 1484 1264
rect 1606 1268 1612 1269
rect 1606 1264 1607 1268
rect 1611 1264 1612 1268
rect 1606 1263 1612 1264
rect 1734 1268 1740 1269
rect 1734 1264 1735 1268
rect 1739 1264 1740 1268
rect 1832 1266 1834 1285
rect 1872 1269 1874 1297
rect 2216 1287 2218 1297
rect 2278 1295 2284 1296
rect 2278 1291 2279 1295
rect 2283 1291 2284 1295
rect 2278 1290 2284 1291
rect 2214 1286 2220 1287
rect 2214 1282 2215 1286
rect 2219 1282 2220 1286
rect 2214 1281 2220 1282
rect 1870 1268 1876 1269
rect 1734 1263 1740 1264
rect 1830 1265 1836 1266
rect 1830 1261 1831 1265
rect 1835 1261 1836 1265
rect 1870 1264 1871 1268
rect 1875 1264 1876 1268
rect 1870 1263 1876 1264
rect 1830 1260 1836 1261
rect 2280 1260 2282 1290
rect 2296 1287 2298 1297
rect 2358 1295 2364 1296
rect 2358 1291 2359 1295
rect 2363 1291 2364 1295
rect 2358 1290 2364 1291
rect 2294 1286 2300 1287
rect 2294 1282 2295 1286
rect 2299 1282 2300 1286
rect 2294 1281 2300 1282
rect 2360 1260 2362 1290
rect 2376 1287 2378 1297
rect 2424 1296 2426 1350
rect 2584 1341 2586 1354
rect 2583 1340 2587 1341
rect 2583 1335 2587 1336
rect 2430 1330 2436 1331
rect 2430 1326 2431 1330
rect 2435 1326 2436 1330
rect 2430 1325 2436 1326
rect 2510 1330 2516 1331
rect 2510 1326 2511 1330
rect 2515 1326 2516 1330
rect 2510 1325 2516 1326
rect 2598 1330 2604 1331
rect 2598 1326 2599 1330
rect 2603 1326 2604 1330
rect 2598 1325 2604 1326
rect 2432 1303 2434 1325
rect 2512 1303 2514 1325
rect 2600 1303 2602 1325
rect 2608 1320 2610 1390
rect 2695 1385 2699 1386
rect 2727 1390 2731 1391
rect 2727 1385 2731 1386
rect 2807 1390 2811 1391
rect 2807 1385 2811 1386
rect 2887 1390 2891 1391
rect 2887 1385 2891 1386
rect 2919 1390 2923 1391
rect 2919 1385 2923 1386
rect 3039 1390 3043 1391
rect 3039 1385 3043 1386
rect 3071 1390 3075 1391
rect 3071 1385 3075 1386
rect 3159 1390 3163 1391
rect 3159 1385 3163 1386
rect 3271 1390 3275 1391
rect 3271 1385 3275 1386
rect 3279 1390 3283 1391
rect 3279 1385 3283 1386
rect 3399 1390 3403 1391
rect 3414 1390 3420 1391
rect 3471 1390 3475 1391
rect 3399 1385 3403 1386
rect 2696 1369 2698 1385
rect 2808 1369 2810 1385
rect 2920 1369 2922 1385
rect 3040 1369 3042 1385
rect 3160 1369 3162 1385
rect 3280 1369 3282 1385
rect 3400 1369 3402 1385
rect 2694 1368 2700 1369
rect 2694 1364 2695 1368
rect 2699 1364 2700 1368
rect 2694 1363 2700 1364
rect 2806 1368 2812 1369
rect 2806 1364 2807 1368
rect 2811 1364 2812 1368
rect 2806 1363 2812 1364
rect 2918 1368 2924 1369
rect 2918 1364 2919 1368
rect 2923 1364 2924 1368
rect 2918 1363 2924 1364
rect 3038 1368 3044 1369
rect 3038 1364 3039 1368
rect 3043 1364 3044 1368
rect 3038 1363 3044 1364
rect 3158 1368 3164 1369
rect 3158 1364 3159 1368
rect 3163 1364 3164 1368
rect 3158 1363 3164 1364
rect 3278 1368 3284 1369
rect 3278 1364 3279 1368
rect 3283 1364 3284 1368
rect 3278 1363 3284 1364
rect 3398 1368 3404 1369
rect 3398 1364 3399 1368
rect 3403 1364 3404 1368
rect 3398 1363 3404 1364
rect 2658 1359 2664 1360
rect 2658 1355 2659 1359
rect 2663 1355 2664 1359
rect 2658 1354 2664 1355
rect 2762 1359 2768 1360
rect 2762 1355 2763 1359
rect 2767 1355 2768 1359
rect 2762 1354 2768 1355
rect 2770 1359 2776 1360
rect 2770 1355 2771 1359
rect 2775 1355 2776 1359
rect 2770 1354 2776 1355
rect 2986 1359 2992 1360
rect 2986 1355 2987 1359
rect 2991 1355 2992 1359
rect 3226 1359 3232 1360
rect 2986 1354 2992 1355
rect 3038 1355 3044 1356
rect 2660 1320 2662 1354
rect 2702 1330 2708 1331
rect 2702 1326 2703 1330
rect 2707 1326 2708 1330
rect 2702 1325 2708 1326
rect 2606 1319 2612 1320
rect 2606 1315 2607 1319
rect 2611 1315 2612 1319
rect 2606 1314 2612 1315
rect 2658 1319 2664 1320
rect 2658 1315 2659 1319
rect 2663 1315 2664 1319
rect 2658 1314 2664 1315
rect 2670 1303 2676 1304
rect 2704 1303 2706 1325
rect 2764 1320 2766 1354
rect 2772 1340 2774 1354
rect 2839 1340 2843 1341
rect 2770 1339 2776 1340
rect 2770 1335 2771 1339
rect 2775 1335 2776 1339
rect 2839 1335 2843 1336
rect 2770 1334 2776 1335
rect 2814 1330 2820 1331
rect 2814 1326 2815 1330
rect 2819 1326 2820 1330
rect 2814 1325 2820 1326
rect 2762 1319 2768 1320
rect 2762 1315 2763 1319
rect 2767 1315 2768 1319
rect 2762 1314 2768 1315
rect 2816 1303 2818 1325
rect 2840 1320 2842 1335
rect 2926 1330 2932 1331
rect 2926 1326 2927 1330
rect 2931 1326 2932 1330
rect 2926 1325 2932 1326
rect 2838 1319 2844 1320
rect 2838 1315 2839 1319
rect 2843 1315 2844 1319
rect 2838 1314 2844 1315
rect 2928 1303 2930 1325
rect 2988 1320 2990 1354
rect 3038 1351 3039 1355
rect 3043 1351 3044 1355
rect 3226 1355 3227 1359
rect 3231 1355 3232 1359
rect 3226 1354 3232 1355
rect 3234 1359 3240 1360
rect 3234 1355 3235 1359
rect 3239 1355 3240 1359
rect 3234 1354 3240 1355
rect 3346 1359 3352 1360
rect 3346 1355 3347 1359
rect 3351 1355 3352 1359
rect 3346 1354 3352 1355
rect 3038 1350 3044 1351
rect 2986 1319 2992 1320
rect 2986 1315 2987 1319
rect 2991 1315 2992 1319
rect 2986 1314 2992 1315
rect 2431 1302 2435 1303
rect 2431 1297 2435 1298
rect 2455 1302 2459 1303
rect 2455 1297 2459 1298
rect 2511 1302 2515 1303
rect 2511 1297 2515 1298
rect 2551 1302 2555 1303
rect 2551 1297 2555 1298
rect 2599 1302 2603 1303
rect 2599 1297 2603 1298
rect 2663 1302 2667 1303
rect 2670 1299 2671 1303
rect 2675 1299 2676 1303
rect 2670 1298 2676 1299
rect 2703 1302 2707 1303
rect 2663 1297 2667 1298
rect 2422 1295 2428 1296
rect 2422 1291 2423 1295
rect 2427 1291 2428 1295
rect 2422 1290 2428 1291
rect 2456 1287 2458 1297
rect 2552 1287 2554 1297
rect 2654 1295 2660 1296
rect 2654 1291 2655 1295
rect 2659 1291 2660 1295
rect 2654 1290 2660 1291
rect 2374 1286 2380 1287
rect 2374 1282 2375 1286
rect 2379 1282 2380 1286
rect 2374 1281 2380 1282
rect 2454 1286 2460 1287
rect 2454 1282 2455 1286
rect 2459 1282 2460 1286
rect 2454 1281 2460 1282
rect 2550 1286 2556 1287
rect 2550 1282 2551 1286
rect 2555 1282 2556 1286
rect 2550 1281 2556 1282
rect 2656 1260 2658 1290
rect 2664 1287 2666 1297
rect 2662 1286 2668 1287
rect 2662 1282 2663 1286
rect 2667 1282 2668 1286
rect 2662 1281 2668 1282
rect 2672 1260 2674 1298
rect 2703 1297 2707 1298
rect 2791 1302 2795 1303
rect 2791 1297 2795 1298
rect 2815 1302 2819 1303
rect 2815 1297 2819 1298
rect 2927 1302 2931 1303
rect 2927 1297 2931 1298
rect 2792 1287 2794 1297
rect 2850 1295 2856 1296
rect 2850 1291 2851 1295
rect 2855 1291 2856 1295
rect 2850 1290 2856 1291
rect 2790 1286 2796 1287
rect 2790 1282 2791 1286
rect 2795 1282 2796 1286
rect 2790 1281 2796 1282
rect 2852 1260 2854 1290
rect 2928 1287 2930 1297
rect 3040 1296 3042 1350
rect 3046 1330 3052 1331
rect 3046 1326 3047 1330
rect 3051 1326 3052 1330
rect 3046 1325 3052 1326
rect 3166 1330 3172 1331
rect 3166 1326 3167 1330
rect 3171 1326 3172 1330
rect 3166 1325 3172 1326
rect 3048 1303 3050 1325
rect 3168 1303 3170 1325
rect 3047 1302 3051 1303
rect 3047 1297 3051 1298
rect 3071 1302 3075 1303
rect 3071 1297 3075 1298
rect 3167 1302 3171 1303
rect 3167 1297 3171 1298
rect 3215 1302 3219 1303
rect 3215 1297 3219 1298
rect 2998 1295 3004 1296
rect 2998 1291 2999 1295
rect 3003 1291 3004 1295
rect 2998 1290 3004 1291
rect 3038 1295 3044 1296
rect 3038 1291 3039 1295
rect 3043 1291 3044 1295
rect 3038 1290 3044 1291
rect 2926 1286 2932 1287
rect 2926 1282 2927 1286
rect 2931 1282 2932 1286
rect 2926 1281 2932 1282
rect 3000 1260 3002 1290
rect 3072 1287 3074 1297
rect 3216 1287 3218 1297
rect 3228 1296 3230 1354
rect 3236 1320 3238 1354
rect 3286 1330 3292 1331
rect 3286 1326 3287 1330
rect 3291 1326 3292 1330
rect 3286 1325 3292 1326
rect 3234 1319 3240 1320
rect 3234 1315 3235 1319
rect 3239 1315 3240 1319
rect 3234 1314 3240 1315
rect 3288 1303 3290 1325
rect 3348 1320 3350 1354
rect 3406 1330 3412 1331
rect 3406 1326 3407 1330
rect 3411 1326 3412 1330
rect 3406 1325 3412 1326
rect 3346 1319 3352 1320
rect 3346 1315 3347 1319
rect 3351 1315 3352 1319
rect 3346 1314 3352 1315
rect 3408 1303 3410 1325
rect 3416 1320 3418 1390
rect 3471 1385 3475 1386
rect 3488 1360 3490 1614
rect 3512 1611 3514 1621
rect 3510 1610 3516 1611
rect 3510 1606 3511 1610
rect 3515 1606 3516 1610
rect 3510 1605 3516 1606
rect 3528 1584 3530 1798
rect 3592 1787 3594 1827
rect 3591 1786 3595 1787
rect 3591 1781 3595 1782
rect 3592 1753 3594 1781
rect 3590 1752 3596 1753
rect 3590 1748 3591 1752
rect 3595 1748 3596 1752
rect 3590 1747 3596 1748
rect 3590 1735 3596 1736
rect 3590 1731 3591 1735
rect 3595 1731 3596 1735
rect 3590 1730 3596 1731
rect 3592 1707 3594 1730
rect 3591 1706 3595 1707
rect 3591 1701 3595 1702
rect 3592 1682 3594 1701
rect 3590 1681 3596 1682
rect 3590 1677 3591 1681
rect 3595 1677 3596 1681
rect 3590 1676 3596 1677
rect 3590 1664 3596 1665
rect 3590 1660 3591 1664
rect 3595 1660 3596 1664
rect 3590 1659 3596 1660
rect 3592 1627 3594 1659
rect 3591 1626 3595 1627
rect 3591 1621 3595 1622
rect 3592 1593 3594 1621
rect 3590 1592 3596 1593
rect 3590 1588 3591 1592
rect 3595 1588 3596 1592
rect 3590 1587 3596 1588
rect 3526 1583 3532 1584
rect 3526 1579 3527 1583
rect 3531 1579 3532 1583
rect 3526 1578 3532 1579
rect 3590 1575 3596 1576
rect 3502 1572 3508 1573
rect 3502 1568 3503 1572
rect 3507 1568 3508 1572
rect 3590 1571 3591 1575
rect 3595 1571 3596 1575
rect 3590 1570 3596 1571
rect 3502 1567 3508 1568
rect 3504 1547 3506 1567
rect 3592 1547 3594 1570
rect 3495 1546 3499 1547
rect 3495 1541 3499 1542
rect 3503 1546 3507 1547
rect 3503 1541 3507 1542
rect 3591 1546 3595 1547
rect 3591 1541 3595 1542
rect 3496 1525 3498 1541
rect 3494 1524 3500 1525
rect 3494 1520 3495 1524
rect 3499 1520 3500 1524
rect 3592 1522 3594 1541
rect 3494 1519 3500 1520
rect 3590 1521 3596 1522
rect 3590 1517 3591 1521
rect 3595 1517 3596 1521
rect 3590 1516 3596 1517
rect 3590 1504 3596 1505
rect 3590 1500 3591 1504
rect 3595 1500 3596 1504
rect 3590 1499 3596 1500
rect 3502 1486 3508 1487
rect 3502 1482 3503 1486
rect 3507 1482 3508 1486
rect 3502 1481 3508 1482
rect 3504 1467 3506 1481
rect 3592 1467 3594 1499
rect 3503 1466 3507 1467
rect 3503 1461 3507 1462
rect 3591 1466 3595 1467
rect 3591 1461 3595 1462
rect 3592 1433 3594 1461
rect 3590 1432 3596 1433
rect 3590 1428 3591 1432
rect 3595 1428 3596 1432
rect 3590 1427 3596 1428
rect 3590 1415 3596 1416
rect 3590 1411 3591 1415
rect 3595 1411 3596 1415
rect 3590 1410 3596 1411
rect 3592 1391 3594 1410
rect 3503 1390 3507 1391
rect 3503 1385 3507 1386
rect 3591 1390 3595 1391
rect 3591 1385 3595 1386
rect 3504 1369 3506 1385
rect 3502 1368 3508 1369
rect 3502 1364 3503 1368
rect 3507 1364 3508 1368
rect 3592 1366 3594 1385
rect 3502 1363 3508 1364
rect 3590 1365 3596 1366
rect 3590 1361 3591 1365
rect 3595 1361 3596 1365
rect 3590 1360 3596 1361
rect 3486 1359 3492 1360
rect 3486 1355 3487 1359
rect 3491 1355 3492 1359
rect 3486 1354 3492 1355
rect 3590 1348 3596 1349
rect 3590 1344 3591 1348
rect 3595 1344 3596 1348
rect 3590 1343 3596 1344
rect 3510 1330 3516 1331
rect 3510 1326 3511 1330
rect 3515 1326 3516 1330
rect 3510 1325 3516 1326
rect 3414 1319 3420 1320
rect 3414 1315 3415 1319
rect 3419 1315 3420 1319
rect 3414 1314 3420 1315
rect 3512 1303 3514 1325
rect 3518 1319 3524 1320
rect 3518 1315 3519 1319
rect 3523 1315 3524 1319
rect 3518 1314 3524 1315
rect 3287 1302 3291 1303
rect 3287 1297 3291 1298
rect 3367 1302 3371 1303
rect 3367 1297 3371 1298
rect 3407 1302 3411 1303
rect 3407 1297 3411 1298
rect 3511 1302 3515 1303
rect 3511 1297 3515 1298
rect 3226 1295 3232 1296
rect 3226 1291 3227 1295
rect 3231 1291 3232 1295
rect 3226 1290 3232 1291
rect 3266 1295 3272 1296
rect 3266 1291 3267 1295
rect 3271 1291 3272 1295
rect 3266 1290 3272 1291
rect 3070 1286 3076 1287
rect 3070 1282 3071 1286
rect 3075 1282 3076 1286
rect 3070 1281 3076 1282
rect 3214 1286 3220 1287
rect 3214 1282 3215 1286
rect 3219 1282 3220 1286
rect 3214 1281 3220 1282
rect 3268 1260 3270 1290
rect 3368 1287 3370 1297
rect 3512 1287 3514 1297
rect 3366 1286 3372 1287
rect 3366 1282 3367 1286
rect 3371 1282 3372 1286
rect 3366 1281 3372 1282
rect 3510 1286 3516 1287
rect 3510 1282 3511 1286
rect 3515 1282 3516 1286
rect 3510 1281 3516 1282
rect 3520 1260 3522 1314
rect 3592 1303 3594 1343
rect 3591 1302 3595 1303
rect 3591 1297 3595 1298
rect 3592 1269 3594 1297
rect 3590 1268 3596 1269
rect 3590 1264 3591 1268
rect 3595 1264 3596 1268
rect 3590 1263 3596 1264
rect 1550 1259 1556 1260
rect 1550 1255 1551 1259
rect 1555 1255 1556 1259
rect 1550 1254 1556 1255
rect 2278 1259 2284 1260
rect 2278 1255 2279 1259
rect 2283 1255 2284 1259
rect 2278 1254 2284 1255
rect 2358 1259 2364 1260
rect 2358 1255 2359 1259
rect 2363 1255 2364 1259
rect 2358 1254 2364 1255
rect 2654 1259 2660 1260
rect 2654 1255 2655 1259
rect 2659 1255 2660 1259
rect 2654 1254 2660 1255
rect 2670 1259 2676 1260
rect 2670 1255 2671 1259
rect 2675 1255 2676 1259
rect 2670 1254 2676 1255
rect 2850 1259 2856 1260
rect 2850 1255 2851 1259
rect 2855 1255 2856 1259
rect 2850 1254 2856 1255
rect 2998 1259 3004 1260
rect 2998 1255 2999 1259
rect 3003 1255 3004 1259
rect 2998 1254 3004 1255
rect 3266 1259 3272 1260
rect 3266 1255 3267 1259
rect 3271 1255 3272 1259
rect 3266 1254 3272 1255
rect 3518 1259 3524 1260
rect 3518 1255 3519 1259
rect 3523 1255 3524 1259
rect 3518 1254 3524 1255
rect 1538 1251 1544 1252
rect 1538 1247 1539 1251
rect 1543 1247 1544 1251
rect 1538 1246 1544 1247
rect 1358 1230 1364 1231
rect 1358 1226 1359 1230
rect 1363 1226 1364 1230
rect 1358 1225 1364 1226
rect 1486 1230 1492 1231
rect 1486 1226 1487 1230
rect 1491 1226 1492 1230
rect 1486 1225 1492 1226
rect 1342 1219 1348 1220
rect 1342 1215 1343 1219
rect 1347 1215 1348 1219
rect 1342 1214 1348 1215
rect 1302 1207 1308 1208
rect 1360 1207 1362 1225
rect 1488 1207 1490 1225
rect 1540 1220 1542 1246
rect 1552 1220 1554 1254
rect 1870 1251 1876 1252
rect 1830 1248 1836 1249
rect 1830 1244 1831 1248
rect 1835 1244 1836 1248
rect 1870 1247 1871 1251
rect 1875 1247 1876 1251
rect 3590 1251 3596 1252
rect 1870 1246 1876 1247
rect 2206 1248 2212 1249
rect 1830 1243 1836 1244
rect 1614 1230 1620 1231
rect 1614 1226 1615 1230
rect 1619 1226 1620 1230
rect 1614 1225 1620 1226
rect 1742 1230 1748 1231
rect 1742 1226 1743 1230
rect 1747 1226 1748 1230
rect 1742 1225 1748 1226
rect 1538 1219 1544 1220
rect 1538 1215 1539 1219
rect 1543 1215 1544 1219
rect 1538 1214 1544 1215
rect 1550 1219 1556 1220
rect 1550 1215 1551 1219
rect 1555 1215 1556 1219
rect 1550 1214 1556 1215
rect 1570 1207 1576 1208
rect 1616 1207 1618 1225
rect 1744 1207 1746 1225
rect 1758 1219 1764 1220
rect 1758 1215 1759 1219
rect 1763 1215 1764 1219
rect 1758 1214 1764 1215
rect 1295 1206 1299 1207
rect 1302 1203 1303 1207
rect 1307 1203 1308 1207
rect 1302 1202 1308 1203
rect 1359 1206 1363 1207
rect 1295 1201 1299 1202
rect 1282 1199 1288 1200
rect 1282 1195 1283 1199
rect 1287 1195 1288 1199
rect 1282 1194 1288 1195
rect 1296 1191 1298 1201
rect 1158 1190 1164 1191
rect 1158 1186 1159 1190
rect 1163 1186 1164 1190
rect 1158 1185 1164 1186
rect 1294 1190 1300 1191
rect 1294 1186 1295 1190
rect 1299 1186 1300 1190
rect 1294 1185 1300 1186
rect 1304 1164 1306 1202
rect 1359 1201 1363 1202
rect 1415 1206 1419 1207
rect 1415 1201 1419 1202
rect 1487 1206 1491 1207
rect 1487 1201 1491 1202
rect 1535 1206 1539 1207
rect 1570 1203 1571 1207
rect 1575 1203 1576 1207
rect 1570 1202 1576 1203
rect 1615 1206 1619 1207
rect 1535 1201 1539 1202
rect 1416 1191 1418 1201
rect 1466 1199 1472 1200
rect 1466 1195 1467 1199
rect 1471 1195 1472 1199
rect 1466 1194 1472 1195
rect 1414 1190 1420 1191
rect 1414 1186 1415 1190
rect 1419 1186 1420 1190
rect 1414 1185 1420 1186
rect 1468 1164 1470 1194
rect 1536 1191 1538 1201
rect 1534 1190 1540 1191
rect 1534 1186 1535 1190
rect 1539 1186 1540 1190
rect 1534 1185 1540 1186
rect 898 1163 904 1164
rect 898 1159 899 1163
rect 903 1159 904 1163
rect 898 1158 904 1159
rect 1058 1163 1064 1164
rect 1058 1159 1059 1163
rect 1063 1159 1064 1163
rect 1058 1158 1064 1159
rect 1210 1163 1216 1164
rect 1210 1159 1211 1163
rect 1215 1159 1216 1163
rect 1210 1158 1216 1159
rect 1302 1163 1308 1164
rect 1302 1159 1303 1163
rect 1307 1159 1308 1163
rect 1302 1158 1308 1159
rect 1466 1163 1472 1164
rect 1466 1159 1467 1163
rect 1471 1159 1472 1163
rect 1466 1158 1472 1159
rect 998 1152 1004 1153
rect 998 1148 999 1152
rect 1003 1148 1004 1152
rect 998 1147 1004 1148
rect 1150 1152 1156 1153
rect 1150 1148 1151 1152
rect 1155 1148 1156 1152
rect 1150 1147 1156 1148
rect 1000 1131 1002 1147
rect 1152 1131 1154 1147
rect 895 1130 899 1131
rect 895 1125 899 1126
rect 999 1130 1003 1131
rect 999 1125 1003 1126
rect 1015 1130 1019 1131
rect 1015 1125 1019 1126
rect 1135 1130 1139 1131
rect 1135 1125 1139 1126
rect 1151 1130 1155 1131
rect 1151 1125 1155 1126
rect 896 1109 898 1125
rect 1016 1109 1018 1125
rect 1136 1109 1138 1125
rect 894 1108 900 1109
rect 894 1104 895 1108
rect 899 1104 900 1108
rect 894 1103 900 1104
rect 1014 1108 1020 1109
rect 1014 1104 1015 1108
rect 1019 1104 1020 1108
rect 1014 1103 1020 1104
rect 1134 1108 1140 1109
rect 1134 1104 1135 1108
rect 1139 1104 1140 1108
rect 1134 1103 1140 1104
rect 314 1099 320 1100
rect 314 1095 315 1099
rect 319 1095 320 1099
rect 314 1094 320 1095
rect 458 1099 464 1100
rect 458 1095 459 1099
rect 463 1095 464 1099
rect 458 1094 464 1095
rect 718 1099 724 1100
rect 718 1095 719 1099
rect 723 1095 724 1099
rect 718 1094 724 1095
rect 854 1099 860 1100
rect 854 1095 855 1099
rect 859 1095 860 1099
rect 854 1094 860 1095
rect 962 1099 968 1100
rect 962 1095 963 1099
rect 967 1095 968 1099
rect 962 1094 968 1095
rect 1082 1099 1088 1100
rect 1082 1095 1083 1099
rect 1087 1095 1088 1099
rect 1082 1094 1088 1095
rect 316 1060 318 1094
rect 390 1070 396 1071
rect 390 1066 391 1070
rect 395 1066 396 1070
rect 390 1065 396 1066
rect 262 1059 268 1060
rect 262 1055 263 1059
rect 267 1055 268 1059
rect 262 1054 268 1055
rect 314 1059 320 1060
rect 314 1055 315 1059
rect 319 1055 320 1059
rect 314 1054 320 1055
rect 392 1043 394 1065
rect 460 1060 462 1094
rect 526 1070 532 1071
rect 526 1066 527 1070
rect 531 1066 532 1070
rect 526 1065 532 1066
rect 654 1070 660 1071
rect 654 1066 655 1070
rect 659 1066 660 1070
rect 654 1065 660 1066
rect 458 1059 464 1060
rect 458 1055 459 1059
rect 463 1055 464 1059
rect 458 1054 464 1055
rect 528 1043 530 1065
rect 626 1059 632 1060
rect 626 1055 627 1059
rect 631 1055 632 1059
rect 626 1054 632 1055
rect 239 1042 243 1043
rect 239 1037 243 1038
rect 255 1042 259 1043
rect 255 1037 259 1038
rect 359 1042 363 1043
rect 359 1037 363 1038
rect 391 1042 395 1043
rect 391 1037 395 1038
rect 471 1042 475 1043
rect 471 1037 475 1038
rect 527 1042 531 1043
rect 527 1037 531 1038
rect 575 1042 579 1043
rect 575 1037 579 1038
rect 240 1027 242 1037
rect 298 1035 304 1036
rect 298 1031 299 1035
rect 303 1031 304 1035
rect 298 1030 304 1031
rect 238 1026 244 1027
rect 238 1022 239 1026
rect 243 1022 244 1026
rect 238 1021 244 1022
rect 300 1000 302 1030
rect 360 1027 362 1037
rect 472 1027 474 1037
rect 534 1035 540 1036
rect 534 1031 535 1035
rect 539 1031 540 1035
rect 534 1030 540 1031
rect 358 1026 364 1027
rect 358 1022 359 1026
rect 363 1022 364 1026
rect 358 1021 364 1022
rect 470 1026 476 1027
rect 470 1022 471 1026
rect 475 1022 476 1026
rect 470 1021 476 1022
rect 536 1000 538 1030
rect 576 1027 578 1037
rect 574 1026 580 1027
rect 574 1022 575 1026
rect 579 1022 580 1026
rect 574 1021 580 1022
rect 628 1000 630 1054
rect 656 1043 658 1065
rect 720 1060 722 1094
rect 782 1070 788 1071
rect 782 1066 783 1070
rect 787 1066 788 1070
rect 782 1065 788 1066
rect 902 1070 908 1071
rect 902 1066 903 1070
rect 907 1066 908 1070
rect 902 1065 908 1066
rect 718 1059 724 1060
rect 718 1055 719 1059
rect 723 1055 724 1059
rect 718 1054 724 1055
rect 678 1043 684 1044
rect 784 1043 786 1065
rect 904 1043 906 1065
rect 964 1060 966 1094
rect 1022 1070 1028 1071
rect 1022 1066 1023 1070
rect 1027 1066 1028 1070
rect 1022 1065 1028 1066
rect 962 1059 968 1060
rect 962 1055 963 1059
rect 967 1055 968 1059
rect 962 1054 968 1055
rect 1024 1043 1026 1065
rect 1084 1060 1086 1094
rect 1194 1091 1200 1092
rect 1194 1087 1195 1091
rect 1199 1087 1200 1091
rect 1194 1086 1200 1087
rect 1142 1070 1148 1071
rect 1142 1066 1143 1070
rect 1147 1066 1148 1070
rect 1142 1065 1148 1066
rect 1082 1059 1088 1060
rect 1082 1055 1083 1059
rect 1087 1055 1088 1059
rect 1082 1054 1088 1055
rect 1144 1043 1146 1065
rect 1196 1060 1198 1086
rect 1212 1060 1214 1158
rect 1286 1152 1292 1153
rect 1286 1148 1287 1152
rect 1291 1148 1292 1152
rect 1286 1147 1292 1148
rect 1406 1152 1412 1153
rect 1406 1148 1407 1152
rect 1411 1148 1412 1152
rect 1406 1147 1412 1148
rect 1526 1152 1532 1153
rect 1526 1148 1527 1152
rect 1531 1148 1532 1152
rect 1526 1147 1532 1148
rect 1288 1131 1290 1147
rect 1408 1131 1410 1147
rect 1528 1131 1530 1147
rect 1255 1130 1259 1131
rect 1255 1125 1259 1126
rect 1287 1130 1291 1131
rect 1287 1125 1291 1126
rect 1375 1130 1379 1131
rect 1375 1125 1379 1126
rect 1407 1130 1411 1131
rect 1407 1125 1411 1126
rect 1503 1130 1507 1131
rect 1503 1125 1507 1126
rect 1527 1130 1531 1131
rect 1527 1125 1531 1126
rect 1256 1109 1258 1125
rect 1376 1109 1378 1125
rect 1504 1109 1506 1125
rect 1254 1108 1260 1109
rect 1254 1104 1255 1108
rect 1259 1104 1260 1108
rect 1254 1103 1260 1104
rect 1374 1108 1380 1109
rect 1374 1104 1375 1108
rect 1379 1104 1380 1108
rect 1374 1103 1380 1104
rect 1502 1108 1508 1109
rect 1502 1104 1503 1108
rect 1507 1104 1508 1108
rect 1502 1103 1508 1104
rect 1572 1100 1574 1202
rect 1615 1201 1619 1202
rect 1655 1206 1659 1207
rect 1655 1201 1659 1202
rect 1743 1206 1747 1207
rect 1743 1201 1747 1202
rect 1751 1206 1755 1207
rect 1751 1201 1755 1202
rect 1586 1199 1592 1200
rect 1586 1195 1587 1199
rect 1591 1195 1592 1199
rect 1586 1194 1592 1195
rect 1588 1164 1590 1194
rect 1656 1191 1658 1201
rect 1706 1199 1712 1200
rect 1706 1195 1707 1199
rect 1711 1195 1712 1199
rect 1706 1194 1712 1195
rect 1654 1190 1660 1191
rect 1654 1186 1655 1190
rect 1659 1186 1660 1190
rect 1654 1185 1660 1186
rect 1708 1164 1710 1194
rect 1752 1191 1754 1201
rect 1750 1190 1756 1191
rect 1750 1186 1751 1190
rect 1755 1186 1756 1190
rect 1750 1185 1756 1186
rect 1760 1164 1762 1214
rect 1832 1207 1834 1243
rect 1872 1223 1874 1246
rect 2206 1244 2207 1248
rect 2211 1244 2212 1248
rect 2206 1243 2212 1244
rect 2286 1248 2292 1249
rect 2286 1244 2287 1248
rect 2291 1244 2292 1248
rect 2286 1243 2292 1244
rect 2366 1248 2372 1249
rect 2366 1244 2367 1248
rect 2371 1244 2372 1248
rect 2366 1243 2372 1244
rect 2446 1248 2452 1249
rect 2446 1244 2447 1248
rect 2451 1244 2452 1248
rect 2446 1243 2452 1244
rect 2542 1248 2548 1249
rect 2542 1244 2543 1248
rect 2547 1244 2548 1248
rect 2542 1243 2548 1244
rect 2654 1248 2660 1249
rect 2654 1244 2655 1248
rect 2659 1244 2660 1248
rect 2654 1243 2660 1244
rect 2782 1248 2788 1249
rect 2782 1244 2783 1248
rect 2787 1244 2788 1248
rect 2782 1243 2788 1244
rect 2918 1248 2924 1249
rect 2918 1244 2919 1248
rect 2923 1244 2924 1248
rect 2918 1243 2924 1244
rect 3062 1248 3068 1249
rect 3062 1244 3063 1248
rect 3067 1244 3068 1248
rect 3062 1243 3068 1244
rect 3206 1248 3212 1249
rect 3206 1244 3207 1248
rect 3211 1244 3212 1248
rect 3206 1243 3212 1244
rect 3358 1248 3364 1249
rect 3358 1244 3359 1248
rect 3363 1244 3364 1248
rect 3358 1243 3364 1244
rect 3502 1248 3508 1249
rect 3502 1244 3503 1248
rect 3507 1244 3508 1248
rect 3590 1247 3591 1251
rect 3595 1247 3596 1251
rect 3590 1246 3596 1247
rect 3502 1243 3508 1244
rect 2126 1231 2132 1232
rect 2126 1227 2127 1231
rect 2131 1227 2132 1231
rect 2126 1226 2132 1227
rect 1871 1222 1875 1223
rect 1871 1217 1875 1218
rect 2111 1222 2115 1223
rect 2111 1217 2115 1218
rect 1831 1206 1835 1207
rect 1831 1201 1835 1202
rect 1832 1173 1834 1201
rect 1872 1198 1874 1217
rect 2112 1201 2114 1217
rect 2110 1200 2116 1201
rect 1870 1197 1876 1198
rect 1870 1193 1871 1197
rect 1875 1193 1876 1197
rect 2110 1196 2111 1200
rect 2115 1196 2116 1200
rect 2110 1195 2116 1196
rect 1870 1192 1876 1193
rect 1870 1180 1876 1181
rect 1870 1176 1871 1180
rect 1875 1176 1876 1180
rect 1870 1175 1876 1176
rect 1830 1172 1836 1173
rect 1830 1168 1831 1172
rect 1835 1168 1836 1172
rect 1830 1167 1836 1168
rect 1586 1163 1592 1164
rect 1586 1159 1587 1163
rect 1591 1159 1592 1163
rect 1586 1158 1592 1159
rect 1706 1163 1712 1164
rect 1706 1159 1707 1163
rect 1711 1159 1712 1163
rect 1706 1158 1712 1159
rect 1758 1163 1764 1164
rect 1758 1159 1759 1163
rect 1763 1159 1764 1163
rect 1758 1158 1764 1159
rect 1830 1155 1836 1156
rect 1646 1152 1652 1153
rect 1646 1148 1647 1152
rect 1651 1148 1652 1152
rect 1646 1147 1652 1148
rect 1742 1152 1748 1153
rect 1742 1148 1743 1152
rect 1747 1148 1748 1152
rect 1830 1151 1831 1155
rect 1835 1151 1836 1155
rect 1830 1150 1836 1151
rect 1742 1147 1748 1148
rect 1648 1131 1650 1147
rect 1744 1131 1746 1147
rect 1832 1131 1834 1150
rect 1872 1139 1874 1175
rect 2118 1162 2124 1163
rect 2118 1158 2119 1162
rect 2123 1158 2124 1162
rect 2118 1157 2124 1158
rect 2120 1139 2122 1157
rect 2128 1152 2130 1226
rect 2208 1223 2210 1243
rect 2288 1223 2290 1243
rect 2368 1223 2370 1243
rect 2448 1223 2450 1243
rect 2544 1223 2546 1243
rect 2656 1223 2658 1243
rect 2662 1231 2668 1232
rect 2662 1227 2663 1231
rect 2667 1227 2668 1231
rect 2662 1226 2668 1227
rect 2207 1222 2211 1223
rect 2207 1217 2211 1218
rect 2287 1222 2291 1223
rect 2287 1217 2291 1218
rect 2303 1222 2307 1223
rect 2303 1217 2307 1218
rect 2367 1222 2371 1223
rect 2367 1217 2371 1218
rect 2407 1222 2411 1223
rect 2407 1217 2411 1218
rect 2447 1222 2451 1223
rect 2447 1217 2451 1218
rect 2527 1222 2531 1223
rect 2527 1217 2531 1218
rect 2543 1222 2547 1223
rect 2543 1217 2547 1218
rect 2647 1222 2651 1223
rect 2647 1217 2651 1218
rect 2655 1222 2659 1223
rect 2655 1217 2659 1218
rect 2208 1201 2210 1217
rect 2304 1201 2306 1217
rect 2408 1201 2410 1217
rect 2528 1201 2530 1217
rect 2648 1201 2650 1217
rect 2206 1200 2212 1201
rect 2206 1196 2207 1200
rect 2211 1196 2212 1200
rect 2206 1195 2212 1196
rect 2302 1200 2308 1201
rect 2302 1196 2303 1200
rect 2307 1196 2308 1200
rect 2302 1195 2308 1196
rect 2406 1200 2412 1201
rect 2406 1196 2407 1200
rect 2411 1196 2412 1200
rect 2406 1195 2412 1196
rect 2526 1200 2532 1201
rect 2526 1196 2527 1200
rect 2531 1196 2532 1200
rect 2526 1195 2532 1196
rect 2646 1200 2652 1201
rect 2646 1196 2647 1200
rect 2651 1196 2652 1200
rect 2646 1195 2652 1196
rect 2178 1191 2184 1192
rect 2178 1187 2179 1191
rect 2183 1187 2184 1191
rect 2178 1186 2184 1187
rect 2274 1191 2280 1192
rect 2274 1187 2275 1191
rect 2279 1187 2280 1191
rect 2274 1186 2280 1187
rect 2370 1191 2376 1192
rect 2370 1187 2371 1191
rect 2375 1187 2376 1191
rect 2370 1186 2376 1187
rect 2474 1191 2480 1192
rect 2474 1187 2475 1191
rect 2479 1187 2480 1191
rect 2474 1186 2480 1187
rect 2482 1191 2488 1192
rect 2482 1187 2483 1191
rect 2487 1187 2488 1191
rect 2482 1186 2488 1187
rect 2180 1152 2182 1186
rect 2214 1162 2220 1163
rect 2214 1158 2215 1162
rect 2219 1158 2220 1162
rect 2214 1157 2220 1158
rect 2126 1151 2132 1152
rect 2126 1147 2127 1151
rect 2131 1147 2132 1151
rect 2126 1146 2132 1147
rect 2178 1151 2184 1152
rect 2178 1147 2179 1151
rect 2183 1147 2184 1151
rect 2178 1146 2184 1147
rect 2216 1139 2218 1157
rect 2276 1152 2278 1186
rect 2310 1162 2316 1163
rect 2310 1158 2311 1162
rect 2315 1158 2316 1162
rect 2310 1157 2316 1158
rect 2274 1151 2280 1152
rect 2274 1147 2275 1151
rect 2279 1147 2280 1151
rect 2274 1146 2280 1147
rect 2312 1139 2314 1157
rect 2372 1152 2374 1186
rect 2414 1162 2420 1163
rect 2414 1158 2415 1162
rect 2419 1158 2420 1162
rect 2414 1157 2420 1158
rect 2370 1151 2376 1152
rect 2370 1147 2371 1151
rect 2375 1147 2376 1151
rect 2370 1146 2376 1147
rect 2416 1139 2418 1157
rect 2476 1152 2478 1186
rect 2474 1151 2480 1152
rect 2474 1147 2475 1151
rect 2479 1147 2480 1151
rect 2474 1146 2480 1147
rect 1871 1138 1875 1139
rect 1871 1133 1875 1134
rect 1903 1138 1907 1139
rect 1903 1133 1907 1134
rect 2119 1138 2123 1139
rect 2119 1133 2123 1134
rect 2127 1138 2131 1139
rect 2127 1133 2131 1134
rect 2215 1138 2219 1139
rect 2215 1133 2219 1134
rect 2311 1138 2315 1139
rect 2311 1133 2315 1134
rect 2359 1138 2363 1139
rect 2359 1133 2363 1134
rect 2415 1138 2419 1139
rect 2415 1133 2419 1134
rect 1631 1130 1635 1131
rect 1631 1125 1635 1126
rect 1647 1130 1651 1131
rect 1647 1125 1651 1126
rect 1743 1130 1747 1131
rect 1743 1125 1747 1126
rect 1831 1130 1835 1131
rect 1831 1125 1835 1126
rect 1632 1109 1634 1125
rect 1744 1109 1746 1125
rect 1630 1108 1636 1109
rect 1630 1104 1631 1108
rect 1635 1104 1636 1108
rect 1630 1103 1636 1104
rect 1742 1108 1748 1109
rect 1742 1104 1743 1108
rect 1747 1104 1748 1108
rect 1832 1106 1834 1125
rect 1742 1103 1748 1104
rect 1830 1105 1836 1106
rect 1872 1105 1874 1133
rect 1904 1123 1906 1133
rect 2128 1123 2130 1133
rect 2360 1123 2362 1133
rect 2484 1132 2486 1186
rect 2583 1164 2587 1165
rect 2534 1162 2540 1163
rect 2534 1158 2535 1162
rect 2539 1158 2540 1162
rect 2583 1159 2587 1160
rect 2654 1162 2660 1163
rect 2534 1157 2540 1158
rect 2536 1139 2538 1157
rect 2535 1138 2539 1139
rect 2535 1133 2539 1134
rect 2575 1138 2579 1139
rect 2575 1133 2579 1134
rect 2482 1131 2488 1132
rect 2482 1127 2483 1131
rect 2487 1127 2488 1131
rect 2482 1126 2488 1127
rect 2576 1123 2578 1133
rect 2584 1132 2586 1159
rect 2654 1158 2655 1162
rect 2659 1158 2660 1162
rect 2654 1157 2660 1158
rect 2656 1139 2658 1157
rect 2664 1152 2666 1226
rect 2784 1223 2786 1243
rect 2920 1223 2922 1243
rect 3064 1223 3066 1243
rect 3208 1223 3210 1243
rect 3360 1223 3362 1243
rect 3366 1231 3372 1232
rect 3366 1227 3367 1231
rect 3371 1227 3372 1231
rect 3366 1226 3372 1227
rect 2775 1222 2779 1223
rect 2775 1217 2779 1218
rect 2783 1222 2787 1223
rect 2783 1217 2787 1218
rect 2911 1222 2915 1223
rect 2911 1217 2915 1218
rect 2919 1222 2923 1223
rect 2919 1217 2923 1218
rect 3055 1222 3059 1223
rect 3055 1217 3059 1218
rect 3063 1222 3067 1223
rect 3063 1217 3067 1218
rect 3199 1222 3203 1223
rect 3199 1217 3203 1218
rect 3207 1222 3211 1223
rect 3207 1217 3211 1218
rect 3343 1222 3347 1223
rect 3343 1217 3347 1218
rect 3359 1222 3363 1223
rect 3359 1217 3363 1218
rect 2776 1201 2778 1217
rect 2912 1201 2914 1217
rect 3056 1201 3058 1217
rect 3200 1201 3202 1217
rect 3344 1201 3346 1217
rect 2774 1200 2780 1201
rect 2774 1196 2775 1200
rect 2779 1196 2780 1200
rect 2774 1195 2780 1196
rect 2910 1200 2916 1201
rect 2910 1196 2911 1200
rect 2915 1196 2916 1200
rect 2910 1195 2916 1196
rect 3054 1200 3060 1201
rect 3054 1196 3055 1200
rect 3059 1196 3060 1200
rect 3054 1195 3060 1196
rect 3198 1200 3204 1201
rect 3198 1196 3199 1200
rect 3203 1196 3204 1200
rect 3198 1195 3204 1196
rect 3342 1200 3348 1201
rect 3342 1196 3343 1200
rect 3347 1196 3348 1200
rect 3342 1195 3348 1196
rect 2718 1191 2724 1192
rect 2718 1187 2719 1191
rect 2723 1187 2724 1191
rect 2718 1186 2724 1187
rect 2850 1191 2856 1192
rect 2850 1187 2851 1191
rect 2855 1187 2856 1191
rect 2850 1186 2856 1187
rect 2990 1191 2996 1192
rect 2990 1187 2991 1191
rect 2995 1187 2996 1191
rect 2990 1186 2996 1187
rect 2998 1191 3004 1192
rect 2998 1187 2999 1191
rect 3003 1187 3004 1191
rect 2998 1186 3004 1187
rect 3274 1191 3280 1192
rect 3274 1187 3275 1191
rect 3279 1187 3280 1191
rect 3274 1186 3280 1187
rect 3282 1191 3288 1192
rect 3282 1187 3283 1191
rect 3287 1187 3288 1191
rect 3282 1186 3288 1187
rect 2720 1152 2722 1186
rect 2782 1162 2788 1163
rect 2782 1158 2783 1162
rect 2787 1158 2788 1162
rect 2782 1157 2788 1158
rect 2662 1151 2668 1152
rect 2662 1147 2663 1151
rect 2667 1147 2668 1151
rect 2662 1146 2668 1147
rect 2718 1151 2724 1152
rect 2718 1147 2719 1151
rect 2723 1147 2724 1151
rect 2718 1146 2724 1147
rect 2784 1139 2786 1157
rect 2852 1152 2854 1186
rect 2918 1162 2924 1163
rect 2918 1158 2919 1162
rect 2923 1158 2924 1162
rect 2918 1157 2924 1158
rect 2850 1151 2856 1152
rect 2850 1147 2851 1151
rect 2855 1147 2856 1151
rect 2850 1146 2856 1147
rect 2920 1139 2922 1157
rect 2992 1152 2994 1186
rect 3000 1165 3002 1186
rect 2999 1164 3003 1165
rect 2999 1159 3003 1160
rect 3062 1162 3068 1163
rect 3062 1158 3063 1162
rect 3067 1158 3068 1162
rect 3062 1157 3068 1158
rect 3206 1162 3212 1163
rect 3206 1158 3207 1162
rect 3211 1158 3212 1162
rect 3206 1157 3212 1158
rect 2990 1151 2996 1152
rect 2990 1147 2991 1151
rect 2995 1147 2996 1151
rect 2990 1146 2996 1147
rect 3064 1139 3066 1157
rect 3208 1139 3210 1157
rect 2655 1138 2659 1139
rect 2655 1133 2659 1134
rect 2775 1138 2779 1139
rect 2775 1133 2779 1134
rect 2783 1138 2787 1139
rect 2783 1133 2787 1134
rect 2919 1138 2923 1139
rect 2919 1133 2923 1134
rect 2967 1138 2971 1139
rect 2967 1133 2971 1134
rect 3063 1138 3067 1139
rect 3063 1133 3067 1134
rect 3159 1138 3163 1139
rect 3159 1133 3163 1134
rect 3207 1138 3211 1139
rect 3207 1133 3211 1134
rect 2582 1131 2588 1132
rect 2582 1127 2583 1131
rect 2587 1127 2588 1131
rect 2582 1126 2588 1127
rect 2626 1131 2632 1132
rect 2626 1127 2627 1131
rect 2631 1127 2632 1131
rect 2626 1126 2632 1127
rect 1902 1122 1908 1123
rect 1902 1118 1903 1122
rect 1907 1118 1908 1122
rect 1902 1117 1908 1118
rect 2126 1122 2132 1123
rect 2126 1118 2127 1122
rect 2131 1118 2132 1122
rect 2126 1117 2132 1118
rect 2358 1122 2364 1123
rect 2358 1118 2359 1122
rect 2363 1118 2364 1122
rect 2358 1117 2364 1118
rect 2574 1122 2580 1123
rect 2574 1118 2575 1122
rect 2579 1118 2580 1122
rect 2574 1117 2580 1118
rect 1830 1101 1831 1105
rect 1835 1101 1836 1105
rect 1830 1100 1836 1101
rect 1870 1104 1876 1105
rect 1870 1100 1871 1104
rect 1875 1100 1876 1104
rect 1322 1099 1328 1100
rect 1322 1095 1323 1099
rect 1327 1095 1328 1099
rect 1322 1094 1328 1095
rect 1442 1099 1448 1100
rect 1442 1095 1443 1099
rect 1447 1095 1448 1099
rect 1442 1094 1448 1095
rect 1570 1099 1576 1100
rect 1570 1095 1571 1099
rect 1575 1095 1576 1099
rect 1570 1094 1576 1095
rect 1698 1099 1704 1100
rect 1870 1099 1876 1100
rect 1698 1095 1699 1099
rect 1703 1095 1704 1099
rect 2628 1096 2630 1126
rect 2776 1123 2778 1133
rect 2826 1131 2832 1132
rect 2826 1127 2827 1131
rect 2831 1127 2832 1131
rect 2826 1126 2832 1127
rect 2774 1122 2780 1123
rect 2774 1118 2775 1122
rect 2779 1118 2780 1122
rect 2774 1117 2780 1118
rect 2828 1096 2830 1126
rect 2968 1123 2970 1133
rect 3160 1123 3162 1133
rect 3276 1132 3278 1186
rect 3284 1152 3286 1186
rect 3350 1162 3356 1163
rect 3350 1158 3351 1162
rect 3355 1158 3356 1162
rect 3350 1157 3356 1158
rect 3282 1151 3288 1152
rect 3282 1147 3283 1151
rect 3287 1147 3288 1151
rect 3282 1146 3288 1147
rect 3352 1139 3354 1157
rect 3368 1152 3370 1226
rect 3504 1223 3506 1243
rect 3592 1223 3594 1246
rect 3495 1222 3499 1223
rect 3495 1217 3499 1218
rect 3503 1222 3507 1223
rect 3503 1217 3507 1218
rect 3591 1222 3595 1223
rect 3591 1217 3595 1218
rect 3496 1201 3498 1217
rect 3494 1200 3500 1201
rect 3494 1196 3495 1200
rect 3499 1196 3500 1200
rect 3592 1198 3594 1217
rect 3494 1195 3500 1196
rect 3590 1197 3596 1198
rect 3590 1193 3591 1197
rect 3595 1193 3596 1197
rect 3590 1192 3596 1193
rect 3590 1180 3596 1181
rect 3590 1176 3591 1180
rect 3595 1176 3596 1180
rect 3590 1175 3596 1176
rect 3502 1162 3508 1163
rect 3502 1158 3503 1162
rect 3507 1158 3508 1162
rect 3502 1157 3508 1158
rect 3366 1151 3372 1152
rect 3366 1147 3367 1151
rect 3371 1147 3372 1151
rect 3366 1146 3372 1147
rect 3504 1139 3506 1157
rect 3518 1151 3524 1152
rect 3518 1147 3519 1151
rect 3523 1147 3524 1151
rect 3518 1146 3524 1147
rect 3343 1138 3347 1139
rect 3343 1133 3347 1134
rect 3351 1138 3355 1139
rect 3351 1133 3355 1134
rect 3503 1138 3507 1139
rect 3503 1133 3507 1134
rect 3511 1138 3515 1139
rect 3511 1133 3515 1134
rect 3254 1131 3260 1132
rect 3254 1127 3255 1131
rect 3259 1127 3260 1131
rect 3254 1126 3260 1127
rect 3274 1131 3280 1132
rect 3274 1127 3275 1131
rect 3279 1127 3280 1131
rect 3274 1126 3280 1127
rect 2966 1122 2972 1123
rect 2966 1118 2967 1122
rect 2971 1118 2972 1122
rect 2966 1117 2972 1118
rect 3158 1122 3164 1123
rect 3158 1118 3159 1122
rect 3163 1118 3164 1122
rect 3158 1117 3164 1118
rect 3256 1096 3258 1126
rect 3344 1123 3346 1133
rect 3512 1123 3514 1133
rect 3342 1122 3348 1123
rect 3342 1118 3343 1122
rect 3347 1118 3348 1122
rect 3342 1117 3348 1118
rect 3510 1122 3516 1123
rect 3510 1118 3511 1122
rect 3515 1118 3516 1122
rect 3510 1117 3516 1118
rect 3520 1096 3522 1146
rect 3592 1139 3594 1175
rect 3591 1138 3595 1139
rect 3591 1133 3595 1134
rect 3592 1105 3594 1133
rect 3590 1104 3596 1105
rect 3590 1100 3591 1104
rect 3595 1100 3596 1104
rect 3590 1099 3596 1100
rect 1698 1094 1704 1095
rect 2214 1095 2220 1096
rect 1262 1070 1268 1071
rect 1262 1066 1263 1070
rect 1267 1066 1268 1070
rect 1262 1065 1268 1066
rect 1194 1059 1200 1060
rect 1194 1055 1195 1059
rect 1199 1055 1200 1059
rect 1194 1054 1200 1055
rect 1210 1059 1216 1060
rect 1210 1055 1211 1059
rect 1215 1055 1216 1059
rect 1210 1054 1216 1055
rect 1264 1043 1266 1065
rect 1324 1060 1326 1094
rect 1382 1070 1388 1071
rect 1382 1066 1383 1070
rect 1387 1066 1388 1070
rect 1382 1065 1388 1066
rect 1322 1059 1328 1060
rect 1322 1055 1323 1059
rect 1327 1055 1328 1059
rect 1322 1054 1328 1055
rect 1384 1043 1386 1065
rect 1444 1060 1446 1094
rect 1510 1070 1516 1071
rect 1510 1066 1511 1070
rect 1515 1066 1516 1070
rect 1510 1065 1516 1066
rect 1638 1070 1644 1071
rect 1638 1066 1639 1070
rect 1643 1066 1644 1070
rect 1638 1065 1644 1066
rect 1442 1059 1448 1060
rect 1442 1055 1443 1059
rect 1447 1055 1448 1059
rect 1442 1054 1448 1055
rect 1512 1043 1514 1065
rect 1640 1043 1642 1065
rect 1700 1060 1702 1094
rect 2214 1091 2215 1095
rect 2219 1091 2220 1095
rect 2214 1090 2220 1091
rect 2626 1095 2632 1096
rect 2626 1091 2627 1095
rect 2631 1091 2632 1095
rect 2626 1090 2632 1091
rect 2826 1095 2832 1096
rect 2826 1091 2827 1095
rect 2831 1091 2832 1095
rect 2826 1090 2832 1091
rect 3018 1095 3024 1096
rect 3018 1091 3019 1095
rect 3023 1091 3024 1095
rect 3018 1090 3024 1091
rect 3210 1095 3216 1096
rect 3210 1091 3211 1095
rect 3215 1091 3216 1095
rect 3210 1090 3216 1091
rect 3254 1095 3260 1096
rect 3254 1091 3255 1095
rect 3259 1091 3260 1095
rect 3254 1090 3260 1091
rect 3518 1095 3524 1096
rect 3518 1091 3519 1095
rect 3523 1091 3524 1095
rect 3518 1090 3524 1091
rect 1830 1088 1836 1089
rect 1830 1084 1831 1088
rect 1835 1084 1836 1088
rect 1830 1083 1836 1084
rect 1870 1087 1876 1088
rect 1870 1083 1871 1087
rect 1875 1083 1876 1087
rect 1750 1070 1756 1071
rect 1750 1066 1751 1070
rect 1755 1066 1756 1070
rect 1750 1065 1756 1066
rect 1698 1059 1704 1060
rect 1698 1055 1699 1059
rect 1703 1055 1704 1059
rect 1698 1054 1704 1055
rect 1752 1043 1754 1065
rect 1832 1043 1834 1083
rect 1870 1082 1876 1083
rect 1894 1084 1900 1085
rect 1872 1063 1874 1082
rect 1894 1080 1895 1084
rect 1899 1080 1900 1084
rect 1894 1079 1900 1080
rect 2118 1084 2124 1085
rect 2118 1080 2119 1084
rect 2123 1080 2124 1084
rect 2118 1079 2124 1080
rect 1896 1063 1898 1079
rect 2120 1063 2122 1079
rect 1871 1062 1875 1063
rect 1871 1057 1875 1058
rect 1895 1062 1899 1063
rect 1895 1057 1899 1058
rect 2015 1062 2019 1063
rect 2015 1057 2019 1058
rect 2119 1062 2123 1063
rect 2119 1057 2123 1058
rect 2167 1062 2171 1063
rect 2167 1057 2171 1058
rect 655 1042 659 1043
rect 655 1037 659 1038
rect 671 1042 675 1043
rect 678 1039 679 1043
rect 683 1039 684 1043
rect 678 1038 684 1039
rect 767 1042 771 1043
rect 671 1037 675 1038
rect 672 1027 674 1037
rect 670 1026 676 1027
rect 670 1022 671 1026
rect 675 1022 676 1026
rect 670 1021 676 1022
rect 680 1000 682 1038
rect 767 1037 771 1038
rect 783 1042 787 1043
rect 783 1037 787 1038
rect 855 1042 859 1043
rect 855 1037 859 1038
rect 903 1042 907 1043
rect 903 1037 907 1038
rect 943 1042 947 1043
rect 943 1037 947 1038
rect 1023 1042 1027 1043
rect 1023 1037 1027 1038
rect 1031 1042 1035 1043
rect 1031 1037 1035 1038
rect 1127 1042 1131 1043
rect 1127 1037 1131 1038
rect 1143 1042 1147 1043
rect 1143 1037 1147 1038
rect 1223 1042 1227 1043
rect 1223 1037 1227 1038
rect 1263 1042 1267 1043
rect 1263 1037 1267 1038
rect 1383 1042 1387 1043
rect 1383 1037 1387 1038
rect 1511 1042 1515 1043
rect 1511 1037 1515 1038
rect 1639 1042 1643 1043
rect 1639 1037 1643 1038
rect 1751 1042 1755 1043
rect 1751 1037 1755 1038
rect 1831 1042 1835 1043
rect 1872 1038 1874 1057
rect 1896 1041 1898 1057
rect 2016 1041 2018 1057
rect 2168 1041 2170 1057
rect 1894 1040 1900 1041
rect 1831 1037 1835 1038
rect 1870 1037 1876 1038
rect 686 1035 692 1036
rect 686 1031 687 1035
rect 691 1031 692 1035
rect 686 1030 692 1031
rect 150 999 156 1000
rect 150 995 151 999
rect 155 995 156 999
rect 150 994 156 995
rect 298 999 304 1000
rect 298 995 299 999
rect 303 995 304 999
rect 298 994 304 995
rect 534 999 540 1000
rect 534 995 535 999
rect 539 995 540 999
rect 534 994 540 995
rect 626 999 632 1000
rect 626 995 627 999
rect 631 995 632 999
rect 626 994 632 995
rect 678 999 684 1000
rect 678 995 679 999
rect 683 995 684 999
rect 678 994 684 995
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 110 986 116 987
rect 134 988 140 989
rect 112 955 114 986
rect 134 984 135 988
rect 139 984 140 988
rect 134 983 140 984
rect 230 988 236 989
rect 230 984 231 988
rect 235 984 236 988
rect 230 983 236 984
rect 350 988 356 989
rect 350 984 351 988
rect 355 984 356 988
rect 350 983 356 984
rect 462 988 468 989
rect 462 984 463 988
rect 467 984 468 988
rect 462 983 468 984
rect 566 988 572 989
rect 566 984 567 988
rect 571 984 572 988
rect 566 983 572 984
rect 662 988 668 989
rect 662 984 663 988
rect 667 984 668 988
rect 662 983 668 984
rect 136 955 138 983
rect 232 955 234 983
rect 352 955 354 983
rect 464 955 466 983
rect 568 955 570 983
rect 664 955 666 983
rect 111 954 115 955
rect 111 949 115 950
rect 135 954 139 955
rect 135 949 139 950
rect 231 954 235 955
rect 231 949 235 950
rect 263 954 267 955
rect 263 949 267 950
rect 351 954 355 955
rect 351 949 355 950
rect 415 954 419 955
rect 415 949 419 950
rect 463 954 467 955
rect 463 949 467 950
rect 559 954 563 955
rect 559 949 563 950
rect 567 954 571 955
rect 567 949 571 950
rect 663 954 667 955
rect 663 949 667 950
rect 112 930 114 949
rect 136 933 138 949
rect 264 933 266 949
rect 416 933 418 949
rect 560 933 562 949
rect 134 932 140 933
rect 110 929 116 930
rect 110 925 111 929
rect 115 925 116 929
rect 134 928 135 932
rect 139 928 140 932
rect 134 927 140 928
rect 262 932 268 933
rect 262 928 263 932
rect 267 928 268 932
rect 262 927 268 928
rect 414 932 420 933
rect 414 928 415 932
rect 419 928 420 932
rect 414 927 420 928
rect 558 932 564 933
rect 558 928 559 932
rect 563 928 564 932
rect 558 927 564 928
rect 110 924 116 925
rect 688 924 690 1030
rect 768 1027 770 1037
rect 818 1035 824 1036
rect 818 1031 819 1035
rect 823 1031 824 1035
rect 818 1030 824 1031
rect 766 1026 772 1027
rect 766 1022 767 1026
rect 771 1022 772 1026
rect 766 1021 772 1022
rect 820 1000 822 1030
rect 856 1027 858 1037
rect 934 1035 940 1036
rect 934 1031 935 1035
rect 939 1031 940 1035
rect 934 1030 940 1031
rect 854 1026 860 1027
rect 854 1022 855 1026
rect 859 1022 860 1026
rect 854 1021 860 1022
rect 936 1000 938 1030
rect 944 1027 946 1037
rect 994 1035 1000 1036
rect 994 1031 995 1035
rect 999 1031 1000 1035
rect 994 1030 1000 1031
rect 942 1026 948 1027
rect 942 1022 943 1026
rect 947 1022 948 1026
rect 942 1021 948 1022
rect 996 1000 998 1030
rect 1032 1027 1034 1037
rect 1082 1035 1088 1036
rect 1082 1031 1083 1035
rect 1087 1031 1088 1035
rect 1082 1030 1088 1031
rect 1030 1026 1036 1027
rect 1030 1022 1031 1026
rect 1035 1022 1036 1026
rect 1030 1021 1036 1022
rect 1084 1000 1086 1030
rect 1128 1027 1130 1037
rect 1178 1035 1184 1036
rect 1178 1031 1179 1035
rect 1183 1031 1184 1035
rect 1178 1030 1184 1031
rect 1126 1026 1132 1027
rect 1126 1022 1127 1026
rect 1131 1022 1132 1026
rect 1126 1021 1132 1022
rect 1180 1000 1182 1030
rect 1224 1027 1226 1037
rect 1222 1026 1228 1027
rect 1222 1022 1223 1026
rect 1227 1022 1228 1026
rect 1222 1021 1228 1022
rect 1832 1009 1834 1037
rect 1870 1033 1871 1037
rect 1875 1033 1876 1037
rect 1894 1036 1895 1040
rect 1899 1036 1900 1040
rect 1894 1035 1900 1036
rect 2014 1040 2020 1041
rect 2014 1036 2015 1040
rect 2019 1036 2020 1040
rect 2014 1035 2020 1036
rect 2166 1040 2172 1041
rect 2166 1036 2167 1040
rect 2171 1036 2172 1040
rect 2166 1035 2172 1036
rect 1870 1032 1876 1033
rect 1962 1031 1968 1032
rect 1962 1027 1963 1031
rect 1967 1027 1968 1031
rect 1962 1026 1968 1027
rect 2082 1031 2088 1032
rect 2082 1027 2083 1031
rect 2087 1027 2088 1031
rect 2082 1026 2088 1027
rect 1870 1020 1876 1021
rect 1870 1016 1871 1020
rect 1875 1016 1876 1020
rect 1870 1015 1876 1016
rect 1830 1008 1836 1009
rect 1830 1004 1831 1008
rect 1835 1004 1836 1008
rect 1830 1003 1836 1004
rect 818 999 824 1000
rect 818 995 819 999
rect 823 995 824 999
rect 818 994 824 995
rect 934 999 940 1000
rect 934 995 935 999
rect 939 995 940 999
rect 934 994 940 995
rect 994 999 1000 1000
rect 994 995 995 999
rect 999 995 1000 999
rect 994 994 1000 995
rect 1082 999 1088 1000
rect 1082 995 1083 999
rect 1087 995 1088 999
rect 1082 994 1088 995
rect 1178 999 1184 1000
rect 1178 995 1179 999
rect 1183 995 1184 999
rect 1178 994 1184 995
rect 1830 991 1836 992
rect 758 988 764 989
rect 758 984 759 988
rect 763 984 764 988
rect 758 983 764 984
rect 846 988 852 989
rect 846 984 847 988
rect 851 984 852 988
rect 846 983 852 984
rect 934 988 940 989
rect 934 984 935 988
rect 939 984 940 988
rect 934 983 940 984
rect 1022 988 1028 989
rect 1022 984 1023 988
rect 1027 984 1028 988
rect 1022 983 1028 984
rect 1118 988 1124 989
rect 1118 984 1119 988
rect 1123 984 1124 988
rect 1118 983 1124 984
rect 1214 988 1220 989
rect 1214 984 1215 988
rect 1219 984 1220 988
rect 1830 987 1831 991
rect 1835 987 1836 991
rect 1830 986 1836 987
rect 1214 983 1220 984
rect 760 955 762 983
rect 848 955 850 983
rect 936 955 938 983
rect 1024 955 1026 983
rect 1120 955 1122 983
rect 1216 955 1218 983
rect 1832 955 1834 986
rect 1872 983 1874 1015
rect 1902 1002 1908 1003
rect 1902 998 1903 1002
rect 1907 998 1908 1002
rect 1902 997 1908 998
rect 1904 983 1906 997
rect 1964 992 1966 1026
rect 2022 1002 2028 1003
rect 2022 998 2023 1002
rect 2027 998 2028 1002
rect 2022 997 2028 998
rect 1962 991 1968 992
rect 1962 987 1963 991
rect 1967 987 1968 991
rect 1962 986 1968 987
rect 2024 983 2026 997
rect 2084 992 2086 1026
rect 2174 1002 2180 1003
rect 2174 998 2175 1002
rect 2179 998 2180 1002
rect 2174 997 2180 998
rect 2082 991 2088 992
rect 2082 987 2083 991
rect 2087 987 2088 991
rect 2082 986 2088 987
rect 2176 983 2178 997
rect 2216 992 2218 1090
rect 2350 1084 2356 1085
rect 2350 1080 2351 1084
rect 2355 1080 2356 1084
rect 2350 1079 2356 1080
rect 2566 1084 2572 1085
rect 2566 1080 2567 1084
rect 2571 1080 2572 1084
rect 2566 1079 2572 1080
rect 2766 1084 2772 1085
rect 2766 1080 2767 1084
rect 2771 1080 2772 1084
rect 2766 1079 2772 1080
rect 2958 1084 2964 1085
rect 2958 1080 2959 1084
rect 2963 1080 2964 1084
rect 2958 1079 2964 1080
rect 2352 1063 2354 1079
rect 2568 1063 2570 1079
rect 2768 1063 2770 1079
rect 2960 1063 2962 1079
rect 2327 1062 2331 1063
rect 2327 1057 2331 1058
rect 2351 1062 2355 1063
rect 2351 1057 2355 1058
rect 2487 1062 2491 1063
rect 2487 1057 2491 1058
rect 2567 1062 2571 1063
rect 2567 1057 2571 1058
rect 2639 1062 2643 1063
rect 2639 1057 2643 1058
rect 2767 1062 2771 1063
rect 2767 1057 2771 1058
rect 2791 1062 2795 1063
rect 2791 1057 2795 1058
rect 2935 1062 2939 1063
rect 2935 1057 2939 1058
rect 2959 1062 2963 1063
rect 2959 1057 2963 1058
rect 2328 1041 2330 1057
rect 2488 1041 2490 1057
rect 2640 1041 2642 1057
rect 2792 1041 2794 1057
rect 2936 1041 2938 1057
rect 2326 1040 2332 1041
rect 2326 1036 2327 1040
rect 2331 1036 2332 1040
rect 2326 1035 2332 1036
rect 2486 1040 2492 1041
rect 2486 1036 2487 1040
rect 2491 1036 2492 1040
rect 2486 1035 2492 1036
rect 2638 1040 2644 1041
rect 2638 1036 2639 1040
rect 2643 1036 2644 1040
rect 2638 1035 2644 1036
rect 2790 1040 2796 1041
rect 2790 1036 2791 1040
rect 2795 1036 2796 1040
rect 2790 1035 2796 1036
rect 2934 1040 2940 1041
rect 2934 1036 2935 1040
rect 2939 1036 2940 1040
rect 2934 1035 2940 1036
rect 2414 1031 2420 1032
rect 2414 1027 2415 1031
rect 2419 1027 2420 1031
rect 2414 1026 2420 1027
rect 2706 1031 2712 1032
rect 2706 1027 2707 1031
rect 2711 1027 2712 1031
rect 2706 1026 2712 1027
rect 2858 1031 2864 1032
rect 2858 1027 2859 1031
rect 2863 1027 2864 1031
rect 2858 1026 2864 1027
rect 3002 1031 3008 1032
rect 3002 1027 3003 1031
rect 3007 1027 3008 1031
rect 3002 1026 3008 1027
rect 2334 1002 2340 1003
rect 2334 998 2335 1002
rect 2339 998 2340 1002
rect 2334 997 2340 998
rect 2206 991 2212 992
rect 2206 987 2207 991
rect 2211 987 2212 991
rect 2206 986 2212 987
rect 2214 991 2220 992
rect 2214 987 2215 991
rect 2219 987 2220 991
rect 2214 986 2220 987
rect 1871 982 1875 983
rect 1871 977 1875 978
rect 1903 982 1907 983
rect 1903 977 1907 978
rect 1983 982 1987 983
rect 1983 977 1987 978
rect 2023 982 2027 983
rect 2023 977 2027 978
rect 2079 982 2083 983
rect 2079 977 2083 978
rect 2175 982 2179 983
rect 2175 977 2179 978
rect 2199 982 2203 983
rect 2199 977 2203 978
rect 703 954 707 955
rect 703 949 707 950
rect 759 954 763 955
rect 759 949 763 950
rect 839 954 843 955
rect 839 949 843 950
rect 847 954 851 955
rect 847 949 851 950
rect 935 954 939 955
rect 935 949 939 950
rect 975 954 979 955
rect 975 949 979 950
rect 1023 954 1027 955
rect 1023 949 1027 950
rect 1103 954 1107 955
rect 1103 949 1107 950
rect 1119 954 1123 955
rect 1119 949 1123 950
rect 1215 954 1219 955
rect 1215 949 1219 950
rect 1223 954 1227 955
rect 1223 949 1227 950
rect 1335 954 1339 955
rect 1335 949 1339 950
rect 1439 954 1443 955
rect 1439 949 1443 950
rect 1543 954 1547 955
rect 1543 949 1547 950
rect 1655 954 1659 955
rect 1655 949 1659 950
rect 1743 954 1747 955
rect 1743 949 1747 950
rect 1831 954 1835 955
rect 1831 949 1835 950
rect 1872 949 1874 977
rect 1904 967 1906 977
rect 1954 975 1960 976
rect 1954 971 1955 975
rect 1959 971 1960 975
rect 1954 970 1960 971
rect 1902 966 1908 967
rect 1902 962 1903 966
rect 1907 962 1908 966
rect 1902 961 1908 962
rect 704 933 706 949
rect 840 933 842 949
rect 976 933 978 949
rect 1104 933 1106 949
rect 1224 933 1226 949
rect 1336 933 1338 949
rect 1440 933 1442 949
rect 1544 933 1546 949
rect 1656 933 1658 949
rect 1744 933 1746 949
rect 702 932 708 933
rect 702 928 703 932
rect 707 928 708 932
rect 702 927 708 928
rect 838 932 844 933
rect 838 928 839 932
rect 843 928 844 932
rect 838 927 844 928
rect 974 932 980 933
rect 974 928 975 932
rect 979 928 980 932
rect 974 927 980 928
rect 1102 932 1108 933
rect 1102 928 1103 932
rect 1107 928 1108 932
rect 1102 927 1108 928
rect 1222 932 1228 933
rect 1222 928 1223 932
rect 1227 928 1228 932
rect 1222 927 1228 928
rect 1334 932 1340 933
rect 1334 928 1335 932
rect 1339 928 1340 932
rect 1334 927 1340 928
rect 1438 932 1444 933
rect 1438 928 1439 932
rect 1443 928 1444 932
rect 1438 927 1444 928
rect 1542 932 1548 933
rect 1542 928 1543 932
rect 1547 928 1548 932
rect 1542 927 1548 928
rect 1654 932 1660 933
rect 1654 928 1655 932
rect 1659 928 1660 932
rect 1654 927 1660 928
rect 1742 932 1748 933
rect 1742 928 1743 932
rect 1747 928 1748 932
rect 1832 930 1834 949
rect 1870 948 1876 949
rect 1870 944 1871 948
rect 1875 944 1876 948
rect 1870 943 1876 944
rect 1956 940 1958 970
rect 1984 967 1986 977
rect 2034 975 2040 976
rect 2034 971 2035 975
rect 2039 971 2040 975
rect 2034 970 2040 971
rect 1982 966 1988 967
rect 1982 962 1983 966
rect 1987 962 1988 966
rect 1982 961 1988 962
rect 2036 940 2038 970
rect 2080 967 2082 977
rect 2130 975 2136 976
rect 2130 971 2131 975
rect 2135 971 2136 975
rect 2130 970 2136 971
rect 2078 966 2084 967
rect 2078 962 2079 966
rect 2083 962 2084 966
rect 2078 961 2084 962
rect 2132 940 2134 970
rect 2200 967 2202 977
rect 2198 966 2204 967
rect 2198 962 2199 966
rect 2203 962 2204 966
rect 2198 961 2204 962
rect 2208 940 2210 986
rect 2336 983 2338 997
rect 2416 992 2418 1026
rect 2494 1002 2500 1003
rect 2494 998 2495 1002
rect 2499 998 2500 1002
rect 2494 997 2500 998
rect 2646 1002 2652 1003
rect 2646 998 2647 1002
rect 2651 998 2652 1002
rect 2646 997 2652 998
rect 2414 991 2420 992
rect 2414 987 2415 991
rect 2419 987 2420 991
rect 2414 986 2420 987
rect 2496 983 2498 997
rect 2648 983 2650 997
rect 2708 992 2710 1026
rect 2798 1002 2804 1003
rect 2798 998 2799 1002
rect 2803 998 2804 1002
rect 2798 997 2804 998
rect 2706 991 2712 992
rect 2706 987 2707 991
rect 2711 987 2712 991
rect 2706 986 2712 987
rect 2800 983 2802 997
rect 2860 992 2862 1026
rect 2942 1002 2948 1003
rect 2942 998 2943 1002
rect 2947 998 2948 1002
rect 2942 997 2948 998
rect 2858 991 2864 992
rect 2858 987 2859 991
rect 2863 987 2864 991
rect 2858 986 2864 987
rect 2944 983 2946 997
rect 3004 992 3006 1026
rect 3020 992 3022 1090
rect 3150 1084 3156 1085
rect 3150 1080 3151 1084
rect 3155 1080 3156 1084
rect 3150 1079 3156 1080
rect 3152 1063 3154 1079
rect 3079 1062 3083 1063
rect 3079 1057 3083 1058
rect 3151 1062 3155 1063
rect 3151 1057 3155 1058
rect 3080 1041 3082 1057
rect 3078 1040 3084 1041
rect 3078 1036 3079 1040
rect 3083 1036 3084 1040
rect 3078 1035 3084 1036
rect 3086 1002 3092 1003
rect 3086 998 3087 1002
rect 3091 998 3092 1002
rect 3086 997 3092 998
rect 3002 991 3008 992
rect 3002 987 3003 991
rect 3007 987 3008 991
rect 3002 986 3008 987
rect 3018 991 3024 992
rect 3018 987 3019 991
rect 3023 987 3024 991
rect 3018 986 3024 987
rect 3088 983 3090 997
rect 3212 992 3214 1090
rect 3590 1087 3596 1088
rect 3334 1084 3340 1085
rect 3334 1080 3335 1084
rect 3339 1080 3340 1084
rect 3334 1079 3340 1080
rect 3502 1084 3508 1085
rect 3502 1080 3503 1084
rect 3507 1080 3508 1084
rect 3590 1083 3591 1087
rect 3595 1083 3596 1087
rect 3590 1082 3596 1083
rect 3502 1079 3508 1080
rect 3336 1063 3338 1079
rect 3504 1063 3506 1079
rect 3592 1063 3594 1082
rect 3223 1062 3227 1063
rect 3223 1057 3227 1058
rect 3335 1062 3339 1063
rect 3335 1057 3339 1058
rect 3375 1062 3379 1063
rect 3375 1057 3379 1058
rect 3503 1062 3507 1063
rect 3503 1057 3507 1058
rect 3591 1062 3595 1063
rect 3591 1057 3595 1058
rect 3224 1041 3226 1057
rect 3376 1041 3378 1057
rect 3504 1041 3506 1057
rect 3222 1040 3228 1041
rect 3222 1036 3223 1040
rect 3227 1036 3228 1040
rect 3222 1035 3228 1036
rect 3374 1040 3380 1041
rect 3374 1036 3375 1040
rect 3379 1036 3380 1040
rect 3374 1035 3380 1036
rect 3502 1040 3508 1041
rect 3502 1036 3503 1040
rect 3507 1036 3508 1040
rect 3592 1038 3594 1057
rect 3502 1035 3508 1036
rect 3590 1037 3596 1038
rect 3590 1033 3591 1037
rect 3595 1033 3596 1037
rect 3590 1032 3596 1033
rect 3306 1031 3312 1032
rect 3306 1027 3307 1031
rect 3311 1027 3312 1031
rect 3306 1026 3312 1027
rect 3230 1002 3236 1003
rect 3230 998 3231 1002
rect 3235 998 3236 1002
rect 3230 997 3236 998
rect 3210 991 3216 992
rect 3210 987 3211 991
rect 3215 987 3216 991
rect 3210 986 3216 987
rect 3232 983 3234 997
rect 3308 992 3310 1026
rect 3590 1020 3596 1021
rect 3590 1016 3591 1020
rect 3595 1016 3596 1020
rect 3590 1015 3596 1016
rect 3382 1002 3388 1003
rect 3382 998 3383 1002
rect 3387 998 3388 1002
rect 3382 997 3388 998
rect 3510 1002 3516 1003
rect 3510 998 3511 1002
rect 3515 998 3516 1002
rect 3510 997 3516 998
rect 3306 991 3312 992
rect 3306 987 3307 991
rect 3311 987 3312 991
rect 3306 986 3312 987
rect 3384 983 3386 997
rect 3512 983 3514 997
rect 3518 991 3524 992
rect 3518 987 3519 991
rect 3523 987 3524 991
rect 3518 986 3524 987
rect 2335 982 2339 983
rect 2335 977 2339 978
rect 2479 982 2483 983
rect 2479 977 2483 978
rect 2495 982 2499 983
rect 2495 977 2499 978
rect 2631 982 2635 983
rect 2631 977 2635 978
rect 2647 982 2651 983
rect 2647 977 2651 978
rect 2791 982 2795 983
rect 2791 977 2795 978
rect 2799 982 2803 983
rect 2799 977 2803 978
rect 2943 982 2947 983
rect 2943 977 2947 978
rect 2967 982 2971 983
rect 2967 977 2971 978
rect 3087 982 3091 983
rect 3087 977 3091 978
rect 3151 982 3155 983
rect 3151 977 3155 978
rect 3231 982 3235 983
rect 3231 977 3235 978
rect 3343 982 3347 983
rect 3343 977 3347 978
rect 3383 982 3387 983
rect 3383 977 3387 978
rect 3511 982 3515 983
rect 3511 977 3515 978
rect 2336 967 2338 977
rect 2406 975 2412 976
rect 2406 971 2407 975
rect 2411 971 2412 975
rect 2406 970 2412 971
rect 2334 966 2340 967
rect 2334 962 2335 966
rect 2339 962 2340 966
rect 2334 961 2340 962
rect 2408 940 2410 970
rect 2480 967 2482 977
rect 2632 967 2634 977
rect 2682 975 2688 976
rect 2682 971 2683 975
rect 2687 971 2688 975
rect 2682 970 2688 971
rect 2478 966 2484 967
rect 2478 962 2479 966
rect 2483 962 2484 966
rect 2478 961 2484 962
rect 2630 966 2636 967
rect 2630 962 2631 966
rect 2635 962 2636 966
rect 2630 961 2636 962
rect 2684 940 2686 970
rect 2792 967 2794 977
rect 2842 975 2848 976
rect 2842 971 2843 975
rect 2847 971 2848 975
rect 2842 970 2848 971
rect 2790 966 2796 967
rect 2790 962 2791 966
rect 2795 962 2796 966
rect 2790 961 2796 962
rect 2844 940 2846 970
rect 2968 967 2970 977
rect 3152 967 3154 977
rect 3210 975 3216 976
rect 3210 971 3211 975
rect 3215 971 3216 975
rect 3210 970 3216 971
rect 2966 966 2972 967
rect 2966 962 2967 966
rect 2971 962 2972 966
rect 2966 961 2972 962
rect 3150 966 3156 967
rect 3150 962 3151 966
rect 3155 962 3156 966
rect 3150 961 3156 962
rect 3212 940 3214 970
rect 3344 967 3346 977
rect 3512 967 3514 977
rect 3342 966 3348 967
rect 3342 962 3343 966
rect 3347 962 3348 966
rect 3342 961 3348 962
rect 3510 966 3516 967
rect 3510 962 3511 966
rect 3515 962 3516 966
rect 3510 961 3516 962
rect 3520 940 3522 986
rect 3592 983 3594 1015
rect 3591 982 3595 983
rect 3591 977 3595 978
rect 3592 949 3594 977
rect 3590 948 3596 949
rect 3590 944 3591 948
rect 3595 944 3596 948
rect 3590 943 3596 944
rect 1954 939 1960 940
rect 1954 935 1955 939
rect 1959 935 1960 939
rect 1954 934 1960 935
rect 2034 939 2040 940
rect 2034 935 2035 939
rect 2039 935 2040 939
rect 2034 934 2040 935
rect 2130 939 2136 940
rect 2130 935 2131 939
rect 2135 935 2136 939
rect 2130 934 2136 935
rect 2206 939 2212 940
rect 2206 935 2207 939
rect 2211 935 2212 939
rect 2206 934 2212 935
rect 2406 939 2412 940
rect 2406 935 2407 939
rect 2411 935 2412 939
rect 2406 934 2412 935
rect 2682 939 2688 940
rect 2682 935 2683 939
rect 2687 935 2688 939
rect 2682 934 2688 935
rect 2842 939 2848 940
rect 2842 935 2843 939
rect 2847 935 2848 939
rect 2842 934 2848 935
rect 3202 939 3208 940
rect 3202 935 3203 939
rect 3207 935 3208 939
rect 3202 934 3208 935
rect 3210 939 3216 940
rect 3210 935 3211 939
rect 3215 935 3216 939
rect 3210 934 3216 935
rect 3518 939 3524 940
rect 3518 935 3519 939
rect 3523 935 3524 939
rect 3518 934 3524 935
rect 1870 931 1876 932
rect 1742 927 1748 928
rect 1830 929 1836 930
rect 1830 925 1831 929
rect 1835 925 1836 929
rect 1870 927 1871 931
rect 1875 927 1876 931
rect 1870 926 1876 927
rect 1894 928 1900 929
rect 1830 924 1836 925
rect 338 923 344 924
rect 338 919 339 923
rect 343 919 344 923
rect 338 918 344 919
rect 494 923 500 924
rect 494 919 495 923
rect 499 919 500 923
rect 494 918 500 919
rect 634 923 640 924
rect 634 919 635 923
rect 639 919 640 923
rect 634 918 640 919
rect 686 923 692 924
rect 686 919 687 923
rect 691 919 692 923
rect 686 918 692 919
rect 778 923 784 924
rect 778 919 779 923
rect 783 919 784 923
rect 778 918 784 919
rect 1042 923 1048 924
rect 1042 919 1043 923
rect 1047 919 1048 923
rect 1042 918 1048 919
rect 1170 923 1176 924
rect 1170 919 1171 923
rect 1175 919 1176 923
rect 1170 918 1176 919
rect 1402 923 1408 924
rect 1402 919 1403 923
rect 1407 919 1408 923
rect 1402 918 1408 919
rect 1506 923 1512 924
rect 1506 919 1507 923
rect 1511 919 1512 923
rect 1506 918 1512 919
rect 1610 923 1616 924
rect 1610 919 1611 923
rect 1615 919 1616 923
rect 1610 918 1616 919
rect 1722 923 1728 924
rect 1722 919 1723 923
rect 1727 919 1728 923
rect 1722 918 1728 919
rect 1742 919 1748 920
rect 110 912 116 913
rect 110 908 111 912
rect 115 908 116 912
rect 110 907 116 908
rect 112 875 114 907
rect 142 894 148 895
rect 142 890 143 894
rect 147 890 148 894
rect 142 889 148 890
rect 270 894 276 895
rect 270 890 271 894
rect 275 890 276 894
rect 270 889 276 890
rect 144 875 146 889
rect 150 883 156 884
rect 150 879 151 883
rect 155 879 156 883
rect 150 878 156 879
rect 111 874 115 875
rect 111 869 115 870
rect 143 874 147 875
rect 143 869 147 870
rect 112 841 114 869
rect 144 859 146 869
rect 142 858 148 859
rect 142 854 143 858
rect 147 854 148 858
rect 142 853 148 854
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 152 832 154 878
rect 272 875 274 889
rect 340 884 342 918
rect 422 894 428 895
rect 422 890 423 894
rect 427 890 428 894
rect 422 889 428 890
rect 338 883 344 884
rect 338 879 339 883
rect 343 879 344 883
rect 338 878 344 879
rect 424 875 426 889
rect 496 884 498 918
rect 566 894 572 895
rect 566 890 567 894
rect 571 890 572 894
rect 566 889 572 890
rect 494 883 500 884
rect 494 879 495 883
rect 499 879 500 883
rect 494 878 500 879
rect 568 875 570 889
rect 247 874 251 875
rect 247 869 251 870
rect 271 874 275 875
rect 271 869 275 870
rect 383 874 387 875
rect 383 869 387 870
rect 423 874 427 875
rect 423 869 427 870
rect 519 874 523 875
rect 519 869 523 870
rect 567 874 571 875
rect 567 869 571 870
rect 202 867 208 868
rect 202 863 203 867
rect 207 863 208 867
rect 202 862 208 863
rect 204 832 206 862
rect 248 859 250 869
rect 258 867 264 868
rect 258 863 259 867
rect 263 863 264 867
rect 258 862 264 863
rect 366 867 372 868
rect 366 863 367 867
rect 371 863 372 867
rect 366 862 372 863
rect 246 858 252 859
rect 246 854 247 858
rect 251 854 252 858
rect 246 853 252 854
rect 260 845 262 862
rect 259 844 263 845
rect 259 839 263 840
rect 150 831 156 832
rect 150 827 151 831
rect 155 827 156 831
rect 150 826 156 827
rect 202 831 208 832
rect 202 827 203 831
rect 207 827 208 831
rect 202 826 208 827
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 110 818 116 819
rect 134 820 140 821
rect 112 787 114 818
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 238 820 244 821
rect 238 816 239 820
rect 243 816 244 820
rect 238 815 244 816
rect 136 787 138 815
rect 240 787 242 815
rect 111 786 115 787
rect 111 781 115 782
rect 135 786 139 787
rect 135 781 139 782
rect 215 786 219 787
rect 215 781 219 782
rect 239 786 243 787
rect 239 781 243 782
rect 303 786 307 787
rect 303 781 307 782
rect 112 762 114 781
rect 136 765 138 781
rect 216 765 218 781
rect 304 765 306 781
rect 134 764 140 765
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 134 760 135 764
rect 139 760 140 764
rect 134 759 140 760
rect 214 764 220 765
rect 214 760 215 764
rect 219 760 220 764
rect 214 759 220 760
rect 302 764 308 765
rect 302 760 303 764
rect 307 760 308 764
rect 302 759 308 760
rect 110 756 116 757
rect 368 756 370 862
rect 384 859 386 869
rect 434 867 440 868
rect 434 863 435 867
rect 439 863 440 867
rect 434 862 440 863
rect 382 858 388 859
rect 382 854 383 858
rect 387 854 388 858
rect 382 853 388 854
rect 436 832 438 862
rect 520 859 522 869
rect 636 868 638 918
rect 710 894 716 895
rect 710 890 711 894
rect 715 890 716 894
rect 710 889 716 890
rect 712 875 714 889
rect 780 884 782 918
rect 846 894 852 895
rect 846 890 847 894
rect 851 890 852 894
rect 846 889 852 890
rect 982 894 988 895
rect 982 890 983 894
rect 987 890 988 894
rect 982 889 988 890
rect 778 883 784 884
rect 778 879 779 883
rect 783 879 784 883
rect 778 878 784 879
rect 838 883 844 884
rect 838 879 839 883
rect 843 879 844 883
rect 838 878 844 879
rect 663 874 667 875
rect 663 869 667 870
rect 711 874 715 875
rect 711 869 715 870
rect 815 874 819 875
rect 815 869 819 870
rect 634 867 640 868
rect 634 863 635 867
rect 639 863 640 867
rect 634 862 640 863
rect 664 859 666 869
rect 816 859 818 869
rect 518 858 524 859
rect 518 854 519 858
rect 523 854 524 858
rect 518 853 524 854
rect 662 858 668 859
rect 662 854 663 858
rect 667 854 668 858
rect 662 853 668 854
rect 814 858 820 859
rect 814 854 815 858
rect 819 854 820 858
rect 814 853 820 854
rect 527 844 531 845
rect 527 839 531 840
rect 528 832 530 839
rect 840 832 842 878
rect 848 875 850 889
rect 984 875 986 889
rect 1044 884 1046 918
rect 1110 894 1116 895
rect 1110 890 1111 894
rect 1115 890 1116 894
rect 1110 889 1116 890
rect 1042 883 1048 884
rect 1042 879 1043 883
rect 1047 879 1048 883
rect 1042 878 1048 879
rect 1112 875 1114 889
rect 1172 884 1174 918
rect 1230 894 1236 895
rect 1230 890 1231 894
rect 1235 890 1236 894
rect 1230 889 1236 890
rect 1342 894 1348 895
rect 1342 890 1343 894
rect 1347 890 1348 894
rect 1342 889 1348 890
rect 1170 883 1176 884
rect 1170 879 1171 883
rect 1175 879 1176 883
rect 1170 878 1176 879
rect 1232 875 1234 889
rect 1344 875 1346 889
rect 1404 884 1406 918
rect 1446 894 1452 895
rect 1446 890 1447 894
rect 1451 890 1452 894
rect 1446 889 1452 890
rect 1390 883 1396 884
rect 1390 879 1391 883
rect 1395 879 1396 883
rect 1390 878 1396 879
rect 1402 883 1408 884
rect 1402 879 1403 883
rect 1407 879 1408 883
rect 1402 878 1408 879
rect 847 874 851 875
rect 847 869 851 870
rect 959 874 963 875
rect 959 869 963 870
rect 983 874 987 875
rect 983 869 987 870
rect 1103 874 1107 875
rect 1103 869 1107 870
rect 1111 874 1115 875
rect 1111 869 1115 870
rect 1231 874 1235 875
rect 1231 869 1235 870
rect 1247 874 1251 875
rect 1247 869 1251 870
rect 1343 874 1347 875
rect 1343 869 1347 870
rect 1383 874 1387 875
rect 1383 869 1387 870
rect 960 859 962 869
rect 1010 867 1016 868
rect 1010 863 1011 867
rect 1015 863 1016 867
rect 1010 862 1016 863
rect 958 858 964 859
rect 958 854 959 858
rect 963 854 964 858
rect 958 853 964 854
rect 1012 832 1014 862
rect 1104 859 1106 869
rect 1154 867 1160 868
rect 1154 863 1155 867
rect 1159 863 1160 867
rect 1154 862 1160 863
rect 1102 858 1108 859
rect 1102 854 1103 858
rect 1107 854 1108 858
rect 1102 853 1108 854
rect 1156 832 1158 862
rect 1248 859 1250 869
rect 1384 859 1386 869
rect 1246 858 1252 859
rect 1246 854 1247 858
rect 1251 854 1252 858
rect 1246 853 1252 854
rect 1382 858 1388 859
rect 1382 854 1383 858
rect 1387 854 1388 858
rect 1382 853 1388 854
rect 1392 832 1394 878
rect 1448 875 1450 889
rect 1508 884 1510 918
rect 1550 894 1556 895
rect 1550 890 1551 894
rect 1555 890 1556 894
rect 1550 889 1556 890
rect 1506 883 1512 884
rect 1506 879 1507 883
rect 1511 879 1512 883
rect 1506 878 1512 879
rect 1552 875 1554 889
rect 1612 884 1614 918
rect 1662 894 1668 895
rect 1662 890 1663 894
rect 1667 890 1668 894
rect 1662 889 1668 890
rect 1610 883 1616 884
rect 1610 879 1611 883
rect 1615 879 1616 883
rect 1610 878 1616 879
rect 1646 875 1652 876
rect 1664 875 1666 889
rect 1724 884 1726 918
rect 1742 915 1743 919
rect 1747 915 1748 919
rect 1742 914 1748 915
rect 1722 883 1728 884
rect 1722 879 1723 883
rect 1727 879 1728 883
rect 1722 878 1728 879
rect 1447 874 1451 875
rect 1447 869 1451 870
rect 1511 874 1515 875
rect 1511 869 1515 870
rect 1551 874 1555 875
rect 1551 869 1555 870
rect 1639 874 1643 875
rect 1646 871 1647 875
rect 1651 871 1652 875
rect 1646 870 1652 871
rect 1663 874 1667 875
rect 1639 869 1643 870
rect 1512 859 1514 869
rect 1518 867 1524 868
rect 1518 863 1519 867
rect 1523 863 1524 867
rect 1518 862 1524 863
rect 1562 867 1568 868
rect 1562 863 1563 867
rect 1567 863 1568 867
rect 1562 862 1568 863
rect 1510 858 1516 859
rect 1510 854 1511 858
rect 1515 854 1516 858
rect 1510 853 1516 854
rect 434 831 440 832
rect 434 827 435 831
rect 439 827 440 831
rect 434 826 440 827
rect 526 831 532 832
rect 526 827 527 831
rect 531 827 532 831
rect 526 826 532 827
rect 838 831 844 832
rect 838 827 839 831
rect 843 827 844 831
rect 838 826 844 827
rect 1010 831 1016 832
rect 1010 827 1011 831
rect 1015 827 1016 831
rect 1010 826 1016 827
rect 1154 831 1160 832
rect 1154 827 1155 831
rect 1159 827 1160 831
rect 1154 826 1160 827
rect 1390 831 1396 832
rect 1390 827 1391 831
rect 1395 827 1396 831
rect 1390 826 1396 827
rect 374 820 380 821
rect 374 816 375 820
rect 379 816 380 820
rect 374 815 380 816
rect 510 820 516 821
rect 510 816 511 820
rect 515 816 516 820
rect 510 815 516 816
rect 654 820 660 821
rect 654 816 655 820
rect 659 816 660 820
rect 654 815 660 816
rect 806 820 812 821
rect 806 816 807 820
rect 811 816 812 820
rect 806 815 812 816
rect 950 820 956 821
rect 950 816 951 820
rect 955 816 956 820
rect 950 815 956 816
rect 1094 820 1100 821
rect 1094 816 1095 820
rect 1099 816 1100 820
rect 1094 815 1100 816
rect 1238 820 1244 821
rect 1238 816 1239 820
rect 1243 816 1244 820
rect 1238 815 1244 816
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1502 820 1508 821
rect 1502 816 1503 820
rect 1507 816 1508 820
rect 1502 815 1508 816
rect 376 787 378 815
rect 512 787 514 815
rect 656 787 658 815
rect 808 787 810 815
rect 952 787 954 815
rect 1096 787 1098 815
rect 1158 803 1164 804
rect 1158 799 1159 803
rect 1163 799 1164 803
rect 1158 798 1164 799
rect 375 786 379 787
rect 375 781 379 782
rect 415 786 419 787
rect 415 781 419 782
rect 511 786 515 787
rect 511 781 515 782
rect 543 786 547 787
rect 543 781 547 782
rect 655 786 659 787
rect 655 781 659 782
rect 687 786 691 787
rect 687 781 691 782
rect 807 786 811 787
rect 807 781 811 782
rect 839 786 843 787
rect 839 781 843 782
rect 951 786 955 787
rect 951 781 955 782
rect 991 786 995 787
rect 991 781 995 782
rect 1095 786 1099 787
rect 1095 781 1099 782
rect 1143 786 1147 787
rect 1143 781 1147 782
rect 416 765 418 781
rect 544 765 546 781
rect 688 765 690 781
rect 840 765 842 781
rect 992 765 994 781
rect 1144 765 1146 781
rect 414 764 420 765
rect 414 760 415 764
rect 419 760 420 764
rect 414 759 420 760
rect 542 764 548 765
rect 542 760 543 764
rect 547 760 548 764
rect 542 759 548 760
rect 686 764 692 765
rect 686 760 687 764
rect 691 760 692 764
rect 686 759 692 760
rect 838 764 844 765
rect 838 760 839 764
rect 843 760 844 764
rect 838 759 844 760
rect 990 764 996 765
rect 990 760 991 764
rect 995 760 996 764
rect 990 759 996 760
rect 1142 764 1148 765
rect 1142 760 1143 764
rect 1147 760 1148 764
rect 1142 759 1148 760
rect 202 755 208 756
rect 202 751 203 755
rect 207 751 208 755
rect 202 750 208 751
rect 282 755 288 756
rect 282 751 283 755
rect 287 751 288 755
rect 368 755 376 756
rect 368 752 371 755
rect 282 750 288 751
rect 370 751 371 752
rect 375 751 376 755
rect 370 750 376 751
rect 486 755 492 756
rect 486 751 487 755
rect 491 751 492 755
rect 486 750 492 751
rect 610 755 616 756
rect 610 751 611 755
rect 615 751 616 755
rect 610 750 616 751
rect 654 755 660 756
rect 654 751 655 755
rect 659 751 660 755
rect 654 750 660 751
rect 906 755 912 756
rect 906 751 907 755
rect 911 751 912 755
rect 906 750 912 751
rect 914 755 920 756
rect 914 751 915 755
rect 919 751 920 755
rect 914 750 920 751
rect 1058 755 1064 756
rect 1058 751 1059 755
rect 1063 751 1064 755
rect 1058 750 1064 751
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 112 703 114 739
rect 142 726 148 727
rect 142 722 143 726
rect 147 722 148 726
rect 142 721 148 722
rect 151 724 155 725
rect 144 703 146 721
rect 151 719 155 720
rect 152 716 154 719
rect 204 716 206 750
rect 222 726 228 727
rect 222 722 223 726
rect 227 722 228 726
rect 222 721 228 722
rect 150 715 156 716
rect 150 711 151 715
rect 155 711 156 715
rect 150 710 156 711
rect 202 715 208 716
rect 202 711 203 715
rect 207 711 208 715
rect 202 710 208 711
rect 224 703 226 721
rect 284 716 286 750
rect 310 726 316 727
rect 310 722 311 726
rect 315 722 316 726
rect 310 721 316 722
rect 422 726 428 727
rect 422 722 423 726
rect 427 722 428 726
rect 422 721 428 722
rect 282 715 288 716
rect 282 711 283 715
rect 287 711 288 715
rect 282 710 288 711
rect 312 703 314 721
rect 424 703 426 721
rect 488 716 490 750
rect 550 726 556 727
rect 550 722 551 726
rect 555 722 556 726
rect 550 721 556 722
rect 430 715 436 716
rect 430 711 431 715
rect 435 711 436 715
rect 430 710 436 711
rect 486 715 492 716
rect 486 711 487 715
rect 491 711 492 715
rect 486 710 492 711
rect 111 702 115 703
rect 111 697 115 698
rect 143 702 147 703
rect 143 697 147 698
rect 223 702 227 703
rect 223 697 227 698
rect 231 702 235 703
rect 231 697 235 698
rect 311 702 315 703
rect 311 697 315 698
rect 319 702 323 703
rect 319 697 323 698
rect 423 702 427 703
rect 423 697 427 698
rect 112 669 114 697
rect 232 687 234 697
rect 274 695 280 696
rect 274 691 275 695
rect 279 691 280 695
rect 274 690 280 691
rect 282 695 288 696
rect 282 691 283 695
rect 287 691 288 695
rect 282 690 288 691
rect 230 686 236 687
rect 230 682 231 686
rect 235 682 236 686
rect 276 685 278 690
rect 230 681 236 682
rect 275 684 279 685
rect 275 679 279 680
rect 110 668 116 669
rect 110 664 111 668
rect 115 664 116 668
rect 110 663 116 664
rect 284 660 286 690
rect 320 687 322 697
rect 370 695 376 696
rect 370 691 371 695
rect 375 691 376 695
rect 370 690 376 691
rect 318 686 324 687
rect 318 682 319 686
rect 323 682 324 686
rect 318 681 324 682
rect 372 660 374 690
rect 424 687 426 697
rect 422 686 428 687
rect 422 682 423 686
rect 427 682 428 686
rect 422 681 428 682
rect 432 660 434 710
rect 552 703 554 721
rect 612 716 614 750
rect 656 725 658 750
rect 694 726 700 727
rect 655 724 659 725
rect 694 722 695 726
rect 699 722 700 726
rect 694 721 700 722
rect 846 726 852 727
rect 846 722 847 726
rect 851 722 852 726
rect 846 721 852 722
rect 655 719 659 720
rect 610 715 616 716
rect 610 711 611 715
rect 615 711 616 715
rect 610 710 616 711
rect 696 703 698 721
rect 848 703 850 721
rect 543 702 547 703
rect 543 697 547 698
rect 551 702 555 703
rect 551 697 555 698
rect 679 702 683 703
rect 679 697 683 698
rect 695 702 699 703
rect 695 697 699 698
rect 815 702 819 703
rect 815 697 819 698
rect 847 702 851 703
rect 847 697 851 698
rect 544 687 546 697
rect 602 695 608 696
rect 602 691 603 695
rect 607 691 608 695
rect 602 690 608 691
rect 542 686 548 687
rect 542 682 543 686
rect 547 682 548 686
rect 542 681 548 682
rect 551 684 555 685
rect 551 679 555 680
rect 552 660 554 679
rect 604 660 606 690
rect 680 687 682 697
rect 738 695 744 696
rect 738 691 739 695
rect 743 691 744 695
rect 738 690 744 691
rect 678 686 684 687
rect 678 682 679 686
rect 683 682 684 686
rect 678 681 684 682
rect 740 660 742 690
rect 816 687 818 697
rect 908 696 910 750
rect 916 716 918 750
rect 998 726 1004 727
rect 998 722 999 726
rect 1003 722 1004 726
rect 998 721 1004 722
rect 914 715 920 716
rect 914 711 915 715
rect 919 711 920 715
rect 914 710 920 711
rect 1000 703 1002 721
rect 1060 716 1062 750
rect 1150 726 1156 727
rect 1150 722 1151 726
rect 1155 722 1156 726
rect 1150 721 1156 722
rect 1058 715 1064 716
rect 1058 711 1059 715
rect 1063 711 1064 715
rect 1058 710 1064 711
rect 1152 703 1154 721
rect 1160 716 1162 798
rect 1240 787 1242 815
rect 1376 787 1378 815
rect 1504 787 1506 815
rect 1239 786 1243 787
rect 1239 781 1243 782
rect 1295 786 1299 787
rect 1295 781 1299 782
rect 1375 786 1379 787
rect 1375 781 1379 782
rect 1447 786 1451 787
rect 1447 781 1451 782
rect 1503 786 1507 787
rect 1503 781 1507 782
rect 1296 765 1298 781
rect 1448 765 1450 781
rect 1294 764 1300 765
rect 1294 760 1295 764
rect 1299 760 1300 764
rect 1294 759 1300 760
rect 1446 764 1452 765
rect 1446 760 1447 764
rect 1451 760 1452 764
rect 1446 759 1452 760
rect 1520 756 1522 862
rect 1564 832 1566 862
rect 1640 859 1642 869
rect 1638 858 1644 859
rect 1638 854 1639 858
rect 1643 854 1644 858
rect 1638 853 1644 854
rect 1648 832 1650 870
rect 1663 869 1667 870
rect 1744 868 1746 914
rect 1830 912 1836 913
rect 1830 908 1831 912
rect 1835 908 1836 912
rect 1830 907 1836 908
rect 1750 894 1756 895
rect 1750 890 1751 894
rect 1755 890 1756 894
rect 1750 889 1756 890
rect 1752 875 1754 889
rect 1832 875 1834 907
rect 1872 895 1874 926
rect 1894 924 1895 928
rect 1899 924 1900 928
rect 1894 923 1900 924
rect 1974 928 1980 929
rect 1974 924 1975 928
rect 1979 924 1980 928
rect 1974 923 1980 924
rect 2070 928 2076 929
rect 2070 924 2071 928
rect 2075 924 2076 928
rect 2070 923 2076 924
rect 2190 928 2196 929
rect 2190 924 2191 928
rect 2195 924 2196 928
rect 2190 923 2196 924
rect 2326 928 2332 929
rect 2326 924 2327 928
rect 2331 924 2332 928
rect 2326 923 2332 924
rect 2470 928 2476 929
rect 2470 924 2471 928
rect 2475 924 2476 928
rect 2470 923 2476 924
rect 2622 928 2628 929
rect 2622 924 2623 928
rect 2627 924 2628 928
rect 2622 923 2628 924
rect 2782 928 2788 929
rect 2782 924 2783 928
rect 2787 924 2788 928
rect 2782 923 2788 924
rect 2958 928 2964 929
rect 2958 924 2959 928
rect 2963 924 2964 928
rect 2958 923 2964 924
rect 3142 928 3148 929
rect 3142 924 3143 928
rect 3147 924 3148 928
rect 3142 923 3148 924
rect 1896 895 1898 923
rect 1976 895 1978 923
rect 2072 895 2074 923
rect 2192 895 2194 923
rect 2310 911 2316 912
rect 2310 907 2311 911
rect 2315 907 2316 911
rect 2310 906 2316 907
rect 1871 894 1875 895
rect 1871 889 1875 890
rect 1895 894 1899 895
rect 1895 889 1899 890
rect 1919 894 1923 895
rect 1919 889 1923 890
rect 1975 894 1979 895
rect 1975 889 1979 890
rect 2071 894 2075 895
rect 2071 889 2075 890
rect 2095 894 2099 895
rect 2095 889 2099 890
rect 2191 894 2195 895
rect 2191 889 2195 890
rect 2271 894 2275 895
rect 2271 889 2275 890
rect 1751 874 1755 875
rect 1751 869 1755 870
rect 1831 874 1835 875
rect 1872 870 1874 889
rect 1920 873 1922 889
rect 2096 873 2098 889
rect 2272 873 2274 889
rect 1918 872 1924 873
rect 1831 869 1835 870
rect 1870 869 1876 870
rect 1742 867 1748 868
rect 1742 863 1743 867
rect 1747 863 1748 867
rect 1742 862 1748 863
rect 1752 859 1754 869
rect 1750 858 1756 859
rect 1750 854 1751 858
rect 1755 854 1756 858
rect 1750 853 1756 854
rect 1832 841 1834 869
rect 1870 865 1871 869
rect 1875 865 1876 869
rect 1918 868 1919 872
rect 1923 868 1924 872
rect 1918 867 1924 868
rect 2094 872 2100 873
rect 2094 868 2095 872
rect 2099 868 2100 872
rect 2094 867 2100 868
rect 2270 872 2276 873
rect 2270 868 2271 872
rect 2275 868 2276 872
rect 2270 867 2276 868
rect 1870 864 1876 865
rect 1986 863 1992 864
rect 1986 859 1987 863
rect 1991 859 1992 863
rect 1986 858 1992 859
rect 1870 852 1876 853
rect 1870 848 1871 852
rect 1875 848 1876 852
rect 1870 847 1876 848
rect 1830 840 1836 841
rect 1830 836 1831 840
rect 1835 836 1836 840
rect 1830 835 1836 836
rect 1562 831 1568 832
rect 1562 827 1563 831
rect 1567 827 1568 831
rect 1562 826 1568 827
rect 1646 831 1652 832
rect 1646 827 1647 831
rect 1651 827 1652 831
rect 1646 826 1652 827
rect 1830 823 1836 824
rect 1630 820 1636 821
rect 1630 816 1631 820
rect 1635 816 1636 820
rect 1630 815 1636 816
rect 1742 820 1748 821
rect 1742 816 1743 820
rect 1747 816 1748 820
rect 1830 819 1831 823
rect 1835 819 1836 823
rect 1872 819 1874 847
rect 1926 834 1932 835
rect 1926 830 1927 834
rect 1931 830 1932 834
rect 1926 829 1932 830
rect 1928 819 1930 829
rect 1988 824 1990 858
rect 2102 834 2108 835
rect 2102 830 2103 834
rect 2107 830 2108 834
rect 2102 829 2108 830
rect 2278 834 2284 835
rect 2278 830 2279 834
rect 2283 830 2284 834
rect 2278 829 2284 830
rect 1986 823 1992 824
rect 1986 819 1987 823
rect 1991 819 1992 823
rect 2104 819 2106 829
rect 2280 819 2282 829
rect 2312 824 2314 906
rect 2328 895 2330 923
rect 2472 895 2474 923
rect 2624 895 2626 923
rect 2784 895 2786 923
rect 2878 911 2884 912
rect 2878 907 2879 911
rect 2883 907 2884 911
rect 2878 906 2884 907
rect 2327 894 2331 895
rect 2327 889 2331 890
rect 2455 894 2459 895
rect 2455 889 2459 890
rect 2471 894 2475 895
rect 2471 889 2475 890
rect 2623 894 2627 895
rect 2623 889 2627 890
rect 2655 894 2659 895
rect 2655 889 2659 890
rect 2783 894 2787 895
rect 2783 889 2787 890
rect 2863 894 2867 895
rect 2863 889 2867 890
rect 2456 873 2458 889
rect 2656 873 2658 889
rect 2864 873 2866 889
rect 2454 872 2460 873
rect 2454 868 2455 872
rect 2459 868 2460 872
rect 2454 867 2460 868
rect 2654 872 2660 873
rect 2654 868 2655 872
rect 2659 868 2660 872
rect 2654 867 2660 868
rect 2862 872 2868 873
rect 2862 868 2863 872
rect 2867 868 2868 872
rect 2862 867 2868 868
rect 2722 863 2728 864
rect 2722 859 2723 863
rect 2727 859 2728 863
rect 2722 858 2728 859
rect 2462 834 2468 835
rect 2462 830 2463 834
rect 2467 830 2468 834
rect 2462 829 2468 830
rect 2662 834 2668 835
rect 2662 830 2663 834
rect 2667 830 2668 834
rect 2662 829 2668 830
rect 2310 823 2316 824
rect 2310 819 2311 823
rect 2315 819 2316 823
rect 2464 819 2466 829
rect 2664 819 2666 829
rect 2724 824 2726 858
rect 2870 834 2876 835
rect 2870 830 2871 834
rect 2875 830 2876 834
rect 2870 829 2876 830
rect 2722 823 2728 824
rect 2722 819 2723 823
rect 2727 819 2728 823
rect 2872 819 2874 829
rect 2880 824 2882 906
rect 2960 895 2962 923
rect 3144 895 3146 923
rect 2959 894 2963 895
rect 2959 889 2963 890
rect 3079 894 3083 895
rect 3079 889 3083 890
rect 3143 894 3147 895
rect 3143 889 3147 890
rect 3080 873 3082 889
rect 3078 872 3084 873
rect 3078 868 3079 872
rect 3083 868 3084 872
rect 3078 867 3084 868
rect 2930 863 2936 864
rect 2930 859 2931 863
rect 2935 859 2936 863
rect 2930 858 2936 859
rect 3194 863 3200 864
rect 3194 859 3195 863
rect 3199 859 3200 863
rect 3194 858 3200 859
rect 2878 823 2884 824
rect 2878 819 2879 823
rect 2883 819 2884 823
rect 1830 818 1836 819
rect 1871 818 1875 819
rect 1742 815 1748 816
rect 1632 787 1634 815
rect 1744 787 1746 815
rect 1832 787 1834 818
rect 1871 813 1875 814
rect 1903 818 1907 819
rect 1903 813 1907 814
rect 1927 818 1931 819
rect 1986 818 1992 819
rect 2015 818 2019 819
rect 1927 813 1931 814
rect 2015 813 2019 814
rect 2103 818 2107 819
rect 2103 813 2107 814
rect 2167 818 2171 819
rect 2167 813 2171 814
rect 2279 818 2283 819
rect 2310 818 2316 819
rect 2327 818 2331 819
rect 2279 813 2283 814
rect 2327 813 2331 814
rect 2463 818 2467 819
rect 2463 813 2467 814
rect 2487 818 2491 819
rect 2487 813 2491 814
rect 2647 818 2651 819
rect 2647 813 2651 814
rect 2663 818 2667 819
rect 2722 818 2728 819
rect 2807 818 2811 819
rect 2663 813 2667 814
rect 2807 813 2811 814
rect 2871 818 2875 819
rect 2878 818 2884 819
rect 2871 813 2875 814
rect 1607 786 1611 787
rect 1607 781 1611 782
rect 1631 786 1635 787
rect 1631 781 1635 782
rect 1743 786 1747 787
rect 1743 781 1747 782
rect 1831 786 1835 787
rect 1872 785 1874 813
rect 1904 803 1906 813
rect 1954 811 1960 812
rect 1954 807 1955 811
rect 1959 807 1960 811
rect 1954 806 1960 807
rect 1902 802 1908 803
rect 1902 798 1903 802
rect 1907 798 1908 802
rect 1902 797 1908 798
rect 1831 781 1835 782
rect 1870 784 1876 785
rect 1608 765 1610 781
rect 1606 764 1612 765
rect 1606 760 1607 764
rect 1611 760 1612 764
rect 1832 762 1834 781
rect 1870 780 1871 784
rect 1875 780 1876 784
rect 1870 779 1876 780
rect 1956 776 1958 806
rect 2016 803 2018 813
rect 2066 811 2072 812
rect 2066 807 2067 811
rect 2071 807 2072 811
rect 2066 806 2072 807
rect 2014 802 2020 803
rect 2014 798 2015 802
rect 2019 798 2020 802
rect 2014 797 2020 798
rect 2068 776 2070 806
rect 2168 803 2170 813
rect 2218 811 2224 812
rect 2218 807 2219 811
rect 2223 807 2224 811
rect 2218 806 2224 807
rect 2166 802 2172 803
rect 2166 798 2167 802
rect 2171 798 2172 802
rect 2166 797 2172 798
rect 2220 776 2222 806
rect 2328 803 2330 813
rect 2378 811 2384 812
rect 2378 807 2379 811
rect 2383 807 2384 811
rect 2378 806 2384 807
rect 2326 802 2332 803
rect 2326 798 2327 802
rect 2331 798 2332 802
rect 2326 797 2332 798
rect 2380 776 2382 806
rect 2488 803 2490 813
rect 2648 803 2650 813
rect 2808 803 2810 813
rect 2932 812 2934 858
rect 3086 834 3092 835
rect 3086 830 3087 834
rect 3091 830 3092 834
rect 3086 829 3092 830
rect 3088 819 3090 829
rect 3196 824 3198 858
rect 3204 824 3206 934
rect 3590 931 3596 932
rect 3334 928 3340 929
rect 3334 924 3335 928
rect 3339 924 3340 928
rect 3334 923 3340 924
rect 3502 928 3508 929
rect 3502 924 3503 928
rect 3507 924 3508 928
rect 3590 927 3591 931
rect 3595 927 3596 931
rect 3590 926 3596 927
rect 3502 923 3508 924
rect 3336 895 3338 923
rect 3504 895 3506 923
rect 3592 895 3594 926
rect 3303 894 3307 895
rect 3303 889 3307 890
rect 3335 894 3339 895
rect 3335 889 3339 890
rect 3503 894 3507 895
rect 3503 889 3507 890
rect 3591 894 3595 895
rect 3591 889 3595 890
rect 3304 873 3306 889
rect 3504 873 3506 889
rect 3302 872 3308 873
rect 3302 868 3303 872
rect 3307 868 3308 872
rect 3302 867 3308 868
rect 3502 872 3508 873
rect 3502 868 3503 872
rect 3507 868 3508 872
rect 3592 870 3594 889
rect 3502 867 3508 868
rect 3590 869 3596 870
rect 3590 865 3591 869
rect 3595 865 3596 869
rect 3590 864 3596 865
rect 3590 852 3596 853
rect 3590 848 3591 852
rect 3595 848 3596 852
rect 3590 847 3596 848
rect 3310 834 3316 835
rect 3310 830 3311 834
rect 3315 830 3316 834
rect 3310 829 3316 830
rect 3510 834 3516 835
rect 3510 830 3511 834
rect 3515 830 3516 834
rect 3510 829 3516 830
rect 3194 823 3200 824
rect 3194 819 3195 823
rect 3199 819 3200 823
rect 2959 818 2963 819
rect 2959 813 2963 814
rect 3087 818 3091 819
rect 3087 813 3091 814
rect 3103 818 3107 819
rect 3194 818 3200 819
rect 3202 823 3208 824
rect 3202 819 3203 823
rect 3207 819 3208 823
rect 3312 819 3314 829
rect 3512 819 3514 829
rect 3518 823 3524 824
rect 3518 819 3519 823
rect 3523 819 3524 823
rect 3592 819 3594 847
rect 3202 818 3208 819
rect 3247 818 3251 819
rect 3103 813 3107 814
rect 3247 813 3251 814
rect 3311 818 3315 819
rect 3311 813 3315 814
rect 3391 818 3395 819
rect 3391 813 3395 814
rect 3511 818 3515 819
rect 3518 818 3524 819
rect 3591 818 3595 819
rect 3511 813 3515 814
rect 2930 811 2936 812
rect 2930 807 2931 811
rect 2935 807 2936 811
rect 2930 806 2936 807
rect 2960 803 2962 813
rect 2978 811 2984 812
rect 2978 807 2979 811
rect 2983 807 2984 811
rect 2978 806 2984 807
rect 3010 811 3016 812
rect 3010 807 3011 811
rect 3015 807 3016 811
rect 3010 806 3016 807
rect 2486 802 2492 803
rect 2486 798 2487 802
rect 2491 798 2492 802
rect 2486 797 2492 798
rect 2646 802 2652 803
rect 2646 798 2647 802
rect 2651 798 2652 802
rect 2646 797 2652 798
rect 2806 802 2812 803
rect 2806 798 2807 802
rect 2811 798 2812 802
rect 2806 797 2812 798
rect 2958 802 2964 803
rect 2958 798 2959 802
rect 2963 798 2964 802
rect 2958 797 2964 798
rect 1954 775 1960 776
rect 1954 771 1955 775
rect 1959 771 1960 775
rect 1954 770 1960 771
rect 2066 775 2072 776
rect 2066 771 2067 775
rect 2071 771 2072 775
rect 2066 770 2072 771
rect 2218 775 2224 776
rect 2218 771 2219 775
rect 2223 771 2224 775
rect 2218 770 2224 771
rect 2378 775 2384 776
rect 2378 771 2379 775
rect 2383 771 2384 775
rect 2378 770 2384 771
rect 2698 775 2704 776
rect 2698 771 2699 775
rect 2703 771 2704 775
rect 2698 770 2704 771
rect 2870 775 2876 776
rect 2870 771 2871 775
rect 2875 771 2876 775
rect 2870 770 2876 771
rect 1870 767 1876 768
rect 1870 763 1871 767
rect 1875 763 1876 767
rect 1870 762 1876 763
rect 1894 764 1900 765
rect 1606 759 1612 760
rect 1830 761 1836 762
rect 1830 757 1831 761
rect 1835 757 1836 761
rect 1830 756 1836 757
rect 1378 755 1384 756
rect 1378 751 1379 755
rect 1383 751 1384 755
rect 1378 750 1384 751
rect 1518 755 1524 756
rect 1518 751 1519 755
rect 1523 751 1524 755
rect 1518 750 1524 751
rect 1530 755 1536 756
rect 1530 751 1531 755
rect 1535 751 1536 755
rect 1530 750 1536 751
rect 1302 726 1308 727
rect 1302 722 1303 726
rect 1307 722 1308 726
rect 1302 721 1308 722
rect 1311 724 1315 725
rect 1158 715 1164 716
rect 1158 711 1159 715
rect 1163 711 1164 715
rect 1158 710 1164 711
rect 1304 703 1306 721
rect 1311 719 1315 720
rect 1312 716 1314 719
rect 1380 716 1382 750
rect 1454 726 1460 727
rect 1454 722 1455 726
rect 1459 722 1460 726
rect 1532 725 1534 750
rect 1830 744 1836 745
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1872 743 1874 762
rect 1894 760 1895 764
rect 1899 760 1900 764
rect 1894 759 1900 760
rect 2006 764 2012 765
rect 2006 760 2007 764
rect 2011 760 2012 764
rect 2006 759 2012 760
rect 2158 764 2164 765
rect 2158 760 2159 764
rect 2163 760 2164 764
rect 2158 759 2164 760
rect 2318 764 2324 765
rect 2318 760 2319 764
rect 2323 760 2324 764
rect 2318 759 2324 760
rect 2478 764 2484 765
rect 2478 760 2479 764
rect 2483 760 2484 764
rect 2478 759 2484 760
rect 2638 764 2644 765
rect 2638 760 2639 764
rect 2643 760 2644 764
rect 2638 759 2644 760
rect 1896 743 1898 759
rect 2008 743 2010 759
rect 2160 743 2162 759
rect 2320 743 2322 759
rect 2418 747 2424 748
rect 2418 743 2419 747
rect 2423 743 2424 747
rect 2480 743 2482 759
rect 2640 743 2642 759
rect 1830 739 1836 740
rect 1871 742 1875 743
rect 1614 726 1620 727
rect 1454 721 1460 722
rect 1531 724 1535 725
rect 1310 715 1316 716
rect 1310 711 1311 715
rect 1315 711 1316 715
rect 1310 710 1316 711
rect 1378 715 1384 716
rect 1378 711 1379 715
rect 1383 711 1384 715
rect 1378 710 1384 711
rect 1456 703 1458 721
rect 1614 722 1615 726
rect 1619 722 1620 726
rect 1614 721 1620 722
rect 1531 719 1535 720
rect 1606 715 1612 716
rect 1606 711 1607 715
rect 1611 711 1612 715
rect 1606 710 1612 711
rect 951 702 955 703
rect 951 697 955 698
rect 999 702 1003 703
rect 999 697 1003 698
rect 1087 702 1091 703
rect 1087 697 1091 698
rect 1151 702 1155 703
rect 1151 697 1155 698
rect 1215 702 1219 703
rect 1215 697 1219 698
rect 1303 702 1307 703
rect 1303 697 1307 698
rect 1335 702 1339 703
rect 1335 697 1339 698
rect 1455 702 1459 703
rect 1455 697 1459 698
rect 1583 702 1587 703
rect 1583 697 1587 698
rect 854 695 860 696
rect 854 691 855 695
rect 859 691 860 695
rect 854 690 860 691
rect 906 695 912 696
rect 906 691 907 695
rect 911 691 912 695
rect 906 690 912 691
rect 814 686 820 687
rect 814 682 815 686
rect 819 682 820 686
rect 814 681 820 682
rect 282 659 288 660
rect 282 655 283 659
rect 287 655 288 659
rect 282 654 288 655
rect 370 659 376 660
rect 370 655 371 659
rect 375 655 376 659
rect 370 654 376 655
rect 430 659 436 660
rect 430 655 431 659
rect 435 655 436 659
rect 430 654 436 655
rect 550 659 556 660
rect 550 655 551 659
rect 555 655 556 659
rect 550 654 556 655
rect 602 659 608 660
rect 602 655 603 659
rect 607 655 608 659
rect 602 654 608 655
rect 738 659 744 660
rect 738 655 739 659
rect 743 655 744 659
rect 738 654 744 655
rect 110 651 116 652
rect 110 647 111 651
rect 115 647 116 651
rect 110 646 116 647
rect 222 648 228 649
rect 112 619 114 646
rect 222 644 223 648
rect 227 644 228 648
rect 222 643 228 644
rect 310 648 316 649
rect 310 644 311 648
rect 315 644 316 648
rect 310 643 316 644
rect 414 648 420 649
rect 414 644 415 648
rect 419 644 420 648
rect 414 643 420 644
rect 534 648 540 649
rect 534 644 535 648
rect 539 644 540 648
rect 534 643 540 644
rect 670 648 676 649
rect 670 644 671 648
rect 675 644 676 648
rect 670 643 676 644
rect 806 648 812 649
rect 806 644 807 648
rect 811 644 812 648
rect 806 643 812 644
rect 224 619 226 643
rect 312 619 314 643
rect 416 619 418 643
rect 536 619 538 643
rect 672 619 674 643
rect 808 619 810 643
rect 111 618 115 619
rect 111 613 115 614
rect 223 618 227 619
rect 223 613 227 614
rect 311 618 315 619
rect 311 613 315 614
rect 415 618 419 619
rect 415 613 419 614
rect 447 618 451 619
rect 447 613 451 614
rect 527 618 531 619
rect 527 613 531 614
rect 535 618 539 619
rect 535 613 539 614
rect 607 618 611 619
rect 607 613 611 614
rect 671 618 675 619
rect 671 613 675 614
rect 687 618 691 619
rect 687 613 691 614
rect 775 618 779 619
rect 775 613 779 614
rect 807 618 811 619
rect 807 613 811 614
rect 112 594 114 613
rect 448 597 450 613
rect 528 597 530 613
rect 608 597 610 613
rect 688 597 690 613
rect 776 597 778 613
rect 446 596 452 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 446 592 447 596
rect 451 592 452 596
rect 446 591 452 592
rect 526 596 532 597
rect 526 592 527 596
rect 531 592 532 596
rect 526 591 532 592
rect 606 596 612 597
rect 606 592 607 596
rect 611 592 612 596
rect 606 591 612 592
rect 686 596 692 597
rect 686 592 687 596
rect 691 592 692 596
rect 686 591 692 592
rect 774 596 780 597
rect 774 592 775 596
rect 779 592 780 596
rect 774 591 780 592
rect 110 588 116 589
rect 856 588 858 690
rect 952 687 954 697
rect 1088 687 1090 697
rect 1094 695 1100 696
rect 1094 691 1095 695
rect 1099 691 1100 695
rect 1094 690 1100 691
rect 1138 695 1144 696
rect 1138 691 1139 695
rect 1143 691 1144 695
rect 1138 690 1144 691
rect 950 686 956 687
rect 950 682 951 686
rect 955 682 956 686
rect 950 681 956 682
rect 1086 686 1092 687
rect 1086 682 1087 686
rect 1091 682 1092 686
rect 1086 681 1092 682
rect 942 648 948 649
rect 942 644 943 648
rect 947 644 948 648
rect 942 643 948 644
rect 1078 648 1084 649
rect 1078 644 1079 648
rect 1083 644 1084 648
rect 1078 643 1084 644
rect 944 619 946 643
rect 1080 619 1082 643
rect 1096 629 1098 690
rect 1140 660 1142 690
rect 1216 687 1218 697
rect 1266 695 1272 696
rect 1266 691 1267 695
rect 1271 691 1272 695
rect 1266 690 1272 691
rect 1214 686 1220 687
rect 1214 682 1215 686
rect 1219 682 1220 686
rect 1214 681 1220 682
rect 1268 660 1270 690
rect 1336 687 1338 697
rect 1386 695 1392 696
rect 1386 691 1387 695
rect 1391 691 1392 695
rect 1386 690 1392 691
rect 1334 686 1340 687
rect 1334 682 1335 686
rect 1339 682 1340 686
rect 1334 681 1340 682
rect 1388 660 1390 690
rect 1456 687 1458 697
rect 1506 695 1512 696
rect 1506 691 1507 695
rect 1511 691 1512 695
rect 1506 690 1512 691
rect 1454 686 1460 687
rect 1454 682 1455 686
rect 1459 682 1460 686
rect 1454 681 1460 682
rect 1508 660 1510 690
rect 1584 687 1586 697
rect 1582 686 1588 687
rect 1582 682 1583 686
rect 1587 682 1588 686
rect 1582 681 1588 682
rect 1608 660 1610 710
rect 1616 703 1618 721
rect 1832 703 1834 739
rect 1871 737 1875 738
rect 1895 742 1899 743
rect 1895 737 1899 738
rect 1967 742 1971 743
rect 1967 737 1971 738
rect 2007 742 2011 743
rect 2007 737 2011 738
rect 2063 742 2067 743
rect 2063 737 2067 738
rect 2159 742 2163 743
rect 2159 737 2163 738
rect 2175 742 2179 743
rect 2175 737 2179 738
rect 2303 742 2307 743
rect 2303 737 2307 738
rect 2319 742 2323 743
rect 2418 742 2424 743
rect 2447 742 2451 743
rect 2319 737 2323 738
rect 1872 718 1874 737
rect 1968 721 1970 737
rect 2064 721 2066 737
rect 2176 721 2178 737
rect 2304 721 2306 737
rect 1966 720 1972 721
rect 1870 717 1876 718
rect 1870 713 1871 717
rect 1875 713 1876 717
rect 1966 716 1967 720
rect 1971 716 1972 720
rect 1966 715 1972 716
rect 2062 720 2068 721
rect 2062 716 2063 720
rect 2067 716 2068 720
rect 2062 715 2068 716
rect 2174 720 2180 721
rect 2174 716 2175 720
rect 2179 716 2180 720
rect 2302 720 2308 721
rect 2174 715 2180 716
rect 2191 716 2195 717
rect 1870 712 1876 713
rect 2302 716 2303 720
rect 2307 716 2308 720
rect 2302 715 2308 716
rect 2034 711 2040 712
rect 2034 707 2035 711
rect 2039 707 2040 711
rect 2034 706 2040 707
rect 2130 711 2136 712
rect 2191 711 2195 712
rect 2246 711 2252 712
rect 2130 707 2131 711
rect 2135 707 2136 711
rect 2130 706 2136 707
rect 1615 702 1619 703
rect 1615 697 1619 698
rect 1831 702 1835 703
rect 1831 697 1835 698
rect 1870 700 1876 701
rect 1832 669 1834 697
rect 1870 696 1871 700
rect 1875 696 1876 700
rect 1870 695 1876 696
rect 1830 668 1836 669
rect 1830 664 1831 668
rect 1835 664 1836 668
rect 1872 667 1874 695
rect 1974 682 1980 683
rect 1974 678 1975 682
rect 1979 678 1980 682
rect 1974 677 1980 678
rect 1976 667 1978 677
rect 1983 676 1987 677
rect 2036 672 2038 706
rect 2070 682 2076 683
rect 2070 678 2071 682
rect 2075 678 2076 682
rect 2070 677 2076 678
rect 1982 671 1988 672
rect 1982 667 1983 671
rect 1987 667 1988 671
rect 1830 663 1836 664
rect 1871 666 1875 667
rect 1871 661 1875 662
rect 1975 666 1979 667
rect 1982 666 1988 667
rect 2034 671 2040 672
rect 2034 667 2035 671
rect 2039 667 2040 671
rect 2072 667 2074 677
rect 2132 672 2134 706
rect 2182 682 2188 683
rect 2182 678 2183 682
rect 2187 678 2188 682
rect 2182 677 2188 678
rect 2130 671 2136 672
rect 2130 667 2131 671
rect 2135 667 2136 671
rect 2184 667 2186 677
rect 2034 666 2040 667
rect 2071 666 2075 667
rect 2130 666 2136 667
rect 2175 666 2179 667
rect 1975 661 1979 662
rect 2071 661 2075 662
rect 2175 661 2179 662
rect 2183 666 2187 667
rect 2183 661 2187 662
rect 1138 659 1144 660
rect 1138 655 1139 659
rect 1143 655 1144 659
rect 1138 654 1144 655
rect 1266 659 1272 660
rect 1266 655 1267 659
rect 1271 655 1272 659
rect 1266 654 1272 655
rect 1386 659 1392 660
rect 1386 655 1387 659
rect 1391 655 1392 659
rect 1386 654 1392 655
rect 1506 659 1512 660
rect 1506 655 1507 659
rect 1511 655 1512 659
rect 1506 654 1512 655
rect 1606 659 1612 660
rect 1606 655 1607 659
rect 1611 655 1612 659
rect 1606 654 1612 655
rect 1830 651 1836 652
rect 1206 648 1212 649
rect 1206 644 1207 648
rect 1211 644 1212 648
rect 1206 643 1212 644
rect 1326 648 1332 649
rect 1326 644 1327 648
rect 1331 644 1332 648
rect 1326 643 1332 644
rect 1446 648 1452 649
rect 1446 644 1447 648
rect 1451 644 1452 648
rect 1446 643 1452 644
rect 1574 648 1580 649
rect 1574 644 1575 648
rect 1579 644 1580 648
rect 1830 647 1831 651
rect 1835 647 1836 651
rect 1830 646 1836 647
rect 1574 643 1580 644
rect 1095 628 1099 629
rect 1095 623 1099 624
rect 1208 619 1210 643
rect 1328 619 1330 643
rect 1411 628 1415 629
rect 1411 623 1415 624
rect 871 618 875 619
rect 871 613 875 614
rect 943 618 947 619
rect 943 613 947 614
rect 959 618 963 619
rect 959 613 963 614
rect 1047 618 1051 619
rect 1047 613 1051 614
rect 1079 618 1083 619
rect 1079 613 1083 614
rect 1143 618 1147 619
rect 1143 613 1147 614
rect 1207 618 1211 619
rect 1207 613 1211 614
rect 1239 618 1243 619
rect 1239 613 1243 614
rect 1327 618 1331 619
rect 1327 613 1331 614
rect 1335 618 1339 619
rect 1335 613 1339 614
rect 872 597 874 613
rect 960 597 962 613
rect 1048 597 1050 613
rect 1144 597 1146 613
rect 1240 597 1242 613
rect 1336 597 1338 613
rect 870 596 876 597
rect 870 592 871 596
rect 875 592 876 596
rect 870 591 876 592
rect 958 596 964 597
rect 958 592 959 596
rect 963 592 964 596
rect 958 591 964 592
rect 1046 596 1052 597
rect 1046 592 1047 596
rect 1051 592 1052 596
rect 1046 591 1052 592
rect 1142 596 1148 597
rect 1142 592 1143 596
rect 1147 592 1148 596
rect 1142 591 1148 592
rect 1238 596 1244 597
rect 1238 592 1239 596
rect 1243 592 1244 596
rect 1238 591 1244 592
rect 1334 596 1340 597
rect 1334 592 1335 596
rect 1339 592 1340 596
rect 1334 591 1340 592
rect 1412 588 1414 623
rect 1448 619 1450 643
rect 1576 619 1578 643
rect 1832 619 1834 646
rect 1872 633 1874 661
rect 2176 651 2178 661
rect 2192 660 2194 711
rect 2246 707 2247 711
rect 2251 707 2252 711
rect 2246 706 2252 707
rect 2382 711 2388 712
rect 2382 707 2383 711
rect 2387 707 2388 711
rect 2382 706 2388 707
rect 2248 672 2250 706
rect 2310 682 2316 683
rect 2310 678 2311 682
rect 2315 678 2316 682
rect 2310 677 2316 678
rect 2246 671 2252 672
rect 2246 667 2247 671
rect 2251 667 2252 671
rect 2312 667 2314 677
rect 2384 672 2386 706
rect 2420 677 2422 742
rect 2447 737 2451 738
rect 2479 742 2483 743
rect 2479 737 2483 738
rect 2599 742 2603 743
rect 2599 737 2603 738
rect 2639 742 2643 743
rect 2639 737 2643 738
rect 2448 721 2450 737
rect 2600 721 2602 737
rect 2446 720 2452 721
rect 2446 716 2447 720
rect 2451 716 2452 720
rect 2446 715 2452 716
rect 2598 720 2604 721
rect 2598 716 2599 720
rect 2603 716 2604 720
rect 2598 715 2604 716
rect 2607 716 2611 717
rect 2607 711 2611 712
rect 2608 708 2610 711
rect 2606 707 2612 708
rect 2606 703 2607 707
rect 2611 703 2612 707
rect 2606 702 2612 703
rect 2454 682 2460 683
rect 2454 678 2455 682
rect 2459 678 2460 682
rect 2454 677 2460 678
rect 2606 682 2612 683
rect 2606 678 2607 682
rect 2611 678 2612 682
rect 2606 677 2612 678
rect 2419 676 2423 677
rect 2382 671 2388 672
rect 2419 671 2423 672
rect 2382 667 2383 671
rect 2387 667 2388 671
rect 2456 667 2458 677
rect 2608 667 2610 677
rect 2700 672 2702 770
rect 2798 764 2804 765
rect 2798 760 2799 764
rect 2803 760 2804 764
rect 2798 759 2804 760
rect 2800 743 2802 759
rect 2751 742 2755 743
rect 2751 737 2755 738
rect 2799 742 2803 743
rect 2799 737 2803 738
rect 2752 721 2754 737
rect 2750 720 2756 721
rect 2750 716 2751 720
rect 2755 716 2756 720
rect 2750 715 2756 716
rect 2818 711 2824 712
rect 2818 707 2819 711
rect 2823 707 2824 711
rect 2818 706 2824 707
rect 2758 682 2764 683
rect 2758 678 2759 682
rect 2763 678 2764 682
rect 2758 677 2764 678
rect 2698 671 2704 672
rect 2698 667 2699 671
rect 2703 667 2704 671
rect 2760 667 2762 677
rect 2246 666 2252 667
rect 2271 666 2275 667
rect 2271 661 2275 662
rect 2311 666 2315 667
rect 2311 661 2315 662
rect 2375 666 2379 667
rect 2382 666 2388 667
rect 2455 666 2459 667
rect 2375 661 2379 662
rect 2455 661 2459 662
rect 2487 666 2491 667
rect 2487 661 2491 662
rect 2607 666 2611 667
rect 2698 666 2704 667
rect 2735 666 2739 667
rect 2607 661 2611 662
rect 2735 661 2739 662
rect 2759 666 2763 667
rect 2759 661 2763 662
rect 2190 659 2196 660
rect 2190 655 2191 659
rect 2195 655 2196 659
rect 2190 654 2196 655
rect 2226 659 2232 660
rect 2226 655 2227 659
rect 2231 655 2232 659
rect 2226 654 2232 655
rect 2174 650 2180 651
rect 2174 646 2175 650
rect 2179 646 2180 650
rect 2174 645 2180 646
rect 1870 632 1876 633
rect 1870 628 1871 632
rect 1875 628 1876 632
rect 1870 627 1876 628
rect 2228 624 2230 654
rect 2272 651 2274 661
rect 2322 659 2328 660
rect 2322 655 2323 659
rect 2327 655 2328 659
rect 2322 654 2328 655
rect 2270 650 2276 651
rect 2270 646 2271 650
rect 2275 646 2276 650
rect 2270 645 2276 646
rect 2324 624 2326 654
rect 2376 651 2378 661
rect 2426 659 2432 660
rect 2426 655 2427 659
rect 2431 655 2432 659
rect 2426 654 2432 655
rect 2374 650 2380 651
rect 2374 646 2375 650
rect 2379 646 2380 650
rect 2374 645 2380 646
rect 2428 624 2430 654
rect 2488 651 2490 661
rect 2538 659 2544 660
rect 2538 655 2539 659
rect 2543 655 2544 659
rect 2538 654 2544 655
rect 2486 650 2492 651
rect 2486 646 2487 650
rect 2491 646 2492 650
rect 2486 645 2492 646
rect 2540 624 2542 654
rect 2608 651 2610 661
rect 2736 651 2738 661
rect 2820 660 2822 706
rect 2872 672 2874 770
rect 2950 764 2956 765
rect 2950 760 2951 764
rect 2955 760 2956 764
rect 2950 759 2956 760
rect 2952 743 2954 759
rect 2903 742 2907 743
rect 2903 737 2907 738
rect 2951 742 2955 743
rect 2951 737 2955 738
rect 2904 721 2906 737
rect 2902 720 2908 721
rect 2902 716 2903 720
rect 2907 716 2908 720
rect 2902 715 2908 716
rect 2980 712 2982 806
rect 3012 776 3014 806
rect 3104 803 3106 813
rect 3154 811 3160 812
rect 3154 807 3155 811
rect 3159 807 3160 811
rect 3154 806 3160 807
rect 3102 802 3108 803
rect 3102 798 3103 802
rect 3107 798 3108 802
rect 3102 797 3108 798
rect 3156 776 3158 806
rect 3248 803 3250 813
rect 3298 811 3304 812
rect 3298 807 3299 811
rect 3303 807 3304 811
rect 3298 806 3304 807
rect 3246 802 3252 803
rect 3246 798 3247 802
rect 3251 798 3252 802
rect 3246 797 3252 798
rect 3300 776 3302 806
rect 3392 803 3394 813
rect 3512 803 3514 813
rect 3390 802 3396 803
rect 3390 798 3391 802
rect 3395 798 3396 802
rect 3390 797 3396 798
rect 3510 802 3516 803
rect 3510 798 3511 802
rect 3515 798 3516 802
rect 3510 797 3516 798
rect 3520 776 3522 818
rect 3591 813 3595 814
rect 3592 785 3594 813
rect 3590 784 3596 785
rect 3590 780 3591 784
rect 3595 780 3596 784
rect 3590 779 3596 780
rect 3010 775 3016 776
rect 3010 771 3011 775
rect 3015 771 3016 775
rect 3010 770 3016 771
rect 3154 775 3160 776
rect 3154 771 3155 775
rect 3159 771 3160 775
rect 3154 770 3160 771
rect 3298 775 3304 776
rect 3298 771 3299 775
rect 3303 771 3304 775
rect 3298 770 3304 771
rect 3518 775 3524 776
rect 3518 771 3519 775
rect 3523 771 3524 775
rect 3518 770 3524 771
rect 3590 767 3596 768
rect 3094 764 3100 765
rect 3094 760 3095 764
rect 3099 760 3100 764
rect 3094 759 3100 760
rect 3238 764 3244 765
rect 3238 760 3239 764
rect 3243 760 3244 764
rect 3238 759 3244 760
rect 3382 764 3388 765
rect 3382 760 3383 764
rect 3387 760 3388 764
rect 3382 759 3388 760
rect 3502 764 3508 765
rect 3502 760 3503 764
rect 3507 760 3508 764
rect 3590 763 3591 767
rect 3595 763 3596 767
rect 3590 762 3596 763
rect 3502 759 3508 760
rect 3096 743 3098 759
rect 3240 743 3242 759
rect 3374 747 3380 748
rect 3374 743 3375 747
rect 3379 743 3380 747
rect 3384 743 3386 759
rect 3504 743 3506 759
rect 3592 743 3594 762
rect 3055 742 3059 743
rect 3055 737 3059 738
rect 3095 742 3099 743
rect 3095 737 3099 738
rect 3207 742 3211 743
rect 3207 737 3211 738
rect 3239 742 3243 743
rect 3239 737 3243 738
rect 3359 742 3363 743
rect 3374 742 3380 743
rect 3383 742 3387 743
rect 3359 737 3363 738
rect 3056 721 3058 737
rect 3208 721 3210 737
rect 3360 721 3362 737
rect 3054 720 3060 721
rect 3054 716 3055 720
rect 3059 716 3060 720
rect 3054 715 3060 716
rect 3206 720 3212 721
rect 3206 716 3207 720
rect 3211 716 3212 720
rect 3206 715 3212 716
rect 3358 720 3364 721
rect 3358 716 3359 720
rect 3363 716 3364 720
rect 3358 715 3364 716
rect 2978 711 2984 712
rect 2978 707 2979 711
rect 2983 707 2984 711
rect 2978 706 2984 707
rect 3274 711 3280 712
rect 3274 707 3275 711
rect 3279 707 3280 711
rect 3274 706 3280 707
rect 3266 703 3272 704
rect 3266 699 3267 703
rect 3271 699 3272 703
rect 3266 698 3272 699
rect 2910 682 2916 683
rect 2910 678 2911 682
rect 2915 678 2916 682
rect 2910 677 2916 678
rect 3062 682 3068 683
rect 3062 678 3063 682
rect 3067 678 3068 682
rect 3062 677 3068 678
rect 3214 682 3220 683
rect 3214 678 3215 682
rect 3219 678 3220 682
rect 3214 677 3220 678
rect 2870 671 2876 672
rect 2870 667 2871 671
rect 2875 667 2876 671
rect 2912 667 2914 677
rect 3064 667 3066 677
rect 3126 671 3132 672
rect 3126 667 3127 671
rect 3131 667 3132 671
rect 3216 667 3218 677
rect 2863 666 2867 667
rect 2870 666 2876 667
rect 2911 666 2915 667
rect 2863 661 2867 662
rect 2911 661 2915 662
rect 2991 666 2995 667
rect 2991 661 2995 662
rect 3063 666 3067 667
rect 3063 661 3067 662
rect 3119 666 3123 667
rect 3126 666 3132 667
rect 3215 666 3219 667
rect 3119 661 3123 662
rect 2818 659 2824 660
rect 2818 655 2819 659
rect 2823 655 2824 659
rect 2818 654 2824 655
rect 2864 651 2866 661
rect 2982 659 2988 660
rect 2982 655 2983 659
rect 2987 655 2988 659
rect 2982 654 2988 655
rect 2606 650 2612 651
rect 2606 646 2607 650
rect 2611 646 2612 650
rect 2606 645 2612 646
rect 2734 650 2740 651
rect 2734 646 2735 650
rect 2739 646 2740 650
rect 2734 645 2740 646
rect 2862 650 2868 651
rect 2862 646 2863 650
rect 2867 646 2868 650
rect 2862 645 2868 646
rect 2984 624 2986 654
rect 2992 651 2994 661
rect 3120 651 3122 661
rect 2990 650 2996 651
rect 2990 646 2991 650
rect 2995 646 2996 650
rect 2990 645 2996 646
rect 3118 650 3124 651
rect 3118 646 3119 650
rect 3123 646 3124 650
rect 3118 645 3124 646
rect 3128 624 3130 666
rect 3215 661 3219 662
rect 3247 666 3251 667
rect 3247 661 3251 662
rect 3248 651 3250 661
rect 3268 660 3270 698
rect 3276 672 3278 706
rect 3366 682 3372 683
rect 3366 678 3367 682
rect 3371 678 3372 682
rect 3366 677 3372 678
rect 3274 671 3280 672
rect 3274 667 3275 671
rect 3279 667 3280 671
rect 3368 667 3370 677
rect 3376 676 3378 742
rect 3383 737 3387 738
rect 3503 742 3507 743
rect 3503 737 3507 738
rect 3591 742 3595 743
rect 3591 737 3595 738
rect 3504 721 3506 737
rect 3502 720 3508 721
rect 3502 716 3503 720
rect 3507 716 3508 720
rect 3592 718 3594 737
rect 3502 715 3508 716
rect 3590 717 3596 718
rect 3590 713 3591 717
rect 3595 713 3596 717
rect 3590 712 3596 713
rect 3590 700 3596 701
rect 3590 696 3591 700
rect 3595 696 3596 700
rect 3590 695 3596 696
rect 3510 682 3516 683
rect 3510 678 3511 682
rect 3515 678 3516 682
rect 3510 677 3516 678
rect 3374 675 3380 676
rect 3374 671 3375 675
rect 3379 671 3380 675
rect 3374 670 3380 671
rect 3512 667 3514 677
rect 3518 671 3524 672
rect 3518 667 3519 671
rect 3523 667 3524 671
rect 3592 667 3594 695
rect 3274 666 3280 667
rect 3367 666 3371 667
rect 3367 661 3371 662
rect 3375 666 3379 667
rect 3375 661 3379 662
rect 3511 666 3515 667
rect 3518 666 3524 667
rect 3591 666 3595 667
rect 3511 661 3515 662
rect 3266 659 3272 660
rect 3266 655 3267 659
rect 3271 655 3272 659
rect 3266 654 3272 655
rect 3298 659 3304 660
rect 3298 655 3299 659
rect 3303 655 3304 659
rect 3298 654 3304 655
rect 3246 650 3252 651
rect 3246 646 3247 650
rect 3251 646 3252 650
rect 3246 645 3252 646
rect 3300 624 3302 654
rect 3376 651 3378 661
rect 3512 651 3514 661
rect 3374 650 3380 651
rect 3374 646 3375 650
rect 3379 646 3380 650
rect 3374 645 3380 646
rect 3510 650 3516 651
rect 3510 646 3511 650
rect 3515 646 3516 650
rect 3510 645 3516 646
rect 3520 624 3522 666
rect 3591 661 3595 662
rect 3526 659 3532 660
rect 3526 655 3527 659
rect 3531 655 3532 659
rect 3526 654 3532 655
rect 2226 623 2232 624
rect 2226 619 2227 623
rect 2231 619 2232 623
rect 1431 618 1435 619
rect 1431 613 1435 614
rect 1447 618 1451 619
rect 1447 613 1451 614
rect 1575 618 1579 619
rect 1575 613 1579 614
rect 1831 618 1835 619
rect 2226 618 2232 619
rect 2322 623 2328 624
rect 2322 619 2323 623
rect 2327 619 2328 623
rect 2322 618 2328 619
rect 2426 623 2432 624
rect 2426 619 2427 623
rect 2431 619 2432 623
rect 2426 618 2432 619
rect 2538 623 2544 624
rect 2538 619 2539 623
rect 2543 619 2544 623
rect 2538 618 2544 619
rect 2786 623 2792 624
rect 2786 619 2787 623
rect 2791 619 2792 623
rect 2786 618 2792 619
rect 2982 623 2988 624
rect 2982 619 2983 623
rect 2987 619 2988 623
rect 2982 618 2988 619
rect 3042 623 3048 624
rect 3042 619 3043 623
rect 3047 619 3048 623
rect 3042 618 3048 619
rect 3126 623 3132 624
rect 3126 619 3127 623
rect 3131 619 3132 623
rect 3126 618 3132 619
rect 3298 623 3304 624
rect 3298 619 3299 623
rect 3303 619 3304 623
rect 3298 618 3304 619
rect 3426 623 3432 624
rect 3426 619 3427 623
rect 3431 619 3432 623
rect 3426 618 3432 619
rect 3518 623 3524 624
rect 3518 619 3519 623
rect 3523 619 3524 623
rect 3518 618 3524 619
rect 1831 613 1835 614
rect 1870 615 1876 616
rect 1432 597 1434 613
rect 1430 596 1436 597
rect 1430 592 1431 596
rect 1435 592 1436 596
rect 1832 594 1834 613
rect 1870 611 1871 615
rect 1875 611 1876 615
rect 1870 610 1876 611
rect 2166 612 2172 613
rect 1430 591 1436 592
rect 1830 593 1836 594
rect 1830 589 1831 593
rect 1835 589 1836 593
rect 1872 591 1874 610
rect 2166 608 2167 612
rect 2171 608 2172 612
rect 2166 607 2172 608
rect 2262 612 2268 613
rect 2262 608 2263 612
rect 2267 608 2268 612
rect 2262 607 2268 608
rect 2366 612 2372 613
rect 2366 608 2367 612
rect 2371 608 2372 612
rect 2366 607 2372 608
rect 2478 612 2484 613
rect 2478 608 2479 612
rect 2483 608 2484 612
rect 2478 607 2484 608
rect 2598 612 2604 613
rect 2598 608 2599 612
rect 2603 608 2604 612
rect 2598 607 2604 608
rect 2726 612 2732 613
rect 2726 608 2727 612
rect 2731 608 2732 612
rect 2726 607 2732 608
rect 2168 591 2170 607
rect 2264 591 2266 607
rect 2368 591 2370 607
rect 2480 591 2482 607
rect 2538 595 2544 596
rect 2538 591 2539 595
rect 2543 591 2544 595
rect 2600 591 2602 607
rect 2728 591 2730 607
rect 1830 588 1836 589
rect 1871 590 1875 591
rect 514 587 520 588
rect 514 583 515 587
rect 519 583 520 587
rect 514 582 520 583
rect 594 587 600 588
rect 594 583 595 587
rect 599 583 600 587
rect 594 582 600 583
rect 674 587 680 588
rect 674 583 675 587
rect 679 583 680 587
rect 674 582 680 583
rect 754 587 760 588
rect 754 583 755 587
rect 759 583 760 587
rect 754 582 760 583
rect 854 587 860 588
rect 854 583 855 587
rect 859 583 860 587
rect 854 582 860 583
rect 862 587 868 588
rect 862 583 863 587
rect 867 583 868 587
rect 862 582 868 583
rect 938 587 944 588
rect 938 583 939 587
rect 943 583 944 587
rect 938 582 944 583
rect 1114 587 1120 588
rect 1114 583 1115 587
rect 1119 583 1120 587
rect 1114 582 1120 583
rect 1210 587 1216 588
rect 1210 583 1211 587
rect 1215 583 1216 587
rect 1210 582 1216 583
rect 1306 587 1312 588
rect 1306 583 1307 587
rect 1311 583 1312 587
rect 1306 582 1312 583
rect 1402 587 1408 588
rect 1402 583 1403 587
rect 1407 583 1408 587
rect 1402 582 1408 583
rect 1410 587 1416 588
rect 1410 583 1411 587
rect 1415 583 1416 587
rect 1871 585 1875 586
rect 2167 590 2171 591
rect 2167 585 2171 586
rect 2263 590 2267 591
rect 2263 585 2267 586
rect 2343 590 2347 591
rect 2343 585 2347 586
rect 2367 590 2371 591
rect 2367 585 2371 586
rect 2423 590 2427 591
rect 2423 585 2427 586
rect 2479 590 2483 591
rect 2479 585 2483 586
rect 2503 590 2507 591
rect 2538 590 2544 591
rect 2591 590 2595 591
rect 2503 585 2507 586
rect 1410 582 1416 583
rect 110 576 116 577
rect 110 572 111 576
rect 115 572 116 576
rect 110 571 116 572
rect 112 531 114 571
rect 454 558 460 559
rect 454 554 455 558
rect 459 554 460 558
rect 454 553 460 554
rect 456 531 458 553
rect 516 548 518 582
rect 534 558 540 559
rect 534 554 535 558
rect 539 554 540 558
rect 534 553 540 554
rect 514 547 520 548
rect 514 543 515 547
rect 519 543 520 547
rect 514 542 520 543
rect 536 531 538 553
rect 596 548 598 582
rect 614 558 620 559
rect 614 554 615 558
rect 619 554 620 558
rect 614 553 620 554
rect 594 547 600 548
rect 594 543 595 547
rect 599 543 600 547
rect 594 542 600 543
rect 598 539 604 540
rect 598 535 599 539
rect 603 535 604 539
rect 598 534 604 535
rect 111 530 115 531
rect 111 525 115 526
rect 335 530 339 531
rect 335 525 339 526
rect 423 530 427 531
rect 423 525 427 526
rect 455 530 459 531
rect 455 525 459 526
rect 511 530 515 531
rect 511 525 515 526
rect 535 530 539 531
rect 535 525 539 526
rect 591 530 595 531
rect 591 525 595 526
rect 112 497 114 525
rect 290 523 296 524
rect 290 519 291 523
rect 295 519 296 523
rect 290 518 296 519
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 112 447 114 474
rect 111 446 115 447
rect 111 441 115 442
rect 223 446 227 447
rect 223 441 227 442
rect 112 422 114 441
rect 224 425 226 441
rect 222 424 228 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 222 420 223 424
rect 227 420 228 424
rect 222 419 228 420
rect 110 416 116 417
rect 292 416 294 518
rect 336 515 338 525
rect 386 523 392 524
rect 386 519 387 523
rect 391 519 392 523
rect 386 518 392 519
rect 334 514 340 515
rect 334 510 335 514
rect 339 510 340 514
rect 334 509 340 510
rect 388 488 390 518
rect 424 515 426 525
rect 474 523 480 524
rect 474 519 475 523
rect 479 519 480 523
rect 474 518 480 519
rect 422 514 428 515
rect 422 510 423 514
rect 427 510 428 514
rect 422 509 428 510
rect 476 488 478 518
rect 512 515 514 525
rect 562 523 568 524
rect 562 519 563 523
rect 567 519 568 523
rect 562 518 568 519
rect 510 514 516 515
rect 510 510 511 514
rect 515 510 516 514
rect 510 509 516 510
rect 564 488 566 518
rect 592 515 594 525
rect 590 514 596 515
rect 590 510 591 514
rect 595 510 596 514
rect 590 509 596 510
rect 600 488 602 534
rect 616 531 618 553
rect 676 548 678 582
rect 694 558 700 559
rect 694 554 695 558
rect 699 554 700 558
rect 694 553 700 554
rect 674 547 680 548
rect 674 543 675 547
rect 679 543 680 547
rect 674 542 680 543
rect 696 531 698 553
rect 756 548 758 582
rect 782 558 788 559
rect 782 554 783 558
rect 787 554 788 558
rect 782 553 788 554
rect 754 547 760 548
rect 754 543 755 547
rect 759 543 760 547
rect 754 542 760 543
rect 784 531 786 553
rect 864 532 866 582
rect 878 558 884 559
rect 878 554 879 558
rect 883 554 884 558
rect 878 553 884 554
rect 862 531 868 532
rect 880 531 882 553
rect 940 548 942 582
rect 966 558 972 559
rect 966 554 967 558
rect 971 554 972 558
rect 966 553 972 554
rect 1054 558 1060 559
rect 1054 554 1055 558
rect 1059 554 1060 558
rect 1054 553 1060 554
rect 938 547 944 548
rect 938 543 939 547
rect 943 543 944 547
rect 938 542 944 543
rect 968 531 970 553
rect 1056 531 1058 553
rect 1116 548 1118 582
rect 1150 558 1156 559
rect 1150 554 1151 558
rect 1155 554 1156 558
rect 1150 553 1156 554
rect 1114 547 1120 548
rect 1114 543 1115 547
rect 1119 543 1120 547
rect 1114 542 1120 543
rect 1152 531 1154 553
rect 1212 548 1214 582
rect 1246 558 1252 559
rect 1246 554 1247 558
rect 1251 554 1252 558
rect 1246 553 1252 554
rect 1210 547 1216 548
rect 1210 543 1211 547
rect 1215 543 1216 547
rect 1210 542 1216 543
rect 1248 531 1250 553
rect 1308 548 1310 582
rect 1342 558 1348 559
rect 1342 554 1343 558
rect 1347 554 1348 558
rect 1342 553 1348 554
rect 1306 547 1312 548
rect 1306 543 1307 547
rect 1311 543 1312 547
rect 1306 542 1312 543
rect 1286 539 1292 540
rect 1286 535 1287 539
rect 1291 535 1292 539
rect 1286 534 1292 535
rect 615 530 619 531
rect 615 525 619 526
rect 671 530 675 531
rect 671 525 675 526
rect 695 530 699 531
rect 695 525 699 526
rect 751 530 755 531
rect 751 525 755 526
rect 783 530 787 531
rect 783 525 787 526
rect 839 530 843 531
rect 862 527 863 531
rect 867 527 868 531
rect 862 526 868 527
rect 879 530 883 531
rect 839 525 843 526
rect 879 525 883 526
rect 927 530 931 531
rect 927 525 931 526
rect 967 530 971 531
rect 967 525 971 526
rect 1015 530 1019 531
rect 1015 525 1019 526
rect 1055 530 1059 531
rect 1055 525 1059 526
rect 1103 530 1107 531
rect 1103 525 1107 526
rect 1151 530 1155 531
rect 1151 525 1155 526
rect 1191 530 1195 531
rect 1191 525 1195 526
rect 1247 530 1251 531
rect 1247 525 1251 526
rect 1279 530 1283 531
rect 1279 525 1283 526
rect 672 515 674 525
rect 722 523 728 524
rect 722 519 723 523
rect 727 519 728 523
rect 722 518 728 519
rect 670 514 676 515
rect 670 510 671 514
rect 675 510 676 514
rect 670 509 676 510
rect 724 488 726 518
rect 752 515 754 525
rect 840 515 842 525
rect 854 523 860 524
rect 854 519 855 523
rect 859 519 860 523
rect 854 518 860 519
rect 890 523 896 524
rect 890 519 891 523
rect 895 519 896 523
rect 890 518 896 519
rect 750 514 756 515
rect 750 510 751 514
rect 755 510 756 514
rect 750 509 756 510
rect 838 514 844 515
rect 838 510 839 514
rect 843 510 844 514
rect 838 509 844 510
rect 386 487 392 488
rect 386 483 387 487
rect 391 483 392 487
rect 386 482 392 483
rect 474 487 480 488
rect 474 483 475 487
rect 479 483 480 487
rect 474 482 480 483
rect 562 487 568 488
rect 562 483 563 487
rect 567 483 568 487
rect 562 482 568 483
rect 598 487 604 488
rect 598 483 599 487
rect 603 483 604 487
rect 598 482 604 483
rect 722 487 728 488
rect 722 483 723 487
rect 727 483 728 487
rect 722 482 728 483
rect 326 476 332 477
rect 326 472 327 476
rect 331 472 332 476
rect 326 471 332 472
rect 414 476 420 477
rect 414 472 415 476
rect 419 472 420 476
rect 414 471 420 472
rect 502 476 508 477
rect 502 472 503 476
rect 507 472 508 476
rect 502 471 508 472
rect 582 476 588 477
rect 582 472 583 476
rect 587 472 588 476
rect 582 471 588 472
rect 662 476 668 477
rect 662 472 663 476
rect 667 472 668 476
rect 662 471 668 472
rect 742 476 748 477
rect 742 472 743 476
rect 747 472 748 476
rect 742 471 748 472
rect 830 476 836 477
rect 830 472 831 476
rect 835 472 836 476
rect 830 471 836 472
rect 328 447 330 471
rect 416 447 418 471
rect 504 447 506 471
rect 584 447 586 471
rect 664 447 666 471
rect 744 447 746 471
rect 832 447 834 471
rect 327 446 331 447
rect 327 441 331 442
rect 335 446 339 447
rect 335 441 339 442
rect 415 446 419 447
rect 415 441 419 442
rect 447 446 451 447
rect 447 441 451 442
rect 503 446 507 447
rect 503 441 507 442
rect 559 446 563 447
rect 559 441 563 442
rect 583 446 587 447
rect 583 441 587 442
rect 663 446 667 447
rect 663 441 667 442
rect 743 446 747 447
rect 743 441 747 442
rect 759 446 763 447
rect 759 441 763 442
rect 831 446 835 447
rect 831 441 835 442
rect 847 446 851 447
rect 847 441 851 442
rect 336 425 338 441
rect 448 425 450 441
rect 560 425 562 441
rect 664 425 666 441
rect 760 425 762 441
rect 848 425 850 441
rect 334 424 340 425
rect 334 420 335 424
rect 339 420 340 424
rect 334 419 340 420
rect 446 424 452 425
rect 446 420 447 424
rect 451 420 452 424
rect 446 419 452 420
rect 558 424 564 425
rect 558 420 559 424
rect 563 420 564 424
rect 558 419 564 420
rect 662 424 668 425
rect 662 420 663 424
rect 667 420 668 424
rect 662 419 668 420
rect 758 424 764 425
rect 758 420 759 424
rect 763 420 764 424
rect 758 419 764 420
rect 846 424 852 425
rect 846 420 847 424
rect 851 420 852 424
rect 846 419 852 420
rect 290 415 296 416
rect 290 411 291 415
rect 295 411 296 415
rect 290 410 296 411
rect 298 415 304 416
rect 298 411 299 415
rect 303 411 304 415
rect 298 410 304 411
rect 402 415 408 416
rect 402 411 403 415
rect 407 411 408 415
rect 402 410 408 411
rect 730 415 736 416
rect 730 411 731 415
rect 735 411 736 415
rect 856 412 858 518
rect 892 488 894 518
rect 928 515 930 525
rect 978 523 984 524
rect 978 519 979 523
rect 983 519 984 523
rect 978 518 984 519
rect 926 514 932 515
rect 926 510 927 514
rect 931 510 932 514
rect 926 509 932 510
rect 980 488 982 518
rect 1016 515 1018 525
rect 1066 523 1072 524
rect 1066 519 1067 523
rect 1071 519 1072 523
rect 1066 518 1072 519
rect 1014 514 1020 515
rect 1014 510 1015 514
rect 1019 510 1020 514
rect 1014 509 1020 510
rect 1068 488 1070 518
rect 1104 515 1106 525
rect 1182 523 1188 524
rect 1182 519 1183 523
rect 1187 519 1188 523
rect 1182 518 1188 519
rect 1102 514 1108 515
rect 1102 510 1103 514
rect 1107 510 1108 514
rect 1102 509 1108 510
rect 1184 488 1186 518
rect 1192 515 1194 525
rect 1270 523 1276 524
rect 1270 519 1271 523
rect 1275 519 1276 523
rect 1270 518 1276 519
rect 1190 514 1196 515
rect 1190 510 1191 514
rect 1195 510 1196 514
rect 1190 509 1196 510
rect 1272 488 1274 518
rect 1280 515 1282 525
rect 1278 514 1284 515
rect 1278 510 1279 514
rect 1283 510 1284 514
rect 1278 509 1284 510
rect 1288 488 1290 534
rect 1344 531 1346 553
rect 1404 548 1406 582
rect 1830 576 1836 577
rect 1830 572 1831 576
rect 1835 572 1836 576
rect 1830 571 1836 572
rect 1438 558 1444 559
rect 1438 554 1439 558
rect 1443 554 1444 558
rect 1438 553 1444 554
rect 1402 547 1408 548
rect 1402 543 1403 547
rect 1407 543 1408 547
rect 1402 542 1408 543
rect 1440 531 1442 553
rect 1832 531 1834 571
rect 1872 566 1874 585
rect 2264 569 2266 585
rect 2344 569 2346 585
rect 2424 569 2426 585
rect 2504 569 2506 585
rect 2262 568 2268 569
rect 1870 565 1876 566
rect 1870 561 1871 565
rect 1875 561 1876 565
rect 2262 564 2263 568
rect 2267 564 2268 568
rect 2262 563 2268 564
rect 2342 568 2348 569
rect 2342 564 2343 568
rect 2347 564 2348 568
rect 2342 563 2348 564
rect 2422 568 2428 569
rect 2422 564 2423 568
rect 2427 564 2428 568
rect 2422 563 2428 564
rect 2502 568 2508 569
rect 2502 564 2503 568
rect 2507 564 2508 568
rect 2502 563 2508 564
rect 1870 560 1876 561
rect 2330 559 2336 560
rect 2330 555 2331 559
rect 2335 555 2336 559
rect 2330 554 2336 555
rect 2410 559 2416 560
rect 2410 555 2411 559
rect 2415 555 2416 559
rect 2410 554 2416 555
rect 2490 559 2496 560
rect 2490 555 2491 559
rect 2495 555 2496 559
rect 2490 554 2496 555
rect 1870 548 1876 549
rect 1870 544 1871 548
rect 1875 544 1876 548
rect 1870 543 1876 544
rect 2283 548 2287 549
rect 2283 543 2287 544
rect 1343 530 1347 531
rect 1343 525 1347 526
rect 1439 530 1443 531
rect 1439 525 1443 526
rect 1831 530 1835 531
rect 1831 525 1835 526
rect 1832 497 1834 525
rect 1872 507 1874 543
rect 2270 530 2276 531
rect 2270 526 2271 530
rect 2275 526 2276 530
rect 2270 525 2276 526
rect 2272 507 2274 525
rect 2284 520 2286 543
rect 2332 520 2334 554
rect 2350 530 2356 531
rect 2350 526 2351 530
rect 2355 526 2356 530
rect 2350 525 2356 526
rect 2282 519 2288 520
rect 2282 515 2283 519
rect 2287 515 2288 519
rect 2282 514 2288 515
rect 2330 519 2336 520
rect 2330 515 2331 519
rect 2335 515 2336 519
rect 2330 514 2336 515
rect 2352 507 2354 525
rect 2412 520 2414 554
rect 2430 530 2436 531
rect 2430 526 2431 530
rect 2435 526 2436 530
rect 2430 525 2436 526
rect 2410 519 2416 520
rect 2410 515 2411 519
rect 2415 515 2416 519
rect 2410 514 2416 515
rect 2432 507 2434 525
rect 2492 520 2494 554
rect 2540 549 2542 590
rect 2591 585 2595 586
rect 2599 590 2603 591
rect 2599 585 2603 586
rect 2695 590 2699 591
rect 2695 585 2699 586
rect 2727 590 2731 591
rect 2727 585 2731 586
rect 2592 569 2594 585
rect 2696 569 2698 585
rect 2590 568 2596 569
rect 2590 564 2591 568
rect 2595 564 2596 568
rect 2590 563 2596 564
rect 2694 568 2700 569
rect 2694 564 2695 568
rect 2699 564 2700 568
rect 2694 563 2700 564
rect 2570 559 2576 560
rect 2570 555 2571 559
rect 2575 555 2576 559
rect 2570 554 2576 555
rect 2658 559 2664 560
rect 2658 555 2659 559
rect 2663 555 2664 559
rect 2658 554 2664 555
rect 2562 551 2568 552
rect 2539 548 2543 549
rect 2562 547 2563 551
rect 2567 547 2568 551
rect 2562 546 2568 547
rect 2539 543 2543 544
rect 2510 530 2516 531
rect 2510 526 2511 530
rect 2515 526 2516 530
rect 2510 525 2516 526
rect 2490 519 2496 520
rect 2490 515 2491 519
rect 2495 515 2496 519
rect 2490 514 2496 515
rect 2512 507 2514 525
rect 1871 506 1875 507
rect 1871 501 1875 502
rect 2191 506 2195 507
rect 2191 501 2195 502
rect 2271 506 2275 507
rect 2271 501 2275 502
rect 2287 506 2291 507
rect 2287 501 2291 502
rect 2351 506 2355 507
rect 2351 501 2355 502
rect 2383 506 2387 507
rect 2383 501 2387 502
rect 2431 506 2435 507
rect 2431 501 2435 502
rect 2487 506 2491 507
rect 2487 501 2491 502
rect 2511 506 2515 507
rect 2511 501 2515 502
rect 1830 496 1836 497
rect 1830 492 1831 496
rect 1835 492 1836 496
rect 1830 491 1836 492
rect 890 487 896 488
rect 890 483 891 487
rect 895 483 896 487
rect 890 482 896 483
rect 978 487 984 488
rect 978 483 979 487
rect 983 483 984 487
rect 978 482 984 483
rect 1066 487 1072 488
rect 1066 483 1067 487
rect 1071 483 1072 487
rect 1066 482 1072 483
rect 1182 487 1188 488
rect 1182 483 1183 487
rect 1187 483 1188 487
rect 1182 482 1188 483
rect 1270 487 1276 488
rect 1270 483 1271 487
rect 1275 483 1276 487
rect 1270 482 1276 483
rect 1286 487 1292 488
rect 1286 483 1287 487
rect 1291 483 1292 487
rect 1286 482 1292 483
rect 1830 479 1836 480
rect 918 476 924 477
rect 918 472 919 476
rect 923 472 924 476
rect 918 471 924 472
rect 1006 476 1012 477
rect 1006 472 1007 476
rect 1011 472 1012 476
rect 1006 471 1012 472
rect 1094 476 1100 477
rect 1094 472 1095 476
rect 1099 472 1100 476
rect 1094 471 1100 472
rect 1182 476 1188 477
rect 1182 472 1183 476
rect 1187 472 1188 476
rect 1182 471 1188 472
rect 1270 476 1276 477
rect 1270 472 1271 476
rect 1275 472 1276 476
rect 1830 475 1831 479
rect 1835 475 1836 479
rect 1830 474 1836 475
rect 1270 471 1276 472
rect 920 447 922 471
rect 1008 447 1010 471
rect 1096 447 1098 471
rect 1184 447 1186 471
rect 1272 447 1274 471
rect 1832 447 1834 474
rect 1872 473 1874 501
rect 2192 491 2194 501
rect 2250 499 2256 500
rect 2250 495 2251 499
rect 2255 495 2256 499
rect 2250 494 2256 495
rect 2190 490 2196 491
rect 2190 486 2191 490
rect 2195 486 2196 490
rect 2190 485 2196 486
rect 1870 472 1876 473
rect 1870 468 1871 472
rect 1875 468 1876 472
rect 1870 467 1876 468
rect 2252 464 2254 494
rect 2288 491 2290 501
rect 2384 491 2386 501
rect 2442 499 2448 500
rect 2442 495 2443 499
rect 2447 495 2448 499
rect 2442 494 2448 495
rect 2286 490 2292 491
rect 2286 486 2287 490
rect 2291 486 2292 490
rect 2286 485 2292 486
rect 2382 490 2388 491
rect 2382 486 2383 490
rect 2387 486 2388 490
rect 2382 485 2388 486
rect 2444 464 2446 494
rect 2488 491 2490 501
rect 2564 500 2566 546
rect 2572 520 2574 554
rect 2598 530 2604 531
rect 2598 526 2599 530
rect 2603 526 2604 530
rect 2598 525 2604 526
rect 2570 519 2576 520
rect 2570 515 2571 519
rect 2575 515 2576 519
rect 2570 514 2576 515
rect 2600 507 2602 525
rect 2660 520 2662 554
rect 2754 551 2760 552
rect 2754 547 2755 551
rect 2759 547 2760 551
rect 2754 546 2760 547
rect 2702 530 2708 531
rect 2702 526 2703 530
rect 2707 526 2708 530
rect 2702 525 2708 526
rect 2658 519 2664 520
rect 2658 515 2659 519
rect 2663 515 2664 519
rect 2658 514 2664 515
rect 2704 507 2706 525
rect 2583 506 2587 507
rect 2583 501 2587 502
rect 2599 506 2603 507
rect 2599 501 2603 502
rect 2687 506 2691 507
rect 2687 501 2691 502
rect 2703 506 2707 507
rect 2703 501 2707 502
rect 2562 499 2568 500
rect 2562 495 2563 499
rect 2567 495 2568 499
rect 2562 494 2568 495
rect 2584 491 2586 501
rect 2642 499 2648 500
rect 2642 495 2643 499
rect 2647 495 2648 499
rect 2642 494 2648 495
rect 2486 490 2492 491
rect 2486 486 2487 490
rect 2491 486 2492 490
rect 2486 485 2492 486
rect 2582 490 2588 491
rect 2582 486 2583 490
rect 2587 486 2588 490
rect 2582 485 2588 486
rect 2644 464 2646 494
rect 2688 491 2690 501
rect 2756 500 2758 546
rect 2788 520 2790 618
rect 2854 612 2860 613
rect 2854 608 2855 612
rect 2859 608 2860 612
rect 2854 607 2860 608
rect 2982 612 2988 613
rect 2982 608 2983 612
rect 2987 608 2988 612
rect 2982 607 2988 608
rect 2856 591 2858 607
rect 2984 591 2986 607
rect 2815 590 2819 591
rect 2815 585 2819 586
rect 2855 590 2859 591
rect 2855 585 2859 586
rect 2959 590 2963 591
rect 2959 585 2963 586
rect 2983 590 2987 591
rect 2983 585 2987 586
rect 2816 569 2818 585
rect 2960 569 2962 585
rect 2814 568 2820 569
rect 2814 564 2815 568
rect 2819 564 2820 568
rect 2814 563 2820 564
rect 2958 568 2964 569
rect 2958 564 2959 568
rect 2963 564 2964 568
rect 2958 563 2964 564
rect 2894 559 2900 560
rect 2894 555 2895 559
rect 2899 555 2900 559
rect 2894 554 2900 555
rect 3026 559 3032 560
rect 3026 555 3027 559
rect 3031 555 3032 559
rect 3026 554 3032 555
rect 2822 530 2828 531
rect 2822 526 2823 530
rect 2827 526 2828 530
rect 2822 525 2828 526
rect 2786 519 2792 520
rect 2786 515 2787 519
rect 2791 515 2792 519
rect 2786 514 2792 515
rect 2824 507 2826 525
rect 2896 520 2898 554
rect 2966 530 2972 531
rect 2966 526 2967 530
rect 2971 526 2972 530
rect 2966 525 2972 526
rect 2894 519 2900 520
rect 2894 515 2895 519
rect 2899 515 2900 519
rect 2894 514 2900 515
rect 2968 507 2970 525
rect 3028 508 3030 554
rect 3044 520 3046 618
rect 3110 612 3116 613
rect 3110 608 3111 612
rect 3115 608 3116 612
rect 3110 607 3116 608
rect 3238 612 3244 613
rect 3238 608 3239 612
rect 3243 608 3244 612
rect 3238 607 3244 608
rect 3366 612 3372 613
rect 3366 608 3367 612
rect 3371 608 3372 612
rect 3366 607 3372 608
rect 3112 591 3114 607
rect 3240 591 3242 607
rect 3368 591 3370 607
rect 3111 590 3115 591
rect 3111 585 3115 586
rect 3239 590 3243 591
rect 3239 585 3243 586
rect 3279 590 3283 591
rect 3279 585 3283 586
rect 3367 590 3371 591
rect 3367 585 3371 586
rect 3112 569 3114 585
rect 3280 569 3282 585
rect 3110 568 3116 569
rect 3110 564 3111 568
rect 3115 564 3116 568
rect 3110 563 3116 564
rect 3278 568 3284 569
rect 3278 564 3279 568
rect 3283 564 3284 568
rect 3278 563 3284 564
rect 3118 530 3124 531
rect 3118 526 3119 530
rect 3123 526 3124 530
rect 3118 525 3124 526
rect 3286 530 3292 531
rect 3286 526 3287 530
rect 3291 526 3292 530
rect 3286 525 3292 526
rect 3042 519 3048 520
rect 3042 515 3043 519
rect 3047 515 3048 519
rect 3042 514 3048 515
rect 3026 507 3032 508
rect 3120 507 3122 525
rect 3288 507 3290 525
rect 3428 520 3430 618
rect 3502 612 3508 613
rect 3502 608 3503 612
rect 3507 608 3508 612
rect 3502 607 3508 608
rect 3504 591 3506 607
rect 3447 590 3451 591
rect 3447 585 3451 586
rect 3503 590 3507 591
rect 3503 585 3507 586
rect 3448 569 3450 585
rect 3446 568 3452 569
rect 3446 564 3447 568
rect 3451 564 3452 568
rect 3446 563 3452 564
rect 3528 560 3530 654
rect 3592 633 3594 661
rect 3590 632 3596 633
rect 3590 628 3591 632
rect 3595 628 3596 632
rect 3590 627 3596 628
rect 3590 615 3596 616
rect 3590 611 3591 615
rect 3595 611 3596 615
rect 3590 610 3596 611
rect 3592 591 3594 610
rect 3591 590 3595 591
rect 3591 585 3595 586
rect 3592 566 3594 585
rect 3590 565 3596 566
rect 3590 561 3591 565
rect 3595 561 3596 565
rect 3590 560 3596 561
rect 3526 559 3532 560
rect 3526 555 3527 559
rect 3531 555 3532 559
rect 3526 554 3532 555
rect 3590 548 3596 549
rect 3590 544 3591 548
rect 3595 544 3596 548
rect 3590 543 3596 544
rect 3454 530 3460 531
rect 3454 526 3455 530
rect 3459 526 3460 530
rect 3454 525 3460 526
rect 3326 519 3332 520
rect 3326 515 3327 519
rect 3331 515 3332 519
rect 3326 514 3332 515
rect 3426 519 3432 520
rect 3426 515 3427 519
rect 3431 515 3432 519
rect 3426 514 3432 515
rect 2791 506 2795 507
rect 2791 501 2795 502
rect 2823 506 2827 507
rect 2823 501 2827 502
rect 2911 506 2915 507
rect 2911 501 2915 502
rect 2967 506 2971 507
rect 3026 503 3027 507
rect 3031 503 3032 507
rect 3026 502 3032 503
rect 3039 506 3043 507
rect 2967 501 2971 502
rect 3039 501 3043 502
rect 3119 506 3123 507
rect 3119 501 3123 502
rect 3175 506 3179 507
rect 3175 501 3179 502
rect 3287 506 3291 507
rect 3287 501 3291 502
rect 3319 506 3323 507
rect 3319 501 3323 502
rect 2754 499 2760 500
rect 2754 495 2755 499
rect 2759 495 2760 499
rect 2754 494 2760 495
rect 2792 491 2794 501
rect 2842 499 2848 500
rect 2842 495 2843 499
rect 2847 495 2848 499
rect 2842 494 2848 495
rect 2686 490 2692 491
rect 2686 486 2687 490
rect 2691 486 2692 490
rect 2686 485 2692 486
rect 2790 490 2796 491
rect 2790 486 2791 490
rect 2795 486 2796 490
rect 2790 485 2796 486
rect 2844 464 2846 494
rect 2912 491 2914 501
rect 3030 499 3036 500
rect 3030 495 3031 499
rect 3035 495 3036 499
rect 3030 494 3036 495
rect 2910 490 2916 491
rect 2910 486 2911 490
rect 2915 486 2916 490
rect 2910 485 2916 486
rect 3032 464 3034 494
rect 3040 491 3042 501
rect 3090 499 3096 500
rect 3090 495 3091 499
rect 3095 495 3096 499
rect 3090 494 3096 495
rect 3038 490 3044 491
rect 3038 486 3039 490
rect 3043 486 3044 490
rect 3038 485 3044 486
rect 3092 464 3094 494
rect 3176 491 3178 501
rect 3226 499 3232 500
rect 3226 495 3227 499
rect 3231 495 3232 499
rect 3226 494 3232 495
rect 3174 490 3180 491
rect 3174 486 3175 490
rect 3179 486 3180 490
rect 3174 485 3180 486
rect 3228 464 3230 494
rect 3320 491 3322 501
rect 3318 490 3324 491
rect 3318 486 3319 490
rect 3323 486 3324 490
rect 3318 485 3324 486
rect 3328 464 3330 514
rect 3456 507 3458 525
rect 3592 507 3594 543
rect 3455 506 3459 507
rect 3455 501 3459 502
rect 3471 506 3475 507
rect 3471 501 3475 502
rect 3591 506 3595 507
rect 3591 501 3595 502
rect 3390 499 3396 500
rect 3390 495 3391 499
rect 3395 495 3396 499
rect 3390 494 3396 495
rect 2250 463 2256 464
rect 2250 459 2251 463
rect 2255 459 2256 463
rect 2250 458 2256 459
rect 2442 463 2448 464
rect 2442 459 2443 463
rect 2447 459 2448 463
rect 2442 458 2448 459
rect 2642 463 2648 464
rect 2642 459 2643 463
rect 2647 459 2648 463
rect 2642 458 2648 459
rect 2842 463 2848 464
rect 2842 459 2843 463
rect 2847 459 2848 463
rect 2842 458 2848 459
rect 3030 463 3036 464
rect 3030 459 3031 463
rect 3035 459 3036 463
rect 3030 458 3036 459
rect 3090 463 3096 464
rect 3090 459 3091 463
rect 3095 459 3096 463
rect 3090 458 3096 459
rect 3226 463 3232 464
rect 3226 459 3227 463
rect 3231 459 3232 463
rect 3226 458 3232 459
rect 3326 463 3332 464
rect 3326 459 3327 463
rect 3331 459 3332 463
rect 3326 458 3332 459
rect 1870 455 1876 456
rect 1870 451 1871 455
rect 1875 451 1876 455
rect 1870 450 1876 451
rect 2182 452 2188 453
rect 919 446 923 447
rect 919 441 923 442
rect 935 446 939 447
rect 935 441 939 442
rect 1007 446 1011 447
rect 1007 441 1011 442
rect 1023 446 1027 447
rect 1023 441 1027 442
rect 1095 446 1099 447
rect 1095 441 1099 442
rect 1111 446 1115 447
rect 1111 441 1115 442
rect 1183 446 1187 447
rect 1183 441 1187 442
rect 1199 446 1203 447
rect 1199 441 1203 442
rect 1271 446 1275 447
rect 1271 441 1275 442
rect 1295 446 1299 447
rect 1295 441 1299 442
rect 1831 446 1835 447
rect 1831 441 1835 442
rect 936 425 938 441
rect 1024 425 1026 441
rect 1112 425 1114 441
rect 1200 425 1202 441
rect 1296 425 1298 441
rect 934 424 940 425
rect 934 420 935 424
rect 939 420 940 424
rect 934 419 940 420
rect 1022 424 1028 425
rect 1022 420 1023 424
rect 1027 420 1028 424
rect 1022 419 1028 420
rect 1110 424 1116 425
rect 1110 420 1111 424
rect 1115 420 1116 424
rect 1110 419 1116 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1294 424 1300 425
rect 1294 420 1295 424
rect 1299 420 1300 424
rect 1832 422 1834 441
rect 1872 427 1874 450
rect 2182 448 2183 452
rect 2187 448 2188 452
rect 2182 447 2188 448
rect 2278 452 2284 453
rect 2278 448 2279 452
rect 2283 448 2284 452
rect 2278 447 2284 448
rect 2374 452 2380 453
rect 2374 448 2375 452
rect 2379 448 2380 452
rect 2374 447 2380 448
rect 2478 452 2484 453
rect 2478 448 2479 452
rect 2483 448 2484 452
rect 2478 447 2484 448
rect 2574 452 2580 453
rect 2574 448 2575 452
rect 2579 448 2580 452
rect 2574 447 2580 448
rect 2678 452 2684 453
rect 2678 448 2679 452
rect 2683 448 2684 452
rect 2678 447 2684 448
rect 2782 452 2788 453
rect 2782 448 2783 452
rect 2787 448 2788 452
rect 2782 447 2788 448
rect 2902 452 2908 453
rect 2902 448 2903 452
rect 2907 448 2908 452
rect 2902 447 2908 448
rect 3030 452 3036 453
rect 3030 448 3031 452
rect 3035 448 3036 452
rect 3030 447 3036 448
rect 3166 452 3172 453
rect 3166 448 3167 452
rect 3171 448 3172 452
rect 3166 447 3172 448
rect 3310 452 3316 453
rect 3310 448 3311 452
rect 3315 448 3316 452
rect 3310 447 3316 448
rect 1990 435 1996 436
rect 1990 431 1991 435
rect 1995 431 1996 435
rect 1990 430 1996 431
rect 1871 426 1875 427
rect 1294 419 1300 420
rect 1830 421 1836 422
rect 1871 421 1875 422
rect 1975 426 1979 427
rect 1975 421 1979 422
rect 1830 417 1831 421
rect 1835 417 1836 421
rect 1830 416 1836 417
rect 914 415 920 416
rect 730 410 736 411
rect 854 411 860 412
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 112 359 114 399
rect 230 386 236 387
rect 230 382 231 386
rect 235 382 236 386
rect 230 381 236 382
rect 232 359 234 381
rect 300 376 302 410
rect 342 386 348 387
rect 342 382 343 386
rect 347 382 348 386
rect 342 381 348 382
rect 298 375 304 376
rect 298 371 299 375
rect 303 371 304 375
rect 298 370 304 371
rect 344 359 346 381
rect 404 376 406 410
rect 454 386 460 387
rect 454 382 455 386
rect 459 382 460 386
rect 454 381 460 382
rect 566 386 572 387
rect 566 382 567 386
rect 571 382 572 386
rect 566 381 572 382
rect 670 386 676 387
rect 670 382 671 386
rect 675 382 676 386
rect 670 381 676 382
rect 402 375 408 376
rect 402 371 403 375
rect 407 371 408 375
rect 402 370 408 371
rect 446 375 452 376
rect 446 371 447 375
rect 451 371 452 375
rect 446 370 452 371
rect 111 358 115 359
rect 111 353 115 354
rect 143 358 147 359
rect 143 353 147 354
rect 231 358 235 359
rect 231 353 235 354
rect 263 358 267 359
rect 263 353 267 354
rect 343 358 347 359
rect 343 353 347 354
rect 399 358 403 359
rect 399 353 403 354
rect 112 325 114 353
rect 144 343 146 353
rect 194 351 200 352
rect 194 347 195 351
rect 199 347 200 351
rect 194 346 200 347
rect 142 342 148 343
rect 142 338 143 342
rect 147 338 148 342
rect 142 337 148 338
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 110 319 116 320
rect 196 316 198 346
rect 264 343 266 353
rect 314 351 320 352
rect 314 347 315 351
rect 319 347 320 351
rect 314 346 320 347
rect 262 342 268 343
rect 262 338 263 342
rect 267 338 268 342
rect 262 337 268 338
rect 316 316 318 346
rect 400 343 402 353
rect 398 342 404 343
rect 398 338 399 342
rect 403 338 404 342
rect 398 337 404 338
rect 448 316 450 370
rect 456 359 458 381
rect 568 359 570 381
rect 672 359 674 381
rect 732 376 734 410
rect 854 407 855 411
rect 859 407 860 411
rect 914 411 915 415
rect 919 411 920 415
rect 914 410 920 411
rect 1002 415 1008 416
rect 1002 411 1003 415
rect 1007 411 1008 415
rect 1002 410 1008 411
rect 1090 415 1096 416
rect 1090 411 1091 415
rect 1095 411 1096 415
rect 1090 410 1096 411
rect 1266 415 1272 416
rect 1266 411 1267 415
rect 1271 411 1272 415
rect 1266 410 1272 411
rect 854 406 860 407
rect 766 386 772 387
rect 766 382 767 386
rect 771 382 772 386
rect 766 381 772 382
rect 854 386 860 387
rect 854 382 855 386
rect 859 382 860 386
rect 854 381 860 382
rect 730 375 736 376
rect 730 371 731 375
rect 735 371 736 375
rect 730 370 736 371
rect 768 359 770 381
rect 856 359 858 381
rect 916 376 918 410
rect 942 386 948 387
rect 942 382 943 386
rect 947 382 948 386
rect 942 381 948 382
rect 914 375 920 376
rect 914 371 915 375
rect 919 371 920 375
rect 914 370 920 371
rect 944 359 946 381
rect 1004 376 1006 410
rect 1030 386 1036 387
rect 1030 382 1031 386
rect 1035 382 1036 386
rect 1030 381 1036 382
rect 1002 375 1008 376
rect 1002 371 1003 375
rect 1007 371 1008 375
rect 1002 370 1008 371
rect 1032 359 1034 381
rect 1092 376 1094 410
rect 1170 407 1176 408
rect 1170 403 1171 407
rect 1175 403 1176 407
rect 1170 402 1176 403
rect 1118 386 1124 387
rect 1118 382 1119 386
rect 1123 382 1124 386
rect 1118 381 1124 382
rect 1090 375 1096 376
rect 1090 371 1091 375
rect 1095 371 1096 375
rect 1090 370 1096 371
rect 1120 359 1122 381
rect 1172 376 1174 402
rect 1206 386 1212 387
rect 1206 382 1207 386
rect 1211 382 1212 386
rect 1206 381 1212 382
rect 1170 375 1176 376
rect 1170 371 1171 375
rect 1175 371 1176 375
rect 1170 370 1176 371
rect 1178 375 1184 376
rect 1178 371 1179 375
rect 1183 371 1184 375
rect 1178 370 1184 371
rect 455 358 459 359
rect 455 353 459 354
rect 535 358 539 359
rect 535 353 539 354
rect 567 358 571 359
rect 567 353 571 354
rect 671 358 675 359
rect 671 353 675 354
rect 767 358 771 359
rect 767 353 771 354
rect 791 358 795 359
rect 791 353 795 354
rect 855 358 859 359
rect 855 353 859 354
rect 911 358 915 359
rect 911 353 915 354
rect 943 358 947 359
rect 943 353 947 354
rect 1023 358 1027 359
rect 1023 353 1027 354
rect 1031 358 1035 359
rect 1031 353 1035 354
rect 1119 358 1123 359
rect 1119 353 1123 354
rect 1127 358 1131 359
rect 1127 353 1131 354
rect 536 343 538 353
rect 586 351 592 352
rect 586 347 587 351
rect 591 347 592 351
rect 586 346 592 347
rect 534 342 540 343
rect 534 338 535 342
rect 539 338 540 342
rect 534 337 540 338
rect 588 316 590 346
rect 672 343 674 353
rect 722 351 728 352
rect 722 347 723 351
rect 727 347 728 351
rect 722 346 728 347
rect 670 342 676 343
rect 670 338 671 342
rect 675 338 676 342
rect 670 337 676 338
rect 724 316 726 346
rect 792 343 794 353
rect 912 343 914 353
rect 962 351 968 352
rect 962 347 963 351
rect 967 347 968 351
rect 962 346 968 347
rect 790 342 796 343
rect 790 338 791 342
rect 795 338 796 342
rect 790 337 796 338
rect 910 342 916 343
rect 910 338 911 342
rect 915 338 916 342
rect 910 337 916 338
rect 964 316 966 346
rect 1024 343 1026 353
rect 1074 351 1080 352
rect 1074 347 1075 351
rect 1079 347 1080 351
rect 1074 346 1080 347
rect 1022 342 1028 343
rect 1022 338 1023 342
rect 1027 338 1028 342
rect 1022 337 1028 338
rect 1076 316 1078 346
rect 1128 343 1130 353
rect 1126 342 1132 343
rect 1126 338 1127 342
rect 1131 338 1132 342
rect 1126 337 1132 338
rect 1180 316 1182 370
rect 1208 359 1210 381
rect 1268 376 1270 410
rect 1830 404 1836 405
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 1872 402 1874 421
rect 1976 405 1978 421
rect 1974 404 1980 405
rect 1830 399 1836 400
rect 1870 401 1876 402
rect 1302 386 1308 387
rect 1302 382 1303 386
rect 1307 382 1308 386
rect 1302 381 1308 382
rect 1266 375 1272 376
rect 1266 371 1267 375
rect 1271 371 1272 375
rect 1266 370 1272 371
rect 1238 359 1244 360
rect 1304 359 1306 381
rect 1446 359 1452 360
rect 1832 359 1834 399
rect 1870 397 1871 401
rect 1875 397 1876 401
rect 1974 400 1975 404
rect 1979 400 1980 404
rect 1974 399 1980 400
rect 1870 396 1876 397
rect 1870 384 1876 385
rect 1870 380 1871 384
rect 1875 380 1876 384
rect 1870 379 1876 380
rect 1207 358 1211 359
rect 1207 353 1211 354
rect 1231 358 1235 359
rect 1238 355 1239 359
rect 1243 355 1244 359
rect 1238 354 1244 355
rect 1303 358 1307 359
rect 1231 353 1235 354
rect 1232 343 1234 353
rect 1230 342 1236 343
rect 1230 338 1231 342
rect 1235 338 1236 342
rect 1230 337 1236 338
rect 1240 316 1242 354
rect 1303 353 1307 354
rect 1335 358 1339 359
rect 1335 353 1339 354
rect 1439 358 1443 359
rect 1446 355 1447 359
rect 1451 355 1452 359
rect 1446 354 1452 355
rect 1831 358 1835 359
rect 1439 353 1443 354
rect 1310 351 1316 352
rect 1310 347 1311 351
rect 1315 347 1316 351
rect 1310 346 1316 347
rect 194 315 200 316
rect 194 311 195 315
rect 199 311 200 315
rect 194 310 200 311
rect 314 315 320 316
rect 314 311 315 315
rect 319 311 320 315
rect 314 310 320 311
rect 446 315 452 316
rect 446 311 447 315
rect 451 311 452 315
rect 446 310 452 311
rect 586 315 592 316
rect 586 311 587 315
rect 591 311 592 315
rect 586 310 592 311
rect 722 315 728 316
rect 722 311 723 315
rect 727 311 728 315
rect 722 310 728 311
rect 838 315 844 316
rect 838 311 839 315
rect 843 311 844 315
rect 838 310 844 311
rect 962 315 968 316
rect 962 311 963 315
rect 967 311 968 315
rect 962 310 968 311
rect 1074 315 1080 316
rect 1074 311 1075 315
rect 1079 311 1080 315
rect 1074 310 1080 311
rect 1178 315 1184 316
rect 1178 311 1179 315
rect 1183 311 1184 315
rect 1178 310 1184 311
rect 1238 315 1244 316
rect 1238 311 1239 315
rect 1243 311 1244 315
rect 1238 310 1244 311
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 110 302 116 303
rect 134 304 140 305
rect 112 275 114 302
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 254 304 260 305
rect 254 300 255 304
rect 259 300 260 304
rect 254 299 260 300
rect 390 304 396 305
rect 390 300 391 304
rect 395 300 396 304
rect 390 299 396 300
rect 526 304 532 305
rect 526 300 527 304
rect 531 300 532 304
rect 526 299 532 300
rect 662 304 668 305
rect 662 300 663 304
rect 667 300 668 304
rect 662 299 668 300
rect 782 304 788 305
rect 782 300 783 304
rect 787 300 788 304
rect 782 299 788 300
rect 136 275 138 299
rect 256 275 258 299
rect 392 275 394 299
rect 528 275 530 299
rect 664 275 666 299
rect 784 275 786 299
rect 111 274 115 275
rect 111 269 115 270
rect 135 274 139 275
rect 135 269 139 270
rect 247 274 251 275
rect 247 269 251 270
rect 255 274 259 275
rect 255 269 259 270
rect 391 274 395 275
rect 391 269 395 270
rect 527 274 531 275
rect 527 269 531 270
rect 543 274 547 275
rect 543 269 547 270
rect 663 274 667 275
rect 663 269 667 270
rect 695 274 699 275
rect 695 269 699 270
rect 783 274 787 275
rect 783 269 787 270
rect 112 250 114 269
rect 136 253 138 269
rect 248 253 250 269
rect 392 253 394 269
rect 544 253 546 269
rect 696 253 698 269
rect 134 252 140 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 246 252 252 253
rect 246 248 247 252
rect 251 248 252 252
rect 246 247 252 248
rect 390 252 396 253
rect 390 248 391 252
rect 395 248 396 252
rect 390 247 396 248
rect 542 252 548 253
rect 542 248 543 252
rect 547 248 548 252
rect 542 247 548 248
rect 694 252 700 253
rect 694 248 695 252
rect 699 248 700 252
rect 694 247 700 248
rect 110 244 116 245
rect 202 243 208 244
rect 202 239 203 243
rect 207 239 208 243
rect 202 238 208 239
rect 314 243 320 244
rect 314 239 315 243
rect 319 239 320 243
rect 314 238 320 239
rect 610 243 616 244
rect 610 239 611 243
rect 615 239 616 243
rect 610 238 616 239
rect 762 243 768 244
rect 762 239 763 243
rect 767 239 768 243
rect 762 238 768 239
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 110 227 116 228
rect 112 163 114 227
rect 142 214 148 215
rect 142 210 143 214
rect 147 210 148 214
rect 142 209 148 210
rect 144 163 146 209
rect 204 204 206 238
rect 254 214 260 215
rect 254 210 255 214
rect 259 210 260 214
rect 254 209 260 210
rect 202 203 208 204
rect 202 199 203 203
rect 207 199 208 203
rect 202 198 208 199
rect 256 163 258 209
rect 316 204 318 238
rect 398 214 404 215
rect 398 210 399 214
rect 403 210 404 214
rect 398 209 404 210
rect 550 214 556 215
rect 550 210 551 214
rect 555 210 556 214
rect 550 209 556 210
rect 314 203 320 204
rect 314 199 315 203
rect 319 199 320 203
rect 314 198 320 199
rect 354 203 360 204
rect 354 199 355 203
rect 359 199 360 203
rect 354 198 360 199
rect 111 162 115 163
rect 111 157 115 158
rect 143 162 147 163
rect 143 157 147 158
rect 223 162 227 163
rect 223 157 227 158
rect 255 162 259 163
rect 255 157 259 158
rect 303 162 307 163
rect 303 157 307 158
rect 112 129 114 157
rect 144 147 146 157
rect 194 155 200 156
rect 194 151 195 155
rect 199 151 200 155
rect 194 150 200 151
rect 142 146 148 147
rect 142 142 143 146
rect 147 142 148 146
rect 142 141 148 142
rect 110 128 116 129
rect 110 124 111 128
rect 115 124 116 128
rect 110 123 116 124
rect 196 120 198 150
rect 224 147 226 157
rect 274 155 280 156
rect 274 151 275 155
rect 279 151 280 155
rect 274 150 280 151
rect 222 146 228 147
rect 222 142 223 146
rect 227 142 228 146
rect 222 141 228 142
rect 276 120 278 150
rect 304 147 306 157
rect 302 146 308 147
rect 302 142 303 146
rect 307 142 308 146
rect 302 141 308 142
rect 356 120 358 198
rect 390 163 396 164
rect 400 163 402 209
rect 552 163 554 209
rect 383 162 387 163
rect 390 159 391 163
rect 395 159 396 163
rect 390 158 396 159
rect 399 162 403 163
rect 383 157 387 158
rect 384 147 386 157
rect 382 146 388 147
rect 382 142 383 146
rect 387 142 388 146
rect 382 141 388 142
rect 392 120 394 158
rect 399 157 403 158
rect 463 162 467 163
rect 463 157 467 158
rect 543 162 547 163
rect 543 157 547 158
rect 551 162 555 163
rect 551 157 555 158
rect 442 155 448 156
rect 442 151 443 155
rect 447 151 448 155
rect 442 150 448 151
rect 444 120 446 150
rect 464 147 466 157
rect 522 155 528 156
rect 522 151 523 155
rect 527 151 528 155
rect 522 150 528 151
rect 462 146 468 147
rect 462 142 463 146
rect 467 142 468 146
rect 462 141 468 142
rect 524 120 526 150
rect 544 147 546 157
rect 612 156 614 238
rect 702 214 708 215
rect 702 210 703 214
rect 707 210 708 214
rect 702 209 708 210
rect 704 163 706 209
rect 764 204 766 238
rect 840 204 842 310
rect 902 304 908 305
rect 902 300 903 304
rect 907 300 908 304
rect 902 299 908 300
rect 1014 304 1020 305
rect 1014 300 1015 304
rect 1019 300 1020 304
rect 1014 299 1020 300
rect 1118 304 1124 305
rect 1118 300 1119 304
rect 1123 300 1124 304
rect 1118 299 1124 300
rect 1222 304 1228 305
rect 1222 300 1223 304
rect 1227 300 1228 304
rect 1222 299 1228 300
rect 904 275 906 299
rect 1016 275 1018 299
rect 1120 275 1122 299
rect 1224 275 1226 299
rect 847 274 851 275
rect 847 269 851 270
rect 903 274 907 275
rect 903 269 907 270
rect 991 274 995 275
rect 991 269 995 270
rect 1015 274 1019 275
rect 1015 269 1019 270
rect 1119 274 1123 275
rect 1119 269 1123 270
rect 1223 274 1227 275
rect 1223 269 1227 270
rect 1239 274 1243 275
rect 1239 269 1243 270
rect 848 253 850 269
rect 992 253 994 269
rect 1120 253 1122 269
rect 1240 253 1242 269
rect 846 252 852 253
rect 846 248 847 252
rect 851 248 852 252
rect 846 247 852 248
rect 990 252 996 253
rect 990 248 991 252
rect 995 248 996 252
rect 990 247 996 248
rect 1118 252 1124 253
rect 1118 248 1119 252
rect 1123 248 1124 252
rect 1118 247 1124 248
rect 1238 252 1244 253
rect 1238 248 1239 252
rect 1243 248 1244 252
rect 1238 247 1244 248
rect 1312 244 1314 346
rect 1336 343 1338 353
rect 1386 351 1392 352
rect 1386 347 1387 351
rect 1391 347 1392 351
rect 1386 346 1392 347
rect 1334 342 1340 343
rect 1334 338 1335 342
rect 1339 338 1340 342
rect 1334 337 1340 338
rect 1388 316 1390 346
rect 1440 343 1442 353
rect 1438 342 1444 343
rect 1438 338 1439 342
rect 1443 338 1444 342
rect 1438 337 1444 338
rect 1448 316 1450 354
rect 1831 353 1835 354
rect 1832 325 1834 353
rect 1872 347 1874 379
rect 1982 366 1988 367
rect 1982 362 1983 366
rect 1987 362 1988 366
rect 1982 361 1988 362
rect 1984 347 1986 361
rect 1992 356 1994 430
rect 2184 427 2186 447
rect 2280 427 2282 447
rect 2376 427 2378 447
rect 2480 427 2482 447
rect 2486 435 2492 436
rect 2486 431 2487 435
rect 2491 431 2492 435
rect 2486 430 2492 431
rect 2063 426 2067 427
rect 2063 421 2067 422
rect 2159 426 2163 427
rect 2159 421 2163 422
rect 2183 426 2187 427
rect 2183 421 2187 422
rect 2255 426 2259 427
rect 2255 421 2259 422
rect 2279 426 2283 427
rect 2279 421 2283 422
rect 2359 426 2363 427
rect 2359 421 2363 422
rect 2375 426 2379 427
rect 2375 421 2379 422
rect 2471 426 2475 427
rect 2471 421 2475 422
rect 2479 426 2483 427
rect 2479 421 2483 422
rect 2064 405 2066 421
rect 2160 405 2162 421
rect 2256 405 2258 421
rect 2360 405 2362 421
rect 2472 405 2474 421
rect 2062 404 2068 405
rect 2062 400 2063 404
rect 2067 400 2068 404
rect 2062 399 2068 400
rect 2158 404 2164 405
rect 2158 400 2159 404
rect 2163 400 2164 404
rect 2158 399 2164 400
rect 2254 404 2260 405
rect 2254 400 2255 404
rect 2259 400 2260 404
rect 2254 399 2260 400
rect 2358 404 2364 405
rect 2358 400 2359 404
rect 2363 400 2364 404
rect 2358 399 2364 400
rect 2470 404 2476 405
rect 2470 400 2471 404
rect 2475 400 2476 404
rect 2470 399 2476 400
rect 2042 395 2048 396
rect 2042 391 2043 395
rect 2047 391 2048 395
rect 2042 390 2048 391
rect 2130 395 2136 396
rect 2130 391 2131 395
rect 2135 391 2136 395
rect 2130 390 2136 391
rect 2226 395 2232 396
rect 2226 391 2227 395
rect 2231 391 2232 395
rect 2226 390 2232 391
rect 2044 356 2046 390
rect 2070 366 2076 367
rect 2070 362 2071 366
rect 2075 362 2076 366
rect 2070 361 2076 362
rect 1990 355 1996 356
rect 1990 351 1991 355
rect 1995 351 1996 355
rect 1990 350 1996 351
rect 2042 355 2048 356
rect 2042 351 2043 355
rect 2047 351 2048 355
rect 2042 350 2048 351
rect 2072 347 2074 361
rect 2132 356 2134 390
rect 2166 366 2172 367
rect 2166 362 2167 366
rect 2171 362 2172 366
rect 2166 361 2172 362
rect 2130 355 2136 356
rect 2130 351 2131 355
rect 2135 351 2136 355
rect 2130 350 2136 351
rect 2168 347 2170 361
rect 2228 356 2230 390
rect 2262 366 2268 367
rect 2262 362 2263 366
rect 2267 362 2268 366
rect 2262 361 2268 362
rect 2366 366 2372 367
rect 2366 362 2367 366
rect 2371 362 2372 366
rect 2366 361 2372 362
rect 2478 366 2484 367
rect 2478 362 2479 366
rect 2483 362 2484 366
rect 2478 361 2484 362
rect 2226 355 2232 356
rect 2226 351 2227 355
rect 2231 351 2232 355
rect 2226 350 2232 351
rect 2264 347 2266 361
rect 2368 347 2370 361
rect 2480 347 2482 361
rect 2488 356 2490 430
rect 2576 427 2578 447
rect 2680 427 2682 447
rect 2784 427 2786 447
rect 2904 427 2906 447
rect 3032 427 3034 447
rect 3168 427 3170 447
rect 3312 427 3314 447
rect 2575 426 2579 427
rect 2575 421 2579 422
rect 2607 426 2611 427
rect 2607 421 2611 422
rect 2679 426 2683 427
rect 2679 421 2683 422
rect 2759 426 2763 427
rect 2759 421 2763 422
rect 2783 426 2787 427
rect 2783 421 2787 422
rect 2903 426 2907 427
rect 2903 421 2907 422
rect 2927 426 2931 427
rect 2927 421 2931 422
rect 3031 426 3035 427
rect 3031 421 3035 422
rect 3111 426 3115 427
rect 3111 421 3115 422
rect 3167 426 3171 427
rect 3167 421 3171 422
rect 3303 426 3307 427
rect 3303 421 3307 422
rect 3311 426 3315 427
rect 3311 421 3315 422
rect 2608 405 2610 421
rect 2760 405 2762 421
rect 2928 405 2930 421
rect 3112 405 3114 421
rect 3304 405 3306 421
rect 2606 404 2612 405
rect 2606 400 2607 404
rect 2611 400 2612 404
rect 2606 399 2612 400
rect 2758 404 2764 405
rect 2758 400 2759 404
rect 2763 400 2764 404
rect 2758 399 2764 400
rect 2926 404 2932 405
rect 2926 400 2927 404
rect 2931 400 2932 404
rect 2926 399 2932 400
rect 3110 404 3116 405
rect 3110 400 3111 404
rect 3115 400 3116 404
rect 3110 399 3116 400
rect 3302 404 3308 405
rect 3302 400 3303 404
rect 3307 400 3308 404
rect 3302 399 3308 400
rect 3392 396 3394 494
rect 3472 491 3474 501
rect 3470 490 3476 491
rect 3470 486 3471 490
rect 3475 486 3476 490
rect 3470 485 3476 486
rect 3592 473 3594 501
rect 3590 472 3596 473
rect 3590 468 3591 472
rect 3595 468 3596 472
rect 3590 467 3596 468
rect 3590 455 3596 456
rect 3462 452 3468 453
rect 3462 448 3463 452
rect 3467 448 3468 452
rect 3590 451 3591 455
rect 3595 451 3596 455
rect 3590 450 3596 451
rect 3462 447 3468 448
rect 3464 427 3466 447
rect 3592 427 3594 450
rect 3463 426 3467 427
rect 3463 421 3467 422
rect 3495 426 3499 427
rect 3495 421 3499 422
rect 3591 426 3595 427
rect 3591 421 3595 422
rect 3496 405 3498 421
rect 3494 404 3500 405
rect 3494 400 3495 404
rect 3499 400 3500 404
rect 3592 402 3594 421
rect 3494 399 3500 400
rect 3590 401 3596 402
rect 3590 397 3591 401
rect 3595 397 3596 401
rect 3590 396 3596 397
rect 2538 395 2544 396
rect 2538 391 2539 395
rect 2543 391 2544 395
rect 2538 390 2544 391
rect 2682 395 2688 396
rect 2682 391 2683 395
rect 2687 391 2688 395
rect 2682 390 2688 391
rect 2850 395 2856 396
rect 2850 391 2851 395
rect 2855 391 2856 395
rect 2850 390 2856 391
rect 3026 395 3032 396
rect 3026 391 3027 395
rect 3031 391 3032 395
rect 3026 390 3032 391
rect 3034 395 3040 396
rect 3034 391 3035 395
rect 3039 391 3040 395
rect 3034 390 3040 391
rect 3390 395 3396 396
rect 3390 391 3391 395
rect 3395 391 3396 395
rect 3390 390 3396 391
rect 3494 391 3500 392
rect 2540 356 2542 390
rect 2614 366 2620 367
rect 2614 362 2615 366
rect 2619 362 2620 366
rect 2614 361 2620 362
rect 2486 355 2492 356
rect 2486 351 2487 355
rect 2491 351 2492 355
rect 2486 350 2492 351
rect 2538 355 2544 356
rect 2538 351 2539 355
rect 2543 351 2544 355
rect 2538 350 2544 351
rect 2616 347 2618 361
rect 2684 356 2686 390
rect 2766 366 2772 367
rect 2766 362 2767 366
rect 2771 362 2772 366
rect 2766 361 2772 362
rect 2682 355 2688 356
rect 2682 351 2683 355
rect 2687 351 2688 355
rect 2682 350 2688 351
rect 2768 347 2770 361
rect 2852 356 2854 390
rect 2934 366 2940 367
rect 2934 362 2935 366
rect 2939 362 2940 366
rect 2934 361 2940 362
rect 2850 355 2856 356
rect 2850 351 2851 355
rect 2855 351 2856 355
rect 2850 350 2856 351
rect 2936 347 2938 361
rect 3028 356 3030 390
rect 3026 355 3032 356
rect 3026 351 3027 355
rect 3031 351 3032 355
rect 3026 350 3032 351
rect 1871 346 1875 347
rect 1871 341 1875 342
rect 1983 346 1987 347
rect 1983 341 1987 342
rect 2071 346 2075 347
rect 2071 341 2075 342
rect 2167 346 2171 347
rect 2167 341 2171 342
rect 2215 346 2219 347
rect 2215 341 2219 342
rect 2263 346 2267 347
rect 2263 341 2267 342
rect 2295 346 2299 347
rect 2295 341 2299 342
rect 2367 346 2371 347
rect 2367 341 2371 342
rect 2383 346 2387 347
rect 2383 341 2387 342
rect 2479 346 2483 347
rect 2479 341 2483 342
rect 2591 346 2595 347
rect 2591 341 2595 342
rect 2615 346 2619 347
rect 2615 341 2619 342
rect 2719 346 2723 347
rect 2719 341 2723 342
rect 2767 346 2771 347
rect 2767 341 2771 342
rect 2847 346 2851 347
rect 2847 341 2851 342
rect 2935 346 2939 347
rect 2935 341 2939 342
rect 2983 346 2987 347
rect 2983 341 2987 342
rect 1830 324 1836 325
rect 1830 320 1831 324
rect 1835 320 1836 324
rect 1830 319 1836 320
rect 1386 315 1392 316
rect 1386 311 1387 315
rect 1391 311 1392 315
rect 1386 310 1392 311
rect 1446 315 1452 316
rect 1446 311 1447 315
rect 1451 311 1452 315
rect 1872 313 1874 341
rect 2216 331 2218 341
rect 2274 339 2280 340
rect 2274 335 2275 339
rect 2279 335 2280 339
rect 2274 334 2280 335
rect 2214 330 2220 331
rect 2214 326 2215 330
rect 2219 326 2220 330
rect 2214 325 2220 326
rect 1446 310 1452 311
rect 1870 312 1876 313
rect 1870 308 1871 312
rect 1875 308 1876 312
rect 1830 307 1836 308
rect 1870 307 1876 308
rect 1326 304 1332 305
rect 1326 300 1327 304
rect 1331 300 1332 304
rect 1326 299 1332 300
rect 1430 304 1436 305
rect 1430 300 1431 304
rect 1435 300 1436 304
rect 1830 303 1831 307
rect 1835 303 1836 307
rect 2276 304 2278 334
rect 2296 331 2298 341
rect 2346 339 2352 340
rect 2346 335 2347 339
rect 2351 335 2352 339
rect 2346 334 2352 335
rect 2294 330 2300 331
rect 2294 326 2295 330
rect 2299 326 2300 330
rect 2294 325 2300 326
rect 2348 304 2350 334
rect 2384 331 2386 341
rect 2434 339 2440 340
rect 2434 335 2435 339
rect 2439 335 2440 339
rect 2434 334 2440 335
rect 2382 330 2388 331
rect 2382 326 2383 330
rect 2387 326 2388 330
rect 2382 325 2388 326
rect 2436 304 2438 334
rect 2480 331 2482 341
rect 2530 339 2536 340
rect 2530 335 2531 339
rect 2535 335 2536 339
rect 2530 334 2536 335
rect 2478 330 2484 331
rect 2478 326 2479 330
rect 2483 326 2484 330
rect 2478 325 2484 326
rect 2532 304 2534 334
rect 2592 331 2594 341
rect 2642 339 2648 340
rect 2642 335 2643 339
rect 2647 335 2648 339
rect 2642 334 2648 335
rect 2590 330 2596 331
rect 2590 326 2591 330
rect 2595 326 2596 330
rect 2590 325 2596 326
rect 2644 304 2646 334
rect 2720 331 2722 341
rect 2848 331 2850 341
rect 2906 339 2912 340
rect 2906 335 2907 339
rect 2911 335 2912 339
rect 2906 334 2912 335
rect 2718 330 2724 331
rect 2718 326 2719 330
rect 2723 326 2724 330
rect 2718 325 2724 326
rect 2846 330 2852 331
rect 2846 326 2847 330
rect 2851 326 2852 330
rect 2846 325 2852 326
rect 2908 304 2910 334
rect 2984 331 2986 341
rect 3036 340 3038 390
rect 3494 387 3495 391
rect 3499 387 3500 391
rect 3494 386 3500 387
rect 3118 366 3124 367
rect 3118 362 3119 366
rect 3123 362 3124 366
rect 3118 361 3124 362
rect 3310 366 3316 367
rect 3310 362 3311 366
rect 3315 362 3316 366
rect 3310 361 3316 362
rect 3120 347 3122 361
rect 3312 347 3314 361
rect 3398 355 3404 356
rect 3398 351 3399 355
rect 3403 351 3404 355
rect 3398 350 3404 351
rect 3119 346 3123 347
rect 3119 341 3123 342
rect 3255 346 3259 347
rect 3255 341 3259 342
rect 3311 346 3315 347
rect 3311 341 3315 342
rect 3391 346 3395 347
rect 3391 341 3395 342
rect 3034 339 3040 340
rect 3034 335 3035 339
rect 3039 335 3040 339
rect 3034 334 3040 335
rect 3102 339 3108 340
rect 3102 335 3103 339
rect 3107 335 3108 339
rect 3102 334 3108 335
rect 2982 330 2988 331
rect 2982 326 2983 330
rect 2987 326 2988 330
rect 2982 325 2988 326
rect 1830 302 1836 303
rect 2274 303 2280 304
rect 1430 299 1436 300
rect 1328 275 1330 299
rect 1432 275 1434 299
rect 1832 275 1834 302
rect 2274 299 2275 303
rect 2279 299 2280 303
rect 2274 298 2280 299
rect 2346 303 2352 304
rect 2346 299 2347 303
rect 2351 299 2352 303
rect 2346 298 2352 299
rect 2434 303 2440 304
rect 2434 299 2435 303
rect 2439 299 2440 303
rect 2434 298 2440 299
rect 2530 303 2536 304
rect 2530 299 2531 303
rect 2535 299 2536 303
rect 2530 298 2536 299
rect 2642 303 2648 304
rect 2642 299 2643 303
rect 2647 299 2648 303
rect 2642 298 2648 299
rect 2898 303 2904 304
rect 2898 299 2899 303
rect 2903 299 2904 303
rect 2898 298 2904 299
rect 2906 303 2912 304
rect 2906 299 2907 303
rect 2911 299 2912 303
rect 2906 298 2912 299
rect 1870 295 1876 296
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 1870 290 1876 291
rect 2206 292 2212 293
rect 1327 274 1331 275
rect 1327 269 1331 270
rect 1359 274 1363 275
rect 1359 269 1363 270
rect 1431 274 1435 275
rect 1431 269 1435 270
rect 1479 274 1483 275
rect 1479 269 1483 270
rect 1599 274 1603 275
rect 1599 269 1603 270
rect 1831 274 1835 275
rect 1831 269 1835 270
rect 1360 253 1362 269
rect 1480 253 1482 269
rect 1600 253 1602 269
rect 1358 252 1364 253
rect 1358 248 1359 252
rect 1363 248 1364 252
rect 1358 247 1364 248
rect 1478 252 1484 253
rect 1478 248 1479 252
rect 1483 248 1484 252
rect 1478 247 1484 248
rect 1598 252 1604 253
rect 1598 248 1599 252
rect 1603 248 1604 252
rect 1832 250 1834 269
rect 1872 267 1874 290
rect 2206 288 2207 292
rect 2211 288 2212 292
rect 2206 287 2212 288
rect 2286 292 2292 293
rect 2286 288 2287 292
rect 2291 288 2292 292
rect 2286 287 2292 288
rect 2374 292 2380 293
rect 2374 288 2375 292
rect 2379 288 2380 292
rect 2374 287 2380 288
rect 2470 292 2476 293
rect 2470 288 2471 292
rect 2475 288 2476 292
rect 2470 287 2476 288
rect 2582 292 2588 293
rect 2582 288 2583 292
rect 2587 288 2588 292
rect 2582 287 2588 288
rect 2710 292 2716 293
rect 2710 288 2711 292
rect 2715 288 2716 292
rect 2710 287 2716 288
rect 2838 292 2844 293
rect 2838 288 2839 292
rect 2843 288 2844 292
rect 2838 287 2844 288
rect 2208 267 2210 287
rect 2288 267 2290 287
rect 2376 267 2378 287
rect 2472 267 2474 287
rect 2550 275 2556 276
rect 2550 271 2551 275
rect 2555 271 2556 275
rect 2550 270 2556 271
rect 1871 266 1875 267
rect 1871 261 1875 262
rect 1991 266 1995 267
rect 1991 261 1995 262
rect 2119 266 2123 267
rect 2119 261 2123 262
rect 2207 266 2211 267
rect 2207 261 2211 262
rect 2255 266 2259 267
rect 2255 261 2259 262
rect 2287 266 2291 267
rect 2287 261 2291 262
rect 2375 266 2379 267
rect 2375 261 2379 262
rect 2391 266 2395 267
rect 2391 261 2395 262
rect 2471 266 2475 267
rect 2471 261 2475 262
rect 2535 266 2539 267
rect 2535 261 2539 262
rect 1598 247 1604 248
rect 1830 249 1836 250
rect 1830 245 1831 249
rect 1835 245 1836 249
rect 1830 244 1836 245
rect 1062 243 1068 244
rect 1062 239 1063 243
rect 1067 239 1068 243
rect 1062 238 1068 239
rect 1186 243 1192 244
rect 1186 239 1187 243
rect 1191 239 1192 243
rect 1186 238 1192 239
rect 1310 243 1316 244
rect 1310 239 1311 243
rect 1315 239 1316 243
rect 1310 238 1316 239
rect 1426 243 1432 244
rect 1426 239 1427 243
rect 1431 239 1432 243
rect 1426 238 1432 239
rect 1546 243 1552 244
rect 1546 239 1547 243
rect 1551 239 1552 243
rect 1872 242 1874 261
rect 1992 245 1994 261
rect 2120 245 2122 261
rect 2256 245 2258 261
rect 2392 245 2394 261
rect 2536 245 2538 261
rect 1990 244 1996 245
rect 1546 238 1552 239
rect 1870 241 1876 242
rect 1050 235 1056 236
rect 1050 231 1051 235
rect 1055 231 1056 235
rect 1050 230 1056 231
rect 854 214 860 215
rect 854 210 855 214
rect 859 210 860 214
rect 854 209 860 210
rect 998 214 1004 215
rect 998 210 999 214
rect 1003 210 1004 214
rect 998 209 1004 210
rect 762 203 768 204
rect 762 199 763 203
rect 767 199 768 203
rect 762 198 768 199
rect 838 203 844 204
rect 838 199 839 203
rect 843 199 844 203
rect 838 198 844 199
rect 790 163 796 164
rect 856 163 858 209
rect 1000 163 1002 209
rect 1052 204 1054 230
rect 1064 204 1066 238
rect 1126 214 1132 215
rect 1126 210 1127 214
rect 1131 210 1132 214
rect 1126 209 1132 210
rect 1050 203 1056 204
rect 1050 199 1051 203
rect 1055 199 1056 203
rect 1050 198 1056 199
rect 1062 203 1068 204
rect 1062 199 1063 203
rect 1067 199 1068 203
rect 1062 198 1068 199
rect 1075 172 1079 173
rect 1075 167 1079 168
rect 623 162 627 163
rect 623 157 627 158
rect 703 162 707 163
rect 703 157 707 158
rect 783 162 787 163
rect 790 159 791 163
rect 795 159 796 163
rect 790 158 796 159
rect 855 162 859 163
rect 783 157 787 158
rect 610 155 616 156
rect 610 151 611 155
rect 615 151 616 155
rect 610 150 616 151
rect 624 147 626 157
rect 674 155 680 156
rect 674 151 675 155
rect 679 151 680 155
rect 674 150 680 151
rect 542 146 548 147
rect 542 142 543 146
rect 547 142 548 146
rect 542 141 548 142
rect 622 146 628 147
rect 622 142 623 146
rect 627 142 628 146
rect 622 141 628 142
rect 676 120 678 150
rect 704 147 706 157
rect 754 155 760 156
rect 754 151 755 155
rect 759 151 760 155
rect 754 150 760 151
rect 702 146 708 147
rect 702 142 703 146
rect 707 142 708 146
rect 702 141 708 142
rect 756 120 758 150
rect 784 147 786 157
rect 782 146 788 147
rect 782 142 783 146
rect 787 142 788 146
rect 782 141 788 142
rect 792 120 794 158
rect 855 157 859 158
rect 863 162 867 163
rect 863 157 867 158
rect 943 162 947 163
rect 943 157 947 158
rect 999 162 1003 163
rect 999 157 1003 158
rect 1023 162 1027 163
rect 1023 157 1027 158
rect 864 147 866 157
rect 914 155 920 156
rect 914 151 915 155
rect 919 151 920 155
rect 914 150 920 151
rect 862 146 868 147
rect 862 142 863 146
rect 867 142 868 146
rect 862 141 868 142
rect 916 120 918 150
rect 944 147 946 157
rect 1006 155 1012 156
rect 1006 151 1007 155
rect 1011 151 1012 155
rect 1006 150 1012 151
rect 942 146 948 147
rect 942 142 943 146
rect 947 142 948 146
rect 942 141 948 142
rect 1008 120 1010 150
rect 1024 147 1026 157
rect 1022 146 1028 147
rect 1022 142 1023 146
rect 1027 142 1028 146
rect 1022 141 1028 142
rect 1076 120 1078 167
rect 1110 163 1116 164
rect 1128 163 1130 209
rect 1188 204 1190 238
rect 1246 214 1252 215
rect 1246 210 1247 214
rect 1251 210 1252 214
rect 1246 209 1252 210
rect 1366 214 1372 215
rect 1366 210 1367 214
rect 1371 210 1372 214
rect 1366 209 1372 210
rect 1186 203 1192 204
rect 1186 199 1187 203
rect 1191 199 1192 203
rect 1186 198 1192 199
rect 1248 163 1250 209
rect 1358 203 1364 204
rect 1358 199 1359 203
rect 1363 199 1364 203
rect 1358 198 1364 199
rect 1360 173 1362 198
rect 1359 172 1363 173
rect 1359 167 1363 168
rect 1368 163 1370 209
rect 1428 204 1430 238
rect 1486 214 1492 215
rect 1486 210 1487 214
rect 1491 210 1492 214
rect 1486 209 1492 210
rect 1426 203 1432 204
rect 1426 199 1427 203
rect 1431 199 1432 203
rect 1426 198 1432 199
rect 1488 163 1490 209
rect 1548 204 1550 238
rect 1870 237 1871 241
rect 1875 237 1876 241
rect 1990 240 1991 244
rect 1995 240 1996 244
rect 1990 239 1996 240
rect 2118 244 2124 245
rect 2118 240 2119 244
rect 2123 240 2124 244
rect 2118 239 2124 240
rect 2254 244 2260 245
rect 2254 240 2255 244
rect 2259 240 2260 244
rect 2254 239 2260 240
rect 2390 244 2396 245
rect 2390 240 2391 244
rect 2395 240 2396 244
rect 2390 239 2396 240
rect 2534 244 2540 245
rect 2534 240 2535 244
rect 2539 240 2540 244
rect 2534 239 2540 240
rect 1870 236 1876 237
rect 2062 235 2068 236
rect 1830 232 1836 233
rect 1830 228 1831 232
rect 1835 228 1836 232
rect 2062 231 2063 235
rect 2067 231 2068 235
rect 2062 230 2068 231
rect 2186 235 2192 236
rect 2186 231 2187 235
rect 2191 231 2192 235
rect 2186 230 2192 231
rect 2334 235 2340 236
rect 2334 231 2335 235
rect 2339 231 2340 235
rect 2334 230 2340 231
rect 2458 235 2464 236
rect 2458 231 2459 235
rect 2463 231 2464 235
rect 2458 230 2464 231
rect 1830 227 1836 228
rect 2050 227 2056 228
rect 1606 214 1612 215
rect 1606 210 1607 214
rect 1611 210 1612 214
rect 1606 209 1612 210
rect 1546 203 1552 204
rect 1546 199 1547 203
rect 1551 199 1552 203
rect 1546 198 1552 199
rect 1608 163 1610 209
rect 1832 163 1834 227
rect 1870 224 1876 225
rect 1870 220 1871 224
rect 1875 220 1876 224
rect 2050 223 2051 227
rect 2055 223 2056 227
rect 2050 222 2056 223
rect 1870 219 1876 220
rect 1872 179 1874 219
rect 1998 206 2004 207
rect 1998 202 1999 206
rect 2003 202 2004 206
rect 1998 201 2004 202
rect 2000 179 2002 201
rect 2052 196 2054 222
rect 2064 196 2066 230
rect 2126 206 2132 207
rect 2126 202 2127 206
rect 2131 202 2132 206
rect 2126 201 2132 202
rect 2050 195 2056 196
rect 2050 191 2051 195
rect 2055 191 2056 195
rect 2050 190 2056 191
rect 2062 195 2068 196
rect 2062 191 2063 195
rect 2067 191 2068 195
rect 2062 190 2068 191
rect 2128 179 2130 201
rect 1871 178 1875 179
rect 1871 173 1875 174
rect 1903 178 1907 179
rect 1903 173 1907 174
rect 1983 178 1987 179
rect 1983 173 1987 174
rect 1999 178 2003 179
rect 1999 173 2003 174
rect 2087 178 2091 179
rect 2087 173 2091 174
rect 2127 178 2131 179
rect 2127 173 2131 174
rect 1103 162 1107 163
rect 1110 159 1111 163
rect 1115 159 1116 163
rect 1110 158 1116 159
rect 1127 162 1131 163
rect 1103 157 1107 158
rect 1104 147 1106 157
rect 1102 146 1108 147
rect 1102 142 1103 146
rect 1107 142 1108 146
rect 1102 141 1108 142
rect 1112 120 1114 158
rect 1127 157 1131 158
rect 1183 162 1187 163
rect 1183 157 1187 158
rect 1247 162 1251 163
rect 1247 157 1251 158
rect 1263 162 1267 163
rect 1263 157 1267 158
rect 1343 162 1347 163
rect 1343 157 1347 158
rect 1367 162 1371 163
rect 1367 157 1371 158
rect 1423 162 1427 163
rect 1423 157 1427 158
rect 1487 162 1491 163
rect 1487 157 1491 158
rect 1511 162 1515 163
rect 1511 157 1515 158
rect 1591 162 1595 163
rect 1591 157 1595 158
rect 1607 162 1611 163
rect 1607 157 1611 158
rect 1671 162 1675 163
rect 1671 157 1675 158
rect 1751 162 1755 163
rect 1751 157 1755 158
rect 1831 162 1835 163
rect 1831 157 1835 158
rect 1162 155 1168 156
rect 1162 151 1163 155
rect 1167 151 1168 155
rect 1162 150 1168 151
rect 1164 120 1166 150
rect 1184 147 1186 157
rect 1264 147 1266 157
rect 1322 155 1328 156
rect 1322 151 1323 155
rect 1327 151 1328 155
rect 1322 150 1328 151
rect 1182 146 1188 147
rect 1182 142 1183 146
rect 1187 142 1188 146
rect 1182 141 1188 142
rect 1262 146 1268 147
rect 1262 142 1263 146
rect 1267 142 1268 146
rect 1262 141 1268 142
rect 1324 120 1326 150
rect 1344 147 1346 157
rect 1402 155 1408 156
rect 1402 151 1403 155
rect 1407 151 1408 155
rect 1402 150 1408 151
rect 1342 146 1348 147
rect 1342 142 1343 146
rect 1347 142 1348 146
rect 1342 141 1348 142
rect 1404 120 1406 150
rect 1424 147 1426 157
rect 1512 147 1514 157
rect 1570 155 1576 156
rect 1570 151 1571 155
rect 1575 151 1576 155
rect 1570 150 1576 151
rect 1422 146 1428 147
rect 1422 142 1423 146
rect 1427 142 1428 146
rect 1422 141 1428 142
rect 1510 146 1516 147
rect 1510 142 1511 146
rect 1515 142 1516 146
rect 1510 141 1516 142
rect 1572 120 1574 150
rect 1592 147 1594 157
rect 1650 155 1656 156
rect 1650 151 1651 155
rect 1655 151 1656 155
rect 1650 150 1656 151
rect 1590 146 1596 147
rect 1590 142 1591 146
rect 1595 142 1596 146
rect 1590 141 1596 142
rect 1652 120 1654 150
rect 1672 147 1674 157
rect 1730 155 1736 156
rect 1730 151 1731 155
rect 1735 151 1736 155
rect 1730 150 1736 151
rect 1670 146 1676 147
rect 1670 142 1671 146
rect 1675 142 1676 146
rect 1670 141 1676 142
rect 1732 120 1734 150
rect 1752 147 1754 157
rect 1802 155 1808 156
rect 1802 151 1803 155
rect 1807 151 1808 155
rect 1802 150 1808 151
rect 1750 146 1756 147
rect 1750 142 1751 146
rect 1755 142 1756 146
rect 1750 141 1756 142
rect 1804 136 1806 150
rect 1802 135 1808 136
rect 1802 131 1803 135
rect 1807 131 1808 135
rect 1802 130 1808 131
rect 1832 129 1834 157
rect 1872 145 1874 173
rect 1904 163 1906 173
rect 1962 171 1968 172
rect 1962 167 1963 171
rect 1967 167 1968 171
rect 1962 166 1968 167
rect 1902 162 1908 163
rect 1902 158 1903 162
rect 1907 158 1908 162
rect 1902 157 1908 158
rect 1870 144 1876 145
rect 1870 140 1871 144
rect 1875 140 1876 144
rect 1870 139 1876 140
rect 1964 136 1966 166
rect 1984 163 1986 173
rect 2042 171 2048 172
rect 2042 167 2043 171
rect 2047 167 2048 171
rect 2042 166 2048 167
rect 1982 162 1988 163
rect 1982 158 1983 162
rect 1987 158 1988 162
rect 1982 157 1988 158
rect 2044 136 2046 166
rect 2088 163 2090 173
rect 2188 172 2190 230
rect 2262 206 2268 207
rect 2262 202 2263 206
rect 2267 202 2268 206
rect 2262 201 2268 202
rect 2264 179 2266 201
rect 2336 196 2338 230
rect 2398 206 2404 207
rect 2398 202 2399 206
rect 2403 202 2404 206
rect 2398 201 2404 202
rect 2334 195 2340 196
rect 2334 191 2335 195
rect 2339 191 2340 195
rect 2334 190 2340 191
rect 2400 179 2402 201
rect 2460 196 2462 230
rect 2542 206 2548 207
rect 2542 202 2543 206
rect 2547 202 2548 206
rect 2542 201 2548 202
rect 2458 195 2464 196
rect 2458 191 2459 195
rect 2463 191 2464 195
rect 2458 190 2464 191
rect 2494 179 2500 180
rect 2544 179 2546 201
rect 2552 196 2554 270
rect 2584 267 2586 287
rect 2712 267 2714 287
rect 2840 267 2842 287
rect 2583 266 2587 267
rect 2583 261 2587 262
rect 2679 266 2683 267
rect 2679 261 2683 262
rect 2711 266 2715 267
rect 2711 261 2715 262
rect 2815 266 2819 267
rect 2815 261 2819 262
rect 2839 266 2843 267
rect 2839 261 2843 262
rect 2680 245 2682 261
rect 2816 245 2818 261
rect 2678 244 2684 245
rect 2678 240 2679 244
rect 2683 240 2684 244
rect 2678 239 2684 240
rect 2814 244 2820 245
rect 2814 240 2815 244
rect 2819 240 2820 244
rect 2814 239 2820 240
rect 2746 235 2752 236
rect 2746 231 2747 235
rect 2751 231 2752 235
rect 2746 230 2752 231
rect 2882 235 2888 236
rect 2882 231 2883 235
rect 2887 231 2888 235
rect 2882 230 2888 231
rect 2686 206 2692 207
rect 2686 202 2687 206
rect 2691 202 2692 206
rect 2686 201 2692 202
rect 2550 195 2556 196
rect 2550 191 2551 195
rect 2555 191 2556 195
rect 2550 190 2556 191
rect 2688 179 2690 201
rect 2748 196 2750 230
rect 2822 206 2828 207
rect 2822 202 2823 206
rect 2827 202 2828 206
rect 2822 201 2828 202
rect 2746 195 2752 196
rect 2746 191 2747 195
rect 2751 191 2752 195
rect 2746 190 2752 191
rect 2824 179 2826 201
rect 2884 196 2886 230
rect 2900 196 2902 298
rect 2974 292 2980 293
rect 2974 288 2975 292
rect 2979 288 2980 292
rect 2974 287 2980 288
rect 2976 267 2978 287
rect 2951 266 2955 267
rect 2951 261 2955 262
rect 2975 266 2979 267
rect 2975 261 2979 262
rect 3095 266 3099 267
rect 3095 261 3099 262
rect 2952 245 2954 261
rect 3096 245 3098 261
rect 2950 244 2956 245
rect 2950 240 2951 244
rect 2955 240 2956 244
rect 2950 239 2956 240
rect 3094 244 3100 245
rect 3094 240 3095 244
rect 3099 240 3100 244
rect 3094 239 3100 240
rect 3104 232 3106 334
rect 3120 331 3122 341
rect 3170 339 3176 340
rect 3170 335 3171 339
rect 3175 335 3176 339
rect 3170 334 3176 335
rect 3118 330 3124 331
rect 3118 326 3119 330
rect 3123 326 3124 330
rect 3118 325 3124 326
rect 3172 304 3174 334
rect 3256 331 3258 341
rect 3370 339 3376 340
rect 3370 335 3371 339
rect 3375 335 3376 339
rect 3370 334 3376 335
rect 3254 330 3260 331
rect 3254 326 3255 330
rect 3259 326 3260 330
rect 3254 325 3260 326
rect 3372 304 3374 334
rect 3392 331 3394 341
rect 3390 330 3396 331
rect 3390 326 3391 330
rect 3395 326 3396 330
rect 3390 325 3396 326
rect 3400 304 3402 350
rect 3496 340 3498 386
rect 3590 384 3596 385
rect 3590 380 3591 384
rect 3595 380 3596 384
rect 3590 379 3596 380
rect 3502 366 3508 367
rect 3502 362 3503 366
rect 3507 362 3508 366
rect 3502 361 3508 362
rect 3504 347 3506 361
rect 3592 347 3594 379
rect 3503 346 3507 347
rect 3503 341 3507 342
rect 3511 346 3515 347
rect 3511 341 3515 342
rect 3591 346 3595 347
rect 3591 341 3595 342
rect 3494 339 3500 340
rect 3494 335 3495 339
rect 3499 335 3500 339
rect 3494 334 3500 335
rect 3512 331 3514 341
rect 3510 330 3516 331
rect 3510 326 3511 330
rect 3515 326 3516 330
rect 3510 325 3516 326
rect 3592 313 3594 341
rect 3590 312 3596 313
rect 3590 308 3591 312
rect 3595 308 3596 312
rect 3590 307 3596 308
rect 3170 303 3176 304
rect 3170 299 3171 303
rect 3175 299 3176 303
rect 3170 298 3176 299
rect 3370 303 3376 304
rect 3370 299 3371 303
rect 3375 299 3376 303
rect 3370 298 3376 299
rect 3398 303 3404 304
rect 3398 299 3399 303
rect 3403 299 3404 303
rect 3398 298 3404 299
rect 3590 295 3596 296
rect 3110 292 3116 293
rect 3110 288 3111 292
rect 3115 288 3116 292
rect 3110 287 3116 288
rect 3246 292 3252 293
rect 3246 288 3247 292
rect 3251 288 3252 292
rect 3246 287 3252 288
rect 3382 292 3388 293
rect 3382 288 3383 292
rect 3387 288 3388 292
rect 3382 287 3388 288
rect 3502 292 3508 293
rect 3502 288 3503 292
rect 3507 288 3508 292
rect 3590 291 3591 295
rect 3595 291 3596 295
rect 3590 290 3596 291
rect 3502 287 3508 288
rect 3112 267 3114 287
rect 3248 267 3250 287
rect 3384 267 3386 287
rect 3504 267 3506 287
rect 3518 275 3524 276
rect 3518 271 3519 275
rect 3523 271 3524 275
rect 3518 270 3524 271
rect 3111 266 3115 267
rect 3111 261 3115 262
rect 3239 266 3243 267
rect 3239 261 3243 262
rect 3247 266 3251 267
rect 3247 261 3251 262
rect 3383 266 3387 267
rect 3383 261 3387 262
rect 3503 266 3507 267
rect 3503 261 3507 262
rect 3240 245 3242 261
rect 3384 245 3386 261
rect 3504 245 3506 261
rect 3238 244 3244 245
rect 3238 240 3239 244
rect 3243 240 3244 244
rect 3238 239 3244 240
rect 3382 244 3388 245
rect 3382 240 3383 244
rect 3387 240 3388 244
rect 3382 239 3388 240
rect 3502 244 3508 245
rect 3502 240 3503 244
rect 3507 240 3508 244
rect 3502 239 3508 240
rect 3194 235 3200 236
rect 3102 231 3108 232
rect 3102 227 3103 231
rect 3107 227 3108 231
rect 3194 231 3195 235
rect 3199 231 3200 235
rect 3194 230 3200 231
rect 3306 235 3312 236
rect 3306 231 3307 235
rect 3311 231 3312 235
rect 3306 230 3312 231
rect 3502 231 3508 232
rect 3102 226 3108 227
rect 2958 206 2964 207
rect 2958 202 2959 206
rect 2963 202 2964 206
rect 2958 201 2964 202
rect 3102 206 3108 207
rect 3102 202 3103 206
rect 3107 202 3108 206
rect 3102 201 3108 202
rect 2882 195 2888 196
rect 2882 191 2883 195
rect 2887 191 2888 195
rect 2882 190 2888 191
rect 2898 195 2904 196
rect 2898 191 2899 195
rect 2903 191 2904 195
rect 2898 190 2904 191
rect 2960 179 2962 201
rect 3104 179 3106 201
rect 3196 196 3198 230
rect 3246 206 3252 207
rect 3246 202 3247 206
rect 3251 202 3252 206
rect 3246 201 3252 202
rect 3194 195 3200 196
rect 3194 191 3195 195
rect 3199 191 3200 195
rect 3194 190 3200 191
rect 3248 179 3250 201
rect 3308 196 3310 230
rect 3502 227 3503 231
rect 3507 227 3508 231
rect 3502 226 3508 227
rect 3390 206 3396 207
rect 3390 202 3391 206
rect 3395 202 3396 206
rect 3390 201 3396 202
rect 3306 195 3312 196
rect 3306 191 3307 195
rect 3311 191 3312 195
rect 3306 190 3312 191
rect 3382 195 3388 196
rect 3382 191 3383 195
rect 3387 191 3388 195
rect 3382 190 3388 191
rect 2215 178 2219 179
rect 2215 173 2219 174
rect 2263 178 2267 179
rect 2263 173 2267 174
rect 2351 178 2355 179
rect 2351 173 2355 174
rect 2399 178 2403 179
rect 2399 173 2403 174
rect 2487 178 2491 179
rect 2494 175 2495 179
rect 2499 175 2500 179
rect 2494 174 2500 175
rect 2543 178 2547 179
rect 2487 173 2491 174
rect 2186 171 2192 172
rect 2186 167 2187 171
rect 2191 167 2192 171
rect 2186 166 2192 167
rect 2216 163 2218 173
rect 2318 171 2324 172
rect 2318 167 2319 171
rect 2323 167 2324 171
rect 2318 166 2324 167
rect 2086 162 2092 163
rect 2086 158 2087 162
rect 2091 158 2092 162
rect 2086 157 2092 158
rect 2214 162 2220 163
rect 2214 158 2215 162
rect 2219 158 2220 162
rect 2214 157 2220 158
rect 2320 136 2322 166
rect 2352 163 2354 173
rect 2478 171 2484 172
rect 2478 167 2479 171
rect 2483 167 2484 171
rect 2478 166 2484 167
rect 2350 162 2356 163
rect 2350 158 2351 162
rect 2355 158 2356 162
rect 2350 157 2356 158
rect 2480 136 2482 166
rect 2488 163 2490 173
rect 2486 162 2492 163
rect 2486 158 2487 162
rect 2491 158 2492 162
rect 2486 157 2492 158
rect 2496 136 2498 174
rect 2543 173 2547 174
rect 2623 178 2627 179
rect 2623 173 2627 174
rect 2687 178 2691 179
rect 2687 173 2691 174
rect 2743 178 2747 179
rect 2743 173 2747 174
rect 2823 178 2827 179
rect 2823 173 2827 174
rect 2855 178 2859 179
rect 2855 173 2859 174
rect 2959 178 2963 179
rect 2959 173 2963 174
rect 3063 178 3067 179
rect 3063 173 3067 174
rect 3103 178 3107 179
rect 3103 173 3107 174
rect 3159 178 3163 179
rect 3159 173 3163 174
rect 3247 178 3251 179
rect 3247 173 3251 174
rect 3343 178 3347 179
rect 3343 173 3347 174
rect 2624 163 2626 173
rect 2674 171 2680 172
rect 2674 167 2675 171
rect 2679 167 2680 171
rect 2674 166 2680 167
rect 2622 162 2628 163
rect 2622 158 2623 162
rect 2627 158 2628 162
rect 2622 157 2628 158
rect 2676 136 2678 166
rect 2744 163 2746 173
rect 2794 171 2800 172
rect 2794 167 2795 171
rect 2799 167 2800 171
rect 2794 166 2800 167
rect 2742 162 2748 163
rect 2742 158 2743 162
rect 2747 158 2748 162
rect 2742 157 2748 158
rect 2796 136 2798 166
rect 2856 163 2858 173
rect 2906 171 2912 172
rect 2906 167 2907 171
rect 2911 167 2912 171
rect 2906 166 2912 167
rect 2854 162 2860 163
rect 2854 158 2855 162
rect 2859 158 2860 162
rect 2854 157 2860 158
rect 2908 136 2910 166
rect 2960 163 2962 173
rect 3010 171 3016 172
rect 3010 167 3011 171
rect 3015 167 3016 171
rect 3010 166 3016 167
rect 2958 162 2964 163
rect 2958 158 2959 162
rect 2963 158 2964 162
rect 2958 157 2964 158
rect 3012 136 3014 166
rect 3064 163 3066 173
rect 3114 171 3120 172
rect 3114 167 3115 171
rect 3119 167 3120 171
rect 3114 166 3120 167
rect 3062 162 3068 163
rect 3062 158 3063 162
rect 3067 158 3068 162
rect 3062 157 3068 158
rect 3116 136 3118 166
rect 3160 163 3162 173
rect 3210 171 3216 172
rect 3210 167 3211 171
rect 3215 167 3216 171
rect 3210 166 3216 167
rect 3158 162 3164 163
rect 3158 158 3159 162
rect 3163 158 3164 162
rect 3158 157 3164 158
rect 3212 136 3214 166
rect 3248 163 3250 173
rect 3298 171 3304 172
rect 3298 167 3299 171
rect 3303 167 3304 171
rect 3298 166 3304 167
rect 3246 162 3252 163
rect 3246 158 3247 162
rect 3251 158 3252 162
rect 3246 157 3252 158
rect 3300 136 3302 166
rect 3344 163 3346 173
rect 3342 162 3348 163
rect 3342 158 3343 162
rect 3347 158 3348 162
rect 3342 157 3348 158
rect 3384 136 3386 190
rect 3392 179 3394 201
rect 3391 178 3395 179
rect 3391 173 3395 174
rect 3431 178 3435 179
rect 3431 173 3435 174
rect 3432 163 3434 173
rect 3504 172 3506 226
rect 3510 206 3516 207
rect 3510 202 3511 206
rect 3515 202 3516 206
rect 3510 201 3516 202
rect 3512 179 3514 201
rect 3520 196 3522 270
rect 3592 267 3594 290
rect 3591 266 3595 267
rect 3591 261 3595 262
rect 3592 242 3594 261
rect 3590 241 3596 242
rect 3590 237 3591 241
rect 3595 237 3596 241
rect 3590 236 3596 237
rect 3590 224 3596 225
rect 3590 220 3591 224
rect 3595 220 3596 224
rect 3590 219 3596 220
rect 3518 195 3524 196
rect 3518 191 3519 195
rect 3523 191 3524 195
rect 3518 190 3524 191
rect 3592 179 3594 219
rect 3511 178 3515 179
rect 3511 173 3515 174
rect 3591 178 3595 179
rect 3591 173 3595 174
rect 3490 171 3496 172
rect 3490 167 3491 171
rect 3495 167 3496 171
rect 3490 166 3496 167
rect 3502 171 3508 172
rect 3502 167 3503 171
rect 3507 167 3508 171
rect 3502 166 3508 167
rect 3430 162 3436 163
rect 3430 158 3431 162
rect 3435 158 3436 162
rect 3430 157 3436 158
rect 3492 136 3494 166
rect 3512 163 3514 173
rect 3510 162 3516 163
rect 3510 158 3511 162
rect 3515 158 3516 162
rect 3510 157 3516 158
rect 3592 145 3594 173
rect 3590 144 3596 145
rect 3590 140 3591 144
rect 3595 140 3596 144
rect 3590 139 3596 140
rect 1962 135 1968 136
rect 1962 131 1963 135
rect 1967 131 1968 135
rect 1962 130 1968 131
rect 2042 135 2048 136
rect 2042 131 2043 135
rect 2047 131 2048 135
rect 2042 130 2048 131
rect 2318 135 2324 136
rect 2318 131 2319 135
rect 2323 131 2324 135
rect 2318 130 2324 131
rect 2478 135 2484 136
rect 2478 131 2479 135
rect 2483 131 2484 135
rect 2478 130 2484 131
rect 2494 135 2500 136
rect 2494 131 2495 135
rect 2499 131 2500 135
rect 2494 130 2500 131
rect 2674 135 2680 136
rect 2674 131 2675 135
rect 2679 131 2680 135
rect 2674 130 2680 131
rect 2794 135 2800 136
rect 2794 131 2795 135
rect 2799 131 2800 135
rect 2794 130 2800 131
rect 2906 135 2912 136
rect 2906 131 2907 135
rect 2911 131 2912 135
rect 2906 130 2912 131
rect 3010 135 3016 136
rect 3010 131 3011 135
rect 3015 131 3016 135
rect 3010 130 3016 131
rect 3114 135 3120 136
rect 3114 131 3115 135
rect 3119 131 3120 135
rect 3114 130 3120 131
rect 3210 135 3216 136
rect 3210 131 3211 135
rect 3215 131 3216 135
rect 3210 130 3216 131
rect 3298 135 3304 136
rect 3298 131 3299 135
rect 3303 131 3304 135
rect 3298 130 3304 131
rect 3382 135 3388 136
rect 3382 131 3383 135
rect 3387 131 3388 135
rect 3382 130 3388 131
rect 3490 135 3496 136
rect 3490 131 3491 135
rect 3495 131 3496 135
rect 3490 130 3496 131
rect 1830 128 1836 129
rect 1830 124 1831 128
rect 1835 124 1836 128
rect 1830 123 1836 124
rect 1870 127 1876 128
rect 1870 123 1871 127
rect 1875 123 1876 127
rect 3590 127 3596 128
rect 1870 122 1876 123
rect 1894 124 1900 125
rect 194 119 200 120
rect 194 115 195 119
rect 199 115 200 119
rect 194 114 200 115
rect 274 119 280 120
rect 274 115 275 119
rect 279 115 280 119
rect 274 114 280 115
rect 354 119 360 120
rect 354 115 355 119
rect 359 115 360 119
rect 354 114 360 115
rect 390 119 396 120
rect 390 115 391 119
rect 395 115 396 119
rect 390 114 396 115
rect 442 119 448 120
rect 442 115 443 119
rect 447 115 448 119
rect 442 114 448 115
rect 522 119 528 120
rect 522 115 523 119
rect 527 115 528 119
rect 522 114 528 115
rect 674 119 680 120
rect 674 115 675 119
rect 679 115 680 119
rect 674 114 680 115
rect 754 119 760 120
rect 754 115 755 119
rect 759 115 760 119
rect 754 114 760 115
rect 790 119 796 120
rect 790 115 791 119
rect 795 115 796 119
rect 790 114 796 115
rect 914 119 920 120
rect 914 115 915 119
rect 919 115 920 119
rect 914 114 920 115
rect 1006 119 1012 120
rect 1006 115 1007 119
rect 1011 115 1012 119
rect 1006 114 1012 115
rect 1074 119 1080 120
rect 1074 115 1075 119
rect 1079 115 1080 119
rect 1074 114 1080 115
rect 1110 119 1116 120
rect 1110 115 1111 119
rect 1115 115 1116 119
rect 1110 114 1116 115
rect 1162 119 1168 120
rect 1162 115 1163 119
rect 1167 115 1168 119
rect 1162 114 1168 115
rect 1322 119 1328 120
rect 1322 115 1323 119
rect 1327 115 1328 119
rect 1322 114 1328 115
rect 1402 119 1408 120
rect 1402 115 1403 119
rect 1407 115 1408 119
rect 1402 114 1408 115
rect 1570 119 1576 120
rect 1570 115 1571 119
rect 1575 115 1576 119
rect 1570 114 1576 115
rect 1650 119 1656 120
rect 1650 115 1651 119
rect 1655 115 1656 119
rect 1650 114 1656 115
rect 1730 119 1736 120
rect 1730 115 1731 119
rect 1735 115 1736 119
rect 1730 114 1736 115
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 1830 111 1836 112
rect 110 106 116 107
rect 134 108 140 109
rect 112 87 114 106
rect 134 104 135 108
rect 139 104 140 108
rect 134 103 140 104
rect 214 108 220 109
rect 214 104 215 108
rect 219 104 220 108
rect 214 103 220 104
rect 294 108 300 109
rect 294 104 295 108
rect 299 104 300 108
rect 294 103 300 104
rect 374 108 380 109
rect 374 104 375 108
rect 379 104 380 108
rect 374 103 380 104
rect 454 108 460 109
rect 454 104 455 108
rect 459 104 460 108
rect 454 103 460 104
rect 534 108 540 109
rect 534 104 535 108
rect 539 104 540 108
rect 534 103 540 104
rect 614 108 620 109
rect 614 104 615 108
rect 619 104 620 108
rect 614 103 620 104
rect 694 108 700 109
rect 694 104 695 108
rect 699 104 700 108
rect 694 103 700 104
rect 774 108 780 109
rect 774 104 775 108
rect 779 104 780 108
rect 774 103 780 104
rect 854 108 860 109
rect 854 104 855 108
rect 859 104 860 108
rect 854 103 860 104
rect 934 108 940 109
rect 934 104 935 108
rect 939 104 940 108
rect 934 103 940 104
rect 1014 108 1020 109
rect 1014 104 1015 108
rect 1019 104 1020 108
rect 1014 103 1020 104
rect 1094 108 1100 109
rect 1094 104 1095 108
rect 1099 104 1100 108
rect 1094 103 1100 104
rect 1174 108 1180 109
rect 1174 104 1175 108
rect 1179 104 1180 108
rect 1174 103 1180 104
rect 1254 108 1260 109
rect 1254 104 1255 108
rect 1259 104 1260 108
rect 1254 103 1260 104
rect 1334 108 1340 109
rect 1334 104 1335 108
rect 1339 104 1340 108
rect 1334 103 1340 104
rect 1414 108 1420 109
rect 1414 104 1415 108
rect 1419 104 1420 108
rect 1414 103 1420 104
rect 1502 108 1508 109
rect 1502 104 1503 108
rect 1507 104 1508 108
rect 1502 103 1508 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1662 108 1668 109
rect 1662 104 1663 108
rect 1667 104 1668 108
rect 1662 103 1668 104
rect 1742 108 1748 109
rect 1742 104 1743 108
rect 1747 104 1748 108
rect 1830 107 1831 111
rect 1835 107 1836 111
rect 1830 106 1836 107
rect 1742 103 1748 104
rect 136 87 138 103
rect 216 87 218 103
rect 296 87 298 103
rect 376 87 378 103
rect 456 87 458 103
rect 536 87 538 103
rect 616 87 618 103
rect 696 87 698 103
rect 776 87 778 103
rect 856 87 858 103
rect 936 87 938 103
rect 1016 87 1018 103
rect 1096 87 1098 103
rect 1176 87 1178 103
rect 1256 87 1258 103
rect 1336 87 1338 103
rect 1416 87 1418 103
rect 1504 87 1506 103
rect 1584 87 1586 103
rect 1664 87 1666 103
rect 1744 87 1746 103
rect 1832 87 1834 106
rect 1872 103 1874 122
rect 1894 120 1895 124
rect 1899 120 1900 124
rect 1894 119 1900 120
rect 1974 124 1980 125
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 2078 124 2084 125
rect 2078 120 2079 124
rect 2083 120 2084 124
rect 2078 119 2084 120
rect 2206 124 2212 125
rect 2206 120 2207 124
rect 2211 120 2212 124
rect 2206 119 2212 120
rect 2342 124 2348 125
rect 2342 120 2343 124
rect 2347 120 2348 124
rect 2342 119 2348 120
rect 2478 124 2484 125
rect 2478 120 2479 124
rect 2483 120 2484 124
rect 2478 119 2484 120
rect 2614 124 2620 125
rect 2614 120 2615 124
rect 2619 120 2620 124
rect 2614 119 2620 120
rect 2734 124 2740 125
rect 2734 120 2735 124
rect 2739 120 2740 124
rect 2734 119 2740 120
rect 2846 124 2852 125
rect 2846 120 2847 124
rect 2851 120 2852 124
rect 2846 119 2852 120
rect 2950 124 2956 125
rect 2950 120 2951 124
rect 2955 120 2956 124
rect 2950 119 2956 120
rect 3054 124 3060 125
rect 3054 120 3055 124
rect 3059 120 3060 124
rect 3054 119 3060 120
rect 3150 124 3156 125
rect 3150 120 3151 124
rect 3155 120 3156 124
rect 3150 119 3156 120
rect 3238 124 3244 125
rect 3238 120 3239 124
rect 3243 120 3244 124
rect 3238 119 3244 120
rect 3334 124 3340 125
rect 3334 120 3335 124
rect 3339 120 3340 124
rect 3334 119 3340 120
rect 3422 124 3428 125
rect 3422 120 3423 124
rect 3427 120 3428 124
rect 3422 119 3428 120
rect 3502 124 3508 125
rect 3502 120 3503 124
rect 3507 120 3508 124
rect 3590 123 3591 127
rect 3595 123 3596 127
rect 3590 122 3596 123
rect 3502 119 3508 120
rect 1896 103 1898 119
rect 1976 103 1978 119
rect 2080 103 2082 119
rect 2208 103 2210 119
rect 2344 103 2346 119
rect 2480 103 2482 119
rect 2616 103 2618 119
rect 2736 103 2738 119
rect 2848 103 2850 119
rect 2952 103 2954 119
rect 3056 103 3058 119
rect 3152 103 3154 119
rect 3240 103 3242 119
rect 3336 103 3338 119
rect 3424 103 3426 119
rect 3504 103 3506 119
rect 3592 103 3594 122
rect 1871 102 1875 103
rect 1871 97 1875 98
rect 1895 102 1899 103
rect 1895 97 1899 98
rect 1975 102 1979 103
rect 1975 97 1979 98
rect 2079 102 2083 103
rect 2079 97 2083 98
rect 2207 102 2211 103
rect 2207 97 2211 98
rect 2343 102 2347 103
rect 2343 97 2347 98
rect 2479 102 2483 103
rect 2479 97 2483 98
rect 2615 102 2619 103
rect 2615 97 2619 98
rect 2735 102 2739 103
rect 2735 97 2739 98
rect 2847 102 2851 103
rect 2847 97 2851 98
rect 2951 102 2955 103
rect 2951 97 2955 98
rect 3055 102 3059 103
rect 3055 97 3059 98
rect 3151 102 3155 103
rect 3151 97 3155 98
rect 3239 102 3243 103
rect 3239 97 3243 98
rect 3335 102 3339 103
rect 3335 97 3339 98
rect 3423 102 3427 103
rect 3423 97 3427 98
rect 3503 102 3507 103
rect 3503 97 3507 98
rect 3591 102 3595 103
rect 3591 97 3595 98
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 215 86 219 87
rect 215 81 219 82
rect 295 86 299 87
rect 295 81 299 82
rect 375 86 379 87
rect 375 81 379 82
rect 455 86 459 87
rect 455 81 459 82
rect 535 86 539 87
rect 535 81 539 82
rect 615 86 619 87
rect 615 81 619 82
rect 695 86 699 87
rect 695 81 699 82
rect 775 86 779 87
rect 775 81 779 82
rect 855 86 859 87
rect 855 81 859 82
rect 935 86 939 87
rect 935 81 939 82
rect 1015 86 1019 87
rect 1015 81 1019 82
rect 1095 86 1099 87
rect 1095 81 1099 82
rect 1175 86 1179 87
rect 1175 81 1179 82
rect 1255 86 1259 87
rect 1255 81 1259 82
rect 1335 86 1339 87
rect 1335 81 1339 82
rect 1415 86 1419 87
rect 1415 81 1419 82
rect 1503 86 1507 87
rect 1503 81 1507 82
rect 1583 86 1587 87
rect 1583 81 1587 82
rect 1663 86 1667 87
rect 1663 81 1667 82
rect 1743 86 1747 87
rect 1743 81 1747 82
rect 1831 86 1835 87
rect 1831 81 1835 82
<< m4c >>
rect 111 3666 115 3670
rect 135 3666 139 3670
rect 215 3666 219 3670
rect 295 3666 299 3670
rect 1831 3666 1835 3670
rect 111 3590 115 3594
rect 1871 3598 1875 3602
rect 2063 3598 2067 3602
rect 2151 3598 2155 3602
rect 2255 3598 2259 3602
rect 2367 3598 2371 3602
rect 2479 3598 2483 3602
rect 2591 3598 2595 3602
rect 2703 3598 2707 3602
rect 2815 3598 2819 3602
rect 2919 3598 2923 3602
rect 143 3590 147 3594
rect 223 3590 227 3594
rect 303 3590 307 3594
rect 343 3590 347 3594
rect 471 3590 475 3594
rect 607 3590 611 3594
rect 743 3590 747 3594
rect 879 3590 883 3594
rect 999 3590 1003 3594
rect 1111 3590 1115 3594
rect 1223 3590 1227 3594
rect 1327 3590 1331 3594
rect 1423 3590 1427 3594
rect 1527 3590 1531 3594
rect 1631 3590 1635 3594
rect 1831 3590 1835 3594
rect 111 3514 115 3518
rect 135 3514 139 3518
rect 191 3514 195 3518
rect 215 3514 219 3518
rect 327 3514 331 3518
rect 335 3514 339 3518
rect 463 3514 467 3518
rect 471 3514 475 3518
rect 599 3514 603 3518
rect 623 3514 627 3518
rect 735 3514 739 3518
rect 775 3514 779 3518
rect 871 3514 875 3518
rect 1871 3522 1875 3526
rect 2055 3522 2059 3526
rect 919 3514 923 3518
rect 991 3514 995 3518
rect 1055 3514 1059 3518
rect 1103 3514 1107 3518
rect 1183 3514 1187 3518
rect 1215 3514 1219 3518
rect 1311 3514 1315 3518
rect 1319 3514 1323 3518
rect 1415 3514 1419 3518
rect 1439 3514 1443 3518
rect 1519 3514 1523 3518
rect 1567 3514 1571 3518
rect 111 3438 115 3442
rect 151 3438 155 3442
rect 199 3438 203 3442
rect 295 3438 299 3442
rect 335 3438 339 3442
rect 455 3438 459 3442
rect 479 3438 483 3442
rect 623 3438 627 3442
rect 631 3438 635 3442
rect 783 3438 787 3442
rect 791 3438 795 3442
rect 927 3438 931 3442
rect 959 3438 963 3442
rect 1063 3438 1067 3442
rect 1623 3514 1627 3518
rect 1831 3514 1835 3518
rect 2087 3522 2091 3526
rect 2143 3522 2147 3526
rect 2167 3522 2171 3526
rect 2247 3522 2251 3526
rect 2263 3522 2267 3526
rect 2359 3522 2363 3526
rect 2367 3522 2371 3526
rect 1119 3438 1123 3442
rect 1191 3438 1195 3442
rect 1271 3438 1275 3442
rect 1319 3438 1323 3442
rect 1415 3438 1419 3442
rect 1447 3438 1451 3442
rect 1559 3438 1563 3442
rect 1575 3438 1579 3442
rect 1711 3438 1715 3442
rect 1831 3438 1835 3442
rect 1871 3438 1875 3442
rect 2095 3438 2099 3442
rect 2111 3438 2115 3442
rect 2175 3438 2179 3442
rect 2199 3438 2203 3442
rect 111 3362 115 3366
rect 143 3362 147 3366
rect 207 3362 211 3366
rect 287 3362 291 3366
rect 335 3362 339 3366
rect 447 3362 451 3366
rect 471 3362 475 3366
rect 615 3362 619 3366
rect 623 3362 627 3366
rect 223 3296 227 3300
rect 111 3282 115 3286
rect 215 3282 219 3286
rect 343 3282 347 3286
rect 351 3282 355 3286
rect 783 3362 787 3366
rect 943 3362 947 3366
rect 951 3362 955 3366
rect 1103 3362 1107 3366
rect 1111 3362 1115 3366
rect 1263 3362 1267 3366
rect 1407 3362 1411 3366
rect 1423 3362 1427 3366
rect 1551 3362 1555 3366
rect 1583 3362 1587 3366
rect 1703 3362 1707 3366
rect 679 3296 683 3300
rect 455 3282 459 3286
rect 479 3282 483 3286
rect 575 3282 579 3286
rect 631 3282 635 3286
rect 703 3282 707 3286
rect 791 3282 795 3286
rect 839 3282 843 3286
rect 951 3282 955 3286
rect 983 3282 987 3286
rect 1111 3282 1115 3286
rect 1119 3282 1123 3286
rect 1255 3282 1259 3286
rect 111 3206 115 3210
rect 343 3206 347 3210
rect 447 3206 451 3210
rect 487 3206 491 3210
rect 567 3206 571 3210
rect 575 3206 579 3210
rect 663 3206 667 3210
rect 695 3206 699 3210
rect 767 3206 771 3210
rect 831 3206 835 3210
rect 887 3206 891 3210
rect 975 3206 979 3210
rect 1743 3362 1747 3366
rect 1831 3362 1835 3366
rect 2471 3522 2475 3526
rect 2487 3522 2491 3526
rect 2583 3522 2587 3526
rect 2615 3522 2619 3526
rect 2695 3522 2699 3526
rect 2743 3522 2747 3526
rect 2807 3522 2811 3526
rect 3015 3598 3019 3602
rect 3111 3598 3115 3602
rect 3207 3598 3211 3602
rect 3303 3598 3307 3602
rect 3399 3598 3403 3602
rect 3591 3598 3595 3602
rect 2871 3522 2875 3526
rect 2911 3522 2915 3526
rect 2991 3522 2995 3526
rect 3007 3522 3011 3526
rect 3103 3522 3107 3526
rect 3119 3522 3123 3526
rect 2271 3438 2275 3442
rect 2303 3438 2307 3442
rect 2375 3438 2379 3442
rect 2415 3438 2419 3442
rect 2495 3438 2499 3442
rect 2543 3438 2547 3442
rect 2623 3438 2627 3442
rect 2679 3438 2683 3442
rect 2751 3438 2755 3442
rect 2815 3438 2819 3442
rect 2879 3438 2883 3442
rect 2959 3438 2963 3442
rect 1871 3358 1875 3362
rect 2103 3358 2107 3362
rect 2127 3358 2131 3362
rect 2191 3358 2195 3362
rect 2223 3358 2227 3362
rect 2295 3358 2299 3362
rect 2335 3358 2339 3362
rect 2407 3358 2411 3362
rect 3199 3522 3203 3526
rect 3247 3522 3251 3526
rect 3295 3522 3299 3526
rect 3375 3522 3379 3526
rect 3391 3522 3395 3526
rect 3591 3522 3595 3526
rect 2999 3438 3003 3442
rect 3111 3438 3115 3442
rect 3127 3438 3131 3442
rect 3255 3438 3259 3442
rect 3263 3438 3267 3442
rect 3383 3438 3387 3442
rect 3423 3438 3427 3442
rect 2455 3358 2459 3362
rect 2535 3358 2539 3362
rect 1271 3282 1275 3286
rect 1383 3282 1387 3286
rect 1431 3282 1435 3286
rect 1511 3282 1515 3286
rect 1591 3282 1595 3286
rect 1639 3282 1643 3286
rect 1751 3282 1755 3286
rect 1831 3282 1835 3286
rect 1871 3270 1875 3274
rect 2135 3270 2139 3274
rect 2583 3358 2587 3362
rect 2671 3358 2675 3362
rect 2719 3358 2723 3362
rect 2807 3358 2811 3362
rect 2863 3358 2867 3362
rect 2951 3358 2955 3362
rect 3007 3358 3011 3362
rect 3103 3358 3107 3362
rect 3591 3438 3595 3442
rect 3159 3358 3163 3362
rect 3255 3358 3259 3362
rect 2231 3270 2235 3274
rect 2279 3270 2283 3274
rect 2343 3270 2347 3274
rect 2415 3270 2419 3274
rect 2463 3270 2467 3274
rect 1023 3206 1027 3210
rect 1111 3206 1115 3210
rect 1191 3206 1195 3210
rect 1247 3206 1251 3210
rect 1375 3206 1379 3210
rect 1503 3206 1507 3210
rect 1567 3206 1571 3210
rect 1631 3206 1635 3210
rect 1743 3206 1747 3210
rect 635 3144 639 3148
rect 111 3126 115 3130
rect 495 3126 499 3130
rect 583 3126 587 3130
rect 591 3126 595 3130
rect 843 3144 847 3148
rect 1207 3144 1211 3148
rect 1487 3144 1491 3148
rect 671 3126 675 3130
rect 759 3126 763 3130
rect 775 3126 779 3130
rect 847 3126 851 3130
rect 895 3126 899 3130
rect 935 3126 939 3130
rect 1023 3126 1027 3130
rect 1031 3126 1035 3130
rect 1111 3126 1115 3130
rect 1199 3126 1203 3130
rect 1287 3126 1291 3130
rect 1375 3126 1379 3130
rect 1383 3126 1387 3130
rect 111 3046 115 3050
rect 543 3046 547 3050
rect 583 3046 587 3050
rect 623 3046 627 3050
rect 663 3046 667 3050
rect 711 3046 715 3050
rect 751 3046 755 3050
rect 807 3046 811 3050
rect 839 3046 843 3050
rect 903 3046 907 3050
rect 927 3046 931 3050
rect 111 2970 115 2974
rect 471 2970 475 2974
rect 551 2970 555 2974
rect 575 2970 579 2974
rect 631 2970 635 2974
rect 687 2970 691 2974
rect 999 3046 1003 3050
rect 1015 3046 1019 3050
rect 1831 3206 1835 3210
rect 1871 3190 1875 3194
rect 1895 3190 1899 3194
rect 1991 3190 1995 3194
rect 2119 3190 2123 3194
rect 2127 3190 2131 3194
rect 2247 3190 2251 3194
rect 1575 3126 1579 3130
rect 1751 3126 1755 3130
rect 2551 3270 2555 3274
rect 2591 3270 2595 3274
rect 2687 3270 2691 3274
rect 2727 3270 2731 3274
rect 2823 3270 2827 3274
rect 2871 3270 2875 3274
rect 2959 3270 2963 3274
rect 3311 3358 3315 3362
rect 3415 3358 3419 3362
rect 3471 3358 3475 3362
rect 3591 3358 3595 3362
rect 3015 3270 3019 3274
rect 3095 3270 3099 3274
rect 3167 3270 3171 3274
rect 3231 3270 3235 3274
rect 3319 3270 3323 3274
rect 3375 3270 3379 3274
rect 3479 3270 3483 3274
rect 3511 3270 3515 3274
rect 2271 3190 2275 3194
rect 2383 3190 2387 3194
rect 2407 3190 2411 3194
rect 2511 3190 2515 3194
rect 2543 3190 2547 3194
rect 1831 3126 1835 3130
rect 1871 3098 1875 3102
rect 1903 3098 1907 3102
rect 1999 3098 2003 3102
rect 2015 3098 2019 3102
rect 2127 3098 2131 3102
rect 1911 3091 1915 3092
rect 1911 3088 1915 3091
rect 2191 3098 2195 3102
rect 2255 3098 2259 3102
rect 2391 3098 2395 3102
rect 2407 3098 2411 3102
rect 2199 3088 2203 3092
rect 1087 3046 1091 3050
rect 1103 3046 1107 3050
rect 1183 3046 1187 3050
rect 1191 3046 1195 3050
rect 1279 3046 1283 3050
rect 1367 3046 1371 3050
rect 1375 3046 1379 3050
rect 1471 3046 1475 3050
rect 1831 3046 1835 3050
rect 1871 3014 1875 3018
rect 719 2970 723 2974
rect 807 2970 811 2974
rect 815 2970 819 2974
rect 911 2970 915 2974
rect 1895 3014 1899 3018
rect 2007 3014 2011 3018
rect 943 2970 947 2974
rect 1007 2970 1011 2974
rect 1087 2970 1091 2974
rect 1095 2970 1099 2974
rect 1191 2970 1195 2974
rect 1247 2970 1251 2974
rect 1287 2970 1291 2974
rect 1383 2970 1387 2974
rect 1415 2970 1419 2974
rect 1479 2970 1483 2974
rect 1591 2970 1595 2974
rect 655 2944 659 2948
rect 951 2944 955 2948
rect 1103 2944 1107 2948
rect 1307 2944 1311 2948
rect 111 2894 115 2898
rect 311 2894 315 2898
rect 431 2894 435 2898
rect 463 2894 467 2898
rect 327 2832 331 2836
rect 111 2818 115 2822
rect 167 2818 171 2822
rect 303 2818 307 2822
rect 319 2818 323 2822
rect 551 2894 555 2898
rect 567 2894 571 2898
rect 679 2894 683 2898
rect 799 2894 803 2898
rect 815 2894 819 2898
rect 935 2894 939 2898
rect 951 2894 955 2898
rect 1079 2894 1083 2898
rect 1087 2894 1091 2898
rect 1223 2894 1227 2898
rect 1239 2894 1243 2898
rect 1751 2970 1755 2974
rect 1831 2970 1835 2974
rect 1871 2938 1875 2942
rect 1359 2894 1363 2898
rect 1407 2894 1411 2898
rect 1495 2894 1499 2898
rect 1583 2894 1587 2898
rect 1631 2894 1635 2898
rect 2047 3014 2051 3018
rect 2183 3014 2187 3018
rect 2223 3014 2227 3018
rect 2639 3190 2643 3194
rect 2679 3190 2683 3194
rect 2767 3190 2771 3194
rect 2815 3190 2819 3194
rect 2895 3190 2899 3194
rect 2951 3190 2955 3194
rect 3031 3190 3035 3194
rect 3087 3190 3091 3194
rect 3175 3190 3179 3194
rect 3223 3190 3227 3194
rect 3591 3270 3595 3274
rect 3327 3190 3331 3194
rect 3367 3190 3371 3194
rect 2519 3098 2523 3102
rect 2647 3098 2651 3102
rect 2655 3098 2659 3102
rect 2775 3098 2779 3102
rect 2903 3098 2907 3102
rect 2935 3098 2939 3102
rect 3039 3098 3043 3102
rect 3183 3098 3187 3102
rect 3231 3098 3235 3102
rect 2415 3088 2419 3092
rect 2943 3088 2947 3092
rect 3487 3190 3491 3194
rect 3503 3190 3507 3194
rect 3591 3190 3595 3194
rect 3335 3098 3339 3102
rect 3495 3098 3499 3102
rect 3511 3098 3515 3102
rect 3591 3098 3595 3102
rect 2391 3014 2395 3018
rect 2399 3014 2403 3018
rect 2543 3014 2547 3018
rect 2647 3014 2651 3018
rect 2687 3014 2691 3018
rect 2815 3014 2819 3018
rect 2927 3014 2931 3018
rect 3039 3014 3043 3018
rect 3143 3014 3147 3018
rect 3223 3014 3227 3018
rect 3239 3014 3243 3018
rect 3335 3014 3339 3018
rect 3423 3014 3427 3018
rect 3503 3014 3507 3018
rect 2567 2952 2571 2956
rect 1903 2938 1907 2942
rect 2055 2938 2059 2942
rect 2087 2938 2091 2942
rect 2231 2938 2235 2942
rect 2295 2938 2299 2942
rect 2399 2938 2403 2942
rect 2487 2938 2491 2942
rect 1743 2894 1747 2898
rect 763 2832 767 2836
rect 439 2818 443 2822
rect 447 2818 451 2822
rect 559 2818 563 2822
rect 607 2818 611 2822
rect 687 2818 691 2822
rect 783 2818 787 2822
rect 823 2818 827 2822
rect 959 2818 963 2822
rect 1095 2818 1099 2822
rect 1143 2818 1147 2822
rect 1231 2818 1235 2822
rect 1335 2818 1339 2822
rect 1367 2818 1371 2822
rect 1503 2818 1507 2822
rect 1535 2818 1539 2822
rect 111 2738 115 2742
rect 135 2738 139 2742
rect 159 2738 163 2742
rect 247 2738 251 2742
rect 295 2738 299 2742
rect 111 2662 115 2666
rect 263 2672 267 2676
rect 391 2738 395 2742
rect 439 2738 443 2742
rect 551 2738 555 2742
rect 599 2738 603 2742
rect 711 2738 715 2742
rect 775 2738 779 2742
rect 879 2738 883 2742
rect 951 2738 955 2742
rect 1039 2738 1043 2742
rect 1135 2738 1139 2742
rect 1199 2738 1203 2742
rect 1831 2894 1835 2898
rect 1871 2854 1875 2858
rect 1895 2854 1899 2858
rect 2079 2854 2083 2858
rect 2551 2938 2555 2942
rect 2671 2938 2675 2942
rect 2695 2938 2699 2942
rect 2823 2938 2827 2942
rect 2839 2938 2843 2942
rect 2715 2931 2719 2932
rect 2715 2928 2719 2931
rect 2919 2952 2923 2956
rect 2935 2938 2939 2942
rect 2999 2938 3003 2942
rect 3047 2938 3051 2942
rect 3151 2938 3155 2942
rect 3247 2938 3251 2942
rect 3303 2938 3307 2942
rect 3343 2938 3347 2942
rect 3591 3014 3595 3018
rect 3431 2938 3435 2942
rect 3455 2938 3459 2942
rect 3511 2938 3515 2942
rect 3591 2938 3595 2942
rect 3311 2928 3315 2932
rect 2135 2854 2139 2858
rect 2263 2854 2267 2858
rect 2287 2854 2291 2858
rect 2391 2854 2395 2858
rect 2479 2854 2483 2858
rect 2519 2854 2523 2858
rect 2647 2854 2651 2858
rect 2663 2854 2667 2858
rect 2767 2854 2771 2858
rect 2831 2854 2835 2858
rect 1639 2818 1643 2822
rect 1735 2818 1739 2822
rect 1751 2818 1755 2822
rect 1831 2818 1835 2822
rect 2663 2800 2667 2804
rect 1871 2770 1875 2774
rect 2143 2770 2147 2774
rect 2231 2770 2235 2774
rect 2271 2770 2275 2774
rect 2311 2770 2315 2774
rect 2391 2770 2395 2774
rect 2399 2770 2403 2774
rect 2471 2770 2475 2774
rect 2527 2770 2531 2774
rect 2551 2770 2555 2774
rect 1327 2738 1331 2742
rect 1359 2738 1363 2742
rect 1519 2738 1523 2742
rect 1527 2738 1531 2742
rect 1687 2738 1691 2742
rect 651 2672 655 2676
rect 143 2662 147 2666
rect 255 2662 259 2666
rect 399 2662 403 2666
rect 551 2662 555 2666
rect 559 2662 563 2666
rect 711 2662 715 2666
rect 719 2662 723 2666
rect 879 2662 883 2666
rect 887 2662 891 2666
rect 1047 2662 1051 2666
rect 1207 2662 1211 2666
rect 1215 2662 1219 2666
rect 111 2582 115 2586
rect 135 2582 139 2586
rect 159 2582 163 2586
rect 247 2582 251 2586
rect 279 2582 283 2586
rect 391 2582 395 2586
rect 415 2582 419 2586
rect 543 2582 547 2586
rect 559 2582 563 2586
rect 703 2582 707 2586
rect 847 2582 851 2586
rect 871 2582 875 2586
rect 983 2582 987 2586
rect 1039 2582 1043 2586
rect 1119 2582 1123 2586
rect 1727 2738 1731 2742
rect 1831 2738 1835 2742
rect 2639 2770 2643 2774
rect 2655 2770 2659 2774
rect 2727 2770 2731 2774
rect 2775 2770 2779 2774
rect 2815 2770 2819 2774
rect 2647 2763 2651 2764
rect 2647 2760 2651 2763
rect 2887 2854 2891 2858
rect 2991 2854 2995 2858
rect 3007 2854 3011 2858
rect 3135 2854 3139 2858
rect 3143 2854 3147 2858
rect 3295 2854 3299 2858
rect 3447 2854 3451 2858
rect 3591 2854 3595 2858
rect 3087 2800 3091 2804
rect 2895 2770 2899 2774
rect 2903 2770 2907 2774
rect 2991 2770 2995 2774
rect 3015 2770 3019 2774
rect 3143 2770 3147 2774
rect 3591 2770 3595 2774
rect 2999 2760 3003 2764
rect 1871 2694 1875 2698
rect 2223 2694 2227 2698
rect 2239 2694 2243 2698
rect 2303 2694 2307 2698
rect 2319 2694 2323 2698
rect 2383 2694 2387 2698
rect 2399 2694 2403 2698
rect 2463 2694 2467 2698
rect 2479 2694 2483 2698
rect 2543 2694 2547 2698
rect 2559 2694 2563 2698
rect 2631 2694 2635 2698
rect 2639 2694 2643 2698
rect 2719 2694 2723 2698
rect 1367 2662 1371 2666
rect 1391 2662 1395 2666
rect 1527 2662 1531 2666
rect 1567 2662 1571 2666
rect 1695 2662 1699 2666
rect 1831 2662 1835 2666
rect 1871 2610 1875 2614
rect 1207 2582 1211 2586
rect 1255 2582 1259 2586
rect 1383 2582 1387 2586
rect 1391 2582 1395 2586
rect 1527 2582 1531 2586
rect 175 2552 179 2556
rect 643 2552 647 2556
rect 355 2520 359 2524
rect 111 2502 115 2506
rect 167 2502 171 2506
rect 287 2502 291 2506
rect 335 2502 339 2506
rect 667 2520 671 2524
rect 415 2502 419 2506
rect 423 2502 427 2506
rect 503 2502 507 2506
rect 567 2502 571 2506
rect 599 2502 603 2506
rect 703 2502 707 2506
rect 711 2502 715 2506
rect 815 2502 819 2506
rect 855 2502 859 2506
rect 935 2502 939 2506
rect 991 2502 995 2506
rect 1063 2502 1067 2506
rect 1127 2502 1131 2506
rect 1191 2502 1195 2506
rect 1263 2502 1267 2506
rect 2191 2610 2195 2614
rect 2247 2610 2251 2614
rect 2271 2610 2275 2614
rect 2327 2610 2331 2614
rect 2351 2610 2355 2614
rect 2407 2610 2411 2614
rect 2431 2610 2435 2614
rect 2487 2610 2491 2614
rect 1559 2582 1563 2586
rect 1831 2582 1835 2586
rect 1871 2526 1875 2530
rect 2119 2526 2123 2530
rect 2183 2526 2187 2530
rect 2207 2526 2211 2530
rect 2263 2526 2267 2530
rect 2303 2526 2307 2530
rect 2343 2526 2347 2530
rect 2399 2526 2403 2530
rect 2423 2526 2427 2530
rect 1327 2502 1331 2506
rect 1399 2502 1403 2506
rect 1471 2502 1475 2506
rect 1535 2502 1539 2506
rect 1831 2502 1835 2506
rect 111 2418 115 2422
rect 327 2418 331 2422
rect 383 2418 387 2422
rect 407 2418 411 2422
rect 463 2418 467 2422
rect 495 2418 499 2422
rect 543 2418 547 2422
rect 591 2418 595 2422
rect 623 2418 627 2422
rect 695 2418 699 2422
rect 703 2418 707 2422
rect 783 2418 787 2422
rect 111 2342 115 2346
rect 391 2342 395 2346
rect 471 2342 475 2346
rect 551 2342 555 2346
rect 631 2342 635 2346
rect 711 2342 715 2346
rect 791 2342 795 2346
rect 807 2418 811 2422
rect 863 2418 867 2422
rect 927 2418 931 2422
rect 943 2418 947 2422
rect 1023 2418 1027 2422
rect 1055 2418 1059 2422
rect 1103 2418 1107 2422
rect 1183 2418 1187 2422
rect 1263 2418 1267 2422
rect 2511 2610 2515 2614
rect 2567 2610 2571 2614
rect 2591 2610 2595 2614
rect 2799 2694 2803 2698
rect 2807 2694 2811 2698
rect 2879 2694 2883 2698
rect 2895 2694 2899 2698
rect 2959 2694 2963 2698
rect 2983 2694 2987 2698
rect 3591 2694 3595 2698
rect 2647 2610 2651 2614
rect 2671 2610 2675 2614
rect 2727 2610 2731 2614
rect 2751 2610 2755 2614
rect 2807 2610 2811 2614
rect 2831 2610 2835 2614
rect 2887 2610 2891 2614
rect 2911 2610 2915 2614
rect 2967 2610 2971 2614
rect 2991 2610 2995 2614
rect 3591 2610 3595 2614
rect 2495 2526 2499 2530
rect 2503 2526 2507 2530
rect 2583 2526 2587 2530
rect 2591 2526 2595 2530
rect 1319 2418 1323 2422
rect 1351 2418 1355 2422
rect 1439 2418 1443 2422
rect 1463 2418 1467 2422
rect 871 2342 875 2346
rect 951 2342 955 2346
rect 1031 2342 1035 2346
rect 1111 2342 1115 2346
rect 1191 2342 1195 2346
rect 1271 2342 1275 2346
rect 1359 2342 1363 2346
rect 1407 2342 1411 2346
rect 1871 2446 1875 2450
rect 1903 2446 1907 2450
rect 1991 2446 1995 2450
rect 2111 2446 2115 2450
rect 2127 2446 2131 2450
rect 1527 2418 1531 2422
rect 1831 2418 1835 2422
rect 1947 2408 1951 2412
rect 2663 2526 2667 2530
rect 2687 2526 2691 2530
rect 2743 2526 2747 2530
rect 2783 2526 2787 2530
rect 2823 2526 2827 2530
rect 2879 2526 2883 2530
rect 2903 2526 2907 2530
rect 2975 2526 2979 2530
rect 2983 2526 2987 2530
rect 3079 2526 3083 2530
rect 3591 2526 3595 2530
rect 2703 2464 2707 2468
rect 2215 2446 2219 2450
rect 2247 2446 2251 2450
rect 2311 2446 2315 2450
rect 2391 2446 2395 2450
rect 2407 2446 2411 2450
rect 2503 2446 2507 2450
rect 2535 2446 2539 2450
rect 2599 2446 2603 2450
rect 2671 2446 2675 2450
rect 2695 2446 2699 2450
rect 2179 2432 2183 2436
rect 2543 2432 2547 2436
rect 3051 2464 3055 2468
rect 2791 2446 2795 2450
rect 2807 2446 2811 2450
rect 2887 2446 2891 2450
rect 2943 2446 2947 2450
rect 2983 2446 2987 2450
rect 3079 2446 3083 2450
rect 3087 2446 3091 2450
rect 3215 2446 3219 2450
rect 3591 2446 3595 2450
rect 2459 2408 2463 2412
rect 1447 2342 1451 2346
rect 1871 2362 1875 2366
rect 1895 2362 1899 2366
rect 1983 2362 1987 2366
rect 2015 2362 2019 2366
rect 2103 2362 2107 2366
rect 2175 2362 2179 2366
rect 2239 2362 2243 2366
rect 2343 2362 2347 2366
rect 2383 2362 2387 2366
rect 1487 2342 1491 2346
rect 1535 2342 1539 2346
rect 1567 2342 1571 2346
rect 1647 2342 1651 2346
rect 1831 2342 1835 2346
rect 2511 2362 2515 2366
rect 2527 2362 2531 2366
rect 2663 2362 2667 2366
rect 2671 2362 2675 2366
rect 2799 2362 2803 2366
rect 2823 2362 2827 2366
rect 2935 2362 2939 2366
rect 2959 2362 2963 2366
rect 3071 2362 3075 2366
rect 3079 2362 3083 2366
rect 111 2258 115 2262
rect 135 2258 139 2262
rect 215 2258 219 2262
rect 295 2258 299 2262
rect 383 2258 387 2262
rect 519 2258 523 2262
rect 671 2258 675 2262
rect 831 2258 835 2262
rect 999 2258 1003 2262
rect 1159 2258 1163 2262
rect 1311 2258 1315 2262
rect 1399 2258 1403 2262
rect 1455 2258 1459 2262
rect 1479 2258 1483 2262
rect 1559 2258 1563 2262
rect 1175 2240 1179 2244
rect 1871 2286 1875 2290
rect 2687 2296 2691 2300
rect 1903 2286 1907 2290
rect 1607 2258 1611 2262
rect 1639 2258 1643 2262
rect 1743 2258 1747 2262
rect 1831 2258 1835 2262
rect 111 2178 115 2182
rect 143 2178 147 2182
rect 191 2178 195 2182
rect 223 2178 227 2182
rect 303 2178 307 2182
rect 311 2178 315 2182
rect 391 2178 395 2182
rect 463 2178 467 2182
rect 527 2178 531 2182
rect 639 2178 643 2182
rect 679 2178 683 2182
rect 823 2178 827 2182
rect 839 2178 843 2182
rect 199 2171 203 2172
rect 199 2168 203 2171
rect 111 2098 115 2102
rect 183 2098 187 2102
rect 215 2098 219 2102
rect 471 2168 475 2172
rect 647 2171 651 2172
rect 647 2168 651 2171
rect 1579 2240 1583 2244
rect 2023 2286 2027 2290
rect 2031 2286 2035 2290
rect 2183 2286 2187 2290
rect 2351 2286 2355 2290
rect 2367 2286 2371 2290
rect 2519 2286 2523 2290
rect 2575 2286 2579 2290
rect 3191 2362 3195 2366
rect 3207 2362 3211 2366
rect 3303 2362 3307 2366
rect 3415 2362 3419 2366
rect 3503 2362 3507 2366
rect 3591 2362 3595 2366
rect 3139 2296 3143 2300
rect 2679 2286 2683 2290
rect 2791 2286 2795 2290
rect 2831 2286 2835 2290
rect 2967 2286 2971 2290
rect 3023 2286 3027 2290
rect 3087 2286 3091 2290
rect 3199 2286 3203 2290
rect 3255 2286 3259 2290
rect 3311 2286 3315 2290
rect 1207 2192 1211 2196
rect 1007 2178 1011 2182
rect 1015 2178 1019 2182
rect 1167 2178 1171 2182
rect 1199 2178 1203 2182
rect 1023 2168 1027 2172
rect 1691 2192 1695 2196
rect 1871 2190 1875 2194
rect 1895 2190 1899 2194
rect 2023 2190 2027 2194
rect 2175 2190 2179 2194
rect 2199 2190 2203 2194
rect 2295 2190 2299 2194
rect 2359 2190 2363 2194
rect 2399 2190 2403 2194
rect 1319 2178 1323 2182
rect 1391 2178 1395 2182
rect 1463 2178 1467 2182
rect 1583 2178 1587 2182
rect 1615 2178 1619 2182
rect 1751 2178 1755 2182
rect 1831 2178 1835 2182
rect 3423 2286 3427 2290
rect 3495 2286 3499 2290
rect 3511 2286 3515 2290
rect 3591 2286 3595 2290
rect 2519 2190 2523 2194
rect 2567 2190 2571 2194
rect 2639 2190 2643 2194
rect 2759 2190 2763 2194
rect 2783 2190 2787 2194
rect 2879 2190 2883 2194
rect 2991 2190 2995 2194
rect 3015 2190 3019 2194
rect 3095 2190 3099 2194
rect 3199 2190 3203 2194
rect 3247 2190 3251 2194
rect 3303 2190 3307 2194
rect 303 2098 307 2102
rect 359 2098 363 2102
rect 455 2098 459 2102
rect 519 2098 523 2102
rect 631 2098 635 2102
rect 703 2098 707 2102
rect 815 2098 819 2102
rect 895 2098 899 2102
rect 1007 2098 1011 2102
rect 1103 2098 1107 2102
rect 1191 2098 1195 2102
rect 1311 2098 1315 2102
rect 1383 2098 1387 2102
rect 1527 2098 1531 2102
rect 1575 2098 1579 2102
rect 1743 2098 1747 2102
rect 111 2022 115 2026
rect 143 2022 147 2026
rect 223 2022 227 2026
rect 263 2022 267 2026
rect 367 2022 371 2026
rect 383 2022 387 2026
rect 111 1938 115 1942
rect 135 1938 139 1942
rect 495 2022 499 2026
rect 527 2022 531 2026
rect 607 2022 611 2026
rect 711 2022 715 2026
rect 719 2022 723 2026
rect 823 2022 827 2026
rect 903 2022 907 2026
rect 927 2022 931 2026
rect 1023 2022 1027 2026
rect 167 1938 171 1942
rect 255 1938 259 1942
rect 327 1938 331 1942
rect 375 1938 379 1942
rect 487 1938 491 1942
rect 599 1938 603 1942
rect 647 1938 651 1942
rect 711 1938 715 1942
rect 111 1862 115 1866
rect 159 1862 163 1866
rect 175 1862 179 1866
rect 303 1862 307 1866
rect 183 1840 187 1844
rect 335 1862 339 1866
rect 447 1862 451 1866
rect 495 1862 499 1866
rect 111 1782 115 1786
rect 151 1782 155 1786
rect 247 1782 251 1786
rect 295 1782 299 1786
rect 423 1782 427 1786
rect 799 1938 803 1942
rect 815 1938 819 1942
rect 1111 2022 1115 2026
rect 1207 2022 1211 2026
rect 1295 2022 1299 2026
rect 1319 2022 1323 2026
rect 1391 2022 1395 2026
rect 1487 2022 1491 2026
rect 1535 2022 1539 2026
rect 1583 2022 1587 2026
rect 2215 2128 2219 2132
rect 2487 2128 2491 2132
rect 1831 2098 1835 2102
rect 1871 2102 1875 2106
rect 2175 2102 2179 2106
rect 2207 2102 2211 2106
rect 2271 2102 2275 2106
rect 2303 2102 2307 2106
rect 2375 2102 2379 2106
rect 2407 2102 2411 2106
rect 2487 2102 2491 2106
rect 1671 2022 1675 2026
rect 1751 2022 1755 2026
rect 1831 2022 1835 2026
rect 1871 2022 1875 2026
rect 2071 2022 2075 2026
rect 2167 2022 2171 2026
rect 2207 2022 2211 2026
rect 2263 2022 2267 2026
rect 2359 2022 2363 2026
rect 2367 2022 2371 2026
rect 2527 2102 2531 2106
rect 2607 2102 2611 2106
rect 2647 2102 2651 2106
rect 2727 2102 2731 2106
rect 3407 2190 3411 2194
rect 3487 2190 3491 2194
rect 3503 2190 3507 2194
rect 3591 2190 3595 2194
rect 2767 2102 2771 2106
rect 2847 2102 2851 2106
rect 2887 2102 2891 2106
rect 2967 2102 2971 2106
rect 2999 2102 3003 2106
rect 3079 2102 3083 2106
rect 3103 2102 3107 2106
rect 3191 2102 3195 2106
rect 3207 2102 3211 2106
rect 3303 2102 3307 2106
rect 3311 2102 3315 2106
rect 3415 2102 3419 2106
rect 3511 2102 3515 2106
rect 3591 2102 3595 2106
rect 2479 2022 2483 2026
rect 2519 2022 2523 2026
rect 2599 2022 2603 2026
rect 2679 2022 2683 2026
rect 2719 2022 2723 2026
rect 2839 2022 2843 2026
rect 2847 2022 2851 2026
rect 2959 2022 2963 2026
rect 3015 2022 3019 2026
rect 919 1938 923 1942
rect 943 1938 947 1942
rect 1015 1938 1019 1942
rect 1079 1938 1083 1942
rect 1103 1938 1107 1942
rect 1199 1938 1203 1942
rect 1215 1938 1219 1942
rect 1287 1938 1291 1942
rect 1351 1938 1355 1942
rect 1383 1938 1387 1942
rect 1479 1938 1483 1942
rect 1487 1938 1491 1942
rect 1575 1938 1579 1942
rect 1623 1938 1627 1942
rect 1663 1938 1667 1942
rect 1743 1938 1747 1942
rect 599 1862 603 1866
rect 655 1862 659 1866
rect 751 1862 755 1866
rect 807 1862 811 1866
rect 903 1862 907 1866
rect 951 1862 955 1866
rect 1055 1862 1059 1866
rect 455 1840 459 1844
rect 1087 1862 1091 1866
rect 1207 1862 1211 1866
rect 1223 1862 1227 1866
rect 2383 1968 2387 1972
rect 1871 1946 1875 1950
rect 1903 1946 1907 1950
rect 2007 1946 2011 1950
rect 1831 1938 1835 1942
rect 2079 1946 2083 1950
rect 2135 1946 2139 1950
rect 2215 1946 2219 1950
rect 2255 1946 2259 1950
rect 2367 1946 2371 1950
rect 2375 1946 2379 1950
rect 1871 1870 1875 1874
rect 1895 1870 1899 1874
rect 1351 1862 1355 1866
rect 1359 1862 1363 1866
rect 1487 1862 1491 1866
rect 1495 1862 1499 1866
rect 1631 1862 1635 1866
rect 1751 1862 1755 1866
rect 1831 1862 1835 1866
rect 439 1782 443 1786
rect 591 1782 595 1786
rect 743 1782 747 1786
rect 751 1782 755 1786
rect 111 1702 115 1706
rect 191 1702 195 1706
rect 255 1702 259 1706
rect 311 1702 315 1706
rect 431 1702 435 1706
rect 447 1702 451 1706
rect 111 1618 115 1622
rect 167 1618 171 1622
rect 895 1782 899 1786
rect 1023 1782 1027 1786
rect 1047 1782 1051 1786
rect 1143 1782 1147 1786
rect 1199 1782 1203 1786
rect 1991 1870 1995 1874
rect 1999 1870 2003 1874
rect 2119 1870 2123 1874
rect 2127 1870 2131 1874
rect 2247 1870 2251 1874
rect 2599 1968 2603 1972
rect 3071 2022 3075 2026
rect 3183 2022 3187 2026
rect 3295 2022 3299 2026
rect 3351 2022 3355 2026
rect 3407 2022 3411 2026
rect 3503 2022 3507 2026
rect 2487 1946 2491 1950
rect 2527 1946 2531 1950
rect 2599 1946 2603 1950
rect 2687 1946 2691 1950
rect 2719 1946 2723 1950
rect 2839 1946 2843 1950
rect 3591 2022 3595 2026
rect 2855 1946 2859 1950
rect 3023 1946 3027 1950
rect 3191 1946 3195 1950
rect 3359 1946 3363 1950
rect 3511 1946 3515 1950
rect 3591 1946 3595 1950
rect 2367 1870 2371 1874
rect 2383 1870 2387 1874
rect 2479 1870 2483 1874
rect 2519 1870 2523 1874
rect 2591 1870 2595 1874
rect 2655 1870 2659 1874
rect 2711 1870 2715 1874
rect 2807 1870 2811 1874
rect 2831 1870 2835 1874
rect 2975 1870 2979 1874
rect 3151 1870 3155 1874
rect 3335 1870 3339 1874
rect 3503 1870 3507 1874
rect 3591 1870 3595 1874
rect 2695 1792 2699 1796
rect 1263 1782 1267 1786
rect 1343 1782 1347 1786
rect 1391 1782 1395 1786
rect 1479 1782 1483 1786
rect 1623 1782 1627 1786
rect 1743 1782 1747 1786
rect 1831 1782 1835 1786
rect 1871 1782 1875 1786
rect 1903 1782 1907 1786
rect 1999 1782 2003 1786
rect 2031 1782 2035 1786
rect 2127 1782 2131 1786
rect 2191 1782 2195 1786
rect 2255 1782 2259 1786
rect 2359 1782 2363 1786
rect 2391 1782 2395 1786
rect 2527 1782 2531 1786
rect 2663 1782 2667 1786
rect 2687 1782 2691 1786
rect 911 1720 915 1724
rect 591 1702 595 1706
rect 599 1702 603 1706
rect 743 1702 747 1706
rect 759 1702 763 1706
rect 895 1702 899 1706
rect 903 1702 907 1706
rect 1031 1702 1035 1706
rect 1039 1702 1043 1706
rect 1151 1702 1155 1706
rect 1183 1702 1187 1706
rect 3259 1792 3263 1796
rect 2815 1782 2819 1786
rect 2839 1782 2843 1786
rect 2983 1782 2987 1786
rect 3119 1782 3123 1786
rect 3159 1782 3163 1786
rect 3255 1782 3259 1786
rect 3343 1782 3347 1786
rect 3391 1782 3395 1786
rect 3511 1782 3515 1786
rect 1343 1720 1347 1724
rect 1271 1702 1275 1706
rect 1319 1702 1323 1706
rect 1399 1702 1403 1706
rect 1447 1702 1451 1706
rect 1575 1702 1579 1706
rect 1711 1702 1715 1706
rect 1831 1702 1835 1706
rect 1871 1702 1875 1706
rect 1895 1702 1899 1706
rect 1991 1702 1995 1706
rect 2023 1702 2027 1706
rect 2135 1702 2139 1706
rect 2183 1702 2187 1706
rect 2295 1702 2299 1706
rect 2351 1702 2355 1706
rect 183 1618 187 1622
rect 303 1618 307 1622
rect 351 1618 355 1622
rect 439 1618 443 1622
rect 543 1618 547 1622
rect 583 1618 587 1622
rect 727 1618 731 1622
rect 735 1618 739 1622
rect 887 1618 891 1622
rect 903 1618 907 1622
rect 111 1538 115 1542
rect 143 1538 147 1542
rect 175 1538 179 1542
rect 247 1538 251 1542
rect 359 1538 363 1542
rect 383 1538 387 1542
rect 1031 1618 1035 1622
rect 1071 1618 1075 1622
rect 1175 1618 1179 1622
rect 1223 1618 1227 1622
rect 1311 1618 1315 1622
rect 1359 1618 1363 1622
rect 1439 1618 1443 1622
rect 1495 1618 1499 1622
rect 1567 1618 1571 1622
rect 1623 1618 1627 1622
rect 1703 1618 1707 1622
rect 1911 1688 1915 1692
rect 2471 1702 2475 1706
rect 2519 1702 2523 1706
rect 2647 1702 2651 1706
rect 2679 1702 2683 1706
rect 2815 1702 2819 1706
rect 2831 1702 2835 1706
rect 2967 1702 2971 1706
rect 2975 1702 2979 1706
rect 3111 1702 3115 1706
rect 3247 1702 3251 1706
rect 3383 1702 3387 1706
rect 2419 1688 2423 1692
rect 2831 1640 2835 1644
rect 1743 1618 1747 1622
rect 1831 1618 1835 1622
rect 1871 1622 1875 1626
rect 1903 1622 1907 1626
rect 1975 1622 1979 1626
rect 1999 1622 2003 1626
rect 2095 1622 2099 1626
rect 2143 1622 2147 1626
rect 2231 1622 2235 1626
rect 2303 1622 2307 1626
rect 2367 1622 2371 1626
rect 2479 1622 2483 1626
rect 2503 1622 2507 1626
rect 2639 1622 2643 1626
rect 2655 1622 2659 1626
rect 2775 1622 2779 1626
rect 2823 1622 2827 1626
rect 2911 1622 2915 1626
rect 2975 1622 2979 1626
rect 3055 1622 3059 1626
rect 3119 1622 3123 1626
rect 3187 1640 3191 1644
rect 3503 1702 3507 1706
rect 3207 1622 3211 1626
rect 3255 1622 3259 1626
rect 3367 1622 3371 1626
rect 3391 1622 3395 1626
rect 3511 1622 3515 1626
rect 527 1538 531 1542
rect 551 1538 555 1542
rect 671 1538 675 1542
rect 735 1538 739 1542
rect 815 1538 819 1542
rect 911 1538 915 1542
rect 951 1538 955 1542
rect 1079 1538 1083 1542
rect 1207 1538 1211 1542
rect 1231 1538 1235 1542
rect 1335 1538 1339 1542
rect 1367 1538 1371 1542
rect 1471 1538 1475 1542
rect 1503 1538 1507 1542
rect 111 1458 115 1462
rect 135 1458 139 1462
rect 231 1458 235 1462
rect 239 1458 243 1462
rect 359 1458 363 1462
rect 375 1458 379 1462
rect 479 1458 483 1462
rect 519 1458 523 1462
rect 599 1458 603 1462
rect 111 1366 115 1370
rect 143 1366 147 1370
rect 239 1366 243 1370
rect 287 1366 291 1370
rect 1631 1538 1635 1542
rect 1751 1538 1755 1542
rect 1831 1538 1835 1542
rect 1871 1542 1875 1546
rect 1967 1542 1971 1546
rect 2087 1542 2091 1546
rect 2167 1542 2171 1546
rect 2223 1542 2227 1546
rect 2255 1542 2259 1546
rect 2343 1542 2347 1546
rect 2359 1542 2363 1546
rect 2103 1528 2107 1532
rect 959 1472 963 1476
rect 1219 1472 1223 1476
rect 663 1458 667 1462
rect 719 1458 723 1462
rect 807 1458 811 1462
rect 831 1458 835 1462
rect 935 1458 939 1462
rect 943 1458 947 1462
rect 1039 1458 1043 1462
rect 1071 1458 1075 1462
rect 1143 1458 1147 1462
rect 1199 1458 1203 1462
rect 2439 1542 2443 1546
rect 2495 1542 2499 1546
rect 2535 1542 2539 1546
rect 2631 1542 2635 1546
rect 2647 1542 2651 1546
rect 2767 1542 2771 1546
rect 2783 1542 2787 1546
rect 2903 1542 2907 1546
rect 2419 1528 2423 1532
rect 2271 1472 2275 1476
rect 1255 1458 1259 1462
rect 1327 1458 1331 1462
rect 1463 1458 1467 1462
rect 1831 1458 1835 1462
rect 1871 1462 1875 1466
rect 2095 1462 2099 1466
rect 2175 1462 2179 1466
rect 2263 1462 2267 1466
rect 2515 1472 2519 1476
rect 2663 1480 2667 1484
rect 2343 1462 2347 1466
rect 2351 1462 2355 1466
rect 2423 1462 2427 1466
rect 2447 1462 2451 1466
rect 2503 1462 2507 1466
rect 2543 1462 2547 1466
rect 2607 1462 2611 1466
rect 2655 1462 2659 1466
rect 2735 1462 2739 1466
rect 2791 1462 2795 1466
rect 2943 1542 2947 1546
rect 3047 1542 3051 1546
rect 3119 1542 3123 1546
rect 3199 1542 3203 1546
rect 3303 1542 3307 1546
rect 3359 1542 3363 1546
rect 3203 1480 3207 1484
rect 2895 1462 2899 1466
rect 2951 1462 2955 1466
rect 3079 1462 3083 1466
rect 3127 1462 3131 1466
rect 3279 1462 3283 1466
rect 3311 1462 3315 1466
rect 3479 1462 3483 1466
rect 2843 1432 2847 1436
rect 3287 1432 3291 1436
rect 367 1366 371 1370
rect 431 1366 435 1370
rect 487 1366 491 1370
rect 583 1366 587 1370
rect 607 1366 611 1370
rect 727 1366 731 1370
rect 735 1366 739 1370
rect 839 1366 843 1370
rect 879 1366 883 1370
rect 943 1366 947 1370
rect 1023 1366 1027 1370
rect 1047 1366 1051 1370
rect 1151 1366 1155 1370
rect 1167 1366 1171 1370
rect 111 1286 115 1290
rect 135 1286 139 1290
rect 263 1286 267 1290
rect 279 1286 283 1290
rect 423 1286 427 1290
rect 111 1202 115 1206
rect 143 1202 147 1206
rect 575 1286 579 1290
rect 591 1286 595 1290
rect 1871 1386 1875 1390
rect 2255 1386 2259 1390
rect 2263 1386 2267 1390
rect 2335 1386 2339 1390
rect 2343 1386 2347 1390
rect 2415 1386 2419 1390
rect 2423 1386 2427 1390
rect 2495 1386 2499 1390
rect 2503 1386 2507 1390
rect 2591 1386 2595 1390
rect 2599 1386 2603 1390
rect 1263 1366 1267 1370
rect 1319 1366 1323 1370
rect 1471 1366 1475 1370
rect 1623 1366 1627 1370
rect 1831 1366 1835 1370
rect 727 1286 731 1290
rect 759 1286 763 1290
rect 871 1286 875 1290
rect 927 1286 931 1290
rect 1015 1286 1019 1290
rect 1079 1286 1083 1290
rect 1159 1286 1163 1290
rect 1223 1286 1227 1290
rect 1311 1286 1315 1290
rect 271 1202 275 1206
rect 311 1202 315 1206
rect 431 1202 435 1206
rect 487 1202 491 1206
rect 423 1195 427 1196
rect 423 1192 427 1195
rect 599 1202 603 1206
rect 671 1202 675 1206
rect 767 1202 771 1206
rect 847 1202 851 1206
rect 679 1192 683 1196
rect 111 1126 115 1130
rect 135 1126 139 1130
rect 247 1126 251 1130
rect 111 1038 115 1042
rect 143 1038 147 1042
rect 303 1126 307 1130
rect 383 1126 387 1130
rect 479 1126 483 1130
rect 519 1126 523 1130
rect 647 1126 651 1130
rect 663 1126 667 1130
rect 775 1126 779 1130
rect 839 1126 843 1130
rect 1095 1224 1099 1228
rect 935 1202 939 1206
rect 1007 1202 1011 1206
rect 1087 1202 1091 1206
rect 1159 1202 1163 1206
rect 1231 1202 1235 1206
rect 1291 1224 1295 1228
rect 1871 1298 1875 1302
rect 2215 1298 2219 1302
rect 2271 1298 2275 1302
rect 2295 1298 2299 1302
rect 2351 1298 2355 1302
rect 2375 1298 2379 1302
rect 1351 1286 1355 1290
rect 1463 1286 1467 1290
rect 1479 1286 1483 1290
rect 1607 1286 1611 1290
rect 1615 1286 1619 1290
rect 1735 1286 1739 1290
rect 1831 1286 1835 1290
rect 2583 1336 2587 1340
rect 2695 1386 2699 1390
rect 2727 1386 2731 1390
rect 2807 1386 2811 1390
rect 2887 1386 2891 1390
rect 2919 1386 2923 1390
rect 3039 1386 3043 1390
rect 3071 1386 3075 1390
rect 3159 1386 3163 1390
rect 3271 1386 3275 1390
rect 3279 1386 3283 1390
rect 3399 1386 3403 1390
rect 2839 1336 2843 1340
rect 2431 1298 2435 1302
rect 2455 1298 2459 1302
rect 2511 1298 2515 1302
rect 2551 1298 2555 1302
rect 2599 1298 2603 1302
rect 2663 1298 2667 1302
rect 2703 1298 2707 1302
rect 2791 1298 2795 1302
rect 2815 1298 2819 1302
rect 2927 1298 2931 1302
rect 3047 1298 3051 1302
rect 3071 1298 3075 1302
rect 3167 1298 3171 1302
rect 3215 1298 3219 1302
rect 3471 1386 3475 1390
rect 3591 1782 3595 1786
rect 3591 1702 3595 1706
rect 3591 1622 3595 1626
rect 3495 1542 3499 1546
rect 3503 1542 3507 1546
rect 3591 1542 3595 1546
rect 3503 1462 3507 1466
rect 3591 1462 3595 1466
rect 3503 1386 3507 1390
rect 3591 1386 3595 1390
rect 3287 1298 3291 1302
rect 3367 1298 3371 1302
rect 3407 1298 3411 1302
rect 3511 1298 3515 1302
rect 3591 1298 3595 1302
rect 1295 1202 1299 1206
rect 1359 1202 1363 1206
rect 1415 1202 1419 1206
rect 1487 1202 1491 1206
rect 1535 1202 1539 1206
rect 1615 1202 1619 1206
rect 895 1126 899 1130
rect 999 1126 1003 1130
rect 1015 1126 1019 1130
rect 1135 1126 1139 1130
rect 1151 1126 1155 1130
rect 239 1038 243 1042
rect 255 1038 259 1042
rect 359 1038 363 1042
rect 391 1038 395 1042
rect 471 1038 475 1042
rect 527 1038 531 1042
rect 575 1038 579 1042
rect 1255 1126 1259 1130
rect 1287 1126 1291 1130
rect 1375 1126 1379 1130
rect 1407 1126 1411 1130
rect 1503 1126 1507 1130
rect 1527 1126 1531 1130
rect 1655 1202 1659 1206
rect 1743 1202 1747 1206
rect 1751 1202 1755 1206
rect 1871 1218 1875 1222
rect 2111 1218 2115 1222
rect 1831 1202 1835 1206
rect 2207 1218 2211 1222
rect 2287 1218 2291 1222
rect 2303 1218 2307 1222
rect 2367 1218 2371 1222
rect 2407 1218 2411 1222
rect 2447 1218 2451 1222
rect 2527 1218 2531 1222
rect 2543 1218 2547 1222
rect 2647 1218 2651 1222
rect 2655 1218 2659 1222
rect 1871 1134 1875 1138
rect 1903 1134 1907 1138
rect 2119 1134 2123 1138
rect 2127 1134 2131 1138
rect 2215 1134 2219 1138
rect 2311 1134 2315 1138
rect 2359 1134 2363 1138
rect 2415 1134 2419 1138
rect 1631 1126 1635 1130
rect 1647 1126 1651 1130
rect 1743 1126 1747 1130
rect 1831 1126 1835 1130
rect 2583 1160 2587 1164
rect 2535 1134 2539 1138
rect 2575 1134 2579 1138
rect 2775 1218 2779 1222
rect 2783 1218 2787 1222
rect 2911 1218 2915 1222
rect 2919 1218 2923 1222
rect 3055 1218 3059 1222
rect 3063 1218 3067 1222
rect 3199 1218 3203 1222
rect 3207 1218 3211 1222
rect 3343 1218 3347 1222
rect 3359 1218 3363 1222
rect 2999 1160 3003 1164
rect 2655 1134 2659 1138
rect 2775 1134 2779 1138
rect 2783 1134 2787 1138
rect 2919 1134 2923 1138
rect 2967 1134 2971 1138
rect 3063 1134 3067 1138
rect 3159 1134 3163 1138
rect 3207 1134 3211 1138
rect 3495 1218 3499 1222
rect 3503 1218 3507 1222
rect 3591 1218 3595 1222
rect 3343 1134 3347 1138
rect 3351 1134 3355 1138
rect 3503 1134 3507 1138
rect 3511 1134 3515 1138
rect 3591 1134 3595 1138
rect 1871 1058 1875 1062
rect 1895 1058 1899 1062
rect 2015 1058 2019 1062
rect 2119 1058 2123 1062
rect 2167 1058 2171 1062
rect 655 1038 659 1042
rect 671 1038 675 1042
rect 767 1038 771 1042
rect 783 1038 787 1042
rect 855 1038 859 1042
rect 903 1038 907 1042
rect 943 1038 947 1042
rect 1023 1038 1027 1042
rect 1031 1038 1035 1042
rect 1127 1038 1131 1042
rect 1143 1038 1147 1042
rect 1223 1038 1227 1042
rect 1263 1038 1267 1042
rect 1383 1038 1387 1042
rect 1511 1038 1515 1042
rect 1639 1038 1643 1042
rect 1751 1038 1755 1042
rect 1831 1038 1835 1042
rect 111 950 115 954
rect 135 950 139 954
rect 231 950 235 954
rect 263 950 267 954
rect 351 950 355 954
rect 415 950 419 954
rect 463 950 467 954
rect 559 950 563 954
rect 567 950 571 954
rect 663 950 667 954
rect 2327 1058 2331 1062
rect 2351 1058 2355 1062
rect 2487 1058 2491 1062
rect 2567 1058 2571 1062
rect 2639 1058 2643 1062
rect 2767 1058 2771 1062
rect 2791 1058 2795 1062
rect 2935 1058 2939 1062
rect 2959 1058 2963 1062
rect 1871 978 1875 982
rect 1903 978 1907 982
rect 1983 978 1987 982
rect 2023 978 2027 982
rect 2079 978 2083 982
rect 2175 978 2179 982
rect 2199 978 2203 982
rect 703 950 707 954
rect 759 950 763 954
rect 839 950 843 954
rect 847 950 851 954
rect 935 950 939 954
rect 975 950 979 954
rect 1023 950 1027 954
rect 1103 950 1107 954
rect 1119 950 1123 954
rect 1215 950 1219 954
rect 1223 950 1227 954
rect 1335 950 1339 954
rect 1439 950 1443 954
rect 1543 950 1547 954
rect 1655 950 1659 954
rect 1743 950 1747 954
rect 1831 950 1835 954
rect 3079 1058 3083 1062
rect 3151 1058 3155 1062
rect 3223 1058 3227 1062
rect 3335 1058 3339 1062
rect 3375 1058 3379 1062
rect 3503 1058 3507 1062
rect 3591 1058 3595 1062
rect 2335 978 2339 982
rect 2479 978 2483 982
rect 2495 978 2499 982
rect 2631 978 2635 982
rect 2647 978 2651 982
rect 2791 978 2795 982
rect 2799 978 2803 982
rect 2943 978 2947 982
rect 2967 978 2971 982
rect 3087 978 3091 982
rect 3151 978 3155 982
rect 3231 978 3235 982
rect 3343 978 3347 982
rect 3383 978 3387 982
rect 3511 978 3515 982
rect 3591 978 3595 982
rect 111 870 115 874
rect 143 870 147 874
rect 247 870 251 874
rect 271 870 275 874
rect 383 870 387 874
rect 423 870 427 874
rect 519 870 523 874
rect 567 870 571 874
rect 259 840 263 844
rect 111 782 115 786
rect 135 782 139 786
rect 215 782 219 786
rect 239 782 243 786
rect 303 782 307 786
rect 663 870 667 874
rect 711 870 715 874
rect 815 870 819 874
rect 527 840 531 844
rect 847 870 851 874
rect 959 870 963 874
rect 983 870 987 874
rect 1103 870 1107 874
rect 1111 870 1115 874
rect 1231 870 1235 874
rect 1247 870 1251 874
rect 1343 870 1347 874
rect 1383 870 1387 874
rect 1447 870 1451 874
rect 1511 870 1515 874
rect 1551 870 1555 874
rect 1639 870 1643 874
rect 1663 870 1667 874
rect 375 782 379 786
rect 415 782 419 786
rect 511 782 515 786
rect 543 782 547 786
rect 655 782 659 786
rect 687 782 691 786
rect 807 782 811 786
rect 839 782 843 786
rect 951 782 955 786
rect 991 782 995 786
rect 1095 782 1099 786
rect 1143 782 1147 786
rect 151 720 155 724
rect 111 698 115 702
rect 143 698 147 702
rect 223 698 227 702
rect 231 698 235 702
rect 311 698 315 702
rect 319 698 323 702
rect 423 698 427 702
rect 275 680 279 684
rect 655 720 659 724
rect 543 698 547 702
rect 551 698 555 702
rect 679 698 683 702
rect 695 698 699 702
rect 815 698 819 702
rect 847 698 851 702
rect 551 680 555 684
rect 1239 782 1243 786
rect 1295 782 1299 786
rect 1375 782 1379 786
rect 1447 782 1451 786
rect 1503 782 1507 786
rect 1871 890 1875 894
rect 1895 890 1899 894
rect 1919 890 1923 894
rect 1975 890 1979 894
rect 2071 890 2075 894
rect 2095 890 2099 894
rect 2191 890 2195 894
rect 2271 890 2275 894
rect 1751 870 1755 874
rect 1831 870 1835 874
rect 2327 890 2331 894
rect 2455 890 2459 894
rect 2471 890 2475 894
rect 2623 890 2627 894
rect 2655 890 2659 894
rect 2783 890 2787 894
rect 2863 890 2867 894
rect 2959 890 2963 894
rect 3079 890 3083 894
rect 3143 890 3147 894
rect 1871 814 1875 818
rect 1903 814 1907 818
rect 1927 814 1931 818
rect 2015 814 2019 818
rect 2103 814 2107 818
rect 2167 814 2171 818
rect 2279 814 2283 818
rect 2327 814 2331 818
rect 2463 814 2467 818
rect 2487 814 2491 818
rect 2647 814 2651 818
rect 2663 814 2667 818
rect 2807 814 2811 818
rect 2871 814 2875 818
rect 1607 782 1611 786
rect 1631 782 1635 786
rect 1743 782 1747 786
rect 1831 782 1835 786
rect 3303 890 3307 894
rect 3335 890 3339 894
rect 3503 890 3507 894
rect 3591 890 3595 894
rect 2959 814 2963 818
rect 3087 814 3091 818
rect 3103 814 3107 818
rect 3247 814 3251 818
rect 3311 814 3315 818
rect 3391 814 3395 818
rect 3511 814 3515 818
rect 1311 720 1315 724
rect 1531 720 1535 724
rect 951 698 955 702
rect 999 698 1003 702
rect 1087 698 1091 702
rect 1151 698 1155 702
rect 1215 698 1219 702
rect 1303 698 1307 702
rect 1335 698 1339 702
rect 1455 698 1459 702
rect 1583 698 1587 702
rect 111 614 115 618
rect 223 614 227 618
rect 311 614 315 618
rect 415 614 419 618
rect 447 614 451 618
rect 527 614 531 618
rect 535 614 539 618
rect 607 614 611 618
rect 671 614 675 618
rect 687 614 691 618
rect 775 614 779 618
rect 807 614 811 618
rect 1871 738 1875 742
rect 1895 738 1899 742
rect 1967 738 1971 742
rect 2007 738 2011 742
rect 2063 738 2067 742
rect 2159 738 2163 742
rect 2175 738 2179 742
rect 2303 738 2307 742
rect 2319 738 2323 742
rect 2191 712 2195 716
rect 1615 698 1619 702
rect 1831 698 1835 702
rect 1983 672 1987 676
rect 1871 662 1875 666
rect 1975 662 1979 666
rect 2071 662 2075 666
rect 2175 662 2179 666
rect 2183 662 2187 666
rect 1095 624 1099 628
rect 1411 624 1415 628
rect 871 614 875 618
rect 943 614 947 618
rect 959 614 963 618
rect 1047 614 1051 618
rect 1079 614 1083 618
rect 1143 614 1147 618
rect 1207 614 1211 618
rect 1239 614 1243 618
rect 1327 614 1331 618
rect 1335 614 1339 618
rect 2447 738 2451 742
rect 2479 738 2483 742
rect 2599 738 2603 742
rect 2639 738 2643 742
rect 2607 712 2611 716
rect 2419 672 2423 676
rect 2751 738 2755 742
rect 2799 738 2803 742
rect 2271 662 2275 666
rect 2311 662 2315 666
rect 2375 662 2379 666
rect 2455 662 2459 666
rect 2487 662 2491 666
rect 2607 662 2611 666
rect 2735 662 2739 666
rect 2759 662 2763 666
rect 2903 738 2907 742
rect 2951 738 2955 742
rect 3591 814 3595 818
rect 3055 738 3059 742
rect 3095 738 3099 742
rect 3207 738 3211 742
rect 3239 738 3243 742
rect 3359 738 3363 742
rect 2863 662 2867 666
rect 2911 662 2915 666
rect 2991 662 2995 666
rect 3063 662 3067 666
rect 3119 662 3123 666
rect 3215 662 3219 666
rect 3247 662 3251 666
rect 3383 738 3387 742
rect 3503 738 3507 742
rect 3591 738 3595 742
rect 3367 662 3371 666
rect 3375 662 3379 666
rect 3511 662 3515 666
rect 3591 662 3595 666
rect 1431 614 1435 618
rect 1447 614 1451 618
rect 1575 614 1579 618
rect 1831 614 1835 618
rect 1871 586 1875 590
rect 2167 586 2171 590
rect 2263 586 2267 590
rect 2343 586 2347 590
rect 2367 586 2371 590
rect 2423 586 2427 590
rect 2479 586 2483 590
rect 2503 586 2507 590
rect 111 526 115 530
rect 335 526 339 530
rect 423 526 427 530
rect 455 526 459 530
rect 511 526 515 530
rect 535 526 539 530
rect 591 526 595 530
rect 111 442 115 446
rect 223 442 227 446
rect 615 526 619 530
rect 671 526 675 530
rect 695 526 699 530
rect 751 526 755 530
rect 783 526 787 530
rect 839 526 843 530
rect 879 526 883 530
rect 927 526 931 530
rect 967 526 971 530
rect 1015 526 1019 530
rect 1055 526 1059 530
rect 1103 526 1107 530
rect 1151 526 1155 530
rect 1191 526 1195 530
rect 1247 526 1251 530
rect 1279 526 1283 530
rect 327 442 331 446
rect 335 442 339 446
rect 415 442 419 446
rect 447 442 451 446
rect 503 442 507 446
rect 559 442 563 446
rect 583 442 587 446
rect 663 442 667 446
rect 743 442 747 446
rect 759 442 763 446
rect 831 442 835 446
rect 847 442 851 446
rect 2283 544 2287 548
rect 1343 526 1347 530
rect 1439 526 1443 530
rect 1831 526 1835 530
rect 2591 586 2595 590
rect 2599 586 2603 590
rect 2695 586 2699 590
rect 2727 586 2731 590
rect 2539 544 2543 548
rect 1871 502 1875 506
rect 2191 502 2195 506
rect 2271 502 2275 506
rect 2287 502 2291 506
rect 2351 502 2355 506
rect 2383 502 2387 506
rect 2431 502 2435 506
rect 2487 502 2491 506
rect 2511 502 2515 506
rect 2583 502 2587 506
rect 2599 502 2603 506
rect 2687 502 2691 506
rect 2703 502 2707 506
rect 2815 586 2819 590
rect 2855 586 2859 590
rect 2959 586 2963 590
rect 2983 586 2987 590
rect 3111 586 3115 590
rect 3239 586 3243 590
rect 3279 586 3283 590
rect 3367 586 3371 590
rect 3447 586 3451 590
rect 3503 586 3507 590
rect 3591 586 3595 590
rect 2791 502 2795 506
rect 2823 502 2827 506
rect 2911 502 2915 506
rect 2967 502 2971 506
rect 3039 502 3043 506
rect 3119 502 3123 506
rect 3175 502 3179 506
rect 3287 502 3291 506
rect 3319 502 3323 506
rect 3455 502 3459 506
rect 3471 502 3475 506
rect 3591 502 3595 506
rect 919 442 923 446
rect 935 442 939 446
rect 1007 442 1011 446
rect 1023 442 1027 446
rect 1095 442 1099 446
rect 1111 442 1115 446
rect 1183 442 1187 446
rect 1199 442 1203 446
rect 1271 442 1275 446
rect 1295 442 1299 446
rect 1831 442 1835 446
rect 1871 422 1875 426
rect 1975 422 1979 426
rect 111 354 115 358
rect 143 354 147 358
rect 231 354 235 358
rect 263 354 267 358
rect 343 354 347 358
rect 399 354 403 358
rect 455 354 459 358
rect 535 354 539 358
rect 567 354 571 358
rect 671 354 675 358
rect 767 354 771 358
rect 791 354 795 358
rect 855 354 859 358
rect 911 354 915 358
rect 943 354 947 358
rect 1023 354 1027 358
rect 1031 354 1035 358
rect 1119 354 1123 358
rect 1127 354 1131 358
rect 1207 354 1211 358
rect 1231 354 1235 358
rect 1303 354 1307 358
rect 1335 354 1339 358
rect 1439 354 1443 358
rect 1831 354 1835 358
rect 111 270 115 274
rect 135 270 139 274
rect 247 270 251 274
rect 255 270 259 274
rect 391 270 395 274
rect 527 270 531 274
rect 543 270 547 274
rect 663 270 667 274
rect 695 270 699 274
rect 783 270 787 274
rect 111 158 115 162
rect 143 158 147 162
rect 223 158 227 162
rect 255 158 259 162
rect 303 158 307 162
rect 383 158 387 162
rect 399 158 403 162
rect 463 158 467 162
rect 543 158 547 162
rect 551 158 555 162
rect 847 270 851 274
rect 903 270 907 274
rect 991 270 995 274
rect 1015 270 1019 274
rect 1119 270 1123 274
rect 1223 270 1227 274
rect 1239 270 1243 274
rect 2063 422 2067 426
rect 2159 422 2163 426
rect 2183 422 2187 426
rect 2255 422 2259 426
rect 2279 422 2283 426
rect 2359 422 2363 426
rect 2375 422 2379 426
rect 2471 422 2475 426
rect 2479 422 2483 426
rect 2575 422 2579 426
rect 2607 422 2611 426
rect 2679 422 2683 426
rect 2759 422 2763 426
rect 2783 422 2787 426
rect 2903 422 2907 426
rect 2927 422 2931 426
rect 3031 422 3035 426
rect 3111 422 3115 426
rect 3167 422 3171 426
rect 3303 422 3307 426
rect 3311 422 3315 426
rect 3463 422 3467 426
rect 3495 422 3499 426
rect 3591 422 3595 426
rect 1871 342 1875 346
rect 1983 342 1987 346
rect 2071 342 2075 346
rect 2167 342 2171 346
rect 2215 342 2219 346
rect 2263 342 2267 346
rect 2295 342 2299 346
rect 2367 342 2371 346
rect 2383 342 2387 346
rect 2479 342 2483 346
rect 2591 342 2595 346
rect 2615 342 2619 346
rect 2719 342 2723 346
rect 2767 342 2771 346
rect 2847 342 2851 346
rect 2935 342 2939 346
rect 2983 342 2987 346
rect 3119 342 3123 346
rect 3255 342 3259 346
rect 3311 342 3315 346
rect 3391 342 3395 346
rect 1327 270 1331 274
rect 1359 270 1363 274
rect 1431 270 1435 274
rect 1479 270 1483 274
rect 1599 270 1603 274
rect 1831 270 1835 274
rect 1871 262 1875 266
rect 1991 262 1995 266
rect 2119 262 2123 266
rect 2207 262 2211 266
rect 2255 262 2259 266
rect 2287 262 2291 266
rect 2375 262 2379 266
rect 2391 262 2395 266
rect 2471 262 2475 266
rect 2535 262 2539 266
rect 1075 168 1079 172
rect 623 158 627 162
rect 703 158 707 162
rect 783 158 787 162
rect 855 158 859 162
rect 863 158 867 162
rect 943 158 947 162
rect 999 158 1003 162
rect 1023 158 1027 162
rect 1359 168 1363 172
rect 1871 174 1875 178
rect 1903 174 1907 178
rect 1983 174 1987 178
rect 1999 174 2003 178
rect 2087 174 2091 178
rect 2127 174 2131 178
rect 1103 158 1107 162
rect 1127 158 1131 162
rect 1183 158 1187 162
rect 1247 158 1251 162
rect 1263 158 1267 162
rect 1343 158 1347 162
rect 1367 158 1371 162
rect 1423 158 1427 162
rect 1487 158 1491 162
rect 1511 158 1515 162
rect 1591 158 1595 162
rect 1607 158 1611 162
rect 1671 158 1675 162
rect 1751 158 1755 162
rect 1831 158 1835 162
rect 2583 262 2587 266
rect 2679 262 2683 266
rect 2711 262 2715 266
rect 2815 262 2819 266
rect 2839 262 2843 266
rect 2951 262 2955 266
rect 2975 262 2979 266
rect 3095 262 3099 266
rect 3503 342 3507 346
rect 3511 342 3515 346
rect 3591 342 3595 346
rect 3111 262 3115 266
rect 3239 262 3243 266
rect 3247 262 3251 266
rect 3383 262 3387 266
rect 3503 262 3507 266
rect 2215 174 2219 178
rect 2263 174 2267 178
rect 2351 174 2355 178
rect 2399 174 2403 178
rect 2487 174 2491 178
rect 2543 174 2547 178
rect 2623 174 2627 178
rect 2687 174 2691 178
rect 2743 174 2747 178
rect 2823 174 2827 178
rect 2855 174 2859 178
rect 2959 174 2963 178
rect 3063 174 3067 178
rect 3103 174 3107 178
rect 3159 174 3163 178
rect 3247 174 3251 178
rect 3343 174 3347 178
rect 3391 174 3395 178
rect 3431 174 3435 178
rect 3591 262 3595 266
rect 3511 174 3515 178
rect 3591 174 3595 178
rect 1871 98 1875 102
rect 1895 98 1899 102
rect 1975 98 1979 102
rect 2079 98 2083 102
rect 2207 98 2211 102
rect 2343 98 2347 102
rect 2479 98 2483 102
rect 2615 98 2619 102
rect 2735 98 2739 102
rect 2847 98 2851 102
rect 2951 98 2955 102
rect 3055 98 3059 102
rect 3151 98 3155 102
rect 3239 98 3243 102
rect 3335 98 3339 102
rect 3423 98 3427 102
rect 3503 98 3507 102
rect 3591 98 3595 102
rect 111 82 115 86
rect 135 82 139 86
rect 215 82 219 86
rect 295 82 299 86
rect 375 82 379 86
rect 455 82 459 86
rect 535 82 539 86
rect 615 82 619 86
rect 695 82 699 86
rect 775 82 779 86
rect 855 82 859 86
rect 935 82 939 86
rect 1015 82 1019 86
rect 1095 82 1099 86
rect 1175 82 1179 86
rect 1255 82 1259 86
rect 1335 82 1339 86
rect 1415 82 1419 86
rect 1503 82 1507 86
rect 1583 82 1587 86
rect 1663 82 1667 86
rect 1743 82 1747 86
rect 1831 82 1835 86
<< m4 >>
rect 84 3665 85 3671
rect 91 3670 1843 3671
rect 91 3666 111 3670
rect 115 3666 135 3670
rect 139 3666 215 3670
rect 219 3666 295 3670
rect 299 3666 1831 3670
rect 1835 3666 1843 3670
rect 91 3665 1843 3666
rect 1849 3665 1850 3671
rect 1854 3597 1855 3603
rect 1861 3602 3631 3603
rect 1861 3598 1871 3602
rect 1875 3598 2063 3602
rect 2067 3598 2151 3602
rect 2155 3598 2255 3602
rect 2259 3598 2367 3602
rect 2371 3598 2479 3602
rect 2483 3598 2591 3602
rect 2595 3598 2703 3602
rect 2707 3598 2815 3602
rect 2819 3598 2919 3602
rect 2923 3598 3015 3602
rect 3019 3598 3111 3602
rect 3115 3598 3207 3602
rect 3211 3598 3303 3602
rect 3307 3598 3399 3602
rect 3403 3598 3591 3602
rect 3595 3598 3631 3602
rect 1861 3597 3631 3598
rect 3637 3597 3638 3603
rect 1854 3595 1862 3597
rect 96 3589 97 3595
rect 103 3594 1855 3595
rect 103 3590 111 3594
rect 115 3590 143 3594
rect 147 3590 223 3594
rect 227 3590 303 3594
rect 307 3590 343 3594
rect 347 3590 471 3594
rect 475 3590 607 3594
rect 611 3590 743 3594
rect 747 3590 879 3594
rect 883 3590 999 3594
rect 1003 3590 1111 3594
rect 1115 3590 1223 3594
rect 1227 3590 1327 3594
rect 1331 3590 1423 3594
rect 1427 3590 1527 3594
rect 1531 3590 1631 3594
rect 1635 3590 1831 3594
rect 1835 3590 1855 3594
rect 103 3589 1855 3590
rect 1861 3589 1862 3595
rect 1842 3521 1843 3527
rect 1849 3526 3619 3527
rect 1849 3522 1871 3526
rect 1875 3522 2055 3526
rect 2059 3522 2087 3526
rect 2091 3522 2143 3526
rect 2147 3522 2167 3526
rect 2171 3522 2247 3526
rect 2251 3522 2263 3526
rect 2267 3522 2359 3526
rect 2363 3522 2367 3526
rect 2371 3522 2471 3526
rect 2475 3522 2487 3526
rect 2491 3522 2583 3526
rect 2587 3522 2615 3526
rect 2619 3522 2695 3526
rect 2699 3522 2743 3526
rect 2747 3522 2807 3526
rect 2811 3522 2871 3526
rect 2875 3522 2911 3526
rect 2915 3522 2991 3526
rect 2995 3522 3007 3526
rect 3011 3522 3103 3526
rect 3107 3522 3119 3526
rect 3123 3522 3199 3526
rect 3203 3522 3247 3526
rect 3251 3522 3295 3526
rect 3299 3522 3375 3526
rect 3379 3522 3391 3526
rect 3395 3522 3591 3526
rect 3595 3522 3619 3526
rect 1849 3521 3619 3522
rect 3625 3521 3626 3527
rect 1842 3519 1850 3521
rect 84 3513 85 3519
rect 91 3518 1843 3519
rect 91 3514 111 3518
rect 115 3514 135 3518
rect 139 3514 191 3518
rect 195 3514 215 3518
rect 219 3514 327 3518
rect 331 3514 335 3518
rect 339 3514 463 3518
rect 467 3514 471 3518
rect 475 3514 599 3518
rect 603 3514 623 3518
rect 627 3514 735 3518
rect 739 3514 775 3518
rect 779 3514 871 3518
rect 875 3514 919 3518
rect 923 3514 991 3518
rect 995 3514 1055 3518
rect 1059 3514 1103 3518
rect 1107 3514 1183 3518
rect 1187 3514 1215 3518
rect 1219 3514 1311 3518
rect 1315 3514 1319 3518
rect 1323 3514 1415 3518
rect 1419 3514 1439 3518
rect 1443 3514 1519 3518
rect 1523 3514 1567 3518
rect 1571 3514 1623 3518
rect 1627 3514 1831 3518
rect 1835 3514 1843 3518
rect 91 3513 1843 3514
rect 1849 3513 1850 3519
rect 96 3437 97 3443
rect 103 3442 1855 3443
rect 103 3438 111 3442
rect 115 3438 151 3442
rect 155 3438 199 3442
rect 203 3438 295 3442
rect 299 3438 335 3442
rect 339 3438 455 3442
rect 459 3438 479 3442
rect 483 3438 623 3442
rect 627 3438 631 3442
rect 635 3438 783 3442
rect 787 3438 791 3442
rect 795 3438 927 3442
rect 931 3438 959 3442
rect 963 3438 1063 3442
rect 1067 3438 1119 3442
rect 1123 3438 1191 3442
rect 1195 3438 1271 3442
rect 1275 3438 1319 3442
rect 1323 3438 1415 3442
rect 1419 3438 1447 3442
rect 1451 3438 1559 3442
rect 1563 3438 1575 3442
rect 1579 3438 1711 3442
rect 1715 3438 1831 3442
rect 1835 3438 1855 3442
rect 103 3437 1855 3438
rect 1861 3442 3638 3443
rect 1861 3438 1871 3442
rect 1875 3438 2095 3442
rect 2099 3438 2111 3442
rect 2115 3438 2175 3442
rect 2179 3438 2199 3442
rect 2203 3438 2271 3442
rect 2275 3438 2303 3442
rect 2307 3438 2375 3442
rect 2379 3438 2415 3442
rect 2419 3438 2495 3442
rect 2499 3438 2543 3442
rect 2547 3438 2623 3442
rect 2627 3438 2679 3442
rect 2683 3438 2751 3442
rect 2755 3438 2815 3442
rect 2819 3438 2879 3442
rect 2883 3438 2959 3442
rect 2963 3438 2999 3442
rect 3003 3438 3111 3442
rect 3115 3438 3127 3442
rect 3131 3438 3255 3442
rect 3259 3438 3263 3442
rect 3267 3438 3383 3442
rect 3387 3438 3423 3442
rect 3427 3438 3591 3442
rect 3595 3438 3638 3442
rect 1861 3437 3638 3438
rect 84 3361 85 3367
rect 91 3366 1843 3367
rect 91 3362 111 3366
rect 115 3362 143 3366
rect 147 3362 207 3366
rect 211 3362 287 3366
rect 291 3362 335 3366
rect 339 3362 447 3366
rect 451 3362 471 3366
rect 475 3362 615 3366
rect 619 3362 623 3366
rect 627 3362 783 3366
rect 787 3362 943 3366
rect 947 3362 951 3366
rect 955 3362 1103 3366
rect 1107 3362 1111 3366
rect 1115 3362 1263 3366
rect 1267 3362 1407 3366
rect 1411 3362 1423 3366
rect 1427 3362 1551 3366
rect 1555 3362 1583 3366
rect 1587 3362 1703 3366
rect 1707 3362 1743 3366
rect 1747 3362 1831 3366
rect 1835 3362 1843 3366
rect 91 3361 1843 3362
rect 1849 3363 1850 3367
rect 1849 3362 3626 3363
rect 1849 3361 1871 3362
rect 1842 3358 1871 3361
rect 1875 3358 2103 3362
rect 2107 3358 2127 3362
rect 2131 3358 2191 3362
rect 2195 3358 2223 3362
rect 2227 3358 2295 3362
rect 2299 3358 2335 3362
rect 2339 3358 2407 3362
rect 2411 3358 2455 3362
rect 2459 3358 2535 3362
rect 2539 3358 2583 3362
rect 2587 3358 2671 3362
rect 2675 3358 2719 3362
rect 2723 3358 2807 3362
rect 2811 3358 2863 3362
rect 2867 3358 2951 3362
rect 2955 3358 3007 3362
rect 3011 3358 3103 3362
rect 3107 3358 3159 3362
rect 3163 3358 3255 3362
rect 3259 3358 3311 3362
rect 3315 3358 3415 3362
rect 3419 3358 3471 3362
rect 3475 3358 3591 3362
rect 3595 3358 3626 3362
rect 1842 3357 3626 3358
rect 222 3300 228 3301
rect 678 3300 684 3301
rect 222 3296 223 3300
rect 227 3296 679 3300
rect 683 3296 684 3300
rect 222 3295 228 3296
rect 678 3295 684 3296
rect 96 3281 97 3287
rect 103 3286 1855 3287
rect 103 3282 111 3286
rect 115 3282 215 3286
rect 219 3282 343 3286
rect 347 3282 351 3286
rect 355 3282 455 3286
rect 459 3282 479 3286
rect 483 3282 575 3286
rect 579 3282 631 3286
rect 635 3282 703 3286
rect 707 3282 791 3286
rect 795 3282 839 3286
rect 843 3282 951 3286
rect 955 3282 983 3286
rect 987 3282 1111 3286
rect 1115 3282 1119 3286
rect 1123 3282 1255 3286
rect 1259 3282 1271 3286
rect 1275 3282 1383 3286
rect 1387 3282 1431 3286
rect 1435 3282 1511 3286
rect 1515 3282 1591 3286
rect 1595 3282 1639 3286
rect 1643 3282 1751 3286
rect 1755 3282 1831 3286
rect 1835 3282 1855 3286
rect 103 3281 1855 3282
rect 1861 3281 1862 3287
rect 1854 3269 1855 3275
rect 1861 3274 3631 3275
rect 1861 3270 1871 3274
rect 1875 3270 2135 3274
rect 2139 3270 2231 3274
rect 2235 3270 2279 3274
rect 2283 3270 2343 3274
rect 2347 3270 2415 3274
rect 2419 3270 2463 3274
rect 2467 3270 2551 3274
rect 2555 3270 2591 3274
rect 2595 3270 2687 3274
rect 2691 3270 2727 3274
rect 2731 3270 2823 3274
rect 2827 3270 2871 3274
rect 2875 3270 2959 3274
rect 2963 3270 3015 3274
rect 3019 3270 3095 3274
rect 3099 3270 3167 3274
rect 3171 3270 3231 3274
rect 3235 3270 3319 3274
rect 3323 3270 3375 3274
rect 3379 3270 3479 3274
rect 3483 3270 3511 3274
rect 3515 3270 3591 3274
rect 3595 3270 3631 3274
rect 1861 3269 3631 3270
rect 3637 3269 3638 3275
rect 84 3205 85 3211
rect 91 3210 1843 3211
rect 91 3206 111 3210
rect 115 3206 343 3210
rect 347 3206 447 3210
rect 451 3206 487 3210
rect 491 3206 567 3210
rect 571 3206 575 3210
rect 579 3206 663 3210
rect 667 3206 695 3210
rect 699 3206 767 3210
rect 771 3206 831 3210
rect 835 3206 887 3210
rect 891 3206 975 3210
rect 979 3206 1023 3210
rect 1027 3206 1111 3210
rect 1115 3206 1191 3210
rect 1195 3206 1247 3210
rect 1251 3206 1375 3210
rect 1379 3206 1503 3210
rect 1507 3206 1567 3210
rect 1571 3206 1631 3210
rect 1635 3206 1743 3210
rect 1747 3206 1831 3210
rect 1835 3206 1843 3210
rect 91 3205 1843 3206
rect 1849 3205 1850 3211
rect 1842 3189 1843 3195
rect 1849 3194 3619 3195
rect 1849 3190 1871 3194
rect 1875 3190 1895 3194
rect 1899 3190 1991 3194
rect 1995 3190 2119 3194
rect 2123 3190 2127 3194
rect 2131 3190 2247 3194
rect 2251 3190 2271 3194
rect 2275 3190 2383 3194
rect 2387 3190 2407 3194
rect 2411 3190 2511 3194
rect 2515 3190 2543 3194
rect 2547 3190 2639 3194
rect 2643 3190 2679 3194
rect 2683 3190 2767 3194
rect 2771 3190 2815 3194
rect 2819 3190 2895 3194
rect 2899 3190 2951 3194
rect 2955 3190 3031 3194
rect 3035 3190 3087 3194
rect 3091 3190 3175 3194
rect 3179 3190 3223 3194
rect 3227 3190 3327 3194
rect 3331 3190 3367 3194
rect 3371 3190 3487 3194
rect 3491 3190 3503 3194
rect 3507 3190 3591 3194
rect 3595 3190 3619 3194
rect 1849 3189 3619 3190
rect 3625 3189 3626 3195
rect 634 3148 640 3149
rect 842 3148 848 3149
rect 634 3144 635 3148
rect 639 3144 843 3148
rect 847 3144 848 3148
rect 634 3143 640 3144
rect 842 3143 848 3144
rect 1206 3148 1212 3149
rect 1486 3148 1492 3149
rect 1206 3144 1207 3148
rect 1211 3144 1487 3148
rect 1491 3144 1492 3148
rect 1206 3143 1212 3144
rect 1486 3143 1492 3144
rect 96 3125 97 3131
rect 103 3130 1855 3131
rect 103 3126 111 3130
rect 115 3126 495 3130
rect 499 3126 583 3130
rect 587 3126 591 3130
rect 595 3126 671 3130
rect 675 3126 759 3130
rect 763 3126 775 3130
rect 779 3126 847 3130
rect 851 3126 895 3130
rect 899 3126 935 3130
rect 939 3126 1023 3130
rect 1027 3126 1031 3130
rect 1035 3126 1111 3130
rect 1115 3126 1199 3130
rect 1203 3126 1287 3130
rect 1291 3126 1375 3130
rect 1379 3126 1383 3130
rect 1387 3126 1575 3130
rect 1579 3126 1751 3130
rect 1755 3126 1831 3130
rect 1835 3126 1855 3130
rect 103 3125 1855 3126
rect 1861 3125 1862 3131
rect 1854 3097 1855 3103
rect 1861 3102 3631 3103
rect 1861 3098 1871 3102
rect 1875 3098 1903 3102
rect 1907 3098 1999 3102
rect 2003 3098 2015 3102
rect 2019 3098 2127 3102
rect 2131 3098 2191 3102
rect 2195 3098 2255 3102
rect 2259 3098 2391 3102
rect 2395 3098 2407 3102
rect 2411 3098 2519 3102
rect 2523 3098 2647 3102
rect 2651 3098 2655 3102
rect 2659 3098 2775 3102
rect 2779 3098 2903 3102
rect 2907 3098 2935 3102
rect 2939 3098 3039 3102
rect 3043 3098 3183 3102
rect 3187 3098 3231 3102
rect 3235 3098 3335 3102
rect 3339 3098 3495 3102
rect 3499 3098 3511 3102
rect 3515 3098 3591 3102
rect 3595 3098 3631 3102
rect 1861 3097 3631 3098
rect 3637 3097 3638 3103
rect 1910 3092 1916 3093
rect 2198 3092 2204 3093
rect 1910 3088 1911 3092
rect 1915 3088 2199 3092
rect 2203 3088 2204 3092
rect 1910 3087 1916 3088
rect 2198 3087 2204 3088
rect 2414 3092 2420 3093
rect 2942 3092 2948 3093
rect 2414 3088 2415 3092
rect 2419 3088 2943 3092
rect 2947 3088 2948 3092
rect 2414 3087 2420 3088
rect 2942 3087 2948 3088
rect 84 3045 85 3051
rect 91 3050 1843 3051
rect 91 3046 111 3050
rect 115 3046 543 3050
rect 547 3046 583 3050
rect 587 3046 623 3050
rect 627 3046 663 3050
rect 667 3046 711 3050
rect 715 3046 751 3050
rect 755 3046 807 3050
rect 811 3046 839 3050
rect 843 3046 903 3050
rect 907 3046 927 3050
rect 931 3046 999 3050
rect 1003 3046 1015 3050
rect 1019 3046 1087 3050
rect 1091 3046 1103 3050
rect 1107 3046 1183 3050
rect 1187 3046 1191 3050
rect 1195 3046 1279 3050
rect 1283 3046 1367 3050
rect 1371 3046 1375 3050
rect 1379 3046 1471 3050
rect 1475 3046 1831 3050
rect 1835 3046 1843 3050
rect 91 3045 1843 3046
rect 1849 3045 1850 3051
rect 1842 3013 1843 3019
rect 1849 3018 3619 3019
rect 1849 3014 1871 3018
rect 1875 3014 1895 3018
rect 1899 3014 2007 3018
rect 2011 3014 2047 3018
rect 2051 3014 2183 3018
rect 2187 3014 2223 3018
rect 2227 3014 2391 3018
rect 2395 3014 2399 3018
rect 2403 3014 2543 3018
rect 2547 3014 2647 3018
rect 2651 3014 2687 3018
rect 2691 3014 2815 3018
rect 2819 3014 2927 3018
rect 2931 3014 3039 3018
rect 3043 3014 3143 3018
rect 3147 3014 3223 3018
rect 3227 3014 3239 3018
rect 3243 3014 3335 3018
rect 3339 3014 3423 3018
rect 3427 3014 3503 3018
rect 3507 3014 3591 3018
rect 3595 3014 3619 3018
rect 1849 3013 3619 3014
rect 3625 3013 3626 3019
rect 96 2969 97 2975
rect 103 2974 1855 2975
rect 103 2970 111 2974
rect 115 2970 471 2974
rect 475 2970 551 2974
rect 555 2970 575 2974
rect 579 2970 631 2974
rect 635 2970 687 2974
rect 691 2970 719 2974
rect 723 2970 807 2974
rect 811 2970 815 2974
rect 819 2970 911 2974
rect 915 2970 943 2974
rect 947 2970 1007 2974
rect 1011 2970 1087 2974
rect 1091 2970 1095 2974
rect 1099 2970 1191 2974
rect 1195 2970 1247 2974
rect 1251 2970 1287 2974
rect 1291 2970 1383 2974
rect 1387 2970 1415 2974
rect 1419 2970 1479 2974
rect 1483 2970 1591 2974
rect 1595 2970 1751 2974
rect 1755 2970 1831 2974
rect 1835 2970 1855 2974
rect 103 2969 1855 2970
rect 1861 2969 1862 2975
rect 2566 2956 2572 2957
rect 2918 2956 2924 2957
rect 2566 2952 2567 2956
rect 2571 2952 2919 2956
rect 2923 2952 2924 2956
rect 2566 2951 2572 2952
rect 2918 2951 2924 2952
rect 654 2948 660 2949
rect 950 2948 956 2949
rect 654 2944 655 2948
rect 659 2944 951 2948
rect 955 2944 956 2948
rect 654 2943 660 2944
rect 950 2943 956 2944
rect 1102 2948 1108 2949
rect 1306 2948 1312 2949
rect 1102 2944 1103 2948
rect 1107 2944 1307 2948
rect 1311 2944 1312 2948
rect 1102 2943 1108 2944
rect 1306 2943 1312 2944
rect 1854 2937 1855 2943
rect 1861 2942 3631 2943
rect 1861 2938 1871 2942
rect 1875 2938 1903 2942
rect 1907 2938 2055 2942
rect 2059 2938 2087 2942
rect 2091 2938 2231 2942
rect 2235 2938 2295 2942
rect 2299 2938 2399 2942
rect 2403 2938 2487 2942
rect 2491 2938 2551 2942
rect 2555 2938 2671 2942
rect 2675 2938 2695 2942
rect 2699 2938 2823 2942
rect 2827 2938 2839 2942
rect 2843 2938 2935 2942
rect 2939 2938 2999 2942
rect 3003 2938 3047 2942
rect 3051 2938 3151 2942
rect 3155 2938 3247 2942
rect 3251 2938 3303 2942
rect 3307 2938 3343 2942
rect 3347 2938 3431 2942
rect 3435 2938 3455 2942
rect 3459 2938 3511 2942
rect 3515 2938 3591 2942
rect 3595 2938 3631 2942
rect 1861 2937 3631 2938
rect 3637 2937 3638 2943
rect 2714 2932 2720 2933
rect 3310 2932 3316 2933
rect 2714 2928 2715 2932
rect 2719 2928 3311 2932
rect 3315 2928 3316 2932
rect 2714 2927 2720 2928
rect 3310 2927 3316 2928
rect 84 2893 85 2899
rect 91 2898 1843 2899
rect 91 2894 111 2898
rect 115 2894 311 2898
rect 315 2894 431 2898
rect 435 2894 463 2898
rect 467 2894 551 2898
rect 555 2894 567 2898
rect 571 2894 679 2898
rect 683 2894 799 2898
rect 803 2894 815 2898
rect 819 2894 935 2898
rect 939 2894 951 2898
rect 955 2894 1079 2898
rect 1083 2894 1087 2898
rect 1091 2894 1223 2898
rect 1227 2894 1239 2898
rect 1243 2894 1359 2898
rect 1363 2894 1407 2898
rect 1411 2894 1495 2898
rect 1499 2894 1583 2898
rect 1587 2894 1631 2898
rect 1635 2894 1743 2898
rect 1747 2894 1831 2898
rect 1835 2894 1843 2898
rect 91 2893 1843 2894
rect 1849 2893 1850 2899
rect 1842 2853 1843 2859
rect 1849 2858 3619 2859
rect 1849 2854 1871 2858
rect 1875 2854 1895 2858
rect 1899 2854 2079 2858
rect 2083 2854 2135 2858
rect 2139 2854 2263 2858
rect 2267 2854 2287 2858
rect 2291 2854 2391 2858
rect 2395 2854 2479 2858
rect 2483 2854 2519 2858
rect 2523 2854 2647 2858
rect 2651 2854 2663 2858
rect 2667 2854 2767 2858
rect 2771 2854 2831 2858
rect 2835 2854 2887 2858
rect 2891 2854 2991 2858
rect 2995 2854 3007 2858
rect 3011 2854 3135 2858
rect 3139 2854 3143 2858
rect 3147 2854 3295 2858
rect 3299 2854 3447 2858
rect 3451 2854 3591 2858
rect 3595 2854 3619 2858
rect 1849 2853 3619 2854
rect 3625 2853 3626 2859
rect 326 2836 332 2837
rect 762 2836 768 2837
rect 326 2832 327 2836
rect 331 2832 763 2836
rect 767 2832 768 2836
rect 326 2831 332 2832
rect 762 2831 768 2832
rect 96 2817 97 2823
rect 103 2822 1855 2823
rect 103 2818 111 2822
rect 115 2818 167 2822
rect 171 2818 303 2822
rect 307 2818 319 2822
rect 323 2818 439 2822
rect 443 2818 447 2822
rect 451 2818 559 2822
rect 563 2818 607 2822
rect 611 2818 687 2822
rect 691 2818 783 2822
rect 787 2818 823 2822
rect 827 2818 959 2822
rect 963 2818 1095 2822
rect 1099 2818 1143 2822
rect 1147 2818 1231 2822
rect 1235 2818 1335 2822
rect 1339 2818 1367 2822
rect 1371 2818 1503 2822
rect 1507 2818 1535 2822
rect 1539 2818 1639 2822
rect 1643 2818 1735 2822
rect 1739 2818 1751 2822
rect 1755 2818 1831 2822
rect 1835 2818 1855 2822
rect 103 2817 1855 2818
rect 1861 2817 1862 2823
rect 2662 2804 2668 2805
rect 3086 2804 3092 2805
rect 2662 2800 2663 2804
rect 2667 2800 3087 2804
rect 3091 2800 3092 2804
rect 2662 2799 2668 2800
rect 3086 2799 3092 2800
rect 1854 2769 1855 2775
rect 1861 2774 3631 2775
rect 1861 2770 1871 2774
rect 1875 2770 2143 2774
rect 2147 2770 2231 2774
rect 2235 2770 2271 2774
rect 2275 2770 2311 2774
rect 2315 2770 2391 2774
rect 2395 2770 2399 2774
rect 2403 2770 2471 2774
rect 2475 2770 2527 2774
rect 2531 2770 2551 2774
rect 2555 2770 2639 2774
rect 2643 2770 2655 2774
rect 2659 2770 2727 2774
rect 2731 2770 2775 2774
rect 2779 2770 2815 2774
rect 2819 2770 2895 2774
rect 2899 2770 2903 2774
rect 2907 2770 2991 2774
rect 2995 2770 3015 2774
rect 3019 2770 3143 2774
rect 3147 2770 3591 2774
rect 3595 2770 3631 2774
rect 1861 2769 3631 2770
rect 3637 2769 3638 2775
rect 2646 2764 2652 2765
rect 2998 2764 3004 2765
rect 2646 2760 2647 2764
rect 2651 2760 2999 2764
rect 3003 2760 3004 2764
rect 2646 2759 2652 2760
rect 2998 2759 3004 2760
rect 84 2737 85 2743
rect 91 2742 1843 2743
rect 91 2738 111 2742
rect 115 2738 135 2742
rect 139 2738 159 2742
rect 163 2738 247 2742
rect 251 2738 295 2742
rect 299 2738 391 2742
rect 395 2738 439 2742
rect 443 2738 551 2742
rect 555 2738 599 2742
rect 603 2738 711 2742
rect 715 2738 775 2742
rect 779 2738 879 2742
rect 883 2738 951 2742
rect 955 2738 1039 2742
rect 1043 2738 1135 2742
rect 1139 2738 1199 2742
rect 1203 2738 1327 2742
rect 1331 2738 1359 2742
rect 1363 2738 1519 2742
rect 1523 2738 1527 2742
rect 1531 2738 1687 2742
rect 1691 2738 1727 2742
rect 1731 2738 1831 2742
rect 1835 2738 1843 2742
rect 91 2737 1843 2738
rect 1849 2737 1850 2743
rect 1842 2693 1843 2699
rect 1849 2698 3619 2699
rect 1849 2694 1871 2698
rect 1875 2694 2223 2698
rect 2227 2694 2239 2698
rect 2243 2694 2303 2698
rect 2307 2694 2319 2698
rect 2323 2694 2383 2698
rect 2387 2694 2399 2698
rect 2403 2694 2463 2698
rect 2467 2694 2479 2698
rect 2483 2694 2543 2698
rect 2547 2694 2559 2698
rect 2563 2694 2631 2698
rect 2635 2694 2639 2698
rect 2643 2694 2719 2698
rect 2723 2694 2799 2698
rect 2803 2694 2807 2698
rect 2811 2694 2879 2698
rect 2883 2694 2895 2698
rect 2899 2694 2959 2698
rect 2963 2694 2983 2698
rect 2987 2694 3591 2698
rect 3595 2694 3619 2698
rect 1849 2693 3619 2694
rect 3625 2693 3626 2699
rect 262 2676 268 2677
rect 650 2676 656 2677
rect 262 2672 263 2676
rect 267 2672 651 2676
rect 655 2672 656 2676
rect 262 2671 268 2672
rect 650 2671 656 2672
rect 96 2661 97 2667
rect 103 2666 1855 2667
rect 103 2662 111 2666
rect 115 2662 143 2666
rect 147 2662 255 2666
rect 259 2662 399 2666
rect 403 2662 551 2666
rect 555 2662 559 2666
rect 563 2662 711 2666
rect 715 2662 719 2666
rect 723 2662 879 2666
rect 883 2662 887 2666
rect 891 2662 1047 2666
rect 1051 2662 1207 2666
rect 1211 2662 1215 2666
rect 1219 2662 1367 2666
rect 1371 2662 1391 2666
rect 1395 2662 1527 2666
rect 1531 2662 1567 2666
rect 1571 2662 1695 2666
rect 1699 2662 1831 2666
rect 1835 2662 1855 2666
rect 103 2661 1855 2662
rect 1861 2661 1862 2667
rect 1854 2609 1855 2615
rect 1861 2614 3631 2615
rect 1861 2610 1871 2614
rect 1875 2610 2191 2614
rect 2195 2610 2247 2614
rect 2251 2610 2271 2614
rect 2275 2610 2327 2614
rect 2331 2610 2351 2614
rect 2355 2610 2407 2614
rect 2411 2610 2431 2614
rect 2435 2610 2487 2614
rect 2491 2610 2511 2614
rect 2515 2610 2567 2614
rect 2571 2610 2591 2614
rect 2595 2610 2647 2614
rect 2651 2610 2671 2614
rect 2675 2610 2727 2614
rect 2731 2610 2751 2614
rect 2755 2610 2807 2614
rect 2811 2610 2831 2614
rect 2835 2610 2887 2614
rect 2891 2610 2911 2614
rect 2915 2610 2967 2614
rect 2971 2610 2991 2614
rect 2995 2610 3591 2614
rect 3595 2610 3631 2614
rect 1861 2609 3631 2610
rect 3637 2609 3638 2615
rect 84 2581 85 2587
rect 91 2586 1843 2587
rect 91 2582 111 2586
rect 115 2582 135 2586
rect 139 2582 159 2586
rect 163 2582 247 2586
rect 251 2582 279 2586
rect 283 2582 391 2586
rect 395 2582 415 2586
rect 419 2582 543 2586
rect 547 2582 559 2586
rect 563 2582 703 2586
rect 707 2582 847 2586
rect 851 2582 871 2586
rect 875 2582 983 2586
rect 987 2582 1039 2586
rect 1043 2582 1119 2586
rect 1123 2582 1207 2586
rect 1211 2582 1255 2586
rect 1259 2582 1383 2586
rect 1387 2582 1391 2586
rect 1395 2582 1527 2586
rect 1531 2582 1559 2586
rect 1563 2582 1831 2586
rect 1835 2582 1843 2586
rect 91 2581 1843 2582
rect 1849 2581 1850 2587
rect 174 2556 180 2557
rect 642 2556 648 2557
rect 174 2552 175 2556
rect 179 2552 643 2556
rect 647 2552 648 2556
rect 174 2551 180 2552
rect 642 2551 648 2552
rect 1842 2525 1843 2531
rect 1849 2530 3619 2531
rect 1849 2526 1871 2530
rect 1875 2526 2119 2530
rect 2123 2526 2183 2530
rect 2187 2526 2207 2530
rect 2211 2526 2263 2530
rect 2267 2526 2303 2530
rect 2307 2526 2343 2530
rect 2347 2526 2399 2530
rect 2403 2526 2423 2530
rect 2427 2526 2495 2530
rect 2499 2526 2503 2530
rect 2507 2526 2583 2530
rect 2587 2526 2591 2530
rect 2595 2526 2663 2530
rect 2667 2526 2687 2530
rect 2691 2526 2743 2530
rect 2747 2526 2783 2530
rect 2787 2526 2823 2530
rect 2827 2526 2879 2530
rect 2883 2526 2903 2530
rect 2907 2526 2975 2530
rect 2979 2526 2983 2530
rect 2987 2526 3079 2530
rect 3083 2526 3591 2530
rect 3595 2526 3619 2530
rect 1849 2525 3619 2526
rect 3625 2525 3626 2531
rect 354 2524 360 2525
rect 666 2524 672 2525
rect 354 2520 355 2524
rect 359 2520 667 2524
rect 671 2520 672 2524
rect 354 2519 360 2520
rect 666 2519 672 2520
rect 96 2501 97 2507
rect 103 2506 1855 2507
rect 103 2502 111 2506
rect 115 2502 167 2506
rect 171 2502 287 2506
rect 291 2502 335 2506
rect 339 2502 415 2506
rect 419 2502 423 2506
rect 427 2502 503 2506
rect 507 2502 567 2506
rect 571 2502 599 2506
rect 603 2502 703 2506
rect 707 2502 711 2506
rect 715 2502 815 2506
rect 819 2502 855 2506
rect 859 2502 935 2506
rect 939 2502 991 2506
rect 995 2502 1063 2506
rect 1067 2502 1127 2506
rect 1131 2502 1191 2506
rect 1195 2502 1263 2506
rect 1267 2502 1327 2506
rect 1331 2502 1399 2506
rect 1403 2502 1471 2506
rect 1475 2502 1535 2506
rect 1539 2502 1831 2506
rect 1835 2502 1855 2506
rect 103 2501 1855 2502
rect 1861 2501 1862 2507
rect 2702 2468 2708 2469
rect 3050 2468 3056 2469
rect 2702 2464 2703 2468
rect 2707 2464 3051 2468
rect 3055 2464 3056 2468
rect 2702 2463 2708 2464
rect 3050 2463 3056 2464
rect 1854 2445 1855 2451
rect 1861 2450 3631 2451
rect 1861 2446 1871 2450
rect 1875 2446 1903 2450
rect 1907 2446 1991 2450
rect 1995 2446 2111 2450
rect 2115 2446 2127 2450
rect 2131 2446 2215 2450
rect 2219 2446 2247 2450
rect 2251 2446 2311 2450
rect 2315 2446 2391 2450
rect 2395 2446 2407 2450
rect 2411 2446 2503 2450
rect 2507 2446 2535 2450
rect 2539 2446 2599 2450
rect 2603 2446 2671 2450
rect 2675 2446 2695 2450
rect 2699 2446 2791 2450
rect 2795 2446 2807 2450
rect 2811 2446 2887 2450
rect 2891 2446 2943 2450
rect 2947 2446 2983 2450
rect 2987 2446 3079 2450
rect 3083 2446 3087 2450
rect 3091 2446 3215 2450
rect 3219 2446 3591 2450
rect 3595 2446 3631 2450
rect 1861 2445 3631 2446
rect 3637 2445 3638 2451
rect 2178 2436 2184 2437
rect 2542 2436 2548 2437
rect 2178 2432 2179 2436
rect 2183 2432 2543 2436
rect 2547 2432 2548 2436
rect 2178 2431 2184 2432
rect 2542 2431 2548 2432
rect 84 2417 85 2423
rect 91 2422 1843 2423
rect 91 2418 111 2422
rect 115 2418 327 2422
rect 331 2418 383 2422
rect 387 2418 407 2422
rect 411 2418 463 2422
rect 467 2418 495 2422
rect 499 2418 543 2422
rect 547 2418 591 2422
rect 595 2418 623 2422
rect 627 2418 695 2422
rect 699 2418 703 2422
rect 707 2418 783 2422
rect 787 2418 807 2422
rect 811 2418 863 2422
rect 867 2418 927 2422
rect 931 2418 943 2422
rect 947 2418 1023 2422
rect 1027 2418 1055 2422
rect 1059 2418 1103 2422
rect 1107 2418 1183 2422
rect 1187 2418 1263 2422
rect 1267 2418 1319 2422
rect 1323 2418 1351 2422
rect 1355 2418 1439 2422
rect 1443 2418 1463 2422
rect 1467 2418 1527 2422
rect 1531 2418 1831 2422
rect 1835 2418 1843 2422
rect 91 2417 1843 2418
rect 1849 2417 1850 2423
rect 1946 2412 1952 2413
rect 2458 2412 2464 2413
rect 1946 2408 1947 2412
rect 1951 2408 2459 2412
rect 2463 2408 2464 2412
rect 1946 2407 1952 2408
rect 2458 2407 2464 2408
rect 1842 2361 1843 2367
rect 1849 2366 3619 2367
rect 1849 2362 1871 2366
rect 1875 2362 1895 2366
rect 1899 2362 1983 2366
rect 1987 2362 2015 2366
rect 2019 2362 2103 2366
rect 2107 2362 2175 2366
rect 2179 2362 2239 2366
rect 2243 2362 2343 2366
rect 2347 2362 2383 2366
rect 2387 2362 2511 2366
rect 2515 2362 2527 2366
rect 2531 2362 2663 2366
rect 2667 2362 2671 2366
rect 2675 2362 2799 2366
rect 2803 2362 2823 2366
rect 2827 2362 2935 2366
rect 2939 2362 2959 2366
rect 2963 2362 3071 2366
rect 3075 2362 3079 2366
rect 3083 2362 3191 2366
rect 3195 2362 3207 2366
rect 3211 2362 3303 2366
rect 3307 2362 3415 2366
rect 3419 2362 3503 2366
rect 3507 2362 3591 2366
rect 3595 2362 3619 2366
rect 1849 2361 3619 2362
rect 3625 2361 3626 2367
rect 96 2341 97 2347
rect 103 2346 1855 2347
rect 103 2342 111 2346
rect 115 2342 391 2346
rect 395 2342 471 2346
rect 475 2342 551 2346
rect 555 2342 631 2346
rect 635 2342 711 2346
rect 715 2342 791 2346
rect 795 2342 871 2346
rect 875 2342 951 2346
rect 955 2342 1031 2346
rect 1035 2342 1111 2346
rect 1115 2342 1191 2346
rect 1195 2342 1271 2346
rect 1275 2342 1359 2346
rect 1363 2342 1407 2346
rect 1411 2342 1447 2346
rect 1451 2342 1487 2346
rect 1491 2342 1535 2346
rect 1539 2342 1567 2346
rect 1571 2342 1647 2346
rect 1651 2342 1831 2346
rect 1835 2342 1855 2346
rect 103 2341 1855 2342
rect 1861 2341 1862 2347
rect 2686 2300 2692 2301
rect 3138 2300 3144 2301
rect 2686 2296 2687 2300
rect 2691 2296 3139 2300
rect 3143 2296 3144 2300
rect 2686 2295 2692 2296
rect 3138 2295 3144 2296
rect 1854 2285 1855 2291
rect 1861 2290 3631 2291
rect 1861 2286 1871 2290
rect 1875 2286 1903 2290
rect 1907 2286 2023 2290
rect 2027 2286 2031 2290
rect 2035 2286 2183 2290
rect 2187 2286 2351 2290
rect 2355 2286 2367 2290
rect 2371 2286 2519 2290
rect 2523 2286 2575 2290
rect 2579 2286 2679 2290
rect 2683 2286 2791 2290
rect 2795 2286 2831 2290
rect 2835 2286 2967 2290
rect 2971 2286 3023 2290
rect 3027 2286 3087 2290
rect 3091 2286 3199 2290
rect 3203 2286 3255 2290
rect 3259 2286 3311 2290
rect 3315 2286 3423 2290
rect 3427 2286 3495 2290
rect 3499 2286 3511 2290
rect 3515 2286 3591 2290
rect 3595 2286 3631 2290
rect 1861 2285 3631 2286
rect 3637 2285 3638 2291
rect 84 2257 85 2263
rect 91 2262 1843 2263
rect 91 2258 111 2262
rect 115 2258 135 2262
rect 139 2258 215 2262
rect 219 2258 295 2262
rect 299 2258 383 2262
rect 387 2258 519 2262
rect 523 2258 671 2262
rect 675 2258 831 2262
rect 835 2258 999 2262
rect 1003 2258 1159 2262
rect 1163 2258 1311 2262
rect 1315 2258 1399 2262
rect 1403 2258 1455 2262
rect 1459 2258 1479 2262
rect 1483 2258 1559 2262
rect 1563 2258 1607 2262
rect 1611 2258 1639 2262
rect 1643 2258 1743 2262
rect 1747 2258 1831 2262
rect 1835 2258 1843 2262
rect 91 2257 1843 2258
rect 1849 2257 1850 2263
rect 1174 2244 1180 2245
rect 1578 2244 1584 2245
rect 1174 2240 1175 2244
rect 1179 2240 1579 2244
rect 1583 2240 1584 2244
rect 1174 2239 1180 2240
rect 1578 2239 1584 2240
rect 1206 2196 1212 2197
rect 1690 2196 1696 2197
rect 1206 2192 1207 2196
rect 1211 2192 1691 2196
rect 1695 2192 1696 2196
rect 1206 2191 1212 2192
rect 1690 2191 1696 2192
rect 1842 2189 1843 2195
rect 1849 2194 3619 2195
rect 1849 2190 1871 2194
rect 1875 2190 1895 2194
rect 1899 2190 2023 2194
rect 2027 2190 2175 2194
rect 2179 2190 2199 2194
rect 2203 2190 2295 2194
rect 2299 2190 2359 2194
rect 2363 2190 2399 2194
rect 2403 2190 2519 2194
rect 2523 2190 2567 2194
rect 2571 2190 2639 2194
rect 2643 2190 2759 2194
rect 2763 2190 2783 2194
rect 2787 2190 2879 2194
rect 2883 2190 2991 2194
rect 2995 2190 3015 2194
rect 3019 2190 3095 2194
rect 3099 2190 3199 2194
rect 3203 2190 3247 2194
rect 3251 2190 3303 2194
rect 3307 2190 3407 2194
rect 3411 2190 3487 2194
rect 3491 2190 3503 2194
rect 3507 2190 3591 2194
rect 3595 2190 3619 2194
rect 1849 2189 3619 2190
rect 3625 2189 3626 2195
rect 96 2177 97 2183
rect 103 2182 1855 2183
rect 103 2178 111 2182
rect 115 2178 143 2182
rect 147 2178 191 2182
rect 195 2178 223 2182
rect 227 2178 303 2182
rect 307 2178 311 2182
rect 315 2178 391 2182
rect 395 2178 463 2182
rect 467 2178 527 2182
rect 531 2178 639 2182
rect 643 2178 679 2182
rect 683 2178 823 2182
rect 827 2178 839 2182
rect 843 2178 1007 2182
rect 1011 2178 1015 2182
rect 1019 2178 1167 2182
rect 1171 2178 1199 2182
rect 1203 2178 1319 2182
rect 1323 2178 1391 2182
rect 1395 2178 1463 2182
rect 1467 2178 1583 2182
rect 1587 2178 1615 2182
rect 1619 2178 1751 2182
rect 1755 2178 1831 2182
rect 1835 2178 1855 2182
rect 103 2177 1855 2178
rect 1861 2177 1862 2183
rect 198 2172 204 2173
rect 470 2172 476 2173
rect 198 2168 199 2172
rect 203 2168 471 2172
rect 475 2168 476 2172
rect 198 2167 204 2168
rect 470 2167 476 2168
rect 646 2172 652 2173
rect 1022 2172 1028 2173
rect 646 2168 647 2172
rect 651 2168 1023 2172
rect 1027 2168 1028 2172
rect 646 2167 652 2168
rect 1022 2167 1028 2168
rect 2214 2132 2220 2133
rect 2486 2132 2492 2133
rect 2214 2128 2215 2132
rect 2219 2128 2487 2132
rect 2491 2128 2492 2132
rect 2214 2127 2220 2128
rect 2486 2127 2492 2128
rect 84 2097 85 2103
rect 91 2102 1843 2103
rect 91 2098 111 2102
rect 115 2098 183 2102
rect 187 2098 215 2102
rect 219 2098 303 2102
rect 307 2098 359 2102
rect 363 2098 455 2102
rect 459 2098 519 2102
rect 523 2098 631 2102
rect 635 2098 703 2102
rect 707 2098 815 2102
rect 819 2098 895 2102
rect 899 2098 1007 2102
rect 1011 2098 1103 2102
rect 1107 2098 1191 2102
rect 1195 2098 1311 2102
rect 1315 2098 1383 2102
rect 1387 2098 1527 2102
rect 1531 2098 1575 2102
rect 1579 2098 1743 2102
rect 1747 2098 1831 2102
rect 1835 2098 1843 2102
rect 91 2097 1843 2098
rect 1849 2097 1850 2103
rect 1854 2101 1855 2107
rect 1861 2106 3631 2107
rect 1861 2102 1871 2106
rect 1875 2102 2175 2106
rect 2179 2102 2207 2106
rect 2211 2102 2271 2106
rect 2275 2102 2303 2106
rect 2307 2102 2375 2106
rect 2379 2102 2407 2106
rect 2411 2102 2487 2106
rect 2491 2102 2527 2106
rect 2531 2102 2607 2106
rect 2611 2102 2647 2106
rect 2651 2102 2727 2106
rect 2731 2102 2767 2106
rect 2771 2102 2847 2106
rect 2851 2102 2887 2106
rect 2891 2102 2967 2106
rect 2971 2102 2999 2106
rect 3003 2102 3079 2106
rect 3083 2102 3103 2106
rect 3107 2102 3191 2106
rect 3195 2102 3207 2106
rect 3211 2102 3303 2106
rect 3307 2102 3311 2106
rect 3315 2102 3415 2106
rect 3419 2102 3511 2106
rect 3515 2102 3591 2106
rect 3595 2102 3631 2106
rect 1861 2101 3631 2102
rect 3637 2101 3638 2107
rect 1842 2031 1843 2037
rect 1849 2031 1874 2037
rect 1868 2027 1874 2031
rect 96 2021 97 2027
rect 103 2026 1855 2027
rect 103 2022 111 2026
rect 115 2022 143 2026
rect 147 2022 223 2026
rect 227 2022 263 2026
rect 267 2022 367 2026
rect 371 2022 383 2026
rect 387 2022 495 2026
rect 499 2022 527 2026
rect 531 2022 607 2026
rect 611 2022 711 2026
rect 715 2022 719 2026
rect 723 2022 823 2026
rect 827 2022 903 2026
rect 907 2022 927 2026
rect 931 2022 1023 2026
rect 1027 2022 1111 2026
rect 1115 2022 1207 2026
rect 1211 2022 1295 2026
rect 1299 2022 1319 2026
rect 1323 2022 1391 2026
rect 1395 2022 1487 2026
rect 1491 2022 1535 2026
rect 1539 2022 1583 2026
rect 1587 2022 1671 2026
rect 1675 2022 1751 2026
rect 1755 2022 1831 2026
rect 1835 2022 1855 2026
rect 103 2021 1855 2022
rect 1861 2021 1862 2027
rect 1868 2026 3619 2027
rect 1868 2022 1871 2026
rect 1875 2022 2071 2026
rect 2075 2022 2167 2026
rect 2171 2022 2207 2026
rect 2211 2022 2263 2026
rect 2267 2022 2359 2026
rect 2363 2022 2367 2026
rect 2371 2022 2479 2026
rect 2483 2022 2519 2026
rect 2523 2022 2599 2026
rect 2603 2022 2679 2026
rect 2683 2022 2719 2026
rect 2723 2022 2839 2026
rect 2843 2022 2847 2026
rect 2851 2022 2959 2026
rect 2963 2022 3015 2026
rect 3019 2022 3071 2026
rect 3075 2022 3183 2026
rect 3187 2022 3295 2026
rect 3299 2022 3351 2026
rect 3355 2022 3407 2026
rect 3411 2022 3503 2026
rect 3507 2022 3591 2026
rect 3595 2022 3619 2026
rect 1868 2021 3619 2022
rect 3625 2021 3626 2027
rect 2382 1972 2388 1973
rect 2598 1972 2604 1973
rect 2382 1968 2383 1972
rect 2387 1968 2599 1972
rect 2603 1968 2604 1972
rect 2382 1967 2388 1968
rect 2598 1967 2604 1968
rect 1854 1945 1855 1951
rect 1861 1950 3631 1951
rect 1861 1946 1871 1950
rect 1875 1946 1903 1950
rect 1907 1946 2007 1950
rect 2011 1946 2079 1950
rect 2083 1946 2135 1950
rect 2139 1946 2215 1950
rect 2219 1946 2255 1950
rect 2259 1946 2367 1950
rect 2371 1946 2375 1950
rect 2379 1946 2487 1950
rect 2491 1946 2527 1950
rect 2531 1946 2599 1950
rect 2603 1946 2687 1950
rect 2691 1946 2719 1950
rect 2723 1946 2839 1950
rect 2843 1946 2855 1950
rect 2859 1946 3023 1950
rect 3027 1946 3191 1950
rect 3195 1946 3359 1950
rect 3363 1946 3511 1950
rect 3515 1946 3591 1950
rect 3595 1946 3631 1950
rect 1861 1945 3631 1946
rect 3637 1945 3638 1951
rect 84 1937 85 1943
rect 91 1942 1843 1943
rect 91 1938 111 1942
rect 115 1938 135 1942
rect 139 1938 167 1942
rect 171 1938 255 1942
rect 259 1938 327 1942
rect 331 1938 375 1942
rect 379 1938 487 1942
rect 491 1938 599 1942
rect 603 1938 647 1942
rect 651 1938 711 1942
rect 715 1938 799 1942
rect 803 1938 815 1942
rect 819 1938 919 1942
rect 923 1938 943 1942
rect 947 1938 1015 1942
rect 1019 1938 1079 1942
rect 1083 1938 1103 1942
rect 1107 1938 1199 1942
rect 1203 1938 1215 1942
rect 1219 1938 1287 1942
rect 1291 1938 1351 1942
rect 1355 1938 1383 1942
rect 1387 1938 1479 1942
rect 1483 1938 1487 1942
rect 1491 1938 1575 1942
rect 1579 1938 1623 1942
rect 1627 1938 1663 1942
rect 1667 1938 1743 1942
rect 1747 1938 1831 1942
rect 1835 1938 1843 1942
rect 91 1937 1843 1938
rect 1849 1937 1850 1943
rect 1842 1871 1843 1877
rect 1849 1875 1874 1877
rect 1849 1874 3619 1875
rect 1849 1871 1871 1874
rect 1868 1870 1871 1871
rect 1875 1870 1895 1874
rect 1899 1870 1991 1874
rect 1995 1870 1999 1874
rect 2003 1870 2119 1874
rect 2123 1870 2127 1874
rect 2131 1870 2247 1874
rect 2251 1870 2367 1874
rect 2371 1870 2383 1874
rect 2387 1870 2479 1874
rect 2483 1870 2519 1874
rect 2523 1870 2591 1874
rect 2595 1870 2655 1874
rect 2659 1870 2711 1874
rect 2715 1870 2807 1874
rect 2811 1870 2831 1874
rect 2835 1870 2975 1874
rect 2979 1870 3151 1874
rect 3155 1870 3335 1874
rect 3339 1870 3503 1874
rect 3507 1870 3591 1874
rect 3595 1870 3619 1874
rect 1868 1869 3619 1870
rect 3625 1869 3626 1875
rect 96 1861 97 1867
rect 103 1866 1855 1867
rect 103 1862 111 1866
rect 115 1862 159 1866
rect 163 1862 175 1866
rect 179 1862 303 1866
rect 307 1862 335 1866
rect 339 1862 447 1866
rect 451 1862 495 1866
rect 499 1862 599 1866
rect 603 1862 655 1866
rect 659 1862 751 1866
rect 755 1862 807 1866
rect 811 1862 903 1866
rect 907 1862 951 1866
rect 955 1862 1055 1866
rect 1059 1862 1087 1866
rect 1091 1862 1207 1866
rect 1211 1862 1223 1866
rect 1227 1862 1351 1866
rect 1355 1862 1359 1866
rect 1363 1862 1487 1866
rect 1491 1862 1495 1866
rect 1499 1862 1631 1866
rect 1635 1862 1751 1866
rect 1755 1862 1831 1866
rect 1835 1862 1855 1866
rect 103 1861 1855 1862
rect 1861 1861 1862 1867
rect 182 1844 188 1845
rect 454 1844 460 1845
rect 182 1840 183 1844
rect 187 1840 455 1844
rect 459 1840 460 1844
rect 182 1839 188 1840
rect 454 1839 460 1840
rect 2694 1796 2700 1797
rect 3258 1796 3264 1797
rect 2694 1792 2695 1796
rect 2699 1792 3259 1796
rect 3263 1792 3264 1796
rect 2694 1791 2700 1792
rect 3258 1791 3264 1792
rect 84 1781 85 1787
rect 91 1786 1843 1787
rect 91 1782 111 1786
rect 115 1782 151 1786
rect 155 1782 247 1786
rect 251 1782 295 1786
rect 299 1782 423 1786
rect 427 1782 439 1786
rect 443 1782 591 1786
rect 595 1782 743 1786
rect 747 1782 751 1786
rect 755 1782 895 1786
rect 899 1782 1023 1786
rect 1027 1782 1047 1786
rect 1051 1782 1143 1786
rect 1147 1782 1199 1786
rect 1203 1782 1263 1786
rect 1267 1782 1343 1786
rect 1347 1782 1391 1786
rect 1395 1782 1479 1786
rect 1483 1782 1623 1786
rect 1627 1782 1743 1786
rect 1747 1782 1831 1786
rect 1835 1782 1843 1786
rect 91 1781 1843 1782
rect 1849 1781 1850 1787
rect 1854 1781 1855 1787
rect 1861 1786 3631 1787
rect 1861 1782 1871 1786
rect 1875 1782 1903 1786
rect 1907 1782 1999 1786
rect 2003 1782 2031 1786
rect 2035 1782 2127 1786
rect 2131 1782 2191 1786
rect 2195 1782 2255 1786
rect 2259 1782 2359 1786
rect 2363 1782 2391 1786
rect 2395 1782 2527 1786
rect 2531 1782 2663 1786
rect 2667 1782 2687 1786
rect 2691 1782 2815 1786
rect 2819 1782 2839 1786
rect 2843 1782 2983 1786
rect 2987 1782 3119 1786
rect 3123 1782 3159 1786
rect 3163 1782 3255 1786
rect 3259 1782 3343 1786
rect 3347 1782 3391 1786
rect 3395 1782 3511 1786
rect 3515 1782 3591 1786
rect 3595 1782 3631 1786
rect 1861 1781 3631 1782
rect 3637 1781 3638 1787
rect 910 1724 916 1725
rect 1342 1724 1348 1725
rect 910 1720 911 1724
rect 915 1720 1343 1724
rect 1347 1720 1348 1724
rect 910 1719 916 1720
rect 1342 1719 1348 1720
rect 1842 1711 1843 1717
rect 1849 1711 1874 1717
rect 1868 1707 1874 1711
rect 96 1701 97 1707
rect 103 1706 1855 1707
rect 103 1702 111 1706
rect 115 1702 191 1706
rect 195 1702 255 1706
rect 259 1702 311 1706
rect 315 1702 431 1706
rect 435 1702 447 1706
rect 451 1702 591 1706
rect 595 1702 599 1706
rect 603 1702 743 1706
rect 747 1702 759 1706
rect 763 1702 895 1706
rect 899 1702 903 1706
rect 907 1702 1031 1706
rect 1035 1702 1039 1706
rect 1043 1702 1151 1706
rect 1155 1702 1183 1706
rect 1187 1702 1271 1706
rect 1275 1702 1319 1706
rect 1323 1702 1399 1706
rect 1403 1702 1447 1706
rect 1451 1702 1575 1706
rect 1579 1702 1711 1706
rect 1715 1702 1831 1706
rect 1835 1702 1855 1706
rect 103 1701 1855 1702
rect 1861 1701 1862 1707
rect 1868 1706 3619 1707
rect 1868 1702 1871 1706
rect 1875 1702 1895 1706
rect 1899 1702 1991 1706
rect 1995 1702 2023 1706
rect 2027 1702 2135 1706
rect 2139 1702 2183 1706
rect 2187 1702 2295 1706
rect 2299 1702 2351 1706
rect 2355 1702 2471 1706
rect 2475 1702 2519 1706
rect 2523 1702 2647 1706
rect 2651 1702 2679 1706
rect 2683 1702 2815 1706
rect 2819 1702 2831 1706
rect 2835 1702 2967 1706
rect 2971 1702 2975 1706
rect 2979 1702 3111 1706
rect 3115 1702 3247 1706
rect 3251 1702 3383 1706
rect 3387 1702 3503 1706
rect 3507 1702 3591 1706
rect 3595 1702 3619 1706
rect 1868 1701 3619 1702
rect 3625 1701 3626 1707
rect 1910 1692 1916 1693
rect 2418 1692 2424 1693
rect 1910 1688 1911 1692
rect 1915 1688 2419 1692
rect 2423 1688 2424 1692
rect 1910 1687 1916 1688
rect 2418 1687 2424 1688
rect 2830 1644 2836 1645
rect 3186 1644 3192 1645
rect 2830 1640 2831 1644
rect 2835 1640 3187 1644
rect 3191 1640 3192 1644
rect 2830 1639 2836 1640
rect 3186 1639 3192 1640
rect 84 1617 85 1623
rect 91 1622 1843 1623
rect 91 1618 111 1622
rect 115 1618 167 1622
rect 171 1618 183 1622
rect 187 1618 303 1622
rect 307 1618 351 1622
rect 355 1618 439 1622
rect 443 1618 543 1622
rect 547 1618 583 1622
rect 587 1618 727 1622
rect 731 1618 735 1622
rect 739 1618 887 1622
rect 891 1618 903 1622
rect 907 1618 1031 1622
rect 1035 1618 1071 1622
rect 1075 1618 1175 1622
rect 1179 1618 1223 1622
rect 1227 1618 1311 1622
rect 1315 1618 1359 1622
rect 1363 1618 1439 1622
rect 1443 1618 1495 1622
rect 1499 1618 1567 1622
rect 1571 1618 1623 1622
rect 1627 1618 1703 1622
rect 1707 1618 1743 1622
rect 1747 1618 1831 1622
rect 1835 1618 1843 1622
rect 91 1617 1843 1618
rect 1849 1617 1850 1623
rect 1854 1621 1855 1627
rect 1861 1626 3631 1627
rect 1861 1622 1871 1626
rect 1875 1622 1903 1626
rect 1907 1622 1975 1626
rect 1979 1622 1999 1626
rect 2003 1622 2095 1626
rect 2099 1622 2143 1626
rect 2147 1622 2231 1626
rect 2235 1622 2303 1626
rect 2307 1622 2367 1626
rect 2371 1622 2479 1626
rect 2483 1622 2503 1626
rect 2507 1622 2639 1626
rect 2643 1622 2655 1626
rect 2659 1622 2775 1626
rect 2779 1622 2823 1626
rect 2827 1622 2911 1626
rect 2915 1622 2975 1626
rect 2979 1622 3055 1626
rect 3059 1622 3119 1626
rect 3123 1622 3207 1626
rect 3211 1622 3255 1626
rect 3259 1622 3367 1626
rect 3371 1622 3391 1626
rect 3395 1622 3511 1626
rect 3515 1622 3591 1626
rect 3595 1622 3631 1626
rect 1861 1621 3631 1622
rect 3637 1621 3638 1627
rect 1842 1547 1843 1553
rect 1849 1547 1874 1553
rect 1868 1546 3619 1547
rect 96 1537 97 1543
rect 103 1542 1855 1543
rect 103 1538 111 1542
rect 115 1538 143 1542
rect 147 1538 175 1542
rect 179 1538 247 1542
rect 251 1538 359 1542
rect 363 1538 383 1542
rect 387 1538 527 1542
rect 531 1538 551 1542
rect 555 1538 671 1542
rect 675 1538 735 1542
rect 739 1538 815 1542
rect 819 1538 911 1542
rect 915 1538 951 1542
rect 955 1538 1079 1542
rect 1083 1538 1207 1542
rect 1211 1538 1231 1542
rect 1235 1538 1335 1542
rect 1339 1538 1367 1542
rect 1371 1538 1471 1542
rect 1475 1538 1503 1542
rect 1507 1538 1631 1542
rect 1635 1538 1751 1542
rect 1755 1538 1831 1542
rect 1835 1538 1855 1542
rect 103 1537 1855 1538
rect 1861 1537 1862 1543
rect 1868 1542 1871 1546
rect 1875 1542 1967 1546
rect 1971 1542 2087 1546
rect 2091 1542 2167 1546
rect 2171 1542 2223 1546
rect 2227 1542 2255 1546
rect 2259 1542 2343 1546
rect 2347 1542 2359 1546
rect 2363 1542 2439 1546
rect 2443 1542 2495 1546
rect 2499 1542 2535 1546
rect 2539 1542 2631 1546
rect 2635 1542 2647 1546
rect 2651 1542 2767 1546
rect 2771 1542 2783 1546
rect 2787 1542 2903 1546
rect 2907 1542 2943 1546
rect 2947 1542 3047 1546
rect 3051 1542 3119 1546
rect 3123 1542 3199 1546
rect 3203 1542 3303 1546
rect 3307 1542 3359 1546
rect 3363 1542 3495 1546
rect 3499 1542 3503 1546
rect 3507 1542 3591 1546
rect 3595 1542 3619 1546
rect 1868 1541 3619 1542
rect 3625 1541 3626 1547
rect 2102 1532 2108 1533
rect 2418 1532 2424 1533
rect 2102 1528 2103 1532
rect 2107 1528 2419 1532
rect 2423 1528 2424 1532
rect 2102 1527 2108 1528
rect 2418 1527 2424 1528
rect 2662 1484 2668 1485
rect 3202 1484 3208 1485
rect 2662 1480 2663 1484
rect 2667 1480 3203 1484
rect 3207 1480 3208 1484
rect 2662 1479 2668 1480
rect 3202 1479 3208 1480
rect 958 1476 964 1477
rect 1218 1476 1224 1477
rect 958 1472 959 1476
rect 963 1472 1219 1476
rect 1223 1472 1224 1476
rect 958 1471 964 1472
rect 1218 1471 1224 1472
rect 2270 1476 2276 1477
rect 2514 1476 2520 1477
rect 2270 1472 2271 1476
rect 2275 1472 2515 1476
rect 2519 1472 2520 1476
rect 2270 1471 2276 1472
rect 2514 1471 2520 1472
rect 84 1457 85 1463
rect 91 1462 1843 1463
rect 91 1458 111 1462
rect 115 1458 135 1462
rect 139 1458 231 1462
rect 235 1458 239 1462
rect 243 1458 359 1462
rect 363 1458 375 1462
rect 379 1458 479 1462
rect 483 1458 519 1462
rect 523 1458 599 1462
rect 603 1458 663 1462
rect 667 1458 719 1462
rect 723 1458 807 1462
rect 811 1458 831 1462
rect 835 1458 935 1462
rect 939 1458 943 1462
rect 947 1458 1039 1462
rect 1043 1458 1071 1462
rect 1075 1458 1143 1462
rect 1147 1458 1199 1462
rect 1203 1458 1255 1462
rect 1259 1458 1327 1462
rect 1331 1458 1463 1462
rect 1467 1458 1831 1462
rect 1835 1458 1843 1462
rect 91 1457 1843 1458
rect 1849 1457 1850 1463
rect 1854 1461 1855 1467
rect 1861 1466 3631 1467
rect 1861 1462 1871 1466
rect 1875 1462 2095 1466
rect 2099 1462 2175 1466
rect 2179 1462 2263 1466
rect 2267 1462 2343 1466
rect 2347 1462 2351 1466
rect 2355 1462 2423 1466
rect 2427 1462 2447 1466
rect 2451 1462 2503 1466
rect 2507 1462 2543 1466
rect 2547 1462 2607 1466
rect 2611 1462 2655 1466
rect 2659 1462 2735 1466
rect 2739 1462 2791 1466
rect 2795 1462 2895 1466
rect 2899 1462 2951 1466
rect 2955 1462 3079 1466
rect 3083 1462 3127 1466
rect 3131 1462 3279 1466
rect 3283 1462 3311 1466
rect 3315 1462 3479 1466
rect 3483 1462 3503 1466
rect 3507 1462 3591 1466
rect 3595 1462 3631 1466
rect 1861 1461 3631 1462
rect 3637 1461 3638 1467
rect 2842 1436 2848 1437
rect 3286 1436 3292 1437
rect 2842 1432 2843 1436
rect 2847 1432 3287 1436
rect 3291 1432 3292 1436
rect 2842 1431 2848 1432
rect 3286 1431 3292 1432
rect 1842 1385 1843 1391
rect 1849 1390 3619 1391
rect 1849 1386 1871 1390
rect 1875 1386 2255 1390
rect 2259 1386 2263 1390
rect 2267 1386 2335 1390
rect 2339 1386 2343 1390
rect 2347 1386 2415 1390
rect 2419 1386 2423 1390
rect 2427 1386 2495 1390
rect 2499 1386 2503 1390
rect 2507 1386 2591 1390
rect 2595 1386 2599 1390
rect 2603 1386 2695 1390
rect 2699 1386 2727 1390
rect 2731 1386 2807 1390
rect 2811 1386 2887 1390
rect 2891 1386 2919 1390
rect 2923 1386 3039 1390
rect 3043 1386 3071 1390
rect 3075 1386 3159 1390
rect 3163 1386 3271 1390
rect 3275 1386 3279 1390
rect 3283 1386 3399 1390
rect 3403 1386 3471 1390
rect 3475 1386 3503 1390
rect 3507 1386 3591 1390
rect 3595 1386 3619 1390
rect 1849 1385 3619 1386
rect 3625 1385 3626 1391
rect 96 1365 97 1371
rect 103 1370 1855 1371
rect 103 1366 111 1370
rect 115 1366 143 1370
rect 147 1366 239 1370
rect 243 1366 287 1370
rect 291 1366 367 1370
rect 371 1366 431 1370
rect 435 1366 487 1370
rect 491 1366 583 1370
rect 587 1366 607 1370
rect 611 1366 727 1370
rect 731 1366 735 1370
rect 739 1366 839 1370
rect 843 1366 879 1370
rect 883 1366 943 1370
rect 947 1366 1023 1370
rect 1027 1366 1047 1370
rect 1051 1366 1151 1370
rect 1155 1366 1167 1370
rect 1171 1366 1263 1370
rect 1267 1366 1319 1370
rect 1323 1366 1471 1370
rect 1475 1366 1623 1370
rect 1627 1366 1831 1370
rect 1835 1366 1855 1370
rect 103 1365 1855 1366
rect 1861 1365 1862 1371
rect 2582 1340 2588 1341
rect 2838 1340 2844 1341
rect 2582 1336 2583 1340
rect 2587 1336 2839 1340
rect 2843 1336 2844 1340
rect 2582 1335 2588 1336
rect 2838 1335 2844 1336
rect 1854 1297 1855 1303
rect 1861 1302 3631 1303
rect 1861 1298 1871 1302
rect 1875 1298 2215 1302
rect 2219 1298 2271 1302
rect 2275 1298 2295 1302
rect 2299 1298 2351 1302
rect 2355 1298 2375 1302
rect 2379 1298 2431 1302
rect 2435 1298 2455 1302
rect 2459 1298 2511 1302
rect 2515 1298 2551 1302
rect 2555 1298 2599 1302
rect 2603 1298 2663 1302
rect 2667 1298 2703 1302
rect 2707 1298 2791 1302
rect 2795 1298 2815 1302
rect 2819 1298 2927 1302
rect 2931 1298 3047 1302
rect 3051 1298 3071 1302
rect 3075 1298 3167 1302
rect 3171 1298 3215 1302
rect 3219 1298 3287 1302
rect 3291 1298 3367 1302
rect 3371 1298 3407 1302
rect 3411 1298 3511 1302
rect 3515 1298 3591 1302
rect 3595 1298 3631 1302
rect 1861 1297 3631 1298
rect 3637 1297 3638 1303
rect 84 1285 85 1291
rect 91 1290 1843 1291
rect 91 1286 111 1290
rect 115 1286 135 1290
rect 139 1286 263 1290
rect 267 1286 279 1290
rect 283 1286 423 1290
rect 427 1286 575 1290
rect 579 1286 591 1290
rect 595 1286 727 1290
rect 731 1286 759 1290
rect 763 1286 871 1290
rect 875 1286 927 1290
rect 931 1286 1015 1290
rect 1019 1286 1079 1290
rect 1083 1286 1159 1290
rect 1163 1286 1223 1290
rect 1227 1286 1311 1290
rect 1315 1286 1351 1290
rect 1355 1286 1463 1290
rect 1467 1286 1479 1290
rect 1483 1286 1607 1290
rect 1611 1286 1615 1290
rect 1619 1286 1735 1290
rect 1739 1286 1831 1290
rect 1835 1286 1843 1290
rect 91 1285 1843 1286
rect 1849 1285 1850 1291
rect 1094 1228 1100 1229
rect 1290 1228 1296 1229
rect 1094 1224 1095 1228
rect 1099 1224 1291 1228
rect 1295 1224 1296 1228
rect 1094 1223 1100 1224
rect 1290 1223 1296 1224
rect 1842 1217 1843 1223
rect 1849 1222 3619 1223
rect 1849 1218 1871 1222
rect 1875 1218 2111 1222
rect 2115 1218 2207 1222
rect 2211 1218 2287 1222
rect 2291 1218 2303 1222
rect 2307 1218 2367 1222
rect 2371 1218 2407 1222
rect 2411 1218 2447 1222
rect 2451 1218 2527 1222
rect 2531 1218 2543 1222
rect 2547 1218 2647 1222
rect 2651 1218 2655 1222
rect 2659 1218 2775 1222
rect 2779 1218 2783 1222
rect 2787 1218 2911 1222
rect 2915 1218 2919 1222
rect 2923 1218 3055 1222
rect 3059 1218 3063 1222
rect 3067 1218 3199 1222
rect 3203 1218 3207 1222
rect 3211 1218 3343 1222
rect 3347 1218 3359 1222
rect 3363 1218 3495 1222
rect 3499 1218 3503 1222
rect 3507 1218 3591 1222
rect 3595 1218 3619 1222
rect 1849 1217 3619 1218
rect 3625 1217 3626 1223
rect 96 1201 97 1207
rect 103 1206 1855 1207
rect 103 1202 111 1206
rect 115 1202 143 1206
rect 147 1202 271 1206
rect 275 1202 311 1206
rect 315 1202 431 1206
rect 435 1202 487 1206
rect 491 1202 599 1206
rect 603 1202 671 1206
rect 675 1202 767 1206
rect 771 1202 847 1206
rect 851 1202 935 1206
rect 939 1202 1007 1206
rect 1011 1202 1087 1206
rect 1091 1202 1159 1206
rect 1163 1202 1231 1206
rect 1235 1202 1295 1206
rect 1299 1202 1359 1206
rect 1363 1202 1415 1206
rect 1419 1202 1487 1206
rect 1491 1202 1535 1206
rect 1539 1202 1615 1206
rect 1619 1202 1655 1206
rect 1659 1202 1743 1206
rect 1747 1202 1751 1206
rect 1755 1202 1831 1206
rect 1835 1202 1855 1206
rect 103 1201 1855 1202
rect 1861 1201 1862 1207
rect 422 1196 428 1197
rect 678 1196 684 1197
rect 422 1192 423 1196
rect 427 1192 679 1196
rect 683 1192 684 1196
rect 422 1191 428 1192
rect 678 1191 684 1192
rect 2582 1164 2588 1165
rect 2998 1164 3004 1165
rect 2582 1160 2583 1164
rect 2587 1160 2999 1164
rect 3003 1160 3004 1164
rect 2582 1159 2588 1160
rect 2998 1159 3004 1160
rect 1854 1133 1855 1139
rect 1861 1138 3631 1139
rect 1861 1134 1871 1138
rect 1875 1134 1903 1138
rect 1907 1134 2119 1138
rect 2123 1134 2127 1138
rect 2131 1134 2215 1138
rect 2219 1134 2311 1138
rect 2315 1134 2359 1138
rect 2363 1134 2415 1138
rect 2419 1134 2535 1138
rect 2539 1134 2575 1138
rect 2579 1134 2655 1138
rect 2659 1134 2775 1138
rect 2779 1134 2783 1138
rect 2787 1134 2919 1138
rect 2923 1134 2967 1138
rect 2971 1134 3063 1138
rect 3067 1134 3159 1138
rect 3163 1134 3207 1138
rect 3211 1134 3343 1138
rect 3347 1134 3351 1138
rect 3355 1134 3503 1138
rect 3507 1134 3511 1138
rect 3515 1134 3591 1138
rect 3595 1134 3631 1138
rect 1861 1133 3631 1134
rect 3637 1133 3638 1139
rect 84 1125 85 1131
rect 91 1130 1843 1131
rect 91 1126 111 1130
rect 115 1126 135 1130
rect 139 1126 247 1130
rect 251 1126 303 1130
rect 307 1126 383 1130
rect 387 1126 479 1130
rect 483 1126 519 1130
rect 523 1126 647 1130
rect 651 1126 663 1130
rect 667 1126 775 1130
rect 779 1126 839 1130
rect 843 1126 895 1130
rect 899 1126 999 1130
rect 1003 1126 1015 1130
rect 1019 1126 1135 1130
rect 1139 1126 1151 1130
rect 1155 1126 1255 1130
rect 1259 1126 1287 1130
rect 1291 1126 1375 1130
rect 1379 1126 1407 1130
rect 1411 1126 1503 1130
rect 1507 1126 1527 1130
rect 1531 1126 1631 1130
rect 1635 1126 1647 1130
rect 1651 1126 1743 1130
rect 1747 1126 1831 1130
rect 1835 1126 1843 1130
rect 91 1125 1843 1126
rect 1849 1125 1850 1131
rect 1842 1057 1843 1063
rect 1849 1062 3619 1063
rect 1849 1058 1871 1062
rect 1875 1058 1895 1062
rect 1899 1058 2015 1062
rect 2019 1058 2119 1062
rect 2123 1058 2167 1062
rect 2171 1058 2327 1062
rect 2331 1058 2351 1062
rect 2355 1058 2487 1062
rect 2491 1058 2567 1062
rect 2571 1058 2639 1062
rect 2643 1058 2767 1062
rect 2771 1058 2791 1062
rect 2795 1058 2935 1062
rect 2939 1058 2959 1062
rect 2963 1058 3079 1062
rect 3083 1058 3151 1062
rect 3155 1058 3223 1062
rect 3227 1058 3335 1062
rect 3339 1058 3375 1062
rect 3379 1058 3503 1062
rect 3507 1058 3591 1062
rect 3595 1058 3619 1062
rect 1849 1057 3619 1058
rect 3625 1057 3626 1063
rect 96 1037 97 1043
rect 103 1042 1855 1043
rect 103 1038 111 1042
rect 115 1038 143 1042
rect 147 1038 239 1042
rect 243 1038 255 1042
rect 259 1038 359 1042
rect 363 1038 391 1042
rect 395 1038 471 1042
rect 475 1038 527 1042
rect 531 1038 575 1042
rect 579 1038 655 1042
rect 659 1038 671 1042
rect 675 1038 767 1042
rect 771 1038 783 1042
rect 787 1038 855 1042
rect 859 1038 903 1042
rect 907 1038 943 1042
rect 947 1038 1023 1042
rect 1027 1038 1031 1042
rect 1035 1038 1127 1042
rect 1131 1038 1143 1042
rect 1147 1038 1223 1042
rect 1227 1038 1263 1042
rect 1267 1038 1383 1042
rect 1387 1038 1511 1042
rect 1515 1038 1639 1042
rect 1643 1038 1751 1042
rect 1755 1038 1831 1042
rect 1835 1038 1855 1042
rect 103 1037 1855 1038
rect 1861 1037 1862 1043
rect 1854 977 1855 983
rect 1861 982 3631 983
rect 1861 978 1871 982
rect 1875 978 1903 982
rect 1907 978 1983 982
rect 1987 978 2023 982
rect 2027 978 2079 982
rect 2083 978 2175 982
rect 2179 978 2199 982
rect 2203 978 2335 982
rect 2339 978 2479 982
rect 2483 978 2495 982
rect 2499 978 2631 982
rect 2635 978 2647 982
rect 2651 978 2791 982
rect 2795 978 2799 982
rect 2803 978 2943 982
rect 2947 978 2967 982
rect 2971 978 3087 982
rect 3091 978 3151 982
rect 3155 978 3231 982
rect 3235 978 3343 982
rect 3347 978 3383 982
rect 3387 978 3511 982
rect 3515 978 3591 982
rect 3595 978 3631 982
rect 1861 977 3631 978
rect 3637 977 3638 983
rect 84 949 85 955
rect 91 954 1843 955
rect 91 950 111 954
rect 115 950 135 954
rect 139 950 231 954
rect 235 950 263 954
rect 267 950 351 954
rect 355 950 415 954
rect 419 950 463 954
rect 467 950 559 954
rect 563 950 567 954
rect 571 950 663 954
rect 667 950 703 954
rect 707 950 759 954
rect 763 950 839 954
rect 843 950 847 954
rect 851 950 935 954
rect 939 950 975 954
rect 979 950 1023 954
rect 1027 950 1103 954
rect 1107 950 1119 954
rect 1123 950 1215 954
rect 1219 950 1223 954
rect 1227 950 1335 954
rect 1339 950 1439 954
rect 1443 950 1543 954
rect 1547 950 1655 954
rect 1659 950 1743 954
rect 1747 950 1831 954
rect 1835 950 1843 954
rect 91 949 1843 950
rect 1849 949 1850 955
rect 1842 889 1843 895
rect 1849 894 3619 895
rect 1849 890 1871 894
rect 1875 890 1895 894
rect 1899 890 1919 894
rect 1923 890 1975 894
rect 1979 890 2071 894
rect 2075 890 2095 894
rect 2099 890 2191 894
rect 2195 890 2271 894
rect 2275 890 2327 894
rect 2331 890 2455 894
rect 2459 890 2471 894
rect 2475 890 2623 894
rect 2627 890 2655 894
rect 2659 890 2783 894
rect 2787 890 2863 894
rect 2867 890 2959 894
rect 2963 890 3079 894
rect 3083 890 3143 894
rect 3147 890 3303 894
rect 3307 890 3335 894
rect 3339 890 3503 894
rect 3507 890 3591 894
rect 3595 890 3619 894
rect 1849 889 3619 890
rect 3625 889 3626 895
rect 96 869 97 875
rect 103 874 1855 875
rect 103 870 111 874
rect 115 870 143 874
rect 147 870 247 874
rect 251 870 271 874
rect 275 870 383 874
rect 387 870 423 874
rect 427 870 519 874
rect 523 870 567 874
rect 571 870 663 874
rect 667 870 711 874
rect 715 870 815 874
rect 819 870 847 874
rect 851 870 959 874
rect 963 870 983 874
rect 987 870 1103 874
rect 1107 870 1111 874
rect 1115 870 1231 874
rect 1235 870 1247 874
rect 1251 870 1343 874
rect 1347 870 1383 874
rect 1387 870 1447 874
rect 1451 870 1511 874
rect 1515 870 1551 874
rect 1555 870 1639 874
rect 1643 870 1663 874
rect 1667 870 1751 874
rect 1755 870 1831 874
rect 1835 870 1855 874
rect 103 869 1855 870
rect 1861 869 1862 875
rect 258 844 264 845
rect 526 844 532 845
rect 258 840 259 844
rect 263 840 527 844
rect 531 840 532 844
rect 258 839 264 840
rect 526 839 532 840
rect 1854 813 1855 819
rect 1861 818 3631 819
rect 1861 814 1871 818
rect 1875 814 1903 818
rect 1907 814 1927 818
rect 1931 814 2015 818
rect 2019 814 2103 818
rect 2107 814 2167 818
rect 2171 814 2279 818
rect 2283 814 2327 818
rect 2331 814 2463 818
rect 2467 814 2487 818
rect 2491 814 2647 818
rect 2651 814 2663 818
rect 2667 814 2807 818
rect 2811 814 2871 818
rect 2875 814 2959 818
rect 2963 814 3087 818
rect 3091 814 3103 818
rect 3107 814 3247 818
rect 3251 814 3311 818
rect 3315 814 3391 818
rect 3395 814 3511 818
rect 3515 814 3591 818
rect 3595 814 3631 818
rect 1861 813 3631 814
rect 3637 813 3638 819
rect 84 781 85 787
rect 91 786 1843 787
rect 91 782 111 786
rect 115 782 135 786
rect 139 782 215 786
rect 219 782 239 786
rect 243 782 303 786
rect 307 782 375 786
rect 379 782 415 786
rect 419 782 511 786
rect 515 782 543 786
rect 547 782 655 786
rect 659 782 687 786
rect 691 782 807 786
rect 811 782 839 786
rect 843 782 951 786
rect 955 782 991 786
rect 995 782 1095 786
rect 1099 782 1143 786
rect 1147 782 1239 786
rect 1243 782 1295 786
rect 1299 782 1375 786
rect 1379 782 1447 786
rect 1451 782 1503 786
rect 1507 782 1607 786
rect 1611 782 1631 786
rect 1635 782 1743 786
rect 1747 782 1831 786
rect 1835 782 1843 786
rect 91 781 1843 782
rect 1849 781 1850 787
rect 1842 737 1843 743
rect 1849 742 3619 743
rect 1849 738 1871 742
rect 1875 738 1895 742
rect 1899 738 1967 742
rect 1971 738 2007 742
rect 2011 738 2063 742
rect 2067 738 2159 742
rect 2163 738 2175 742
rect 2179 738 2303 742
rect 2307 738 2319 742
rect 2323 738 2447 742
rect 2451 738 2479 742
rect 2483 738 2599 742
rect 2603 738 2639 742
rect 2643 738 2751 742
rect 2755 738 2799 742
rect 2803 738 2903 742
rect 2907 738 2951 742
rect 2955 738 3055 742
rect 3059 738 3095 742
rect 3099 738 3207 742
rect 3211 738 3239 742
rect 3243 738 3359 742
rect 3363 738 3383 742
rect 3387 738 3503 742
rect 3507 738 3591 742
rect 3595 738 3619 742
rect 1849 737 3619 738
rect 3625 737 3626 743
rect 150 724 156 725
rect 654 724 660 725
rect 150 720 151 724
rect 155 720 655 724
rect 659 720 660 724
rect 150 719 156 720
rect 654 719 660 720
rect 1310 724 1316 725
rect 1530 724 1536 725
rect 1310 720 1311 724
rect 1315 720 1531 724
rect 1535 720 1536 724
rect 1310 719 1316 720
rect 1530 719 1536 720
rect 2190 716 2196 717
rect 2606 716 2612 717
rect 2190 712 2191 716
rect 2195 712 2607 716
rect 2611 712 2612 716
rect 2190 711 2196 712
rect 2606 711 2612 712
rect 96 697 97 703
rect 103 702 1855 703
rect 103 698 111 702
rect 115 698 143 702
rect 147 698 223 702
rect 227 698 231 702
rect 235 698 311 702
rect 315 698 319 702
rect 323 698 423 702
rect 427 698 543 702
rect 547 698 551 702
rect 555 698 679 702
rect 683 698 695 702
rect 699 698 815 702
rect 819 698 847 702
rect 851 698 951 702
rect 955 698 999 702
rect 1003 698 1087 702
rect 1091 698 1151 702
rect 1155 698 1215 702
rect 1219 698 1303 702
rect 1307 698 1335 702
rect 1339 698 1455 702
rect 1459 698 1583 702
rect 1587 698 1615 702
rect 1619 698 1831 702
rect 1835 698 1855 702
rect 103 697 1855 698
rect 1861 697 1862 703
rect 274 684 280 685
rect 550 684 556 685
rect 274 680 275 684
rect 279 680 551 684
rect 555 680 556 684
rect 274 679 280 680
rect 550 679 556 680
rect 1982 676 1988 677
rect 2418 676 2424 677
rect 1982 672 1983 676
rect 1987 672 2419 676
rect 2423 672 2424 676
rect 1982 671 1988 672
rect 2418 671 2424 672
rect 1854 661 1855 667
rect 1861 666 3631 667
rect 1861 662 1871 666
rect 1875 662 1975 666
rect 1979 662 2071 666
rect 2075 662 2175 666
rect 2179 662 2183 666
rect 2187 662 2271 666
rect 2275 662 2311 666
rect 2315 662 2375 666
rect 2379 662 2455 666
rect 2459 662 2487 666
rect 2491 662 2607 666
rect 2611 662 2735 666
rect 2739 662 2759 666
rect 2763 662 2863 666
rect 2867 662 2911 666
rect 2915 662 2991 666
rect 2995 662 3063 666
rect 3067 662 3119 666
rect 3123 662 3215 666
rect 3219 662 3247 666
rect 3251 662 3367 666
rect 3371 662 3375 666
rect 3379 662 3511 666
rect 3515 662 3591 666
rect 3595 662 3631 666
rect 1861 661 3631 662
rect 3637 661 3638 667
rect 1094 628 1100 629
rect 1410 628 1416 629
rect 1094 624 1095 628
rect 1099 624 1411 628
rect 1415 624 1416 628
rect 1094 623 1100 624
rect 1410 623 1416 624
rect 84 613 85 619
rect 91 618 1843 619
rect 91 614 111 618
rect 115 614 223 618
rect 227 614 311 618
rect 315 614 415 618
rect 419 614 447 618
rect 451 614 527 618
rect 531 614 535 618
rect 539 614 607 618
rect 611 614 671 618
rect 675 614 687 618
rect 691 614 775 618
rect 779 614 807 618
rect 811 614 871 618
rect 875 614 943 618
rect 947 614 959 618
rect 963 614 1047 618
rect 1051 614 1079 618
rect 1083 614 1143 618
rect 1147 614 1207 618
rect 1211 614 1239 618
rect 1243 614 1327 618
rect 1331 614 1335 618
rect 1339 614 1431 618
rect 1435 614 1447 618
rect 1451 614 1575 618
rect 1579 614 1831 618
rect 1835 614 1843 618
rect 91 613 1843 614
rect 1849 613 1850 619
rect 1842 585 1843 591
rect 1849 590 3619 591
rect 1849 586 1871 590
rect 1875 586 2167 590
rect 2171 586 2263 590
rect 2267 586 2343 590
rect 2347 586 2367 590
rect 2371 586 2423 590
rect 2427 586 2479 590
rect 2483 586 2503 590
rect 2507 586 2591 590
rect 2595 586 2599 590
rect 2603 586 2695 590
rect 2699 586 2727 590
rect 2731 586 2815 590
rect 2819 586 2855 590
rect 2859 586 2959 590
rect 2963 586 2983 590
rect 2987 586 3111 590
rect 3115 586 3239 590
rect 3243 586 3279 590
rect 3283 586 3367 590
rect 3371 586 3447 590
rect 3451 586 3503 590
rect 3507 586 3591 590
rect 3595 586 3619 590
rect 1849 585 3619 586
rect 3625 585 3626 591
rect 2282 548 2288 549
rect 2538 548 2544 549
rect 2282 544 2283 548
rect 2287 544 2539 548
rect 2543 544 2544 548
rect 2282 543 2288 544
rect 2538 543 2544 544
rect 96 525 97 531
rect 103 530 1855 531
rect 103 526 111 530
rect 115 526 335 530
rect 339 526 423 530
rect 427 526 455 530
rect 459 526 511 530
rect 515 526 535 530
rect 539 526 591 530
rect 595 526 615 530
rect 619 526 671 530
rect 675 526 695 530
rect 699 526 751 530
rect 755 526 783 530
rect 787 526 839 530
rect 843 526 879 530
rect 883 526 927 530
rect 931 526 967 530
rect 971 526 1015 530
rect 1019 526 1055 530
rect 1059 526 1103 530
rect 1107 526 1151 530
rect 1155 526 1191 530
rect 1195 526 1247 530
rect 1251 526 1279 530
rect 1283 526 1343 530
rect 1347 526 1439 530
rect 1443 526 1831 530
rect 1835 526 1855 530
rect 103 525 1855 526
rect 1861 525 1862 531
rect 1854 501 1855 507
rect 1861 506 3631 507
rect 1861 502 1871 506
rect 1875 502 2191 506
rect 2195 502 2271 506
rect 2275 502 2287 506
rect 2291 502 2351 506
rect 2355 502 2383 506
rect 2387 502 2431 506
rect 2435 502 2487 506
rect 2491 502 2511 506
rect 2515 502 2583 506
rect 2587 502 2599 506
rect 2603 502 2687 506
rect 2691 502 2703 506
rect 2707 502 2791 506
rect 2795 502 2823 506
rect 2827 502 2911 506
rect 2915 502 2967 506
rect 2971 502 3039 506
rect 3043 502 3119 506
rect 3123 502 3175 506
rect 3179 502 3287 506
rect 3291 502 3319 506
rect 3323 502 3455 506
rect 3459 502 3471 506
rect 3475 502 3591 506
rect 3595 502 3631 506
rect 1861 501 3631 502
rect 3637 501 3638 507
rect 84 441 85 447
rect 91 446 1843 447
rect 91 442 111 446
rect 115 442 223 446
rect 227 442 327 446
rect 331 442 335 446
rect 339 442 415 446
rect 419 442 447 446
rect 451 442 503 446
rect 507 442 559 446
rect 563 442 583 446
rect 587 442 663 446
rect 667 442 743 446
rect 747 442 759 446
rect 763 442 831 446
rect 835 442 847 446
rect 851 442 919 446
rect 923 442 935 446
rect 939 442 1007 446
rect 1011 442 1023 446
rect 1027 442 1095 446
rect 1099 442 1111 446
rect 1115 442 1183 446
rect 1187 442 1199 446
rect 1203 442 1271 446
rect 1275 442 1295 446
rect 1299 442 1831 446
rect 1835 442 1843 446
rect 91 441 1843 442
rect 1849 441 1850 447
rect 1842 421 1843 427
rect 1849 426 3619 427
rect 1849 422 1871 426
rect 1875 422 1975 426
rect 1979 422 2063 426
rect 2067 422 2159 426
rect 2163 422 2183 426
rect 2187 422 2255 426
rect 2259 422 2279 426
rect 2283 422 2359 426
rect 2363 422 2375 426
rect 2379 422 2471 426
rect 2475 422 2479 426
rect 2483 422 2575 426
rect 2579 422 2607 426
rect 2611 422 2679 426
rect 2683 422 2759 426
rect 2763 422 2783 426
rect 2787 422 2903 426
rect 2907 422 2927 426
rect 2931 422 3031 426
rect 3035 422 3111 426
rect 3115 422 3167 426
rect 3171 422 3303 426
rect 3307 422 3311 426
rect 3315 422 3463 426
rect 3467 422 3495 426
rect 3499 422 3591 426
rect 3595 422 3619 426
rect 1849 421 3619 422
rect 3625 421 3626 427
rect 96 353 97 359
rect 103 358 1855 359
rect 103 354 111 358
rect 115 354 143 358
rect 147 354 231 358
rect 235 354 263 358
rect 267 354 343 358
rect 347 354 399 358
rect 403 354 455 358
rect 459 354 535 358
rect 539 354 567 358
rect 571 354 671 358
rect 675 354 767 358
rect 771 354 791 358
rect 795 354 855 358
rect 859 354 911 358
rect 915 354 943 358
rect 947 354 1023 358
rect 1027 354 1031 358
rect 1035 354 1119 358
rect 1123 354 1127 358
rect 1131 354 1207 358
rect 1211 354 1231 358
rect 1235 354 1303 358
rect 1307 354 1335 358
rect 1339 354 1439 358
rect 1443 354 1831 358
rect 1835 354 1855 358
rect 103 353 1855 354
rect 1861 353 1862 359
rect 1854 341 1855 347
rect 1861 346 3631 347
rect 1861 342 1871 346
rect 1875 342 1983 346
rect 1987 342 2071 346
rect 2075 342 2167 346
rect 2171 342 2215 346
rect 2219 342 2263 346
rect 2267 342 2295 346
rect 2299 342 2367 346
rect 2371 342 2383 346
rect 2387 342 2479 346
rect 2483 342 2591 346
rect 2595 342 2615 346
rect 2619 342 2719 346
rect 2723 342 2767 346
rect 2771 342 2847 346
rect 2851 342 2935 346
rect 2939 342 2983 346
rect 2987 342 3119 346
rect 3123 342 3255 346
rect 3259 342 3311 346
rect 3315 342 3391 346
rect 3395 342 3503 346
rect 3507 342 3511 346
rect 3515 342 3591 346
rect 3595 342 3631 346
rect 1861 341 3631 342
rect 3637 341 3638 347
rect 84 269 85 275
rect 91 274 1843 275
rect 91 270 111 274
rect 115 270 135 274
rect 139 270 247 274
rect 251 270 255 274
rect 259 270 391 274
rect 395 270 527 274
rect 531 270 543 274
rect 547 270 663 274
rect 667 270 695 274
rect 699 270 783 274
rect 787 270 847 274
rect 851 270 903 274
rect 907 270 991 274
rect 995 270 1015 274
rect 1019 270 1119 274
rect 1123 270 1223 274
rect 1227 270 1239 274
rect 1243 270 1327 274
rect 1331 270 1359 274
rect 1363 270 1431 274
rect 1435 270 1479 274
rect 1483 270 1599 274
rect 1603 270 1831 274
rect 1835 270 1843 274
rect 91 269 1843 270
rect 1849 269 1850 275
rect 1842 267 1850 269
rect 1842 261 1843 267
rect 1849 266 3619 267
rect 1849 262 1871 266
rect 1875 262 1991 266
rect 1995 262 2119 266
rect 2123 262 2207 266
rect 2211 262 2255 266
rect 2259 262 2287 266
rect 2291 262 2375 266
rect 2379 262 2391 266
rect 2395 262 2471 266
rect 2475 262 2535 266
rect 2539 262 2583 266
rect 2587 262 2679 266
rect 2683 262 2711 266
rect 2715 262 2815 266
rect 2819 262 2839 266
rect 2843 262 2951 266
rect 2955 262 2975 266
rect 2979 262 3095 266
rect 3099 262 3111 266
rect 3115 262 3239 266
rect 3243 262 3247 266
rect 3251 262 3383 266
rect 3387 262 3503 266
rect 3507 262 3591 266
rect 3595 262 3619 266
rect 1849 261 3619 262
rect 3625 261 3626 267
rect 1854 173 1855 179
rect 1861 178 3631 179
rect 1861 174 1871 178
rect 1875 174 1903 178
rect 1907 174 1983 178
rect 1987 174 1999 178
rect 2003 174 2087 178
rect 2091 174 2127 178
rect 2131 174 2215 178
rect 2219 174 2263 178
rect 2267 174 2351 178
rect 2355 174 2399 178
rect 2403 174 2487 178
rect 2491 174 2543 178
rect 2547 174 2623 178
rect 2627 174 2687 178
rect 2691 174 2743 178
rect 2747 174 2823 178
rect 2827 174 2855 178
rect 2859 174 2959 178
rect 2963 174 3063 178
rect 3067 174 3103 178
rect 3107 174 3159 178
rect 3163 174 3247 178
rect 3251 174 3343 178
rect 3347 174 3391 178
rect 3395 174 3431 178
rect 3435 174 3511 178
rect 3515 174 3591 178
rect 3595 174 3631 178
rect 1861 173 3631 174
rect 3637 173 3638 179
rect 1074 172 1080 173
rect 1358 172 1364 173
rect 1074 168 1075 172
rect 1079 168 1359 172
rect 1363 168 1364 172
rect 1074 167 1080 168
rect 1358 167 1364 168
rect 96 157 97 163
rect 103 162 1855 163
rect 103 158 111 162
rect 115 158 143 162
rect 147 158 223 162
rect 227 158 255 162
rect 259 158 303 162
rect 307 158 383 162
rect 387 158 399 162
rect 403 158 463 162
rect 467 158 543 162
rect 547 158 551 162
rect 555 158 623 162
rect 627 158 703 162
rect 707 158 783 162
rect 787 158 855 162
rect 859 158 863 162
rect 867 158 943 162
rect 947 158 999 162
rect 1003 158 1023 162
rect 1027 158 1103 162
rect 1107 158 1127 162
rect 1131 158 1183 162
rect 1187 158 1247 162
rect 1251 158 1263 162
rect 1267 158 1343 162
rect 1347 158 1367 162
rect 1371 158 1423 162
rect 1427 158 1487 162
rect 1491 158 1511 162
rect 1515 158 1591 162
rect 1595 158 1607 162
rect 1611 158 1671 162
rect 1675 158 1751 162
rect 1755 158 1831 162
rect 1835 158 1855 162
rect 103 157 1855 158
rect 1861 157 1862 163
rect 1842 97 1843 103
rect 1849 102 3619 103
rect 1849 98 1871 102
rect 1875 98 1895 102
rect 1899 98 1975 102
rect 1979 98 2079 102
rect 2083 98 2207 102
rect 2211 98 2343 102
rect 2347 98 2479 102
rect 2483 98 2615 102
rect 2619 98 2735 102
rect 2739 98 2847 102
rect 2851 98 2951 102
rect 2955 98 3055 102
rect 3059 98 3151 102
rect 3155 98 3239 102
rect 3243 98 3335 102
rect 3339 98 3423 102
rect 3427 98 3503 102
rect 3507 98 3591 102
rect 3595 98 3619 102
rect 1849 97 3619 98
rect 3625 97 3626 103
rect 84 81 85 87
rect 91 86 1843 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 215 86
rect 219 82 295 86
rect 299 82 375 86
rect 379 82 455 86
rect 459 82 535 86
rect 539 82 615 86
rect 619 82 695 86
rect 699 82 775 86
rect 779 82 855 86
rect 859 82 935 86
rect 939 82 1015 86
rect 1019 82 1095 86
rect 1099 82 1175 86
rect 1179 82 1255 86
rect 1259 82 1335 86
rect 1339 82 1415 86
rect 1419 82 1503 86
rect 1507 82 1583 86
rect 1587 82 1663 86
rect 1667 82 1743 86
rect 1747 82 1831 86
rect 1835 82 1843 86
rect 91 81 1843 82
rect 1849 81 1850 87
<< m5c >>
rect 85 3665 91 3671
rect 1843 3665 1849 3671
rect 1855 3597 1861 3603
rect 3631 3597 3637 3603
rect 97 3589 103 3595
rect 1855 3589 1861 3595
rect 1843 3521 1849 3527
rect 3619 3521 3625 3527
rect 85 3513 91 3519
rect 1843 3513 1849 3519
rect 97 3437 103 3443
rect 1855 3437 1861 3443
rect 85 3361 91 3367
rect 1843 3361 1849 3367
rect 97 3281 103 3287
rect 1855 3281 1861 3287
rect 1855 3269 1861 3275
rect 3631 3269 3637 3275
rect 85 3205 91 3211
rect 1843 3205 1849 3211
rect 1843 3189 1849 3195
rect 3619 3189 3625 3195
rect 97 3125 103 3131
rect 1855 3125 1861 3131
rect 1855 3097 1861 3103
rect 3631 3097 3637 3103
rect 85 3045 91 3051
rect 1843 3045 1849 3051
rect 1843 3013 1849 3019
rect 3619 3013 3625 3019
rect 97 2969 103 2975
rect 1855 2969 1861 2975
rect 1855 2937 1861 2943
rect 3631 2937 3637 2943
rect 85 2893 91 2899
rect 1843 2893 1849 2899
rect 1843 2853 1849 2859
rect 3619 2853 3625 2859
rect 97 2817 103 2823
rect 1855 2817 1861 2823
rect 1855 2769 1861 2775
rect 3631 2769 3637 2775
rect 85 2737 91 2743
rect 1843 2737 1849 2743
rect 1843 2693 1849 2699
rect 3619 2693 3625 2699
rect 97 2661 103 2667
rect 1855 2661 1861 2667
rect 1855 2609 1861 2615
rect 3631 2609 3637 2615
rect 85 2581 91 2587
rect 1843 2581 1849 2587
rect 1843 2525 1849 2531
rect 3619 2525 3625 2531
rect 97 2501 103 2507
rect 1855 2501 1861 2507
rect 1855 2445 1861 2451
rect 3631 2445 3637 2451
rect 85 2417 91 2423
rect 1843 2417 1849 2423
rect 1843 2361 1849 2367
rect 3619 2361 3625 2367
rect 97 2341 103 2347
rect 1855 2341 1861 2347
rect 1855 2285 1861 2291
rect 3631 2285 3637 2291
rect 85 2257 91 2263
rect 1843 2257 1849 2263
rect 1843 2189 1849 2195
rect 3619 2189 3625 2195
rect 97 2177 103 2183
rect 1855 2177 1861 2183
rect 85 2097 91 2103
rect 1843 2097 1849 2103
rect 1855 2101 1861 2107
rect 3631 2101 3637 2107
rect 1843 2031 1849 2037
rect 97 2021 103 2027
rect 1855 2021 1861 2027
rect 3619 2021 3625 2027
rect 1855 1945 1861 1951
rect 3631 1945 3637 1951
rect 85 1937 91 1943
rect 1843 1937 1849 1943
rect 1843 1871 1849 1877
rect 3619 1869 3625 1875
rect 97 1861 103 1867
rect 1855 1861 1861 1867
rect 85 1781 91 1787
rect 1843 1781 1849 1787
rect 1855 1781 1861 1787
rect 3631 1781 3637 1787
rect 1843 1711 1849 1717
rect 97 1701 103 1707
rect 1855 1701 1861 1707
rect 3619 1701 3625 1707
rect 85 1617 91 1623
rect 1843 1617 1849 1623
rect 1855 1621 1861 1627
rect 3631 1621 3637 1627
rect 1843 1547 1849 1553
rect 97 1537 103 1543
rect 1855 1537 1861 1543
rect 3619 1541 3625 1547
rect 85 1457 91 1463
rect 1843 1457 1849 1463
rect 1855 1461 1861 1467
rect 3631 1461 3637 1467
rect 1843 1385 1849 1391
rect 3619 1385 3625 1391
rect 97 1365 103 1371
rect 1855 1365 1861 1371
rect 1855 1297 1861 1303
rect 3631 1297 3637 1303
rect 85 1285 91 1291
rect 1843 1285 1849 1291
rect 1843 1217 1849 1223
rect 3619 1217 3625 1223
rect 97 1201 103 1207
rect 1855 1201 1861 1207
rect 1855 1133 1861 1139
rect 3631 1133 3637 1139
rect 85 1125 91 1131
rect 1843 1125 1849 1131
rect 1843 1057 1849 1063
rect 3619 1057 3625 1063
rect 97 1037 103 1043
rect 1855 1037 1861 1043
rect 1855 977 1861 983
rect 3631 977 3637 983
rect 85 949 91 955
rect 1843 949 1849 955
rect 1843 889 1849 895
rect 3619 889 3625 895
rect 97 869 103 875
rect 1855 869 1861 875
rect 1855 813 1861 819
rect 3631 813 3637 819
rect 85 781 91 787
rect 1843 781 1849 787
rect 1843 737 1849 743
rect 3619 737 3625 743
rect 97 697 103 703
rect 1855 697 1861 703
rect 1855 661 1861 667
rect 3631 661 3637 667
rect 85 613 91 619
rect 1843 613 1849 619
rect 1843 585 1849 591
rect 3619 585 3625 591
rect 97 525 103 531
rect 1855 525 1861 531
rect 1855 501 1861 507
rect 3631 501 3637 507
rect 85 441 91 447
rect 1843 441 1849 447
rect 1843 421 1849 427
rect 3619 421 3625 427
rect 97 353 103 359
rect 1855 353 1861 359
rect 1855 341 1861 347
rect 3631 341 3637 347
rect 85 269 91 275
rect 1843 269 1849 275
rect 1843 261 1849 267
rect 3619 261 3625 267
rect 1855 173 1861 179
rect 3631 173 3637 179
rect 97 157 103 163
rect 1855 157 1861 163
rect 1843 97 1849 103
rect 3619 97 3625 103
rect 85 81 91 87
rect 1843 81 1849 87
<< m5 >>
rect 84 3671 92 3672
rect 84 3665 85 3671
rect 91 3665 92 3671
rect 84 3519 92 3665
rect 84 3513 85 3519
rect 91 3513 92 3519
rect 84 3367 92 3513
rect 84 3361 85 3367
rect 91 3361 92 3367
rect 84 3211 92 3361
rect 84 3205 85 3211
rect 91 3205 92 3211
rect 84 3051 92 3205
rect 84 3045 85 3051
rect 91 3045 92 3051
rect 84 2899 92 3045
rect 84 2893 85 2899
rect 91 2893 92 2899
rect 84 2743 92 2893
rect 84 2737 85 2743
rect 91 2737 92 2743
rect 84 2587 92 2737
rect 84 2581 85 2587
rect 91 2581 92 2587
rect 84 2423 92 2581
rect 84 2417 85 2423
rect 91 2417 92 2423
rect 84 2263 92 2417
rect 84 2257 85 2263
rect 91 2257 92 2263
rect 84 2103 92 2257
rect 84 2097 85 2103
rect 91 2097 92 2103
rect 84 1943 92 2097
rect 84 1937 85 1943
rect 91 1937 92 1943
rect 84 1787 92 1937
rect 84 1781 85 1787
rect 91 1781 92 1787
rect 84 1623 92 1781
rect 84 1617 85 1623
rect 91 1617 92 1623
rect 84 1463 92 1617
rect 84 1457 85 1463
rect 91 1457 92 1463
rect 84 1291 92 1457
rect 84 1285 85 1291
rect 91 1285 92 1291
rect 84 1131 92 1285
rect 84 1125 85 1131
rect 91 1125 92 1131
rect 84 955 92 1125
rect 84 949 85 955
rect 91 949 92 955
rect 84 787 92 949
rect 84 781 85 787
rect 91 781 92 787
rect 84 619 92 781
rect 84 613 85 619
rect 91 613 92 619
rect 84 447 92 613
rect 84 441 85 447
rect 91 441 92 447
rect 84 275 92 441
rect 84 269 85 275
rect 91 269 92 275
rect 84 87 92 269
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 3595 104 3672
rect 96 3589 97 3595
rect 103 3589 104 3595
rect 96 3443 104 3589
rect 96 3437 97 3443
rect 103 3437 104 3443
rect 96 3287 104 3437
rect 96 3281 97 3287
rect 103 3281 104 3287
rect 96 3131 104 3281
rect 96 3125 97 3131
rect 103 3125 104 3131
rect 96 2975 104 3125
rect 96 2969 97 2975
rect 103 2969 104 2975
rect 96 2823 104 2969
rect 96 2817 97 2823
rect 103 2817 104 2823
rect 96 2667 104 2817
rect 96 2661 97 2667
rect 103 2661 104 2667
rect 96 2507 104 2661
rect 96 2501 97 2507
rect 103 2501 104 2507
rect 96 2347 104 2501
rect 96 2341 97 2347
rect 103 2341 104 2347
rect 96 2183 104 2341
rect 96 2177 97 2183
rect 103 2177 104 2183
rect 96 2027 104 2177
rect 96 2021 97 2027
rect 103 2021 104 2027
rect 96 1867 104 2021
rect 96 1861 97 1867
rect 103 1861 104 1867
rect 96 1707 104 1861
rect 96 1701 97 1707
rect 103 1701 104 1707
rect 96 1543 104 1701
rect 96 1537 97 1543
rect 103 1537 104 1543
rect 96 1371 104 1537
rect 96 1365 97 1371
rect 103 1365 104 1371
rect 96 1207 104 1365
rect 96 1201 97 1207
rect 103 1201 104 1207
rect 96 1043 104 1201
rect 96 1037 97 1043
rect 103 1037 104 1043
rect 96 875 104 1037
rect 96 869 97 875
rect 103 869 104 875
rect 96 703 104 869
rect 96 697 97 703
rect 103 697 104 703
rect 96 531 104 697
rect 96 525 97 531
rect 103 525 104 531
rect 96 359 104 525
rect 96 353 97 359
rect 103 353 104 359
rect 96 163 104 353
rect 96 157 97 163
rect 103 157 104 163
rect 96 72 104 157
rect 1842 3671 1850 3672
rect 1842 3665 1843 3671
rect 1849 3665 1850 3671
rect 1842 3527 1850 3665
rect 1842 3521 1843 3527
rect 1849 3521 1850 3527
rect 1842 3519 1850 3521
rect 1842 3513 1843 3519
rect 1849 3513 1850 3519
rect 1842 3367 1850 3513
rect 1842 3361 1843 3367
rect 1849 3361 1850 3367
rect 1842 3211 1850 3361
rect 1842 3205 1843 3211
rect 1849 3205 1850 3211
rect 1842 3195 1850 3205
rect 1842 3189 1843 3195
rect 1849 3189 1850 3195
rect 1842 3051 1850 3189
rect 1842 3045 1843 3051
rect 1849 3045 1850 3051
rect 1842 3019 1850 3045
rect 1842 3013 1843 3019
rect 1849 3013 1850 3019
rect 1842 2899 1850 3013
rect 1842 2893 1843 2899
rect 1849 2893 1850 2899
rect 1842 2859 1850 2893
rect 1842 2853 1843 2859
rect 1849 2853 1850 2859
rect 1842 2743 1850 2853
rect 1842 2737 1843 2743
rect 1849 2737 1850 2743
rect 1842 2699 1850 2737
rect 1842 2693 1843 2699
rect 1849 2693 1850 2699
rect 1842 2587 1850 2693
rect 1842 2581 1843 2587
rect 1849 2581 1850 2587
rect 1842 2531 1850 2581
rect 1842 2525 1843 2531
rect 1849 2525 1850 2531
rect 1842 2423 1850 2525
rect 1842 2417 1843 2423
rect 1849 2417 1850 2423
rect 1842 2367 1850 2417
rect 1842 2361 1843 2367
rect 1849 2361 1850 2367
rect 1842 2263 1850 2361
rect 1842 2257 1843 2263
rect 1849 2257 1850 2263
rect 1842 2195 1850 2257
rect 1842 2189 1843 2195
rect 1849 2189 1850 2195
rect 1842 2103 1850 2189
rect 1842 2097 1843 2103
rect 1849 2097 1850 2103
rect 1842 2037 1850 2097
rect 1842 2031 1843 2037
rect 1849 2031 1850 2037
rect 1842 1943 1850 2031
rect 1842 1937 1843 1943
rect 1849 1937 1850 1943
rect 1842 1877 1850 1937
rect 1842 1871 1843 1877
rect 1849 1871 1850 1877
rect 1842 1787 1850 1871
rect 1842 1781 1843 1787
rect 1849 1781 1850 1787
rect 1842 1717 1850 1781
rect 1842 1711 1843 1717
rect 1849 1711 1850 1717
rect 1842 1623 1850 1711
rect 1842 1617 1843 1623
rect 1849 1617 1850 1623
rect 1842 1553 1850 1617
rect 1842 1547 1843 1553
rect 1849 1547 1850 1553
rect 1842 1463 1850 1547
rect 1842 1457 1843 1463
rect 1849 1457 1850 1463
rect 1842 1391 1850 1457
rect 1842 1385 1843 1391
rect 1849 1385 1850 1391
rect 1842 1291 1850 1385
rect 1842 1285 1843 1291
rect 1849 1285 1850 1291
rect 1842 1223 1850 1285
rect 1842 1217 1843 1223
rect 1849 1217 1850 1223
rect 1842 1131 1850 1217
rect 1842 1125 1843 1131
rect 1849 1125 1850 1131
rect 1842 1063 1850 1125
rect 1842 1057 1843 1063
rect 1849 1057 1850 1063
rect 1842 955 1850 1057
rect 1842 949 1843 955
rect 1849 949 1850 955
rect 1842 895 1850 949
rect 1842 889 1843 895
rect 1849 889 1850 895
rect 1842 787 1850 889
rect 1842 781 1843 787
rect 1849 781 1850 787
rect 1842 743 1850 781
rect 1842 737 1843 743
rect 1849 737 1850 743
rect 1842 619 1850 737
rect 1842 613 1843 619
rect 1849 613 1850 619
rect 1842 591 1850 613
rect 1842 585 1843 591
rect 1849 585 1850 591
rect 1842 447 1850 585
rect 1842 441 1843 447
rect 1849 441 1850 447
rect 1842 427 1850 441
rect 1842 421 1843 427
rect 1849 421 1850 427
rect 1842 275 1850 421
rect 1842 269 1843 275
rect 1849 269 1850 275
rect 1842 267 1850 269
rect 1842 261 1843 267
rect 1849 261 1850 267
rect 1842 103 1850 261
rect 1842 97 1843 103
rect 1849 97 1850 103
rect 1842 87 1850 97
rect 1842 81 1843 87
rect 1849 81 1850 87
rect 1842 72 1850 81
rect 1854 3603 1862 3672
rect 1854 3597 1855 3603
rect 1861 3597 1862 3603
rect 1854 3595 1862 3597
rect 1854 3589 1855 3595
rect 1861 3589 1862 3595
rect 1854 3443 1862 3589
rect 1854 3437 1855 3443
rect 1861 3437 1862 3443
rect 1854 3287 1862 3437
rect 1854 3281 1855 3287
rect 1861 3281 1862 3287
rect 1854 3275 1862 3281
rect 1854 3269 1855 3275
rect 1861 3269 1862 3275
rect 1854 3131 1862 3269
rect 1854 3125 1855 3131
rect 1861 3125 1862 3131
rect 1854 3103 1862 3125
rect 1854 3097 1855 3103
rect 1861 3097 1862 3103
rect 1854 2975 1862 3097
rect 1854 2969 1855 2975
rect 1861 2969 1862 2975
rect 1854 2943 1862 2969
rect 1854 2937 1855 2943
rect 1861 2937 1862 2943
rect 1854 2823 1862 2937
rect 1854 2817 1855 2823
rect 1861 2817 1862 2823
rect 1854 2775 1862 2817
rect 1854 2769 1855 2775
rect 1861 2769 1862 2775
rect 1854 2667 1862 2769
rect 1854 2661 1855 2667
rect 1861 2661 1862 2667
rect 1854 2615 1862 2661
rect 1854 2609 1855 2615
rect 1861 2609 1862 2615
rect 1854 2507 1862 2609
rect 1854 2501 1855 2507
rect 1861 2501 1862 2507
rect 1854 2451 1862 2501
rect 1854 2445 1855 2451
rect 1861 2445 1862 2451
rect 1854 2347 1862 2445
rect 1854 2341 1855 2347
rect 1861 2341 1862 2347
rect 1854 2291 1862 2341
rect 1854 2285 1855 2291
rect 1861 2285 1862 2291
rect 1854 2183 1862 2285
rect 1854 2177 1855 2183
rect 1861 2177 1862 2183
rect 1854 2107 1862 2177
rect 1854 2101 1855 2107
rect 1861 2101 1862 2107
rect 1854 2027 1862 2101
rect 1854 2021 1855 2027
rect 1861 2021 1862 2027
rect 1854 1951 1862 2021
rect 1854 1945 1855 1951
rect 1861 1945 1862 1951
rect 1854 1867 1862 1945
rect 1854 1861 1855 1867
rect 1861 1861 1862 1867
rect 1854 1787 1862 1861
rect 1854 1781 1855 1787
rect 1861 1781 1862 1787
rect 1854 1707 1862 1781
rect 1854 1701 1855 1707
rect 1861 1701 1862 1707
rect 1854 1627 1862 1701
rect 1854 1621 1855 1627
rect 1861 1621 1862 1627
rect 1854 1543 1862 1621
rect 1854 1537 1855 1543
rect 1861 1537 1862 1543
rect 1854 1467 1862 1537
rect 1854 1461 1855 1467
rect 1861 1461 1862 1467
rect 1854 1371 1862 1461
rect 1854 1365 1855 1371
rect 1861 1365 1862 1371
rect 1854 1303 1862 1365
rect 1854 1297 1855 1303
rect 1861 1297 1862 1303
rect 1854 1207 1862 1297
rect 1854 1201 1855 1207
rect 1861 1201 1862 1207
rect 1854 1139 1862 1201
rect 1854 1133 1855 1139
rect 1861 1133 1862 1139
rect 1854 1043 1862 1133
rect 1854 1037 1855 1043
rect 1861 1037 1862 1043
rect 1854 983 1862 1037
rect 1854 977 1855 983
rect 1861 977 1862 983
rect 1854 875 1862 977
rect 1854 869 1855 875
rect 1861 869 1862 875
rect 1854 819 1862 869
rect 1854 813 1855 819
rect 1861 813 1862 819
rect 1854 703 1862 813
rect 1854 697 1855 703
rect 1861 697 1862 703
rect 1854 667 1862 697
rect 1854 661 1855 667
rect 1861 661 1862 667
rect 1854 531 1862 661
rect 1854 525 1855 531
rect 1861 525 1862 531
rect 1854 507 1862 525
rect 1854 501 1855 507
rect 1861 501 1862 507
rect 1854 359 1862 501
rect 1854 353 1855 359
rect 1861 353 1862 359
rect 1854 347 1862 353
rect 1854 341 1855 347
rect 1861 341 1862 347
rect 1854 179 1862 341
rect 1854 173 1855 179
rect 1861 173 1862 179
rect 1854 163 1862 173
rect 1854 157 1855 163
rect 1861 157 1862 163
rect 1854 72 1862 157
rect 3618 3527 3626 3672
rect 3618 3521 3619 3527
rect 3625 3521 3626 3527
rect 3618 3195 3626 3521
rect 3618 3189 3619 3195
rect 3625 3189 3626 3195
rect 3618 3019 3626 3189
rect 3618 3013 3619 3019
rect 3625 3013 3626 3019
rect 3618 2859 3626 3013
rect 3618 2853 3619 2859
rect 3625 2853 3626 2859
rect 3618 2699 3626 2853
rect 3618 2693 3619 2699
rect 3625 2693 3626 2699
rect 3618 2531 3626 2693
rect 3618 2525 3619 2531
rect 3625 2525 3626 2531
rect 3618 2367 3626 2525
rect 3618 2361 3619 2367
rect 3625 2361 3626 2367
rect 3618 2195 3626 2361
rect 3618 2189 3619 2195
rect 3625 2189 3626 2195
rect 3618 2027 3626 2189
rect 3618 2021 3619 2027
rect 3625 2021 3626 2027
rect 3618 1875 3626 2021
rect 3618 1869 3619 1875
rect 3625 1869 3626 1875
rect 3618 1707 3626 1869
rect 3618 1701 3619 1707
rect 3625 1701 3626 1707
rect 3618 1547 3626 1701
rect 3618 1541 3619 1547
rect 3625 1541 3626 1547
rect 3618 1391 3626 1541
rect 3618 1385 3619 1391
rect 3625 1385 3626 1391
rect 3618 1223 3626 1385
rect 3618 1217 3619 1223
rect 3625 1217 3626 1223
rect 3618 1063 3626 1217
rect 3618 1057 3619 1063
rect 3625 1057 3626 1063
rect 3618 895 3626 1057
rect 3618 889 3619 895
rect 3625 889 3626 895
rect 3618 743 3626 889
rect 3618 737 3619 743
rect 3625 737 3626 743
rect 3618 591 3626 737
rect 3618 585 3619 591
rect 3625 585 3626 591
rect 3618 427 3626 585
rect 3618 421 3619 427
rect 3625 421 3626 427
rect 3618 267 3626 421
rect 3618 261 3619 267
rect 3625 261 3626 267
rect 3618 103 3626 261
rect 3618 97 3619 103
rect 3625 97 3626 103
rect 3618 72 3626 97
rect 3630 3603 3638 3672
rect 3630 3597 3631 3603
rect 3637 3597 3638 3603
rect 3630 3275 3638 3597
rect 3630 3269 3631 3275
rect 3637 3269 3638 3275
rect 3630 3103 3638 3269
rect 3630 3097 3631 3103
rect 3637 3097 3638 3103
rect 3630 2943 3638 3097
rect 3630 2937 3631 2943
rect 3637 2937 3638 2943
rect 3630 2775 3638 2937
rect 3630 2769 3631 2775
rect 3637 2769 3638 2775
rect 3630 2615 3638 2769
rect 3630 2609 3631 2615
rect 3637 2609 3638 2615
rect 3630 2451 3638 2609
rect 3630 2445 3631 2451
rect 3637 2445 3638 2451
rect 3630 2291 3638 2445
rect 3630 2285 3631 2291
rect 3637 2285 3638 2291
rect 3630 2107 3638 2285
rect 3630 2101 3631 2107
rect 3637 2101 3638 2107
rect 3630 1951 3638 2101
rect 3630 1945 3631 1951
rect 3637 1945 3638 1951
rect 3630 1787 3638 1945
rect 3630 1781 3631 1787
rect 3637 1781 3638 1787
rect 3630 1627 3638 1781
rect 3630 1621 3631 1627
rect 3637 1621 3638 1627
rect 3630 1467 3638 1621
rect 3630 1461 3631 1467
rect 3637 1461 3638 1467
rect 3630 1303 3638 1461
rect 3630 1297 3631 1303
rect 3637 1297 3638 1303
rect 3630 1139 3638 1297
rect 3630 1133 3631 1139
rect 3637 1133 3638 1139
rect 3630 983 3638 1133
rect 3630 977 3631 983
rect 3637 977 3638 983
rect 3630 819 3638 977
rect 3630 813 3631 819
rect 3637 813 3638 819
rect 3630 667 3638 813
rect 3630 661 3631 667
rect 3637 661 3638 667
rect 3630 507 3638 661
rect 3630 501 3631 507
rect 3637 501 3638 507
rect 3630 347 3638 501
rect 3630 341 3631 347
rect 3637 341 3638 347
rect 3630 179 3638 341
rect 3630 173 3631 179
rect 3637 173 3638 179
rect 3630 72 3638 173
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__173
timestamp 1731220575
transform 1 0 3584 0 1 3544
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220575
transform 1 0 1864 0 1 3544
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220575
transform 1 0 3584 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220575
transform 1 0 1864 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220575
transform 1 0 3584 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220575
transform 1 0 1864 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220575
transform 1 0 3584 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220575
transform 1 0 1864 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220575
transform 1 0 3584 0 1 3216
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220575
transform 1 0 1864 0 1 3216
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220575
transform 1 0 3584 0 -1 3172
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220575
transform 1 0 1864 0 -1 3172
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220575
transform 1 0 3584 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220575
transform 1 0 1864 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220575
transform 1 0 3584 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220575
transform 1 0 1864 0 -1 2996
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220575
transform 1 0 3584 0 1 2884
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220575
transform 1 0 1864 0 1 2884
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220575
transform 1 0 3584 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220575
transform 1 0 1864 0 -1 2836
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220575
transform 1 0 3584 0 1 2716
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220575
transform 1 0 1864 0 1 2716
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220575
transform 1 0 3584 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220575
transform 1 0 1864 0 -1 2676
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220575
transform 1 0 3584 0 1 2556
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220575
transform 1 0 1864 0 1 2556
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220575
transform 1 0 3584 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220575
transform 1 0 1864 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220575
transform 1 0 3584 0 1 2392
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220575
transform 1 0 1864 0 1 2392
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220575
transform 1 0 3584 0 -1 2344
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220575
transform 1 0 1864 0 -1 2344
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220575
transform 1 0 3584 0 1 2232
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220575
transform 1 0 1864 0 1 2232
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220575
transform 1 0 3584 0 -1 2172
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220575
transform 1 0 1864 0 -1 2172
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220575
transform 1 0 3584 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220575
transform 1 0 1864 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220575
transform 1 0 3584 0 -1 2004
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220575
transform 1 0 1864 0 -1 2004
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220575
transform 1 0 3584 0 1 1892
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220575
transform 1 0 1864 0 1 1892
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220575
transform 1 0 3584 0 -1 1852
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220575
transform 1 0 1864 0 -1 1852
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220575
transform 1 0 3584 0 1 1728
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220575
transform 1 0 1864 0 1 1728
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220575
transform 1 0 3584 0 -1 1684
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220575
transform 1 0 1864 0 -1 1684
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220575
transform 1 0 3584 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220575
transform 1 0 1864 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220575
transform 1 0 3584 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220575
transform 1 0 1864 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220575
transform 1 0 3584 0 1 1408
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220575
transform 1 0 1864 0 1 1408
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220575
transform 1 0 3584 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220575
transform 1 0 1864 0 -1 1368
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220575
transform 1 0 3584 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220575
transform 1 0 1864 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220575
transform 1 0 3584 0 -1 1200
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220575
transform 1 0 1864 0 -1 1200
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220575
transform 1 0 3584 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220575
transform 1 0 1864 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220575
transform 1 0 3584 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220575
transform 1 0 1864 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220575
transform 1 0 3584 0 1 924
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220575
transform 1 0 1864 0 1 924
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220575
transform 1 0 3584 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220575
transform 1 0 1864 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220575
transform 1 0 3584 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220575
transform 1 0 1864 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220575
transform 1 0 3584 0 -1 720
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220575
transform 1 0 1864 0 -1 720
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220575
transform 1 0 3584 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220575
transform 1 0 1864 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220575
transform 1 0 3584 0 -1 568
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220575
transform 1 0 1864 0 -1 568
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220575
transform 1 0 3584 0 1 448
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220575
transform 1 0 1864 0 1 448
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220575
transform 1 0 3584 0 -1 404
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220575
transform 1 0 1864 0 -1 404
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220575
transform 1 0 3584 0 1 288
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220575
transform 1 0 1864 0 1 288
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220575
transform 1 0 3584 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220575
transform 1 0 1864 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220575
transform 1 0 3584 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220575
transform 1 0 1864 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220575
transform 1 0 1824 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220575
transform 1 0 104 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220575
transform 1 0 1824 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220575
transform 1 0 104 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220575
transform 1 0 1824 0 -1 3496
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220575
transform 1 0 104 0 -1 3496
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220575
transform 1 0 1824 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220575
transform 1 0 104 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220575
transform 1 0 1824 0 -1 3344
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220575
transform 1 0 104 0 -1 3344
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220575
transform 1 0 1824 0 1 3228
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220575
transform 1 0 104 0 1 3228
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220575
transform 1 0 1824 0 -1 3188
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220575
transform 1 0 104 0 -1 3188
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220575
transform 1 0 1824 0 1 3072
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220575
transform 1 0 104 0 1 3072
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220575
transform 1 0 1824 0 -1 3028
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220575
transform 1 0 104 0 -1 3028
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220575
transform 1 0 1824 0 1 2916
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220575
transform 1 0 104 0 1 2916
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220575
transform 1 0 1824 0 -1 2876
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220575
transform 1 0 104 0 -1 2876
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220575
transform 1 0 1824 0 1 2764
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220575
transform 1 0 104 0 1 2764
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220575
transform 1 0 1824 0 -1 2720
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220575
transform 1 0 104 0 -1 2720
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220575
transform 1 0 1824 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220575
transform 1 0 104 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220575
transform 1 0 1824 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220575
transform 1 0 104 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220575
transform 1 0 1824 0 1 2448
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220575
transform 1 0 104 0 1 2448
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220575
transform 1 0 1824 0 -1 2400
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220575
transform 1 0 104 0 -1 2400
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220575
transform 1 0 1824 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220575
transform 1 0 104 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220575
transform 1 0 1824 0 -1 2240
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220575
transform 1 0 104 0 -1 2240
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220575
transform 1 0 1824 0 1 2124
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220575
transform 1 0 104 0 1 2124
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220575
transform 1 0 1824 0 -1 2080
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220575
transform 1 0 104 0 -1 2080
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220575
transform 1 0 1824 0 1 1968
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220575
transform 1 0 104 0 1 1968
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220575
transform 1 0 1824 0 -1 1920
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220575
transform 1 0 104 0 -1 1920
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220575
transform 1 0 1824 0 1 1808
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220575
transform 1 0 104 0 1 1808
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220575
transform 1 0 1824 0 -1 1764
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220575
transform 1 0 104 0 -1 1764
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220575
transform 1 0 1824 0 1 1648
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220575
transform 1 0 104 0 1 1648
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220575
transform 1 0 1824 0 -1 1600
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220575
transform 1 0 104 0 -1 1600
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220575
transform 1 0 1824 0 1 1484
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220575
transform 1 0 104 0 1 1484
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220575
transform 1 0 1824 0 -1 1440
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220575
transform 1 0 104 0 -1 1440
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220575
transform 1 0 1824 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220575
transform 1 0 104 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220575
transform 1 0 1824 0 -1 1268
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220575
transform 1 0 104 0 -1 1268
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220575
transform 1 0 1824 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220575
transform 1 0 104 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220575
transform 1 0 1824 0 -1 1108
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220575
transform 1 0 104 0 -1 1108
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220575
transform 1 0 1824 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220575
transform 1 0 104 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220575
transform 1 0 1824 0 -1 932
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220575
transform 1 0 104 0 -1 932
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220575
transform 1 0 1824 0 1 816
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220575
transform 1 0 104 0 1 816
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220575
transform 1 0 1824 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220575
transform 1 0 104 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220575
transform 1 0 1824 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220575
transform 1 0 104 0 1 644
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220575
transform 1 0 1824 0 -1 596
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220575
transform 1 0 104 0 -1 596
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220575
transform 1 0 1824 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220575
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220575
transform 1 0 1824 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220575
transform 1 0 104 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220575
transform 1 0 1824 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220575
transform 1 0 104 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220575
transform 1 0 1824 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220575
transform 1 0 104 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220575
transform 1 0 1824 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220575
transform 1 0 104 0 1 104
box 7 3 12 24
use _0_0std_0_0cells_0_0LATCHINV  tst_5999_6
timestamp 1731220575
transform 1 0 3416 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5998_6
timestamp 1731220575
transform 1 0 3496 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5997_6
timestamp 1731220575
transform 1 0 3496 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5996_6
timestamp 1731220575
transform 1 0 3496 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5995_6
timestamp 1731220575
transform 1 0 3488 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5994_6
timestamp 1731220575
transform 1 0 3456 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5993_6
timestamp 1731220575
transform 1 0 3296 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5992_6
timestamp 1731220575
transform 1 0 3376 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5991_6
timestamp 1731220575
transform 1 0 3240 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5990_6
timestamp 1731220575
transform 1 0 3104 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5989_6
timestamp 1731220575
transform 1 0 3088 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5988_6
timestamp 1731220575
transform 1 0 3232 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5987_6
timestamp 1731220575
transform 1 0 3376 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5986_6
timestamp 1731220575
transform 1 0 3328 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5985_6
timestamp 1731220575
transform 1 0 3232 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5984_6
timestamp 1731220575
transform 1 0 3144 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5983_6
timestamp 1731220575
transform 1 0 3048 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5982_6
timestamp 1731220575
transform 1 0 2944 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5981_6
timestamp 1731220575
transform 1 0 2840 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5980_6
timestamp 1731220575
transform 1 0 2728 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5979_6
timestamp 1731220575
transform 1 0 2608 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5978_6
timestamp 1731220575
transform 1 0 2672 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5977_6
timestamp 1731220575
transform 1 0 2808 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5976_6
timestamp 1731220575
transform 1 0 2944 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5975_6
timestamp 1731220575
transform 1 0 2832 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5974_6
timestamp 1731220575
transform 1 0 2968 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5973_6
timestamp 1731220575
transform 1 0 3104 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5972_6
timestamp 1731220575
transform 1 0 2920 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5971_6
timestamp 1731220575
transform 1 0 2752 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5970_6
timestamp 1731220575
transform 1 0 2600 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5969_6
timestamp 1731220575
transform 1 0 2464 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5968_6
timestamp 1731220575
transform 1 0 2568 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5967_6
timestamp 1731220575
transform 1 0 2672 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5966_6
timestamp 1731220575
transform 1 0 2952 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5965_6
timestamp 1731220575
transform 1 0 2808 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5964_6
timestamp 1731220575
transform 1 0 2720 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5963_6
timestamp 1731220575
transform 1 0 2896 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5962_6
timestamp 1731220575
transform 1 0 2792 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5961_6
timestamp 1731220575
transform 1 0 3072 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5960_6
timestamp 1731220575
transform 1 0 3296 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5959_6
timestamp 1731220575
transform 1 0 3136 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5958_6
timestamp 1731220575
transform 1 0 3328 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5957_6
timestamp 1731220575
transform 1 0 3368 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5956_6
timestamp 1731220575
transform 1 0 3216 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5955_6
timestamp 1731220575
transform 1 0 3144 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5954_6
timestamp 1731220575
transform 1 0 3328 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5953_6
timestamp 1731220575
transform 1 0 3192 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5952_6
timestamp 1731220575
transform 1 0 3336 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5951_6
timestamp 1731220575
transform 1 0 3352 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5950_6
timestamp 1731220575
transform 1 0 3200 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5949_6
timestamp 1731220575
transform 1 0 3152 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5948_6
timestamp 1731220575
transform 1 0 3272 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5947_6
timestamp 1731220575
transform 1 0 3392 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5946_6
timestamp 1731220575
transform 1 0 3464 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5945_6
timestamp 1731220575
transform 1 0 3488 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5944_6
timestamp 1731220575
transform 1 0 3496 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5943_6
timestamp 1731220575
transform 1 0 3496 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5942_6
timestamp 1731220575
transform 1 0 3496 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5941_6
timestamp 1731220575
transform 1 0 3496 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5940_6
timestamp 1731220575
transform 1 0 3496 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5939_6
timestamp 1731220575
transform 1 0 3496 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5938_6
timestamp 1731220575
transform 1 0 3488 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5937_6
timestamp 1731220575
transform 1 0 3496 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5936_6
timestamp 1731220575
transform 1 0 3496 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5935_6
timestamp 1731220575
transform 1 0 3496 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5934_6
timestamp 1731220575
transform 1 0 3496 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5933_6
timestamp 1731220575
transform 1 0 3496 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5932_6
timestamp 1731220575
transform 1 0 3496 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5931_6
timestamp 1731220575
transform 1 0 3496 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5930_6
timestamp 1731220575
transform 1 0 3440 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5929_6
timestamp 1731220575
transform 1 0 3360 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5928_6
timestamp 1731220575
transform 1 0 3232 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5927_6
timestamp 1731220575
transform 1 0 3200 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5926_6
timestamp 1731220575
transform 1 0 3352 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5925_6
timestamp 1731220575
transform 1 0 3376 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5924_6
timestamp 1731220575
transform 1 0 3232 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5923_6
timestamp 1731220575
transform 1 0 3088 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5922_6
timestamp 1731220575
transform 1 0 2944 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5921_6
timestamp 1731220575
transform 1 0 3048 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5920_6
timestamp 1731220575
transform 1 0 3104 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5919_6
timestamp 1731220575
transform 1 0 3272 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5918_6
timestamp 1731220575
transform 1 0 3304 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5917_6
timestamp 1731220575
transform 1 0 3160 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5916_6
timestamp 1731220575
transform 1 0 3024 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5915_6
timestamp 1731220575
transform 1 0 2896 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5914_6
timestamp 1731220575
transform 1 0 2776 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5913_6
timestamp 1731220575
transform 1 0 3104 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5912_6
timestamp 1731220575
transform 1 0 2976 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5911_6
timestamp 1731220575
transform 1 0 2848 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5910_6
timestamp 1731220575
transform 1 0 2744 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5909_6
timestamp 1731220575
transform 1 0 2632 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5908_6
timestamp 1731220575
transform 1 0 2448 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5907_6
timestamp 1731220575
transform 1 0 2648 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5906_6
timestamp 1731220575
transform 1 0 2856 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5905_6
timestamp 1731220575
transform 1 0 2952 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5904_6
timestamp 1731220575
transform 1 0 2776 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5903_6
timestamp 1731220575
transform 1 0 2616 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5902_6
timestamp 1731220575
transform 1 0 2632 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5901_6
timestamp 1731220575
transform 1 0 2784 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5900_6
timestamp 1731220575
transform 1 0 2928 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5899_6
timestamp 1731220575
transform 1 0 3072 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5898_6
timestamp 1731220575
transform 1 0 2952 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5897_6
timestamp 1731220575
transform 1 0 2760 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5896_6
timestamp 1731220575
transform 1 0 2560 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5895_6
timestamp 1731220575
transform 1 0 3048 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5894_6
timestamp 1731220575
transform 1 0 2904 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5893_6
timestamp 1731220575
transform 1 0 2768 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5892_6
timestamp 1731220575
transform 1 0 2640 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5891_6
timestamp 1731220575
transform 1 0 2776 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5890_6
timestamp 1731220575
transform 1 0 2912 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5889_6
timestamp 1731220575
transform 1 0 3056 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5888_6
timestamp 1731220575
transform 1 0 3032 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5887_6
timestamp 1731220575
transform 1 0 2912 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5886_6
timestamp 1731220575
transform 1 0 2496 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5885_6
timestamp 1731220575
transform 1 0 2336 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5884_6
timestamp 1731220575
transform 1 0 2256 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5883_6
timestamp 1731220575
transform 1 0 2800 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5882_6
timestamp 1731220575
transform 1 0 2688 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5881_6
timestamp 1731220575
transform 1 0 2584 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5880_6
timestamp 1731220575
transform 1 0 2592 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5879_6
timestamp 1731220575
transform 1 0 2720 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5878_6
timestamp 1731220575
transform 1 0 3264 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5877_6
timestamp 1731220575
transform 1 0 3064 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5876_6
timestamp 1731220575
transform 1 0 2880 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5875_6
timestamp 1731220575
transform 1 0 2776 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5874_6
timestamp 1731220575
transform 1 0 2640 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5873_6
timestamp 1731220575
transform 1 0 3296 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5872_6
timestamp 1731220575
transform 1 0 3112 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5871_6
timestamp 1731220575
transform 1 0 2936 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5870_6
timestamp 1731220575
transform 1 0 2896 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5869_6
timestamp 1731220575
transform 1 0 2760 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5868_6
timestamp 1731220575
transform 1 0 2624 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5867_6
timestamp 1731220575
transform 1 0 3040 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5866_6
timestamp 1731220575
transform 1 0 3352 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5865_6
timestamp 1731220575
transform 1 0 3192 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5864_6
timestamp 1731220575
transform 1 0 3104 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5863_6
timestamp 1731220575
transform 1 0 2960 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5862_6
timestamp 1731220575
transform 1 0 2808 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5861_6
timestamp 1731220575
transform 1 0 3240 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5860_6
timestamp 1731220575
transform 1 0 3376 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5859_6
timestamp 1731220575
transform 1 0 3376 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5858_6
timestamp 1731220575
transform 1 0 3240 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5857_6
timestamp 1731220575
transform 1 0 3104 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5856_6
timestamp 1731220575
transform 1 0 2968 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5855_6
timestamp 1731220575
transform 1 0 2824 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5854_6
timestamp 1731220575
transform 1 0 2672 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5853_6
timestamp 1731220575
transform 1 0 3328 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5852_6
timestamp 1731220575
transform 1 0 3144 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5851_6
timestamp 1731220575
transform 1 0 2968 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5850_6
timestamp 1731220575
transform 1 0 2800 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5849_6
timestamp 1731220575
transform 1 0 2648 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5848_6
timestamp 1731220575
transform 1 0 2512 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5847_6
timestamp 1731220575
transform 1 0 2824 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5846_6
timestamp 1731220575
transform 1 0 2704 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5845_6
timestamp 1731220575
transform 1 0 2584 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5844_6
timestamp 1731220575
transform 1 0 2472 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5843_6
timestamp 1731220575
transform 1 0 2360 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5842_6
timestamp 1731220575
transform 1 0 2672 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5841_6
timestamp 1731220575
transform 1 0 2840 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5840_6
timestamp 1731220575
transform 1 0 3008 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5839_6
timestamp 1731220575
transform 1 0 3064 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5838_6
timestamp 1731220575
transform 1 0 2952 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5837_6
timestamp 1731220575
transform 1 0 2832 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5836_6
timestamp 1731220575
transform 1 0 2872 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5835_6
timestamp 1731220575
transform 1 0 2984 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5834_6
timestamp 1731220575
transform 1 0 3088 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5833_6
timestamp 1731220575
transform 1 0 3192 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5832_6
timestamp 1731220575
transform 1 0 3296 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5831_6
timestamp 1731220575
transform 1 0 3288 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5830_6
timestamp 1731220575
transform 1 0 3176 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5829_6
timestamp 1731220575
transform 1 0 3400 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5828_6
timestamp 1731220575
transform 1 0 3344 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5827_6
timestamp 1731220575
transform 1 0 3176 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5826_6
timestamp 1731220575
transform 1 0 3496 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5825_6
timestamp 1731220575
transform 1 0 3496 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5824_6
timestamp 1731220575
transform 1 0 3496 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5823_6
timestamp 1731220575
transform 1 0 3400 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5822_6
timestamp 1731220575
transform 1 0 3240 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5821_6
timestamp 1731220575
transform 1 0 3008 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5820_6
timestamp 1731220575
transform 1 0 3480 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5819_6
timestamp 1731220575
transform 1 0 3496 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5818_6
timestamp 1731220575
transform 1 0 3408 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5817_6
timestamp 1731220575
transform 1 0 3296 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5816_6
timestamp 1731220575
transform 1 0 3184 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5815_6
timestamp 1731220575
transform 1 0 3072 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5814_6
timestamp 1731220575
transform 1 0 2952 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5813_6
timestamp 1731220575
transform 1 0 2816 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5812_6
timestamp 1731220575
transform 1 0 2664 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5811_6
timestamp 1731220575
transform 1 0 3200 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5810_6
timestamp 1731220575
transform 1 0 3064 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5809_6
timestamp 1731220575
transform 1 0 2928 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5808_6
timestamp 1731220575
transform 1 0 2792 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5807_6
timestamp 1731220575
transform 1 0 2656 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5806_6
timestamp 1731220575
transform 1 0 3072 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5805_6
timestamp 1731220575
transform 1 0 2968 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5804_6
timestamp 1731220575
transform 1 0 2872 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5803_6
timestamp 1731220575
transform 1 0 2776 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5802_6
timestamp 1731220575
transform 1 0 2680 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5801_6
timestamp 1731220575
transform 1 0 2584 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5800_6
timestamp 1731220575
transform 1 0 2976 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5799_6
timestamp 1731220575
transform 1 0 2896 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5798_6
timestamp 1731220575
transform 1 0 2816 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5797_6
timestamp 1731220575
transform 1 0 2736 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5796_6
timestamp 1731220575
transform 1 0 2656 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5795_6
timestamp 1731220575
transform 1 0 2632 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5794_6
timestamp 1731220575
transform 1 0 2712 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5793_6
timestamp 1731220575
transform 1 0 2952 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5792_6
timestamp 1731220575
transform 1 0 2872 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5791_6
timestamp 1731220575
transform 1 0 2792 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5790_6
timestamp 1731220575
transform 1 0 2712 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5789_6
timestamp 1731220575
transform 1 0 2624 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5788_6
timestamp 1731220575
transform 1 0 2976 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5787_6
timestamp 1731220575
transform 1 0 2888 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5786_6
timestamp 1731220575
transform 1 0 2800 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5785_6
timestamp 1731220575
transform 1 0 2760 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5784_6
timestamp 1731220575
transform 1 0 2640 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5783_6
timestamp 1731220575
transform 1 0 3128 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5782_6
timestamp 1731220575
transform 1 0 3000 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5781_6
timestamp 1731220575
transform 1 0 2880 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5780_6
timestamp 1731220575
transform 1 0 2824 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5779_6
timestamp 1731220575
transform 1 0 2656 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5778_6
timestamp 1731220575
transform 1 0 3288 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5777_6
timestamp 1731220575
transform 1 0 3136 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5776_6
timestamp 1731220575
transform 1 0 2984 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5775_6
timestamp 1731220575
transform 1 0 2808 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5774_6
timestamp 1731220575
transform 1 0 2680 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5773_6
timestamp 1731220575
transform 1 0 2536 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5772_6
timestamp 1731220575
transform 1 0 2920 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5771_6
timestamp 1731220575
transform 1 0 3032 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5770_6
timestamp 1731220575
transform 1 0 3136 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5769_6
timestamp 1731220575
transform 1 0 3232 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5768_6
timestamp 1731220575
transform 1 0 3440 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5767_6
timestamp 1731220575
transform 1 0 3416 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5766_6
timestamp 1731220575
transform 1 0 3328 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5765_6
timestamp 1731220575
transform 1 0 3496 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5764_6
timestamp 1731220575
transform 1 0 3496 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5763_6
timestamp 1731220575
transform 1 0 3216 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5762_6
timestamp 1731220575
transform 1 0 3480 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5761_6
timestamp 1731220575
transform 1 0 3360 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5760_6
timestamp 1731220575
transform 1 0 3496 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5759_6
timestamp 1731220575
transform 1 0 3464 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5758_6
timestamp 1731220575
transform 1 0 3304 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5757_6
timestamp 1731220575
transform 1 0 3248 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5756_6
timestamp 1731220575
transform 1 0 3408 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5755_6
timestamp 1731220575
transform 1 0 3368 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5754_6
timestamp 1731220575
transform 1 0 3240 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5753_6
timestamp 1731220575
transform 1 0 3112 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5752_6
timestamp 1731220575
transform 1 0 3384 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5751_6
timestamp 1731220575
transform 1 0 3288 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5750_6
timestamp 1731220575
transform 1 0 3192 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5749_6
timestamp 1731220575
transform 1 0 3096 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5748_6
timestamp 1731220575
transform 1 0 3000 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5747_6
timestamp 1731220575
transform 1 0 2904 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5746_6
timestamp 1731220575
transform 1 0 2800 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5745_6
timestamp 1731220575
transform 1 0 2688 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5744_6
timestamp 1731220575
transform 1 0 2864 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5743_6
timestamp 1731220575
transform 1 0 2984 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5742_6
timestamp 1731220575
transform 1 0 2944 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5741_6
timestamp 1731220575
transform 1 0 3096 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5740_6
timestamp 1731220575
transform 1 0 3152 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5739_6
timestamp 1731220575
transform 1 0 3000 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5738_6
timestamp 1731220575
transform 1 0 2944 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5737_6
timestamp 1731220575
transform 1 0 3080 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5736_6
timestamp 1731220575
transform 1 0 3216 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5735_6
timestamp 1731220575
transform 1 0 3320 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5734_6
timestamp 1731220575
transform 1 0 3168 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5733_6
timestamp 1731220575
transform 1 0 3024 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5732_6
timestamp 1731220575
transform 1 0 2888 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5731_6
timestamp 1731220575
transform 1 0 2760 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5730_6
timestamp 1731220575
transform 1 0 2632 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5729_6
timestamp 1731220575
transform 1 0 2504 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5728_6
timestamp 1731220575
transform 1 0 2536 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5727_6
timestamp 1731220575
transform 1 0 2672 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5726_6
timestamp 1731220575
transform 1 0 2808 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5725_6
timestamp 1731220575
transform 1 0 2856 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5724_6
timestamp 1731220575
transform 1 0 2712 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5723_6
timestamp 1731220575
transform 1 0 2576 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5722_6
timestamp 1731220575
transform 1 0 2528 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5721_6
timestamp 1731220575
transform 1 0 2664 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5720_6
timestamp 1731220575
transform 1 0 2800 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5719_6
timestamp 1731220575
transform 1 0 2736 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5718_6
timestamp 1731220575
transform 1 0 2608 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5717_6
timestamp 1731220575
transform 1 0 2480 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5716_6
timestamp 1731220575
transform 1 0 2360 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5715_6
timestamp 1731220575
transform 1 0 2576 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5714_6
timestamp 1731220575
transform 1 0 2464 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5713_6
timestamp 1731220575
transform 1 0 2352 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5712_6
timestamp 1731220575
transform 1 0 2240 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5711_6
timestamp 1731220575
transform 1 0 2136 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5710_6
timestamp 1731220575
transform 1 0 2048 0 1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5709_6
timestamp 1731220575
transform 1 0 2080 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5708_6
timestamp 1731220575
transform 1 0 2160 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5707_6
timestamp 1731220575
transform 1 0 2256 0 -1 3524
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5706_6
timestamp 1731220575
transform 1 0 2184 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5705_6
timestamp 1731220575
transform 1 0 2096 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5704_6
timestamp 1731220575
transform 1 0 2288 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5703_6
timestamp 1731220575
transform 1 0 2400 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5702_6
timestamp 1731220575
transform 1 0 2448 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5701_6
timestamp 1731220575
transform 1 0 2328 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5700_6
timestamp 1731220575
transform 1 0 2216 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5699_6
timestamp 1731220575
transform 1 0 2120 0 -1 3360
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5698_6
timestamp 1731220575
transform 1 0 2120 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5697_6
timestamp 1731220575
transform 1 0 2400 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5696_6
timestamp 1731220575
transform 1 0 2264 0 1 3196
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5695_6
timestamp 1731220575
transform 1 0 2240 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5694_6
timestamp 1731220575
transform 1 0 2376 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5693_6
timestamp 1731220575
transform 1 0 2920 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5692_6
timestamp 1731220575
transform 1 0 2640 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5691_6
timestamp 1731220575
transform 1 0 2392 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5690_6
timestamp 1731220575
transform 1 0 2216 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5689_6
timestamp 1731220575
transform 1 0 2384 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5688_6
timestamp 1731220575
transform 1 0 2472 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5687_6
timestamp 1731220575
transform 1 0 2280 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5686_6
timestamp 1731220575
transform 1 0 2072 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5685_6
timestamp 1731220575
transform 1 0 2128 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5684_6
timestamp 1731220575
transform 1 0 2256 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5683_6
timestamp 1731220575
transform 1 0 2384 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5682_6
timestamp 1731220575
transform 1 0 2512 0 -1 2856
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5681_6
timestamp 1731220575
transform 1 0 2536 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5680_6
timestamp 1731220575
transform 1 0 2456 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5679_6
timestamp 1731220575
transform 1 0 2376 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5678_6
timestamp 1731220575
transform 1 0 2296 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5677_6
timestamp 1731220575
transform 1 0 2216 0 1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5676_6
timestamp 1731220575
transform 1 0 2232 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5675_6
timestamp 1731220575
transform 1 0 2312 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5674_6
timestamp 1731220575
transform 1 0 2392 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5673_6
timestamp 1731220575
transform 1 0 2472 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5672_6
timestamp 1731220575
transform 1 0 2552 0 -1 2696
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5671_6
timestamp 1731220575
transform 1 0 2576 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5670_6
timestamp 1731220575
transform 1 0 2496 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5669_6
timestamp 1731220575
transform 1 0 2416 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5668_6
timestamp 1731220575
transform 1 0 2336 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5667_6
timestamp 1731220575
transform 1 0 2256 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5666_6
timestamp 1731220575
transform 1 0 2176 0 1 2536
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5665_6
timestamp 1731220575
transform 1 0 2488 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5664_6
timestamp 1731220575
transform 1 0 2392 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5663_6
timestamp 1731220575
transform 1 0 2296 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5662_6
timestamp 1731220575
transform 1 0 2200 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5661_6
timestamp 1731220575
transform 1 0 2112 0 -1 2528
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5660_6
timestamp 1731220575
transform 1 0 2520 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5659_6
timestamp 1731220575
transform 1 0 2376 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5658_6
timestamp 1731220575
transform 1 0 2232 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5657_6
timestamp 1731220575
transform 1 0 2096 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5656_6
timestamp 1731220575
transform 1 0 1976 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5655_6
timestamp 1731220575
transform 1 0 1888 0 1 2372
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5654_6
timestamp 1731220575
transform 1 0 2504 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5653_6
timestamp 1731220575
transform 1 0 2336 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5652_6
timestamp 1731220575
transform 1 0 2168 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5651_6
timestamp 1731220575
transform 1 0 2008 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5650_6
timestamp 1731220575
transform 1 0 1888 0 -1 2364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5649_6
timestamp 1731220575
transform 1 0 1888 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5648_6
timestamp 1731220575
transform 1 0 2016 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5647_6
timestamp 1731220575
transform 1 0 2168 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5646_6
timestamp 1731220575
transform 1 0 2352 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5645_6
timestamp 1731220575
transform 1 0 2776 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5644_6
timestamp 1731220575
transform 1 0 2560 0 1 2212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5643_6
timestamp 1731220575
transform 1 0 2392 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5642_6
timestamp 1731220575
transform 1 0 2288 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5641_6
timestamp 1731220575
transform 1 0 2192 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5640_6
timestamp 1731220575
transform 1 0 2512 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5639_6
timestamp 1731220575
transform 1 0 2632 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5638_6
timestamp 1731220575
transform 1 0 2752 0 -1 2192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5637_6
timestamp 1731220575
transform 1 0 2712 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5636_6
timestamp 1731220575
transform 1 0 2592 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5635_6
timestamp 1731220575
transform 1 0 2472 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5634_6
timestamp 1731220575
transform 1 0 2360 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5633_6
timestamp 1731220575
transform 1 0 2256 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5632_6
timestamp 1731220575
transform 1 0 2160 0 1 2028
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5631_6
timestamp 1731220575
transform 1 0 2512 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5630_6
timestamp 1731220575
transform 1 0 2352 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5629_6
timestamp 1731220575
transform 1 0 2200 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5628_6
timestamp 1731220575
transform 1 0 2064 0 -1 2024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5627_6
timestamp 1731220575
transform 1 0 1992 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5626_6
timestamp 1731220575
transform 1 0 2120 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5625_6
timestamp 1731220575
transform 1 0 2240 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5624_6
timestamp 1731220575
transform 1 0 2376 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5623_6
timestamp 1731220575
transform 1 0 2240 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5622_6
timestamp 1731220575
transform 1 0 2112 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5621_6
timestamp 1731220575
transform 1 0 1736 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5620_6
timestamp 1731220575
transform 1 0 1616 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5619_6
timestamp 1731220575
transform 1 0 1472 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5618_6
timestamp 1731220575
transform 1 0 1336 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5617_6
timestamp 1731220575
transform 1 0 1616 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5616_6
timestamp 1731220575
transform 1 0 1480 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5615_6
timestamp 1731220575
transform 1 0 1344 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5614_6
timestamp 1731220575
transform 1 0 1208 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5613_6
timestamp 1731220575
transform 1 0 1472 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5612_6
timestamp 1731220575
transform 1 0 1376 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5611_6
timestamp 1731220575
transform 1 0 1280 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5610_6
timestamp 1731220575
transform 1 0 1192 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5609_6
timestamp 1731220575
transform 1 0 1096 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5608_6
timestamp 1731220575
transform 1 0 1304 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5607_6
timestamp 1731220575
transform 1 0 1096 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5606_6
timestamp 1731220575
transform 1 0 1008 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5605_6
timestamp 1731220575
transform 1 0 912 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5604_6
timestamp 1731220575
transform 1 0 808 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5603_6
timestamp 1731220575
transform 1 0 936 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5602_6
timestamp 1731220575
transform 1 0 1072 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5601_6
timestamp 1731220575
transform 1 0 1040 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5600_6
timestamp 1731220575
transform 1 0 1192 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5599_6
timestamp 1731220575
transform 1 0 1136 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5598_6
timestamp 1731220575
transform 1 0 1016 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5597_6
timestamp 1731220575
transform 1 0 888 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5596_6
timestamp 1731220575
transform 1 0 1384 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5595_6
timestamp 1731220575
transform 1 0 1256 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5594_6
timestamp 1731220575
transform 1 0 1168 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5593_6
timestamp 1731220575
transform 1 0 1304 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5592_6
timestamp 1731220575
transform 1 0 1432 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5591_6
timestamp 1731220575
transform 1 0 1560 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5590_6
timestamp 1731220575
transform 1 0 1696 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5589_6
timestamp 1731220575
transform 1 0 1736 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5588_6
timestamp 1731220575
transform 1 0 1616 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5587_6
timestamp 1731220575
transform 1 0 1488 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5586_6
timestamp 1731220575
transform 1 0 1352 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5585_6
timestamp 1731220575
transform 1 0 1216 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5584_6
timestamp 1731220575
transform 1 0 1064 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5583_6
timestamp 1731220575
transform 1 0 1456 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5582_6
timestamp 1731220575
transform 1 0 1320 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5581_6
timestamp 1731220575
transform 1 0 1192 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5580_6
timestamp 1731220575
transform 1 0 1064 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5579_6
timestamp 1731220575
transform 1 0 936 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5578_6
timestamp 1731220575
transform 1 0 1248 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5577_6
timestamp 1731220575
transform 1 0 1136 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5576_6
timestamp 1731220575
transform 1 0 1032 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5575_6
timestamp 1731220575
transform 1 0 928 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5574_6
timestamp 1731220575
transform 1 0 824 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5573_6
timestamp 1731220575
transform 1 0 712 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5572_6
timestamp 1731220575
transform 1 0 1152 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5571_6
timestamp 1731220575
transform 1 0 1008 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5570_6
timestamp 1731220575
transform 1 0 864 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5569_6
timestamp 1731220575
transform 1 0 720 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5568_6
timestamp 1731220575
transform 1 0 568 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5567_6
timestamp 1731220575
transform 1 0 752 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5566_6
timestamp 1731220575
transform 1 0 920 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5565_6
timestamp 1731220575
transform 1 0 832 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5564_6
timestamp 1731220575
transform 1 0 768 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5563_6
timestamp 1731220575
transform 1 0 640 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5562_6
timestamp 1731220575
transform 1 0 560 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5561_6
timestamp 1731220575
transform 1 0 456 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5560_6
timestamp 1731220575
transform 1 0 656 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5559_6
timestamp 1731220575
transform 1 0 696 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5558_6
timestamp 1731220575
transform 1 0 832 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5557_6
timestamp 1731220575
transform 1 0 800 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5556_6
timestamp 1731220575
transform 1 0 648 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5555_6
timestamp 1731220575
transform 1 0 552 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5554_6
timestamp 1731220575
transform 1 0 408 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5553_6
timestamp 1731220575
transform 1 0 256 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5552_6
timestamp 1731220575
transform 1 0 224 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5551_6
timestamp 1731220575
transform 1 0 344 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5550_6
timestamp 1731220575
transform 1 0 512 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5549_6
timestamp 1731220575
transform 1 0 376 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5548_6
timestamp 1731220575
transform 1 0 240 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5547_6
timestamp 1731220575
transform 1 0 296 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5546_6
timestamp 1731220575
transform 1 0 656 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5545_6
timestamp 1731220575
transform 1 0 472 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5544_6
timestamp 1731220575
transform 1 0 584 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5543_6
timestamp 1731220575
transform 1 0 416 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5542_6
timestamp 1731220575
transform 1 0 416 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5541_6
timestamp 1731220575
transform 1 0 272 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5540_6
timestamp 1731220575
transform 1 0 352 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5539_6
timestamp 1731220575
transform 1 0 472 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5538_6
timestamp 1731220575
transform 1 0 592 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5537_6
timestamp 1731220575
transform 1 0 800 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5536_6
timestamp 1731220575
transform 1 0 656 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5535_6
timestamp 1731220575
transform 1 0 512 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5534_6
timestamp 1731220575
transform 1 0 368 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5533_6
timestamp 1731220575
transform 1 0 536 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5532_6
timestamp 1731220575
transform 1 0 720 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5531_6
timestamp 1731220575
transform 1 0 896 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5530_6
timestamp 1731220575
transform 1 0 1024 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5529_6
timestamp 1731220575
transform 1 0 880 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5528_6
timestamp 1731220575
transform 1 0 728 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5527_6
timestamp 1731220575
transform 1 0 576 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5526_6
timestamp 1731220575
transform 1 0 584 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5525_6
timestamp 1731220575
transform 1 0 744 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5524_6
timestamp 1731220575
transform 1 0 888 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5523_6
timestamp 1731220575
transform 1 0 736 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5522_6
timestamp 1731220575
transform 1 0 584 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5521_6
timestamp 1731220575
transform 1 0 480 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5520_6
timestamp 1731220575
transform 1 0 640 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5519_6
timestamp 1731220575
transform 1 0 792 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5518_6
timestamp 1731220575
transform 1 0 704 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5517_6
timestamp 1731220575
transform 1 0 592 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5516_6
timestamp 1731220575
transform 1 0 480 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5515_6
timestamp 1731220575
transform 1 0 512 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5514_6
timestamp 1731220575
transform 1 0 696 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5513_6
timestamp 1731220575
transform 1 0 888 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5512_6
timestamp 1731220575
transform 1 0 808 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5511_6
timestamp 1731220575
transform 1 0 624 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5510_6
timestamp 1731220575
transform 1 0 1000 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5509_6
timestamp 1731220575
transform 1 0 992 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5508_6
timestamp 1731220575
transform 1 0 824 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5507_6
timestamp 1731220575
transform 1 0 664 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5506_6
timestamp 1731220575
transform 1 0 512 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5505_6
timestamp 1731220575
transform 1 0 376 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5504_6
timestamp 1731220575
transform 1 0 288 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5503_6
timestamp 1731220575
transform 1 0 208 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5502_6
timestamp 1731220575
transform 1 0 128 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5501_6
timestamp 1731220575
transform 1 0 176 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5500_6
timestamp 1731220575
transform 1 0 448 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5499_6
timestamp 1731220575
transform 1 0 296 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5498_6
timestamp 1731220575
transform 1 0 208 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5497_6
timestamp 1731220575
transform 1 0 352 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5496_6
timestamp 1731220575
transform 1 0 368 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5495_6
timestamp 1731220575
transform 1 0 248 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5494_6
timestamp 1731220575
transform 1 0 128 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5493_6
timestamp 1731220575
transform 1 0 160 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5492_6
timestamp 1731220575
transform 1 0 320 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5491_6
timestamp 1731220575
transform 1 0 288 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5490_6
timestamp 1731220575
transform 1 0 144 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5489_6
timestamp 1731220575
transform 1 0 432 0 1 1788
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5488_6
timestamp 1731220575
transform 1 0 416 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5487_6
timestamp 1731220575
transform 1 0 240 0 -1 1784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5486_6
timestamp 1731220575
transform 1 0 432 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5485_6
timestamp 1731220575
transform 1 0 296 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5484_6
timestamp 1731220575
transform 1 0 176 0 1 1628
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5483_6
timestamp 1731220575
transform 1 0 160 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5482_6
timestamp 1731220575
transform 1 0 344 0 -1 1620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5481_6
timestamp 1731220575
transform 1 0 232 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5480_6
timestamp 1731220575
transform 1 0 128 0 1 1464
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5479_6
timestamp 1731220575
transform 1 0 128 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5478_6
timestamp 1731220575
transform 1 0 224 0 -1 1460
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5477_6
timestamp 1731220575
transform 1 0 128 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5476_6
timestamp 1731220575
transform 1 0 128 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5475_6
timestamp 1731220575
transform 1 0 256 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5474_6
timestamp 1731220575
transform 1 0 128 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5473_6
timestamp 1731220575
transform 1 0 128 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5472_6
timestamp 1731220575
transform 1 0 128 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5471_6
timestamp 1731220575
transform 1 0 128 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5470_6
timestamp 1731220575
transform 1 0 128 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5469_6
timestamp 1731220575
transform 1 0 232 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5468_6
timestamp 1731220575
transform 1 0 504 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5467_6
timestamp 1731220575
transform 1 0 368 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5466_6
timestamp 1731220575
transform 1 0 296 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5465_6
timestamp 1731220575
transform 1 0 208 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5464_6
timestamp 1731220575
transform 1 0 128 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5463_6
timestamp 1731220575
transform 1 0 680 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5462_6
timestamp 1731220575
transform 1 0 536 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5461_6
timestamp 1731220575
transform 1 0 408 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5460_6
timestamp 1731220575
transform 1 0 408 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5459_6
timestamp 1731220575
transform 1 0 304 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5458_6
timestamp 1731220575
transform 1 0 216 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5457_6
timestamp 1731220575
transform 1 0 528 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5456_6
timestamp 1731220575
transform 1 0 664 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5455_6
timestamp 1731220575
transform 1 0 800 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5454_6
timestamp 1731220575
transform 1 0 768 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5453_6
timestamp 1731220575
transform 1 0 680 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5452_6
timestamp 1731220575
transform 1 0 600 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5451_6
timestamp 1731220575
transform 1 0 520 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5450_6
timestamp 1731220575
transform 1 0 440 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5449_6
timestamp 1731220575
transform 1 0 576 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5448_6
timestamp 1731220575
transform 1 0 496 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5447_6
timestamp 1731220575
transform 1 0 408 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5446_6
timestamp 1731220575
transform 1 0 320 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5445_6
timestamp 1731220575
transform 1 0 216 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5444_6
timestamp 1731220575
transform 1 0 328 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5443_6
timestamp 1731220575
transform 1 0 440 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5442_6
timestamp 1731220575
transform 1 0 384 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5441_6
timestamp 1731220575
transform 1 0 248 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5440_6
timestamp 1731220575
transform 1 0 128 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5439_6
timestamp 1731220575
transform 1 0 128 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5438_6
timestamp 1731220575
transform 1 0 240 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5437_6
timestamp 1731220575
transform 1 0 384 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5436_6
timestamp 1731220575
transform 1 0 288 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5435_6
timestamp 1731220575
transform 1 0 208 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5434_6
timestamp 1731220575
transform 1 0 128 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5433_6
timestamp 1731220575
transform 1 0 368 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5432_6
timestamp 1731220575
transform 1 0 448 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5431_6
timestamp 1731220575
transform 1 0 528 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5430_6
timestamp 1731220575
transform 1 0 768 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5429_6
timestamp 1731220575
transform 1 0 688 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5428_6
timestamp 1731220575
transform 1 0 608 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5427_6
timestamp 1731220575
transform 1 0 536 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5426_6
timestamp 1731220575
transform 1 0 688 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5425_6
timestamp 1731220575
transform 1 0 840 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5424_6
timestamp 1731220575
transform 1 0 776 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5423_6
timestamp 1731220575
transform 1 0 656 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5422_6
timestamp 1731220575
transform 1 0 520 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5421_6
timestamp 1731220575
transform 1 0 552 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5420_6
timestamp 1731220575
transform 1 0 656 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5419_6
timestamp 1731220575
transform 1 0 752 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5418_6
timestamp 1731220575
transform 1 0 736 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5417_6
timestamp 1731220575
transform 1 0 656 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5416_6
timestamp 1731220575
transform 1 0 864 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5415_6
timestamp 1731220575
transform 1 0 952 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5414_6
timestamp 1731220575
transform 1 0 936 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5413_6
timestamp 1731220575
transform 1 0 832 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5412_6
timestamp 1731220575
transform 1 0 984 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5411_6
timestamp 1731220575
transform 1 0 1136 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5410_6
timestamp 1731220575
transform 1 0 1232 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5409_6
timestamp 1731220575
transform 1 0 1088 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5408_6
timestamp 1731220575
transform 1 0 944 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5407_6
timestamp 1731220575
transform 1 0 968 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5406_6
timestamp 1731220575
transform 1 0 1096 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5405_6
timestamp 1731220575
transform 1 0 1216 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5404_6
timestamp 1731220575
transform 1 0 1208 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5403_6
timestamp 1731220575
transform 1 0 1112 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5402_6
timestamp 1731220575
transform 1 0 1016 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5401_6
timestamp 1731220575
transform 1 0 928 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5400_6
timestamp 1731220575
transform 1 0 840 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5399_6
timestamp 1731220575
transform 1 0 752 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5398_6
timestamp 1731220575
transform 1 0 888 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5397_6
timestamp 1731220575
transform 1 0 1008 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5396_6
timestamp 1731220575
transform 1 0 1128 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5395_6
timestamp 1731220575
transform 1 0 1496 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5394_6
timestamp 1731220575
transform 1 0 1368 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5393_6
timestamp 1731220575
transform 1 0 1248 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5392_6
timestamp 1731220575
transform 1 0 1144 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5391_6
timestamp 1731220575
transform 1 0 992 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5390_6
timestamp 1731220575
transform 1 0 1280 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5389_6
timestamp 1731220575
transform 1 0 1216 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5388_6
timestamp 1731220575
transform 1 0 1072 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5387_6
timestamp 1731220575
transform 1 0 1344 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5386_6
timestamp 1731220575
transform 1 0 1304 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5385_6
timestamp 1731220575
transform 1 0 1456 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5384_6
timestamp 1731220575
transform 1 0 1608 0 1 1292
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5383_6
timestamp 1731220575
transform 1 0 1600 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5382_6
timestamp 1731220575
transform 1 0 1472 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5381_6
timestamp 1731220575
transform 1 0 1728 0 -1 1288
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5380_6
timestamp 1731220575
transform 1 0 1736 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5379_6
timestamp 1731220575
transform 1 0 1640 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5378_6
timestamp 1731220575
transform 1 0 1520 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5377_6
timestamp 1731220575
transform 1 0 1400 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5376_6
timestamp 1731220575
transform 1 0 1624 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5375_6
timestamp 1731220575
transform 1 0 1736 0 -1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5374_6
timestamp 1731220575
transform 1 0 1888 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5373_6
timestamp 1731220575
transform 1 0 1888 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5372_6
timestamp 1731220575
transform 1 0 2008 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5371_6
timestamp 1731220575
transform 1 0 2160 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5370_6
timestamp 1731220575
transform 1 0 2184 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5369_6
timestamp 1731220575
transform 1 0 2064 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5368_6
timestamp 1731220575
transform 1 0 1968 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5367_6
timestamp 1731220575
transform 1 0 1888 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5366_6
timestamp 1731220575
transform 1 0 1736 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5365_6
timestamp 1731220575
transform 1 0 1736 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5364_6
timestamp 1731220575
transform 1 0 1648 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5363_6
timestamp 1731220575
transform 1 0 1536 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5362_6
timestamp 1731220575
transform 1 0 1432 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5361_6
timestamp 1731220575
transform 1 0 1328 0 -1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5360_6
timestamp 1731220575
transform 1 0 1368 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5359_6
timestamp 1731220575
transform 1 0 1624 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5358_6
timestamp 1731220575
transform 1 0 1496 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5357_6
timestamp 1731220575
transform 1 0 1440 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5356_6
timestamp 1731220575
transform 1 0 1288 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5355_6
timestamp 1731220575
transform 1 0 1600 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5354_6
timestamp 1731220575
transform 1 0 1568 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5353_6
timestamp 1731220575
transform 1 0 1440 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5352_6
timestamp 1731220575
transform 1 0 1320 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5351_6
timestamp 1731220575
transform 1 0 1200 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5350_6
timestamp 1731220575
transform 1 0 1072 0 1 624
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5349_6
timestamp 1731220575
transform 1 0 1424 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5348_6
timestamp 1731220575
transform 1 0 1328 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5347_6
timestamp 1731220575
transform 1 0 1232 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5346_6
timestamp 1731220575
transform 1 0 1136 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5345_6
timestamp 1731220575
transform 1 0 1040 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5344_6
timestamp 1731220575
transform 1 0 1264 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5343_6
timestamp 1731220575
transform 1 0 1176 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5342_6
timestamp 1731220575
transform 1 0 1088 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5341_6
timestamp 1731220575
transform 1 0 1000 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5340_6
timestamp 1731220575
transform 1 0 912 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5339_6
timestamp 1731220575
transform 1 0 824 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5338_6
timestamp 1731220575
transform 1 0 840 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5337_6
timestamp 1731220575
transform 1 0 928 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5336_6
timestamp 1731220575
transform 1 0 1016 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5335_6
timestamp 1731220575
transform 1 0 1104 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5334_6
timestamp 1731220575
transform 1 0 1288 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5333_6
timestamp 1731220575
transform 1 0 1192 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5332_6
timestamp 1731220575
transform 1 0 1112 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5331_6
timestamp 1731220575
transform 1 0 1008 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5330_6
timestamp 1731220575
transform 1 0 896 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5329_6
timestamp 1731220575
transform 1 0 1216 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5328_6
timestamp 1731220575
transform 1 0 1424 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5327_6
timestamp 1731220575
transform 1 0 1320 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5326_6
timestamp 1731220575
transform 1 0 1232 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5325_6
timestamp 1731220575
transform 1 0 1112 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5324_6
timestamp 1731220575
transform 1 0 984 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5323_6
timestamp 1731220575
transform 1 0 1592 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5322_6
timestamp 1731220575
transform 1 0 1472 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5321_6
timestamp 1731220575
transform 1 0 1352 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5320_6
timestamp 1731220575
transform 1 0 1008 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5319_6
timestamp 1731220575
transform 1 0 928 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5318_6
timestamp 1731220575
transform 1 0 848 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5317_6
timestamp 1731220575
transform 1 0 1088 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5316_6
timestamp 1731220575
transform 1 0 1168 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5315_6
timestamp 1731220575
transform 1 0 1248 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5314_6
timestamp 1731220575
transform 1 0 1328 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5313_6
timestamp 1731220575
transform 1 0 1408 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5312_6
timestamp 1731220575
transform 1 0 1496 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5311_6
timestamp 1731220575
transform 1 0 1576 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5310_6
timestamp 1731220575
transform 1 0 1656 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5309_6
timestamp 1731220575
transform 1 0 1736 0 1 84
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5308_6
timestamp 1731220575
transform 1 0 1888 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5307_6
timestamp 1731220575
transform 1 0 1968 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5306_6
timestamp 1731220575
transform 1 0 2072 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5305_6
timestamp 1731220575
transform 1 0 2472 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5304_6
timestamp 1731220575
transform 1 0 2336 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5303_6
timestamp 1731220575
transform 1 0 2200 0 1 100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5302_6
timestamp 1731220575
transform 1 0 2112 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5301_6
timestamp 1731220575
transform 1 0 1984 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5300_6
timestamp 1731220575
transform 1 0 2248 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5299_6
timestamp 1731220575
transform 1 0 2384 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5298_6
timestamp 1731220575
transform 1 0 2528 0 -1 264
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5297_6
timestamp 1731220575
transform 1 0 2704 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5296_6
timestamp 1731220575
transform 1 0 2576 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5295_6
timestamp 1731220575
transform 1 0 2464 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5294_6
timestamp 1731220575
transform 1 0 2368 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5293_6
timestamp 1731220575
transform 1 0 2280 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5292_6
timestamp 1731220575
transform 1 0 2200 0 1 268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5291_6
timestamp 1731220575
transform 1 0 2352 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5290_6
timestamp 1731220575
transform 1 0 2248 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5289_6
timestamp 1731220575
transform 1 0 2152 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5288_6
timestamp 1731220575
transform 1 0 2056 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5287_6
timestamp 1731220575
transform 1 0 1968 0 -1 424
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5286_6
timestamp 1731220575
transform 1 0 2176 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5285_6
timestamp 1731220575
transform 1 0 2272 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5284_6
timestamp 1731220575
transform 1 0 2368 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5283_6
timestamp 1731220575
transform 1 0 2472 0 1 428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5282_6
timestamp 1731220575
transform 1 0 2688 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5281_6
timestamp 1731220575
transform 1 0 2584 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5280_6
timestamp 1731220575
transform 1 0 2496 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5279_6
timestamp 1731220575
transform 1 0 2416 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5278_6
timestamp 1731220575
transform 1 0 2336 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5277_6
timestamp 1731220575
transform 1 0 2256 0 -1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5276_6
timestamp 1731220575
transform 1 0 2592 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5275_6
timestamp 1731220575
transform 1 0 2472 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5274_6
timestamp 1731220575
transform 1 0 2360 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5273_6
timestamp 1731220575
transform 1 0 2256 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5272_6
timestamp 1731220575
transform 1 0 2160 0 1 588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5271_6
timestamp 1731220575
transform 1 0 2592 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5270_6
timestamp 1731220575
transform 1 0 2440 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5269_6
timestamp 1731220575
transform 1 0 2296 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5268_6
timestamp 1731220575
transform 1 0 2168 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5267_6
timestamp 1731220575
transform 1 0 2056 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5266_6
timestamp 1731220575
transform 1 0 1960 0 -1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5265_6
timestamp 1731220575
transform 1 0 2472 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5264_6
timestamp 1731220575
transform 1 0 2312 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5263_6
timestamp 1731220575
transform 1 0 2152 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5262_6
timestamp 1731220575
transform 1 0 2000 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5261_6
timestamp 1731220575
transform 1 0 1888 0 1 740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5260_6
timestamp 1731220575
transform 1 0 1912 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5259_6
timestamp 1731220575
transform 1 0 2088 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5258_6
timestamp 1731220575
transform 1 0 2264 0 -1 892
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5257_6
timestamp 1731220575
transform 1 0 2320 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5256_6
timestamp 1731220575
transform 1 0 2464 0 1 904
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5255_6
timestamp 1731220575
transform 1 0 2480 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5254_6
timestamp 1731220575
transform 1 0 2320 0 -1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5253_6
timestamp 1731220575
transform 1 0 2112 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5252_6
timestamp 1731220575
transform 1 0 2344 0 1 1060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5251_6
timestamp 1731220575
transform 1 0 2520 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5250_6
timestamp 1731220575
transform 1 0 2400 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5249_6
timestamp 1731220575
transform 1 0 2296 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5248_6
timestamp 1731220575
transform 1 0 2200 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5247_6
timestamp 1731220575
transform 1 0 2104 0 -1 1220
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5246_6
timestamp 1731220575
transform 1 0 2200 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5245_6
timestamp 1731220575
transform 1 0 2280 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5244_6
timestamp 1731220575
transform 1 0 2360 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5243_6
timestamp 1731220575
transform 1 0 2648 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5242_6
timestamp 1731220575
transform 1 0 2536 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5241_6
timestamp 1731220575
transform 1 0 2440 0 1 1224
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5240_6
timestamp 1731220575
transform 1 0 2416 0 -1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5239_6
timestamp 1731220575
transform 1 0 2488 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5238_6
timestamp 1731220575
transform 1 0 2408 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5237_6
timestamp 1731220575
transform 1 0 2328 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5236_6
timestamp 1731220575
transform 1 0 2248 0 1 1388
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5235_6
timestamp 1731220575
transform 1 0 2528 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5234_6
timestamp 1731220575
transform 1 0 2432 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5233_6
timestamp 1731220575
transform 1 0 2336 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5232_6
timestamp 1731220575
transform 1 0 2248 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5231_6
timestamp 1731220575
transform 1 0 2160 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5230_6
timestamp 1731220575
transform 1 0 2080 0 -1 1544
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5229_6
timestamp 1731220575
transform 1 0 2488 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5228_6
timestamp 1731220575
transform 1 0 2352 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5227_6
timestamp 1731220575
transform 1 0 2216 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5226_6
timestamp 1731220575
transform 1 0 2080 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5225_6
timestamp 1731220575
transform 1 0 1960 0 1 1548
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5224_6
timestamp 1731220575
transform 1 0 2640 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5223_6
timestamp 1731220575
transform 1 0 2464 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5222_6
timestamp 1731220575
transform 1 0 2288 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5221_6
timestamp 1731220575
transform 1 0 2128 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5220_6
timestamp 1731220575
transform 1 0 1984 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5219_6
timestamp 1731220575
transform 1 0 1888 0 -1 1704
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5218_6
timestamp 1731220575
transform 1 0 2512 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5217_6
timestamp 1731220575
transform 1 0 2344 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5216_6
timestamp 1731220575
transform 1 0 2176 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5215_6
timestamp 1731220575
transform 1 0 2016 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5214_6
timestamp 1731220575
transform 1 0 1888 0 1 1708
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5213_6
timestamp 1731220575
transform 1 0 1984 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5212_6
timestamp 1731220575
transform 1 0 1888 0 -1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5211_6
timestamp 1731220575
transform 1 0 1888 0 1 1872
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5210_6
timestamp 1731220575
transform 1 0 1736 0 -1 1940
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5209_6
timestamp 1731220575
transform 1 0 1736 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5208_6
timestamp 1731220575
transform 1 0 1656 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5207_6
timestamp 1731220575
transform 1 0 1568 0 1 1948
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5206_6
timestamp 1731220575
transform 1 0 1520 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5205_6
timestamp 1731220575
transform 1 0 1736 0 -1 2100
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5204_6
timestamp 1731220575
transform 1 0 1736 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5203_6
timestamp 1731220575
transform 1 0 1568 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5202_6
timestamp 1731220575
transform 1 0 1376 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5201_6
timestamp 1731220575
transform 1 0 1184 0 1 2104
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5200_6
timestamp 1731220575
transform 1 0 1736 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5199_6
timestamp 1731220575
transform 1 0 1600 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5198_6
timestamp 1731220575
transform 1 0 1448 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5197_6
timestamp 1731220575
transform 1 0 1304 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5196_6
timestamp 1731220575
transform 1 0 1152 0 -1 2260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5195_6
timestamp 1731220575
transform 1 0 1632 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5194_6
timestamp 1731220575
transform 1 0 1552 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5193_6
timestamp 1731220575
transform 1 0 1472 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5192_6
timestamp 1731220575
transform 1 0 1392 0 1 2268
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5191_6
timestamp 1731220575
transform 1 0 1344 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5190_6
timestamp 1731220575
transform 1 0 1432 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5189_6
timestamp 1731220575
transform 1 0 1520 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5188_6
timestamp 1731220575
transform 1 0 1456 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5187_6
timestamp 1731220575
transform 1 0 1312 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5186_6
timestamp 1731220575
transform 1 0 1248 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5185_6
timestamp 1731220575
transform 1 0 1384 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5184_6
timestamp 1731220575
transform 1 0 1520 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5183_6
timestamp 1731220575
transform 1 0 1552 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5182_6
timestamp 1731220575
transform 1 0 1376 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5181_6
timestamp 1731220575
transform 1 0 1352 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5180_6
timestamp 1731220575
transform 1 0 1512 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5179_6
timestamp 1731220575
transform 1 0 1680 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5178_6
timestamp 1731220575
transform 1 0 1720 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5177_6
timestamp 1731220575
transform 1 0 1520 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5176_6
timestamp 1731220575
transform 1 0 1488 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5175_6
timestamp 1731220575
transform 1 0 1624 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5174_6
timestamp 1731220575
transform 1 0 1736 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5173_6
timestamp 1731220575
transform 1 0 1736 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5172_6
timestamp 1731220575
transform 1 0 1888 0 1 2864
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5171_6
timestamp 1731220575
transform 1 0 1888 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5170_6
timestamp 1731220575
transform 1 0 2040 0 -1 3016
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5169_6
timestamp 1731220575
transform 1 0 2000 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5168_6
timestamp 1731220575
transform 1 0 1888 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5167_6
timestamp 1731220575
transform 1 0 2176 0 1 3024
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5166_6
timestamp 1731220575
transform 1 0 2112 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5165_6
timestamp 1731220575
transform 1 0 1984 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5164_6
timestamp 1731220575
transform 1 0 1888 0 -1 3192
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5163_6
timestamp 1731220575
transform 1 0 1736 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5162_6
timestamp 1731220575
transform 1 0 1736 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5161_6
timestamp 1731220575
transform 1 0 1624 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5160_6
timestamp 1731220575
transform 1 0 1496 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5159_6
timestamp 1731220575
transform 1 0 1368 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5158_6
timestamp 1731220575
transform 1 0 1416 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5157_6
timestamp 1731220575
transform 1 0 1576 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5156_6
timestamp 1731220575
transform 1 0 1736 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5155_6
timestamp 1731220575
transform 1 0 1696 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5154_6
timestamp 1731220575
transform 1 0 1544 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5153_6
timestamp 1731220575
transform 1 0 1400 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5152_6
timestamp 1731220575
transform 1 0 1256 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5151_6
timestamp 1731220575
transform 1 0 1304 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5150_6
timestamp 1731220575
transform 1 0 1432 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5149_6
timestamp 1731220575
transform 1 0 1560 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5148_6
timestamp 1731220575
transform 1 0 1616 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5147_6
timestamp 1731220575
transform 1 0 1512 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5146_6
timestamp 1731220575
transform 1 0 1408 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5145_6
timestamp 1731220575
transform 1 0 1312 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5144_6
timestamp 1731220575
transform 1 0 1208 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5143_6
timestamp 1731220575
transform 1 0 1096 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5142_6
timestamp 1731220575
transform 1 0 984 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5141_6
timestamp 1731220575
transform 1 0 864 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5140_6
timestamp 1731220575
transform 1 0 912 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5139_6
timestamp 1731220575
transform 1 0 1048 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5138_6
timestamp 1731220575
transform 1 0 1176 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5137_6
timestamp 1731220575
transform 1 0 1104 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5136_6
timestamp 1731220575
transform 1 0 944 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5135_6
timestamp 1731220575
transform 1 0 936 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5134_6
timestamp 1731220575
transform 1 0 1096 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5133_6
timestamp 1731220575
transform 1 0 1256 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5132_6
timestamp 1731220575
transform 1 0 1240 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5131_6
timestamp 1731220575
transform 1 0 1104 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5130_6
timestamp 1731220575
transform 1 0 968 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5129_6
timestamp 1731220575
transform 1 0 1016 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5128_6
timestamp 1731220575
transform 1 0 1184 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5127_6
timestamp 1731220575
transform 1 0 1560 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5126_6
timestamp 1731220575
transform 1 0 1368 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5125_6
timestamp 1731220575
transform 1 0 1360 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5124_6
timestamp 1731220575
transform 1 0 1272 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5123_6
timestamp 1731220575
transform 1 0 1184 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5122_6
timestamp 1731220575
transform 1 0 1096 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5121_6
timestamp 1731220575
transform 1 0 1008 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5120_6
timestamp 1731220575
transform 1 0 1080 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5119_6
timestamp 1731220575
transform 1 0 1176 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5118_6
timestamp 1731220575
transform 1 0 1272 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5117_6
timestamp 1731220575
transform 1 0 1368 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5116_6
timestamp 1731220575
transform 1 0 1464 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5115_6
timestamp 1731220575
transform 1 0 1576 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5114_6
timestamp 1731220575
transform 1 0 1400 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5113_6
timestamp 1731220575
transform 1 0 1232 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5112_6
timestamp 1731220575
transform 1 0 1072 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5111_6
timestamp 1731220575
transform 1 0 1352 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5110_6
timestamp 1731220575
transform 1 0 1216 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5109_6
timestamp 1731220575
transform 1 0 1080 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5108_6
timestamp 1731220575
transform 1 0 944 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5107_6
timestamp 1731220575
transform 1 0 944 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5106_6
timestamp 1731220575
transform 1 0 1128 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5105_6
timestamp 1731220575
transform 1 0 1320 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5104_6
timestamp 1731220575
transform 1 0 1192 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5103_6
timestamp 1731220575
transform 1 0 1032 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5102_6
timestamp 1731220575
transform 1 0 872 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5101_6
timestamp 1731220575
transform 1 0 864 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5100_6
timestamp 1731220575
transform 1 0 1032 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_599_6
timestamp 1731220575
transform 1 0 1200 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_598_6
timestamp 1731220575
transform 1 0 1112 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_597_6
timestamp 1731220575
transform 1 0 976 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_596_6
timestamp 1731220575
transform 1 0 840 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_595_6
timestamp 1731220575
transform 1 0 920 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_594_6
timestamp 1731220575
transform 1 0 1048 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_593_6
timestamp 1731220575
transform 1 0 1176 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_592_6
timestamp 1731220575
transform 1 0 1256 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_591_6
timestamp 1731220575
transform 1 0 1176 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_590_6
timestamp 1731220575
transform 1 0 1096 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_589_6
timestamp 1731220575
transform 1 0 1016 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_588_6
timestamp 1731220575
transform 1 0 936 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_587_6
timestamp 1731220575
transform 1 0 856 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_586_6
timestamp 1731220575
transform 1 0 776 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_585_6
timestamp 1731220575
transform 1 0 696 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_584_6
timestamp 1731220575
transform 1 0 616 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_583_6
timestamp 1731220575
transform 1 0 536 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_582_6
timestamp 1731220575
transform 1 0 456 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_581_6
timestamp 1731220575
transform 1 0 376 0 -1 2420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_580_6
timestamp 1731220575
transform 1 0 800 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_579_6
timestamp 1731220575
transform 1 0 688 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_578_6
timestamp 1731220575
transform 1 0 584 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_577_6
timestamp 1731220575
transform 1 0 488 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_576_6
timestamp 1731220575
transform 1 0 400 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_575_6
timestamp 1731220575
transform 1 0 320 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_574_6
timestamp 1731220575
transform 1 0 696 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_573_6
timestamp 1731220575
transform 1 0 552 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_572_6
timestamp 1731220575
transform 1 0 408 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_571_6
timestamp 1731220575
transform 1 0 272 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_570_6
timestamp 1731220575
transform 1 0 152 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_569_6
timestamp 1731220575
transform 1 0 696 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_568_6
timestamp 1731220575
transform 1 0 536 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_567_6
timestamp 1731220575
transform 1 0 384 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_566_6
timestamp 1731220575
transform 1 0 240 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_565_6
timestamp 1731220575
transform 1 0 128 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_564_6
timestamp 1731220575
transform 1 0 128 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_563_6
timestamp 1731220575
transform 1 0 240 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_562_6
timestamp 1731220575
transform 1 0 704 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_561_6
timestamp 1731220575
transform 1 0 544 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_560_6
timestamp 1731220575
transform 1 0 384 0 -1 2740
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_559_6
timestamp 1731220575
transform 1 0 288 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_558_6
timestamp 1731220575
transform 1 0 152 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_557_6
timestamp 1731220575
transform 1 0 768 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_556_6
timestamp 1731220575
transform 1 0 592 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_555_6
timestamp 1731220575
transform 1 0 432 0 1 2744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_554_6
timestamp 1731220575
transform 1 0 424 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_553_6
timestamp 1731220575
transform 1 0 304 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_552_6
timestamp 1731220575
transform 1 0 808 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_551_6
timestamp 1731220575
transform 1 0 672 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_550_6
timestamp 1731220575
transform 1 0 544 0 -1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_549_6
timestamp 1731220575
transform 1 0 456 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_548_6
timestamp 1731220575
transform 1 0 560 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_547_6
timestamp 1731220575
transform 1 0 928 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_546_6
timestamp 1731220575
transform 1 0 792 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_545_6
timestamp 1731220575
transform 1 0 672 0 1 2896
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_544_6
timestamp 1731220575
transform 1 0 616 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_543_6
timestamp 1731220575
transform 1 0 536 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_542_6
timestamp 1731220575
transform 1 0 704 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_541_6
timestamp 1731220575
transform 1 0 800 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_540_6
timestamp 1731220575
transform 1 0 896 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_539_6
timestamp 1731220575
transform 1 0 992 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_538_6
timestamp 1731220575
transform 1 0 920 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_537_6
timestamp 1731220575
transform 1 0 832 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_536_6
timestamp 1731220575
transform 1 0 744 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_535_6
timestamp 1731220575
transform 1 0 656 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_534_6
timestamp 1731220575
transform 1 0 576 0 1 3052
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_533_6
timestamp 1731220575
transform 1 0 880 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_532_6
timestamp 1731220575
transform 1 0 760 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_531_6
timestamp 1731220575
transform 1 0 656 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_530_6
timestamp 1731220575
transform 1 0 568 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_529_6
timestamp 1731220575
transform 1 0 480 0 -1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_528_6
timestamp 1731220575
transform 1 0 824 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_527_6
timestamp 1731220575
transform 1 0 688 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_526_6
timestamp 1731220575
transform 1 0 560 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_525_6
timestamp 1731220575
transform 1 0 440 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_524_6
timestamp 1731220575
transform 1 0 336 0 1 3208
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_523_6
timestamp 1731220575
transform 1 0 776 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_522_6
timestamp 1731220575
transform 1 0 616 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_521_6
timestamp 1731220575
transform 1 0 464 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_520_6
timestamp 1731220575
transform 1 0 328 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_519_6
timestamp 1731220575
transform 1 0 200 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_518_6
timestamp 1731220575
transform 1 0 776 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_517_6
timestamp 1731220575
transform 1 0 608 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_516_6
timestamp 1731220575
transform 1 0 440 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_515_6
timestamp 1731220575
transform 1 0 280 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_514_6
timestamp 1731220575
transform 1 0 136 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_513_6
timestamp 1731220575
transform 1 0 184 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_512_6
timestamp 1731220575
transform 1 0 320 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_511_6
timestamp 1731220575
transform 1 0 464 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_510_6
timestamp 1731220575
transform 1 0 616 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_59_6
timestamp 1731220575
transform 1 0 768 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_58_6
timestamp 1731220575
transform 1 0 728 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_57_6
timestamp 1731220575
transform 1 0 592 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_56_6
timestamp 1731220575
transform 1 0 456 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_55_6
timestamp 1731220575
transform 1 0 328 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_54_6
timestamp 1731220575
transform 1 0 208 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_53_6
timestamp 1731220575
transform 1 0 128 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_52_6
timestamp 1731220575
transform 1 0 128 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_51_6
timestamp 1731220575
transform 1 0 208 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_50_6
timestamp 1731220575
transform 1 0 288 0 -1 3668
box 8 4 70 72
<< end >>
