magic
tech sky130l
timestamp 1730593880
<< m1 >>
rect 240 643 244 667
rect 224 587 228 619
rect 344 295 348 319
rect 448 203 452 263
rect 680 231 684 259
<< m2c >>
rect 194 851 198 855
rect 242 851 246 855
rect 290 851 294 855
rect 338 851 342 855
rect 111 841 115 845
rect 775 841 779 845
rect 111 823 115 827
rect 775 823 779 827
rect 111 781 115 785
rect 775 781 779 785
rect 111 763 115 767
rect 775 763 779 767
rect 322 751 326 755
rect 370 751 374 755
rect 418 751 422 755
rect 466 751 470 755
rect 514 753 518 757
rect 490 743 494 747
rect 250 739 254 743
rect 298 739 302 743
rect 346 739 350 743
rect 394 739 398 743
rect 442 739 446 743
rect 538 739 542 743
rect 586 739 590 743
rect 634 739 638 743
rect 682 739 686 743
rect 730 739 734 743
rect 111 729 115 733
rect 775 729 779 733
rect 111 711 115 715
rect 775 711 779 715
rect 240 667 244 671
rect 111 661 115 665
rect 111 643 115 647
rect 775 661 779 665
rect 775 643 779 647
rect 240 639 244 643
rect 146 633 150 637
rect 202 633 206 637
rect 290 633 294 637
rect 394 631 398 635
rect 506 631 510 635
rect 626 631 630 635
rect 730 631 734 635
rect 146 623 150 627
rect 730 623 734 627
rect 194 619 198 623
rect 224 619 228 623
rect 266 619 270 623
rect 370 619 374 623
rect 490 619 494 623
rect 618 619 622 623
rect 111 609 115 613
rect 111 591 115 595
rect 775 609 779 613
rect 775 591 779 595
rect 224 583 228 587
rect 111 549 115 553
rect 775 549 779 553
rect 111 531 115 535
rect 775 531 779 535
rect 146 519 150 523
rect 194 519 198 523
rect 250 519 254 523
rect 330 519 334 523
rect 426 519 430 523
rect 530 519 534 523
rect 642 519 646 523
rect 730 519 734 523
rect 274 503 278 507
rect 730 503 734 507
rect 322 499 326 503
rect 378 499 382 503
rect 442 499 446 503
rect 506 499 510 503
rect 578 499 582 503
rect 658 499 662 503
rect 111 489 115 493
rect 775 489 779 493
rect 111 471 115 475
rect 775 471 779 475
rect 111 425 115 429
rect 775 425 779 429
rect 111 407 115 411
rect 775 407 779 411
rect 426 397 430 401
rect 474 397 478 401
rect 522 395 526 399
rect 570 395 574 399
rect 618 395 622 399
rect 666 395 670 399
rect 722 397 726 401
rect 706 387 710 391
rect 298 383 302 387
rect 346 383 350 387
rect 394 383 398 387
rect 442 383 446 387
rect 498 383 502 387
rect 562 383 566 387
rect 634 383 638 387
rect 111 373 115 377
rect 775 373 779 377
rect 111 355 115 359
rect 775 355 779 359
rect 344 319 348 323
rect 111 313 115 317
rect 111 295 115 299
rect 775 313 779 317
rect 775 295 779 299
rect 344 291 348 295
rect 146 285 150 289
rect 226 285 230 289
rect 314 285 318 289
rect 410 283 414 287
rect 506 283 510 287
rect 602 283 606 287
rect 698 285 702 289
rect 146 267 150 271
rect 730 267 734 271
rect 202 263 206 267
rect 290 263 294 267
rect 378 263 382 267
rect 448 263 452 267
rect 466 263 470 267
rect 554 263 558 267
rect 642 263 646 267
rect 111 253 115 257
rect 111 235 115 239
rect 680 259 684 263
rect 775 253 779 257
rect 775 235 779 239
rect 680 227 684 231
rect 448 199 452 203
rect 111 189 115 193
rect 775 189 779 193
rect 111 171 115 175
rect 775 171 779 175
rect 194 161 198 165
rect 282 161 286 165
rect 370 161 374 165
rect 466 161 470 165
rect 562 159 566 163
rect 658 159 662 163
rect 730 159 734 163
rect 202 143 206 147
rect 730 143 734 147
rect 250 139 254 143
rect 298 139 302 143
rect 346 139 350 143
rect 394 139 398 143
rect 442 139 446 143
rect 490 139 494 143
rect 538 139 542 143
rect 586 139 590 143
rect 634 139 638 143
rect 682 139 686 143
rect 111 129 115 133
rect 775 129 779 133
rect 111 111 115 115
rect 775 111 779 115
<< m2 >>
rect 154 857 160 858
rect 154 853 155 857
rect 159 853 160 857
rect 202 857 208 858
rect 154 852 160 853
rect 166 855 172 856
rect 166 851 167 855
rect 171 854 172 855
rect 193 855 199 856
rect 193 854 194 855
rect 171 852 194 854
rect 171 851 172 852
rect 166 850 172 851
rect 193 851 194 852
rect 198 851 199 855
rect 202 853 203 857
rect 207 853 208 857
rect 250 857 256 858
rect 202 852 208 853
rect 214 855 220 856
rect 193 850 199 851
rect 214 851 215 855
rect 219 854 220 855
rect 241 855 247 856
rect 241 854 242 855
rect 219 852 242 854
rect 219 851 220 852
rect 214 850 220 851
rect 241 851 242 852
rect 246 851 247 855
rect 250 853 251 857
rect 255 853 256 857
rect 298 857 304 858
rect 250 852 256 853
rect 262 855 268 856
rect 241 850 247 851
rect 262 851 263 855
rect 267 854 268 855
rect 289 855 295 856
rect 289 854 290 855
rect 267 852 290 854
rect 267 851 268 852
rect 262 850 268 851
rect 289 851 290 852
rect 294 851 295 855
rect 298 853 299 857
rect 303 853 304 857
rect 346 857 352 858
rect 298 852 304 853
rect 310 855 316 856
rect 289 850 295 851
rect 310 851 311 855
rect 315 854 316 855
rect 337 855 343 856
rect 337 854 338 855
rect 315 852 338 854
rect 315 851 316 852
rect 310 850 316 851
rect 337 851 338 852
rect 342 851 343 855
rect 346 853 347 857
rect 351 853 352 857
rect 346 852 352 853
rect 337 850 343 851
rect 110 845 116 846
rect 110 841 111 845
rect 115 841 116 845
rect 110 840 116 841
rect 774 845 780 846
rect 774 841 775 845
rect 779 841 780 845
rect 774 840 780 841
rect 110 827 116 828
rect 110 823 111 827
rect 115 823 116 827
rect 110 822 116 823
rect 134 827 140 828
rect 134 823 135 827
rect 139 823 140 827
rect 134 822 140 823
rect 182 827 188 828
rect 182 823 183 827
rect 187 823 188 827
rect 182 822 188 823
rect 230 827 236 828
rect 230 823 231 827
rect 235 823 236 827
rect 230 822 236 823
rect 278 827 284 828
rect 278 823 279 827
rect 283 823 284 827
rect 278 822 284 823
rect 326 827 332 828
rect 326 823 327 827
rect 331 823 332 827
rect 326 822 332 823
rect 774 827 780 828
rect 774 823 775 827
rect 779 823 780 827
rect 774 822 780 823
rect 166 819 172 820
rect 166 815 167 819
rect 171 815 172 819
rect 166 814 172 815
rect 214 819 220 820
rect 214 815 215 819
rect 219 815 220 819
rect 214 814 220 815
rect 262 819 268 820
rect 262 815 263 819
rect 267 815 268 819
rect 262 814 268 815
rect 310 819 316 820
rect 310 815 311 819
rect 315 815 316 819
rect 310 814 316 815
rect 318 819 324 820
rect 318 815 319 819
rect 323 818 324 819
rect 323 816 329 818
rect 323 815 324 816
rect 318 814 324 815
rect 342 795 348 796
rect 342 791 343 795
rect 347 791 348 795
rect 342 790 348 791
rect 390 795 396 796
rect 390 791 391 795
rect 395 791 396 795
rect 390 790 396 791
rect 438 795 444 796
rect 438 791 439 795
rect 443 791 444 795
rect 438 790 444 791
rect 486 795 492 796
rect 486 791 487 795
rect 491 791 492 795
rect 486 790 492 791
rect 494 791 500 792
rect 494 787 495 791
rect 499 790 500 791
rect 499 788 505 790
rect 499 787 500 788
rect 494 786 500 787
rect 110 785 116 786
rect 110 781 111 785
rect 115 781 116 785
rect 110 780 116 781
rect 310 785 316 786
rect 310 781 311 785
rect 315 781 316 785
rect 310 780 316 781
rect 358 785 364 786
rect 358 781 359 785
rect 363 781 364 785
rect 358 780 364 781
rect 406 785 412 786
rect 406 781 407 785
rect 411 781 412 785
rect 406 780 412 781
rect 454 785 460 786
rect 454 781 455 785
rect 459 781 460 785
rect 454 780 460 781
rect 502 785 508 786
rect 502 781 503 785
rect 507 781 508 785
rect 502 780 508 781
rect 774 785 780 786
rect 774 781 775 785
rect 779 781 780 785
rect 774 780 780 781
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 774 767 780 768
rect 110 762 116 763
rect 486 763 492 764
rect 486 759 487 763
rect 491 762 492 763
rect 774 763 775 767
rect 779 763 780 767
rect 774 762 780 763
rect 491 760 518 762
rect 491 759 492 760
rect 486 758 492 759
rect 516 758 518 760
rect 513 757 519 758
rect 318 755 327 756
rect 318 751 319 755
rect 326 751 327 755
rect 318 750 327 751
rect 330 755 336 756
rect 330 751 331 755
rect 335 751 336 755
rect 330 750 336 751
rect 342 755 348 756
rect 342 751 343 755
rect 347 754 348 755
rect 369 755 375 756
rect 369 754 370 755
rect 347 752 370 754
rect 347 751 348 752
rect 342 750 348 751
rect 369 751 370 752
rect 374 751 375 755
rect 369 750 375 751
rect 378 755 384 756
rect 378 751 379 755
rect 383 751 384 755
rect 378 750 384 751
rect 390 755 396 756
rect 390 751 391 755
rect 395 754 396 755
rect 417 755 423 756
rect 417 754 418 755
rect 395 752 418 754
rect 395 751 396 752
rect 390 750 396 751
rect 417 751 418 752
rect 422 751 423 755
rect 417 750 423 751
rect 426 755 432 756
rect 426 751 427 755
rect 431 751 432 755
rect 426 750 432 751
rect 438 755 444 756
rect 438 751 439 755
rect 443 754 444 755
rect 465 755 471 756
rect 465 754 466 755
rect 443 752 466 754
rect 443 751 444 752
rect 438 750 444 751
rect 465 751 466 752
rect 470 751 471 755
rect 465 750 471 751
rect 474 755 480 756
rect 474 751 475 755
rect 479 751 480 755
rect 513 753 514 757
rect 518 753 519 757
rect 513 752 519 753
rect 522 755 528 756
rect 474 750 480 751
rect 522 751 523 755
rect 527 751 528 755
rect 522 750 528 751
rect 486 747 495 748
rect 258 745 264 746
rect 249 743 255 744
rect 249 739 250 743
rect 254 739 255 743
rect 258 741 259 745
rect 263 741 264 745
rect 306 745 312 746
rect 258 740 264 741
rect 270 743 276 744
rect 249 738 255 739
rect 270 739 271 743
rect 275 742 276 743
rect 297 743 303 744
rect 297 742 298 743
rect 275 740 298 742
rect 275 739 276 740
rect 270 738 276 739
rect 297 739 298 740
rect 302 739 303 743
rect 306 741 307 745
rect 311 741 312 745
rect 354 745 360 746
rect 306 740 312 741
rect 318 743 324 744
rect 297 738 303 739
rect 318 739 319 743
rect 323 742 324 743
rect 345 743 351 744
rect 345 742 346 743
rect 323 740 346 742
rect 323 739 324 740
rect 318 738 324 739
rect 345 739 346 740
rect 350 739 351 743
rect 354 741 355 745
rect 359 741 360 745
rect 402 745 408 746
rect 354 740 360 741
rect 393 743 399 744
rect 345 738 351 739
rect 393 739 394 743
rect 398 739 399 743
rect 402 741 403 745
rect 407 741 408 745
rect 450 745 456 746
rect 402 740 408 741
rect 441 743 447 744
rect 393 738 399 739
rect 422 739 428 740
rect 422 738 423 739
rect 252 734 254 738
rect 396 736 423 738
rect 374 735 380 736
rect 374 734 375 735
rect 110 733 116 734
rect 110 729 111 733
rect 115 729 116 733
rect 252 732 375 734
rect 374 731 375 732
rect 379 731 380 735
rect 422 735 423 736
rect 427 735 428 739
rect 441 739 442 743
rect 446 739 447 743
rect 450 741 451 745
rect 455 741 456 745
rect 486 743 487 747
rect 494 743 495 747
rect 486 742 495 743
rect 498 745 504 746
rect 450 740 456 741
rect 498 741 499 745
rect 503 741 504 745
rect 546 745 552 746
rect 498 740 504 741
rect 534 743 543 744
rect 441 738 447 739
rect 470 739 476 740
rect 470 738 471 739
rect 444 736 471 738
rect 422 734 428 735
rect 470 735 471 736
rect 475 735 476 739
rect 534 739 535 743
rect 542 739 543 743
rect 546 741 547 745
rect 551 741 552 745
rect 594 745 600 746
rect 546 740 552 741
rect 558 743 564 744
rect 534 738 543 739
rect 558 739 559 743
rect 563 742 564 743
rect 585 743 591 744
rect 585 742 586 743
rect 563 740 586 742
rect 563 739 564 740
rect 558 738 564 739
rect 585 739 586 740
rect 590 739 591 743
rect 594 741 595 745
rect 599 741 600 745
rect 642 745 648 746
rect 594 740 600 741
rect 606 743 612 744
rect 585 738 591 739
rect 606 739 607 743
rect 611 742 612 743
rect 633 743 639 744
rect 633 742 634 743
rect 611 740 634 742
rect 611 739 612 740
rect 606 738 612 739
rect 633 739 634 740
rect 638 739 639 743
rect 642 741 643 745
rect 647 741 648 745
rect 690 745 696 746
rect 642 740 648 741
rect 654 743 660 744
rect 633 738 639 739
rect 654 739 655 743
rect 659 742 660 743
rect 681 743 687 744
rect 681 742 682 743
rect 659 740 682 742
rect 659 739 660 740
rect 654 738 660 739
rect 681 739 682 740
rect 686 739 687 743
rect 690 741 691 745
rect 695 741 696 745
rect 738 745 744 746
rect 690 740 696 741
rect 702 743 708 744
rect 681 738 687 739
rect 702 739 703 743
rect 707 742 708 743
rect 729 743 735 744
rect 729 742 730 743
rect 707 740 730 742
rect 707 739 708 740
rect 702 738 708 739
rect 729 739 730 740
rect 734 739 735 743
rect 738 741 739 745
rect 743 741 744 745
rect 738 740 744 741
rect 729 738 735 739
rect 470 734 476 735
rect 374 730 380 731
rect 774 733 780 734
rect 110 728 116 729
rect 774 729 775 733
rect 779 729 780 733
rect 774 728 780 729
rect 110 715 116 716
rect 110 711 111 715
rect 115 711 116 715
rect 110 710 116 711
rect 238 715 244 716
rect 238 711 239 715
rect 243 711 244 715
rect 238 710 244 711
rect 286 715 292 716
rect 286 711 287 715
rect 291 711 292 715
rect 286 710 292 711
rect 334 715 340 716
rect 334 711 335 715
rect 339 711 340 715
rect 334 710 340 711
rect 382 715 388 716
rect 382 711 383 715
rect 387 711 388 715
rect 382 710 388 711
rect 430 715 436 716
rect 430 711 431 715
rect 435 711 436 715
rect 430 710 436 711
rect 478 715 484 716
rect 478 711 479 715
rect 483 711 484 715
rect 478 710 484 711
rect 526 715 532 716
rect 526 711 527 715
rect 531 711 532 715
rect 526 710 532 711
rect 574 715 580 716
rect 574 711 575 715
rect 579 711 580 715
rect 574 710 580 711
rect 622 715 628 716
rect 622 711 623 715
rect 627 711 628 715
rect 622 710 628 711
rect 670 715 676 716
rect 670 711 671 715
rect 675 711 676 715
rect 670 710 676 711
rect 718 715 724 716
rect 718 711 719 715
rect 723 711 724 715
rect 718 710 724 711
rect 774 715 780 716
rect 774 711 775 715
rect 779 711 780 715
rect 774 710 780 711
rect 270 707 276 708
rect 270 703 271 707
rect 275 703 276 707
rect 270 702 276 703
rect 318 707 324 708
rect 318 703 319 707
rect 323 703 324 707
rect 318 702 324 703
rect 366 707 372 708
rect 366 703 367 707
rect 371 703 372 707
rect 366 702 372 703
rect 374 707 380 708
rect 374 703 375 707
rect 379 706 380 707
rect 422 707 428 708
rect 379 704 385 706
rect 379 703 380 704
rect 374 702 380 703
rect 422 703 423 707
rect 427 706 428 707
rect 470 707 476 708
rect 427 704 433 706
rect 427 703 428 704
rect 422 702 428 703
rect 470 703 471 707
rect 475 706 476 707
rect 558 707 564 708
rect 475 704 481 706
rect 475 703 476 704
rect 470 702 476 703
rect 558 703 559 707
rect 563 703 564 707
rect 558 702 564 703
rect 606 707 612 708
rect 606 703 607 707
rect 611 703 612 707
rect 606 702 612 703
rect 654 707 660 708
rect 654 703 655 707
rect 659 703 660 707
rect 654 702 660 703
rect 702 707 708 708
rect 702 703 703 707
rect 707 703 708 707
rect 702 702 708 703
rect 726 707 732 708
rect 726 703 727 707
rect 731 703 732 707
rect 726 702 732 703
rect 414 675 420 676
rect 126 671 132 672
rect 126 667 127 671
rect 131 670 132 671
rect 174 671 180 672
rect 131 668 137 670
rect 131 667 132 668
rect 126 666 132 667
rect 174 667 175 671
rect 179 670 180 671
rect 239 671 245 672
rect 179 668 193 670
rect 179 667 180 668
rect 174 666 180 667
rect 239 667 240 671
rect 244 670 245 671
rect 414 671 415 675
rect 419 671 420 675
rect 534 675 540 676
rect 414 670 420 671
rect 422 671 428 672
rect 244 668 281 670
rect 244 667 245 668
rect 239 666 245 667
rect 422 667 423 671
rect 427 670 428 671
rect 534 671 535 675
rect 539 674 540 675
rect 539 672 617 674
rect 539 671 540 672
rect 534 670 540 671
rect 710 671 716 672
rect 427 668 497 670
rect 427 667 428 668
rect 422 666 428 667
rect 710 667 711 671
rect 715 670 716 671
rect 715 668 721 670
rect 715 667 716 668
rect 710 666 716 667
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 110 660 116 661
rect 134 665 140 666
rect 134 661 135 665
rect 139 661 140 665
rect 134 660 140 661
rect 190 665 196 666
rect 190 661 191 665
rect 195 661 196 665
rect 190 660 196 661
rect 278 665 284 666
rect 278 661 279 665
rect 283 661 284 665
rect 278 660 284 661
rect 382 665 388 666
rect 382 661 383 665
rect 387 661 388 665
rect 382 660 388 661
rect 494 665 500 666
rect 494 661 495 665
rect 499 661 500 665
rect 494 660 500 661
rect 614 665 620 666
rect 614 661 615 665
rect 619 661 620 665
rect 614 660 620 661
rect 718 665 724 666
rect 718 661 719 665
rect 723 661 724 665
rect 718 660 724 661
rect 774 665 780 666
rect 774 661 775 665
rect 779 661 780 665
rect 774 660 780 661
rect 110 647 116 648
rect 110 643 111 647
rect 115 643 116 647
rect 774 647 780 648
rect 110 642 116 643
rect 174 643 180 644
rect 174 642 175 643
rect 147 640 175 642
rect 147 638 149 640
rect 174 639 175 640
rect 179 639 180 643
rect 239 643 245 644
rect 239 642 240 643
rect 174 638 180 639
rect 204 640 240 642
rect 204 638 206 640
rect 239 639 240 640
rect 244 639 245 643
rect 422 643 428 644
rect 422 642 423 643
rect 239 638 245 639
rect 292 640 423 642
rect 292 638 294 640
rect 422 639 423 640
rect 427 639 428 643
rect 774 643 775 647
rect 779 643 780 647
rect 774 642 780 643
rect 422 638 428 639
rect 145 637 151 638
rect 145 633 146 637
rect 150 633 151 637
rect 201 637 207 638
rect 145 632 151 633
rect 154 635 160 636
rect 154 631 155 635
rect 159 631 160 635
rect 201 633 202 637
rect 206 633 207 637
rect 289 637 295 638
rect 201 632 207 633
rect 210 635 216 636
rect 154 630 160 631
rect 210 631 211 635
rect 215 631 216 635
rect 289 633 290 637
rect 294 633 295 637
rect 289 632 295 633
rect 298 635 304 636
rect 210 630 216 631
rect 298 631 299 635
rect 303 631 304 635
rect 298 630 304 631
rect 366 635 372 636
rect 366 631 367 635
rect 371 634 372 635
rect 393 635 399 636
rect 393 634 394 635
rect 371 632 394 634
rect 371 631 372 632
rect 366 630 372 631
rect 393 631 394 632
rect 398 631 399 635
rect 393 630 399 631
rect 402 635 408 636
rect 402 631 403 635
rect 407 631 408 635
rect 402 630 408 631
rect 414 635 420 636
rect 414 631 415 635
rect 419 634 420 635
rect 505 635 511 636
rect 505 634 506 635
rect 419 632 506 634
rect 419 631 420 632
rect 414 630 420 631
rect 505 631 506 632
rect 510 631 511 635
rect 505 630 511 631
rect 514 635 520 636
rect 514 631 515 635
rect 519 631 520 635
rect 625 635 631 636
rect 514 630 520 631
rect 614 631 620 632
rect 126 627 132 628
rect 126 623 127 627
rect 131 626 132 627
rect 145 627 151 628
rect 145 626 146 627
rect 131 624 146 626
rect 131 623 132 624
rect 126 622 132 623
rect 145 623 146 624
rect 150 623 151 627
rect 614 627 615 631
rect 619 630 620 631
rect 625 631 626 635
rect 630 631 631 635
rect 625 630 631 631
rect 634 635 640 636
rect 634 631 635 635
rect 639 631 640 635
rect 634 630 640 631
rect 726 635 735 636
rect 726 631 727 635
rect 734 631 735 635
rect 726 630 735 631
rect 738 635 744 636
rect 738 631 739 635
rect 743 631 744 635
rect 738 630 744 631
rect 619 628 629 630
rect 619 627 620 628
rect 614 626 620 627
rect 710 627 716 628
rect 145 622 151 623
rect 154 625 160 626
rect 154 621 155 625
rect 159 621 160 625
rect 202 625 208 626
rect 154 620 160 621
rect 166 623 172 624
rect 166 619 167 623
rect 171 622 172 623
rect 193 623 199 624
rect 193 622 194 623
rect 171 620 194 622
rect 171 619 172 620
rect 166 618 172 619
rect 193 619 194 620
rect 198 619 199 623
rect 202 621 203 625
rect 207 621 208 625
rect 274 625 280 626
rect 202 620 208 621
rect 223 623 229 624
rect 193 618 199 619
rect 223 619 224 623
rect 228 622 229 623
rect 265 623 271 624
rect 265 622 266 623
rect 228 620 266 622
rect 228 619 229 620
rect 223 618 229 619
rect 265 619 266 620
rect 270 619 271 623
rect 274 621 275 625
rect 279 621 280 625
rect 378 625 384 626
rect 274 620 280 621
rect 286 623 292 624
rect 265 618 271 619
rect 286 619 287 623
rect 291 622 292 623
rect 369 623 375 624
rect 369 622 370 623
rect 291 620 370 622
rect 291 619 292 620
rect 286 618 292 619
rect 369 619 370 620
rect 374 619 375 623
rect 378 621 379 625
rect 383 621 384 625
rect 498 625 504 626
rect 378 620 384 621
rect 390 623 396 624
rect 369 618 375 619
rect 390 619 391 623
rect 395 622 396 623
rect 489 623 495 624
rect 489 622 490 623
rect 395 620 490 622
rect 395 619 396 620
rect 390 618 396 619
rect 489 619 490 620
rect 494 619 495 623
rect 498 621 499 625
rect 503 621 504 625
rect 626 625 632 626
rect 498 620 504 621
rect 550 623 556 624
rect 489 618 495 619
rect 550 619 551 623
rect 555 622 556 623
rect 617 623 623 624
rect 617 622 618 623
rect 555 620 618 622
rect 555 619 556 620
rect 550 618 556 619
rect 617 619 618 620
rect 622 619 623 623
rect 626 621 627 625
rect 631 621 632 625
rect 710 623 711 627
rect 715 626 716 627
rect 729 627 735 628
rect 729 626 730 627
rect 715 624 730 626
rect 715 623 716 624
rect 710 622 716 623
rect 729 623 730 624
rect 734 623 735 627
rect 729 622 735 623
rect 738 625 744 626
rect 626 620 632 621
rect 738 621 739 625
rect 743 621 744 625
rect 738 620 744 621
rect 617 618 623 619
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 110 608 116 609
rect 774 613 780 614
rect 774 609 775 613
rect 779 609 780 613
rect 774 608 780 609
rect 110 595 116 596
rect 110 591 111 595
rect 115 591 116 595
rect 110 590 116 591
rect 134 595 140 596
rect 134 591 135 595
rect 139 591 140 595
rect 134 590 140 591
rect 182 595 188 596
rect 182 591 183 595
rect 187 591 188 595
rect 182 590 188 591
rect 254 595 260 596
rect 254 591 255 595
rect 259 591 260 595
rect 254 590 260 591
rect 358 595 364 596
rect 358 591 359 595
rect 363 591 364 595
rect 358 590 364 591
rect 478 595 484 596
rect 478 591 479 595
rect 483 591 484 595
rect 478 590 484 591
rect 606 595 612 596
rect 606 591 607 595
rect 611 591 612 595
rect 606 590 612 591
rect 718 595 724 596
rect 718 591 719 595
rect 723 591 724 595
rect 718 590 724 591
rect 774 595 780 596
rect 774 591 775 595
rect 779 591 780 595
rect 774 590 780 591
rect 166 587 172 588
rect 166 583 167 587
rect 171 583 172 587
rect 223 587 229 588
rect 223 586 224 587
rect 217 584 224 586
rect 166 582 172 583
rect 223 583 224 584
rect 228 583 229 587
rect 223 582 229 583
rect 286 587 292 588
rect 286 583 287 587
rect 291 583 292 587
rect 286 582 292 583
rect 390 587 396 588
rect 390 583 391 587
rect 395 583 396 587
rect 550 587 556 588
rect 550 586 551 587
rect 513 584 551 586
rect 390 582 396 583
rect 550 583 551 584
rect 555 583 556 587
rect 550 582 556 583
rect 558 587 564 588
rect 558 583 559 587
rect 563 586 564 587
rect 726 587 732 588
rect 563 584 609 586
rect 563 583 564 584
rect 558 582 564 583
rect 726 583 727 587
rect 731 583 732 587
rect 726 582 732 583
rect 458 567 464 568
rect 458 563 459 567
rect 463 566 464 567
rect 463 564 522 566
rect 463 563 464 564
rect 458 562 464 563
rect 520 561 522 564
rect 614 563 620 564
rect 174 559 180 560
rect 174 558 175 559
rect 169 556 175 558
rect 174 555 175 556
rect 179 555 180 559
rect 230 559 236 560
rect 230 558 231 559
rect 217 556 231 558
rect 174 554 180 555
rect 230 555 231 556
rect 235 555 236 559
rect 294 559 300 560
rect 294 558 295 559
rect 273 556 295 558
rect 230 554 236 555
rect 294 555 295 556
rect 299 555 300 559
rect 406 559 412 560
rect 406 558 407 559
rect 353 556 407 558
rect 294 554 300 555
rect 406 555 407 556
rect 411 555 412 559
rect 510 559 516 560
rect 510 558 511 559
rect 449 556 511 558
rect 406 554 412 555
rect 510 555 511 556
rect 515 555 516 559
rect 614 559 615 563
rect 619 562 620 563
rect 619 560 633 562
rect 619 559 620 560
rect 614 558 620 559
rect 710 559 716 560
rect 510 554 516 555
rect 710 555 711 559
rect 715 558 716 559
rect 715 556 721 558
rect 715 555 716 556
rect 710 554 716 555
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 110 548 116 549
rect 134 553 140 554
rect 134 549 135 553
rect 139 549 140 553
rect 134 548 140 549
rect 182 553 188 554
rect 182 549 183 553
rect 187 549 188 553
rect 182 548 188 549
rect 238 553 244 554
rect 238 549 239 553
rect 243 549 244 553
rect 238 548 244 549
rect 318 553 324 554
rect 318 549 319 553
rect 323 549 324 553
rect 318 548 324 549
rect 414 553 420 554
rect 414 549 415 553
rect 419 549 420 553
rect 414 548 420 549
rect 518 553 524 554
rect 518 549 519 553
rect 523 549 524 553
rect 518 548 524 549
rect 630 553 636 554
rect 630 549 631 553
rect 635 549 636 553
rect 630 548 636 549
rect 718 553 724 554
rect 718 549 719 553
rect 723 549 724 553
rect 718 548 724 549
rect 774 553 780 554
rect 774 549 775 553
rect 779 549 780 553
rect 774 548 780 549
rect 110 535 116 536
rect 110 531 111 535
rect 115 531 116 535
rect 110 530 116 531
rect 774 535 780 536
rect 774 531 775 535
rect 779 531 780 535
rect 774 530 780 531
rect 142 523 151 524
rect 142 519 143 523
rect 150 519 151 523
rect 142 518 151 519
rect 154 523 160 524
rect 154 519 155 523
rect 159 519 160 523
rect 154 518 160 519
rect 174 523 180 524
rect 174 519 175 523
rect 179 522 180 523
rect 193 523 199 524
rect 193 522 194 523
rect 179 520 194 522
rect 179 519 180 520
rect 174 518 180 519
rect 193 519 194 520
rect 198 519 199 523
rect 193 518 199 519
rect 202 523 208 524
rect 202 519 203 523
rect 207 519 208 523
rect 202 518 208 519
rect 230 523 236 524
rect 230 519 231 523
rect 235 522 236 523
rect 249 523 255 524
rect 249 522 250 523
rect 235 520 250 522
rect 235 519 236 520
rect 230 518 236 519
rect 249 519 250 520
rect 254 519 255 523
rect 249 518 255 519
rect 258 523 264 524
rect 258 519 259 523
rect 263 519 264 523
rect 258 518 264 519
rect 294 523 300 524
rect 294 519 295 523
rect 299 522 300 523
rect 329 523 335 524
rect 329 522 330 523
rect 299 520 330 522
rect 299 519 300 520
rect 294 518 300 519
rect 329 519 330 520
rect 334 519 335 523
rect 329 518 335 519
rect 338 523 344 524
rect 338 519 339 523
rect 343 519 344 523
rect 338 518 344 519
rect 406 523 412 524
rect 406 519 407 523
rect 411 522 412 523
rect 425 523 431 524
rect 425 522 426 523
rect 411 520 426 522
rect 411 519 412 520
rect 406 518 412 519
rect 425 519 426 520
rect 430 519 431 523
rect 425 518 431 519
rect 434 523 440 524
rect 434 519 435 523
rect 439 519 440 523
rect 434 518 440 519
rect 510 523 516 524
rect 510 519 511 523
rect 515 522 516 523
rect 529 523 535 524
rect 529 522 530 523
rect 515 520 530 522
rect 515 519 516 520
rect 510 518 516 519
rect 529 519 530 520
rect 534 519 535 523
rect 529 518 535 519
rect 538 523 544 524
rect 538 519 539 523
rect 543 519 544 523
rect 538 518 544 519
rect 638 523 647 524
rect 638 519 639 523
rect 646 519 647 523
rect 638 518 647 519
rect 650 523 656 524
rect 650 519 651 523
rect 655 519 656 523
rect 650 518 656 519
rect 726 523 735 524
rect 726 519 727 523
rect 734 519 735 523
rect 726 518 735 519
rect 738 523 744 524
rect 738 519 739 523
rect 743 519 744 523
rect 738 518 744 519
rect 458 511 464 512
rect 458 510 459 511
rect 276 508 459 510
rect 273 507 279 508
rect 273 503 274 507
rect 278 503 279 507
rect 458 507 459 508
rect 463 507 464 511
rect 458 506 464 507
rect 710 507 716 508
rect 273 502 279 503
rect 282 505 288 506
rect 282 501 283 505
rect 287 501 288 505
rect 330 505 336 506
rect 282 500 288 501
rect 294 503 300 504
rect 294 499 295 503
rect 299 502 300 503
rect 321 503 327 504
rect 321 502 322 503
rect 299 500 322 502
rect 299 499 300 500
rect 294 498 300 499
rect 321 499 322 500
rect 326 499 327 503
rect 330 501 331 505
rect 335 501 336 505
rect 386 505 392 506
rect 330 500 336 501
rect 358 503 364 504
rect 321 498 327 499
rect 358 499 359 503
rect 363 502 364 503
rect 377 503 383 504
rect 377 502 378 503
rect 363 500 378 502
rect 363 499 364 500
rect 358 498 364 499
rect 377 499 378 500
rect 382 499 383 503
rect 386 501 387 505
rect 391 501 392 505
rect 450 505 456 506
rect 386 500 392 501
rect 398 503 404 504
rect 377 498 383 499
rect 398 499 399 503
rect 403 502 404 503
rect 441 503 447 504
rect 441 502 442 503
rect 403 500 442 502
rect 403 499 404 500
rect 398 498 404 499
rect 441 499 442 500
rect 446 499 447 503
rect 450 501 451 505
rect 455 501 456 505
rect 514 505 520 506
rect 450 500 456 501
rect 462 503 468 504
rect 441 498 447 499
rect 462 499 463 503
rect 467 502 468 503
rect 505 503 511 504
rect 505 502 506 503
rect 467 500 506 502
rect 467 499 468 500
rect 462 498 468 499
rect 505 499 506 500
rect 510 499 511 503
rect 514 501 515 505
rect 519 501 520 505
rect 586 505 592 506
rect 514 500 520 501
rect 526 503 532 504
rect 505 498 511 499
rect 526 499 527 503
rect 531 502 532 503
rect 577 503 583 504
rect 577 502 578 503
rect 531 500 578 502
rect 531 499 532 500
rect 526 498 532 499
rect 577 499 578 500
rect 582 499 583 503
rect 586 501 587 505
rect 591 501 592 505
rect 666 505 672 506
rect 586 500 592 501
rect 657 503 663 504
rect 577 498 583 499
rect 657 499 658 503
rect 662 499 663 503
rect 666 501 667 505
rect 671 501 672 505
rect 710 503 711 507
rect 715 506 716 507
rect 729 507 735 508
rect 729 506 730 507
rect 715 504 730 506
rect 715 503 716 504
rect 710 502 716 503
rect 729 503 730 504
rect 734 503 735 507
rect 729 502 735 503
rect 738 505 744 506
rect 666 500 672 501
rect 738 501 739 505
rect 743 501 744 505
rect 738 500 744 501
rect 657 498 663 499
rect 686 499 692 500
rect 686 498 687 499
rect 660 496 687 498
rect 686 495 687 496
rect 691 495 692 499
rect 686 494 692 495
rect 110 493 116 494
rect 110 489 111 493
rect 115 489 116 493
rect 110 488 116 489
rect 774 493 780 494
rect 774 489 775 493
rect 779 489 780 493
rect 774 488 780 489
rect 110 475 116 476
rect 110 471 111 475
rect 115 471 116 475
rect 110 470 116 471
rect 262 475 268 476
rect 262 471 263 475
rect 267 471 268 475
rect 262 470 268 471
rect 310 475 316 476
rect 310 471 311 475
rect 315 471 316 475
rect 310 470 316 471
rect 366 475 372 476
rect 366 471 367 475
rect 371 471 372 475
rect 366 470 372 471
rect 430 475 436 476
rect 430 471 431 475
rect 435 471 436 475
rect 430 470 436 471
rect 494 475 500 476
rect 494 471 495 475
rect 499 471 500 475
rect 494 470 500 471
rect 566 475 572 476
rect 566 471 567 475
rect 571 471 572 475
rect 566 470 572 471
rect 646 475 652 476
rect 646 471 647 475
rect 651 471 652 475
rect 646 470 652 471
rect 718 475 724 476
rect 718 471 719 475
rect 723 471 724 475
rect 718 470 724 471
rect 774 475 780 476
rect 774 471 775 475
rect 779 471 780 475
rect 774 470 780 471
rect 294 467 300 468
rect 294 463 295 467
rect 299 463 300 467
rect 358 467 364 468
rect 358 466 359 467
rect 345 464 359 466
rect 294 462 300 463
rect 358 463 359 464
rect 363 463 364 467
rect 358 462 364 463
rect 398 467 404 468
rect 398 463 399 467
rect 403 463 404 467
rect 398 462 404 463
rect 462 467 468 468
rect 462 463 463 467
rect 467 463 468 467
rect 462 462 468 463
rect 526 467 532 468
rect 526 463 527 467
rect 531 463 532 467
rect 526 462 532 463
rect 534 467 540 468
rect 534 463 535 467
rect 539 466 540 467
rect 638 467 644 468
rect 539 464 569 466
rect 539 463 540 464
rect 534 462 540 463
rect 638 463 639 467
rect 643 466 644 467
rect 726 467 732 468
rect 643 464 649 466
rect 643 463 644 464
rect 638 462 644 463
rect 726 463 727 467
rect 731 463 732 467
rect 726 462 732 463
rect 494 439 500 440
rect 454 435 460 436
rect 454 434 455 435
rect 449 432 455 434
rect 454 431 455 432
rect 459 431 460 435
rect 494 435 495 439
rect 499 435 500 439
rect 590 439 596 440
rect 494 434 500 435
rect 550 435 556 436
rect 550 434 551 435
rect 545 432 551 434
rect 454 430 460 431
rect 550 431 551 432
rect 555 431 556 435
rect 590 435 591 439
rect 595 435 596 439
rect 686 439 692 440
rect 590 434 596 435
rect 598 435 604 436
rect 550 430 556 431
rect 598 431 599 435
rect 603 434 604 435
rect 686 435 687 439
rect 691 435 692 439
rect 686 434 692 435
rect 702 435 708 436
rect 603 432 609 434
rect 603 431 604 432
rect 598 430 604 431
rect 702 431 703 435
rect 707 434 708 435
rect 707 432 713 434
rect 707 431 708 432
rect 702 430 708 431
rect 110 429 116 430
rect 110 425 111 429
rect 115 425 116 429
rect 110 424 116 425
rect 414 429 420 430
rect 414 425 415 429
rect 419 425 420 429
rect 414 424 420 425
rect 462 429 468 430
rect 462 425 463 429
rect 467 425 468 429
rect 462 424 468 425
rect 510 429 516 430
rect 510 425 511 429
rect 515 425 516 429
rect 510 424 516 425
rect 558 429 564 430
rect 558 425 559 429
rect 563 425 564 429
rect 558 424 564 425
rect 606 429 612 430
rect 606 425 607 429
rect 611 425 612 429
rect 606 424 612 425
rect 654 429 660 430
rect 654 425 655 429
rect 659 425 660 429
rect 654 424 660 425
rect 710 429 716 430
rect 710 425 711 429
rect 715 425 716 429
rect 710 424 716 425
rect 774 429 780 430
rect 774 425 775 429
rect 779 425 780 429
rect 774 424 780 425
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 534 411 540 412
rect 534 410 535 411
rect 110 406 116 407
rect 428 408 535 410
rect 428 402 430 408
rect 534 407 535 408
rect 539 407 540 411
rect 774 411 780 412
rect 534 406 540 407
rect 726 407 732 408
rect 726 406 727 407
rect 454 403 460 404
rect 425 401 431 402
rect 425 397 426 401
rect 430 397 431 401
rect 425 396 431 397
rect 434 399 440 400
rect 434 395 435 399
rect 439 395 440 399
rect 454 399 455 403
rect 459 402 460 403
rect 724 403 727 406
rect 731 403 732 407
rect 774 407 775 411
rect 779 407 780 411
rect 774 406 780 407
rect 724 402 732 403
rect 459 401 479 402
rect 459 400 474 401
rect 459 399 460 400
rect 454 398 460 399
rect 473 397 474 400
rect 478 397 479 401
rect 721 401 727 402
rect 473 396 479 397
rect 482 399 488 400
rect 434 394 440 395
rect 482 395 483 399
rect 487 395 488 399
rect 482 394 488 395
rect 494 399 500 400
rect 494 395 495 399
rect 499 398 500 399
rect 521 399 527 400
rect 521 398 522 399
rect 499 396 522 398
rect 499 395 500 396
rect 494 394 500 395
rect 521 395 522 396
rect 526 395 527 399
rect 521 394 527 395
rect 530 399 536 400
rect 530 395 531 399
rect 535 395 536 399
rect 530 394 536 395
rect 550 399 556 400
rect 550 395 551 399
rect 555 398 556 399
rect 569 399 575 400
rect 569 398 570 399
rect 555 396 570 398
rect 555 395 556 396
rect 550 394 556 395
rect 569 395 570 396
rect 574 395 575 399
rect 569 394 575 395
rect 578 399 584 400
rect 578 395 579 399
rect 583 395 584 399
rect 578 394 584 395
rect 590 399 596 400
rect 590 395 591 399
rect 595 398 596 399
rect 617 399 623 400
rect 617 398 618 399
rect 595 396 618 398
rect 595 395 596 396
rect 590 394 596 395
rect 617 395 618 396
rect 622 395 623 399
rect 617 394 623 395
rect 626 399 632 400
rect 626 395 627 399
rect 631 395 632 399
rect 626 394 632 395
rect 654 399 660 400
rect 654 395 655 399
rect 659 398 660 399
rect 665 399 671 400
rect 665 398 666 399
rect 659 396 666 398
rect 659 395 660 396
rect 654 394 660 395
rect 665 395 666 396
rect 670 395 671 399
rect 665 394 671 395
rect 674 399 680 400
rect 674 395 675 399
rect 679 395 680 399
rect 721 397 722 401
rect 726 397 727 401
rect 721 396 727 397
rect 730 399 736 400
rect 674 394 680 395
rect 730 395 731 399
rect 735 395 736 399
rect 730 394 736 395
rect 702 391 711 392
rect 306 389 312 390
rect 297 387 303 388
rect 297 383 298 387
rect 302 383 303 387
rect 306 385 307 389
rect 311 385 312 389
rect 354 389 360 390
rect 306 384 312 385
rect 318 387 324 388
rect 297 382 303 383
rect 318 383 319 387
rect 323 386 324 387
rect 345 387 351 388
rect 345 386 346 387
rect 323 384 346 386
rect 323 383 324 384
rect 318 382 324 383
rect 345 383 346 384
rect 350 383 351 387
rect 354 385 355 389
rect 359 385 360 389
rect 402 389 408 390
rect 354 384 360 385
rect 366 387 372 388
rect 345 382 351 383
rect 366 383 367 387
rect 371 386 372 387
rect 393 387 399 388
rect 393 386 394 387
rect 371 384 394 386
rect 371 383 372 384
rect 366 382 372 383
rect 393 383 394 384
rect 398 383 399 387
rect 402 385 403 389
rect 407 385 408 389
rect 450 389 456 390
rect 402 384 408 385
rect 441 387 447 388
rect 393 382 399 383
rect 441 383 442 387
rect 446 383 447 387
rect 450 385 451 389
rect 455 385 456 389
rect 506 389 512 390
rect 450 384 456 385
rect 497 387 503 388
rect 441 382 447 383
rect 470 383 476 384
rect 470 382 471 383
rect 300 378 302 382
rect 444 380 471 382
rect 422 379 428 380
rect 422 378 423 379
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 300 376 423 378
rect 422 375 423 376
rect 427 375 428 379
rect 470 379 471 380
rect 475 379 476 383
rect 497 383 498 387
rect 502 383 503 387
rect 506 385 507 389
rect 511 385 512 389
rect 570 389 576 390
rect 506 384 512 385
rect 561 387 567 388
rect 497 382 503 383
rect 526 383 532 384
rect 526 382 527 383
rect 500 380 527 382
rect 470 378 476 379
rect 526 379 527 380
rect 531 379 532 383
rect 561 383 562 387
rect 566 383 567 387
rect 570 385 571 389
rect 575 385 576 389
rect 642 389 648 390
rect 633 387 639 388
rect 633 386 634 387
rect 570 384 576 385
rect 632 384 634 386
rect 561 382 567 383
rect 598 383 604 384
rect 598 382 599 383
rect 564 380 599 382
rect 526 378 532 379
rect 598 379 599 380
rect 603 379 604 383
rect 598 378 604 379
rect 630 383 634 384
rect 638 383 639 387
rect 642 385 643 389
rect 647 385 648 389
rect 702 387 703 391
rect 710 387 711 391
rect 702 386 711 387
rect 714 389 720 390
rect 642 384 648 385
rect 714 385 715 389
rect 719 385 720 389
rect 714 384 720 385
rect 630 379 631 383
rect 635 382 639 383
rect 635 379 636 382
rect 630 378 636 379
rect 422 374 428 375
rect 774 377 780 378
rect 110 372 116 373
rect 774 373 775 377
rect 779 373 780 377
rect 774 372 780 373
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 286 359 292 360
rect 286 355 287 359
rect 291 355 292 359
rect 286 354 292 355
rect 334 359 340 360
rect 334 355 335 359
rect 339 355 340 359
rect 334 354 340 355
rect 382 359 388 360
rect 382 355 383 359
rect 387 355 388 359
rect 382 354 388 355
rect 430 359 436 360
rect 430 355 431 359
rect 435 355 436 359
rect 430 354 436 355
rect 486 359 492 360
rect 486 355 487 359
rect 491 355 492 359
rect 486 354 492 355
rect 550 359 556 360
rect 550 355 551 359
rect 555 355 556 359
rect 550 354 556 355
rect 622 359 628 360
rect 622 355 623 359
rect 627 355 628 359
rect 622 354 628 355
rect 694 359 700 360
rect 694 355 695 359
rect 699 355 700 359
rect 694 354 700 355
rect 774 359 780 360
rect 774 355 775 359
rect 779 355 780 359
rect 774 354 780 355
rect 318 351 324 352
rect 318 347 319 351
rect 323 347 324 351
rect 318 346 324 347
rect 366 351 372 352
rect 366 347 367 351
rect 371 347 372 351
rect 366 346 372 347
rect 406 351 412 352
rect 406 347 407 351
rect 411 347 412 351
rect 406 346 412 347
rect 422 351 428 352
rect 422 347 423 351
rect 427 350 428 351
rect 470 351 476 352
rect 427 348 433 350
rect 427 347 428 348
rect 422 346 428 347
rect 470 347 471 351
rect 475 350 476 351
rect 526 351 532 352
rect 475 348 489 350
rect 475 347 476 348
rect 470 346 476 347
rect 526 347 527 351
rect 531 350 532 351
rect 654 351 660 352
rect 531 348 553 350
rect 531 347 532 348
rect 526 346 532 347
rect 654 347 655 351
rect 659 347 660 351
rect 654 346 660 347
rect 702 351 708 352
rect 702 347 703 351
rect 707 347 708 351
rect 702 346 708 347
rect 630 327 636 328
rect 630 326 631 327
rect 625 324 631 326
rect 126 323 132 324
rect 126 319 127 323
rect 131 322 132 323
rect 182 323 188 324
rect 131 320 137 322
rect 131 319 132 320
rect 126 318 132 319
rect 182 319 183 323
rect 187 322 188 323
rect 254 323 260 324
rect 187 320 217 322
rect 187 319 188 320
rect 182 318 188 319
rect 254 319 255 323
rect 259 322 260 323
rect 343 323 349 324
rect 259 320 305 322
rect 259 319 260 320
rect 254 318 260 319
rect 343 319 344 323
rect 348 322 349 323
rect 582 323 588 324
rect 582 322 583 323
rect 348 320 401 322
rect 529 320 583 322
rect 348 319 349 320
rect 343 318 349 319
rect 582 319 583 320
rect 587 319 588 323
rect 630 323 631 324
rect 635 323 636 327
rect 630 322 636 323
rect 726 323 732 324
rect 726 322 727 323
rect 721 320 727 322
rect 582 318 588 319
rect 726 319 727 320
rect 731 319 732 323
rect 726 318 732 319
rect 110 317 116 318
rect 110 313 111 317
rect 115 313 116 317
rect 110 312 116 313
rect 134 317 140 318
rect 134 313 135 317
rect 139 313 140 317
rect 134 312 140 313
rect 214 317 220 318
rect 214 313 215 317
rect 219 313 220 317
rect 214 312 220 313
rect 302 317 308 318
rect 302 313 303 317
rect 307 313 308 317
rect 302 312 308 313
rect 398 317 404 318
rect 398 313 399 317
rect 403 313 404 317
rect 398 312 404 313
rect 494 317 500 318
rect 494 313 495 317
rect 499 313 500 317
rect 494 312 500 313
rect 590 317 596 318
rect 590 313 591 317
rect 595 313 596 317
rect 590 312 596 313
rect 686 317 692 318
rect 686 313 687 317
rect 691 313 692 317
rect 686 312 692 313
rect 774 317 780 318
rect 774 313 775 317
rect 779 313 780 317
rect 774 312 780 313
rect 110 299 116 300
rect 110 295 111 299
rect 115 295 116 299
rect 774 299 780 300
rect 110 294 116 295
rect 182 295 188 296
rect 182 294 183 295
rect 148 292 183 294
rect 148 290 150 292
rect 182 291 183 292
rect 187 291 188 295
rect 254 295 260 296
rect 254 294 255 295
rect 182 290 188 291
rect 228 292 255 294
rect 228 290 230 292
rect 254 291 255 292
rect 259 291 260 295
rect 343 295 349 296
rect 343 294 344 295
rect 254 290 260 291
rect 316 292 344 294
rect 316 290 318 292
rect 343 291 344 292
rect 348 291 349 295
rect 702 295 708 296
rect 702 294 703 295
rect 343 290 349 291
rect 700 291 703 294
rect 707 291 708 295
rect 774 295 775 299
rect 779 295 780 299
rect 774 294 780 295
rect 700 290 708 291
rect 145 289 151 290
rect 145 285 146 289
rect 150 285 151 289
rect 225 289 231 290
rect 145 284 151 285
rect 154 287 160 288
rect 154 283 155 287
rect 159 283 160 287
rect 225 285 226 289
rect 230 285 231 289
rect 313 289 319 290
rect 225 284 231 285
rect 234 287 240 288
rect 154 282 160 283
rect 234 283 235 287
rect 239 283 240 287
rect 313 285 314 289
rect 318 285 319 289
rect 697 289 703 290
rect 313 284 319 285
rect 322 287 328 288
rect 234 282 240 283
rect 322 283 323 287
rect 327 283 328 287
rect 322 282 328 283
rect 406 287 415 288
rect 406 283 407 287
rect 414 283 415 287
rect 406 282 415 283
rect 418 287 424 288
rect 418 283 419 287
rect 423 283 424 287
rect 418 282 424 283
rect 502 287 511 288
rect 502 283 503 287
rect 510 283 511 287
rect 502 282 511 283
rect 514 287 520 288
rect 514 283 515 287
rect 519 283 520 287
rect 514 282 520 283
rect 582 287 588 288
rect 582 283 583 287
rect 587 286 588 287
rect 601 287 607 288
rect 601 286 602 287
rect 587 284 602 286
rect 587 283 588 284
rect 582 282 588 283
rect 601 283 602 284
rect 606 283 607 287
rect 601 282 607 283
rect 610 287 616 288
rect 610 283 611 287
rect 615 283 616 287
rect 697 285 698 289
rect 702 285 703 289
rect 697 284 703 285
rect 706 287 712 288
rect 610 282 616 283
rect 706 283 707 287
rect 711 283 712 287
rect 706 282 712 283
rect 126 271 132 272
rect 126 267 127 271
rect 131 270 132 271
rect 145 271 151 272
rect 145 270 146 271
rect 131 268 146 270
rect 131 267 132 268
rect 126 266 132 267
rect 145 267 146 268
rect 150 267 151 271
rect 726 271 735 272
rect 145 266 151 267
rect 154 269 160 270
rect 154 265 155 269
rect 159 265 160 269
rect 210 269 216 270
rect 154 264 160 265
rect 166 267 172 268
rect 166 263 167 267
rect 171 266 172 267
rect 201 267 207 268
rect 201 266 202 267
rect 171 264 202 266
rect 171 263 172 264
rect 166 262 172 263
rect 201 263 202 264
rect 206 263 207 267
rect 210 265 211 269
rect 215 265 216 269
rect 298 269 304 270
rect 210 264 216 265
rect 222 267 228 268
rect 201 262 207 263
rect 222 263 223 267
rect 227 266 228 267
rect 289 267 295 268
rect 289 266 290 267
rect 227 264 290 266
rect 227 263 228 264
rect 222 262 228 263
rect 289 263 290 264
rect 294 263 295 267
rect 298 265 299 269
rect 303 265 304 269
rect 386 269 392 270
rect 298 264 304 265
rect 310 267 316 268
rect 289 262 295 263
rect 310 263 311 267
rect 315 266 316 267
rect 377 267 383 268
rect 377 266 378 267
rect 315 264 378 266
rect 315 263 316 264
rect 310 262 316 263
rect 377 263 378 264
rect 382 263 383 267
rect 386 265 387 269
rect 391 265 392 269
rect 474 269 480 270
rect 386 264 392 265
rect 447 267 453 268
rect 377 262 383 263
rect 447 263 448 267
rect 452 266 453 267
rect 465 267 471 268
rect 465 266 466 267
rect 452 264 466 266
rect 452 263 453 264
rect 447 262 453 263
rect 465 263 466 264
rect 470 263 471 267
rect 474 265 475 269
rect 479 265 480 269
rect 562 269 568 270
rect 474 264 480 265
rect 486 267 492 268
rect 465 262 471 263
rect 486 263 487 267
rect 491 266 492 267
rect 553 267 559 268
rect 553 266 554 267
rect 491 264 554 266
rect 491 263 492 264
rect 486 262 492 263
rect 553 263 554 264
rect 558 263 559 267
rect 562 265 563 269
rect 567 265 568 269
rect 650 269 656 270
rect 562 264 568 265
rect 641 267 647 268
rect 553 262 559 263
rect 641 263 642 267
rect 646 263 647 267
rect 650 265 651 269
rect 655 265 656 269
rect 726 267 727 271
rect 734 267 735 271
rect 726 266 735 267
rect 738 269 744 270
rect 650 264 656 265
rect 738 265 739 269
rect 743 265 744 269
rect 738 264 744 265
rect 641 262 647 263
rect 679 263 685 264
rect 679 262 680 263
rect 644 260 680 262
rect 679 259 680 260
rect 684 259 685 263
rect 679 258 685 259
rect 110 257 116 258
rect 110 253 111 257
rect 115 253 116 257
rect 110 252 116 253
rect 774 257 780 258
rect 774 253 775 257
rect 779 253 780 257
rect 774 252 780 253
rect 110 239 116 240
rect 110 235 111 239
rect 115 235 116 239
rect 110 234 116 235
rect 134 239 140 240
rect 134 235 135 239
rect 139 235 140 239
rect 134 234 140 235
rect 190 239 196 240
rect 190 235 191 239
rect 195 235 196 239
rect 190 234 196 235
rect 278 239 284 240
rect 278 235 279 239
rect 283 235 284 239
rect 278 234 284 235
rect 366 239 372 240
rect 366 235 367 239
rect 371 235 372 239
rect 366 234 372 235
rect 454 239 460 240
rect 454 235 455 239
rect 459 235 460 239
rect 454 234 460 235
rect 542 239 548 240
rect 542 235 543 239
rect 547 235 548 239
rect 542 234 548 235
rect 630 239 636 240
rect 630 235 631 239
rect 635 235 636 239
rect 630 234 636 235
rect 718 239 724 240
rect 718 235 719 239
rect 723 235 724 239
rect 718 234 724 235
rect 774 239 780 240
rect 774 235 775 239
rect 779 235 780 239
rect 774 234 780 235
rect 166 231 172 232
rect 166 227 167 231
rect 171 227 172 231
rect 166 226 172 227
rect 222 231 228 232
rect 222 227 223 231
rect 227 227 228 231
rect 222 226 228 227
rect 310 231 316 232
rect 310 227 311 231
rect 315 227 316 231
rect 310 226 316 227
rect 374 231 380 232
rect 374 227 375 231
rect 379 227 380 231
rect 374 226 380 227
rect 486 231 492 232
rect 486 227 487 231
rect 491 227 492 231
rect 486 226 492 227
rect 502 231 508 232
rect 502 227 503 231
rect 507 230 508 231
rect 654 231 660 232
rect 507 228 545 230
rect 507 227 508 228
rect 502 226 508 227
rect 654 227 655 231
rect 659 227 660 231
rect 654 226 660 227
rect 679 231 685 232
rect 679 227 680 231
rect 684 230 685 231
rect 684 228 721 230
rect 684 227 685 228
rect 679 226 685 227
rect 447 203 453 204
rect 174 199 180 200
rect 174 195 175 199
rect 179 198 180 199
rect 234 199 240 200
rect 179 196 185 198
rect 179 195 180 196
rect 174 194 180 195
rect 234 195 235 199
rect 239 198 240 199
rect 338 199 344 200
rect 239 196 273 198
rect 239 195 240 196
rect 234 194 240 195
rect 338 195 339 199
rect 343 198 344 199
rect 447 199 448 203
rect 452 202 453 203
rect 452 200 457 202
rect 452 199 453 200
rect 447 198 453 199
rect 494 199 500 200
rect 343 196 361 198
rect 343 195 344 196
rect 338 194 344 195
rect 494 195 495 199
rect 499 198 500 199
rect 702 199 708 200
rect 702 198 703 199
rect 499 196 553 198
rect 681 196 703 198
rect 499 195 500 196
rect 494 194 500 195
rect 702 195 703 196
rect 707 195 708 199
rect 702 194 708 195
rect 710 199 716 200
rect 710 195 711 199
rect 715 198 716 199
rect 715 196 721 198
rect 715 195 716 196
rect 710 194 716 195
rect 110 193 116 194
rect 110 189 111 193
rect 115 189 116 193
rect 110 188 116 189
rect 182 193 188 194
rect 182 189 183 193
rect 187 189 188 193
rect 182 188 188 189
rect 270 193 276 194
rect 270 189 271 193
rect 275 189 276 193
rect 270 188 276 189
rect 358 193 364 194
rect 358 189 359 193
rect 363 189 364 193
rect 358 188 364 189
rect 454 193 460 194
rect 454 189 455 193
rect 459 189 460 193
rect 454 188 460 189
rect 550 193 556 194
rect 550 189 551 193
rect 555 189 556 193
rect 550 188 556 189
rect 646 193 652 194
rect 646 189 647 193
rect 651 189 652 193
rect 646 188 652 189
rect 718 193 724 194
rect 718 189 719 193
rect 723 189 724 193
rect 718 188 724 189
rect 774 193 780 194
rect 774 189 775 193
rect 779 189 780 193
rect 774 188 780 189
rect 110 175 116 176
rect 110 171 111 175
rect 115 171 116 175
rect 774 175 780 176
rect 110 170 116 171
rect 234 171 240 172
rect 234 170 235 171
rect 196 168 235 170
rect 196 166 198 168
rect 234 167 235 168
rect 239 167 240 171
rect 338 171 344 172
rect 338 170 339 171
rect 234 166 240 167
rect 284 168 339 170
rect 284 166 286 168
rect 338 167 339 168
rect 343 167 344 171
rect 374 171 380 172
rect 374 170 375 171
rect 338 166 344 167
rect 372 167 375 170
rect 379 167 380 171
rect 494 171 500 172
rect 494 170 495 171
rect 372 166 380 167
rect 468 168 495 170
rect 468 166 470 168
rect 494 167 495 168
rect 499 167 500 171
rect 774 171 775 175
rect 779 171 780 175
rect 774 170 780 171
rect 494 166 500 167
rect 193 165 199 166
rect 193 161 194 165
rect 198 161 199 165
rect 281 165 287 166
rect 193 160 199 161
rect 202 163 208 164
rect 202 159 203 163
rect 207 159 208 163
rect 281 161 282 165
rect 286 161 287 165
rect 369 165 375 166
rect 281 160 287 161
rect 290 163 296 164
rect 202 158 208 159
rect 290 159 291 163
rect 295 159 296 163
rect 369 161 370 165
rect 374 161 375 165
rect 465 165 471 166
rect 369 160 375 161
rect 378 163 384 164
rect 290 158 296 159
rect 378 159 379 163
rect 383 159 384 163
rect 465 161 466 165
rect 470 161 471 165
rect 465 160 471 161
rect 474 163 480 164
rect 378 158 384 159
rect 474 159 475 163
rect 479 159 480 163
rect 474 158 480 159
rect 561 163 567 164
rect 561 159 562 163
rect 566 159 567 163
rect 561 158 567 159
rect 570 163 576 164
rect 570 159 571 163
rect 575 159 576 163
rect 570 158 576 159
rect 654 163 663 164
rect 654 159 655 163
rect 662 159 663 163
rect 654 158 663 159
rect 666 163 672 164
rect 666 159 667 163
rect 671 159 672 163
rect 666 158 672 159
rect 702 163 708 164
rect 702 159 703 163
rect 707 162 708 163
rect 729 163 735 164
rect 729 162 730 163
rect 707 160 730 162
rect 707 159 708 160
rect 702 158 708 159
rect 729 159 730 160
rect 734 159 735 163
rect 729 158 735 159
rect 738 163 744 164
rect 738 159 739 163
rect 743 159 744 163
rect 738 158 744 159
rect 564 154 566 158
rect 582 155 588 156
rect 582 154 583 155
rect 564 152 583 154
rect 582 151 583 152
rect 587 151 588 155
rect 582 150 588 151
rect 174 147 180 148
rect 174 143 175 147
rect 179 146 180 147
rect 201 147 207 148
rect 201 146 202 147
rect 179 144 202 146
rect 179 143 180 144
rect 174 142 180 143
rect 201 143 202 144
rect 206 143 207 147
rect 710 147 716 148
rect 201 142 207 143
rect 210 145 216 146
rect 210 141 211 145
rect 215 141 216 145
rect 258 145 264 146
rect 210 140 216 141
rect 222 143 228 144
rect 222 139 223 143
rect 227 142 228 143
rect 249 143 255 144
rect 249 142 250 143
rect 227 140 250 142
rect 227 139 228 140
rect 222 138 228 139
rect 249 139 250 140
rect 254 139 255 143
rect 258 141 259 145
rect 263 141 264 145
rect 306 145 312 146
rect 258 140 264 141
rect 270 143 276 144
rect 249 138 255 139
rect 270 139 271 143
rect 275 142 276 143
rect 297 143 303 144
rect 297 142 298 143
rect 275 140 298 142
rect 275 139 276 140
rect 270 138 276 139
rect 297 139 298 140
rect 302 139 303 143
rect 306 141 307 145
rect 311 141 312 145
rect 354 145 360 146
rect 306 140 312 141
rect 318 143 324 144
rect 297 138 303 139
rect 318 139 319 143
rect 323 142 324 143
rect 345 143 351 144
rect 345 142 346 143
rect 323 140 346 142
rect 323 139 324 140
rect 318 138 324 139
rect 345 139 346 140
rect 350 139 351 143
rect 354 141 355 145
rect 359 141 360 145
rect 402 145 408 146
rect 354 140 360 141
rect 366 143 372 144
rect 345 138 351 139
rect 366 139 367 143
rect 371 142 372 143
rect 393 143 399 144
rect 393 142 394 143
rect 371 140 394 142
rect 371 139 372 140
rect 366 138 372 139
rect 393 139 394 140
rect 398 139 399 143
rect 402 141 403 145
rect 407 141 408 145
rect 450 145 456 146
rect 402 140 408 141
rect 414 143 420 144
rect 393 138 399 139
rect 414 139 415 143
rect 419 142 420 143
rect 441 143 447 144
rect 441 142 442 143
rect 419 140 442 142
rect 419 139 420 140
rect 414 138 420 139
rect 441 139 442 140
rect 446 139 447 143
rect 450 141 451 145
rect 455 141 456 145
rect 498 145 504 146
rect 450 140 456 141
rect 462 143 468 144
rect 441 138 447 139
rect 462 139 463 143
rect 467 142 468 143
rect 489 143 495 144
rect 489 142 490 143
rect 467 140 490 142
rect 467 139 468 140
rect 462 138 468 139
rect 489 139 490 140
rect 494 139 495 143
rect 498 141 499 145
rect 503 141 504 145
rect 546 145 552 146
rect 498 140 504 141
rect 510 143 516 144
rect 489 138 495 139
rect 510 139 511 143
rect 515 142 516 143
rect 537 143 543 144
rect 537 142 538 143
rect 515 140 538 142
rect 515 139 516 140
rect 510 138 516 139
rect 537 139 538 140
rect 542 139 543 143
rect 546 141 547 145
rect 551 141 552 145
rect 594 145 600 146
rect 546 140 552 141
rect 558 143 564 144
rect 537 138 543 139
rect 558 139 559 143
rect 563 142 564 143
rect 585 143 591 144
rect 585 142 586 143
rect 563 140 586 142
rect 563 139 564 140
rect 558 138 564 139
rect 585 139 586 140
rect 590 139 591 143
rect 594 141 595 145
rect 599 141 600 145
rect 642 145 648 146
rect 594 140 600 141
rect 633 143 639 144
rect 585 138 591 139
rect 633 139 634 143
rect 638 139 639 143
rect 642 141 643 145
rect 647 141 648 145
rect 690 145 696 146
rect 642 140 648 141
rect 681 143 687 144
rect 633 138 639 139
rect 662 139 668 140
rect 662 138 663 139
rect 636 136 663 138
rect 662 135 663 136
rect 667 135 668 139
rect 681 139 682 143
rect 686 139 687 143
rect 690 141 691 145
rect 695 141 696 145
rect 710 143 711 147
rect 715 146 716 147
rect 729 147 735 148
rect 729 146 730 147
rect 715 144 730 146
rect 715 143 716 144
rect 710 142 716 143
rect 729 143 730 144
rect 734 143 735 147
rect 729 142 735 143
rect 738 145 744 146
rect 690 140 696 141
rect 738 141 739 145
rect 743 141 744 145
rect 738 140 744 141
rect 681 138 687 139
rect 710 139 716 140
rect 710 138 711 139
rect 684 136 711 138
rect 662 134 668 135
rect 710 135 711 136
rect 715 135 716 139
rect 710 134 716 135
rect 110 133 116 134
rect 110 129 111 133
rect 115 129 116 133
rect 110 128 116 129
rect 774 133 780 134
rect 774 129 775 133
rect 779 129 780 133
rect 774 128 780 129
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 110 110 116 111
rect 190 115 196 116
rect 190 111 191 115
rect 195 111 196 115
rect 190 110 196 111
rect 238 115 244 116
rect 238 111 239 115
rect 243 111 244 115
rect 238 110 244 111
rect 286 115 292 116
rect 286 111 287 115
rect 291 111 292 115
rect 286 110 292 111
rect 334 115 340 116
rect 334 111 335 115
rect 339 111 340 115
rect 334 110 340 111
rect 382 115 388 116
rect 382 111 383 115
rect 387 111 388 115
rect 382 110 388 111
rect 430 115 436 116
rect 430 111 431 115
rect 435 111 436 115
rect 430 110 436 111
rect 478 115 484 116
rect 478 111 479 115
rect 483 111 484 115
rect 478 110 484 111
rect 526 115 532 116
rect 526 111 527 115
rect 531 111 532 115
rect 526 110 532 111
rect 574 115 580 116
rect 574 111 575 115
rect 579 111 580 115
rect 574 110 580 111
rect 622 115 628 116
rect 622 111 623 115
rect 627 111 628 115
rect 622 110 628 111
rect 670 115 676 116
rect 670 111 671 115
rect 675 111 676 115
rect 670 110 676 111
rect 718 115 724 116
rect 718 111 719 115
rect 723 111 724 115
rect 718 110 724 111
rect 774 115 780 116
rect 774 111 775 115
rect 779 111 780 115
rect 774 110 780 111
rect 222 107 228 108
rect 222 103 223 107
rect 227 103 228 107
rect 222 102 228 103
rect 270 107 276 108
rect 270 103 271 107
rect 275 103 276 107
rect 270 102 276 103
rect 318 107 324 108
rect 318 103 319 107
rect 323 103 324 107
rect 318 102 324 103
rect 366 107 372 108
rect 366 103 367 107
rect 371 103 372 107
rect 366 102 372 103
rect 414 107 420 108
rect 414 103 415 107
rect 419 103 420 107
rect 414 102 420 103
rect 462 107 468 108
rect 462 103 463 107
rect 467 103 468 107
rect 462 102 468 103
rect 510 107 516 108
rect 510 103 511 107
rect 515 103 516 107
rect 510 102 516 103
rect 558 107 564 108
rect 558 103 559 107
rect 563 103 564 107
rect 558 102 564 103
rect 582 107 588 108
rect 582 103 583 107
rect 587 103 588 107
rect 582 102 588 103
rect 662 107 668 108
rect 662 103 663 107
rect 667 106 668 107
rect 710 107 716 108
rect 667 104 673 106
rect 667 103 668 104
rect 662 102 668 103
rect 710 103 711 107
rect 715 106 716 107
rect 715 104 721 106
rect 715 103 716 104
rect 710 102 716 103
<< m3c >>
rect 155 853 159 857
rect 167 851 171 855
rect 203 853 207 857
rect 215 851 219 855
rect 251 853 255 857
rect 263 851 267 855
rect 299 853 303 857
rect 311 851 315 855
rect 347 853 351 857
rect 111 841 115 845
rect 775 841 779 845
rect 111 823 115 827
rect 135 823 139 827
rect 183 823 187 827
rect 231 823 235 827
rect 279 823 283 827
rect 327 823 331 827
rect 775 823 779 827
rect 167 815 171 819
rect 215 815 219 819
rect 263 815 267 819
rect 311 815 315 819
rect 319 815 323 819
rect 343 791 347 795
rect 391 791 395 795
rect 439 791 443 795
rect 487 791 491 795
rect 495 787 499 791
rect 111 781 115 785
rect 311 781 315 785
rect 359 781 363 785
rect 407 781 411 785
rect 455 781 459 785
rect 503 781 507 785
rect 775 781 779 785
rect 111 763 115 767
rect 487 759 491 763
rect 775 763 779 767
rect 319 751 322 755
rect 322 751 323 755
rect 331 751 335 755
rect 343 751 347 755
rect 379 751 383 755
rect 391 751 395 755
rect 427 751 431 755
rect 439 751 443 755
rect 475 751 479 755
rect 523 751 527 755
rect 259 741 263 745
rect 271 739 275 743
rect 307 741 311 745
rect 319 739 323 743
rect 355 741 359 745
rect 403 741 407 745
rect 111 729 115 733
rect 375 731 379 735
rect 423 735 427 739
rect 451 741 455 745
rect 487 743 490 747
rect 490 743 491 747
rect 499 741 503 745
rect 471 735 475 739
rect 535 739 538 743
rect 538 739 539 743
rect 547 741 551 745
rect 559 739 563 743
rect 595 741 599 745
rect 607 739 611 743
rect 643 741 647 745
rect 655 739 659 743
rect 691 741 695 745
rect 703 739 707 743
rect 739 741 743 745
rect 775 729 779 733
rect 111 711 115 715
rect 239 711 243 715
rect 287 711 291 715
rect 335 711 339 715
rect 383 711 387 715
rect 431 711 435 715
rect 479 711 483 715
rect 527 711 531 715
rect 575 711 579 715
rect 623 711 627 715
rect 671 711 675 715
rect 719 711 723 715
rect 775 711 779 715
rect 271 703 275 707
rect 319 703 323 707
rect 367 703 371 707
rect 375 703 379 707
rect 423 703 427 707
rect 471 703 475 707
rect 559 703 563 707
rect 607 703 611 707
rect 655 703 659 707
rect 703 703 707 707
rect 727 703 731 707
rect 127 667 131 671
rect 175 667 179 671
rect 415 671 419 675
rect 423 667 427 671
rect 535 671 539 675
rect 711 667 715 671
rect 111 661 115 665
rect 135 661 139 665
rect 191 661 195 665
rect 279 661 283 665
rect 383 661 387 665
rect 495 661 499 665
rect 615 661 619 665
rect 719 661 723 665
rect 775 661 779 665
rect 111 643 115 647
rect 175 639 179 643
rect 423 639 427 643
rect 775 643 779 647
rect 155 631 159 635
rect 211 631 215 635
rect 299 631 303 635
rect 367 631 371 635
rect 403 631 407 635
rect 415 631 419 635
rect 515 631 519 635
rect 127 623 131 627
rect 615 627 619 631
rect 635 631 639 635
rect 727 631 730 635
rect 730 631 731 635
rect 739 631 743 635
rect 155 621 159 625
rect 167 619 171 623
rect 203 621 207 625
rect 275 621 279 625
rect 287 619 291 623
rect 379 621 383 625
rect 391 619 395 623
rect 499 621 503 625
rect 551 619 555 623
rect 627 621 631 625
rect 711 623 715 627
rect 739 621 743 625
rect 111 609 115 613
rect 775 609 779 613
rect 111 591 115 595
rect 135 591 139 595
rect 183 591 187 595
rect 255 591 259 595
rect 359 591 363 595
rect 479 591 483 595
rect 607 591 611 595
rect 719 591 723 595
rect 775 591 779 595
rect 167 583 171 587
rect 287 583 291 587
rect 391 583 395 587
rect 551 583 555 587
rect 559 583 563 587
rect 727 583 731 587
rect 459 563 463 567
rect 175 555 179 559
rect 231 555 235 559
rect 295 555 299 559
rect 407 555 411 559
rect 511 555 515 559
rect 615 559 619 563
rect 711 555 715 559
rect 111 549 115 553
rect 135 549 139 553
rect 183 549 187 553
rect 239 549 243 553
rect 319 549 323 553
rect 415 549 419 553
rect 519 549 523 553
rect 631 549 635 553
rect 719 549 723 553
rect 775 549 779 553
rect 111 531 115 535
rect 775 531 779 535
rect 143 519 146 523
rect 146 519 147 523
rect 155 519 159 523
rect 175 519 179 523
rect 203 519 207 523
rect 231 519 235 523
rect 259 519 263 523
rect 295 519 299 523
rect 339 519 343 523
rect 407 519 411 523
rect 435 519 439 523
rect 511 519 515 523
rect 539 519 543 523
rect 639 519 642 523
rect 642 519 643 523
rect 651 519 655 523
rect 727 519 730 523
rect 730 519 731 523
rect 739 519 743 523
rect 459 507 463 511
rect 283 501 287 505
rect 295 499 299 503
rect 331 501 335 505
rect 359 499 363 503
rect 387 501 391 505
rect 399 499 403 503
rect 451 501 455 505
rect 463 499 467 503
rect 515 501 519 505
rect 527 499 531 503
rect 587 501 591 505
rect 667 501 671 505
rect 711 503 715 507
rect 739 501 743 505
rect 687 495 691 499
rect 111 489 115 493
rect 775 489 779 493
rect 111 471 115 475
rect 263 471 267 475
rect 311 471 315 475
rect 367 471 371 475
rect 431 471 435 475
rect 495 471 499 475
rect 567 471 571 475
rect 647 471 651 475
rect 719 471 723 475
rect 775 471 779 475
rect 295 463 299 467
rect 359 463 363 467
rect 399 463 403 467
rect 463 463 467 467
rect 527 463 531 467
rect 535 463 539 467
rect 639 463 643 467
rect 727 463 731 467
rect 455 431 459 435
rect 495 435 499 439
rect 551 431 555 435
rect 591 435 595 439
rect 599 431 603 435
rect 687 435 691 439
rect 703 431 707 435
rect 111 425 115 429
rect 415 425 419 429
rect 463 425 467 429
rect 511 425 515 429
rect 559 425 563 429
rect 607 425 611 429
rect 655 425 659 429
rect 711 425 715 429
rect 775 425 779 429
rect 111 407 115 411
rect 535 407 539 411
rect 435 395 439 399
rect 455 399 459 403
rect 727 403 731 407
rect 775 407 779 411
rect 483 395 487 399
rect 495 395 499 399
rect 531 395 535 399
rect 551 395 555 399
rect 579 395 583 399
rect 591 395 595 399
rect 627 395 631 399
rect 655 395 659 399
rect 675 395 679 399
rect 731 395 735 399
rect 307 385 311 389
rect 319 383 323 387
rect 355 385 359 389
rect 367 383 371 387
rect 403 385 407 389
rect 451 385 455 389
rect 111 373 115 377
rect 423 375 427 379
rect 471 379 475 383
rect 507 385 511 389
rect 527 379 531 383
rect 571 385 575 389
rect 599 379 603 383
rect 643 385 647 389
rect 703 387 706 391
rect 706 387 707 391
rect 715 385 719 389
rect 631 379 635 383
rect 775 373 779 377
rect 111 355 115 359
rect 287 355 291 359
rect 335 355 339 359
rect 383 355 387 359
rect 431 355 435 359
rect 487 355 491 359
rect 551 355 555 359
rect 623 355 627 359
rect 695 355 699 359
rect 775 355 779 359
rect 319 347 323 351
rect 367 347 371 351
rect 407 347 411 351
rect 423 347 427 351
rect 471 347 475 351
rect 527 347 531 351
rect 655 347 659 351
rect 703 347 707 351
rect 127 319 131 323
rect 183 319 187 323
rect 255 319 259 323
rect 583 319 587 323
rect 631 323 635 327
rect 727 319 731 323
rect 111 313 115 317
rect 135 313 139 317
rect 215 313 219 317
rect 303 313 307 317
rect 399 313 403 317
rect 495 313 499 317
rect 591 313 595 317
rect 687 313 691 317
rect 775 313 779 317
rect 111 295 115 299
rect 183 291 187 295
rect 255 291 259 295
rect 703 291 707 295
rect 775 295 779 299
rect 155 283 159 287
rect 235 283 239 287
rect 323 283 327 287
rect 407 283 410 287
rect 410 283 411 287
rect 419 283 423 287
rect 503 283 506 287
rect 506 283 507 287
rect 515 283 519 287
rect 583 283 587 287
rect 611 283 615 287
rect 707 283 711 287
rect 127 267 131 271
rect 155 265 159 269
rect 167 263 171 267
rect 211 265 215 269
rect 223 263 227 267
rect 299 265 303 269
rect 311 263 315 267
rect 387 265 391 269
rect 475 265 479 269
rect 487 263 491 267
rect 563 265 567 269
rect 651 265 655 269
rect 727 267 730 271
rect 730 267 731 271
rect 739 265 743 269
rect 111 253 115 257
rect 775 253 779 257
rect 111 235 115 239
rect 135 235 139 239
rect 191 235 195 239
rect 279 235 283 239
rect 367 235 371 239
rect 455 235 459 239
rect 543 235 547 239
rect 631 235 635 239
rect 719 235 723 239
rect 775 235 779 239
rect 167 227 171 231
rect 223 227 227 231
rect 311 227 315 231
rect 375 227 379 231
rect 487 227 491 231
rect 503 227 507 231
rect 655 227 659 231
rect 175 195 179 199
rect 235 195 239 199
rect 339 195 343 199
rect 495 195 499 199
rect 703 195 707 199
rect 711 195 715 199
rect 111 189 115 193
rect 183 189 187 193
rect 271 189 275 193
rect 359 189 363 193
rect 455 189 459 193
rect 551 189 555 193
rect 647 189 651 193
rect 719 189 723 193
rect 775 189 779 193
rect 111 171 115 175
rect 235 167 239 171
rect 339 167 343 171
rect 375 167 379 171
rect 495 167 499 171
rect 775 171 779 175
rect 203 159 207 163
rect 291 159 295 163
rect 379 159 383 163
rect 475 159 479 163
rect 571 159 575 163
rect 655 159 658 163
rect 658 159 659 163
rect 667 159 671 163
rect 703 159 707 163
rect 739 159 743 163
rect 583 151 587 155
rect 175 143 179 147
rect 211 141 215 145
rect 223 139 227 143
rect 259 141 263 145
rect 271 139 275 143
rect 307 141 311 145
rect 319 139 323 143
rect 355 141 359 145
rect 367 139 371 143
rect 403 141 407 145
rect 415 139 419 143
rect 451 141 455 145
rect 463 139 467 143
rect 499 141 503 145
rect 511 139 515 143
rect 547 141 551 145
rect 559 139 563 143
rect 595 141 599 145
rect 643 141 647 145
rect 663 135 667 139
rect 691 141 695 145
rect 711 143 715 147
rect 739 141 743 145
rect 711 135 715 139
rect 111 129 115 133
rect 775 129 779 133
rect 111 111 115 115
rect 191 111 195 115
rect 239 111 243 115
rect 287 111 291 115
rect 335 111 339 115
rect 383 111 387 115
rect 431 111 435 115
rect 479 111 483 115
rect 527 111 531 115
rect 575 111 579 115
rect 623 111 627 115
rect 671 111 675 115
rect 719 111 723 115
rect 775 111 779 115
rect 223 103 227 107
rect 271 103 275 107
rect 319 103 323 107
rect 367 103 371 107
rect 415 103 419 107
rect 463 103 467 107
rect 511 103 515 107
rect 559 103 563 107
rect 583 103 587 107
rect 663 103 667 107
rect 711 103 715 107
<< m3 >>
rect 111 862 115 863
rect 155 862 159 863
rect 203 862 207 863
rect 251 862 255 863
rect 299 862 303 863
rect 347 862 351 863
rect 775 862 779 863
rect 111 857 115 858
rect 154 857 160 858
rect 112 846 114 857
rect 154 853 155 857
rect 159 853 160 857
rect 202 857 208 858
rect 154 852 160 853
rect 166 855 172 856
rect 166 851 167 855
rect 171 851 172 855
rect 202 853 203 857
rect 207 853 208 857
rect 250 857 256 858
rect 202 852 208 853
rect 214 855 220 856
rect 166 850 172 851
rect 214 851 215 855
rect 219 851 220 855
rect 250 853 251 857
rect 255 853 256 857
rect 298 857 304 858
rect 250 852 256 853
rect 262 855 268 856
rect 214 850 220 851
rect 262 851 263 855
rect 267 851 268 855
rect 298 853 299 857
rect 303 853 304 857
rect 346 857 352 858
rect 775 857 779 858
rect 298 852 304 853
rect 310 855 316 856
rect 262 850 268 851
rect 310 851 311 855
rect 315 851 316 855
rect 346 853 347 857
rect 351 853 352 857
rect 346 852 352 853
rect 310 850 316 851
rect 110 845 116 846
rect 110 841 111 845
rect 115 841 116 845
rect 110 840 116 841
rect 110 827 116 828
rect 110 823 111 827
rect 115 823 116 827
rect 110 822 116 823
rect 134 827 140 828
rect 134 823 135 827
rect 139 823 140 827
rect 134 822 140 823
rect 112 807 114 822
rect 136 807 138 822
rect 168 820 170 850
rect 182 827 188 828
rect 182 823 183 827
rect 187 823 188 827
rect 182 822 188 823
rect 166 819 172 820
rect 166 815 167 819
rect 171 815 172 819
rect 166 814 172 815
rect 184 807 186 822
rect 216 820 218 850
rect 230 827 236 828
rect 230 823 231 827
rect 235 823 236 827
rect 230 822 236 823
rect 214 819 220 820
rect 214 815 215 819
rect 219 815 220 819
rect 214 814 220 815
rect 232 807 234 822
rect 264 820 266 850
rect 278 827 284 828
rect 278 823 279 827
rect 283 823 284 827
rect 278 822 284 823
rect 262 819 268 820
rect 262 815 263 819
rect 267 815 268 819
rect 262 814 268 815
rect 280 807 282 822
rect 312 820 314 850
rect 776 846 778 857
rect 774 845 780 846
rect 774 841 775 845
rect 779 841 780 845
rect 774 840 780 841
rect 326 827 332 828
rect 326 823 327 827
rect 331 823 332 827
rect 326 822 332 823
rect 774 827 780 828
rect 774 823 775 827
rect 779 823 780 827
rect 774 822 780 823
rect 310 819 316 820
rect 310 815 311 819
rect 315 815 316 819
rect 310 814 316 815
rect 318 819 324 820
rect 318 815 319 819
rect 323 815 324 819
rect 318 814 324 815
rect 111 806 115 807
rect 111 801 115 802
rect 135 806 139 807
rect 135 801 139 802
rect 183 806 187 807
rect 183 801 187 802
rect 231 806 235 807
rect 231 801 235 802
rect 279 806 283 807
rect 279 801 283 802
rect 311 806 315 807
rect 311 801 315 802
rect 112 786 114 801
rect 312 786 314 801
rect 110 785 116 786
rect 110 781 111 785
rect 115 781 116 785
rect 110 780 116 781
rect 310 785 316 786
rect 310 781 311 785
rect 315 781 316 785
rect 310 780 316 781
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 110 762 116 763
rect 112 751 114 762
rect 320 756 322 814
rect 328 807 330 822
rect 776 807 778 822
rect 327 806 331 807
rect 327 801 331 802
rect 359 806 363 807
rect 359 801 363 802
rect 407 806 411 807
rect 407 801 411 802
rect 455 806 459 807
rect 455 801 459 802
rect 503 806 507 807
rect 503 801 507 802
rect 775 806 779 807
rect 775 801 779 802
rect 342 795 348 796
rect 342 791 343 795
rect 347 791 348 795
rect 342 790 348 791
rect 344 756 346 790
rect 360 786 362 801
rect 390 795 396 796
rect 390 791 391 795
rect 395 791 396 795
rect 390 790 396 791
rect 358 785 364 786
rect 358 781 359 785
rect 363 781 364 785
rect 358 780 364 781
rect 392 756 394 790
rect 408 786 410 801
rect 438 795 444 796
rect 438 791 439 795
rect 443 791 444 795
rect 438 790 444 791
rect 406 785 412 786
rect 406 781 407 785
rect 411 781 412 785
rect 406 780 412 781
rect 440 756 442 790
rect 456 786 458 801
rect 486 795 492 796
rect 486 791 487 795
rect 491 791 492 795
rect 486 790 492 791
rect 494 791 500 792
rect 454 785 460 786
rect 454 781 455 785
rect 459 781 460 785
rect 454 780 460 781
rect 488 764 490 790
rect 494 787 495 791
rect 499 787 500 791
rect 494 786 500 787
rect 504 786 506 801
rect 776 786 778 801
rect 486 763 492 764
rect 486 759 487 763
rect 491 759 492 763
rect 486 758 492 759
rect 318 755 324 756
rect 318 751 319 755
rect 323 751 324 755
rect 111 750 115 751
rect 259 750 263 751
rect 307 750 311 751
rect 318 750 324 751
rect 330 755 336 756
rect 330 751 331 755
rect 335 751 336 755
rect 330 750 336 751
rect 342 755 348 756
rect 342 751 343 755
rect 347 751 348 755
rect 378 755 384 756
rect 378 751 379 755
rect 383 751 384 755
rect 342 750 348 751
rect 355 750 359 751
rect 378 750 384 751
rect 390 755 396 756
rect 390 751 391 755
rect 395 751 396 755
rect 426 755 432 756
rect 426 751 427 755
rect 431 751 432 755
rect 390 750 396 751
rect 403 750 407 751
rect 426 750 432 751
rect 438 755 444 756
rect 438 751 439 755
rect 443 751 444 755
rect 474 755 480 756
rect 496 755 498 786
rect 502 785 508 786
rect 502 781 503 785
rect 507 781 508 785
rect 502 780 508 781
rect 774 785 780 786
rect 774 781 775 785
rect 779 781 780 785
rect 774 780 780 781
rect 774 767 780 768
rect 774 763 775 767
rect 779 763 780 767
rect 774 762 780 763
rect 474 751 475 755
rect 479 751 480 755
rect 438 750 444 751
rect 451 750 455 751
rect 474 750 480 751
rect 488 753 498 755
rect 522 755 528 756
rect 488 748 490 753
rect 522 751 523 755
rect 527 751 528 755
rect 776 751 778 762
rect 499 750 503 751
rect 522 750 528 751
rect 547 750 551 751
rect 111 745 115 746
rect 258 745 264 746
rect 112 734 114 745
rect 258 741 259 745
rect 263 741 264 745
rect 306 745 312 746
rect 331 745 335 746
rect 354 745 360 746
rect 379 745 383 746
rect 402 745 408 746
rect 427 745 431 746
rect 450 745 456 746
rect 475 745 479 746
rect 486 747 492 748
rect 258 740 264 741
rect 270 743 276 744
rect 270 739 271 743
rect 275 739 276 743
rect 306 741 307 745
rect 311 741 312 745
rect 306 740 312 741
rect 318 743 324 744
rect 270 738 276 739
rect 318 739 319 743
rect 323 739 324 743
rect 354 741 355 745
rect 359 741 360 745
rect 354 740 360 741
rect 402 741 403 745
rect 407 741 408 745
rect 402 740 408 741
rect 450 741 451 745
rect 455 741 456 745
rect 486 743 487 747
rect 491 743 492 747
rect 595 750 599 751
rect 643 750 647 751
rect 691 750 695 751
rect 739 750 743 751
rect 775 750 779 751
rect 486 742 492 743
rect 498 745 504 746
rect 523 745 527 746
rect 546 745 552 746
rect 450 740 456 741
rect 498 741 499 745
rect 503 741 504 745
rect 498 740 504 741
rect 534 743 540 744
rect 318 738 324 739
rect 422 739 428 740
rect 110 733 116 734
rect 110 729 111 733
rect 115 729 116 733
rect 110 728 116 729
rect 110 715 116 716
rect 110 711 111 715
rect 115 711 116 715
rect 110 710 116 711
rect 238 715 244 716
rect 238 711 239 715
rect 243 711 244 715
rect 238 710 244 711
rect 112 687 114 710
rect 240 687 242 710
rect 272 708 274 738
rect 286 715 292 716
rect 286 711 287 715
rect 291 711 292 715
rect 286 710 292 711
rect 270 707 276 708
rect 270 703 271 707
rect 275 703 276 707
rect 270 702 276 703
rect 288 687 290 710
rect 320 708 322 738
rect 374 735 380 736
rect 374 731 375 735
rect 379 731 380 735
rect 422 735 423 739
rect 427 735 428 739
rect 422 734 428 735
rect 470 739 476 740
rect 470 735 471 739
rect 475 735 476 739
rect 534 739 535 743
rect 539 739 540 743
rect 546 741 547 745
rect 551 741 552 745
rect 594 745 600 746
rect 546 740 552 741
rect 558 743 564 744
rect 534 738 540 739
rect 558 739 559 743
rect 563 739 564 743
rect 594 741 595 745
rect 599 741 600 745
rect 642 745 648 746
rect 594 740 600 741
rect 606 743 612 744
rect 558 738 564 739
rect 606 739 607 743
rect 611 739 612 743
rect 642 741 643 745
rect 647 741 648 745
rect 690 745 696 746
rect 642 740 648 741
rect 654 743 660 744
rect 606 738 612 739
rect 654 739 655 743
rect 659 739 660 743
rect 690 741 691 745
rect 695 741 696 745
rect 738 745 744 746
rect 775 745 779 746
rect 690 740 696 741
rect 702 743 708 744
rect 654 738 660 739
rect 702 739 703 743
rect 707 739 708 743
rect 738 741 739 745
rect 743 741 744 745
rect 738 740 744 741
rect 702 738 708 739
rect 470 734 476 735
rect 374 730 380 731
rect 334 715 340 716
rect 334 711 335 715
rect 339 711 340 715
rect 334 710 340 711
rect 318 707 324 708
rect 318 703 319 707
rect 323 703 324 707
rect 318 702 324 703
rect 336 687 338 710
rect 376 708 378 730
rect 382 715 388 716
rect 382 711 383 715
rect 387 711 388 715
rect 382 710 388 711
rect 366 707 372 708
rect 366 703 367 707
rect 371 703 372 707
rect 366 702 372 703
rect 374 707 380 708
rect 374 703 375 707
rect 379 703 380 707
rect 374 702 380 703
rect 111 686 115 687
rect 111 681 115 682
rect 135 686 139 687
rect 135 681 139 682
rect 191 686 195 687
rect 191 681 195 682
rect 239 686 243 687
rect 239 681 243 682
rect 279 686 283 687
rect 279 681 283 682
rect 287 686 291 687
rect 287 681 291 682
rect 335 686 339 687
rect 335 681 339 682
rect 112 666 114 681
rect 126 671 132 672
rect 126 667 127 671
rect 131 667 132 671
rect 126 666 132 667
rect 136 666 138 681
rect 174 671 180 672
rect 174 667 175 671
rect 179 667 180 671
rect 174 666 180 667
rect 192 666 194 681
rect 280 666 282 681
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 110 660 116 661
rect 110 647 116 648
rect 110 643 111 647
rect 115 643 116 647
rect 110 642 116 643
rect 112 631 114 642
rect 111 630 115 631
rect 128 628 130 666
rect 134 665 140 666
rect 134 661 135 665
rect 139 661 140 665
rect 134 660 140 661
rect 176 644 178 666
rect 190 665 196 666
rect 190 661 191 665
rect 195 661 196 665
rect 190 660 196 661
rect 278 665 284 666
rect 278 661 279 665
rect 283 661 284 665
rect 278 660 284 661
rect 174 643 180 644
rect 174 639 175 643
rect 179 639 180 643
rect 174 638 180 639
rect 368 636 370 702
rect 384 687 386 710
rect 424 708 426 734
rect 430 715 436 716
rect 430 711 431 715
rect 435 711 436 715
rect 430 710 436 711
rect 422 707 428 708
rect 422 703 423 707
rect 427 703 428 707
rect 422 702 428 703
rect 432 687 434 710
rect 472 708 474 734
rect 478 715 484 716
rect 478 711 479 715
rect 483 711 484 715
rect 478 710 484 711
rect 526 715 532 716
rect 526 711 527 715
rect 531 711 532 715
rect 526 710 532 711
rect 470 707 476 708
rect 470 703 471 707
rect 475 703 476 707
rect 470 702 476 703
rect 480 687 482 710
rect 528 687 530 710
rect 383 686 387 687
rect 383 681 387 682
rect 431 686 435 687
rect 431 681 435 682
rect 479 686 483 687
rect 479 681 483 682
rect 495 686 499 687
rect 495 681 499 682
rect 527 686 531 687
rect 527 681 531 682
rect 384 666 386 681
rect 414 675 420 676
rect 414 671 415 675
rect 419 671 420 675
rect 414 670 420 671
rect 422 671 428 672
rect 382 665 388 666
rect 382 661 383 665
rect 387 661 388 665
rect 382 660 388 661
rect 416 636 418 670
rect 422 667 423 671
rect 427 667 428 671
rect 422 666 428 667
rect 496 666 498 681
rect 536 676 538 738
rect 560 708 562 738
rect 574 715 580 716
rect 574 711 575 715
rect 579 711 580 715
rect 574 710 580 711
rect 558 707 564 708
rect 558 703 559 707
rect 563 703 564 707
rect 558 702 564 703
rect 576 687 578 710
rect 608 708 610 738
rect 622 715 628 716
rect 622 711 623 715
rect 627 711 628 715
rect 622 710 628 711
rect 606 707 612 708
rect 606 703 607 707
rect 611 703 612 707
rect 606 702 612 703
rect 624 687 626 710
rect 656 708 658 738
rect 670 715 676 716
rect 670 711 671 715
rect 675 711 676 715
rect 670 710 676 711
rect 654 707 660 708
rect 654 703 655 707
rect 659 703 660 707
rect 654 702 660 703
rect 672 687 674 710
rect 704 708 706 738
rect 776 734 778 745
rect 774 733 780 734
rect 774 729 775 733
rect 779 729 780 733
rect 774 728 780 729
rect 718 715 724 716
rect 718 711 719 715
rect 723 711 724 715
rect 718 710 724 711
rect 774 715 780 716
rect 774 711 775 715
rect 779 711 780 715
rect 774 710 780 711
rect 702 707 708 708
rect 702 703 703 707
rect 707 703 708 707
rect 702 702 708 703
rect 720 687 722 710
rect 726 707 732 708
rect 726 703 727 707
rect 731 703 732 707
rect 726 702 732 703
rect 575 686 579 687
rect 575 681 579 682
rect 615 686 619 687
rect 615 681 619 682
rect 623 686 627 687
rect 623 681 627 682
rect 671 686 675 687
rect 671 681 675 682
rect 719 686 723 687
rect 719 681 723 682
rect 534 675 540 676
rect 534 671 535 675
rect 539 671 540 675
rect 534 670 540 671
rect 616 666 618 681
rect 710 671 716 672
rect 710 667 711 671
rect 715 667 716 671
rect 710 666 716 667
rect 720 666 722 681
rect 424 644 426 666
rect 494 665 500 666
rect 494 661 495 665
rect 499 661 500 665
rect 494 660 500 661
rect 614 665 620 666
rect 614 661 615 665
rect 619 661 620 665
rect 614 660 620 661
rect 422 643 428 644
rect 422 639 423 643
rect 427 639 428 643
rect 422 638 428 639
rect 154 635 160 636
rect 154 631 155 635
rect 159 631 160 635
rect 210 635 216 636
rect 210 631 211 635
rect 215 631 216 635
rect 298 635 304 636
rect 298 631 299 635
rect 303 631 304 635
rect 154 630 160 631
rect 203 630 207 631
rect 210 630 216 631
rect 275 630 279 631
rect 298 630 304 631
rect 366 635 372 636
rect 366 631 367 635
rect 371 631 372 635
rect 402 635 408 636
rect 402 631 403 635
rect 407 631 408 635
rect 366 630 372 631
rect 379 630 383 631
rect 402 630 408 631
rect 414 635 420 636
rect 414 631 415 635
rect 419 631 420 635
rect 514 635 520 636
rect 514 631 515 635
rect 519 631 520 635
rect 634 635 640 636
rect 414 630 420 631
rect 499 630 503 631
rect 514 630 520 631
rect 614 631 620 632
rect 634 631 635 635
rect 639 631 640 635
rect 111 625 115 626
rect 126 627 132 628
rect 112 614 114 625
rect 126 623 127 627
rect 131 623 132 627
rect 614 627 615 631
rect 619 627 620 631
rect 614 626 620 627
rect 627 630 631 631
rect 634 630 640 631
rect 712 628 714 666
rect 718 665 724 666
rect 718 661 719 665
rect 723 661 724 665
rect 718 660 724 661
rect 728 636 730 702
rect 776 687 778 710
rect 775 686 779 687
rect 775 681 779 682
rect 776 666 778 681
rect 774 665 780 666
rect 774 661 775 665
rect 779 661 780 665
rect 774 660 780 661
rect 774 647 780 648
rect 774 643 775 647
rect 779 643 780 647
rect 774 642 780 643
rect 726 635 732 636
rect 726 631 727 635
rect 731 631 732 635
rect 726 630 732 631
rect 738 635 744 636
rect 738 631 739 635
rect 743 631 744 635
rect 776 631 778 642
rect 738 630 744 631
rect 775 630 779 631
rect 126 622 132 623
rect 154 625 160 626
rect 154 621 155 625
rect 159 621 160 625
rect 202 625 208 626
rect 211 625 215 626
rect 274 625 280 626
rect 299 625 303 626
rect 378 625 384 626
rect 403 625 407 626
rect 498 625 504 626
rect 515 625 519 626
rect 154 620 160 621
rect 166 623 172 624
rect 166 619 167 623
rect 171 619 172 623
rect 202 621 203 625
rect 207 621 208 625
rect 202 620 208 621
rect 274 621 275 625
rect 279 621 280 625
rect 274 620 280 621
rect 286 623 292 624
rect 166 618 172 619
rect 286 619 287 623
rect 291 619 292 623
rect 378 621 379 625
rect 383 621 384 625
rect 378 620 384 621
rect 390 623 396 624
rect 286 618 292 619
rect 390 619 391 623
rect 395 619 396 623
rect 498 621 499 625
rect 503 621 504 625
rect 498 620 504 621
rect 550 623 556 624
rect 390 618 396 619
rect 550 619 551 623
rect 555 619 556 623
rect 550 618 556 619
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 110 608 116 609
rect 110 595 116 596
rect 110 591 111 595
rect 115 591 116 595
rect 110 590 116 591
rect 134 595 140 596
rect 134 591 135 595
rect 139 591 140 595
rect 134 590 140 591
rect 112 575 114 590
rect 136 575 138 590
rect 168 588 170 618
rect 182 595 188 596
rect 182 591 183 595
rect 187 591 188 595
rect 182 590 188 591
rect 254 595 260 596
rect 254 591 255 595
rect 259 591 260 595
rect 254 590 260 591
rect 166 587 172 588
rect 166 583 167 587
rect 171 583 172 587
rect 166 582 172 583
rect 184 575 186 590
rect 256 575 258 590
rect 288 588 290 618
rect 358 595 364 596
rect 358 591 359 595
rect 363 591 364 595
rect 358 590 364 591
rect 286 587 292 588
rect 286 583 287 587
rect 291 583 292 587
rect 286 582 292 583
rect 360 575 362 590
rect 392 588 394 618
rect 478 595 484 596
rect 478 591 479 595
rect 483 591 484 595
rect 478 590 484 591
rect 390 587 396 588
rect 390 583 391 587
rect 395 583 396 587
rect 390 582 396 583
rect 480 575 482 590
rect 552 588 554 618
rect 606 595 612 596
rect 606 591 607 595
rect 611 591 612 595
rect 606 590 612 591
rect 550 587 556 588
rect 550 583 551 587
rect 555 583 556 587
rect 550 582 556 583
rect 558 587 564 588
rect 558 583 559 587
rect 563 583 564 587
rect 558 582 564 583
rect 111 574 115 575
rect 111 569 115 570
rect 135 574 139 575
rect 135 569 139 570
rect 183 574 187 575
rect 183 569 187 570
rect 239 574 243 575
rect 239 569 243 570
rect 255 574 259 575
rect 255 569 259 570
rect 319 574 323 575
rect 319 569 323 570
rect 359 574 363 575
rect 359 569 363 570
rect 415 574 419 575
rect 415 569 419 570
rect 479 574 483 575
rect 479 569 483 570
rect 519 574 523 575
rect 519 569 523 570
rect 112 554 114 569
rect 136 554 138 569
rect 174 559 180 560
rect 174 555 175 559
rect 179 555 180 559
rect 174 554 180 555
rect 184 554 186 569
rect 230 559 236 560
rect 230 555 231 559
rect 235 555 236 559
rect 230 554 236 555
rect 240 554 242 569
rect 294 559 300 560
rect 294 555 295 559
rect 299 555 300 559
rect 294 554 300 555
rect 320 554 322 569
rect 406 559 412 560
rect 406 555 407 559
rect 411 555 412 559
rect 406 554 412 555
rect 416 554 418 569
rect 458 567 464 568
rect 458 563 459 567
rect 463 563 464 567
rect 458 562 464 563
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 110 548 116 549
rect 134 553 140 554
rect 134 549 135 553
rect 139 549 140 553
rect 134 548 140 549
rect 110 535 116 536
rect 110 531 111 535
rect 115 531 116 535
rect 110 530 116 531
rect 112 511 114 530
rect 143 524 147 525
rect 176 524 178 554
rect 182 553 188 554
rect 182 549 183 553
rect 187 549 188 553
rect 182 548 188 549
rect 232 524 234 554
rect 238 553 244 554
rect 238 549 239 553
rect 243 549 244 553
rect 238 548 244 549
rect 296 524 298 554
rect 318 553 324 554
rect 318 549 319 553
rect 323 549 324 553
rect 318 548 324 549
rect 408 524 410 554
rect 414 553 420 554
rect 414 549 415 553
rect 419 549 420 553
rect 414 548 420 549
rect 142 519 143 524
rect 147 519 148 524
rect 142 518 148 519
rect 154 523 160 524
rect 154 519 155 523
rect 159 519 160 523
rect 154 518 160 519
rect 174 523 180 524
rect 174 519 175 523
rect 179 519 180 523
rect 174 518 180 519
rect 202 523 208 524
rect 202 519 203 523
rect 207 519 208 523
rect 202 518 208 519
rect 230 523 236 524
rect 230 519 231 523
rect 235 519 236 523
rect 230 518 236 519
rect 258 523 264 524
rect 258 519 259 523
rect 263 519 264 523
rect 258 518 264 519
rect 294 523 300 524
rect 294 519 295 523
rect 299 519 300 523
rect 294 518 300 519
rect 338 523 344 524
rect 338 519 339 523
rect 343 519 344 523
rect 338 518 344 519
rect 406 523 412 524
rect 406 519 407 523
rect 411 519 412 523
rect 406 518 412 519
rect 434 523 440 524
rect 434 519 435 523
rect 439 519 440 523
rect 434 518 440 519
rect 156 511 158 518
rect 204 511 206 518
rect 260 511 262 518
rect 340 511 342 518
rect 436 511 438 518
rect 460 512 462 562
rect 510 559 516 560
rect 510 555 511 559
rect 515 555 516 559
rect 510 554 516 555
rect 520 554 522 569
rect 512 524 514 554
rect 518 553 524 554
rect 518 549 519 553
rect 523 549 524 553
rect 518 548 524 549
rect 560 525 562 582
rect 608 575 610 590
rect 607 574 611 575
rect 607 569 611 570
rect 616 564 618 626
rect 626 625 632 626
rect 635 625 639 626
rect 710 627 716 628
rect 626 621 627 625
rect 631 621 632 625
rect 710 623 711 627
rect 715 623 716 627
rect 710 622 716 623
rect 738 625 744 626
rect 775 625 779 626
rect 626 620 632 621
rect 738 621 739 625
rect 743 621 744 625
rect 738 620 744 621
rect 776 614 778 625
rect 774 613 780 614
rect 774 609 775 613
rect 779 609 780 613
rect 774 608 780 609
rect 718 595 724 596
rect 718 591 719 595
rect 723 591 724 595
rect 718 590 724 591
rect 774 595 780 596
rect 774 591 775 595
rect 779 591 780 595
rect 774 590 780 591
rect 720 575 722 590
rect 726 587 732 588
rect 726 583 727 587
rect 731 583 732 587
rect 726 582 732 583
rect 631 574 635 575
rect 631 569 635 570
rect 719 574 723 575
rect 719 569 723 570
rect 614 563 620 564
rect 614 559 615 563
rect 619 559 620 563
rect 614 558 620 559
rect 632 554 634 569
rect 710 559 716 560
rect 710 555 711 559
rect 715 555 716 559
rect 710 554 716 555
rect 720 554 722 569
rect 630 553 636 554
rect 630 549 631 553
rect 635 549 636 553
rect 630 548 636 549
rect 559 524 563 525
rect 510 523 516 524
rect 510 519 511 523
rect 515 519 516 523
rect 510 518 516 519
rect 538 523 544 524
rect 538 519 539 523
rect 543 519 544 523
rect 559 519 563 520
rect 638 523 644 524
rect 638 519 639 523
rect 643 519 644 523
rect 538 518 544 519
rect 638 518 644 519
rect 650 523 656 524
rect 650 519 651 523
rect 655 519 656 523
rect 650 518 656 519
rect 458 511 464 512
rect 540 511 542 518
rect 111 510 115 511
rect 111 505 115 506
rect 155 510 159 511
rect 155 505 159 506
rect 203 510 207 511
rect 203 505 207 506
rect 259 510 263 511
rect 283 510 287 511
rect 331 510 335 511
rect 339 510 343 511
rect 387 510 391 511
rect 435 510 439 511
rect 451 510 455 511
rect 458 507 459 511
rect 463 507 464 511
rect 458 506 464 507
rect 515 510 519 511
rect 539 510 543 511
rect 587 510 591 511
rect 259 505 263 506
rect 282 505 288 506
rect 112 494 114 505
rect 282 501 283 505
rect 287 501 288 505
rect 330 505 336 506
rect 339 505 343 506
rect 386 505 392 506
rect 435 505 439 506
rect 450 505 456 506
rect 282 500 288 501
rect 294 503 300 504
rect 294 499 295 503
rect 299 499 300 503
rect 330 501 331 505
rect 335 501 336 505
rect 330 500 336 501
rect 358 503 364 504
rect 294 498 300 499
rect 358 499 359 503
rect 363 499 364 503
rect 386 501 387 505
rect 391 501 392 505
rect 386 500 392 501
rect 398 503 404 504
rect 358 498 364 499
rect 398 499 399 503
rect 403 499 404 503
rect 450 501 451 505
rect 455 501 456 505
rect 514 505 520 506
rect 539 505 543 506
rect 586 505 592 506
rect 450 500 456 501
rect 462 503 468 504
rect 398 498 404 499
rect 462 499 463 503
rect 467 499 468 503
rect 514 501 515 505
rect 519 501 520 505
rect 514 500 520 501
rect 526 503 532 504
rect 462 498 468 499
rect 526 499 527 503
rect 531 499 532 503
rect 586 501 587 505
rect 591 501 592 505
rect 586 500 592 501
rect 526 498 532 499
rect 110 493 116 494
rect 110 489 111 493
rect 115 489 116 493
rect 110 488 116 489
rect 110 475 116 476
rect 110 471 111 475
rect 115 471 116 475
rect 110 470 116 471
rect 262 475 268 476
rect 262 471 263 475
rect 267 471 268 475
rect 262 470 268 471
rect 112 451 114 470
rect 264 451 266 470
rect 296 468 298 498
rect 310 475 316 476
rect 310 471 311 475
rect 315 471 316 475
rect 310 470 316 471
rect 294 467 300 468
rect 294 463 295 467
rect 299 463 300 467
rect 294 462 300 463
rect 312 451 314 470
rect 360 468 362 498
rect 366 475 372 476
rect 366 471 367 475
rect 371 471 372 475
rect 366 470 372 471
rect 358 467 364 468
rect 358 463 359 467
rect 363 463 364 467
rect 358 462 364 463
rect 368 451 370 470
rect 400 468 402 498
rect 430 475 436 476
rect 430 471 431 475
rect 435 471 436 475
rect 430 470 436 471
rect 398 467 404 468
rect 398 463 399 467
rect 403 463 404 467
rect 398 462 404 463
rect 432 451 434 470
rect 464 468 466 498
rect 494 475 500 476
rect 494 471 495 475
rect 499 471 500 475
rect 494 470 500 471
rect 462 467 468 468
rect 462 463 463 467
rect 467 463 468 467
rect 462 462 468 463
rect 496 451 498 470
rect 528 468 530 498
rect 566 475 572 476
rect 566 471 567 475
rect 571 471 572 475
rect 566 470 572 471
rect 526 467 532 468
rect 526 463 527 467
rect 531 463 532 467
rect 526 462 532 463
rect 534 467 540 468
rect 534 463 535 467
rect 539 463 540 467
rect 534 462 540 463
rect 111 450 115 451
rect 111 445 115 446
rect 263 450 267 451
rect 263 445 267 446
rect 311 450 315 451
rect 311 445 315 446
rect 367 450 371 451
rect 367 445 371 446
rect 415 450 419 451
rect 415 445 419 446
rect 431 450 435 451
rect 431 445 435 446
rect 463 450 467 451
rect 463 445 467 446
rect 495 450 499 451
rect 495 445 499 446
rect 511 450 515 451
rect 511 445 515 446
rect 112 430 114 445
rect 416 430 418 445
rect 454 435 460 436
rect 454 431 455 435
rect 459 431 460 435
rect 454 430 460 431
rect 464 430 466 445
rect 494 439 500 440
rect 494 435 495 439
rect 499 435 500 439
rect 494 434 500 435
rect 110 429 116 430
rect 110 425 111 429
rect 115 425 116 429
rect 110 424 116 425
rect 414 429 420 430
rect 414 425 415 429
rect 419 425 420 429
rect 414 424 420 425
rect 110 411 116 412
rect 110 407 111 411
rect 115 407 116 411
rect 110 406 116 407
rect 112 395 114 406
rect 456 404 458 430
rect 462 429 468 430
rect 462 425 463 429
rect 467 425 468 429
rect 462 424 468 425
rect 454 403 460 404
rect 434 399 440 400
rect 434 395 435 399
rect 439 395 440 399
rect 454 399 455 403
rect 459 399 460 403
rect 496 400 498 434
rect 512 430 514 445
rect 510 429 516 430
rect 510 425 511 429
rect 515 425 516 429
rect 510 424 516 425
rect 536 412 538 462
rect 568 451 570 470
rect 640 468 642 518
rect 652 511 654 518
rect 651 510 655 511
rect 667 510 671 511
rect 712 508 714 554
rect 718 553 724 554
rect 718 549 719 553
rect 723 549 724 553
rect 718 548 724 549
rect 728 524 730 582
rect 776 575 778 590
rect 775 574 779 575
rect 775 569 779 570
rect 776 554 778 569
rect 774 553 780 554
rect 774 549 775 553
rect 779 549 780 553
rect 774 548 780 549
rect 774 535 780 536
rect 774 531 775 535
rect 779 531 780 535
rect 774 530 780 531
rect 726 523 732 524
rect 726 519 727 523
rect 731 519 732 523
rect 726 518 732 519
rect 738 523 744 524
rect 738 519 739 523
rect 743 519 744 523
rect 738 518 744 519
rect 740 511 742 518
rect 776 511 778 530
rect 739 510 743 511
rect 710 507 716 508
rect 651 505 655 506
rect 666 505 672 506
rect 666 501 667 505
rect 671 501 672 505
rect 710 503 711 507
rect 715 503 716 507
rect 775 510 779 511
rect 710 502 716 503
rect 738 505 744 506
rect 775 505 779 506
rect 666 500 672 501
rect 738 501 739 505
rect 743 501 744 505
rect 738 500 744 501
rect 686 499 692 500
rect 686 495 687 499
rect 691 495 692 499
rect 686 494 692 495
rect 776 494 778 505
rect 646 475 652 476
rect 646 471 647 475
rect 651 471 652 475
rect 646 470 652 471
rect 638 467 644 468
rect 638 463 639 467
rect 643 463 644 467
rect 638 462 644 463
rect 648 451 650 470
rect 559 450 563 451
rect 559 445 563 446
rect 567 450 571 451
rect 567 445 571 446
rect 607 450 611 451
rect 607 445 611 446
rect 647 450 651 451
rect 647 445 651 446
rect 655 450 659 451
rect 655 445 659 446
rect 550 435 556 436
rect 550 431 551 435
rect 555 431 556 435
rect 550 430 556 431
rect 560 430 562 445
rect 590 439 596 440
rect 590 435 591 439
rect 595 435 596 439
rect 590 434 596 435
rect 598 435 604 436
rect 534 411 540 412
rect 534 407 535 411
rect 539 407 540 411
rect 534 406 540 407
rect 552 400 554 430
rect 558 429 564 430
rect 558 425 559 429
rect 563 425 564 429
rect 558 424 564 425
rect 592 400 594 434
rect 598 431 599 435
rect 603 431 604 435
rect 598 430 604 431
rect 608 430 610 445
rect 656 430 658 445
rect 688 440 690 494
rect 774 493 780 494
rect 774 489 775 493
rect 779 489 780 493
rect 774 488 780 489
rect 718 475 724 476
rect 718 471 719 475
rect 723 471 724 475
rect 718 470 724 471
rect 774 475 780 476
rect 774 471 775 475
rect 779 471 780 475
rect 774 470 780 471
rect 720 451 722 470
rect 726 467 732 468
rect 726 463 727 467
rect 731 463 732 467
rect 726 462 732 463
rect 711 450 715 451
rect 711 445 715 446
rect 719 450 723 451
rect 719 445 723 446
rect 686 439 692 440
rect 686 435 687 439
rect 691 435 692 439
rect 686 434 692 435
rect 702 435 708 436
rect 702 431 703 435
rect 707 431 708 435
rect 702 430 708 431
rect 712 430 714 445
rect 454 398 460 399
rect 482 399 488 400
rect 482 395 483 399
rect 487 395 488 399
rect 111 394 115 395
rect 307 394 311 395
rect 355 394 359 395
rect 403 394 407 395
rect 434 394 440 395
rect 451 394 455 395
rect 482 394 488 395
rect 494 399 500 400
rect 494 395 495 399
rect 499 395 500 399
rect 530 399 536 400
rect 530 395 531 399
rect 535 395 536 399
rect 494 394 500 395
rect 507 394 511 395
rect 530 394 536 395
rect 550 399 556 400
rect 550 395 551 399
rect 555 395 556 399
rect 578 399 584 400
rect 578 395 579 399
rect 583 395 584 399
rect 550 394 556 395
rect 571 394 575 395
rect 578 394 584 395
rect 590 399 596 400
rect 590 395 591 399
rect 595 395 596 399
rect 590 394 596 395
rect 111 389 115 390
rect 306 389 312 390
rect 112 378 114 389
rect 306 385 307 389
rect 311 385 312 389
rect 354 389 360 390
rect 306 384 312 385
rect 318 387 324 388
rect 318 383 319 387
rect 323 383 324 387
rect 354 385 355 389
rect 359 385 360 389
rect 402 389 408 390
rect 435 389 439 390
rect 450 389 456 390
rect 483 389 487 390
rect 506 389 512 390
rect 531 389 535 390
rect 570 389 576 390
rect 579 389 583 390
rect 354 384 360 385
rect 366 387 372 388
rect 318 382 324 383
rect 366 383 367 387
rect 371 383 372 387
rect 402 385 403 389
rect 407 385 408 389
rect 402 384 408 385
rect 450 385 451 389
rect 455 385 456 389
rect 450 384 456 385
rect 506 385 507 389
rect 511 385 512 389
rect 506 384 512 385
rect 570 385 571 389
rect 575 385 576 389
rect 570 384 576 385
rect 600 384 602 430
rect 606 429 612 430
rect 606 425 607 429
rect 611 425 612 429
rect 606 424 612 425
rect 654 429 660 430
rect 654 425 655 429
rect 659 425 660 429
rect 654 424 660 425
rect 626 399 632 400
rect 626 395 627 399
rect 631 395 632 399
rect 654 399 660 400
rect 654 395 655 399
rect 659 395 660 399
rect 626 394 632 395
rect 643 394 647 395
rect 654 394 660 395
rect 674 399 680 400
rect 674 395 675 399
rect 679 395 680 399
rect 674 394 680 395
rect 627 389 631 390
rect 642 389 648 390
rect 642 385 643 389
rect 647 385 648 389
rect 642 384 648 385
rect 366 382 372 383
rect 470 383 476 384
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 110 372 116 373
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 286 359 292 360
rect 286 355 287 359
rect 291 355 292 359
rect 286 354 292 355
rect 112 339 114 354
rect 288 339 290 354
rect 320 352 322 382
rect 334 359 340 360
rect 334 355 335 359
rect 339 355 340 359
rect 334 354 340 355
rect 318 351 324 352
rect 318 347 319 351
rect 323 347 324 351
rect 318 346 324 347
rect 336 339 338 354
rect 368 352 370 382
rect 422 379 428 380
rect 422 375 423 379
rect 427 375 428 379
rect 470 379 471 383
rect 475 379 476 383
rect 470 378 476 379
rect 526 383 532 384
rect 526 379 527 383
rect 531 379 532 383
rect 526 378 532 379
rect 598 383 604 384
rect 598 379 599 383
rect 603 379 604 383
rect 598 378 604 379
rect 630 383 636 384
rect 630 379 631 383
rect 635 379 636 383
rect 630 378 636 379
rect 422 374 428 375
rect 382 359 388 360
rect 382 355 383 359
rect 387 355 388 359
rect 382 354 388 355
rect 366 351 372 352
rect 366 347 367 351
rect 371 347 372 351
rect 366 346 372 347
rect 384 339 386 354
rect 424 352 426 374
rect 430 359 436 360
rect 430 355 431 359
rect 435 355 436 359
rect 430 354 436 355
rect 406 351 412 352
rect 406 347 407 351
rect 411 347 412 351
rect 406 346 412 347
rect 422 351 428 352
rect 422 347 423 351
rect 427 347 428 351
rect 422 346 428 347
rect 111 338 115 339
rect 111 333 115 334
rect 135 338 139 339
rect 135 333 139 334
rect 215 338 219 339
rect 215 333 219 334
rect 287 338 291 339
rect 287 333 291 334
rect 303 338 307 339
rect 303 333 307 334
rect 335 338 339 339
rect 335 333 339 334
rect 383 338 387 339
rect 383 333 387 334
rect 399 338 403 339
rect 399 333 403 334
rect 112 318 114 333
rect 126 323 132 324
rect 126 319 127 323
rect 131 319 132 323
rect 126 318 132 319
rect 136 318 138 333
rect 182 323 188 324
rect 182 319 183 323
rect 187 319 188 323
rect 182 318 188 319
rect 216 318 218 333
rect 254 323 260 324
rect 254 319 255 323
rect 259 319 260 323
rect 254 318 260 319
rect 304 318 306 333
rect 400 318 402 333
rect 110 317 116 318
rect 110 313 111 317
rect 115 313 116 317
rect 110 312 116 313
rect 110 299 116 300
rect 110 295 111 299
rect 115 295 116 299
rect 110 294 116 295
rect 112 275 114 294
rect 111 274 115 275
rect 128 272 130 318
rect 134 317 140 318
rect 134 313 135 317
rect 139 313 140 317
rect 134 312 140 313
rect 184 296 186 318
rect 214 317 220 318
rect 214 313 215 317
rect 219 313 220 317
rect 214 312 220 313
rect 256 296 258 318
rect 302 317 308 318
rect 302 313 303 317
rect 307 313 308 317
rect 302 312 308 313
rect 398 317 404 318
rect 398 313 399 317
rect 403 313 404 317
rect 398 312 404 313
rect 182 295 188 296
rect 182 291 183 295
rect 187 291 188 295
rect 182 290 188 291
rect 254 295 260 296
rect 254 291 255 295
rect 259 291 260 295
rect 254 290 260 291
rect 408 288 410 346
rect 432 339 434 354
rect 472 352 474 378
rect 486 359 492 360
rect 486 355 487 359
rect 491 355 492 359
rect 486 354 492 355
rect 470 351 476 352
rect 470 347 471 351
rect 475 347 476 351
rect 470 346 476 347
rect 488 339 490 354
rect 528 352 530 378
rect 550 359 556 360
rect 550 355 551 359
rect 555 355 556 359
rect 550 354 556 355
rect 622 359 628 360
rect 622 355 623 359
rect 627 355 628 359
rect 622 354 628 355
rect 526 351 532 352
rect 526 347 527 351
rect 531 347 532 351
rect 526 346 532 347
rect 552 339 554 354
rect 624 339 626 354
rect 431 338 435 339
rect 431 333 435 334
rect 487 338 491 339
rect 487 333 491 334
rect 495 338 499 339
rect 495 333 499 334
rect 551 338 555 339
rect 551 333 555 334
rect 591 338 595 339
rect 591 333 595 334
rect 623 338 627 339
rect 623 333 627 334
rect 496 318 498 333
rect 582 323 588 324
rect 582 319 583 323
rect 587 319 588 323
rect 582 318 588 319
rect 592 318 594 333
rect 632 328 634 378
rect 656 352 658 394
rect 704 392 706 430
rect 710 429 716 430
rect 710 425 711 429
rect 715 425 716 429
rect 710 424 716 425
rect 728 408 730 462
rect 776 451 778 470
rect 775 450 779 451
rect 775 445 779 446
rect 776 430 778 445
rect 774 429 780 430
rect 774 425 775 429
rect 779 425 780 429
rect 774 424 780 425
rect 774 411 780 412
rect 726 407 732 408
rect 726 403 727 407
rect 731 403 732 407
rect 774 407 775 411
rect 779 407 780 411
rect 774 406 780 407
rect 726 402 732 403
rect 730 399 736 400
rect 730 395 731 399
rect 735 395 736 399
rect 776 395 778 406
rect 715 394 719 395
rect 730 394 736 395
rect 775 394 779 395
rect 675 389 679 390
rect 702 391 708 392
rect 702 387 703 391
rect 707 387 708 391
rect 702 386 708 387
rect 714 389 720 390
rect 731 389 735 390
rect 775 389 779 390
rect 714 385 715 389
rect 719 385 720 389
rect 714 384 720 385
rect 776 378 778 389
rect 774 377 780 378
rect 774 373 775 377
rect 779 373 780 377
rect 774 372 780 373
rect 694 359 700 360
rect 694 355 695 359
rect 699 355 700 359
rect 694 354 700 355
rect 774 359 780 360
rect 774 355 775 359
rect 779 355 780 359
rect 774 354 780 355
rect 654 351 660 352
rect 654 347 655 351
rect 659 347 660 351
rect 654 346 660 347
rect 696 339 698 354
rect 702 351 708 352
rect 702 347 703 351
rect 707 347 708 351
rect 702 346 708 347
rect 687 338 691 339
rect 687 333 691 334
rect 695 338 699 339
rect 695 333 699 334
rect 630 327 636 328
rect 630 323 631 327
rect 635 323 636 327
rect 630 322 636 323
rect 688 318 690 333
rect 494 317 500 318
rect 494 313 495 317
rect 499 313 500 317
rect 494 312 500 313
rect 584 288 586 318
rect 590 317 596 318
rect 590 313 591 317
rect 595 313 596 317
rect 590 312 596 313
rect 686 317 692 318
rect 686 313 687 317
rect 691 313 692 317
rect 686 312 692 313
rect 704 296 706 346
rect 776 339 778 354
rect 775 338 779 339
rect 775 333 779 334
rect 726 323 732 324
rect 726 319 727 323
rect 731 319 732 323
rect 726 318 732 319
rect 776 318 778 333
rect 702 295 708 296
rect 702 291 703 295
rect 707 291 708 295
rect 702 290 708 291
rect 154 287 160 288
rect 154 283 155 287
rect 159 283 160 287
rect 154 282 160 283
rect 234 287 240 288
rect 234 283 235 287
rect 239 283 240 287
rect 234 282 240 283
rect 322 287 328 288
rect 322 283 323 287
rect 327 283 328 287
rect 322 282 328 283
rect 406 287 412 288
rect 406 283 407 287
rect 411 283 412 287
rect 406 282 412 283
rect 418 287 424 288
rect 418 283 419 287
rect 423 283 424 287
rect 418 282 424 283
rect 502 287 508 288
rect 502 283 503 287
rect 507 283 508 287
rect 502 282 508 283
rect 514 287 520 288
rect 514 283 515 287
rect 519 283 520 287
rect 514 282 520 283
rect 582 287 588 288
rect 582 283 583 287
rect 587 283 588 287
rect 582 282 588 283
rect 610 287 616 288
rect 610 283 611 287
rect 615 283 616 287
rect 610 282 616 283
rect 706 287 712 288
rect 706 283 707 287
rect 711 283 712 287
rect 706 282 712 283
rect 156 275 158 282
rect 236 275 238 282
rect 324 275 326 282
rect 420 275 422 282
rect 155 274 159 275
rect 111 269 115 270
rect 126 271 132 272
rect 112 258 114 269
rect 126 267 127 271
rect 131 267 132 271
rect 211 274 215 275
rect 235 274 239 275
rect 299 274 303 275
rect 323 274 327 275
rect 387 274 391 275
rect 419 274 423 275
rect 475 274 479 275
rect 126 266 132 267
rect 154 269 160 270
rect 154 265 155 269
rect 159 265 160 269
rect 210 269 216 270
rect 235 269 239 270
rect 298 269 304 270
rect 323 269 327 270
rect 386 269 392 270
rect 419 269 423 270
rect 474 269 480 270
rect 154 264 160 265
rect 166 267 172 268
rect 166 263 167 267
rect 171 263 172 267
rect 210 265 211 269
rect 215 265 216 269
rect 210 264 216 265
rect 222 267 228 268
rect 166 262 172 263
rect 222 263 223 267
rect 227 263 228 267
rect 298 265 299 269
rect 303 265 304 269
rect 298 264 304 265
rect 310 267 316 268
rect 222 262 228 263
rect 310 263 311 267
rect 315 263 316 267
rect 386 265 387 269
rect 391 265 392 269
rect 386 264 392 265
rect 474 265 475 269
rect 479 265 480 269
rect 474 264 480 265
rect 486 267 492 268
rect 310 262 316 263
rect 486 263 487 267
rect 491 263 492 267
rect 486 262 492 263
rect 110 257 116 258
rect 110 253 111 257
rect 115 253 116 257
rect 110 252 116 253
rect 110 239 116 240
rect 110 235 111 239
rect 115 235 116 239
rect 110 234 116 235
rect 134 239 140 240
rect 134 235 135 239
rect 139 235 140 239
rect 134 234 140 235
rect 112 215 114 234
rect 136 215 138 234
rect 168 232 170 262
rect 190 239 196 240
rect 190 235 191 239
rect 195 235 196 239
rect 190 234 196 235
rect 166 231 172 232
rect 166 227 167 231
rect 171 227 172 231
rect 166 226 172 227
rect 192 215 194 234
rect 224 232 226 262
rect 278 239 284 240
rect 278 235 279 239
rect 283 235 284 239
rect 278 234 284 235
rect 222 231 228 232
rect 222 227 223 231
rect 227 227 228 231
rect 222 226 228 227
rect 280 215 282 234
rect 312 232 314 262
rect 366 239 372 240
rect 366 235 367 239
rect 371 235 372 239
rect 366 234 372 235
rect 454 239 460 240
rect 454 235 455 239
rect 459 235 460 239
rect 454 234 460 235
rect 310 231 316 232
rect 310 227 311 231
rect 315 227 316 231
rect 310 226 316 227
rect 368 215 370 234
rect 374 231 380 232
rect 374 227 375 231
rect 379 227 380 231
rect 374 226 380 227
rect 111 214 115 215
rect 111 209 115 210
rect 135 214 139 215
rect 135 209 139 210
rect 183 214 187 215
rect 183 209 187 210
rect 191 214 195 215
rect 191 209 195 210
rect 271 214 275 215
rect 271 209 275 210
rect 279 214 283 215
rect 279 209 283 210
rect 359 214 363 215
rect 359 209 363 210
rect 367 214 371 215
rect 367 209 371 210
rect 112 194 114 209
rect 174 199 180 200
rect 174 195 175 199
rect 179 195 180 199
rect 174 194 180 195
rect 184 194 186 209
rect 234 199 240 200
rect 234 195 235 199
rect 239 195 240 199
rect 234 194 240 195
rect 272 194 274 209
rect 338 199 344 200
rect 338 195 339 199
rect 343 195 344 199
rect 338 194 344 195
rect 360 194 362 209
rect 110 193 116 194
rect 110 189 111 193
rect 115 189 116 193
rect 110 188 116 189
rect 110 175 116 176
rect 110 171 111 175
rect 115 171 116 175
rect 110 170 116 171
rect 112 151 114 170
rect 111 150 115 151
rect 176 148 178 194
rect 182 193 188 194
rect 182 189 183 193
rect 187 189 188 193
rect 182 188 188 189
rect 236 172 238 194
rect 270 193 276 194
rect 270 189 271 193
rect 275 189 276 193
rect 270 188 276 189
rect 340 172 342 194
rect 358 193 364 194
rect 358 189 359 193
rect 363 189 364 193
rect 358 188 364 189
rect 376 172 378 226
rect 456 215 458 234
rect 488 232 490 262
rect 504 232 506 282
rect 516 275 518 282
rect 612 275 614 282
rect 708 275 710 282
rect 515 274 519 275
rect 563 274 567 275
rect 611 274 615 275
rect 651 274 655 275
rect 707 274 711 275
rect 728 272 730 318
rect 774 317 780 318
rect 774 313 775 317
rect 779 313 780 317
rect 774 312 780 313
rect 774 299 780 300
rect 774 295 775 299
rect 779 295 780 299
rect 774 294 780 295
rect 776 275 778 294
rect 739 274 743 275
rect 515 269 519 270
rect 562 269 568 270
rect 611 269 615 270
rect 650 269 656 270
rect 707 269 711 270
rect 726 271 732 272
rect 562 265 563 269
rect 567 265 568 269
rect 562 264 568 265
rect 650 265 651 269
rect 655 265 656 269
rect 726 267 727 271
rect 731 267 732 271
rect 775 274 779 275
rect 726 266 732 267
rect 738 269 744 270
rect 775 269 779 270
rect 650 264 656 265
rect 738 265 739 269
rect 743 265 744 269
rect 738 264 744 265
rect 776 258 778 269
rect 774 257 780 258
rect 774 253 775 257
rect 779 253 780 257
rect 774 252 780 253
rect 542 239 548 240
rect 542 235 543 239
rect 547 235 548 239
rect 542 234 548 235
rect 630 239 636 240
rect 630 235 631 239
rect 635 235 636 239
rect 630 234 636 235
rect 718 239 724 240
rect 718 235 719 239
rect 723 235 724 239
rect 718 234 724 235
rect 774 239 780 240
rect 774 235 775 239
rect 779 235 780 239
rect 774 234 780 235
rect 486 231 492 232
rect 486 227 487 231
rect 491 227 492 231
rect 486 226 492 227
rect 502 231 508 232
rect 502 227 503 231
rect 507 227 508 231
rect 502 226 508 227
rect 544 215 546 234
rect 632 215 634 234
rect 654 231 660 232
rect 654 227 655 231
rect 659 227 660 231
rect 654 226 660 227
rect 455 214 459 215
rect 455 209 459 210
rect 543 214 547 215
rect 543 209 547 210
rect 551 214 555 215
rect 551 209 555 210
rect 631 214 635 215
rect 631 209 635 210
rect 647 214 651 215
rect 647 209 651 210
rect 456 194 458 209
rect 494 199 500 200
rect 494 195 495 199
rect 499 195 500 199
rect 494 194 500 195
rect 552 194 554 209
rect 648 194 650 209
rect 454 193 460 194
rect 454 189 455 193
rect 459 189 460 193
rect 454 188 460 189
rect 496 172 498 194
rect 550 193 556 194
rect 550 189 551 193
rect 555 189 556 193
rect 550 188 556 189
rect 646 193 652 194
rect 646 189 647 193
rect 651 189 652 193
rect 646 188 652 189
rect 234 171 240 172
rect 234 167 235 171
rect 239 167 240 171
rect 234 166 240 167
rect 338 171 344 172
rect 338 167 339 171
rect 343 167 344 171
rect 338 166 344 167
rect 374 171 380 172
rect 374 167 375 171
rect 379 167 380 171
rect 374 166 380 167
rect 494 171 500 172
rect 494 167 495 171
rect 499 167 500 171
rect 494 166 500 167
rect 656 164 658 226
rect 720 215 722 234
rect 776 215 778 234
rect 719 214 723 215
rect 719 209 723 210
rect 775 214 779 215
rect 775 209 779 210
rect 702 199 708 200
rect 702 195 703 199
rect 707 195 708 199
rect 702 194 708 195
rect 710 199 716 200
rect 710 195 711 199
rect 715 195 716 199
rect 710 194 716 195
rect 720 194 722 209
rect 776 194 778 209
rect 704 164 706 194
rect 202 163 208 164
rect 202 159 203 163
rect 207 159 208 163
rect 202 158 208 159
rect 290 163 296 164
rect 290 159 291 163
rect 295 159 296 163
rect 290 158 296 159
rect 378 163 384 164
rect 378 159 379 163
rect 383 159 384 163
rect 378 158 384 159
rect 474 163 480 164
rect 474 159 475 163
rect 479 159 480 163
rect 474 158 480 159
rect 570 163 576 164
rect 570 159 571 163
rect 575 159 576 163
rect 570 158 576 159
rect 654 163 660 164
rect 654 159 655 163
rect 659 159 660 163
rect 654 158 660 159
rect 666 163 672 164
rect 666 159 667 163
rect 671 159 672 163
rect 666 158 672 159
rect 702 163 708 164
rect 702 159 703 163
rect 707 159 708 163
rect 702 158 708 159
rect 204 151 206 158
rect 292 151 294 158
rect 380 151 382 158
rect 476 151 478 158
rect 572 151 574 158
rect 582 155 588 156
rect 582 151 583 155
rect 587 151 588 155
rect 668 151 670 158
rect 203 150 207 151
rect 111 145 115 146
rect 174 147 180 148
rect 112 134 114 145
rect 174 143 175 147
rect 179 143 180 147
rect 211 150 215 151
rect 259 150 263 151
rect 291 150 295 151
rect 307 150 311 151
rect 355 150 359 151
rect 379 150 383 151
rect 403 150 407 151
rect 451 150 455 151
rect 475 150 479 151
rect 499 150 503 151
rect 547 150 551 151
rect 571 150 575 151
rect 582 150 588 151
rect 595 150 599 151
rect 203 145 207 146
rect 210 145 216 146
rect 174 142 180 143
rect 210 141 211 145
rect 215 141 216 145
rect 258 145 264 146
rect 291 145 295 146
rect 306 145 312 146
rect 210 140 216 141
rect 222 143 228 144
rect 222 139 223 143
rect 227 139 228 143
rect 258 141 259 145
rect 263 141 264 145
rect 258 140 264 141
rect 270 143 276 144
rect 222 138 228 139
rect 270 139 271 143
rect 275 139 276 143
rect 306 141 307 145
rect 311 141 312 145
rect 354 145 360 146
rect 379 145 383 146
rect 402 145 408 146
rect 306 140 312 141
rect 318 143 324 144
rect 270 138 276 139
rect 318 139 319 143
rect 323 139 324 143
rect 354 141 355 145
rect 359 141 360 145
rect 354 140 360 141
rect 366 143 372 144
rect 318 138 324 139
rect 366 139 367 143
rect 371 139 372 143
rect 402 141 403 145
rect 407 141 408 145
rect 450 145 456 146
rect 475 145 479 146
rect 498 145 504 146
rect 402 140 408 141
rect 414 143 420 144
rect 366 138 372 139
rect 414 139 415 143
rect 419 139 420 143
rect 450 141 451 145
rect 455 141 456 145
rect 450 140 456 141
rect 462 143 468 144
rect 414 138 420 139
rect 462 139 463 143
rect 467 139 468 143
rect 498 141 499 145
rect 503 141 504 145
rect 546 145 552 146
rect 571 145 575 146
rect 498 140 504 141
rect 510 143 516 144
rect 462 138 468 139
rect 510 139 511 143
rect 515 139 516 143
rect 546 141 547 145
rect 551 141 552 145
rect 546 140 552 141
rect 558 143 564 144
rect 510 138 516 139
rect 558 139 559 143
rect 563 139 564 143
rect 558 138 564 139
rect 110 133 116 134
rect 110 129 111 133
rect 115 129 116 133
rect 110 128 116 129
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 110 110 116 111
rect 190 115 196 116
rect 190 111 191 115
rect 195 111 196 115
rect 190 110 196 111
rect 112 95 114 110
rect 192 95 194 110
rect 224 108 226 138
rect 238 115 244 116
rect 238 111 239 115
rect 243 111 244 115
rect 238 110 244 111
rect 222 107 228 108
rect 222 103 223 107
rect 227 103 228 107
rect 222 102 228 103
rect 240 95 242 110
rect 272 108 274 138
rect 286 115 292 116
rect 286 111 287 115
rect 291 111 292 115
rect 286 110 292 111
rect 270 107 276 108
rect 270 103 271 107
rect 275 103 276 107
rect 270 102 276 103
rect 288 95 290 110
rect 320 108 322 138
rect 334 115 340 116
rect 334 111 335 115
rect 339 111 340 115
rect 334 110 340 111
rect 318 107 324 108
rect 318 103 319 107
rect 323 103 324 107
rect 318 102 324 103
rect 336 95 338 110
rect 368 108 370 138
rect 382 115 388 116
rect 382 111 383 115
rect 387 111 388 115
rect 382 110 388 111
rect 366 107 372 108
rect 366 103 367 107
rect 371 103 372 107
rect 366 102 372 103
rect 384 95 386 110
rect 416 108 418 138
rect 430 115 436 116
rect 430 111 431 115
rect 435 111 436 115
rect 430 110 436 111
rect 414 107 420 108
rect 414 103 415 107
rect 419 103 420 107
rect 414 102 420 103
rect 432 95 434 110
rect 464 108 466 138
rect 478 115 484 116
rect 478 111 479 115
rect 483 111 484 115
rect 478 110 484 111
rect 462 107 468 108
rect 462 103 463 107
rect 467 103 468 107
rect 462 102 468 103
rect 480 95 482 110
rect 512 108 514 138
rect 526 115 532 116
rect 526 111 527 115
rect 531 111 532 115
rect 526 110 532 111
rect 510 107 516 108
rect 510 103 511 107
rect 515 103 516 107
rect 510 102 516 103
rect 528 95 530 110
rect 560 108 562 138
rect 574 115 580 116
rect 574 111 575 115
rect 579 111 580 115
rect 574 110 580 111
rect 558 107 564 108
rect 558 103 559 107
rect 563 103 564 107
rect 558 102 564 103
rect 576 95 578 110
rect 584 108 586 150
rect 643 150 647 151
rect 667 150 671 151
rect 691 150 695 151
rect 712 148 714 194
rect 718 193 724 194
rect 718 189 719 193
rect 723 189 724 193
rect 718 188 724 189
rect 774 193 780 194
rect 774 189 775 193
rect 779 189 780 193
rect 774 188 780 189
rect 774 175 780 176
rect 774 171 775 175
rect 779 171 780 175
rect 774 170 780 171
rect 738 163 744 164
rect 738 159 739 163
rect 743 159 744 163
rect 738 158 744 159
rect 740 151 742 158
rect 776 151 778 170
rect 739 150 743 151
rect 710 147 716 148
rect 594 145 600 146
rect 594 141 595 145
rect 599 141 600 145
rect 594 140 600 141
rect 642 145 648 146
rect 667 145 671 146
rect 690 145 696 146
rect 642 141 643 145
rect 647 141 648 145
rect 642 140 648 141
rect 690 141 691 145
rect 695 141 696 145
rect 710 143 711 147
rect 715 143 716 147
rect 775 150 779 151
rect 710 142 716 143
rect 738 145 744 146
rect 775 145 779 146
rect 690 140 696 141
rect 738 141 739 145
rect 743 141 744 145
rect 738 140 744 141
rect 662 139 668 140
rect 662 135 663 139
rect 667 135 668 139
rect 662 134 668 135
rect 710 139 716 140
rect 710 135 711 139
rect 715 135 716 139
rect 710 134 716 135
rect 776 134 778 145
rect 622 115 628 116
rect 622 111 623 115
rect 627 111 628 115
rect 622 110 628 111
rect 582 107 588 108
rect 582 103 583 107
rect 587 103 588 107
rect 582 102 588 103
rect 624 95 626 110
rect 664 108 666 134
rect 670 115 676 116
rect 670 111 671 115
rect 675 111 676 115
rect 670 110 676 111
rect 662 107 668 108
rect 662 103 663 107
rect 667 103 668 107
rect 662 102 668 103
rect 672 95 674 110
rect 712 108 714 134
rect 774 133 780 134
rect 774 129 775 133
rect 779 129 780 133
rect 774 128 780 129
rect 718 115 724 116
rect 718 111 719 115
rect 723 111 724 115
rect 718 110 724 111
rect 774 115 780 116
rect 774 111 775 115
rect 779 111 780 115
rect 774 110 780 111
rect 710 107 716 108
rect 710 103 711 107
rect 715 103 716 107
rect 710 102 716 103
rect 720 95 722 110
rect 776 95 778 110
rect 111 94 115 95
rect 111 89 115 90
rect 191 94 195 95
rect 191 89 195 90
rect 239 94 243 95
rect 239 89 243 90
rect 287 94 291 95
rect 287 89 291 90
rect 335 94 339 95
rect 335 89 339 90
rect 383 94 387 95
rect 383 89 387 90
rect 431 94 435 95
rect 431 89 435 90
rect 479 94 483 95
rect 479 89 483 90
rect 527 94 531 95
rect 527 89 531 90
rect 575 94 579 95
rect 575 89 579 90
rect 623 94 627 95
rect 623 89 627 90
rect 671 94 675 95
rect 671 89 675 90
rect 719 94 723 95
rect 719 89 723 90
rect 775 94 779 95
rect 775 89 779 90
<< m4c >>
rect 111 858 115 862
rect 155 858 159 862
rect 203 858 207 862
rect 251 858 255 862
rect 299 858 303 862
rect 347 858 351 862
rect 775 858 779 862
rect 111 802 115 806
rect 135 802 139 806
rect 183 802 187 806
rect 231 802 235 806
rect 279 802 283 806
rect 311 802 315 806
rect 327 802 331 806
rect 359 802 363 806
rect 407 802 411 806
rect 455 802 459 806
rect 503 802 507 806
rect 775 802 779 806
rect 111 746 115 750
rect 259 746 263 750
rect 307 746 311 750
rect 331 746 335 750
rect 355 746 359 750
rect 379 746 383 750
rect 403 746 407 750
rect 427 746 431 750
rect 451 746 455 750
rect 475 746 479 750
rect 499 746 503 750
rect 523 746 527 750
rect 547 746 551 750
rect 595 746 599 750
rect 643 746 647 750
rect 691 746 695 750
rect 739 746 743 750
rect 775 746 779 750
rect 111 682 115 686
rect 135 682 139 686
rect 191 682 195 686
rect 239 682 243 686
rect 279 682 283 686
rect 287 682 291 686
rect 335 682 339 686
rect 111 626 115 630
rect 383 682 387 686
rect 431 682 435 686
rect 479 682 483 686
rect 495 682 499 686
rect 527 682 531 686
rect 575 682 579 686
rect 615 682 619 686
rect 623 682 627 686
rect 671 682 675 686
rect 719 682 723 686
rect 155 626 159 630
rect 203 626 207 630
rect 211 626 215 630
rect 275 626 279 630
rect 299 626 303 630
rect 379 626 383 630
rect 403 626 407 630
rect 499 626 503 630
rect 515 626 519 630
rect 627 626 631 630
rect 635 626 639 630
rect 775 682 779 686
rect 111 570 115 574
rect 135 570 139 574
rect 183 570 187 574
rect 239 570 243 574
rect 255 570 259 574
rect 319 570 323 574
rect 359 570 363 574
rect 415 570 419 574
rect 479 570 483 574
rect 519 570 523 574
rect 143 523 147 524
rect 143 520 147 523
rect 607 570 611 574
rect 739 626 743 630
rect 775 626 779 630
rect 631 570 635 574
rect 719 570 723 574
rect 559 520 563 524
rect 111 506 115 510
rect 155 506 159 510
rect 203 506 207 510
rect 259 506 263 510
rect 283 506 287 510
rect 331 506 335 510
rect 339 506 343 510
rect 387 506 391 510
rect 435 506 439 510
rect 451 506 455 510
rect 515 506 519 510
rect 539 506 543 510
rect 587 506 591 510
rect 111 446 115 450
rect 263 446 267 450
rect 311 446 315 450
rect 367 446 371 450
rect 415 446 419 450
rect 431 446 435 450
rect 463 446 467 450
rect 495 446 499 450
rect 511 446 515 450
rect 651 506 655 510
rect 667 506 671 510
rect 775 570 779 574
rect 739 506 743 510
rect 775 506 779 510
rect 559 446 563 450
rect 567 446 571 450
rect 607 446 611 450
rect 647 446 651 450
rect 655 446 659 450
rect 711 446 715 450
rect 719 446 723 450
rect 111 390 115 394
rect 307 390 311 394
rect 355 390 359 394
rect 403 390 407 394
rect 435 390 439 394
rect 451 390 455 394
rect 483 390 487 394
rect 507 390 511 394
rect 531 390 535 394
rect 571 390 575 394
rect 579 390 583 394
rect 627 390 631 394
rect 643 390 647 394
rect 111 334 115 338
rect 135 334 139 338
rect 215 334 219 338
rect 287 334 291 338
rect 303 334 307 338
rect 335 334 339 338
rect 383 334 387 338
rect 399 334 403 338
rect 111 270 115 274
rect 431 334 435 338
rect 487 334 491 338
rect 495 334 499 338
rect 551 334 555 338
rect 591 334 595 338
rect 623 334 627 338
rect 675 390 679 394
rect 775 446 779 450
rect 715 390 719 394
rect 731 390 735 394
rect 775 390 779 394
rect 687 334 691 338
rect 695 334 699 338
rect 775 334 779 338
rect 155 270 159 274
rect 211 270 215 274
rect 235 270 239 274
rect 299 270 303 274
rect 323 270 327 274
rect 387 270 391 274
rect 419 270 423 274
rect 475 270 479 274
rect 111 210 115 214
rect 135 210 139 214
rect 183 210 187 214
rect 191 210 195 214
rect 271 210 275 214
rect 279 210 283 214
rect 359 210 363 214
rect 367 210 371 214
rect 111 146 115 150
rect 515 270 519 274
rect 563 270 567 274
rect 611 270 615 274
rect 651 270 655 274
rect 707 270 711 274
rect 739 270 743 274
rect 775 270 779 274
rect 455 210 459 214
rect 543 210 547 214
rect 551 210 555 214
rect 631 210 635 214
rect 647 210 651 214
rect 719 210 723 214
rect 775 210 779 214
rect 203 146 207 150
rect 211 146 215 150
rect 259 146 263 150
rect 291 146 295 150
rect 307 146 311 150
rect 355 146 359 150
rect 379 146 383 150
rect 403 146 407 150
rect 451 146 455 150
rect 475 146 479 150
rect 499 146 503 150
rect 547 146 551 150
rect 571 146 575 150
rect 595 146 599 150
rect 643 146 647 150
rect 667 146 671 150
rect 691 146 695 150
rect 739 146 743 150
rect 775 146 779 150
rect 111 90 115 94
rect 191 90 195 94
rect 239 90 243 94
rect 287 90 291 94
rect 335 90 339 94
rect 383 90 387 94
rect 431 90 435 94
rect 479 90 483 94
rect 527 90 531 94
rect 575 90 579 94
rect 623 90 627 94
rect 671 90 675 94
rect 719 90 723 94
rect 775 90 779 94
<< m4 >>
rect 96 857 97 863
rect 103 862 811 863
rect 103 858 111 862
rect 115 858 155 862
rect 159 858 203 862
rect 207 858 251 862
rect 255 858 299 862
rect 303 858 347 862
rect 351 858 775 862
rect 779 858 811 862
rect 103 857 811 858
rect 817 857 818 863
rect 84 801 85 807
rect 91 806 799 807
rect 91 802 111 806
rect 115 802 135 806
rect 139 802 183 806
rect 187 802 231 806
rect 235 802 279 806
rect 283 802 311 806
rect 315 802 327 806
rect 331 802 359 806
rect 363 802 407 806
rect 411 802 455 806
rect 459 802 503 806
rect 507 802 775 806
rect 779 802 799 806
rect 91 801 799 802
rect 805 801 806 807
rect 96 745 97 751
rect 103 750 811 751
rect 103 746 111 750
rect 115 746 259 750
rect 263 746 307 750
rect 311 746 331 750
rect 335 746 355 750
rect 359 746 379 750
rect 383 746 403 750
rect 407 746 427 750
rect 431 746 451 750
rect 455 746 475 750
rect 479 746 499 750
rect 503 746 523 750
rect 527 746 547 750
rect 551 746 595 750
rect 599 746 643 750
rect 647 746 691 750
rect 695 746 739 750
rect 743 746 775 750
rect 779 746 811 750
rect 103 745 811 746
rect 817 745 818 751
rect 84 681 85 687
rect 91 686 799 687
rect 91 682 111 686
rect 115 682 135 686
rect 139 682 191 686
rect 195 682 239 686
rect 243 682 279 686
rect 283 682 287 686
rect 291 682 335 686
rect 339 682 383 686
rect 387 682 431 686
rect 435 682 479 686
rect 483 682 495 686
rect 499 682 527 686
rect 531 682 575 686
rect 579 682 615 686
rect 619 682 623 686
rect 627 682 671 686
rect 675 682 719 686
rect 723 682 775 686
rect 779 682 799 686
rect 91 681 799 682
rect 805 681 806 687
rect 96 625 97 631
rect 103 630 811 631
rect 103 626 111 630
rect 115 626 155 630
rect 159 626 203 630
rect 207 626 211 630
rect 215 626 275 630
rect 279 626 299 630
rect 303 626 379 630
rect 383 626 403 630
rect 407 626 499 630
rect 503 626 515 630
rect 519 626 627 630
rect 631 626 635 630
rect 639 626 739 630
rect 743 626 775 630
rect 779 626 811 630
rect 103 625 811 626
rect 817 625 818 631
rect 84 569 85 575
rect 91 574 799 575
rect 91 570 111 574
rect 115 570 135 574
rect 139 570 183 574
rect 187 570 239 574
rect 243 570 255 574
rect 259 570 319 574
rect 323 570 359 574
rect 363 570 415 574
rect 419 570 479 574
rect 483 570 519 574
rect 523 570 607 574
rect 611 570 631 574
rect 635 570 719 574
rect 723 570 775 574
rect 779 570 799 574
rect 91 569 799 570
rect 805 569 806 575
rect 142 524 148 525
rect 558 524 564 525
rect 142 520 143 524
rect 147 520 559 524
rect 563 520 564 524
rect 142 519 148 520
rect 558 519 564 520
rect 96 505 97 511
rect 103 510 811 511
rect 103 506 111 510
rect 115 506 155 510
rect 159 506 203 510
rect 207 506 259 510
rect 263 506 283 510
rect 287 506 331 510
rect 335 506 339 510
rect 343 506 387 510
rect 391 506 435 510
rect 439 506 451 510
rect 455 506 515 510
rect 519 506 539 510
rect 543 506 587 510
rect 591 506 651 510
rect 655 506 667 510
rect 671 506 739 510
rect 743 506 775 510
rect 779 506 811 510
rect 103 505 811 506
rect 817 505 818 511
rect 84 445 85 451
rect 91 450 799 451
rect 91 446 111 450
rect 115 446 263 450
rect 267 446 311 450
rect 315 446 367 450
rect 371 446 415 450
rect 419 446 431 450
rect 435 446 463 450
rect 467 446 495 450
rect 499 446 511 450
rect 515 446 559 450
rect 563 446 567 450
rect 571 446 607 450
rect 611 446 647 450
rect 651 446 655 450
rect 659 446 711 450
rect 715 446 719 450
rect 723 446 775 450
rect 779 446 799 450
rect 91 445 799 446
rect 805 445 806 451
rect 96 389 97 395
rect 103 394 811 395
rect 103 390 111 394
rect 115 390 307 394
rect 311 390 355 394
rect 359 390 403 394
rect 407 390 435 394
rect 439 390 451 394
rect 455 390 483 394
rect 487 390 507 394
rect 511 390 531 394
rect 535 390 571 394
rect 575 390 579 394
rect 583 390 627 394
rect 631 390 643 394
rect 647 390 675 394
rect 679 390 715 394
rect 719 390 731 394
rect 735 390 775 394
rect 779 390 811 394
rect 103 389 811 390
rect 817 389 818 395
rect 84 333 85 339
rect 91 338 799 339
rect 91 334 111 338
rect 115 334 135 338
rect 139 334 215 338
rect 219 334 287 338
rect 291 334 303 338
rect 307 334 335 338
rect 339 334 383 338
rect 387 334 399 338
rect 403 334 431 338
rect 435 334 487 338
rect 491 334 495 338
rect 499 334 551 338
rect 555 334 591 338
rect 595 334 623 338
rect 627 334 687 338
rect 691 334 695 338
rect 699 334 775 338
rect 779 334 799 338
rect 91 333 799 334
rect 805 333 806 339
rect 96 269 97 275
rect 103 274 811 275
rect 103 270 111 274
rect 115 270 155 274
rect 159 270 211 274
rect 215 270 235 274
rect 239 270 299 274
rect 303 270 323 274
rect 327 270 387 274
rect 391 270 419 274
rect 423 270 475 274
rect 479 270 515 274
rect 519 270 563 274
rect 567 270 611 274
rect 615 270 651 274
rect 655 270 707 274
rect 711 270 739 274
rect 743 270 775 274
rect 779 270 811 274
rect 103 269 811 270
rect 817 269 818 275
rect 84 209 85 215
rect 91 214 799 215
rect 91 210 111 214
rect 115 210 135 214
rect 139 210 183 214
rect 187 210 191 214
rect 195 210 271 214
rect 275 210 279 214
rect 283 210 359 214
rect 363 210 367 214
rect 371 210 455 214
rect 459 210 543 214
rect 547 210 551 214
rect 555 210 631 214
rect 635 210 647 214
rect 651 210 719 214
rect 723 210 775 214
rect 779 210 799 214
rect 91 209 799 210
rect 805 209 806 215
rect 96 145 97 151
rect 103 150 811 151
rect 103 146 111 150
rect 115 146 203 150
rect 207 146 211 150
rect 215 146 259 150
rect 263 146 291 150
rect 295 146 307 150
rect 311 146 355 150
rect 359 146 379 150
rect 383 146 403 150
rect 407 146 451 150
rect 455 146 475 150
rect 479 146 499 150
rect 503 146 547 150
rect 551 146 571 150
rect 575 146 595 150
rect 599 146 643 150
rect 647 146 667 150
rect 671 146 691 150
rect 695 146 739 150
rect 743 146 775 150
rect 779 146 811 150
rect 103 145 811 146
rect 817 145 818 151
rect 84 89 85 95
rect 91 94 799 95
rect 91 90 111 94
rect 115 90 191 94
rect 195 90 239 94
rect 243 90 287 94
rect 291 90 335 94
rect 339 90 383 94
rect 387 90 431 94
rect 435 90 479 94
rect 483 90 527 94
rect 531 90 575 94
rect 579 90 623 94
rect 627 90 671 94
rect 675 90 719 94
rect 723 90 775 94
rect 779 90 799 94
rect 91 89 799 90
rect 805 89 806 95
<< m5c >>
rect 97 857 103 863
rect 811 857 817 863
rect 85 801 91 807
rect 799 801 805 807
rect 97 745 103 751
rect 811 745 817 751
rect 85 681 91 687
rect 799 681 805 687
rect 97 625 103 631
rect 811 625 817 631
rect 85 569 91 575
rect 799 569 805 575
rect 97 505 103 511
rect 811 505 817 511
rect 85 445 91 451
rect 799 445 805 451
rect 97 389 103 395
rect 811 389 817 395
rect 85 333 91 339
rect 799 333 805 339
rect 97 269 103 275
rect 811 269 817 275
rect 85 209 91 215
rect 799 209 805 215
rect 97 145 103 151
rect 811 145 817 151
rect 85 89 91 95
rect 799 89 805 95
<< m5 >>
rect 84 807 92 864
rect 84 801 85 807
rect 91 801 92 807
rect 84 687 92 801
rect 84 681 85 687
rect 91 681 92 687
rect 84 575 92 681
rect 84 569 85 575
rect 91 569 92 575
rect 84 451 92 569
rect 84 445 85 451
rect 91 445 92 451
rect 84 339 92 445
rect 84 333 85 339
rect 91 333 92 339
rect 84 215 92 333
rect 84 209 85 215
rect 91 209 92 215
rect 84 95 92 209
rect 84 89 85 95
rect 91 89 92 95
rect 84 72 92 89
rect 96 863 104 864
rect 96 857 97 863
rect 103 857 104 863
rect 96 751 104 857
rect 96 745 97 751
rect 103 745 104 751
rect 96 631 104 745
rect 96 625 97 631
rect 103 625 104 631
rect 96 511 104 625
rect 96 505 97 511
rect 103 505 104 511
rect 96 395 104 505
rect 96 389 97 395
rect 103 389 104 395
rect 96 275 104 389
rect 96 269 97 275
rect 103 269 104 275
rect 96 151 104 269
rect 96 145 97 151
rect 103 145 104 151
rect 96 72 104 145
rect 798 807 806 864
rect 798 801 799 807
rect 805 801 806 807
rect 798 687 806 801
rect 798 681 799 687
rect 805 681 806 687
rect 798 575 806 681
rect 798 569 799 575
rect 805 569 806 575
rect 798 451 806 569
rect 798 445 799 451
rect 805 445 806 451
rect 798 339 806 445
rect 798 333 799 339
rect 805 333 806 339
rect 798 215 806 333
rect 798 209 799 215
rect 805 209 806 215
rect 798 95 806 209
rect 798 89 799 95
rect 805 89 806 95
rect 798 72 806 89
rect 810 863 818 864
rect 810 857 811 863
rect 817 857 818 863
rect 810 751 818 857
rect 810 745 811 751
rect 817 745 818 751
rect 810 631 818 745
rect 810 625 811 631
rect 817 625 818 631
rect 810 511 818 625
rect 810 505 811 511
rect 817 505 818 511
rect 810 395 818 505
rect 810 389 811 395
rect 817 389 818 395
rect 810 275 818 389
rect 810 269 811 275
rect 817 269 818 275
rect 810 151 818 269
rect 810 145 811 151
rect 817 145 818 151
rect 810 72 818 145
use welltap_svt  __well_tap__0
timestamp 1730593880
transform 1 0 104 0 1 108
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730593880
transform 1 0 104 0 1 108
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0OR2X1  or_561_6
timestamp 1730593880
transform 1 0 184 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_561_6
timestamp 1730593880
transform 1 0 184 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_562_6
timestamp 1730593880
transform 1 0 232 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_562_6
timestamp 1730593880
transform 1 0 232 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_563_6
timestamp 1730593880
transform 1 0 280 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_563_6
timestamp 1730593880
transform 1 0 280 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_564_6
timestamp 1730593880
transform 1 0 328 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_564_6
timestamp 1730593880
transform 1 0 328 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_565_6
timestamp 1730593880
transform 1 0 376 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_565_6
timestamp 1730593880
transform 1 0 376 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_566_6
timestamp 1730593880
transform 1 0 424 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_566_6
timestamp 1730593880
transform 1 0 424 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_567_6
timestamp 1730593880
transform 1 0 472 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_567_6
timestamp 1730593880
transform 1 0 472 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_568_6
timestamp 1730593880
transform 1 0 520 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_568_6
timestamp 1730593880
transform 1 0 520 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_569_6
timestamp 1730593880
transform 1 0 568 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_569_6
timestamp 1730593880
transform 1 0 568 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_599_6
timestamp 1730593880
transform 1 0 616 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_599_6
timestamp 1730593880
transform 1 0 616 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_598_6
timestamp 1730593880
transform 1 0 664 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_598_6
timestamp 1730593880
transform 1 0 664 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_597_6
timestamp 1730593880
transform 1 0 712 0 1 92
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_597_6
timestamp 1730593880
transform 1 0 712 0 1 92
box 7 3 44 54
use welltap_svt  __well_tap__1
timestamp 1730593880
transform 1 0 768 0 1 108
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730593880
transform 1 0 768 0 1 108
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730593880
transform 1 0 104 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730593880
transform 1 0 104 0 -1 196
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_560_6
timestamp 1730593880
transform 1 0 176 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_560_6
timestamp 1730593880
transform 1 0 176 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_559_6
timestamp 1730593880
transform 1 0 264 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_559_6
timestamp 1730593880
transform 1 0 264 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_558_6
timestamp 1730593880
transform 1 0 352 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_558_6
timestamp 1730593880
transform 1 0 352 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_571_6
timestamp 1730593880
transform 1 0 448 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_571_6
timestamp 1730593880
transform 1 0 448 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_570_6
timestamp 1730593880
transform 1 0 544 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_570_6
timestamp 1730593880
transform 1 0 544 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_595_6
timestamp 1730593880
transform 1 0 640 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_595_6
timestamp 1730593880
transform 1 0 640 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_596_6
timestamp 1730593880
transform 1 0 712 0 -1 212
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_596_6
timestamp 1730593880
transform 1 0 712 0 -1 212
box 7 3 44 54
use welltap_svt  __well_tap__3
timestamp 1730593880
transform 1 0 768 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730593880
transform 1 0 768 0 -1 196
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_554_6
timestamp 1730593880
transform 1 0 128 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_554_6
timestamp 1730593880
transform 1 0 128 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_555_6
timestamp 1730593880
transform 1 0 184 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_555_6
timestamp 1730593880
transform 1 0 184 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_556_6
timestamp 1730593880
transform 1 0 272 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_556_6
timestamp 1730593880
transform 1 0 272 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_557_6
timestamp 1730593880
transform 1 0 360 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_557_6
timestamp 1730593880
transform 1 0 360 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_572_6
timestamp 1730593880
transform 1 0 448 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_572_6
timestamp 1730593880
transform 1 0 448 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_573_6
timestamp 1730593880
transform 1 0 536 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_573_6
timestamp 1730593880
transform 1 0 536 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_594_6
timestamp 1730593880
transform 1 0 624 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_594_6
timestamp 1730593880
transform 1 0 624 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_593_6
timestamp 1730593880
transform 1 0 712 0 1 216
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_593_6
timestamp 1730593880
transform 1 0 712 0 1 216
box 7 3 44 54
use welltap_svt  __well_tap__4
timestamp 1730593880
transform 1 0 104 0 1 232
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730593880
transform 1 0 104 0 1 232
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730593880
transform 1 0 768 0 1 232
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730593880
transform 1 0 768 0 1 232
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730593880
transform 1 0 104 0 -1 320
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730593880
transform 1 0 104 0 -1 320
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_553_6
timestamp 1730593880
transform 1 0 128 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_553_6
timestamp 1730593880
transform 1 0 128 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_552_6
timestamp 1730593880
transform 1 0 208 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_552_6
timestamp 1730593880
transform 1 0 208 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_551_6
timestamp 1730593880
transform 1 0 296 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_551_6
timestamp 1730593880
transform 1 0 296 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_550_6
timestamp 1730593880
transform 1 0 392 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_550_6
timestamp 1730593880
transform 1 0 392 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_574_6
timestamp 1730593880
transform 1 0 488 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_574_6
timestamp 1730593880
transform 1 0 488 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_575_6
timestamp 1730593880
transform 1 0 584 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_575_6
timestamp 1730593880
transform 1 0 584 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_592_6
timestamp 1730593880
transform 1 0 680 0 -1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_592_6
timestamp 1730593880
transform 1 0 680 0 -1 336
box 7 3 44 54
use welltap_svt  __well_tap__7
timestamp 1730593880
transform 1 0 768 0 -1 320
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730593880
transform 1 0 768 0 -1 320
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730593880
transform 1 0 104 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730593880
transform 1 0 104 0 1 352
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_547_6
timestamp 1730593880
transform 1 0 280 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_547_6
timestamp 1730593880
transform 1 0 280 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_548_6
timestamp 1730593880
transform 1 0 328 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_548_6
timestamp 1730593880
transform 1 0 328 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_549_6
timestamp 1730593880
transform 1 0 376 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_549_6
timestamp 1730593880
transform 1 0 376 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_546_6
timestamp 1730593880
transform 1 0 424 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_546_6
timestamp 1730593880
transform 1 0 424 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_545_6
timestamp 1730593880
transform 1 0 480 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_545_6
timestamp 1730593880
transform 1 0 480 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_544_6
timestamp 1730593880
transform 1 0 544 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_544_6
timestamp 1730593880
transform 1 0 544 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_576_6
timestamp 1730593880
transform 1 0 616 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_576_6
timestamp 1730593880
transform 1 0 616 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_591_6
timestamp 1730593880
transform 1 0 688 0 1 336
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_591_6
timestamp 1730593880
transform 1 0 688 0 1 336
box 7 3 44 54
use welltap_svt  __well_tap__9
timestamp 1730593880
transform 1 0 768 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730593880
transform 1 0 768 0 1 352
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730593880
transform 1 0 104 0 -1 432
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730593880
transform 1 0 104 0 -1 432
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_539_6
timestamp 1730593880
transform 1 0 408 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_539_6
timestamp 1730593880
transform 1 0 408 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_540_6
timestamp 1730593880
transform 1 0 456 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_540_6
timestamp 1730593880
transform 1 0 456 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_541_6
timestamp 1730593880
transform 1 0 504 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_541_6
timestamp 1730593880
transform 1 0 504 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_542_6
timestamp 1730593880
transform 1 0 552 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_542_6
timestamp 1730593880
transform 1 0 552 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_543_6
timestamp 1730593880
transform 1 0 600 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_543_6
timestamp 1730593880
transform 1 0 600 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_577_6
timestamp 1730593880
transform 1 0 648 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_577_6
timestamp 1730593880
transform 1 0 648 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_590_6
timestamp 1730593880
transform 1 0 704 0 -1 448
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_590_6
timestamp 1730593880
transform 1 0 704 0 -1 448
box 7 3 44 54
use welltap_svt  __well_tap__11
timestamp 1730593880
transform 1 0 768 0 -1 432
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730593880
transform 1 0 768 0 -1 432
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730593880
transform 1 0 104 0 1 468
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730593880
transform 1 0 104 0 1 468
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_533_6
timestamp 1730593880
transform 1 0 256 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_533_6
timestamp 1730593880
transform 1 0 256 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_534_6
timestamp 1730593880
transform 1 0 304 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_534_6
timestamp 1730593880
transform 1 0 304 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_535_6
timestamp 1730593880
transform 1 0 360 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_535_6
timestamp 1730593880
transform 1 0 360 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_536_6
timestamp 1730593880
transform 1 0 424 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_536_6
timestamp 1730593880
transform 1 0 424 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_537_6
timestamp 1730593880
transform 1 0 488 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_537_6
timestamp 1730593880
transform 1 0 488 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_538_6
timestamp 1730593880
transform 1 0 560 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_538_6
timestamp 1730593880
transform 1 0 560 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_578_6
timestamp 1730593880
transform 1 0 640 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_578_6
timestamp 1730593880
transform 1 0 640 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_589_6
timestamp 1730593880
transform 1 0 712 0 1 452
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_589_6
timestamp 1730593880
transform 1 0 712 0 1 452
box 7 3 44 54
use welltap_svt  __well_tap__13
timestamp 1730593880
transform 1 0 768 0 1 468
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730593880
transform 1 0 768 0 1 468
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730593880
transform 1 0 104 0 -1 556
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730593880
transform 1 0 104 0 -1 556
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_527_6
timestamp 1730593880
transform 1 0 128 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_527_6
timestamp 1730593880
transform 1 0 128 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_528_6
timestamp 1730593880
transform 1 0 176 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_528_6
timestamp 1730593880
transform 1 0 176 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_529_6
timestamp 1730593880
transform 1 0 232 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_529_6
timestamp 1730593880
transform 1 0 232 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_530_6
timestamp 1730593880
transform 1 0 312 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_530_6
timestamp 1730593880
transform 1 0 312 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_531_6
timestamp 1730593880
transform 1 0 408 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_531_6
timestamp 1730593880
transform 1 0 408 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_532_6
timestamp 1730593880
transform 1 0 512 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_532_6
timestamp 1730593880
transform 1 0 512 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_579_6
timestamp 1730593880
transform 1 0 624 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_579_6
timestamp 1730593880
transform 1 0 624 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_588_6
timestamp 1730593880
transform 1 0 712 0 -1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_588_6
timestamp 1730593880
transform 1 0 712 0 -1 572
box 7 3 44 54
use welltap_svt  __well_tap__15
timestamp 1730593880
transform 1 0 768 0 -1 556
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730593880
transform 1 0 768 0 -1 556
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_521_6
timestamp 1730593880
transform 1 0 128 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_521_6
timestamp 1730593880
transform 1 0 128 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_522_6
timestamp 1730593880
transform 1 0 176 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_522_6
timestamp 1730593880
transform 1 0 176 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_523_6
timestamp 1730593880
transform 1 0 248 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_523_6
timestamp 1730593880
transform 1 0 248 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_524_6
timestamp 1730593880
transform 1 0 352 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_524_6
timestamp 1730593880
transform 1 0 352 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_525_6
timestamp 1730593880
transform 1 0 472 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_525_6
timestamp 1730593880
transform 1 0 472 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_526_6
timestamp 1730593880
transform 1 0 600 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_526_6
timestamp 1730593880
transform 1 0 600 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_587_6
timestamp 1730593880
transform 1 0 712 0 1 572
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_587_6
timestamp 1730593880
transform 1 0 712 0 1 572
box 7 3 44 54
use welltap_svt  __well_tap__16
timestamp 1730593880
transform 1 0 104 0 1 588
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730593880
transform 1 0 104 0 1 588
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_520_6
timestamp 1730593880
transform 1 0 128 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_520_6
timestamp 1730593880
transform 1 0 128 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_519_6
timestamp 1730593880
transform 1 0 184 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_519_6
timestamp 1730593880
transform 1 0 184 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_518_6
timestamp 1730593880
transform 1 0 272 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_518_6
timestamp 1730593880
transform 1 0 272 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_516_6
timestamp 1730593880
transform 1 0 376 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_516_6
timestamp 1730593880
transform 1 0 376 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_517_6
timestamp 1730593880
transform 1 0 488 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_517_6
timestamp 1730593880
transform 1 0 488 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_580_6
timestamp 1730593880
transform 1 0 608 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_580_6
timestamp 1730593880
transform 1 0 608 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_586_6
timestamp 1730593880
transform 1 0 712 0 -1 684
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_586_6
timestamp 1730593880
transform 1 0 712 0 -1 684
box 7 3 44 54
use welltap_svt  __well_tap__17
timestamp 1730593880
transform 1 0 768 0 1 588
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730593880
transform 1 0 768 0 1 588
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730593880
transform 1 0 104 0 -1 668
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730593880
transform 1 0 104 0 -1 668
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_513_6
timestamp 1730593880
transform 1 0 232 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_513_6
timestamp 1730593880
transform 1 0 232 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_514_6
timestamp 1730593880
transform 1 0 280 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_514_6
timestamp 1730593880
transform 1 0 280 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_515_6
timestamp 1730593880
transform 1 0 328 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_515_6
timestamp 1730593880
transform 1 0 328 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_512_6
timestamp 1730593880
transform 1 0 376 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_512_6
timestamp 1730593880
transform 1 0 376 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_511_6
timestamp 1730593880
transform 1 0 424 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_511_6
timestamp 1730593880
transform 1 0 424 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_510_6
timestamp 1730593880
transform 1 0 472 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_510_6
timestamp 1730593880
transform 1 0 472 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_581_6
timestamp 1730593880
transform 1 0 520 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_581_6
timestamp 1730593880
transform 1 0 520 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_582_6
timestamp 1730593880
transform 1 0 568 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_582_6
timestamp 1730593880
transform 1 0 568 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_583_6
timestamp 1730593880
transform 1 0 616 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_583_6
timestamp 1730593880
transform 1 0 616 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_584_6
timestamp 1730593880
transform 1 0 664 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_584_6
timestamp 1730593880
transform 1 0 664 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_585_6
timestamp 1730593880
transform 1 0 712 0 1 692
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_585_6
timestamp 1730593880
transform 1 0 712 0 1 692
box 7 3 44 54
use welltap_svt  __well_tap__19
timestamp 1730593880
transform 1 0 768 0 -1 668
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730593880
transform 1 0 768 0 -1 668
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730593880
transform 1 0 104 0 1 708
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730593880
transform 1 0 104 0 1 708
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730593880
transform 1 0 768 0 1 708
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730593880
transform 1 0 768 0 1 708
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730593880
transform 1 0 104 0 -1 788
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730593880
transform 1 0 104 0 -1 788
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_55_6
timestamp 1730593880
transform 1 0 304 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_55_6
timestamp 1730593880
transform 1 0 304 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_56_6
timestamp 1730593880
transform 1 0 352 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_56_6
timestamp 1730593880
transform 1 0 352 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_57_6
timestamp 1730593880
transform 1 0 400 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_57_6
timestamp 1730593880
transform 1 0 400 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_58_6
timestamp 1730593880
transform 1 0 448 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_58_6
timestamp 1730593880
transform 1 0 448 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_59_6
timestamp 1730593880
transform 1 0 496 0 -1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_59_6
timestamp 1730593880
transform 1 0 496 0 -1 804
box 7 3 44 54
use welltap_svt  __well_tap__23
timestamp 1730593880
transform 1 0 768 0 -1 788
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730593880
transform 1 0 768 0 -1 788
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730593880
transform 1 0 104 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730593880
transform 1 0 104 0 1 820
box 8 4 12 24
use _0_0std_0_0cells_0_0OR2X1  or_50_6
timestamp 1730593880
transform 1 0 128 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_50_6
timestamp 1730593880
transform 1 0 128 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_51_6
timestamp 1730593880
transform 1 0 176 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_51_6
timestamp 1730593880
transform 1 0 176 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_52_6
timestamp 1730593880
transform 1 0 224 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_52_6
timestamp 1730593880
transform 1 0 224 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_53_6
timestamp 1730593880
transform 1 0 272 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_53_6
timestamp 1730593880
transform 1 0 272 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_54_6
timestamp 1730593880
transform 1 0 320 0 1 804
box 7 3 44 54
use _0_0std_0_0cells_0_0OR2X1  or_54_6
timestamp 1730593880
transform 1 0 320 0 1 804
box 7 3 44 54
use welltap_svt  __well_tap__25
timestamp 1730593880
transform 1 0 768 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730593880
transform 1 0 768 0 1 820
box 8 4 12 24
<< end >>
