magic
tech TSMC180
timestamp 1734144021
<< m1 >>
rect 1462 4497 1466 4500
rect 2866 4497 2870 4500
rect 4269 4018 4272 4022
rect 4269 3538 4272 3542
rect 4269 3058 4272 3062
rect 4269 2578 4272 2582
rect 4269 2098 4272 2102
rect 4269 1618 4272 1622
rect 4269 1138 4272 1142
rect 4269 658 4272 662
rect 250 180 254 183
rect 442 180 446 183
rect 634 180 638 183
rect 826 180 830 183
rect 1018 180 1022 183
rect 1204 180 1208 183
rect 1396 180 1400 183
rect 1588 180 1592 183
rect 1780 180 1784 183
rect 1972 180 1976 183
rect 2164 180 2168 183
rect 2356 180 2360 183
rect 2548 180 2552 183
rect 2740 180 2744 183
rect 2932 180 2936 183
rect 3124 180 3128 183
rect 3310 180 3314 183
rect 3502 180 3506 183
rect 3694 180 3698 183
rect 3886 180 3890 183
rect 4078 180 4082 183
use welltap_svt  __well_tap__0
timestamp 1734143631
transform 1 0 72 0 1 230
box 6 10 9 20
use welltap_svt  __well_tap__1
timestamp 1734143631
transform 1 0 4230 0 1 230
box 6 10 9 20
use welltap_svt  __well_tap__2
timestamp 1734143631
transform 1 0 72 0 -1 440
box 6 10 9 20
use welltap_svt  __well_tap__3
timestamp 1734143631
transform 1 0 4230 0 -1 440
box 6 10 9 20
use welltap_svt  __well_tap__4
timestamp 1734143631
transform 1 0 72 0 1 500
box 6 10 9 20
use welltap_svt  __well_tap__5
timestamp 1734143631
transform 1 0 4230 0 1 500
box 6 10 9 20
use welltap_svt  __well_tap__6
timestamp 1734143631
transform 1 0 72 0 -1 680
box 6 10 9 20
use welltap_svt  __well_tap__7
timestamp 1734143631
transform 1 0 4230 0 -1 680
box 6 10 9 20
use welltap_svt  __well_tap__8
timestamp 1734143631
transform 1 0 72 0 1 740
box 6 10 9 20
use welltap_svt  __well_tap__9
timestamp 1734143631
transform 1 0 4230 0 1 740
box 6 10 9 20
use welltap_svt  __well_tap__10
timestamp 1734143631
transform 1 0 72 0 -1 920
box 6 10 9 20
use welltap_svt  __well_tap__11
timestamp 1734143631
transform 1 0 4230 0 -1 920
box 6 10 9 20
use welltap_svt  __well_tap__12
timestamp 1734143631
transform 1 0 72 0 1 980
box 6 10 9 20
use welltap_svt  __well_tap__13
timestamp 1734143631
transform 1 0 4230 0 1 980
box 6 10 9 20
use welltap_svt  __well_tap__14
timestamp 1734143631
transform 1 0 72 0 -1 1160
box 6 10 9 20
use welltap_svt  __well_tap__15
timestamp 1734143631
transform 1 0 4230 0 -1 1160
box 6 10 9 20
use welltap_svt  __well_tap__16
timestamp 1734143631
transform 1 0 72 0 1 1220
box 6 10 9 20
use welltap_svt  __well_tap__17
timestamp 1734143631
transform 1 0 4230 0 1 1220
box 6 10 9 20
use welltap_svt  __well_tap__18
timestamp 1734143631
transform 1 0 72 0 -1 1390
box 6 10 9 20
use welltap_svt  __well_tap__19
timestamp 1734143631
transform 1 0 4230 0 -1 1390
box 6 10 9 20
use welltap_svt  __well_tap__20
timestamp 1734143631
transform 1 0 72 0 1 1450
box 6 10 9 20
use welltap_svt  __well_tap__21
timestamp 1734143631
transform 1 0 4230 0 1 1450
box 6 10 9 20
use welltap_svt  __well_tap__22
timestamp 1734143631
transform 1 0 72 0 -1 1630
box 6 10 9 20
use welltap_svt  __well_tap__23
timestamp 1734143631
transform 1 0 4230 0 -1 1630
box 6 10 9 20
use welltap_svt  __well_tap__24
timestamp 1734143631
transform 1 0 72 0 1 1690
box 6 10 9 20
use welltap_svt  __well_tap__25
timestamp 1734143631
transform 1 0 4230 0 1 1690
box 6 10 9 20
use welltap_svt  __well_tap__26
timestamp 1734143631
transform 1 0 72 0 -1 1870
box 6 10 9 20
use welltap_svt  __well_tap__27
timestamp 1734143631
transform 1 0 4230 0 -1 1870
box 6 10 9 20
use welltap_svt  __well_tap__28
timestamp 1734143631
transform 1 0 72 0 1 1930
box 6 10 9 20
use welltap_svt  __well_tap__29
timestamp 1734143631
transform 1 0 4230 0 1 1930
box 6 10 9 20
use welltap_svt  __well_tap__30
timestamp 1734143631
transform 1 0 72 0 -1 2100
box 6 10 9 20
use welltap_svt  __well_tap__31
timestamp 1734143631
transform 1 0 4230 0 -1 2100
box 6 10 9 20
use welltap_svt  __well_tap__32
timestamp 1734143631
transform 1 0 72 0 1 2160
box 6 10 9 20
use welltap_svt  __well_tap__33
timestamp 1734143631
transform 1 0 4230 0 1 2160
box 6 10 9 20
use welltap_svt  __well_tap__34
timestamp 1734143631
transform 1 0 72 0 -1 2340
box 6 10 9 20
use welltap_svt  __well_tap__35
timestamp 1734143631
transform 1 0 4230 0 -1 2340
box 6 10 9 20
use welltap_svt  __well_tap__36
timestamp 1734143631
transform 1 0 72 0 1 2400
box 6 10 9 20
use welltap_svt  __well_tap__37
timestamp 1734143631
transform 1 0 4230 0 1 2400
box 6 10 9 20
use welltap_svt  __well_tap__38
timestamp 1734143631
transform 1 0 72 0 -1 2580
box 6 10 9 20
use welltap_svt  __well_tap__39
timestamp 1734143631
transform 1 0 4230 0 -1 2580
box 6 10 9 20
use welltap_svt  __well_tap__40
timestamp 1734143631
transform 1 0 72 0 1 2640
box 6 10 9 20
use welltap_svt  __well_tap__41
timestamp 1734143631
transform 1 0 4230 0 1 2640
box 6 10 9 20
use welltap_svt  __well_tap__42
timestamp 1734143631
transform 1 0 72 0 -1 2820
box 6 10 9 20
use welltap_svt  __well_tap__43
timestamp 1734143631
transform 1 0 4230 0 -1 2820
box 6 10 9 20
use welltap_svt  __well_tap__44
timestamp 1734143631
transform 1 0 72 0 1 2880
box 6 10 9 20
use welltap_svt  __well_tap__45
timestamp 1734143631
transform 1 0 4230 0 1 2880
box 6 10 9 20
use welltap_svt  __well_tap__46
timestamp 1734143631
transform 1 0 72 0 -1 3060
box 6 10 9 20
use welltap_svt  __well_tap__47
timestamp 1734143631
transform 1 0 4230 0 -1 3060
box 6 10 9 20
use welltap_svt  __well_tap__48
timestamp 1734143631
transform 1 0 72 0 1 3120
box 6 10 9 20
use welltap_svt  __well_tap__49
timestamp 1734143631
transform 1 0 4230 0 1 3120
box 6 10 9 20
use welltap_svt  __well_tap__50
timestamp 1734143631
transform 1 0 72 0 -1 3300
box 6 10 9 20
use welltap_svt  __well_tap__51
timestamp 1734143631
transform 1 0 4230 0 -1 3300
box 6 10 9 20
use welltap_svt  __well_tap__52
timestamp 1734143631
transform 1 0 72 0 1 3360
box 6 10 9 20
use welltap_svt  __well_tap__53
timestamp 1734143631
transform 1 0 4230 0 1 3360
box 6 10 9 20
use welltap_svt  __well_tap__54
timestamp 1734143631
transform 1 0 72 0 -1 3540
box 6 10 9 20
use welltap_svt  __well_tap__55
timestamp 1734143631
transform 1 0 4230 0 -1 3540
box 6 10 9 20
use welltap_svt  __well_tap__56
timestamp 1734143631
transform 1 0 72 0 1 3600
box 6 10 9 20
use welltap_svt  __well_tap__57
timestamp 1734143631
transform 1 0 4230 0 1 3600
box 6 10 9 20
use welltap_svt  __well_tap__58
timestamp 1734143631
transform 1 0 72 0 -1 3770
box 6 10 9 20
use welltap_svt  __well_tap__59
timestamp 1734143631
transform 1 0 4230 0 -1 3770
box 6 10 9 20
use welltap_svt  __well_tap__60
timestamp 1734143631
transform 1 0 72 0 1 3830
box 6 10 9 20
use welltap_svt  __well_tap__61
timestamp 1734143631
transform 1 0 4230 0 1 3830
box 6 10 9 20
use welltap_svt  __well_tap__62
timestamp 1734143631
transform 1 0 72 0 -1 4000
box 6 10 9 20
use welltap_svt  __well_tap__63
timestamp 1734143631
transform 1 0 4230 0 -1 4000
box 6 10 9 20
use welltap_svt  __well_tap__64
timestamp 1734143631
transform 1 0 72 0 1 4060
box 6 10 9 20
use welltap_svt  __well_tap__65
timestamp 1734143631
transform 1 0 4230 0 1 4060
box 6 10 9 20
use welltap_svt  __well_tap__66
timestamp 1734143631
transform 1 0 72 0 -1 4240
box 6 10 9 20
use welltap_svt  __well_tap__67
timestamp 1734143631
transform 1 0 4230 0 -1 4240
box 6 10 9 20
use welltap_svt  __well_tap__68
timestamp 1734143631
transform 1 0 72 0 1 4300
box 6 10 9 20
use welltap_svt  __well_tap__69
timestamp 1734143631
transform 1 0 4230 0 1 4300
box 6 10 9 20
use welltap_svt  __well_tap__70
timestamp 1734143631
transform 1 0 72 0 -1 4460
box 6 10 9 20
use welltap_svt  __well_tap__71
timestamp 1734143631
transform 1 0 4230 0 -1 4460
box 6 10 9 20
use _0_0std_0_0cells_0_0LATCHINV  case__split_actrl__latch_al
timestamp 1734143852
transform 1 0 1962 0 -1 2610
box 0 0 84 100
use _0_0std_0_0cells_0_0NOR2X2  case__split_actrl__latch_anx
timestamp 1734143946
transform 1 0 2130 0 -1 2610
box 0 0 48 100
use _0_0std_0_0cells_0_0LATCH  case__split_adata__latch
timestamp 1734143796
transform 1 0 1878 0 -1 3080
box 0 0 96 80
use _0_0std_0_0cells_0_0AND2X1  case__split_aelem__c_aa1
timestamp 1734143631
transform 1 0 2058 0 1 2850
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  case__split_aelem__c_aa2
timestamp 1734143631
transform 1 0 2274 0 -1 2850
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  case__split_aelem__c_aa3
timestamp 1734143631
transform 1 0 2088 0 -1 2850
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  case__split_aelem__c_aandR1
timestamp 1734143631
transform 1 0 2052 0 1 2610
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  case__split_aelem__c_aandR2
timestamp 1734143631
transform 1 0 2136 0 1 2610
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  case__split_aelem__c_ac1_acx0
timestamp 1734143631
transform 1 0 2178 0 -1 2840
box 6 10 65 70
use _0_0cell_0_0g0n_0x1  case__split_aelem__c_ac1_acx1
timestamp 1734143631
transform 1 0 2166 0 1 2870
box 6 10 21 40
use _0_0std_0_0cells_0_0INVX1  case__split_aelem__c_actrl__inv
timestamp 1734143760
transform 1 0 2070 0 -1 2600
box 0 0 30 70
use _0_0cell_0_0g0n_0x0  case__split_aelem__c_adelay_acx0
timestamp 1734143631
transform 1 0 2088 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  case__split_aelem__c_adelay_acx1
timestamp 1734143631
transform 1 0 2136 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  case__split_aelem__c_adelay_acx2
timestamp 1734143631
transform 1 0 2070 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  case__split_aelem__c_adelay_acx3
timestamp 1734143631
transform 1 0 1980 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  case__split_aelem__c_adelay_acx4
timestamp 1734143631
transform 1 0 1908 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  case__split_aelem__c_adelay_acx5
timestamp 1734143631
transform 1 0 1914 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  case__split_aelem__c_adelay_acx6
timestamp 1734143631
transform 1 0 2028 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  case__split_aelem__c_adelay_acx7
timestamp 1734143631
transform 1 0 2226 0 1 2610
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  case__split_aelem__c_ai1
timestamp 1734143760
transform 1 0 2232 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  case__split_aelem__c_an1
timestamp 1734143909
transform 1 0 1968 0 -1 2850
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  case__split_apulseG_aand
timestamp 1734143631
transform 1 0 1794 0 -1 3090
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai
timestamp 1734143760
transform 1 0 1842 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai1
timestamp 1734143760
transform 1 0 1746 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai2
timestamp 1734143760
transform 1 0 1704 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai3
timestamp 1734143760
transform 1 0 1662 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai4
timestamp 1734143760
transform 1 0 1620 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai5
timestamp 1734143760
transform 1 0 1590 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai6
timestamp 1734143760
transform 1 0 1632 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai7
timestamp 1734143760
transform 1 0 1668 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai8
timestamp 1734143760
transform 1 0 1704 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  case__split_apulseG_ai9
timestamp 1734143760
transform 1 0 1746 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  case__split_apulseG_anor
timestamp 1734143909
transform 1 0 1788 0 1 3090
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  check__caps_aand_aand
timestamp 1734143631
transform 1 0 2340 0 -1 3570
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  check__caps_aand_aelem__c_aa1
timestamp 1734143631
transform 1 0 1482 0 -1 3570
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  check__caps_aand_aelem__c_aa2
timestamp 1734143631
transform 1 0 1326 0 -1 3570
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  check__caps_aand_aelem__c_ac1_acx0
timestamp 1734143631
transform 1 0 1512 0 1 3580
box 6 10 65 70
use _0_0cell_0_0g0n_0x1  check__caps_aand_aelem__c_ac1_acx1
timestamp 1734143631
transform 1 0 1482 0 1 3820
box 6 10 21 40
use _0_0cell_0_0g0n_0x0  check__caps_aand_aelem__c_adelay_acx0
timestamp 1734143631
transform 1 0 1698 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_aand_aelem__c_adelay_acx1
timestamp 1734143631
transform 1 0 1722 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_aand_aelem__c_adelay_acx2
timestamp 1734143631
transform 1 0 1782 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_aand_aelem__c_adelay_acx3
timestamp 1734143631
transform 1 0 1794 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_aand_aelem__c_adelay_acx4
timestamp 1734143631
transform 1 0 1710 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_aand_aelem__c_adelay_acx5
timestamp 1734143631
transform 1 0 1746 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_aand_aelem__c_adelay_acx6
timestamp 1734143631
transform 1 0 1848 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_aand_aelem__c_adelay_acx7
timestamp 1734143631
transform 1 0 1854 0 1 3330
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_aelem__c_ai1
timestamp 1734143760
transform 1 0 1398 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__caps_aand_aelem__c_an1
timestamp 1734143909
transform 1 0 1728 0 1 3570
box 0 0 42 80
use _0_0std_0_0cells_0_0LATCH  check__caps_aand_alatch
timestamp 1734143796
transform 1 0 1950 0 1 3580
box 0 0 96 80
use _0_0std_0_0cells_0_0AND2X1  check__caps_aand_apulseG_aand
timestamp 1734143631
transform 1 0 1806 0 1 4030
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai1
timestamp 1734143760
transform 1 0 1674 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai2
timestamp 1734143760
transform 1 0 1686 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai3
timestamp 1734143760
transform 1 0 1728 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai4
timestamp 1734143760
transform 1 0 1776 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai5
timestamp 1734143760
transform 1 0 1818 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai6
timestamp 1734143760
transform 1 0 1866 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai7
timestamp 1734143760
transform 1 0 1842 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai8
timestamp 1734143760
transform 1 0 1788 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai9
timestamp 1734143760
transform 1 0 1776 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_aand_apulseG_ai
timestamp 1734143760
transform 1 0 1626 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__caps_aand_apulseG_anor
timestamp 1734143909
transform 1 0 1656 0 1 4030
box 0 0 42 80
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp65_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 4164 0 1 2860
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 4110 0 -1 2830
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp65_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 4050 0 1 2850
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 3984 0 1 2870
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp65_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 4068 0 -1 2600
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 4044 0 -1 2590
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp65_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 4128 0 -1 2610
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 4200 0 -1 2590
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp65_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 3996 0 1 2380
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 3852 0 1 2390
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp65_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 3966 0 -1 2370
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 3864 0 -1 2350
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp65_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 3576 0 1 2380
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 3738 0 -1 2830
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp65_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 3648 0 1 2370
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 3660 0 -1 2350
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp65_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 3750 0 1 3100
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 3414 0 1 3110
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp65_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 3762 0 -1 3090
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 3702 0 1 2870
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp65_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 3258 0 -1 3080
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 3204 0 -1 3310
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp65_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 3156 0 -1 3090
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 3192 0 1 2870
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp65_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 3066 0 -1 3080
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 3000 0 1 3110
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp65_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 2970 0 1 2850
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 2916 0 1 2870
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp65_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 2844 0 -1 3320
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 2700 0 -1 3310
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp65_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 2748 0 -1 3330
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp65_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 2742 0 1 3350
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  check__caps_acmp65_acelem_acx0
timestamp 1734143631
transform 1 0 2088 0 1 4040
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay1_acx0
timestamp 1734143631
transform 1 0 2028 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay1_acx1
timestamp 1734143631
transform 1 0 1632 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay1_acx2
timestamp 1734143631
transform 1 0 1644 0 -1 4490
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay1_acx3
timestamp 1734143631
transform 1 0 1506 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay1_acx4
timestamp 1734143631
transform 1 0 1440 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay1_acx5
timestamp 1734143631
transform 1 0 1368 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay1_acx6
timestamp 1734143631
transform 1 0 1296 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay1_acx7
timestamp 1734143631
transform 1 0 1230 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay2_acx0
timestamp 1734143631
transform 1 0 1104 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay2_acx1
timestamp 1734143631
transform 1 0 1050 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay2_acx2
timestamp 1734143631
transform 1 0 996 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay2_acx3
timestamp 1734143631
transform 1 0 978 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay2_acx4
timestamp 1734143631
transform 1 0 924 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay2_acx5
timestamp 1734143631
transform 1 0 870 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay2_acx6
timestamp 1734143631
transform 1 0 858 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay2_acx7
timestamp 1734143631
transform 1 0 792 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay3_acx0
timestamp 1734143631
transform 1 0 930 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay3_acx1
timestamp 1734143631
transform 1 0 996 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay3_acx2
timestamp 1734143631
transform 1 0 1062 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay3_acx3
timestamp 1734143631
transform 1 0 894 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay3_acx4
timestamp 1734143631
transform 1 0 966 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay3_acx5
timestamp 1734143631
transform 1 0 1170 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay3_acx6
timestamp 1734143631
transform 1 0 1242 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp65_adelay3_acx7
timestamp 1734143631
transform 1 0 1308 0 1 3800
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_ainv__l1
timestamp 1734143760
transform 1 0 2196 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_ainv__l2
timestamp 1734143760
transform 1 0 2094 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_ainv__r
timestamp 1734143760
transform 1 0 2058 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al1_50_6
timestamp 1734143796
transform 1 0 4092 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al1_51_6
timestamp 1734143796
transform 1 0 3918 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al1_52_6
timestamp 1734143796
transform 1 0 3948 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al1_53_6
timestamp 1734143796
transform 1 0 3234 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al1_54_6
timestamp 1734143796
transform 1 0 3462 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al1_55_6
timestamp 1734143796
transform 1 0 3246 0 1 2860
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al1_56_6
timestamp 1734143796
transform 1 0 2946 0 -1 3080
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al1_57_6
timestamp 1734143796
transform 1 0 2886 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al2_50_6
timestamp 1734143796
transform 1 0 4038 0 -1 3080
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al2_51_6
timestamp 1734143796
transform 1 0 4026 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al2_52_6
timestamp 1734143796
transform 1 0 3888 0 1 2380
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al2_53_6
timestamp 1734143796
transform 1 0 3330 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al2_54_6
timestamp 1734143796
transform 1 0 3636 0 -1 3320
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al2_55_6
timestamp 1734143796
transform 1 0 3228 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al2_56_6
timestamp 1734143796
transform 1 0 3102 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp65_al2_57_6
timestamp 1734143796
transform 1 0 2982 0 -1 3320
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  check__caps_acmp65_anor
timestamp 1734143909
transform 1 0 1968 0 -1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  check__caps_acmp65_aor__l1
timestamp 1734143975
transform 1 0 2226 0 1 4040
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  check__caps_acmp65_aor__l2
timestamp 1734143975
transform 1 0 2076 0 -1 4260
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  check__caps_acmp65_apulseG_aand
timestamp 1734143631
transform 1 0 2880 0 -1 4270
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai1
timestamp 1734143760
transform 1 0 2802 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai2
timestamp 1734143760
transform 1 0 2760 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai3
timestamp 1734143760
transform 1 0 2742 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai4
timestamp 1734143760
transform 1 0 2898 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai5
timestamp 1734143760
transform 1 0 3078 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai6
timestamp 1734143760
transform 1 0 2994 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai7
timestamp 1734143760
transform 1 0 2892 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai8
timestamp 1734143760
transform 1 0 2940 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai9
timestamp 1734143760
transform 1 0 2958 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp65_apulseG_ai
timestamp 1734143760
transform 1 0 2514 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__caps_acmp65_apulseG_anor
timestamp 1734143909
transform 1 0 2568 0 -1 4270
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  check__caps_acmp65_atoGND
timestamp 1734144021
transform 1 0 4170 0 -1 3070
box 0 0 30 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp91_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 4014 0 1 3100
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 3984 0 -1 3070
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp91_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 3930 0 1 3090
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 3870 0 -1 3070
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp91_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 4014 0 -1 2840
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 3858 0 1 2630
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp91_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 3912 0 -1 2850
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 3888 0 1 2630
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp91_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 3678 0 -1 2600
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 3558 0 -1 2590
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp91_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 3738 0 -1 2610
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 3816 0 1 2390
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp91_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 3498 0 -1 2600
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 3474 0 -1 2830
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp91_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 3426 0 -1 2610
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 3456 0 1 2390
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp91_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 3594 0 1 2860
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 3522 0 1 2870
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp91_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 3522 0 -1 2850
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 3420 0 -1 2830
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp91_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 3108 0 -1 2840
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 3048 0 1 3110
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp91_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 3120 0 1 2610
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 3078 0 1 2630
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp91_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 2766 0 -1 3080
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 2928 0 -1 3310
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp91_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 2850 0 -1 3090
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 2856 0 1 2870
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__caps_acmp91_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 2940 0 -1 3560
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 3042 0 -1 3550
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__caps_acmp91_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 2826 0 -1 3570
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__caps_acmp91_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 2484 0 -1 3550
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  check__caps_acmp91_acelem_acx0
timestamp 1734143631
transform 1 0 1950 0 1 4040
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay1_acx0
timestamp 1734143631
transform 1 0 1728 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay1_acx1
timestamp 1734143631
transform 1 0 1590 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay1_acx2
timestamp 1734143631
transform 1 0 1500 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay1_acx3
timestamp 1734143631
transform 1 0 1284 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay1_acx4
timestamp 1734143631
transform 1 0 1230 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay1_acx5
timestamp 1734143631
transform 1 0 1182 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay1_acx6
timestamp 1734143631
transform 1 0 942 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay1_acx7
timestamp 1734143631
transform 1 0 894 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay2_acx0
timestamp 1734143631
transform 1 0 900 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay2_acx1
timestamp 1734143631
transform 1 0 828 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay2_acx2
timestamp 1734143631
transform 1 0 756 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay2_acx3
timestamp 1734143631
transform 1 0 840 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay2_acx4
timestamp 1734143631
transform 1 0 768 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay2_acx5
timestamp 1734143631
transform 1 0 696 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay2_acx6
timestamp 1734143631
transform 1 0 618 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay2_acx7
timestamp 1734143631
transform 1 0 690 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay3_acx0
timestamp 1734143631
transform 1 0 750 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay3_acx1
timestamp 1734143631
transform 1 0 774 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay3_acx2
timestamp 1734143631
transform 1 0 828 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay3_acx3
timestamp 1734143631
transform 1 0 888 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay3_acx4
timestamp 1734143631
transform 1 0 954 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay3_acx5
timestamp 1734143631
transform 1 0 1080 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay3_acx6
timestamp 1734143631
transform 1 0 1080 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acmp91_adelay3_acx7
timestamp 1734143631
transform 1 0 1146 0 1 3330
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_ainv__l1
timestamp 1734143760
transform 1 0 2028 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_ainv__l2
timestamp 1734143760
transform 1 0 1968 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_ainv__r
timestamp 1734143760
transform 1 0 1866 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al1_50_6
timestamp 1734143796
transform 1 0 3822 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al1_51_6
timestamp 1734143796
transform 1 0 3786 0 -1 2840
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al1_52_6
timestamp 1734143796
transform 1 0 3582 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al1_53_6
timestamp 1734143796
transform 1 0 3420 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al1_54_6
timestamp 1734143796
transform 1 0 3492 0 -1 3080
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al1_55_6
timestamp 1734143796
transform 1 0 3066 0 1 2860
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al1_56_6
timestamp 1734143796
transform 1 0 2886 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al1_57_6
timestamp 1734143796
transform 1 0 2778 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al2_50_6
timestamp 1734143796
transform 1 0 3798 0 -1 3320
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al2_51_6
timestamp 1734143796
transform 1 0 3774 0 1 2860
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al2_52_6
timestamp 1734143796
transform 1 0 3810 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al2_53_6
timestamp 1734143796
transform 1 0 3720 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al2_54_6
timestamp 1734143796
transform 1 0 3630 0 -1 3080
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al2_55_6
timestamp 1734143796
transform 1 0 3216 0 -1 2840
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al2_56_6
timestamp 1734143796
transform 1 0 2772 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acmp91_al2_57_6
timestamp 1734143796
transform 1 0 2898 0 1 3580
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  check__caps_acmp91_anor
timestamp 1734143909
transform 1 0 1734 0 1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  check__caps_acmp91_aor__l1
timestamp 1734143975
transform 1 0 1896 0 1 4040
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  check__caps_acmp91_aor__l2
timestamp 1734143975
transform 1 0 1896 0 -1 4260
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  check__caps_acmp91_apulseG_aand
timestamp 1734143631
transform 1 0 2754 0 -1 4030
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai1
timestamp 1734143760
transform 1 0 2664 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai2
timestamp 1734143760
transform 1 0 2628 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai3
timestamp 1734143760
transform 1 0 2682 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai4
timestamp 1734143760
transform 1 0 2736 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai5
timestamp 1734143760
transform 1 0 2784 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai6
timestamp 1734143760
transform 1 0 2832 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai7
timestamp 1734143760
transform 1 0 2862 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai8
timestamp 1734143760
transform 1 0 2808 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai9
timestamp 1734143760
transform 1 0 2760 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acmp91_apulseG_ai
timestamp 1734143760
transform 1 0 2412 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__caps_acmp91_apulseG_anor
timestamp 1734143909
transform 1 0 2604 0 1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  check__caps_acmp91_atoGND
timestamp 1734144021
transform 1 0 4056 0 -1 3310
box 0 0 30 50
use _0_0cell_0_0g0n1n2naa_012aax0  check__caps_acp_acelem_acx0
timestamp 1734143631
transform 1 0 2616 0 -1 4020
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  check__caps_acp_adelay1_acx0
timestamp 1734143631
transform 1 0 2496 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acp_adelay1_acx1
timestamp 1734143631
transform 1 0 2448 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acp_adelay1_acx2
timestamp 1734143631
transform 1 0 2454 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acp_adelay1_acx3
timestamp 1734143631
transform 1 0 2388 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acp_adelay1_acx4
timestamp 1734143631
transform 1 0 2262 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acp_adelay1_acx5
timestamp 1734143631
transform 1 0 2202 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acp_adelay1_acx6
timestamp 1734143631
transform 1 0 2148 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_acp_adelay1_acx7
timestamp 1734143631
transform 1 0 2160 0 1 4030
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_ainv__1
timestamp 1734143760
transform 1 0 2574 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_ainv__2
timestamp 1734143760
transform 1 0 2466 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_ainv__3
timestamp 1734143760
transform 1 0 2454 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  check__caps_acp_al_50_6
timestamp 1734143796
transform 1 0 3582 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acp_al_51_6
timestamp 1734143796
transform 1 0 3618 0 -1 2840
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acp_al_52_6
timestamp 1734143796
transform 1 0 3618 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acp_al_53_6
timestamp 1734143796
transform 1 0 3516 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acp_al_54_6
timestamp 1734143796
transform 1 0 3354 0 -1 3080
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acp_al_55_6
timestamp 1734143796
transform 1 0 3378 0 1 2860
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acp_al_56_6
timestamp 1734143796
transform 1 0 3288 0 -1 3320
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__caps_acp_al_57_6
timestamp 1734143796
transform 1 0 2988 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  check__caps_acp_anor__2
timestamp 1734143909
transform 1 0 2544 0 1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  check__caps_acp_anor__3
timestamp 1734143909
transform 1 0 2364 0 1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  check__caps_acp_aor__1
timestamp 1734143975
transform 1 0 2508 0 -1 4020
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  check__caps_acp_apulseG_aand
timestamp 1734143631
transform 1 0 3126 0 -1 4030
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai1
timestamp 1734143760
transform 1 0 2982 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai2
timestamp 1734143760
transform 1 0 3006 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai3
timestamp 1734143760
transform 1 0 3048 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai4
timestamp 1734143760
transform 1 0 3084 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai5
timestamp 1734143760
transform 1 0 3120 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai6
timestamp 1734143760
transform 1 0 3156 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai7
timestamp 1734143760
transform 1 0 3192 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai8
timestamp 1734143760
transform 1 0 3156 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai
timestamp 1734143760
transform 1 0 2712 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_acp_apulseG_ai9
timestamp 1734143760
transform 1 0 3192 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__caps_acp_apulseG_anor
timestamp 1734143909
transform 1 0 2916 0 1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  check__caps_ainv_aelem__c_aa1
timestamp 1734143631
transform 1 0 1380 0 1 3800
box 0 0 60 80
use _0_0cell_0_0g0n1na_01ax0  check__caps_ainv_aelem__c_ac1_acx0
timestamp 1734143631
transform 1 0 1500 0 -1 4020
box 6 10 63 60
use _0_0cell_0_0g0n_0x1  check__caps_ainv_aelem__c_ac1_acx1
timestamp 1734143631
transform 1 0 1572 0 -1 4010
box 6 10 21 40
use _0_0cell_0_0g0n_0x0  check__caps_ainv_aelem__c_adelay_acx0
timestamp 1734143631
transform 1 0 1662 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_ainv_aelem__c_adelay_acx1
timestamp 1734143631
transform 1 0 1608 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_ainv_aelem__c_adelay_acx2
timestamp 1734143631
transform 1 0 1626 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_ainv_aelem__c_adelay_acx3
timestamp 1734143631
transform 1 0 1548 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_ainv_aelem__c_adelay_acx4
timestamp 1734143631
transform 1 0 1548 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_ainv_aelem__c_adelay_acx5
timestamp 1734143631
transform 1 0 1470 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_ainv_aelem__c_adelay_acx6
timestamp 1734143631
transform 1 0 1434 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__caps_ainv_aelem__c_adelay_acx7
timestamp 1734143631
transform 1 0 1440 0 -1 3570
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_aelem__c_ai1
timestamp 1734143760
transform 1 0 1338 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__caps_ainv_aelem__c_an1
timestamp 1734143909
transform 1 0 1458 0 -1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_ain
timestamp 1734143760
transform 1 0 2430 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  check__caps_ainv_alatch
timestamp 1734143796
transform 1 0 2292 0 1 3580
box 0 0 96 80
use _0_0std_0_0cells_0_0AND2X1  check__caps_ainv_apulseG_aand
timestamp 1734143631
transform 1 0 2226 0 1 3570
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai1
timestamp 1734143760
transform 1 0 2118 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai2
timestamp 1734143760
transform 1 0 2172 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai3
timestamp 1734143760
transform 1 0 2226 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai
timestamp 1734143760
transform 1 0 2010 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai4
timestamp 1734143760
transform 1 0 2190 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai5
timestamp 1734143760
transform 1 0 2154 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai6
timestamp 1734143760
transform 1 0 2112 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai7
timestamp 1734143760
transform 1 0 2154 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai8
timestamp 1734143760
transform 1 0 2220 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__caps_ainv_apulseG_ai9
timestamp 1734143760
transform 1 0 2280 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__caps_ainv_apulseG_anor
timestamp 1734143909
transform 1 0 2058 0 -1 3800
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  check__caps_asrcNeg65_anor
timestamp 1734143909
transform 1 0 2154 0 1 4270
box 0 0 42 80
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg65_aset0
timestamp 1734144001
transform 1 0 3924 0 -1 3070
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg65_aset1
timestamp 1734144001
transform 1 0 4134 0 1 2630
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg65_aset2
timestamp 1734144001
transform 1 0 4068 0 1 2390
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg65_aset3
timestamp 1734144001
transform 1 0 3732 0 1 2390
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg65_aset4
timestamp 1734144001
transform 1 0 3546 0 -1 3310
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg65_aset5
timestamp 1734144001
transform 1 0 3354 0 1 3110
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__caps_asrcNeg65_aset6
timestamp 1734144021
transform 1 0 3450 0 -1 3310
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg65_aset7
timestamp 1734144001
transform 1 0 3120 0 -1 3310
box 0 0 30 50
use _0_0std_0_0cells_0_0NOR2X1  check__caps_asrcNeg91_anor
timestamp 1734143909
transform 1 0 2016 0 -1 4270
box 0 0 42 80
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg91_asetGND0
timestamp 1734144001
transform 1 0 3960 0 -1 3310
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__caps_asrcNeg91_asetGND1
timestamp 1734144021
transform 1 0 3912 0 1 2870
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg91_asetGND2
timestamp 1734144001
transform 1 0 3912 0 -1 2590
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__caps_asrcNeg91_asetGND3
timestamp 1734144021
transform 1 0 3822 0 1 2630
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__caps_asrcNeg91_asetGND4
timestamp 1734144021
transform 1 0 3702 0 1 3110
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg91_asetGND5
timestamp 1734144001
transform 1 0 3354 0 -1 2830
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__caps_asrcNeg91_asetGND6
timestamp 1734144021
transform 1 0 2652 0 1 3110
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__caps_asrcNeg91_asetGND7
timestamp 1734144001
transform 1 0 3030 0 1 3590
box 0 0 30 50
use _0_0std_0_0cells_0_0AND2X1  check__lower_aand_aand
timestamp 1734143631
transform 1 0 2280 0 -1 3800
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  check__lower_aand_aelem__c_aa1
timestamp 1734143631
transform 1 0 1008 0 -1 3570
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  check__lower_aand_aelem__c_aa2
timestamp 1734143631
transform 1 0 804 0 -1 3570
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  check__lower_aand_aelem__c_ac1_acx0
timestamp 1734143631
transform 1 0 1080 0 -1 3560
box 6 10 65 70
use _0_0cell_0_0g0n_0x1  check__lower_aand_aelem__c_ac1_acx1
timestamp 1734143631
transform 1 0 1050 0 1 3590
box 6 10 21 40
use _0_0cell_0_0g0n_0x0  check__lower_aand_aelem__c_adelay_acx0
timestamp 1734143631
transform 1 0 1098 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_aand_aelem__c_adelay_acx1
timestamp 1734143631
transform 1 0 1098 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_aand_aelem__c_adelay_acx2
timestamp 1734143631
transform 1 0 1152 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_aand_aelem__c_adelay_acx3
timestamp 1734143631
transform 1 0 1170 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_aand_aelem__c_adelay_acx4
timestamp 1734143631
transform 1 0 1224 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_aand_aelem__c_adelay_acx5
timestamp 1734143631
transform 1 0 1212 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_aand_aelem__c_adelay_acx6
timestamp 1734143631
transform 1 0 1272 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_aand_aelem__c_adelay_acx7
timestamp 1734143631
transform 1 0 1332 0 1 3330
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_aelem__c_ai1
timestamp 1734143760
transform 1 0 876 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__lower_aand_aelem__c_an1
timestamp 1734143909
transform 1 0 1272 0 -1 3570
box 0 0 42 80
use _0_0std_0_0cells_0_0LATCH  check__lower_aand_alatch
timestamp 1734143796
transform 1 0 1620 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0AND2X1  check__lower_aand_apulseG_aand
timestamp 1734143631
transform 1 0 1374 0 1 3570
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai1
timestamp 1734143760
transform 1 0 1410 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai2
timestamp 1734143760
transform 1 0 1482 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai3
timestamp 1734143760
transform 1 0 1338 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai4
timestamp 1734143760
transform 1 0 1272 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai
timestamp 1734143760
transform 1 0 1152 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai5
timestamp 1734143760
transform 1 0 1206 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai6
timestamp 1734143760
transform 1 0 1248 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai7
timestamp 1734143760
transform 1 0 1284 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai8
timestamp 1734143760
transform 1 0 1314 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_aand_apulseG_ai9
timestamp 1734143760
transform 1 0 1344 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__lower_aand_apulseG_anor
timestamp 1734143909
transform 1 0 1200 0 -1 3800
box 0 0 42 80
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp97_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 4044 0 -1 4020
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 4140 0 1 3820
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp97_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 4116 0 -1 4030
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 4200 0 -1 4010
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp97_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 4068 0 -1 3790
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 4038 0 -1 3780
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp97_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 4104 0 1 3570
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 4068 0 1 3590
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp97_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 3918 0 1 3580
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 3768 0 -1 4010
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp97_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 3984 0 1 3570
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 4014 0 -1 3550
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp97_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 3660 0 1 4040
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 3672 0 -1 4250
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp97_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 3678 0 -1 4030
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 3630 0 -1 4010
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp97_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 3528 0 -1 4260
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 3498 0 -1 4250
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp97_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 3594 0 -1 4270
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 3594 0 1 4050
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp97_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 3432 0 -1 4260
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 3384 0 1 4050
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp97_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 3432 0 1 4030
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 3534 0 1 4050
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp97_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 3276 0 -1 4020
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 3234 0 -1 4010
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp97_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 3360 0 -1 4030
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 3462 0 -1 4010
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp97_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 3030 0 -1 4020
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 3000 0 -1 4010
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp97_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 2922 0 -1 4030
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp97_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 2790 0 1 3820
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  check__lower_acmp97_acelem_acx0
timestamp 1734143631
transform 1 0 1428 0 1 4040
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay1_acx0
timestamp 1734143631
transform 1 0 1284 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay1_acx1
timestamp 1734143631
transform 1 0 1134 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay1_acx2
timestamp 1734143631
transform 1 0 948 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay1_acx3
timestamp 1734143631
transform 1 0 894 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay1_acx4
timestamp 1734143631
transform 1 0 840 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay1_acx5
timestamp 1734143631
transform 1 0 786 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay1_acx6
timestamp 1734143631
transform 1 0 732 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay1_acx7
timestamp 1734143631
transform 1 0 684 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay2_acx0
timestamp 1734143631
transform 1 0 642 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay2_acx1
timestamp 1734143631
transform 1 0 606 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay2_acx2
timestamp 1734143631
transform 1 0 570 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay2_acx3
timestamp 1734143631
transform 1 0 534 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay2_acx4
timestamp 1734143631
transform 1 0 624 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay2_acx5
timestamp 1734143631
transform 1 0 558 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay2_acx6
timestamp 1734143631
transform 1 0 492 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay2_acx7
timestamp 1734143631
transform 1 0 426 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay3_acx0
timestamp 1734143631
transform 1 0 462 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay3_acx1
timestamp 1734143631
transform 1 0 534 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay3_acx2
timestamp 1734143631
transform 1 0 504 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay3_acx3
timestamp 1734143631
transform 1 0 552 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay3_acx4
timestamp 1734143631
transform 1 0 606 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay3_acx5
timestamp 1734143631
transform 1 0 666 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay3_acx6
timestamp 1734143631
transform 1 0 720 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp97_adelay3_acx7
timestamp 1734143631
transform 1 0 684 0 -1 3800
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_ainv__l1
timestamp 1734143760
transform 1 0 1548 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_ainv__l2
timestamp 1734143760
transform 1 0 1326 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_ainv__r
timestamp 1734143760
transform 1 0 1428 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al1_50_6
timestamp 1734143796
transform 1 0 3936 0 -1 4020
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al1_51_6
timestamp 1734143796
transform 1 0 3930 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al1_52_6
timestamp 1734143796
transform 1 0 3810 0 1 3580
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al1_53_6
timestamp 1734143796
transform 1 0 3696 0 1 3810
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al1_54_6
timestamp 1734143796
transform 1 0 3510 0 -1 4020
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al1_55_6
timestamp 1734143796
transform 1 0 3294 0 1 3810
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al1_56_6
timestamp 1734143796
transform 1 0 3150 0 1 3810
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al1_57_6
timestamp 1734143796
transform 1 0 2820 0 -1 4020
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al2_50_6
timestamp 1734143796
transform 1 0 4086 0 1 4040
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al2_51_6
timestamp 1734143796
transform 1 0 4128 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al2_52_6
timestamp 1734143796
transform 1 0 3774 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al2_53_6
timestamp 1734143796
transform 1 0 3762 0 1 4040
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al2_54_6
timestamp 1734143796
transform 1 0 3552 0 1 4280
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al2_55_6
timestamp 1734143796
transform 1 0 3330 0 -1 4260
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al2_56_6
timestamp 1734143796
transform 1 0 3210 0 1 4040
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp97_al2_57_6
timestamp 1734143796
transform 1 0 3036 0 1 4040
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  check__lower_acmp97_anor
timestamp 1734143909
transform 1 0 1380 0 -1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  check__lower_acmp97_aor__l1
timestamp 1734143975
transform 1 0 1536 0 1 4040
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  check__lower_acmp97_aor__l2
timestamp 1734143975
transform 1 0 1368 0 1 4040
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  check__lower_acmp97_apulseG_aand
timestamp 1734143631
transform 1 0 2748 0 -1 3800
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai
timestamp 1734143760
transform 1 0 2262 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai1
timestamp 1734143760
transform 1 0 2640 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai2
timestamp 1734143760
transform 1 0 2586 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai3
timestamp 1734143760
transform 1 0 2538 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai4
timestamp 1734143760
transform 1 0 2478 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai5
timestamp 1734143760
transform 1 0 2526 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai6
timestamp 1734143760
transform 1 0 2568 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai7
timestamp 1734143760
transform 1 0 2610 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai8
timestamp 1734143760
transform 1 0 2652 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp97_apulseG_ai9
timestamp 1734143760
transform 1 0 2700 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__lower_acmp97_apulseG_anor
timestamp 1734143909
transform 1 0 2358 0 1 3800
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  check__lower_acmp97_atoGND
timestamp 1734144021
transform 1 0 4008 0 1 4050
box 0 0 30 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp123_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 4008 0 1 4280
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 3978 0 -1 4250
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp123_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 4014 0 -1 4270
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 4104 0 -1 4250
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp123_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 3900 0 1 4040
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 3864 0 1 3820
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp123_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 3852 0 -1 4030
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 3810 0 -1 4010
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp123_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 3822 0 -1 3560
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 3774 0 1 3590
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp123_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 3840 0 1 3330
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 3918 0 1 3350
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp123_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 3702 0 1 3580
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 3570 0 -1 3780
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp123_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 3618 0 1 3570
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 3552 0 -1 3550
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp123_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 3372 0 -1 3790
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 3300 0 1 3590
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp123_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 3384 0 1 3570
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 3342 0 1 3590
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp123_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 3342 0 -1 3560
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 3252 0 1 3590
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp123_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 3234 0 -1 3570
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 3198 0 1 3350
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp123_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 3174 0 -1 3790
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 3018 0 -1 3780
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp123_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 3150 0 1 3570
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 3096 0 1 3590
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  check__lower_acmp123_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 2826 0 -1 3790
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 2640 0 1 3590
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  check__lower_acmp123_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 2796 0 1 3570
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  check__lower_acmp123_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 2598 0 1 3590
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  check__lower_acmp123_acelem_acx0
timestamp 1734143631
transform 1 0 1182 0 1 4040
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay1_acx0
timestamp 1734143631
transform 1 0 1164 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay1_acx1
timestamp 1734143631
transform 1 0 1086 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay1_acx2
timestamp 1734143631
transform 1 0 1032 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay1_acx3
timestamp 1734143631
transform 1 0 810 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay1_acx4
timestamp 1734143631
transform 1 0 750 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay1_acx5
timestamp 1734143631
transform 1 0 690 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay1_acx6
timestamp 1734143631
transform 1 0 666 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay1_acx7
timestamp 1734143631
transform 1 0 600 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay2_acx0
timestamp 1734143631
transform 1 0 726 0 1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay2_acx1
timestamp 1734143631
transform 1 0 822 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay2_acx2
timestamp 1734143631
transform 1 0 744 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay2_acx3
timestamp 1734143631
transform 1 0 672 0 -1 4030
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay2_acx4
timestamp 1734143631
transform 1 0 612 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay2_acx5
timestamp 1734143631
transform 1 0 564 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay2_acx6
timestamp 1734143631
transform 1 0 522 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay2_acx7
timestamp 1734143631
transform 1 0 462 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay3_acx0
timestamp 1734143631
transform 1 0 534 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay3_acx1
timestamp 1734143631
transform 1 0 606 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay3_acx2
timestamp 1734143631
transform 1 0 540 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay3_acx3
timestamp 1734143631
transform 1 0 462 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay3_acx4
timestamp 1734143631
transform 1 0 498 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay3_acx5
timestamp 1734143631
transform 1 0 564 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay3_acx6
timestamp 1734143631
transform 1 0 630 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acmp123_adelay3_acx7
timestamp 1734143631
transform 1 0 720 0 1 3330
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_ainv__l1
timestamp 1734143760
transform 1 0 1488 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_ainv__l2
timestamp 1734143760
transform 1 0 1242 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_ainv__r
timestamp 1734143760
transform 1 0 1128 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al1_50_6
timestamp 1734143796
transform 1 0 3876 0 -1 4260
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al1_51_6
timestamp 1734143796
transform 1 0 3966 0 1 3810
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al1_52_6
timestamp 1734143796
transform 1 0 3708 0 -1 3560
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al1_53_6
timestamp 1734143796
transform 1 0 3510 0 1 3580
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al1_54_6
timestamp 1734143796
transform 1 0 3456 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al1_55_6
timestamp 1734143796
transform 1 0 3102 0 -1 3560
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al1_56_6
timestamp 1734143796
transform 1 0 3252 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al1_57_6
timestamp 1734143796
transform 1 0 2904 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al2_50_6
timestamp 1734143796
transform 1 0 3858 0 1 4280
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al2_51_6
timestamp 1734143796
transform 1 0 3702 0 -1 4260
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al2_52_6
timestamp 1734143796
transform 1 0 3900 0 -1 3560
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al2_53_6
timestamp 1734143796
transform 1 0 3612 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al2_54_6
timestamp 1734143796
transform 1 0 3444 0 1 3810
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al2_55_6
timestamp 1734143796
transform 1 0 3432 0 -1 3560
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al2_56_6
timestamp 1734143796
transform 1 0 3060 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acmp123_al2_57_6
timestamp 1734143796
transform 1 0 2862 0 1 3810
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  check__lower_acmp123_anor
timestamp 1734143909
transform 1 0 1098 0 -1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  check__lower_acmp123_aor__l1
timestamp 1734143975
transform 1 0 1404 0 -1 4260
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  check__lower_acmp123_aor__l2
timestamp 1734143975
transform 1 0 1182 0 -1 4260
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  check__lower_acmp123_apulseG_aand
timestamp 1734143631
transform 1 0 2694 0 1 4270
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai1
timestamp 1734143760
transform 1 0 2430 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai2
timestamp 1734143760
transform 1 0 2088 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai3
timestamp 1734143760
transform 1 0 2274 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai4
timestamp 1734143760
transform 1 0 2442 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai5
timestamp 1734143760
transform 1 0 2592 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai6
timestamp 1734143760
transform 1 0 2544 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai7
timestamp 1734143760
transform 1 0 2586 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai8
timestamp 1734143760
transform 1 0 2622 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai9
timestamp 1734143760
transform 1 0 2658 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acmp123_apulseG_ai
timestamp 1734143760
transform 1 0 2370 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__lower_acmp123_apulseG_anor
timestamp 1734143909
transform 1 0 2484 0 1 4270
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  check__lower_acmp123_atoGND
timestamp 1734144021
transform 1 0 4002 0 -1 4470
box 0 0 30 50
use _0_0cell_0_0g0n1n2naa_012aax0  check__lower_acp_acelem_acx0
timestamp 1734143631
transform 1 0 2328 0 -1 4020
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  check__lower_acp_adelay1_acx0
timestamp 1734143631
transform 1 0 2322 0 -1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acp_adelay1_acx1
timestamp 1734143631
transform 1 0 2304 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acp_adelay1_acx2
timestamp 1734143631
transform 1 0 2232 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acp_adelay1_acx3
timestamp 1734143631
transform 1 0 1878 0 -1 4490
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acp_adelay1_acx4
timestamp 1734143631
transform 1 0 1968 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acp_adelay1_acx5
timestamp 1734143631
transform 1 0 1914 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acp_adelay1_acx6
timestamp 1734143631
transform 1 0 1572 0 1 4270
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_acp_adelay1_acx7
timestamp 1734143631
transform 1 0 1608 0 -1 4270
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_ainv__1
timestamp 1734143760
transform 1 0 2292 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_ainv__2
timestamp 1734143760
transform 1 0 2328 0 1 4040
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_ainv__3
timestamp 1734143760
transform 1 0 2412 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  check__lower_acp_al_50_6
timestamp 1734143796
transform 1 0 3594 0 -1 3560
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acp_al_51_6
timestamp 1734143796
transform 1 0 3738 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acp_al_52_6
timestamp 1734143796
transform 1 0 3636 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acp_al_53_6
timestamp 1734143796
transform 1 0 3534 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acp_al_54_6
timestamp 1734143796
transform 1 0 3432 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acp_al_55_6
timestamp 1734143796
transform 1 0 3330 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acp_al_56_6
timestamp 1734143796
transform 1 0 3228 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  check__lower_acp_al_57_6
timestamp 1734143796
transform 1 0 3096 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  check__lower_acp_anor__2
timestamp 1734143909
transform 1 0 2220 0 -1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  check__lower_acp_anor__3
timestamp 1734143909
transform 1 0 2280 0 1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  check__lower_acp_aor__1
timestamp 1734143975
transform 1 0 2406 0 -1 4020
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  check__lower_acp_apulseG_aand
timestamp 1734143631
transform 1 0 3264 0 -1 4270
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai1
timestamp 1734143760
transform 1 0 3120 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai2
timestamp 1734143760
transform 1 0 3180 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai3
timestamp 1734143760
transform 1 0 3288 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai4
timestamp 1734143760
transform 1 0 3516 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai5
timestamp 1734143760
transform 1 0 3756 0 -1 4480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai6
timestamp 1734143760
transform 1 0 3474 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai7
timestamp 1734143760
transform 1 0 3318 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai8
timestamp 1734143760
transform 1 0 3246 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai
timestamp 1734143760
transform 1 0 2844 0 1 4280
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_acp_apulseG_ai9
timestamp 1734143760
transform 1 0 3228 0 -1 4260
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__lower_acp_apulseG_anor
timestamp 1734143909
transform 1 0 3048 0 1 4270
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  check__lower_ainv_aelem__c_aa1
timestamp 1734143631
transform 1 0 822 0 1 3800
box 0 0 60 80
use _0_0cell_0_0g0n1na_01ax0  check__lower_ainv_aelem__c_ac1_acx0
timestamp 1734143631
transform 1 0 990 0 1 3810
box 6 10 63 60
use _0_0cell_0_0g0n_0x1  check__lower_ainv_aelem__c_ac1_acx1
timestamp 1734143631
transform 1 0 1038 0 -1 4010
box 6 10 21 40
use _0_0cell_0_0g0n_0x0  check__lower_ainv_aelem__c_adelay_acx0
timestamp 1734143631
transform 1 0 1068 0 1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_ainv_aelem__c_adelay_acx1
timestamp 1734143631
transform 1 0 1038 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_ainv_aelem__c_adelay_acx2
timestamp 1734143631
transform 1 0 972 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_ainv_aelem__c_adelay_acx3
timestamp 1734143631
transform 1 0 984 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_ainv_aelem__c_adelay_acx4
timestamp 1734143631
transform 1 0 912 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_ainv_aelem__c_adelay_acx5
timestamp 1734143631
transform 1 0 912 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_ainv_aelem__c_adelay_acx6
timestamp 1734143631
transform 1 0 960 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  check__lower_ainv_aelem__c_adelay_acx7
timestamp 1734143631
transform 1 0 1014 0 1 3330
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_aelem__c_ai1
timestamp 1734143760
transform 1 0 774 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__lower_ainv_aelem__c_an1
timestamp 1734143909
transform 1 0 1122 0 1 3800
box 0 0 42 80
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_ain
timestamp 1734143760
transform 1 0 2496 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  check__lower_ainv_alatch
timestamp 1734143796
transform 1 0 2364 0 -1 3790
box 0 0 96 80
use _0_0std_0_0cells_0_0AND2X1  check__lower_ainv_apulseG_aand
timestamp 1734143631
transform 1 0 2070 0 1 3800
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai1
timestamp 1734143760
transform 1 0 2034 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai2
timestamp 1734143760
transform 1 0 2082 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai3
timestamp 1734143760
transform 1 0 2124 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai4
timestamp 1734143760
transform 1 0 2160 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai5
timestamp 1734143760
transform 1 0 2190 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai
timestamp 1734143760
transform 1 0 1848 0 -1 4020
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai6
timestamp 1734143760
transform 1 0 2208 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai7
timestamp 1734143760
transform 1 0 2262 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai8
timestamp 1734143760
transform 1 0 2310 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  check__lower_ainv_apulseG_ai9
timestamp 1734143760
transform 1 0 2154 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  check__lower_ainv_apulseG_anor
timestamp 1734143909
transform 1 0 1902 0 -1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  check__lower_asrcNeg97_anor
timestamp 1734143909
transform 1 0 1272 0 1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg97_asetGND0
timestamp 1734144001
transform 1 0 4152 0 -1 4250
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg97_asetGND1
timestamp 1734144001
transform 1 0 4188 0 1 3590
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg97_asetGND2
timestamp 1734144001
transform 1 0 3888 0 -1 3780
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg97_asetGND3
timestamp 1734144001
transform 1 0 3840 0 -1 4250
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg97_asetGND4
timestamp 1734144001
transform 1 0 3696 0 1 4290
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__lower_asrcNeg97_asetGND5
timestamp 1734144021
transform 1 0 3396 0 1 4290
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__lower_asrcNeg97_asetGND6
timestamp 1734144021
transform 1 0 3330 0 1 4050
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg97_asetGND7
timestamp 1734144001
transform 1 0 3090 0 -1 4010
box 0 0 30 50
use _0_0std_0_0cells_0_0NOR2X1  check__lower_asrcNeg123_anor
timestamp 1734143909
transform 1 0 1338 0 -1 4270
box 0 0 42 80
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg123_asetGND0
timestamp 1734144001
transform 1 0 3774 0 1 4290
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__lower_asrcNeg123_asetGND1
timestamp 1734144021
transform 1 0 3804 0 -1 4250
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg123_asetGND2
timestamp 1734144001
transform 1 0 3954 0 1 3350
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__lower_asrcNeg123_asetGND3
timestamp 1734144021
transform 1 0 3726 0 -1 3780
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__lower_asrcNeg123_asetGND4
timestamp 1734144021
transform 1 0 3600 0 1 3820
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__lower_asrcNeg123_asetGND5
timestamp 1734144021
transform 1 0 3468 0 1 3590
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  check__lower_asrcNeg123_asetGND6
timestamp 1734144021
transform 1 0 3078 0 1 3820
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  check__lower_asrcNeg123_asetGND7
timestamp 1734144001
transform 1 0 3006 0 1 3820
box 0 0 30 50
use _0_0cell_0_0g0n1n2naa_012aax0  copy__ctrl__shift__splits_acelem_acx0
timestamp 1734143631
transform 1 0 2532 0 1 2860
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift__splits_adelay1_acx0
timestamp 1734143631
transform 1 0 2388 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift__splits_adelay1_acx1
timestamp 1734143631
transform 1 0 2460 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift__splits_adelay1_acx2
timestamp 1734143631
transform 1 0 2466 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift__splits_adelay1_acx3
timestamp 1734143631
transform 1 0 2520 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift__splits_adelay1_acx4
timestamp 1734143631
transform 1 0 2496 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift__splits_adelay1_acx5
timestamp 1734143631
transform 1 0 2430 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift__splits_adelay1_acx6
timestamp 1734143631
transform 1 0 2364 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift__splits_adelay1_acx7
timestamp 1734143631
transform 1 0 2298 0 1 2610
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_ainv__1
timestamp 1734143760
transform 1 0 2628 0 1 2620
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_ainv__2
timestamp 1734143760
transform 1 0 2526 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_ainv__3
timestamp 1734143760
transform 1 0 2580 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  copy__ctrl__shift__splits_al_50_6
timestamp 1734143796
transform 1 0 2406 0 1 2380
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  copy__ctrl__shift__splits_anor__2
timestamp 1734143909
transform 1 0 2676 0 1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  copy__ctrl__shift__splits_anor__3
timestamp 1734143909
transform 1 0 2304 0 1 2850
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  copy__ctrl__shift__splits_aor__1
timestamp 1734143975
transform 1 0 2634 0 -1 3080
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  copy__ctrl__shift__splits_apulseG_aand
timestamp 1734143631
transform 1 0 2334 0 1 2370
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai
timestamp 1734143760
transform 1 0 2412 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai1
timestamp 1734143760
transform 1 0 2364 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai2
timestamp 1734143760
transform 1 0 2310 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai3
timestamp 1734143760
transform 1 0 2256 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai4
timestamp 1734143760
transform 1 0 2250 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai5
timestamp 1734143760
transform 1 0 2292 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai6
timestamp 1734143760
transform 1 0 2322 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai7
timestamp 1734143760
transform 1 0 2364 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai8
timestamp 1734143760
transform 1 0 2364 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift__splits_apulseG_ai9
timestamp 1734143760
transform 1 0 2406 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  copy__ctrl__shift__splits_apulseG_anor
timestamp 1734143909
transform 1 0 2412 0 -1 2610
box 0 0 42 80
use _0_0cell_0_0g0n1n2naa_012aax0  copy__ctrl__shift_acelem_acx0
timestamp 1734143631
transform 1 0 2334 0 -1 3080
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift_adelay1_acx0
timestamp 1734143631
transform 1 0 2418 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift_adelay1_acx1
timestamp 1734143631
transform 1 0 2472 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift_adelay1_acx2
timestamp 1734143631
transform 1 0 2526 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift_adelay1_acx3
timestamp 1734143631
transform 1 0 2580 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift_adelay1_acx4
timestamp 1734143631
transform 1 0 2634 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift_adelay1_acx5
timestamp 1734143631
transform 1 0 2634 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift_adelay1_acx6
timestamp 1734143631
transform 1 0 2604 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__ctrl__shift_adelay1_acx7
timestamp 1734143631
transform 1 0 2550 0 1 3090
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_ainv__1
timestamp 1734143760
transform 1 0 2418 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_ainv__2
timestamp 1734143760
transform 1 0 2358 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_ainv__3
timestamp 1734143760
transform 1 0 2250 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  copy__ctrl__shift_al_50_6
timestamp 1734143796
transform 1 0 1980 0 1 3100
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  copy__ctrl__shift_anor__2
timestamp 1734143909
transform 1 0 2466 0 -1 3090
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  copy__ctrl__shift_anor__3
timestamp 1734143909
transform 1 0 2562 0 -1 2610
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  copy__ctrl__shift_aor__1
timestamp 1734143975
transform 1 0 2262 0 -1 3080
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  copy__ctrl__shift_apulseG_aand
timestamp 1734143631
transform 1 0 2472 0 1 3090
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai
timestamp 1734143760
transform 1 0 2310 0 1 3340
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai1
timestamp 1734143760
transform 1 0 2502 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai2
timestamp 1734143760
transform 1 0 2568 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai3
timestamp 1734143760
transform 1 0 2436 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai4
timestamp 1734143760
transform 1 0 2376 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai5
timestamp 1734143760
transform 1 0 2274 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai6
timestamp 1734143760
transform 1 0 2322 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai7
timestamp 1734143760
transform 1 0 2334 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai8
timestamp 1734143760
transform 1 0 2376 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__ctrl__shift_apulseG_ai9
timestamp 1734143760
transform 1 0 2424 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  copy__ctrl__shift_apulseG_anor
timestamp 1734143909
transform 1 0 2358 0 1 3330
box 0 0 42 80
use _0_0cell_0_0g0n1n2naa_012aax0  copy__P__comparisons_acelem_acx0
timestamp 1734143631
transform 1 0 2718 0 -1 3560
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  copy__P__comparisons_adelay1_acx0
timestamp 1734143631
transform 1 0 2688 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P__comparisons_adelay1_acx1
timestamp 1734143631
transform 1 0 2652 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P__comparisons_adelay1_acx2
timestamp 1734143631
transform 1 0 2592 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P__comparisons_adelay1_acx3
timestamp 1734143631
transform 1 0 2532 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P__comparisons_adelay1_acx4
timestamp 1734143631
transform 1 0 2550 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P__comparisons_adelay1_acx5
timestamp 1734143631
transform 1 0 2496 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P__comparisons_adelay1_acx6
timestamp 1734143631
transform 1 0 2442 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P__comparisons_adelay1_acx7
timestamp 1734143631
transform 1 0 2394 0 1 3570
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_ainv__1
timestamp 1734143760
transform 1 0 2682 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_ainv__2
timestamp 1734143760
transform 1 0 2736 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_ainv__3
timestamp 1734143760
transform 1 0 2712 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  copy__P__comparisons_al_50_6
timestamp 1734143796
transform 1 0 3180 0 1 2380
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P__comparisons_al_51_6
timestamp 1734143796
transform 1 0 2946 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P__comparisons_al_52_6
timestamp 1734143796
transform 1 0 3408 0 -1 2360
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P__comparisons_al_53_6
timestamp 1734143796
transform 1 0 3042 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P__comparisons_al_54_6
timestamp 1734143796
transform 1 0 3138 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P__comparisons_al_55_6
timestamp 1734143796
transform 1 0 3318 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P__comparisons_al_56_6
timestamp 1734143796
transform 1 0 2958 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P__comparisons_al_57_6
timestamp 1734143796
transform 1 0 3210 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  copy__P__comparisons_anor__2
timestamp 1734143909
transform 1 0 2706 0 1 3800
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  copy__P__comparisons_anor__3
timestamp 1734143909
transform 1 0 2700 0 -1 4030
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  copy__P__comparisons_aor__1
timestamp 1734143975
transform 1 0 2700 0 1 3100
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  copy__P__comparisons_apulseG_aand
timestamp 1734143631
transform 1 0 3498 0 1 2370
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai
timestamp 1734143760
transform 1 0 2832 0 1 2620
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai1
timestamp 1734143760
transform 1 0 3564 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai2
timestamp 1734143760
transform 1 0 3606 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai3
timestamp 1734143760
transform 1 0 3714 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai4
timestamp 1734143760
transform 1 0 3744 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai5
timestamp 1734143760
transform 1 0 3672 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai6
timestamp 1734143760
transform 1 0 3606 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai7
timestamp 1734143760
transform 1 0 3552 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai8
timestamp 1734143760
transform 1 0 3504 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P__comparisons_apulseG_ai9
timestamp 1734143760
transform 1 0 3504 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  copy__P__comparisons_apulseG_anor
timestamp 1734143909
transform 1 0 3000 0 1 2370
box 0 0 42 80
use _0_0cell_0_0g0n1n2naa_012aax0  copy__P_acelem_acx0
timestamp 1734143631
transform 1 0 2808 0 -1 2600
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  copy__P_adelay1_acx0
timestamp 1734143631
transform 1 0 2880 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P_adelay1_acx1
timestamp 1734143631
transform 1 0 2892 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P_adelay1_acx2
timestamp 1734143631
transform 1 0 3012 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P_adelay1_acx3
timestamp 1734143631
transform 1 0 2916 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P_adelay1_acx4
timestamp 1734143631
transform 1 0 2784 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P_adelay1_acx5
timestamp 1734143631
transform 1 0 2712 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P_adelay1_acx6
timestamp 1734143631
transform 1 0 2724 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  copy__P_adelay1_acx7
timestamp 1734143631
transform 1 0 2820 0 -1 2850
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  copy__P_ainv__1
timestamp 1734143760
transform 1 0 2778 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_ainv__2
timestamp 1734143760
transform 1 0 2916 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_ainv__3
timestamp 1734143760
transform 1 0 2640 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  copy__P_al_50_6
timestamp 1734143796
transform 1 0 3258 0 -1 2360
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P_al_51_6
timestamp 1734143796
transform 1 0 3060 0 1 2380
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P_al_52_6
timestamp 1734143796
transform 1 0 3336 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P_al_53_6
timestamp 1734143796
transform 1 0 3138 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P_al_54_6
timestamp 1734143796
transform 1 0 3180 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P_al_55_6
timestamp 1734143796
transform 1 0 3270 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P_al_56_6
timestamp 1734143796
transform 1 0 3114 0 -1 2360
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  copy__P_al_57_6
timestamp 1734143796
transform 1 0 3294 0 1 2380
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  copy__P_anor__2
timestamp 1734143909
transform 1 0 2760 0 1 2610
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  copy__P_anor__3
timestamp 1734143909
transform 1 0 2934 0 1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  copy__P_aor__1
timestamp 1734143975
transform 1 0 2670 0 -1 2600
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  copy__P_apulseG_aand
timestamp 1734143631
transform 1 0 3276 0 -1 2130
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai
timestamp 1734143760
transform 1 0 2880 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai1
timestamp 1734143760
transform 1 0 3414 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai2
timestamp 1734143760
transform 1 0 3432 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai3
timestamp 1734143760
transform 1 0 3468 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai4
timestamp 1734143760
transform 1 0 3612 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai5
timestamp 1734143760
transform 1 0 3708 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai6
timestamp 1734143760
transform 1 0 3810 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai7
timestamp 1734143760
transform 1 0 3522 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai8
timestamp 1734143760
transform 1 0 3444 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  copy__P_apulseG_ai9
timestamp 1734143760
transform 1 0 3372 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  copy__P_apulseG_anor
timestamp 1734143909
transform 1 0 3030 0 -1 2370
box 0 0 42 80
use _0_0cell_0_0g0n1n2naa_012aax0  cp1_acelem_acx0
timestamp 1734143631
transform 1 0 1800 0 1 2620
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  cp1_adelay1_acx0
timestamp 1734143631
transform 1 0 1884 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  cp1_adelay1_acx1
timestamp 1734143631
transform 1 0 1854 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  cp1_adelay1_acx2
timestamp 1734143631
transform 1 0 1908 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  cp1_adelay1_acx3
timestamp 1734143631
transform 1 0 1890 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  cp1_adelay1_acx4
timestamp 1734143631
transform 1 0 1944 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  cp1_adelay1_acx5
timestamp 1734143631
transform 1 0 1920 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  cp1_adelay1_acx6
timestamp 1734143631
transform 1 0 1860 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  cp1_adelay1_acx7
timestamp 1734143631
transform 1 0 1794 0 -1 2370
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  cp1_ainv__1
timestamp 1734143760
transform 1 0 2202 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_ainv__2
timestamp 1734143760
transform 1 0 1548 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_ainv__3
timestamp 1734143760
transform 1 0 1686 0 1 2620
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  cp1_al_50_6
timestamp 1734143796
transform 1 0 1704 0 -1 2840
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  cp1_anor__2
timestamp 1734143909
transform 1 0 2196 0 1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  cp1_anor__3
timestamp 1734143909
transform 1 0 1494 0 -1 2850
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  cp1_aor__1
timestamp 1734143975
transform 1 0 1734 0 1 2620
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  cp1_apulseG_aand
timestamp 1734143631
transform 1 0 1632 0 -1 2850
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai1
timestamp 1734143760
transform 1 0 1842 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai2
timestamp 1734143760
transform 1 0 1776 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai3
timestamp 1734143760
transform 1 0 1716 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai4
timestamp 1734143760
transform 1 0 1488 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai5
timestamp 1734143760
transform 1 0 1518 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai6
timestamp 1734143760
transform 1 0 1554 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai7
timestamp 1734143760
transform 1 0 1602 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai8
timestamp 1734143760
transform 1 0 1656 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai
timestamp 1734143760
transform 1 0 1866 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  cp1_apulseG_ai9
timestamp 1734143760
transform 1 0 1590 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  cp1_apulseG_anor
timestamp 1734143909
transform 1 0 1812 0 -1 2850
box 0 0 42 80
use _0_0cell_0_0g0n1n2naa_012aax0  ctrl__lower__copy_acelem_acx0
timestamp 1734143631
transform 1 0 1644 0 1 3340
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  ctrl__lower__copy_adelay1_acx0
timestamp 1734143631
transform 1 0 1680 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  ctrl__lower__copy_adelay1_acx1
timestamp 1734143631
transform 1 0 1698 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  ctrl__lower__copy_adelay1_acx2
timestamp 1734143631
transform 1 0 1812 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  ctrl__lower__copy_adelay1_acx3
timestamp 1734143631
transform 1 0 1800 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  ctrl__lower__copy_adelay1_acx4
timestamp 1734143631
transform 1 0 1866 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  ctrl__lower__copy_adelay1_acx5
timestamp 1734143631
transform 1 0 1884 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  ctrl__lower__copy_adelay1_acx6
timestamp 1734143631
transform 1 0 1932 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  ctrl__lower__copy_adelay1_acx7
timestamp 1734143631
transform 1 0 2004 0 -1 3090
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_ainv__1
timestamp 1734143760
transform 1 0 1656 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_ainv__2
timestamp 1734143760
transform 1 0 1662 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_ainv__3
timestamp 1734143760
transform 1 0 1392 0 1 3340
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  ctrl__lower__copy_al_50_6
timestamp 1734143796
transform 1 0 1824 0 -1 3560
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  ctrl__lower__copy_anor__2
timestamp 1734143909
transform 1 0 1788 0 1 3570
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  ctrl__lower__copy_anor__3
timestamp 1734143909
transform 1 0 1728 0 -1 3330
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  ctrl__lower__copy_aor__1
timestamp 1734143975
transform 1 0 1446 0 1 3340
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  ctrl__lower__copy_apulseG_aand
timestamp 1734143631
transform 1 0 1746 0 -1 3570
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai
timestamp 1734143760
transform 1 0 1590 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai1
timestamp 1734143760
transform 1 0 1620 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai2
timestamp 1734143760
transform 1 0 1584 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai3
timestamp 1734143760
transform 1 0 1548 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai4
timestamp 1734143760
transform 1 0 1518 0 1 3340
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai5
timestamp 1734143760
transform 1 0 1560 0 1 3340
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai6
timestamp 1734143760
transform 1 0 1602 0 1 3340
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai7
timestamp 1734143760
transform 1 0 1590 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai8
timestamp 1734143760
transform 1 0 1728 0 1 3340
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  ctrl__lower__copy_apulseG_ai9
timestamp 1734143760
transform 1 0 1770 0 1 3340
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  ctrl__lower__copy_apulseG_anor
timestamp 1734143909
transform 1 0 1626 0 1 3570
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  merge_aand1
timestamp 1734143631
transform 1 0 2400 0 1 2130
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  merge_aand2
timestamp 1734143631
transform 1 0 2496 0 -1 2370
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  merge_acelem1_acx0
timestamp 1734143631
transform 1 0 2562 0 1 2140
box 6 10 65 70
use _0_0cell_0_0g0n1n2naa_012aax0  merge_acelem2_acx0
timestamp 1734143631
transform 1 0 2706 0 -1 2360
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  merge_adelay1_acx0
timestamp 1734143631
transform 1 0 2640 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay1_acx1
timestamp 1734143631
transform 1 0 2640 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay1_acx2
timestamp 1734143631
transform 1 0 2574 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay1_acx3
timestamp 1734143631
transform 1 0 2562 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay1_acx4
timestamp 1734143631
transform 1 0 2604 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay1_acx5
timestamp 1734143631
transform 1 0 2622 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay1_acx6
timestamp 1734143631
transform 1 0 2568 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay1_acx7
timestamp 1734143631
transform 1 0 2448 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay2_acx0
timestamp 1734143631
transform 1 0 2706 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay2_acx1
timestamp 1734143631
transform 1 0 3174 0 1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay2_acx2
timestamp 1734143631
transform 1 0 3570 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay2_acx3
timestamp 1734143631
transform 1 0 3666 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay2_acx4
timestamp 1734143631
transform 1 0 3738 0 1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay2_acx5
timestamp 1734143631
transform 1 0 3858 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay2_acx6
timestamp 1734143631
transform 1 0 3912 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay2_acx7
timestamp 1734143631
transform 1 0 4062 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay3_acx0
timestamp 1734143631
transform 1 0 4140 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay3_acx1
timestamp 1734143631
transform 1 0 4182 0 -1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay3_acx2
timestamp 1734143631
transform 1 0 4188 0 1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay3_acx3
timestamp 1734143631
transform 1 0 4188 0 -1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay3_acx4
timestamp 1734143631
transform 1 0 4188 0 -1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay3_acx5
timestamp 1734143631
transform 1 0 4188 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay3_acx6
timestamp 1734143631
transform 1 0 4188 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  merge_adelay3_acx7
timestamp 1734143631
transform 1 0 4188 0 1 200
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  merge_ainv1__Cd
timestamp 1734143760
transform 1 0 2520 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Cf
timestamp 1734143760
transform 1 0 2658 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Ct
timestamp 1734143760
transform 1 0 2466 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__L1
timestamp 1734143760
transform 1 0 2442 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__L2
timestamp 1734143760
transform 1 0 3150 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Ra
timestamp 1734143760
transform 1 0 2616 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Rd1
timestamp 1734143760
transform 1 0 1992 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Rd2
timestamp 1734143760
transform 1 0 2346 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Rd3
timestamp 1734143760
transform 1 0 2724 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Rd4
timestamp 1734143760
transform 1 0 2052 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Rd5
timestamp 1734143760
transform 1 0 2322 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Rd6
timestamp 1734143760
transform 1 0 1860 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Rd7
timestamp 1734143760
transform 1 0 2106 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_ainv__Rd8
timestamp 1734143760
transform 1 0 2154 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  merge_al_50_6
timestamp 1734143796
transform 1 0 2034 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  merge_al_51_6
timestamp 1734143796
transform 1 0 2388 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  merge_al_52_6
timestamp 1734143796
transform 1 0 2610 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  merge_al_53_6
timestamp 1734143796
transform 1 0 2106 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  merge_al_54_6
timestamp 1734143796
transform 1 0 2358 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  merge_al_55_6
timestamp 1734143796
transform 1 0 1902 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  merge_al_56_6
timestamp 1734143796
transform 1 0 2136 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  merge_al_57_6
timestamp 1734143796
transform 1 0 2226 0 -1 1890
box 0 0 96 80
use _0_0std_0_0cells_0_0MUX2X1  merge_amux_50_6
timestamp 1734143875
transform 1 0 2142 0 1 1900
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  merge_amux_51_6
timestamp 1734143875
transform 1 0 2502 0 1 1900
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  merge_amux_52_6
timestamp 1734143875
transform 1 0 2496 0 1 1660
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  merge_amux_53_6
timestamp 1734143875
transform 1 0 2226 0 1 1660
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  merge_amux_54_6
timestamp 1734143875
transform 1 0 2460 0 -1 1660
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  merge_amux_55_6
timestamp 1734143875
transform 1 0 2010 0 -1 1660
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  merge_amux_56_6
timestamp 1734143875
transform 1 0 2232 0 -1 1660
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  merge_amux_57_6
timestamp 1734143875
transform 1 0 2244 0 1 1900
box 0 0 90 90
use _0_0std_0_0cells_0_0NOR2X1  merge_anor__Ra
timestamp 1734143909
transform 1 0 2568 0 -1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  merge_aor__Cf
timestamp 1734143975
transform 1 0 2700 0 1 2140
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  merge_aor__L2
timestamp 1734143975
transform 1 0 2940 0 1 2140
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  merge_aor
timestamp 1734143975
transform 1 0 2640 0 1 2140
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  merge_aor__Ct
timestamp 1734143975
transform 1 0 2502 0 1 2140
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  merge_aor__L1
timestamp 1734143975
transform 1 0 2502 0 -1 2120
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  merge_apulseG_aand
timestamp 1734143631
transform 1 0 2364 0 -1 1900
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai
timestamp 1734143760
transform 1 0 2652 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai1
timestamp 1734143760
transform 1 0 2610 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai2
timestamp 1734143760
transform 1 0 2664 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai3
timestamp 1734143760
transform 1 0 2718 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai4
timestamp 1734143760
transform 1 0 2628 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai5
timestamp 1734143760
transform 1 0 2544 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai6
timestamp 1734143760
transform 1 0 2466 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai7
timestamp 1734143760
transform 1 0 2448 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai8
timestamp 1734143760
transform 1 0 2394 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  merge_apulseG_ai9
timestamp 1734143760
transform 1 0 2340 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  merge_apulseG_anor
timestamp 1734143909
transform 1 0 2586 0 -1 2130
box 0 0 42 80
use circuitwell  npwells
timestamp 0
transform 1 0 60 0 1 180
box 0 0 1 1
use _0_0std_0_0cells_0_0AND2X1  or_aelem__c_aa1
timestamp 1734143631
transform 1 0 1902 0 1 3330
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  or_aelem__c_aa2
timestamp 1734143631
transform 1 0 1986 0 -1 3330
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  or_aelem__c_ac1_acx0
timestamp 1734143631
transform 1 0 2070 0 -1 3320
box 6 10 65 70
use _0_0cell_0_0g0n_0x1  or_aelem__c_ac1_acx1
timestamp 1734143631
transform 1 0 2040 0 1 3350
box 6 10 21 40
use _0_0cell_0_0g0n_0x0  or_aelem__c_adelay_acx0
timestamp 1734143631
transform 1 0 2202 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  or_aelem__c_adelay_acx1
timestamp 1734143631
transform 1 0 2256 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  or_aelem__c_adelay_acx2
timestamp 1734143631
transform 1 0 2166 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  or_aelem__c_adelay_acx3
timestamp 1734143631
transform 1 0 2130 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  or_aelem__c_adelay_acx4
timestamp 1734143631
transform 1 0 2172 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  or_aelem__c_adelay_acx5
timestamp 1734143631
transform 1 0 2208 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  or_aelem__c_adelay_acx6
timestamp 1734143631
transform 1 0 2202 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  or_aelem__c_adelay_acx7
timestamp 1734143631
transform 1 0 2286 0 1 3090
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  or_aelem__c_ai1
timestamp 1734143760
transform 1 0 1932 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  or_aelem__c_an1
timestamp 1734143909
transform 1 0 2220 0 -1 3330
box 0 0 42 80
use _0_0std_0_0cells_0_0LATCH  or_alatch
timestamp 1734143796
transform 1 0 2082 0 1 3340
box 0 0 96 80
use _0_0std_0_0cells_0_0OR2X1  or_aor
timestamp 1734143975
transform 1 0 1974 0 1 3340
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  or_apulseG_aand
timestamp 1734143631
transform 1 0 1992 0 -1 3570
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai1
timestamp 1734143760
transform 1 0 2010 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai2
timestamp 1734143760
transform 1 0 1962 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai3
timestamp 1734143760
transform 1 0 1944 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai4
timestamp 1734143760
transform 1 0 1872 0 1 3810
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai5
timestamp 1734143760
transform 1 0 1806 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai6
timestamp 1734143760
transform 1 0 1860 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai7
timestamp 1734143760
transform 1 0 1914 0 -1 3790
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai
timestamp 1734143760
transform 1 0 2064 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai8
timestamp 1734143760
transform 1 0 1902 0 1 3580
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  or_apulseG_ai9
timestamp 1734143760
transform 1 0 1938 0 -1 3560
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  or_apulseG_anor
timestamp 1734143909
transform 1 0 2082 0 -1 3570
box 0 0 42 80
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderLeft_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 1422 0 -1 2840
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 1524 0 1 2630
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderLeft_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 1428 0 1 2610
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 1380 0 1 2630
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderLeft_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 1500 0 1 2380
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 1446 0 1 2150
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderLeft_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 1488 0 -1 2370
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 1572 0 -1 2350
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderLeft_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 1248 0 1 1910
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 1152 0 1 1680
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderLeft_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 1182 0 -1 1900
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 1122 0 -1 1880
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderLeft_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 1020 0 1 1200
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 1110 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderLeft_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 1026 0 -1 1190
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 1116 0 1 1210
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderLeft_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 996 0 1 960
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 1044 0 -1 1400
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderLeft_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 1068 0 1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 1152 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderLeft_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 1026 0 -1 1890
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 966 0 1 1920
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderLeft_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 918 0 -1 1900
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 852 0 -1 1880
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderLeft_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 1008 0 -1 2360
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 1008 0 -1 2590
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderLeft_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 1014 0 1 2130
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 1086 0 -1 2110
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderLeft_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 1044 0 1 2620
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 1128 0 1 2630
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderLeft_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 1050 0 -1 2610
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderLeft_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 1092 0 1 2390
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  post_aadderLeft_acelem_acx0
timestamp 1734143631
transform 1 0 678 0 1 2860
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay1_acx0
timestamp 1734143631
transform 1 0 516 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay1_acx1
timestamp 1734143631
transform 1 0 492 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay1_acx2
timestamp 1734143631
transform 1 0 456 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay1_acx3
timestamp 1734143631
transform 1 0 240 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay1_acx4
timestamp 1734143631
transform 1 0 204 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay1_acx5
timestamp 1734143631
transform 1 0 168 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay1_acx6
timestamp 1734143631
transform 1 0 132 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay1_acx7
timestamp 1734143631
transform 1 0 96 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay2_acx0
timestamp 1734143631
transform 1 0 168 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay2_acx1
timestamp 1734143631
transform 1 0 210 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay2_acx2
timestamp 1734143631
transform 1 0 258 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay2_acx3
timestamp 1734143631
transform 1 0 210 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay2_acx4
timestamp 1734143631
transform 1 0 306 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay2_acx5
timestamp 1734143631
transform 1 0 276 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay2_acx6
timestamp 1734143631
transform 1 0 282 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderLeft_adelay2_acx7
timestamp 1734143631
transform 1 0 354 0 1 2610
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_ainv__l1
timestamp 1734143760
transform 1 0 486 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_ainv__l2
timestamp 1734143760
transform 1 0 546 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_ainv__r
timestamp 1734143760
transform 1 0 660 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al1_50_6
timestamp 1734143796
transform 1 0 1314 0 -1 2840
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al1_51_6
timestamp 1734143796
transform 1 0 1380 0 -1 2360
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al1_52_6
timestamp 1734143796
transform 1 0 1122 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al1_53_6
timestamp 1734143796
transform 1 0 882 0 1 1200
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al1_54_6
timestamp 1734143796
transform 1 0 918 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al1_55_6
timestamp 1734143796
transform 1 0 858 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al1_56_6
timestamp 1734143796
transform 1 0 828 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al1_57_6
timestamp 1734143796
transform 1 0 924 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al2_50_6
timestamp 1734143796
transform 1 0 1362 0 1 2860
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al2_51_6
timestamp 1734143796
transform 1 0 1428 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al2_52_6
timestamp 1734143796
transform 1 0 1392 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al2_53_6
timestamp 1734143796
transform 1 0 810 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al2_54_6
timestamp 1734143796
transform 1 0 834 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al2_55_6
timestamp 1734143796
transform 1 0 810 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al2_56_6
timestamp 1734143796
transform 1 0 1080 0 -1 2360
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderLeft_al2_57_6
timestamp 1734143796
transform 1 0 948 0 -1 2840
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  post_aadderLeft_anor
timestamp 1734143909
transform 1 0 642 0 -1 2610
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  post_aadderLeft_aor__l1
timestamp 1734143975
transform 1 0 528 0 -1 3080
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  post_aadderLeft_aor__l2
timestamp 1734143975
transform 1 0 594 0 1 3100
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  post_aadderLeft_apulseG_aand
timestamp 1734143631
transform 1 0 1116 0 -1 2850
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai1
timestamp 1734143760
transform 1 0 978 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai2
timestamp 1734143760
transform 1 0 1008 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai3
timestamp 1734143760
transform 1 0 1038 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai4
timestamp 1734143760
transform 1 0 1068 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai
timestamp 1734143760
transform 1 0 828 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai5
timestamp 1734143760
transform 1 0 1050 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai6
timestamp 1734143760
transform 1 0 948 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai7
timestamp 1734143760
transform 1 0 1002 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai8
timestamp 1734143760
transform 1 0 1092 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderLeft_apulseG_ai9
timestamp 1734143760
transform 1 0 1080 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  post_aadderLeft_apulseG_anor
timestamp 1734143909
transform 1 0 864 0 -1 3090
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  post_aadderLeft_atoGND
timestamp 1734144021
transform 1 0 1458 0 1 2870
box 0 0 30 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderRight_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 1230 0 1 2860
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 1284 0 1 2630
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderRight_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 1290 0 1 2850
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 1332 0 1 2630
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderRight_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 1254 0 -1 2600
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 1284 0 -1 2350
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderRight_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 1236 0 1 2370
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 1314 0 -1 2350
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderRight_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 1266 0 -1 2120
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 1338 0 1 1920
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderRight_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 1362 0 -1 2130
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 1356 0 -1 1880
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderRight_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 1050 0 1 1670
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 894 0 -1 1640
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderRight_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 1026 0 -1 1660
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 960 0 -1 1640
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderRight_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 846 0 1 1430
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 834 0 1 1680
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderRight_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 918 0 1 1420
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 1104 0 -1 1400
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderRight_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 738 0 1 1910
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 834 0 -1 2110
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderRight_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 738 0 -1 1900
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 678 0 -1 1880
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderRight_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 942 0 1 2140
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 972 0 1 2390
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderRight_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 966 0 -1 2130
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 1044 0 -1 2110
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  post_aadderRight_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 876 0 -1 2600
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 960 0 -1 2590
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  post_aadderRight_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 870 0 1 2370
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  post_aadderRight_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 1032 0 1 2390
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  post_aadderRight_acelem_acx0
timestamp 1734143631
transform 1 0 750 0 -1 3080
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay1_acx0
timestamp 1734143631
transform 1 0 708 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay1_acx1
timestamp 1734143631
transform 1 0 672 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay1_acx2
timestamp 1734143631
transform 1 0 624 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay1_acx3
timestamp 1734143631
transform 1 0 576 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay1_acx4
timestamp 1734143631
transform 1 0 528 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay1_acx5
timestamp 1734143631
transform 1 0 348 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay1_acx6
timestamp 1734143631
transform 1 0 312 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay1_acx7
timestamp 1734143631
transform 1 0 276 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay2_acx0
timestamp 1734143631
transform 1 0 354 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay2_acx1
timestamp 1734143631
transform 1 0 306 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay2_acx2
timestamp 1734143631
transform 1 0 282 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay2_acx3
timestamp 1734143631
transform 1 0 354 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay2_acx4
timestamp 1734143631
transform 1 0 360 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay2_acx5
timestamp 1734143631
transform 1 0 366 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay2_acx6
timestamp 1734143631
transform 1 0 390 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_aadderRight_adelay2_acx7
timestamp 1734143631
transform 1 0 486 0 -1 2610
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_ainv__l1
timestamp 1734143760
transform 1 0 654 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_ainv__l2
timestamp 1734143760
transform 1 0 660 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_ainv__r
timestamp 1734143760
transform 1 0 708 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al1_50_6
timestamp 1734143796
transform 1 0 1128 0 1 2860
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al1_51_6
timestamp 1734143796
transform 1 0 1356 0 1 2380
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al1_52_6
timestamp 1734143796
transform 1 0 1140 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al1_53_6
timestamp 1734143796
transform 1 0 1002 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al1_54_6
timestamp 1734143796
transform 1 0 912 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al1_55_6
timestamp 1734143796
transform 1 0 648 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al1_56_6
timestamp 1734143796
transform 1 0 864 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al1_57_6
timestamp 1734143796
transform 1 0 762 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al2_50_6
timestamp 1734143796
transform 1 0 1272 0 -1 3080
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al2_51_6
timestamp 1734143796
transform 1 0 1140 0 -1 2600
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al2_52_6
timestamp 1734143796
transform 1 0 1098 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al2_53_6
timestamp 1734143796
transform 1 0 954 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al2_54_6
timestamp 1734143796
transform 1 0 774 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al2_55_6
timestamp 1734143796
transform 1 0 630 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al2_56_6
timestamp 1734143796
transform 1 0 858 0 -1 2360
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_aadderRight_al2_57_6
timestamp 1734143796
transform 1 0 810 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  post_aadderRight_anor
timestamp 1734143909
transform 1 0 702 0 -1 2610
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  post_aadderRight_aor__l1
timestamp 1734143975
transform 1 0 690 0 -1 3080
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  post_aadderRight_aor__l2
timestamp 1734143975
transform 1 0 696 0 1 3100
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  post_aadderRight_apulseG_aand
timestamp 1734143631
transform 1 0 912 0 -1 3090
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai2
timestamp 1734143760
transform 1 0 774 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai3
timestamp 1734143760
transform 1 0 840 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai4
timestamp 1734143760
transform 1 0 912 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai5
timestamp 1734143760
transform 1 0 996 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai6
timestamp 1734143760
transform 1 0 1176 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai7
timestamp 1734143760
transform 1 0 1146 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai8
timestamp 1734143760
transform 1 0 1062 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai9
timestamp 1734143760
transform 1 0 978 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai
timestamp 1734143760
transform 1 0 816 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_aadderRight_apulseG_ai1
timestamp 1734143760
transform 1 0 762 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  post_aadderRight_apulseG_anor
timestamp 1734143909
transform 1 0 888 0 1 3090
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  post_aadderRight_atoGND
timestamp 1734144021
transform 1 0 1230 0 -1 3070
box 0 0 30 50
use _0_0cell_0_0g0n1n2naa_012aax0  post_acp1_acelem_acx0
timestamp 1734143631
transform 1 0 1230 0 -1 2840
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  post_acp1_adelay1_acx0
timestamp 1734143631
transform 1 0 1188 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_acp1_adelay1_acx1
timestamp 1734143631
transform 1 0 1146 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_acp1_adelay1_acx2
timestamp 1734143631
transform 1 0 1104 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_acp1_adelay1_acx3
timestamp 1734143631
transform 1 0 882 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_acp1_adelay1_acx4
timestamp 1734143631
transform 1 0 852 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_acp1_adelay1_acx5
timestamp 1734143631
transform 1 0 810 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_acp1_adelay1_acx6
timestamp 1734143631
transform 1 0 762 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_acp1_adelay1_acx7
timestamp 1734143631
transform 1 0 588 0 -1 2610
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  post_acp1_ainv__1
timestamp 1734143760
transform 1 0 918 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_ainv__2
timestamp 1734143760
transform 1 0 1188 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_ainv__3
timestamp 1734143760
transform 1 0 1602 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  post_acp1_al_50_6
timestamp 1734143796
transform 1 0 1572 0 1 2620
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  post_acp1_anor__2
timestamp 1734143909
transform 1 0 756 0 -1 2850
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  post_acp1_anor__3
timestamp 1734143909
transform 1 0 1176 0 1 2610
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  post_acp1_aor__1
timestamp 1734143975
transform 1 0 1584 0 -1 2600
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  post_acp1_apulseG_aand
timestamp 1734143631
transform 1 0 1518 0 -1 3090
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai1
timestamp 1734143760
transform 1 0 1572 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai2
timestamp 1734143760
transform 1 0 1518 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai3
timestamp 1734143760
transform 1 0 1440 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai4
timestamp 1734143760
transform 1 0 1356 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai5
timestamp 1734143760
transform 1 0 1266 0 -1 3320
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai6
timestamp 1734143760
transform 1 0 1230 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai7
timestamp 1734143760
transform 1 0 1308 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai9
timestamp 1734143760
transform 1 0 1476 0 -1 3080
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai
timestamp 1734143760
transform 1 0 1446 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_acp1_apulseG_ai8
timestamp 1734143760
transform 1 0 1380 0 1 3100
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  post_acp1_apulseG_anor
timestamp 1734143909
transform 1 0 1506 0 1 3090
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  post_amerge_aand1
timestamp 1734143631
transform 1 0 564 0 -1 2130
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  post_amerge_aand2
timestamp 1734143631
transform 1 0 630 0 -1 2130
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  post_amerge_acelem1_acx0
timestamp 1734143631
transform 1 0 684 0 -1 2360
box 6 10 65 70
use _0_0cell_0_0g0n1n2naa_012aax0  post_amerge_acelem2_acx0
timestamp 1734143631
transform 1 0 774 0 -1 2360
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  post_amerge_adelay1_acx0
timestamp 1734143631
transform 1 0 570 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay1_acx1
timestamp 1734143631
transform 1 0 558 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay1_acx2
timestamp 1734143631
transform 1 0 498 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay1_acx3
timestamp 1734143631
transform 1 0 516 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay1_acx4
timestamp 1734143631
transform 1 0 450 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay1_acx5
timestamp 1734143631
transform 1 0 462 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay1_acx6
timestamp 1734143631
transform 1 0 516 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay1_acx7
timestamp 1734143631
transform 1 0 576 0 1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay2_acx0
timestamp 1734143631
transform 1 0 1656 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay2_acx1
timestamp 1734143631
transform 1 0 1704 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay2_acx2
timestamp 1734143631
transform 1 0 1752 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay2_acx3
timestamp 1734143631
transform 1 0 1800 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay2_acx4
timestamp 1734143631
transform 1 0 1728 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay2_acx5
timestamp 1734143631
transform 1 0 1788 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay2_acx6
timestamp 1734143631
transform 1 0 1842 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay2_acx7
timestamp 1734143631
transform 1 0 1998 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay3_acx0
timestamp 1734143631
transform 1 0 2052 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay3_acx1
timestamp 1734143631
transform 1 0 2100 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay3_acx2
timestamp 1734143631
transform 1 0 2148 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay3_acx3
timestamp 1734143631
transform 1 0 2094 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay3_acx4
timestamp 1734143631
transform 1 0 2274 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay3_acx5
timestamp 1734143631
transform 1 0 2268 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay3_acx6
timestamp 1734143631
transform 1 0 2322 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_amerge_adelay3_acx7
timestamp 1734143631
transform 1 0 2382 0 -1 2130
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv1__Cd
timestamp 1734143760
transform 1 0 642 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Cf
timestamp 1734143760
transform 1 0 696 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Ct
timestamp 1734143760
transform 1 0 582 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__L1
timestamp 1734143760
transform 1 0 492 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__L2
timestamp 1734143760
transform 1 0 540 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Ra
timestamp 1734143760
transform 1 0 1344 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Rd1
timestamp 1734143760
transform 1 0 1986 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Rd2
timestamp 1734143760
transform 1 0 2034 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Rd3
timestamp 1734143760
transform 1 0 2088 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Rd4
timestamp 1734143760
transform 1 0 1968 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Rd5
timestamp 1734143760
transform 1 0 1992 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Rd6
timestamp 1734143760
transform 1 0 1920 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Rd7
timestamp 1734143760
transform 1 0 2022 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_ainv__Rd8
timestamp 1734143760
transform 1 0 1932 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  post_amerge_al_50_6
timestamp 1734143796
transform 1 0 1884 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_amerge_al_51_6
timestamp 1734143796
transform 1 0 1812 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_amerge_al_52_6
timestamp 1734143796
transform 1 0 1878 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_amerge_al_53_6
timestamp 1734143796
transform 1 0 1638 0 -1 1890
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_amerge_al_54_6
timestamp 1734143796
transform 1 0 1524 0 -1 1890
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_amerge_al_55_6
timestamp 1734143796
transform 1 0 1644 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_amerge_al_56_6
timestamp 1734143796
transform 1 0 1518 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_amerge_al_57_6
timestamp 1734143796
transform 1 0 1764 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0MUX2X1  post_amerge_amux_50_6
timestamp 1734143875
transform 1 0 1326 0 -1 2610
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  post_amerge_amux_51_6
timestamp 1734143875
transform 1 0 1482 0 1 2130
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  post_amerge_amux_52_6
timestamp 1734143875
transform 1 0 1410 0 -1 1900
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  post_amerge_amux_53_6
timestamp 1734143875
transform 1 0 1134 0 -1 1660
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  post_amerge_amux_54_6
timestamp 1734143875
transform 1 0 1110 0 1 1420
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  post_amerge_amux_55_6
timestamp 1734143875
transform 1 0 744 0 1 1660
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  post_amerge_amux_56_6
timestamp 1734143875
transform 1 0 1008 0 1 1900
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  post_amerge_amux_57_6
timestamp 1734143875
transform 1 0 1188 0 -1 2370
box 0 0 90 90
use _0_0std_0_0cells_0_0NOR2X1  post_amerge_anor__Ra
timestamp 1734143909
transform 1 0 1980 0 -1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  post_amerge_aor
timestamp 1734143975
transform 1 0 786 0 1 2380
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  post_amerge_aor__Cf
timestamp 1734143975
transform 1 0 750 0 1 2140
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  post_amerge_aor__Ct
timestamp 1734143975
transform 1 0 612 0 -1 2360
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  post_amerge_aor__L1
timestamp 1734143975
transform 1 0 624 0 1 2380
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  post_amerge_aor__L2
timestamp 1734143975
transform 1 0 702 0 1 2380
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  post_amerge_apulseG_aand
timestamp 1734143631
transform 1 0 1680 0 1 2130
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai
timestamp 1734143760
transform 1 0 1668 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai1
timestamp 1734143760
transform 1 0 1668 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai2
timestamp 1734143760
transform 1 0 1614 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai3
timestamp 1734143760
transform 1 0 1632 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai4
timestamp 1734143760
transform 1 0 1584 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai5
timestamp 1734143760
transform 1 0 1530 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai6
timestamp 1734143760
transform 1 0 1590 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai7
timestamp 1734143760
transform 1 0 1644 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai8
timestamp 1734143760
transform 1 0 1698 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_amerge_apulseG_ai9
timestamp 1734143760
transform 1 0 1758 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  post_amerge_apulseG_anor
timestamp 1734143909
transform 1 0 1722 0 -1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  post_asplit_aand1
timestamp 1734143631
transform 1 0 588 0 -1 3090
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  post_asplit_aand2
timestamp 1734143631
transform 1 0 414 0 -1 3090
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  post_asplit_acelem_acx0
timestamp 1734143631
transform 1 0 414 0 1 2380
box 6 10 65 70
use _0_0std_0_0cells_0_0LATCH  post_asplit_acontrolLatch
timestamp 1734143796
transform 1 0 606 0 1 2620
box 0 0 96 80
use _0_0cell_0_0g0n_0x0  post_asplit_adelay1_acx0
timestamp 1734143631
transform 1 0 420 0 1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay1_acx1
timestamp 1734143631
transform 1 0 420 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay1_acx2
timestamp 1734143631
transform 1 0 426 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay1_acx3
timestamp 1734143631
transform 1 0 390 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay1_acx4
timestamp 1734143631
transform 1 0 390 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay1_acx5
timestamp 1734143631
transform 1 0 324 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay1_acx6
timestamp 1734143631
transform 1 0 264 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay1_acx7
timestamp 1734143631
transform 1 0 210 0 -1 3800
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay2_acx0
timestamp 1734143631
transform 1 0 240 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay2_acx1
timestamp 1734143631
transform 1 0 318 0 1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay2_acx2
timestamp 1734143631
transform 1 0 276 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay2_acx3
timestamp 1734143631
transform 1 0 354 0 -1 3570
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay2_acx4
timestamp 1734143631
transform 1 0 384 0 1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay2_acx5
timestamp 1734143631
transform 1 0 402 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay2_acx6
timestamp 1734143631
transform 1 0 456 0 -1 3330
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  post_asplit_adelay2_acx7
timestamp 1734143631
transform 1 0 486 0 1 3090
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  post_asplit_ainv__ctr
timestamp 1734143760
transform 1 0 606 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_ainv__c
timestamp 1734143760
transform 1 0 528 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_ainv__l
timestamp 1734143760
transform 1 0 354 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_ainv__r
timestamp 1734143760
transform 1 0 432 0 1 2620
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  post_asplit_al_50_6
timestamp 1734143796
transform 1 0 1242 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_asplit_al_51_6
timestamp 1734143796
transform 1 0 1344 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_asplit_al_52_6
timestamp 1734143796
transform 1 0 1188 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_asplit_al_53_6
timestamp 1734143796
transform 1 0 1056 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_asplit_al_54_6
timestamp 1734143796
transform 1 0 936 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_asplit_al_55_6
timestamp 1734143796
transform 1 0 822 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_asplit_al_56_6
timestamp 1734143796
transform 1 0 744 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  post_asplit_al_57_6
timestamp 1734143796
transform 1 0 732 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  post_asplit_anor__R
timestamp 1734143909
transform 1 0 708 0 1 2610
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  post_asplit_aor
timestamp 1734143975
transform 1 0 792 0 1 2860
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  post_asplit_aor1
timestamp 1734143975
transform 1 0 408 0 -1 2600
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  post_asplit_aor2
timestamp 1734143975
transform 1 0 354 0 1 2380
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  post_asplit_apulseG_aand
timestamp 1734143631
transform 1 0 540 0 1 2610
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai2
timestamp 1734143760
transform 1 0 534 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai3
timestamp 1734143760
transform 1 0 468 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai4
timestamp 1734143760
transform 1 0 414 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai5
timestamp 1734143760
transform 1 0 324 0 1 2860
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai
timestamp 1734143760
transform 1 0 606 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai1
timestamp 1734143760
transform 1 0 474 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai6
timestamp 1734143760
transform 1 0 348 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai7
timestamp 1734143760
transform 1 0 414 0 -1 2840
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai8
timestamp 1734143760
transform 1 0 468 0 1 2620
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  post_asplit_apulseG_ai9
timestamp 1734143760
transform 1 0 504 0 1 2620
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  post_asplit_apulseG_anor
timestamp 1734143909
transform 1 0 534 0 -1 2850
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  post_asrc65_anor
timestamp 1734143909
transform 1 0 576 0 -1 3330
box 0 0 42 80
use _0_0std_0_0cells_0_0TIEHIX1  post_asrc65_asetGND0
timestamp 1734144001
transform 1 0 1434 0 -1 3070
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc65_asetGND1
timestamp 1734144021
transform 1 0 1536 0 -1 2590
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc65_asetGND2
timestamp 1734144021
transform 1 0 1470 0 -1 2110
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc65_asetGND3
timestamp 1734144021
transform 1 0 960 0 1 970
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc65_asetGND4
timestamp 1734144021
transform 1 0 930 0 1 970
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc65_asetGND5
timestamp 1734144021
transform 1 0 918 0 1 1920
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  post_asrc65_asetGND6
timestamp 1734144001
transform 1 0 1158 0 1 2390
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc65_asetGND7
timestamp 1734144021
transform 1 0 1044 0 -1 2830
box 0 0 30 50
use _0_0std_0_0cells_0_0NOR2X1  post_asrc97_anor
timestamp 1734143909
transform 1 0 642 0 -1 3330
box 0 0 42 80
use _0_0std_0_0cells_0_0TIEHIX1  post_asrc97_asetGND0
timestamp 1734144001
transform 1 0 1386 0 -1 3070
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc97_asetGND1
timestamp 1734144021
transform 1 0 1236 0 1 2630
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc97_asetGND2
timestamp 1734144021
transform 1 0 1206 0 1 2150
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc97_asetGND3
timestamp 1734144021
transform 1 0 1116 0 1 1680
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc97_asetGND4
timestamp 1734144021
transform 1 0 708 0 -1 1400
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  post_asrc97_asetGND5
timestamp 1734144001
transform 1 0 696 0 -1 2110
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  post_asrc97_asetGND6
timestamp 1734144001
transform 1 0 966 0 -1 2350
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  post_asrc97_asetGND7
timestamp 1734144021
transform 1 0 888 0 -1 2830
box 0 0 30 50
use circuitppnp  ppnps
timestamp 0
transform 1 0 60 0 1 180
box 0 0 1 1
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderLeft_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 3012 0 -1 1650
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 2898 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderLeft_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 2928 0 1 1420
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 2868 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderLeft_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 2850 0 -1 1410
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 2814 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderLeft_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 2790 0 1 1190
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 2628 0 1 1210
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderLeft_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 2724 0 -1 1180
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 2808 0 1 970
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderLeft_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 2718 0 1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 2664 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderLeft_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 2754 0 -1 940
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 2856 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderLeft_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 2646 0 -1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 2508 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderLeft_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 2856 0 1 720
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 2952 0 1 970
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderLeft_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 2796 0 -1 710
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 2718 0 1 490
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderLeft_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 3150 0 -1 1180
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 3150 0 1 1210
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderLeft_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 3096 0 1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 3042 0 1 730
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderLeft_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 3186 0 1 1200
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 3318 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderLeft_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 3228 0 -1 1190
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 3156 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderLeft_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 3282 0 1 960
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 3228 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderLeft_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 3294 0 -1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderLeft_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 3132 0 1 730
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  pre_aadderLeft_acelem_acx0
timestamp 1734143631
transform 1 0 3846 0 -1 1180
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay1_acx0
timestamp 1734143631
transform 1 0 3906 0 1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay1_acx1
timestamp 1734143631
transform 1 0 3960 0 1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay1_acx2
timestamp 1734143631
transform 1 0 3972 0 -1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay1_acx3
timestamp 1734143631
transform 1 0 4002 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay1_acx4
timestamp 1734143631
transform 1 0 4068 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay1_acx5
timestamp 1734143631
transform 1 0 4044 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay1_acx6
timestamp 1734143631
transform 1 0 3990 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay1_acx7
timestamp 1734143631
transform 1 0 3996 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay2_acx0
timestamp 1734143631
transform 1 0 4152 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay2_acx1
timestamp 1734143631
transform 1 0 4134 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay2_acx2
timestamp 1734143631
transform 1 0 4140 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay2_acx3
timestamp 1734143631
transform 1 0 4074 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay2_acx4
timestamp 1734143631
transform 1 0 4008 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay2_acx5
timestamp 1734143631
transform 1 0 3948 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay2_acx6
timestamp 1734143631
transform 1 0 3888 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderLeft_adelay2_acx7
timestamp 1734143631
transform 1 0 3828 0 1 200
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_ainv__l1
timestamp 1734143760
transform 1 0 3822 0 -1 1410
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_ainv__l2
timestamp 1734143760
transform 1 0 3960 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_ainv__r
timestamp 1734143760
transform 1 0 3858 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al1_50_6
timestamp 1734143796
transform 1 0 2892 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al1_51_6
timestamp 1734143796
transform 1 0 2766 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al1_52_6
timestamp 1734143796
transform 1 0 2676 0 1 1200
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al1_53_6
timestamp 1734143796
transform 1 0 2844 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al1_54_6
timestamp 1734143796
transform 1 0 2748 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al1_55_6
timestamp 1734143796
transform 1 0 3036 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al1_56_6
timestamp 1734143796
transform 1 0 3126 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al1_57_6
timestamp 1734143796
transform 1 0 3180 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al2_50_6
timestamp 1734143796
transform 1 0 3000 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al2_51_6
timestamp 1734143796
transform 1 0 2880 0 1 1200
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al2_52_6
timestamp 1734143796
transform 1 0 2862 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al2_53_6
timestamp 1734143796
transform 1 0 2928 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al2_54_6
timestamp 1734143796
transform 1 0 2928 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al2_55_6
timestamp 1734143796
transform 1 0 3036 0 1 1200
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al2_56_6
timestamp 1734143796
transform 1 0 3252 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderLeft_al2_57_6
timestamp 1734143796
transform 1 0 3348 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  pre_aadderLeft_anor
timestamp 1734143909
transform 1 0 3858 0 1 710
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  pre_aadderLeft_aor__l1
timestamp 1734143975
transform 1 0 3804 0 1 1200
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  pre_aadderLeft_aor__l2
timestamp 1734143975
transform 1 0 4032 0 1 1200
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  pre_aadderLeft_apulseG_aand
timestamp 1734143631
transform 1 0 3366 0 1 1190
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai
timestamp 1734143760
transform 1 0 3702 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai1
timestamp 1734143760
transform 1 0 3438 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai2
timestamp 1734143760
transform 1 0 3480 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai3
timestamp 1734143760
transform 1 0 3522 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai4
timestamp 1734143760
transform 1 0 3564 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai5
timestamp 1734143760
transform 1 0 3606 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai6
timestamp 1734143760
transform 1 0 3546 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai7
timestamp 1734143760
transform 1 0 3480 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai8
timestamp 1734143760
transform 1 0 3420 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderLeft_apulseG_ai9
timestamp 1734143760
transform 1 0 3366 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  pre_aadderLeft_apulseG_anor
timestamp 1734143909
transform 1 0 3606 0 1 1190
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  pre_aadderLeft_atoGND
timestamp 1734144021
transform 1 0 3072 0 1 1680
box 0 0 30 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderRight_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 2802 0 -1 1890
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 2724 0 1 1680
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderRight_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 2826 0 1 1660
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 2772 0 1 1680
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderRight_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 2694 0 1 1430
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 2562 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderRight_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 2604 0 1 1420
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 2388 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderRight_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 2538 0 1 1200
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 2598 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderRight_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 2484 0 -1 1190
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 2418 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderRight_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 2538 0 1 960
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 2676 0 -1 690
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderRight_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 2550 0 -1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 2460 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderRight_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 2784 0 -1 460
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 2886 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderRight_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 2724 0 1 200
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 2694 0 1 220
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderRight_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 3036 0 -1 700
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 3084 0 1 730
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderRight_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 3006 0 1 470
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 2958 0 1 490
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderRight_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 3360 0 -1 700
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 3264 0 1 490
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderRight_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 3264 0 -1 710
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 3216 0 -1 690
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  pre_aadderRight_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 3198 0 1 480
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 3288 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  pre_aadderRight_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 3198 0 -1 470
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  pre_aadderRight_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 3150 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  pre_aadderRight_acelem_acx0
timestamp 1734143631
transform 1 0 4014 0 1 960
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay1_acx0
timestamp 1734143631
transform 1 0 4104 0 -1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay1_acx1
timestamp 1734143631
transform 1 0 4152 0 -1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay1_acx2
timestamp 1734143631
transform 1 0 4170 0 1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay1_acx3
timestamp 1734143631
transform 1 0 4110 0 1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay1_acx4
timestamp 1734143631
transform 1 0 4050 0 -1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay1_acx5
timestamp 1734143631
transform 1 0 4128 0 -1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay1_acx6
timestamp 1734143631
transform 1 0 4140 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay1_acx7
timestamp 1734143631
transform 1 0 4188 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay2_acx0
timestamp 1734143631
transform 1 0 4188 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay2_acx1
timestamp 1734143631
transform 1 0 4152 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay2_acx2
timestamp 1734143631
transform 1 0 4098 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay2_acx3
timestamp 1734143631
transform 1 0 4104 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay2_acx4
timestamp 1734143631
transform 1 0 4050 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay2_acx5
timestamp 1734143631
transform 1 0 4062 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay2_acx6
timestamp 1734143631
transform 1 0 3990 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_aadderRight_adelay2_acx7
timestamp 1734143631
transform 1 0 3924 0 -1 470
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_ainv__l1
timestamp 1734143760
transform 1 0 4134 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_ainv__l2
timestamp 1734143760
transform 1 0 3930 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_ainv__r
timestamp 1734143760
transform 1 0 3894 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al1_50_6
timestamp 1734143796
transform 1 0 2916 0 -1 1890
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al1_51_6
timestamp 1734143796
transform 1 0 2772 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al1_52_6
timestamp 1734143796
transform 1 0 2610 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al1_53_6
timestamp 1734143796
transform 1 0 2610 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al1_54_6
timestamp 1734143796
transform 1 0 2700 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al1_55_6
timestamp 1734143796
transform 1 0 2988 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al1_56_6
timestamp 1734143796
transform 1 0 3258 0 1 1200
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al1_57_6
timestamp 1734143796
transform 1 0 3180 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al2_50_6
timestamp 1734143796
transform 1 0 2718 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al2_51_6
timestamp 1734143796
transform 1 0 2442 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al2_52_6
timestamp 1734143796
transform 1 0 2424 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al2_53_6
timestamp 1734143796
transform 1 0 2436 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al2_54_6
timestamp 1734143796
transform 1 0 2814 0 1 210
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al2_55_6
timestamp 1734143796
transform 1 0 2868 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al2_56_6
timestamp 1734143796
transform 1 0 3306 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_aadderRight_al2_57_6
timestamp 1734143796
transform 1 0 3294 0 1 480
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  pre_aadderRight_anor
timestamp 1734143909
transform 1 0 3930 0 1 710
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  pre_aadderRight_aor__l1
timestamp 1734143975
transform 1 0 4038 0 -1 1180
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  pre_aadderRight_aor__l2
timestamp 1734143975
transform 1 0 3972 0 -1 1180
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  pre_aadderRight_apulseG_aand
timestamp 1734143631
transform 1 0 3480 0 1 950
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai
timestamp 1734143760
transform 1 0 3732 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai1
timestamp 1734143760
transform 1 0 3546 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai2
timestamp 1734143760
transform 1 0 3582 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai3
timestamp 1734143760
transform 1 0 3630 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai4
timestamp 1734143760
transform 1 0 3678 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai5
timestamp 1734143760
transform 1 0 3726 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai6
timestamp 1734143760
transform 1 0 3642 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai7
timestamp 1734143760
transform 1 0 3558 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai8
timestamp 1734143760
transform 1 0 3408 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_aadderRight_apulseG_ai9
timestamp 1734143760
transform 1 0 3480 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  pre_aadderRight_apulseG_anor
timestamp 1734143909
transform 1 0 3732 0 1 950
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  pre_aadderRight_atoGND
timestamp 1734144021
transform 1 0 2814 0 -1 2110
box 0 0 30 50
use _0_0cell_0_0g0n1n2naa_012aax0  pre_acp1_acelem_acx0
timestamp 1734143631
transform 1 0 2760 0 1 2140
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  pre_acp1_adelay1_acx0
timestamp 1734143631
transform 1 0 2886 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_acp1_adelay1_acx1
timestamp 1734143631
transform 1 0 3108 0 1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_acp1_adelay1_acx2
timestamp 1734143631
transform 1 0 3204 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_acp1_adelay1_acx3
timestamp 1734143631
transform 1 0 3300 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_acp1_adelay1_acx4
timestamp 1734143631
transform 1 0 3510 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_acp1_adelay1_acx5
timestamp 1734143631
transform 1 0 3552 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_acp1_adelay1_acx6
timestamp 1734143631
transform 1 0 3600 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_acp1_adelay1_acx7
timestamp 1734143631
transform 1 0 3696 0 1 1420
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  pre_acp1_ainv__1
timestamp 1734143760
transform 1 0 2844 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_ainv__2
timestamp 1734143760
transform 1 0 3252 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_ainv__3
timestamp 1734143760
transform 1 0 2046 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  pre_acp1_al_50_6
timestamp 1734143796
transform 1 0 2208 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  pre_acp1_anor__2
timestamp 1734143909
transform 1 0 2952 0 -1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  pre_acp1_anor__3
timestamp 1734143909
transform 1 0 3438 0 -1 1420
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  pre_acp1_aor__1
timestamp 1734143975
transform 1 0 2310 0 1 2140
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  pre_acp1_apulseG_aand
timestamp 1734143631
transform 1 0 2202 0 1 2130
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai
timestamp 1734143760
transform 1 0 2232 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai1
timestamp 1734143760
transform 1 0 2142 0 -1 2360
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai2
timestamp 1734143760
transform 1 0 2166 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai3
timestamp 1734143760
transform 1 0 2130 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai4
timestamp 1734143760
transform 1 0 2088 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai5
timestamp 1734143760
transform 1 0 1998 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai6
timestamp 1734143760
transform 1 0 2046 0 1 2140
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai7
timestamp 1734143760
transform 1 0 2082 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai8
timestamp 1734143760
transform 1 0 2124 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_acp1_apulseG_ai9
timestamp 1734143760
transform 1 0 2166 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  pre_acp1_apulseG_anor
timestamp 1734143909
transform 1 0 2178 0 -1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  pre_amerge_aand1
timestamp 1734143631
transform 1 0 3786 0 -1 710
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  pre_amerge_aand2
timestamp 1734143631
transform 1 0 3600 0 -1 710
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  pre_amerge_acelem1_acx0
timestamp 1734143631
transform 1 0 3912 0 1 480
box 6 10 65 70
use _0_0cell_0_0g0n1n2naa_012aax0  pre_amerge_acelem2_acx0
timestamp 1734143631
transform 1 0 3762 0 1 480
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay1_acx0
timestamp 1734143631
transform 1 0 3666 0 -1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay1_acx1
timestamp 1734143631
transform 1 0 3618 0 -1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay1_acx2
timestamp 1734143631
transform 1 0 3660 0 1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay1_acx3
timestamp 1734143631
transform 1 0 3666 0 -1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay1_acx4
timestamp 1734143631
transform 1 0 3798 0 1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay1_acx5
timestamp 1734143631
transform 1 0 3810 0 -1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay1_acx6
timestamp 1734143631
transform 1 0 3696 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay1_acx7
timestamp 1734143631
transform 1 0 3726 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay2_acx0
timestamp 1734143631
transform 1 0 3624 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay2_acx1
timestamp 1734143631
transform 1 0 3552 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay2_acx2
timestamp 1734143631
transform 1 0 3552 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay2_acx3
timestamp 1734143631
transform 1 0 3594 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay2_acx4
timestamp 1734143631
transform 1 0 3654 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay2_acx5
timestamp 1734143631
transform 1 0 3720 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay2_acx6
timestamp 1734143631
transform 1 0 3720 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay2_acx7
timestamp 1734143631
transform 1 0 3660 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay3_acx0
timestamp 1734143631
transform 1 0 3594 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay3_acx1
timestamp 1734143631
transform 1 0 3528 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay3_acx2
timestamp 1734143631
transform 1 0 3462 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay3_acx3
timestamp 1734143631
transform 1 0 3402 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay3_acx4
timestamp 1734143631
transform 1 0 3342 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay3_acx5
timestamp 1734143631
transform 1 0 3276 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay3_acx6
timestamp 1734143631
transform 1 0 3204 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_amerge_adelay3_acx7
timestamp 1734143631
transform 1 0 3000 0 1 200
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv1__Cd
timestamp 1734143760
transform 1 0 3504 0 -1 700
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Cf
timestamp 1734143760
transform 1 0 3678 0 -1 700
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Ct
timestamp 1734143760
transform 1 0 3870 0 -1 700
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__L1
timestamp 1734143760
transform 1 0 3864 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__L2
timestamp 1734143760
transform 1 0 3780 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Ra
timestamp 1734143760
transform 1 0 3642 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Rd1
timestamp 1734143760
transform 1 0 2238 0 -1 1410
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Rd2
timestamp 1734143760
transform 1 0 2214 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Rd3
timestamp 1734143760
transform 1 0 2262 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Rd4
timestamp 1734143760
transform 1 0 2286 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Rd5
timestamp 1734143760
transform 1 0 2340 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Rd6
timestamp 1734143760
transform 1 0 2382 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Rd7
timestamp 1734143760
transform 1 0 2544 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_ainv__Rd8
timestamp 1734143760
transform 1 0 2778 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  pre_amerge_al_50_6
timestamp 1734143796
transform 1 0 2298 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_amerge_al_51_6
timestamp 1734143796
transform 1 0 2280 0 1 1200
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_amerge_al_52_6
timestamp 1734143796
transform 1 0 2286 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_amerge_al_53_6
timestamp 1734143796
transform 1 0 2340 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_amerge_al_54_6
timestamp 1734143796
transform 1 0 2526 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_amerge_al_55_6
timestamp 1734143796
transform 1 0 2634 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_amerge_al_56_6
timestamp 1734143796
transform 1 0 2946 0 -1 460
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_amerge_al_57_6
timestamp 1734143796
transform 1 0 3072 0 1 210
box 0 0 96 80
use _0_0std_0_0cells_0_0MUX2X1  pre_amerge_amux_50_6
timestamp 1734143875
transform 1 0 2736 0 -1 1420
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  pre_amerge_amux_51_6
timestamp 1734143875
transform 1 0 2412 0 1 1190
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  pre_amerge_amux_52_6
timestamp 1734143875
transform 1 0 2304 0 1 950
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  pre_amerge_amux_53_6
timestamp 1734143875
transform 1 0 2424 0 1 710
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  pre_amerge_amux_54_6
timestamp 1734143875
transform 1 0 2658 0 -1 470
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  pre_amerge_amux_55_6
timestamp 1734143875
transform 1 0 2838 0 1 470
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  pre_amerge_amux_56_6
timestamp 1734143875
transform 1 0 3108 0 -1 710
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  pre_amerge_amux_57_6
timestamp 1734143875
transform 1 0 3096 0 1 470
box 0 0 90 90
use _0_0std_0_0cells_0_0NOR2X1  pre_amerge_anor__Ra
timestamp 1734143909
transform 1 0 3078 0 -1 470
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  pre_amerge_aor
timestamp 1734143975
transform 1 0 3768 0 1 720
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  pre_amerge_aor__Cf
timestamp 1734143975
transform 1 0 3690 0 1 480
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  pre_amerge_aor__Ct
timestamp 1734143975
transform 1 0 3918 0 -1 700
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  pre_amerge_aor__L1
timestamp 1734143975
transform 1 0 3846 0 1 480
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  pre_amerge_aor__L2
timestamp 1734143975
transform 1 0 3780 0 -1 460
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  pre_amerge_apulseG_aand
timestamp 1734143631
transform 1 0 3396 0 1 470
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai
timestamp 1734143760
transform 1 0 3492 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai1
timestamp 1734143760
transform 1 0 3468 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai2
timestamp 1734143760
transform 1 0 3510 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai3
timestamp 1734143760
transform 1 0 3552 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai4
timestamp 1734143760
transform 1 0 3594 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai5
timestamp 1734143760
transform 1 0 3540 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai6
timestamp 1734143760
transform 1 0 3492 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai7
timestamp 1734143760
transform 1 0 3450 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai8
timestamp 1734143760
transform 1 0 3408 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_amerge_apulseG_ai9
timestamp 1734143760
transform 1 0 3372 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  pre_amerge_apulseG_anor
timestamp 1734143909
transform 1 0 3444 0 -1 710
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  pre_asplit_aand1
timestamp 1734143631
transform 1 0 4074 0 -1 1420
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  pre_asplit_aand2
timestamp 1734143631
transform 1 0 3888 0 -1 1420
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  pre_asplit_acelem_acx0
timestamp 1734143631
transform 1 0 3768 0 -1 1650
box 6 10 65 70
use _0_0std_0_0cells_0_0LATCH  pre_asplit_acontrolLatch
timestamp 1734143796
transform 1 0 3504 0 -1 1410
box 0 0 96 80
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay1_acx0
timestamp 1734143631
transform 1 0 3828 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay1_acx1
timestamp 1734143631
transform 1 0 3930 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay1_acx2
timestamp 1734143631
transform 1 0 4032 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay1_acx3
timestamp 1734143631
transform 1 0 4038 0 1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay1_acx4
timestamp 1734143631
transform 1 0 3918 0 1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay1_acx5
timestamp 1734143631
transform 1 0 3954 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay1_acx6
timestamp 1734143631
transform 1 0 3996 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay1_acx7
timestamp 1734143631
transform 1 0 4044 0 1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay2_acx0
timestamp 1734143631
transform 1 0 4116 0 1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay2_acx1
timestamp 1734143631
transform 1 0 4074 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay2_acx2
timestamp 1734143631
transform 1 0 4020 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay2_acx3
timestamp 1734143631
transform 1 0 3966 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay2_acx4
timestamp 1734143631
transform 1 0 3906 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay2_acx5
timestamp 1734143631
transform 1 0 3834 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay2_acx6
timestamp 1734143631
transform 1 0 3984 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  pre_asplit_adelay2_acx7
timestamp 1734143631
transform 1 0 3990 0 -1 1420
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  pre_asplit_ainv__c
timestamp 1734143760
transform 1 0 3648 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_ainv__ctr
timestamp 1734143760
transform 1 0 3714 0 -1 1410
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_ainv__l
timestamp 1734143760
transform 1 0 3522 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_ainv__r
timestamp 1734143760
transform 1 0 3768 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  pre_asplit_al_50_6
timestamp 1734143796
transform 1 0 2976 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_asplit_al_51_6
timestamp 1734143796
transform 1 0 2844 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_asplit_al_52_6
timestamp 1734143796
transform 1 0 2934 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_asplit_al_53_6
timestamp 1734143796
transform 1 0 2604 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_asplit_al_54_6
timestamp 1734143796
transform 1 0 2940 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_asplit_al_55_6
timestamp 1734143796
transform 1 0 3096 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_asplit_al_56_6
timestamp 1734143796
transform 1 0 3288 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  pre_asplit_al_57_6
timestamp 1734143796
transform 1 0 3192 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  pre_asplit_anor__R
timestamp 1734143909
transform 1 0 3756 0 -1 1420
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  pre_asplit_aor1
timestamp 1734143975
transform 1 0 3570 0 1 1670
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  pre_asplit_aor2
timestamp 1734143975
transform 1 0 3696 0 -1 1650
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  pre_asplit_aor
timestamp 1734143975
transform 1 0 3738 0 1 1200
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  pre_asplit_apulseG_aand
timestamp 1734143631
transform 1 0 3486 0 1 1660
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai1
timestamp 1734143760
transform 1 0 3798 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai3
timestamp 1734143760
transform 1 0 3876 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai
timestamp 1734143760
transform 1 0 3708 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai2
timestamp 1734143760
transform 1 0 3834 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai4
timestamp 1734143760
transform 1 0 3882 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai5
timestamp 1734143760
transform 1 0 3930 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai6
timestamp 1734143760
transform 1 0 3984 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai7
timestamp 1734143760
transform 1 0 3786 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai8
timestamp 1734143760
transform 1 0 3696 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  pre_asplit_apulseG_ai9
timestamp 1734143760
transform 1 0 3648 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  pre_asplit_apulseG_anor
timestamp 1734143909
transform 1 0 3750 0 -1 1900
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  pre_asrc65_anor
timestamp 1734143909
transform 1 0 3882 0 1 1190
box 0 0 42 80
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc65_aset0
timestamp 1734144001
transform 1 0 3090 0 -1 1640
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc65_aset1
timestamp 1734144001
transform 1 0 2988 0 1 1210
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc65_aset2
timestamp 1734144001
transform 1 0 2982 0 -1 1170
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc65_aset3
timestamp 1734144001
transform 1 0 3078 0 -1 930
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc65_aset4
timestamp 1734144001
transform 1 0 3000 0 -1 690
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc65_aset5
timestamp 1734144001
transform 1 0 3066 0 -1 1400
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  pre_asrc65_aset6
timestamp 1734144021
transform 1 0 3378 0 -1 1400
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc65_aset7
timestamp 1734144001
transform 1 0 3444 0 1 970
box 0 0 30 50
use _0_0std_0_0cells_0_0NOR2X1  pre_asrc97_anor
timestamp 1734143909
transform 1 0 3786 0 -1 1190
box 0 0 42 80
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc97_asetGND0
timestamp 1734144001
transform 1 0 2766 0 -1 2110
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc97_asetGND1
timestamp 1734144001
transform 1 0 2562 0 -1 1640
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc97_asetGND2
timestamp 1734144001
transform 1 0 2550 0 -1 1400
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc97_asetGND3
timestamp 1734144001
transform 1 0 2400 0 1 970
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc97_asetGND4
timestamp 1734144001
transform 1 0 2934 0 1 220
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  pre_asrc97_asetGND5
timestamp 1734144021
transform 1 0 2964 0 -1 690
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  pre_asrc97_asetGND6
timestamp 1734144021
transform 1 0 3432 0 1 730
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  pre_asrc97_asetGND7
timestamp 1734144001
transform 1 0 3330 0 -1 450
box 0 0 30 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_aadd__key_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 1968 0 1 1430
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 2064 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_aadd__key_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 1872 0 1 1420
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 1812 0 -1 1400
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_aadd__key_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 2028 0 -1 1410
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 1914 0 1 1210
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_aadd__key_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 1974 0 1 1190
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 1974 0 -1 1400
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_aadd__key_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 1956 0 -1 1180
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 2034 0 1 970
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_aadd__key_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 1944 0 1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 1902 0 1 970
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_aadd__key_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 2076 0 1 960
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 2118 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_aadd__key_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 2022 0 -1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 1974 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_aadd__key_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 2142 0 1 720
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 2094 0 1 730
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_aadd__key_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 2136 0 -1 710
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 1956 0 -1 690
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_aadd__key_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 1980 0 -1 700
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 2076 0 1 490
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_aadd__key_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 1998 0 1 470
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 1932 0 1 490
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_aadd__key_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 2208 0 1 480
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 2274 0 1 490
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_aadd__key_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 2160 0 -1 470
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 2016 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_aadd__key_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 2316 0 -1 700
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 2400 0 1 490
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_aadd__key_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 2310 0 1 470
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_aadd__key_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 2274 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  shft_aadd__key_acelem_acx0
timestamp 1734143631
transform 1 0 2610 0 1 480
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay1_acx0
timestamp 1734143631
transform 1 0 2334 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay1_acx1
timestamp 1734143631
transform 1 0 2286 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay1_acx2
timestamp 1734143631
transform 1 0 2220 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay1_acx3
timestamp 1734143631
transform 1 0 2154 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay1_acx4
timestamp 1734143631
transform 1 0 1788 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay1_acx5
timestamp 1734143631
transform 1 0 1746 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay1_acx6
timestamp 1734143631
transform 1 0 1704 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay1_acx7
timestamp 1734143631
transform 1 0 1170 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay2_acx0
timestamp 1734143631
transform 1 0 1056 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay2_acx1
timestamp 1734143631
transform 1 0 732 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay2_acx2
timestamp 1734143631
transform 1 0 690 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay2_acx3
timestamp 1734143631
transform 1 0 654 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay2_acx4
timestamp 1734143631
transform 1 0 618 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay2_acx5
timestamp 1734143631
transform 1 0 576 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay2_acx6
timestamp 1734143631
transform 1 0 534 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_aadd__key_adelay2_acx7
timestamp 1734143631
transform 1 0 486 0 1 200
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_ainv__l1
timestamp 1734143760
transform 1 0 2658 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_ainv__l2
timestamp 1734143760
transform 1 0 2586 0 -1 700
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_ainv__r
timestamp 1734143760
transform 1 0 2088 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al1_50_6
timestamp 1734143796
transform 1 0 2124 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al1_51_6
timestamp 1734143796
transform 1 0 2082 0 1 1200
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al1_52_6
timestamp 1734143796
transform 1 0 2160 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al1_53_6
timestamp 1734143796
transform 1 0 2166 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al1_54_6
timestamp 1734143796
transform 1 0 2226 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al1_55_6
timestamp 1734143796
transform 1 0 2040 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al1_56_6
timestamp 1734143796
transform 1 0 2382 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al1_57_6
timestamp 1734143796
transform 1 0 2484 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al2_50_6
timestamp 1734143796
transform 1 0 2256 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al2_51_6
timestamp 1734143796
transform 1 0 2112 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al2_52_6
timestamp 1734143796
transform 1 0 2040 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al2_53_6
timestamp 1734143796
transform 1 0 2154 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al2_54_6
timestamp 1734143796
transform 1 0 1974 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al2_55_6
timestamp 1734143796
transform 1 0 1860 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al2_56_6
timestamp 1734143796
transform 1 0 2106 0 1 480
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_aadd__key_al2_57_6
timestamp 1734143796
transform 1 0 2214 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  shft_aadd__key_anor
timestamp 1734143909
transform 1 0 1956 0 1 470
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  shft_aadd__key_aor__l1
timestamp 1734143975
transform 1 0 2604 0 1 210
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_aadd__key_aor__l2
timestamp 1734143975
transform 1 0 2622 0 -1 700
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  shft_aadd__key_apulseG_aand
timestamp 1734143631
transform 1 0 2454 0 1 470
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai1
timestamp 1734143760
transform 1 0 2532 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai2
timestamp 1734143760
transform 1 0 2592 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai
timestamp 1734143760
transform 1 0 2406 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai3
timestamp 1734143760
transform 1 0 2574 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai4
timestamp 1734143760
transform 1 0 2544 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai5
timestamp 1734143760
transform 1 0 2514 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai6
timestamp 1734143760
transform 1 0 2478 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai7
timestamp 1734143760
transform 1 0 2346 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai8
timestamp 1734143760
transform 1 0 2394 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_aadd__key_apulseG_ai9
timestamp 1734143760
transform 1 0 2436 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  shft_aadd__key_apulseG_anor
timestamp 1734143909
transform 1 0 2466 0 -1 470
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  shft_aadd__key_atoGND
timestamp 1734144021
transform 1 0 1812 0 -1 1640
box 0 0 30 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_acomp_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 1848 0 -1 1890
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 1806 0 1 1680
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_acomp_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 1848 0 1 1660
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 1944 0 1 1680
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_acomp_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 1728 0 -1 1650
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 1728 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_acomp_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 1656 0 1 1420
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 1632 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_acomp_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 1638 0 1 1200
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 1794 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_acomp_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 1734 0 1 1190
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 1848 0 1 1210
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_acomp_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 1662 0 1 960
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 1728 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_acomp_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 1752 0 1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 1854 0 1 970
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_acomp_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 1632 0 -1 940
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 1614 0 -1 690
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_acomp_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 1632 0 1 710
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 1578 0 1 730
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_acomp_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 1518 0 1 480
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 1518 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_acomp_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 1572 0 -1 470
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 1530 0 1 220
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_acomp_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 1458 0 1 210
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 1122 0 1 220
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_acomp_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 1380 0 1 200
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 1344 0 1 220
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_acomp_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 918 0 1 210
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 1002 0 1 220
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_acomp_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 822 0 1 200
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_acomp_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 684 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  shft_acomp_acelem_acx0
timestamp 1734143631
transform 1 0 348 0 1 1670
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay1_acx0
timestamp 1734143631
transform 1 0 408 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay1_acx1
timestamp 1734143631
transform 1 0 372 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay1_acx2
timestamp 1734143631
transform 1 0 318 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay1_acx3
timestamp 1734143631
transform 1 0 240 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay1_acx4
timestamp 1734143631
transform 1 0 216 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay1_acx5
timestamp 1734143631
transform 1 0 174 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay1_acx6
timestamp 1734143631
transform 1 0 228 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay1_acx7
timestamp 1734143631
transform 1 0 252 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay2_acx0
timestamp 1734143631
transform 1 0 204 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay2_acx1
timestamp 1734143631
transform 1 0 168 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay2_acx2
timestamp 1734143631
transform 1 0 132 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay2_acx3
timestamp 1734143631
transform 1 0 96 0 -1 3090
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay2_acx4
timestamp 1734143631
transform 1 0 96 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay2_acx5
timestamp 1734143631
transform 1 0 132 0 1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay2_acx6
timestamp 1734143631
transform 1 0 144 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay2_acx7
timestamp 1734143631
transform 1 0 96 0 -1 2850
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay3_acx0
timestamp 1734143631
transform 1 0 96 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay3_acx1
timestamp 1734143631
transform 1 0 96 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay3_acx2
timestamp 1734143631
transform 1 0 96 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay3_acx3
timestamp 1734143631
transform 1 0 132 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay3_acx4
timestamp 1734143631
transform 1 0 132 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay3_acx5
timestamp 1734143631
transform 1 0 96 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay3_acx6
timestamp 1734143631
transform 1 0 96 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomp_adelay3_acx7
timestamp 1734143631
transform 1 0 138 0 1 2130
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  shft_acomp_ainv__l1
timestamp 1734143760
transform 1 0 240 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_ainv__l2
timestamp 1734143760
transform 1 0 294 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_ainv__r
timestamp 1734143760
transform 1 0 258 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al1_50_6
timestamp 1734143796
transform 1 0 1692 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al1_51_6
timestamp 1734143796
transform 1 0 1758 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al1_52_6
timestamp 1734143796
transform 1 0 1506 0 1 1200
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al1_53_6
timestamp 1734143796
transform 1 0 1536 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al1_54_6
timestamp 1734143796
transform 1 0 1734 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al1_55_6
timestamp 1734143796
transform 1 0 1638 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al1_56_6
timestamp 1734143796
transform 1 0 1230 0 1 210
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al1_57_6
timestamp 1734143796
transform 1 0 840 0 -1 460
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al2_50_6
timestamp 1734143796
transform 1 0 1746 0 -1 1890
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al2_51_6
timestamp 1734143796
transform 1 0 1602 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al2_52_6
timestamp 1734143796
transform 1 0 1548 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al2_53_6
timestamp 1734143796
transform 1 0 1620 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al2_54_6
timestamp 1734143796
transform 1 0 1500 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al2_55_6
timestamp 1734143796
transform 1 0 1674 0 -1 460
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al2_56_6
timestamp 1734143796
transform 1 0 1566 0 1 210
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_acomp_al2_57_6
timestamp 1734143796
transform 1 0 726 0 -1 460
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  shft_acomp_anor
timestamp 1734143909
transform 1 0 204 0 -1 1900
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  shft_acomp_aor__l1
timestamp 1734143975
transform 1 0 282 0 1 1670
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_acomp_aor__l2
timestamp 1734143975
transform 1 0 330 0 -1 1890
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  shft_acomp_apulseG_aand
timestamp 1734143631
transform 1 0 720 0 1 470
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai
timestamp 1734143760
transform 1 0 642 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai1
timestamp 1734143760
transform 1 0 660 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai2
timestamp 1734143760
transform 1 0 600 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai3
timestamp 1734143760
transform 1 0 546 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai4
timestamp 1734143760
transform 1 0 378 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai5
timestamp 1734143760
transform 1 0 432 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai6
timestamp 1734143760
transform 1 0 486 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai7
timestamp 1734143760
transform 1 0 540 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai8
timestamp 1734143760
transform 1 0 588 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomp_apulseG_ai9
timestamp 1734143760
transform 1 0 636 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  shft_acomp_apulseG_anor
timestamp 1734143909
transform 1 0 612 0 -1 950
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  shft_acomp_atoGND
timestamp 1734144021
transform 1 0 1824 0 1 1920
box 0 0 30 50
use _0_0cell_0_0g0n1n2naa_012aax0  shft_acomps_acelem_acx0
timestamp 1734143631
transform 1 0 186 0 1 1910
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  shft_acomps_adelay1_acx0
timestamp 1734143631
transform 1 0 294 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomps_adelay1_acx1
timestamp 1734143631
transform 1 0 318 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomps_adelay1_acx2
timestamp 1734143631
transform 1 0 252 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomps_adelay1_acx3
timestamp 1734143631
transform 1 0 192 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomps_adelay1_acx4
timestamp 1734143631
transform 1 0 132 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomps_adelay1_acx5
timestamp 1734143631
transform 1 0 96 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomps_adelay1_acx6
timestamp 1734143631
transform 1 0 96 0 1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_acomps_adelay1_acx7
timestamp 1734143631
transform 1 0 132 0 1 1900
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  shft_acomps_ainv__1
timestamp 1734143760
transform 1 0 162 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_ainv__2
timestamp 1734143760
transform 1 0 252 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_ainv__3
timestamp 1734143760
transform 1 0 168 0 -1 2120
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  shft_acomps_al_50_6
timestamp 1734143796
transform 1 0 600 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  shft_acomps_anor__2
timestamp 1734143909
transform 1 0 186 0 1 1660
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  shft_acomps_anor__3
timestamp 1734143909
transform 1 0 348 0 -1 2130
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  shft_acomps_aor__1
timestamp 1734143975
transform 1 0 198 0 -1 2120
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  shft_acomps_apulseG_aand
timestamp 1734143631
transform 1 0 462 0 -1 710
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai
timestamp 1734143760
transform 1 0 282 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai1
timestamp 1734143760
transform 1 0 510 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai2
timestamp 1734143760
transform 1 0 540 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai3
timestamp 1734143760
transform 1 0 480 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai4
timestamp 1734143760
transform 1 0 426 0 -1 700
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai5
timestamp 1734143760
transform 1 0 390 0 -1 700
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai6
timestamp 1734143760
transform 1 0 354 0 -1 700
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai7
timestamp 1734143760
transform 1 0 360 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai8
timestamp 1734143760
transform 1 0 402 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_acomps_apulseG_ai9
timestamp 1734143760
transform 1 0 444 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  shft_acomps_apulseG_anor
timestamp 1734143909
transform 1 0 324 0 1 950
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  shft_amerge_aand1
timestamp 1734143631
transform 1 0 414 0 -1 1420
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  shft_amerge_aand2
timestamp 1734143631
transform 1 0 558 0 -1 1420
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  shft_amerge_acelem1_acx0
timestamp 1734143631
transform 1 0 318 0 -1 1410
box 6 10 65 70
use _0_0cell_0_0g0n1n2naa_012aax0  shft_amerge_acelem2_acx0
timestamp 1734143631
transform 1 0 330 0 1 1200
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay1_acx0
timestamp 1734143631
transform 1 0 96 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay1_acx1
timestamp 1734143631
transform 1 0 96 0 1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay1_acx2
timestamp 1734143631
transform 1 0 96 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay1_acx3
timestamp 1734143631
transform 1 0 132 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay1_acx4
timestamp 1734143631
transform 1 0 102 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay1_acx5
timestamp 1734143631
transform 1 0 138 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay1_acx6
timestamp 1734143631
transform 1 0 168 0 -1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay1_acx7
timestamp 1734143631
transform 1 0 180 0 1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay2_acx0
timestamp 1734143631
transform 1 0 384 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay2_acx1
timestamp 1734143631
transform 1 0 312 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay2_acx2
timestamp 1734143631
transform 1 0 252 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay2_acx3
timestamp 1734143631
transform 1 0 192 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay2_acx4
timestamp 1734143631
transform 1 0 180 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay2_acx5
timestamp 1734143631
transform 1 0 228 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay2_acx6
timestamp 1734143631
transform 1 0 276 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay2_acx7
timestamp 1734143631
transform 1 0 186 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay3_acx0
timestamp 1734143631
transform 1 0 132 0 -1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay3_acx1
timestamp 1734143631
transform 1 0 132 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay3_acx2
timestamp 1734143631
transform 1 0 168 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay3_acx3
timestamp 1734143631
transform 1 0 204 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay3_acx4
timestamp 1734143631
transform 1 0 246 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay3_acx5
timestamp 1734143631
transform 1 0 282 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay3_acx6
timestamp 1734143631
transform 1 0 318 0 1 2610
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_amerge_adelay3_acx7
timestamp 1734143631
transform 1 0 294 0 -1 2610
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv1__Cd
timestamp 1734143760
transform 1 0 648 0 -1 1410
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Cf
timestamp 1734143760
transform 1 0 498 0 -1 1410
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Ct
timestamp 1734143760
transform 1 0 414 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__L1
timestamp 1734143760
transform 1 0 372 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__L2
timestamp 1734143760
transform 1 0 318 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Ra
timestamp 1734143760
transform 1 0 336 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Rd1
timestamp 1734143760
transform 1 0 1290 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Rd2
timestamp 1734143760
transform 1 0 1416 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Rd3
timestamp 1734143760
transform 1 0 1260 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Rd4
timestamp 1734143760
transform 1 0 1188 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Rd5
timestamp 1734143760
transform 1 0 948 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Rd6
timestamp 1734143760
transform 1 0 918 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Rd7
timestamp 1734143760
transform 1 0 762 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_ainv__Rd8
timestamp 1734143760
transform 1 0 618 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  shft_amerge_al_50_6
timestamp 1734143796
transform 1 0 1302 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_amerge_al_51_6
timestamp 1734143796
transform 1 0 1470 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_amerge_al_52_6
timestamp 1734143796
transform 1 0 1200 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_amerge_al_53_6
timestamp 1734143796
transform 1 0 1086 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_amerge_al_54_6
timestamp 1734143796
transform 1 0 984 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_amerge_al_55_6
timestamp 1734143796
transform 1 0 822 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_amerge_al_56_6
timestamp 1734143796
transform 1 0 738 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_amerge_al_57_6
timestamp 1734143796
transform 1 0 600 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0MUX2X1  shft_amerge_amux_50_6
timestamp 1734143875
transform 1 0 1278 0 -1 1420
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  shft_amerge_amux_51_6
timestamp 1734143875
transform 1 0 1170 0 1 1190
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  shft_amerge_amux_52_6
timestamp 1734143875
transform 1 0 1158 0 1 950
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  shft_amerge_amux_53_6
timestamp 1734143875
transform 1 0 1140 0 -1 710
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  shft_amerge_amux_54_6
timestamp 1734143875
transform 1 0 1134 0 1 470
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  shft_amerge_amux_55_6
timestamp 1734143875
transform 1 0 804 0 1 470
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  shft_amerge_amux_56_6
timestamp 1734143875
transform 1 0 738 0 -1 710
box 0 0 90 90
use _0_0std_0_0cells_0_0MUX2X1  shft_amerge_amux_57_6
timestamp 1734143875
transform 1 0 648 0 1 950
box 0 0 90 90
use _0_0std_0_0cells_0_0NOR2X1  shft_amerge_anor__Ra
timestamp 1734143909
transform 1 0 432 0 -1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  shft_amerge_aor
timestamp 1734143975
transform 1 0 318 0 1 1430
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_amerge_aor__Cf
timestamp 1734143975
transform 1 0 444 0 1 1200
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_amerge_aor__Ct
timestamp 1734143975
transform 1 0 252 0 -1 1410
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_amerge_aor__L1
timestamp 1734143975
transform 1 0 264 0 1 960
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_amerge_aor__L2
timestamp 1734143975
transform 1 0 288 0 -1 700
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  shft_amerge_apulseG_aand
timestamp 1734143631
transform 1 0 426 0 1 1660
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai1
timestamp 1734143760
transform 1 0 456 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai2
timestamp 1734143760
transform 1 0 432 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai3
timestamp 1734143760
transform 1 0 480 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai4
timestamp 1734143760
transform 1 0 528 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai
timestamp 1734143760
transform 1 0 384 0 1 1910
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai5
timestamp 1734143760
transform 1 0 510 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai6
timestamp 1734143760
transform 1 0 564 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai7
timestamp 1734143760
transform 1 0 618 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai8
timestamp 1734143760
transform 1 0 588 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_amerge_apulseG_ai9
timestamp 1734143760
transform 1 0 492 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  shft_amerge_apulseG_anor
timestamp 1734143909
transform 1 0 396 0 -1 1900
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  shft_asplit_aand1
timestamp 1734143631
transform 1 0 324 0 1 710
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  shft_asplit_aand2
timestamp 1734143631
transform 1 0 234 0 1 710
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  shft_asplit_acelem_acx0
timestamp 1734143631
transform 1 0 198 0 -1 1650
box 6 10 65 70
use _0_0std_0_0cells_0_0LATCH  shft_asplit_acontrolLatch
timestamp 1734143796
transform 1 0 384 0 1 720
box 0 0 96 80
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay1_acx0
timestamp 1734143631
transform 1 0 210 0 -1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay1_acx1
timestamp 1734143631
transform 1 0 102 0 1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay1_acx2
timestamp 1734143631
transform 1 0 96 0 -1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay1_acx3
timestamp 1734143631
transform 1 0 96 0 1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay1_acx4
timestamp 1734143631
transform 1 0 96 0 -1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay1_acx5
timestamp 1734143631
transform 1 0 96 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay1_acx6
timestamp 1734143631
transform 1 0 96 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay1_acx7
timestamp 1734143631
transform 1 0 132 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay2_acx0
timestamp 1734143631
transform 1 0 168 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay2_acx1
timestamp 1734143631
transform 1 0 132 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay2_acx2
timestamp 1734143631
transform 1 0 96 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay2_acx3
timestamp 1734143631
transform 1 0 96 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay2_acx4
timestamp 1734143631
transform 1 0 132 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay2_acx5
timestamp 1734143631
transform 1 0 186 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay2_acx6
timestamp 1734143631
transform 1 0 216 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asplit_adelay2_acx7
timestamp 1734143631
transform 1 0 234 0 -1 710
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  shft_asplit_ainv__c
timestamp 1734143760
transform 1 0 132 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_ainv__ctr
timestamp 1734143760
transform 1 0 204 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_ainv__l
timestamp 1734143760
transform 1 0 330 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_ainv__r
timestamp 1734143760
transform 1 0 168 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  shft_asplit_al_50_6
timestamp 1734143796
transform 1 0 1536 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asplit_al_51_6
timestamp 1734143796
transform 1 0 1212 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asplit_al_52_6
timestamp 1734143796
transform 1 0 1500 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asplit_al_53_6
timestamp 1734143796
transform 1 0 1458 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asplit_al_54_6
timestamp 1734143796
transform 1 0 1512 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asplit_al_55_6
timestamp 1734143796
transform 1 0 1410 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asplit_al_56_6
timestamp 1734143796
transform 1 0 936 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asplit_al_57_6
timestamp 1734143796
transform 1 0 834 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  shft_asplit_anor__R
timestamp 1734143909
transform 1 0 180 0 1 1420
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  shft_asplit_aor1
timestamp 1734143975
transform 1 0 270 0 -1 1650
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_asplit_aor2
timestamp 1734143975
transform 1 0 132 0 1 1670
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_asplit_aor
timestamp 1734143975
transform 1 0 228 0 1 1430
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  shft_asplit_apulseG_aand
timestamp 1734143631
transform 1 0 222 0 -1 1190
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai
timestamp 1734143760
transform 1 0 132 0 -1 1410
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai1
timestamp 1734143760
transform 1 0 192 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai2
timestamp 1734143760
transform 1 0 132 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai3
timestamp 1734143760
transform 1 0 162 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai4
timestamp 1734143760
transform 1 0 162 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai5
timestamp 1734143760
transform 1 0 132 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai6
timestamp 1734143760
transform 1 0 132 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai7
timestamp 1734143760
transform 1 0 174 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai8
timestamp 1734143760
transform 1 0 228 0 -1 940
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asplit_apulseG_ai9
timestamp 1734143760
transform 1 0 228 0 1 960
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  shft_asplit_apulseG_anor
timestamp 1734143909
transform 1 0 138 0 1 1190
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  shft_asrc1_anor
timestamp 1734143909
transform 1 0 276 0 1 1900
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  shft_asrc1_asetGND0
timestamp 1734144021
transform 1 0 1770 0 1 1920
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc1_asetGND1
timestamp 1734144001
transform 1 0 1644 0 1 1680
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc1_asetGND2
timestamp 1734144001
transform 1 0 1656 0 -1 1400
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  shft_asrc1_asetGND3
timestamp 1734144021
transform 1 0 1740 0 -1 1170
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  shft_asrc1_asetGND4
timestamp 1734144021
transform 1 0 1788 0 -1 930
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc1_asetGND5
timestamp 1734144001
transform 1 0 1806 0 -1 450
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc1_asetGND6
timestamp 1734144001
transform 1 0 1668 0 1 220
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc1_asetGND7
timestamp 1734144001
transform 1 0 774 0 1 220
box 0 0 30 50
use _0_0std_0_0cells_0_0NOR2X1  shft_asrc2_anor
timestamp 1734143909
transform 1 0 288 0 1 1190
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  shft_asrc2_asetGND0
timestamp 1734144021
transform 1 0 1542 0 -1 1640
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc2_asetGND1
timestamp 1734144001
transform 1 0 1506 0 -1 1400
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc2_asetGND2
timestamp 1734144001
transform 1 0 1476 0 1 970
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  shft_asrc2_asetGND3
timestamp 1734144021
transform 1 0 1410 0 1 730
box 0 0 30 50
use _0_0std_0_0cells_0_0TIELOX1  shft_asrc2_asetGND4
timestamp 1734144021
transform 1 0 1464 0 -1 450
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc2_asetGND5
timestamp 1734144001
transform 1 0 1008 0 -1 450
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc2_asetGND6
timestamp 1734144001
transform 1 0 780 0 -1 930
box 0 0 30 50
use _0_0std_0_0cells_0_0TIEHIX1  shft_asrc2_asetGND7
timestamp 1734144001
transform 1 0 462 0 -1 1170
box 0 0 30 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_asub_aadd_50_6_acx0
timestamp 1734143631
transform 1 0 1452 0 -1 1650
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_50_6_acx1
timestamp 1734143631
transform 1 0 1440 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_asub_aadd_50_6_acx2
timestamp 1734143631
transform 1 0 1464 0 1 1420
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_50_6_acx3
timestamp 1734143631
transform 1 0 1416 0 1 1440
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_asub_aadd_51_6_acx0
timestamp 1734143631
transform 1 0 1422 0 1 1200
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_51_6_acx1
timestamp 1734143631
transform 1 0 1446 0 -1 1170
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_asub_aadd_51_6_acx2
timestamp 1734143631
transform 1 0 1326 0 1 1190
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_51_6_acx3
timestamp 1734143631
transform 1 0 1284 0 1 1210
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_asub_aadd_52_6_acx0
timestamp 1734143631
transform 1 0 1386 0 1 960
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_52_6_acx1
timestamp 1734143631
transform 1 0 1326 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_asub_aadd_52_6_acx2
timestamp 1734143631
transform 1 0 1392 0 -1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_52_6_acx3
timestamp 1734143631
transform 1 0 1260 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_asub_aadd_53_6_acx0
timestamp 1734143631
transform 1 0 1344 0 -1 700
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_53_6_acx1
timestamp 1734143631
transform 1 0 1344 0 1 490
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_asub_aadd_53_6_acx2
timestamp 1734143631
transform 1 0 1266 0 -1 710
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_53_6_acx3
timestamp 1734143631
transform 1 0 1236 0 -1 690
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_asub_aadd_54_6_acx0
timestamp 1734143631
transform 1 0 1254 0 1 480
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_54_6_acx1
timestamp 1734143631
transform 1 0 1158 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_asub_aadd_54_6_acx2
timestamp 1734143631
transform 1 0 1248 0 -1 470
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_54_6_acx3
timestamp 1734143631
transform 1 0 1206 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_asub_aadd_55_6_acx0
timestamp 1734143631
transform 1 0 1044 0 1 480
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_55_6_acx1
timestamp 1734143631
transform 1 0 708 0 -1 690
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_asub_aadd_55_6_acx2
timestamp 1734143631
transform 1 0 1062 0 -1 470
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_55_6_acx3
timestamp 1734143631
transform 1 0 960 0 -1 450
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_asub_aadd_56_6_acx0
timestamp 1734143631
transform 1 0 666 0 1 720
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_56_6_acx1
timestamp 1734143631
transform 1 0 570 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_asub_aadd_56_6_acx2
timestamp 1734143631
transform 1 0 726 0 1 710
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_56_6_acx3
timestamp 1734143631
transform 1 0 798 0 1 730
box 6 10 21 50
use _0_0cell_0_0g0n1na2no0n1noa_01o2a01aox0  shft_asub_aadd_57_6_acx0
timestamp 1734143631
transform 1 0 468 0 1 960
box 6 10 57 70
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_57_6_acx1
timestamp 1734143631
transform 1 0 432 0 -1 930
box 6 10 21 50
use _0_0cell_0_0g0n1n2noo3na0n1n2naao_012oo3a012aaox0  shft_asub_aadd_57_6_acx2
timestamp 1734143631
transform 1 0 480 0 -1 950
box 6 10 69 110
use _0_0cell_0_0g0n_0x2  shft_asub_aadd_57_6_acx3
timestamp 1734143631
transform 1 0 624 0 1 970
box 6 10 21 50
use _0_0cell_0_0g0n1n2naa_012aax0  shft_asub_acelem_acx0
timestamp 1734143631
transform 1 0 336 0 -1 1180
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  shft_asub_adelay1_acx0
timestamp 1734143631
transform 1 0 192 0 1 950
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay1_acx1
timestamp 1734143631
transform 1 0 132 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay1_acx2
timestamp 1734143631
transform 1 0 168 0 1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay1_acx3
timestamp 1734143631
transform 1 0 180 0 -1 710
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay1_acx4
timestamp 1734143631
transform 1 0 270 0 1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay1_acx5
timestamp 1734143631
transform 1 0 318 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay1_acx6
timestamp 1734143631
transform 1 0 252 0 -1 470
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay1_acx7
timestamp 1734143631
transform 1 0 108 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay2_acx0
timestamp 1734143631
transform 1 0 144 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay2_acx1
timestamp 1734143631
transform 1 0 180 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay2_acx2
timestamp 1734143631
transform 1 0 216 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay2_acx3
timestamp 1734143631
transform 1 0 252 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay2_acx4
timestamp 1734143631
transform 1 0 294 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay2_acx5
timestamp 1734143631
transform 1 0 342 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay2_acx6
timestamp 1734143631
transform 1 0 390 0 1 200
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asub_adelay2_acx7
timestamp 1734143631
transform 1 0 438 0 1 200
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  shft_asub_ainv__l1
timestamp 1734143760
transform 1 0 294 0 1 720
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_ainv__l2
timestamp 1734143760
transform 1 0 258 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_ainv__r
timestamp 1734143760
transform 1 0 420 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  shft_asub_al1_50_6
timestamp 1734143796
transform 1 0 1314 0 1 1430
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al1_51_6
timestamp 1734143796
transform 1 0 1158 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al1_52_6
timestamp 1734143796
transform 1 0 1320 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al1_53_6
timestamp 1734143796
transform 1 0 1194 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al1_54_6
timestamp 1734143796
transform 1 0 1398 0 1 480
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al1_55_6
timestamp 1734143796
transform 1 0 1038 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al1_56_6
timestamp 1734143796
transform 1 0 570 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al1_57_6
timestamp 1734143796
transform 1 0 528 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al2_50_6
timestamp 1734143796
transform 1 0 1320 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al2_51_6
timestamp 1734143796
transform 1 0 1392 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al2_52_6
timestamp 1734143796
transform 1 0 1266 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al2_53_6
timestamp 1734143796
transform 1 0 1302 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al2_54_6
timestamp 1734143796
transform 1 0 1344 0 -1 460
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al2_55_6
timestamp 1734143796
transform 1 0 918 0 1 480
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al2_56_6
timestamp 1734143796
transform 1 0 672 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asub_al2_57_6
timestamp 1734143796
transform 1 0 372 0 1 960
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  shft_asub_anor
timestamp 1734143909
transform 1 0 402 0 1 1190
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  shft_asub_aor__l1
timestamp 1734143975
transform 1 0 288 0 -1 940
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shft_asub_aor__l2
timestamp 1734143975
transform 1 0 282 0 -1 1180
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  shft_asub_apulseG_aand
timestamp 1734143631
transform 1 0 540 0 1 1420
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai1
timestamp 1734143760
transform 1 0 468 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai2
timestamp 1734143760
transform 1 0 510 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai3
timestamp 1734143760
transform 1 0 528 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai4
timestamp 1734143760
transform 1 0 558 0 1 1670
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai5
timestamp 1734143760
transform 1 0 558 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai6
timestamp 1734143760
transform 1 0 618 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai7
timestamp 1734143760
transform 1 0 684 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai8
timestamp 1734143760
transform 1 0 750 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai9
timestamp 1734143760
transform 1 0 822 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asub_apulseG_ai
timestamp 1734143760
transform 1 0 378 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  shft_asub_apulseG_anor
timestamp 1734143909
transform 1 0 450 0 1 1420
box 0 0 42 80
use _0_0std_0_0cells_0_0TIELOX1  shft_asub_atoGND
timestamp 1734144021
transform 1 0 1590 0 1 1680
box 0 0 30 50
use _0_0cell_0_0g0n1n2naa_012aax0  shft_asums_acelem_acx0
timestamp 1734143631
transform 1 0 558 0 -1 1180
box 6 10 65 70
use _0_0cell_0_0g0n_0x0  shft_asums_adelay1_acx0
timestamp 1734143631
transform 1 0 654 0 -1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asums_adelay1_acx1
timestamp 1734143631
transform 1 0 708 0 -1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asums_adelay1_acx2
timestamp 1734143631
transform 1 0 798 0 1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asums_adelay1_acx3
timestamp 1734143631
transform 1 0 714 0 1 1190
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asums_adelay1_acx4
timestamp 1734143631
transform 1 0 702 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asums_adelay1_acx5
timestamp 1734143631
transform 1 0 498 0 1 1420
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asums_adelay1_acx6
timestamp 1734143631
transform 1 0 420 0 -1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shft_asums_adelay1_acx7
timestamp 1734143631
transform 1 0 372 0 -1 1660
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  shft_asums_ainv__1
timestamp 1734143760
transform 1 0 510 0 -1 1180
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_ainv__2
timestamp 1734143760
transform 1 0 576 0 1 1200
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_ainv__3
timestamp 1734143760
transform 1 0 492 0 1 480
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  shft_asums_al_50_6
timestamp 1734143796
transform 1 0 1698 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asums_al_51_6
timestamp 1734143796
transform 1 0 1854 0 -1 1410
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asums_al_52_6
timestamp 1734143796
transform 1 0 1842 0 -1 1180
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asums_al_53_6
timestamp 1734143796
transform 1 0 1848 0 -1 940
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asums_al_54_6
timestamp 1734143796
transform 1 0 1854 0 1 720
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asums_al_55_6
timestamp 1734143796
transform 1 0 1734 0 -1 700
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asums_al_56_6
timestamp 1734143796
transform 1 0 1716 0 1 480
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shft_asums_al_57_6
timestamp 1734143796
transform 1 0 1602 0 1 480
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  shft_asums_anor__2
timestamp 1734143909
transform 1 0 510 0 1 1190
box 0 0 42 80
use _0_0std_0_0cells_0_0NOR2X1  shft_asums_anor__3
timestamp 1734143909
transform 1 0 216 0 1 1190
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  shft_asums_aor__1
timestamp 1734143975
transform 1 0 534 0 -1 700
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  shft_asums_apulseG_aand
timestamp 1734143631
transform 1 0 1824 0 1 470
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai
timestamp 1734143760
transform 1 0 1830 0 -1 700
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai1
timestamp 1734143760
transform 1 0 1872 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai2
timestamp 1734143760
transform 1 0 1944 0 -1 460
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai3
timestamp 1734143760
transform 1 0 1938 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai4
timestamp 1734143760
transform 1 0 1986 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai5
timestamp 1734143760
transform 1 0 2040 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai6
timestamp 1734143760
transform 1 0 2094 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai7
timestamp 1734143760
transform 1 0 1902 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai8
timestamp 1734143760
transform 1 0 1866 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shft_asums_apulseG_ai9
timestamp 1734143760
transform 1 0 1830 0 1 210
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  shft_asums_apulseG_anor
timestamp 1734143909
transform 1 0 1890 0 1 470
box 0 0 42 80
use _0_0std_0_0cells_0_0AND2X1  shift__split_aand1
timestamp 1734143631
transform 1 0 3438 0 -1 1900
box 0 0 60 80
use _0_0std_0_0cells_0_0AND2X1  shift__split_aand2
timestamp 1734143631
transform 1 0 3348 0 -1 1900
box 0 0 60 80
use _0_0cell_0_0g0n1n2naa_012aax0  shift__split_acelem_acx0
timestamp 1734143631
transform 1 0 2736 0 1 2380
box 6 10 65 70
use _0_0std_0_0cells_0_0LATCH  shift__split_acontrolLatch
timestamp 1734143796
transform 1 0 3054 0 -1 2120
box 0 0 96 80
use _0_0cell_0_0g0n_0x0  shift__split_adelay1_acx0
timestamp 1734143631
transform 1 0 3774 0 1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay1_acx1
timestamp 1734143631
transform 1 0 3756 0 -1 2370
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay1_acx2
timestamp 1734143631
transform 1 0 3834 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay1_acx3
timestamp 1734143631
transform 1 0 3960 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay1_acx4
timestamp 1734143631
transform 1 0 4092 0 1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay1_acx5
timestamp 1734143631
transform 1 0 4140 0 -1 2130
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay1_acx6
timestamp 1734143631
transform 1 0 4164 0 1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay1_acx7
timestamp 1734143631
transform 1 0 4152 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay2_acx0
timestamp 1734143631
transform 1 0 4188 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay2_acx1
timestamp 1734143631
transform 1 0 4188 0 1 1660
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay2_acx2
timestamp 1734143631
transform 1 0 4116 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay2_acx3
timestamp 1734143631
transform 1 0 4080 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay2_acx4
timestamp 1734143631
transform 1 0 4038 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay2_acx5
timestamp 1734143631
transform 1 0 3912 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay2_acx6
timestamp 1734143631
transform 1 0 3834 0 -1 1900
box 6 10 33 100
use _0_0cell_0_0g0n_0x0  shift__split_adelay2_acx7
timestamp 1734143631
transform 1 0 3618 0 -1 1900
box 6 10 33 100
use _0_0std_0_0cells_0_0INVX1  shift__split_ainv__c
timestamp 1734143760
transform 1 0 2466 0 -1 2600
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_ainv__ctr
timestamp 1734143760
transform 1 0 3282 0 -1 1890
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_ainv__l
timestamp 1734143760
transform 1 0 2694 0 1 2620
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_ainv__r
timestamp 1734143760
transform 1 0 2826 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0LATCH  shift__split_al_50_6
timestamp 1734143796
transform 1 0 3012 0 1 2140
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shift__split_al_51_6
timestamp 1734143796
transform 1 0 2958 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shift__split_al_52_6
timestamp 1734143796
transform 1 0 3282 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shift__split_al_53_6
timestamp 1734143796
transform 1 0 2856 0 -1 2120
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shift__split_al_54_6
timestamp 1734143796
transform 1 0 3138 0 -1 1650
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shift__split_al_55_6
timestamp 1734143796
transform 1 0 3144 0 1 1670
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shift__split_al_56_6
timestamp 1734143796
transform 1 0 3060 0 -1 1890
box 0 0 96 80
use _0_0std_0_0cells_0_0LATCH  shift__split_al_57_6
timestamp 1734143796
transform 1 0 3240 0 1 1910
box 0 0 96 80
use _0_0std_0_0cells_0_0NOR2X1  shift__split_anor__R
timestamp 1734143909
transform 1 0 2802 0 -1 2370
box 0 0 42 80
use _0_0std_0_0cells_0_0OR2X1  shift__split_aor1
timestamp 1734143975
transform 1 0 2724 0 -1 2600
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shift__split_aor2
timestamp 1734143975
transform 1 0 2502 0 -1 2600
box 0 0 54 70
use _0_0std_0_0cells_0_0OR2X1  shift__split_aor
timestamp 1734143975
transform 1 0 2868 0 -1 2360
box 0 0 54 70
use _0_0std_0_0cells_0_0AND2X1  shift__split_apulseG_aand
timestamp 1734143631
transform 1 0 3348 0 -1 1660
box 0 0 60 80
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai
timestamp 1734143760
transform 1 0 3408 0 1 2380
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai1
timestamp 1734143760
transform 1 0 3414 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai2
timestamp 1734143760
transform 1 0 3444 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai3
timestamp 1734143760
transform 1 0 3474 0 -1 1650
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai4
timestamp 1734143760
transform 1 0 3516 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai5
timestamp 1734143760
transform 1 0 3570 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai6
timestamp 1734143760
transform 1 0 3630 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai7
timestamp 1734143760
transform 1 0 3468 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai8
timestamp 1734143760
transform 1 0 3426 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0INVX1  shift__split_apulseG_ai9
timestamp 1734143760
transform 1 0 3390 0 1 1430
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  shift__split_apulseG_anor
timestamp 1734143909
transform 1 0 3414 0 1 1660
box 0 0 42 80
use _0_0std_0_0cells_0_0INVX1  sink__ctrl__lower_ai
timestamp 1734143760
transform 1 0 1998 0 1 2620
box 0 0 30 70
use _0_0std_0_0cells_0_0NOR2X1  sink__ctrl__lower_an
timestamp 1734143909
transform 1 0 1938 0 1 2610
box 0 0 42 80
<< labels >>
flabel m1 s 4269 2578 4272 2582 0 FreeSans 24 0 0 0 P.d[0]
port 0 nsew signal input
flabel m1 s 4269 3538 4272 3542 0 FreeSans 24 0 0 0 P.d[1]
port 1 nsew signal input
flabel m1 s 4269 658 4272 662 0 FreeSans 24 0 0 0 P.d[2]
port 2 nsew signal input
flabel m1 s 4269 1618 4272 1622 0 FreeSans 24 0 0 0 P.d[3]
port 3 nsew signal input
flabel m1 s 4269 1138 4272 1142 0 FreeSans 24 0 0 0 P.d[4]
port 4 nsew signal input
flabel m1 s 4269 2098 4272 2102 0 FreeSans 24 0 0 0 P.d[5]
port 5 nsew signal input
flabel m1 s 4269 3058 4272 3062 0 FreeSans 24 0 0 0 P.d[6]
port 6 nsew signal input
flabel m1 s 4269 4018 4272 4022 0 FreeSans 24 0 0 0 P.d[7]
port 7 nsew signal input
flabel m1 s 1462 4497 1466 4500 0 FreeSans 24 0 0 0 P.r
port 8 nsew signal input
flabel m1 s 2866 4497 2870 4500 0 FreeSans 24 0 0 0 P.a
port 9 nsew signal output
flabel m1 s 2740 180 2744 183 0 FreeSans 24 0 0 0 K.d[0]
port 10 nsew signal input
flabel m1 s 2164 180 2168 183 0 FreeSans 24 0 0 0 K.d[1]
port 11 nsew signal input
flabel m1 s 1396 180 1400 183 0 FreeSans 24 0 0 0 K.d[2]
port 12 nsew signal input
flabel m1 s 2356 180 2360 183 0 FreeSans 24 0 0 0 K.d[3]
port 13 nsew signal input
flabel m1 s 826 180 830 183 0 FreeSans 24 0 0 0 K.d[4]
port 14 nsew signal input
flabel m1 s 442 180 446 183 0 FreeSans 24 0 0 0 K.d[5]
port 15 nsew signal input
flabel m1 s 1972 180 1976 183 0 FreeSans 24 0 0 0 K.d[6]
port 16 nsew signal input
flabel m1 s 2548 180 2552 183 0 FreeSans 24 0 0 0 K.d[7]
port 17 nsew signal input
flabel m1 s 3502 180 3506 183 0 FreeSans 24 0 0 0 K.r
port 18 nsew signal input
flabel m1 s 3694 180 3698 183 0 FreeSans 24 0 0 0 K.a
port 19 nsew signal output
flabel m1 s 634 180 638 183 0 FreeSans 24 0 0 0 C.d[0]
port 20 nsew signal output
flabel m1 s 3124 180 3128 183 0 FreeSans 24 0 0 0 C.d[1]
port 21 nsew signal output
flabel m1 s 3886 180 3890 183 0 FreeSans 24 0 0 0 C.d[2]
port 22 nsew signal output
flabel m1 s 1018 180 1022 183 0 FreeSans 24 0 0 0 C.d[3]
port 23 nsew signal output
flabel m1 s 2932 180 2936 183 0 FreeSans 24 0 0 0 C.d[4]
port 24 nsew signal output
flabel m1 s 250 180 254 183 0 FreeSans 24 0 0 0 C.d[5]
port 25 nsew signal output
flabel m1 s 1588 180 1592 183 0 FreeSans 24 0 0 0 C.d[6]
port 26 nsew signal output
flabel m1 s 1780 180 1784 183 0 FreeSans 24 0 0 0 C.d[7]
port 27 nsew signal output
flabel m1 s 4078 180 4082 183 0 FreeSans 24 0 0 0 C.r
port 28 nsew signal output
flabel m1 s 3310 180 3314 183 0 FreeSans 24 0 0 0 C.a
port 29 nsew signal output
flabel m1 s 1204 180 1208 183 0 FreeSans 24 0 0 0 Reset
port 30 nsew signal input
<< properties >>
string FIXED_BBOX 60 180 4272 4500
<< end >>
