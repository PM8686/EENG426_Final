magic
tech sky130l
timestamp 1731220350
<< m1 >>
rect 1568 3891 1572 3915
rect 448 3731 452 3767
rect 1600 3731 1604 3767
rect 2272 3743 2276 3767
rect 3672 3743 3676 3795
rect 272 3479 276 3583
rect 1128 3567 1132 3591
rect 2992 3575 2996 3599
rect 3000 3575 3004 3615
rect 1216 3387 1220 3411
rect 1384 3387 1388 3411
rect 3456 3279 3460 3323
rect 3208 3251 3212 3275
rect 256 3219 260 3243
rect 2840 3135 2844 3155
rect 648 2923 652 2951
rect 648 2919 656 2923
rect 664 2883 668 2907
rect 3760 2787 3764 2819
rect 3040 2759 3044 2783
rect 3232 2759 3236 2783
rect 3640 2759 3644 2783
rect 664 2719 668 2743
rect 1512 2719 1516 2743
rect 2720 2627 2724 2655
rect 2904 2579 2908 2603
rect 1296 2551 1300 2575
rect 656 2379 660 2403
rect 1520 2379 1524 2431
rect 888 2263 892 2291
rect 888 2259 896 2263
rect 944 2219 948 2243
rect 240 2099 244 2127
rect 1128 2099 1132 2127
rect 1488 2051 1492 2087
rect 2904 1967 2908 2055
rect 3792 1943 3796 1987
rect 3216 1915 3220 1939
rect 712 1883 716 1907
rect 832 1883 836 1907
rect 952 1883 956 1907
rect 1544 1883 1548 1907
rect 1664 1883 1668 1907
rect 3032 1811 3036 1911
rect 2944 1759 2948 1783
rect 1248 1723 1252 1747
rect 240 1607 244 1635
rect 704 1563 708 1587
rect 392 1455 396 1475
rect 3720 1459 3724 1511
rect 408 1399 412 1443
rect 3120 1431 3124 1455
rect 552 1399 556 1423
rect 800 1399 804 1423
rect 1424 1399 1428 1423
rect 3704 1327 3708 1347
rect 888 1243 892 1275
rect 1640 1243 1644 1267
rect 1136 1087 1140 1111
rect 1504 1087 1508 1119
rect 400 931 404 955
rect 728 931 732 955
rect 3208 787 3212 811
rect 728 467 732 491
rect 1520 467 1524 511
rect 232 311 236 335
rect 896 151 900 223
rect 240 123 244 147
rect 336 123 340 147
rect 1400 123 1404 147
rect 1504 123 1508 147
rect 1608 123 1612 147
rect 2160 135 2164 159
<< m2c >>
rect 2136 3947 2140 3951
rect 2392 3947 2396 3951
rect 2656 3947 2660 3951
rect 2904 3947 2908 3951
rect 3152 3947 3156 3951
rect 3408 3947 3412 3951
rect 2192 3935 2196 3939
rect 2336 3935 2340 3939
rect 2504 3935 2508 3939
rect 2680 3935 2684 3939
rect 2864 3935 2868 3939
rect 3048 3935 3052 3939
rect 3240 3935 3244 3939
rect 3432 3935 3436 3939
rect 3624 3935 3628 3939
rect 376 3927 380 3931
rect 576 3927 580 3931
rect 768 3927 772 3931
rect 952 3927 956 3931
rect 1128 3927 1132 3931
rect 1296 3927 1300 3931
rect 1448 3927 1452 3931
rect 1584 3927 1588 3931
rect 1720 3927 1724 3931
rect 1856 3927 1860 3931
rect 1968 3927 1972 3931
rect 344 3915 348 3919
rect 480 3915 484 3919
rect 632 3915 636 3919
rect 800 3915 804 3919
rect 976 3915 980 3919
rect 1160 3915 1164 3919
rect 1352 3915 1356 3919
rect 1544 3915 1548 3919
rect 1568 3915 1572 3919
rect 1744 3915 1748 3919
rect 1568 3887 1572 3891
rect 2328 3795 2332 3799
rect 2440 3795 2444 3799
rect 2560 3795 2564 3799
rect 2696 3795 2700 3799
rect 2840 3795 2844 3799
rect 2984 3795 2988 3799
rect 3128 3795 3132 3799
rect 3272 3795 3276 3799
rect 3408 3795 3412 3799
rect 3536 3795 3540 3799
rect 3664 3795 3668 3799
rect 3672 3795 3676 3799
rect 3792 3795 3796 3799
rect 3904 3795 3908 3799
rect 296 3767 300 3771
rect 400 3767 404 3771
rect 448 3767 452 3771
rect 504 3767 508 3771
rect 600 3767 604 3771
rect 696 3767 700 3771
rect 792 3767 796 3771
rect 896 3767 900 3771
rect 1000 3767 1004 3771
rect 1104 3767 1108 3771
rect 1216 3767 1220 3771
rect 1328 3767 1332 3771
rect 1448 3767 1452 3771
rect 1568 3767 1572 3771
rect 1600 3767 1604 3771
rect 1696 3767 1700 3771
rect 2136 3767 2140 3771
rect 2248 3767 2252 3771
rect 2272 3767 2276 3771
rect 2392 3767 2396 3771
rect 2544 3767 2548 3771
rect 2704 3767 2708 3771
rect 2872 3767 2876 3771
rect 3048 3767 3052 3771
rect 3224 3767 3228 3771
rect 3400 3767 3404 3771
rect 3576 3767 3580 3771
rect 224 3755 228 3759
rect 416 3755 420 3759
rect 616 3755 620 3759
rect 816 3755 820 3759
rect 1024 3755 1028 3759
rect 1232 3755 1236 3759
rect 1448 3755 1452 3759
rect 448 3727 452 3731
rect 1672 3755 1676 3759
rect 2272 3739 2276 3743
rect 3752 3767 3756 3771
rect 3904 3767 3908 3771
rect 3672 3739 3676 3743
rect 1600 3727 1604 3731
rect 2136 3615 2140 3619
rect 2264 3615 2268 3619
rect 2432 3615 2436 3619
rect 2616 3615 2620 3619
rect 2800 3615 2804 3619
rect 2992 3615 2996 3619
rect 3000 3615 3004 3619
rect 3176 3615 3180 3619
rect 3360 3615 3364 3619
rect 3544 3615 3548 3619
rect 3736 3615 3740 3619
rect 3904 3615 3908 3619
rect 216 3607 220 3611
rect 448 3607 452 3611
rect 680 3607 684 3611
rect 904 3607 908 3611
rect 1120 3607 1124 3611
rect 1328 3607 1332 3611
rect 1544 3607 1548 3611
rect 1760 3607 1764 3611
rect 2168 3599 2172 3603
rect 2344 3599 2348 3603
rect 2536 3599 2540 3603
rect 2736 3599 2740 3603
rect 2936 3599 2940 3603
rect 2992 3599 2996 3603
rect 232 3591 236 3595
rect 424 3591 428 3595
rect 624 3591 628 3595
rect 840 3591 844 3595
rect 1056 3591 1060 3595
rect 1128 3591 1132 3595
rect 1280 3591 1284 3595
rect 1512 3591 1516 3595
rect 1752 3591 1756 3595
rect 272 3583 276 3587
rect 2992 3571 2996 3575
rect 3128 3599 3132 3603
rect 3320 3599 3324 3603
rect 3512 3599 3516 3603
rect 3704 3599 3708 3603
rect 3904 3599 3908 3603
rect 3000 3571 3004 3575
rect 1128 3563 1132 3567
rect 272 3475 276 3479
rect 2392 3455 2396 3459
rect 2512 3455 2516 3459
rect 2648 3455 2652 3459
rect 2800 3455 2804 3459
rect 2976 3455 2980 3459
rect 3176 3455 3180 3459
rect 3400 3455 3404 3459
rect 3632 3455 3636 3459
rect 3872 3455 3876 3459
rect 360 3443 364 3447
rect 496 3443 500 3447
rect 648 3443 652 3447
rect 808 3443 812 3447
rect 976 3443 980 3447
rect 1144 3443 1148 3447
rect 1312 3443 1316 3447
rect 1488 3443 1492 3447
rect 1664 3443 1668 3447
rect 1840 3443 1844 3447
rect 2512 3443 2516 3447
rect 2616 3443 2620 3447
rect 2728 3443 2732 3447
rect 2840 3443 2844 3447
rect 2968 3443 2972 3447
rect 3112 3443 3116 3447
rect 3272 3443 3276 3447
rect 3448 3443 3452 3447
rect 3632 3443 3636 3447
rect 3816 3443 3820 3447
rect 560 3411 564 3415
rect 712 3411 716 3415
rect 864 3411 868 3415
rect 1024 3411 1028 3415
rect 1192 3411 1196 3415
rect 1216 3411 1220 3415
rect 1360 3411 1364 3415
rect 1384 3411 1388 3415
rect 1528 3411 1532 3415
rect 1704 3411 1708 3415
rect 1880 3411 1884 3415
rect 1216 3383 1220 3387
rect 1384 3383 1388 3387
rect 3456 3323 3460 3327
rect 2632 3291 2636 3295
rect 2784 3291 2788 3295
rect 2936 3291 2940 3295
rect 3088 3291 3092 3295
rect 3240 3291 3244 3295
rect 3392 3291 3396 3295
rect 3544 3291 3548 3295
rect 3696 3291 3700 3295
rect 3848 3291 3852 3295
rect 2480 3275 2484 3279
rect 2616 3275 2620 3279
rect 2752 3275 2756 3279
rect 2896 3275 2900 3279
rect 3040 3275 3044 3279
rect 3184 3275 3188 3279
rect 3208 3275 3212 3279
rect 3320 3275 3324 3279
rect 3448 3275 3452 3279
rect 3456 3275 3460 3279
rect 3568 3275 3572 3279
rect 3688 3275 3692 3279
rect 3808 3275 3812 3279
rect 3904 3275 3908 3279
rect 360 3259 364 3263
rect 544 3259 548 3263
rect 736 3259 740 3263
rect 928 3259 932 3263
rect 1120 3259 1124 3263
rect 1312 3259 1316 3263
rect 1504 3259 1508 3263
rect 1696 3259 1700 3263
rect 1888 3259 1892 3263
rect 3208 3247 3212 3251
rect 200 3243 204 3247
rect 256 3243 260 3247
rect 384 3243 388 3247
rect 584 3243 588 3247
rect 784 3243 788 3247
rect 976 3243 980 3247
rect 1160 3243 1164 3247
rect 1336 3243 1340 3247
rect 1512 3243 1516 3247
rect 1688 3243 1692 3247
rect 1864 3243 1868 3247
rect 256 3215 260 3219
rect 2840 3155 2844 3159
rect 2840 3131 2844 3135
rect 2312 3123 2316 3127
rect 2464 3123 2468 3127
rect 2624 3123 2628 3127
rect 2792 3123 2796 3127
rect 2968 3123 2972 3127
rect 3144 3123 3148 3127
rect 3328 3123 3332 3127
rect 3512 3123 3516 3127
rect 3696 3123 3700 3127
rect 3880 3123 3884 3127
rect 2144 3107 2148 3111
rect 2288 3107 2292 3111
rect 2440 3107 2444 3111
rect 2592 3107 2596 3111
rect 2752 3107 2756 3111
rect 2920 3107 2924 3111
rect 3104 3107 3108 3111
rect 3296 3107 3300 3111
rect 3496 3107 3500 3111
rect 3704 3107 3708 3111
rect 3904 3107 3908 3111
rect 208 3095 212 3099
rect 408 3095 412 3099
rect 608 3095 612 3099
rect 808 3095 812 3099
rect 992 3095 996 3099
rect 1168 3095 1172 3099
rect 1328 3095 1332 3099
rect 1488 3095 1492 3099
rect 1640 3095 1644 3099
rect 1800 3095 1804 3099
rect 328 3083 332 3087
rect 504 3083 508 3087
rect 680 3083 684 3087
rect 864 3083 868 3087
rect 1040 3083 1044 3087
rect 1208 3083 1212 3087
rect 1368 3083 1372 3087
rect 1520 3083 1524 3087
rect 1672 3083 1676 3087
rect 1832 3083 1836 3087
rect 2136 2959 2140 2963
rect 2248 2959 2252 2963
rect 2392 2959 2396 2963
rect 2544 2959 2548 2963
rect 2720 2959 2724 2963
rect 2920 2959 2924 2963
rect 3152 2959 3156 2963
rect 3400 2959 3404 2963
rect 3664 2959 3668 2963
rect 3904 2959 3908 2963
rect 648 2951 652 2955
rect 2136 2943 2140 2947
rect 2328 2943 2332 2947
rect 2552 2943 2556 2947
rect 2800 2943 2804 2947
rect 3064 2943 3068 2947
rect 3344 2943 3348 2947
rect 3632 2943 3636 2947
rect 3904 2943 3908 2947
rect 408 2919 412 2923
rect 504 2919 508 2923
rect 608 2919 612 2923
rect 656 2919 660 2923
rect 720 2919 724 2923
rect 848 2919 852 2923
rect 1000 2919 1004 2923
rect 1168 2919 1172 2923
rect 1360 2919 1364 2923
rect 1560 2919 1564 2923
rect 1776 2919 1780 2923
rect 1968 2919 1972 2923
rect 272 2907 276 2911
rect 392 2907 396 2911
rect 512 2907 516 2911
rect 640 2907 644 2911
rect 664 2907 668 2911
rect 768 2907 772 2911
rect 912 2907 916 2911
rect 1064 2907 1068 2911
rect 1232 2907 1236 2911
rect 1416 2907 1420 2911
rect 1600 2907 1604 2911
rect 1792 2907 1796 2911
rect 1968 2907 1972 2911
rect 664 2879 668 2883
rect 3760 2819 3764 2823
rect 2736 2795 2740 2799
rect 2952 2795 2956 2799
rect 3160 2795 3164 2799
rect 3352 2795 3356 2799
rect 3544 2795 3548 2799
rect 3736 2795 3740 2799
rect 3904 2795 3908 2799
rect 2136 2783 2140 2787
rect 2264 2783 2268 2787
rect 2408 2783 2412 2787
rect 2544 2783 2548 2787
rect 2672 2783 2676 2787
rect 2792 2783 2796 2787
rect 2904 2783 2908 2787
rect 3008 2783 3012 2787
rect 3040 2783 3044 2787
rect 3112 2783 3116 2787
rect 3208 2783 3212 2787
rect 3232 2783 3236 2787
rect 3304 2783 3308 2787
rect 3408 2783 3412 2787
rect 3512 2783 3516 2787
rect 3616 2783 3620 2787
rect 3640 2783 3644 2787
rect 3712 2783 3716 2787
rect 3760 2783 3764 2787
rect 3808 2783 3812 2787
rect 3904 2783 3908 2787
rect 200 2763 204 2767
rect 312 2763 316 2767
rect 464 2763 468 2767
rect 616 2763 620 2767
rect 776 2763 780 2767
rect 944 2763 948 2767
rect 1112 2763 1116 2767
rect 1288 2763 1292 2767
rect 1464 2763 1468 2767
rect 1640 2763 1644 2767
rect 1816 2763 1820 2767
rect 1968 2763 1972 2767
rect 3040 2755 3044 2759
rect 3232 2755 3236 2759
rect 3640 2755 3644 2759
rect 200 2743 204 2747
rect 320 2743 324 2747
rect 472 2743 476 2747
rect 640 2743 644 2747
rect 664 2743 668 2747
rect 808 2743 812 2747
rect 984 2743 988 2747
rect 1152 2743 1156 2747
rect 1320 2743 1324 2747
rect 1488 2743 1492 2747
rect 1512 2743 1516 2747
rect 1664 2743 1668 2747
rect 664 2715 668 2719
rect 1512 2715 1516 2719
rect 2720 2655 2724 2659
rect 2160 2623 2164 2627
rect 2328 2623 2332 2627
rect 2504 2623 2508 2627
rect 2680 2623 2684 2627
rect 2720 2623 2724 2627
rect 2848 2623 2852 2627
rect 3008 2623 3012 2627
rect 3160 2623 3164 2627
rect 3304 2623 3308 2627
rect 3448 2623 3452 2627
rect 3600 2623 3604 2627
rect 232 2603 236 2607
rect 424 2603 428 2607
rect 624 2603 628 2607
rect 824 2603 828 2607
rect 1016 2603 1020 2607
rect 1208 2603 1212 2607
rect 1392 2603 1396 2607
rect 1576 2603 1580 2607
rect 1768 2603 1772 2607
rect 2280 2603 2284 2607
rect 2432 2603 2436 2607
rect 2584 2603 2588 2607
rect 2736 2603 2740 2607
rect 2880 2603 2884 2607
rect 2904 2603 2908 2607
rect 3016 2603 3020 2607
rect 3152 2603 3156 2607
rect 3288 2603 3292 2607
rect 3432 2603 3436 2607
rect 640 2575 644 2579
rect 752 2575 756 2579
rect 872 2575 876 2579
rect 1000 2575 1004 2579
rect 1136 2575 1140 2579
rect 1272 2575 1276 2579
rect 1296 2575 1300 2579
rect 1416 2575 1420 2579
rect 1560 2575 1564 2579
rect 1712 2575 1716 2579
rect 1864 2575 1868 2579
rect 2904 2575 2908 2579
rect 1296 2547 1300 2551
rect 2160 2459 2164 2463
rect 2280 2459 2284 2463
rect 2408 2459 2412 2463
rect 2536 2459 2540 2463
rect 2664 2459 2668 2463
rect 2784 2459 2788 2463
rect 2904 2459 2908 2463
rect 3032 2459 3036 2463
rect 3160 2459 3164 2463
rect 3288 2459 3292 2463
rect 2136 2435 2140 2439
rect 2256 2435 2260 2439
rect 2384 2435 2388 2439
rect 2504 2435 2508 2439
rect 2624 2435 2628 2439
rect 2744 2435 2748 2439
rect 2856 2435 2860 2439
rect 2976 2435 2980 2439
rect 3096 2435 3100 2439
rect 3216 2435 3220 2439
rect 568 2431 572 2435
rect 672 2431 676 2435
rect 784 2431 788 2435
rect 912 2431 916 2435
rect 1048 2431 1052 2435
rect 1192 2431 1196 2435
rect 1344 2431 1348 2435
rect 1496 2431 1500 2435
rect 1520 2431 1524 2435
rect 1648 2431 1652 2435
rect 1808 2431 1812 2435
rect 1968 2431 1972 2435
rect 600 2403 604 2407
rect 656 2403 660 2407
rect 736 2403 740 2407
rect 880 2403 884 2407
rect 1024 2403 1028 2407
rect 1168 2403 1172 2407
rect 1312 2403 1316 2407
rect 1456 2403 1460 2407
rect 656 2375 660 2379
rect 1592 2403 1596 2407
rect 1720 2403 1724 2407
rect 1856 2403 1860 2407
rect 1968 2403 1972 2407
rect 1520 2375 1524 2379
rect 888 2291 892 2295
rect 2232 2291 2236 2295
rect 2424 2293 2428 2297
rect 2600 2291 2604 2295
rect 2768 2291 2772 2295
rect 2936 2291 2940 2295
rect 3096 2291 3100 2295
rect 3264 2291 3268 2295
rect 2136 2279 2140 2283
rect 2232 2279 2236 2283
rect 2352 2279 2356 2283
rect 2488 2279 2492 2283
rect 2624 2279 2628 2283
rect 2768 2279 2772 2283
rect 2904 2279 2908 2283
rect 3048 2279 3052 2283
rect 3192 2279 3196 2283
rect 3336 2279 3340 2283
rect 600 2259 604 2263
rect 712 2259 716 2263
rect 832 2259 836 2263
rect 896 2259 900 2263
rect 960 2259 964 2263
rect 1096 2259 1100 2263
rect 1232 2259 1236 2263
rect 1360 2259 1364 2263
rect 1488 2259 1492 2263
rect 1616 2259 1620 2263
rect 1736 2259 1740 2263
rect 1864 2259 1868 2263
rect 1968 2259 1972 2263
rect 480 2243 484 2247
rect 600 2243 604 2247
rect 736 2243 740 2247
rect 888 2243 892 2247
rect 944 2243 948 2247
rect 1056 2243 1060 2247
rect 1240 2243 1244 2247
rect 1432 2243 1436 2247
rect 1632 2243 1636 2247
rect 1832 2243 1836 2247
rect 944 2215 948 2219
rect 2136 2139 2140 2143
rect 2360 2139 2364 2143
rect 2568 2139 2572 2143
rect 2752 2139 2756 2143
rect 2928 2139 2932 2143
rect 3088 2139 3092 2143
rect 3240 2139 3244 2143
rect 3384 2139 3388 2143
rect 3536 2139 3540 2143
rect 240 2127 244 2131
rect 1128 2127 1132 2131
rect 2464 2103 2468 2107
rect 2560 2103 2564 2107
rect 2656 2103 2660 2107
rect 2752 2103 2756 2107
rect 2848 2103 2852 2107
rect 2944 2103 2948 2107
rect 3040 2103 3044 2107
rect 3136 2103 3140 2107
rect 3232 2103 3236 2107
rect 3328 2103 3332 2107
rect 3424 2103 3428 2107
rect 3520 2103 3524 2107
rect 3616 2103 3620 2107
rect 3712 2103 3716 2107
rect 3808 2103 3812 2107
rect 3904 2103 3908 2107
rect 200 2095 204 2099
rect 240 2095 244 2099
rect 312 2095 316 2099
rect 456 2095 460 2099
rect 616 2095 620 2099
rect 776 2095 780 2099
rect 936 2095 940 2099
rect 1096 2095 1100 2099
rect 1128 2095 1132 2099
rect 1256 2095 1260 2099
rect 1416 2095 1420 2099
rect 1576 2095 1580 2099
rect 1744 2095 1748 2099
rect 1488 2087 1492 2091
rect 200 2075 204 2079
rect 312 2075 316 2079
rect 464 2075 468 2079
rect 616 2075 620 2079
rect 768 2075 772 2079
rect 912 2075 916 2079
rect 1056 2075 1060 2079
rect 1192 2075 1196 2079
rect 1320 2075 1324 2079
rect 1448 2075 1452 2079
rect 1584 2075 1588 2079
rect 1488 2047 1492 2051
rect 2904 2055 2908 2059
rect 3792 1987 3796 1991
rect 2256 1963 2260 1967
rect 2464 1963 2468 1967
rect 2712 1963 2716 1967
rect 2904 1963 2908 1967
rect 2984 1963 2988 1967
rect 3280 1963 3284 1967
rect 3592 1963 3596 1967
rect 3904 1963 3908 1967
rect 2136 1939 2140 1943
rect 2304 1939 2308 1943
rect 2512 1939 2516 1943
rect 2736 1939 2740 1943
rect 2960 1939 2964 1943
rect 3192 1939 3196 1943
rect 3216 1939 3220 1943
rect 3424 1939 3428 1943
rect 3656 1939 3660 1943
rect 3792 1939 3796 1943
rect 3896 1939 3900 1943
rect 296 1919 300 1923
rect 456 1919 460 1923
rect 632 1919 636 1923
rect 816 1919 820 1923
rect 1008 1919 1012 1923
rect 1200 1919 1204 1923
rect 1400 1919 1404 1923
rect 1608 1919 1612 1923
rect 3032 1911 3036 1915
rect 3216 1911 3220 1915
rect 576 1907 580 1911
rect 688 1907 692 1911
rect 712 1907 716 1911
rect 808 1907 812 1911
rect 832 1907 836 1911
rect 928 1907 932 1911
rect 952 1907 956 1911
rect 1048 1907 1052 1911
rect 1168 1907 1172 1911
rect 1288 1907 1292 1911
rect 1400 1907 1404 1911
rect 1520 1907 1524 1911
rect 1544 1907 1548 1911
rect 1640 1907 1644 1911
rect 1664 1907 1668 1911
rect 1760 1907 1764 1911
rect 712 1879 716 1883
rect 832 1879 836 1883
rect 952 1879 956 1883
rect 1544 1879 1548 1883
rect 1664 1879 1668 1883
rect 3032 1807 3036 1811
rect 2136 1799 2140 1803
rect 2264 1799 2268 1803
rect 2432 1799 2436 1803
rect 2608 1799 2612 1803
rect 2784 1799 2788 1803
rect 2952 1799 2956 1803
rect 3104 1799 3108 1803
rect 3248 1799 3252 1803
rect 3384 1799 3388 1803
rect 3520 1799 3524 1803
rect 3648 1799 3652 1803
rect 3776 1799 3780 1803
rect 3904 1799 3908 1803
rect 2136 1783 2140 1787
rect 2248 1783 2252 1787
rect 2392 1783 2396 1787
rect 2552 1783 2556 1787
rect 2720 1783 2724 1787
rect 2896 1783 2900 1787
rect 2944 1783 2948 1787
rect 3088 1783 3092 1787
rect 3288 1783 3292 1787
rect 3496 1783 3500 1787
rect 3712 1783 3716 1787
rect 3904 1783 3908 1787
rect 680 1759 684 1763
rect 776 1759 780 1763
rect 880 1759 884 1763
rect 992 1759 996 1763
rect 1104 1759 1108 1763
rect 1224 1759 1228 1763
rect 1344 1759 1348 1763
rect 1464 1759 1468 1763
rect 1584 1759 1588 1763
rect 1704 1759 1708 1763
rect 2944 1755 2948 1759
rect 432 1747 436 1751
rect 560 1747 564 1751
rect 704 1747 708 1751
rect 864 1747 868 1751
rect 1032 1747 1036 1751
rect 1208 1747 1212 1751
rect 1248 1747 1252 1751
rect 1392 1747 1396 1751
rect 1576 1747 1580 1751
rect 1768 1747 1772 1751
rect 1248 1719 1252 1723
rect 240 1635 244 1639
rect 2288 1635 2292 1639
rect 2392 1635 2396 1639
rect 2504 1635 2508 1639
rect 2624 1635 2628 1639
rect 2752 1635 2756 1639
rect 2888 1635 2892 1639
rect 3032 1635 3036 1639
rect 3192 1635 3196 1639
rect 3368 1635 3372 1639
rect 3552 1635 3556 1639
rect 3736 1635 3740 1639
rect 3904 1635 3908 1639
rect 2456 1619 2460 1623
rect 2568 1619 2572 1623
rect 2680 1619 2684 1623
rect 2800 1619 2804 1623
rect 2920 1619 2924 1623
rect 3040 1619 3044 1623
rect 3160 1619 3164 1623
rect 3280 1619 3284 1623
rect 3400 1619 3404 1623
rect 3520 1619 3524 1623
rect 200 1603 204 1607
rect 240 1603 244 1607
rect 312 1603 316 1607
rect 464 1603 468 1607
rect 632 1603 636 1607
rect 808 1603 812 1607
rect 1000 1603 1004 1607
rect 1200 1603 1204 1607
rect 1408 1603 1412 1607
rect 1616 1603 1620 1607
rect 1832 1603 1836 1607
rect 200 1587 204 1591
rect 320 1587 324 1591
rect 488 1587 492 1591
rect 680 1587 684 1591
rect 704 1587 708 1591
rect 896 1587 900 1591
rect 1128 1587 1132 1591
rect 1376 1587 1380 1591
rect 1632 1587 1636 1591
rect 1896 1587 1900 1591
rect 704 1559 708 1563
rect 3720 1511 3724 1515
rect 2608 1479 2612 1483
rect 2736 1479 2740 1483
rect 2864 1479 2868 1483
rect 3000 1479 3004 1483
rect 3136 1479 3140 1483
rect 3272 1479 3276 1483
rect 3400 1479 3404 1483
rect 3528 1479 3532 1483
rect 3656 1479 3660 1483
rect 392 1475 396 1479
rect 3792 1479 3796 1483
rect 3904 1479 3908 1483
rect 2584 1455 2588 1459
rect 2696 1455 2700 1459
rect 2824 1455 2828 1459
rect 2960 1455 2964 1459
rect 3096 1455 3100 1459
rect 3120 1455 3124 1459
rect 3240 1455 3244 1459
rect 3376 1455 3380 1459
rect 3512 1455 3516 1459
rect 3648 1455 3652 1459
rect 3720 1455 3724 1459
rect 3784 1455 3788 1459
rect 3904 1455 3908 1459
rect 392 1451 396 1455
rect 304 1443 308 1447
rect 408 1443 412 1447
rect 472 1443 476 1447
rect 648 1443 652 1447
rect 840 1443 844 1447
rect 1032 1443 1036 1447
rect 1224 1443 1228 1447
rect 1416 1443 1420 1447
rect 1608 1443 1612 1447
rect 1800 1443 1804 1447
rect 1968 1443 1972 1447
rect 3120 1427 3124 1431
rect 528 1423 532 1427
rect 552 1423 556 1427
rect 648 1423 652 1427
rect 776 1423 780 1427
rect 800 1423 804 1427
rect 920 1423 924 1427
rect 1072 1423 1076 1427
rect 1232 1423 1236 1427
rect 1400 1423 1404 1427
rect 1424 1423 1428 1427
rect 1576 1423 1580 1427
rect 1752 1423 1756 1427
rect 1936 1423 1940 1427
rect 408 1395 412 1399
rect 552 1395 556 1399
rect 800 1395 804 1399
rect 1424 1395 1428 1399
rect 3704 1347 3708 1351
rect 3704 1323 3708 1327
rect 2464 1315 2468 1319
rect 2600 1315 2604 1319
rect 2744 1315 2748 1319
rect 2888 1315 2892 1319
rect 3032 1315 3036 1319
rect 3176 1315 3180 1319
rect 3320 1315 3324 1319
rect 3472 1315 3476 1319
rect 3624 1315 3628 1319
rect 3776 1315 3780 1319
rect 3904 1315 3908 1319
rect 2312 1299 2316 1303
rect 2440 1299 2444 1303
rect 2576 1299 2580 1303
rect 2712 1299 2716 1303
rect 2856 1299 2860 1303
rect 3008 1299 3012 1303
rect 3176 1299 3180 1303
rect 3352 1299 3356 1303
rect 3536 1299 3540 1303
rect 3728 1299 3732 1303
rect 3904 1299 3908 1303
rect 720 1283 724 1287
rect 832 1283 836 1287
rect 952 1283 956 1287
rect 1080 1283 1084 1287
rect 1208 1283 1212 1287
rect 1344 1283 1348 1287
rect 1480 1283 1484 1287
rect 1624 1283 1628 1287
rect 1768 1283 1772 1287
rect 1912 1283 1916 1287
rect 888 1275 892 1279
rect 504 1267 508 1271
rect 616 1267 620 1271
rect 736 1267 740 1271
rect 864 1267 868 1271
rect 1000 1267 1004 1271
rect 1144 1267 1148 1271
rect 1296 1267 1300 1271
rect 1456 1267 1460 1271
rect 1616 1267 1620 1271
rect 1640 1267 1644 1271
rect 1784 1267 1788 1271
rect 888 1239 892 1243
rect 1640 1239 1644 1243
rect 2136 1155 2140 1159
rect 2248 1155 2252 1159
rect 2368 1155 2372 1159
rect 2496 1155 2500 1159
rect 2624 1155 2628 1159
rect 2776 1155 2780 1159
rect 2952 1155 2956 1159
rect 3152 1155 3156 1159
rect 3376 1155 3380 1159
rect 3608 1155 3612 1159
rect 3848 1155 3852 1159
rect 2136 1139 2140 1143
rect 2264 1139 2268 1143
rect 2416 1139 2420 1143
rect 2576 1139 2580 1143
rect 2744 1139 2748 1143
rect 2936 1139 2940 1143
rect 3152 1139 3156 1143
rect 3384 1139 3388 1143
rect 3624 1139 3628 1143
rect 3872 1139 3876 1143
rect 232 1127 236 1131
rect 368 1127 372 1131
rect 528 1127 532 1131
rect 696 1127 700 1131
rect 872 1127 876 1131
rect 1048 1127 1052 1131
rect 1224 1127 1228 1131
rect 1400 1127 1404 1131
rect 1576 1127 1580 1131
rect 1760 1127 1764 1131
rect 1504 1119 1508 1123
rect 200 1111 204 1115
rect 304 1111 308 1115
rect 440 1111 444 1115
rect 592 1111 596 1115
rect 760 1111 764 1115
rect 928 1111 932 1115
rect 1104 1111 1108 1115
rect 1136 1111 1140 1115
rect 1280 1111 1284 1115
rect 1456 1111 1460 1115
rect 1136 1083 1140 1087
rect 1632 1111 1636 1115
rect 1808 1111 1812 1115
rect 1968 1111 1972 1115
rect 1504 1083 1508 1087
rect 2136 987 2140 991
rect 2328 987 2332 991
rect 2552 987 2556 991
rect 2768 987 2772 991
rect 2984 987 2988 991
rect 3184 987 3188 991
rect 3376 987 3380 991
rect 3560 987 3564 991
rect 3744 987 3748 991
rect 3904 987 3908 991
rect 200 971 204 975
rect 352 971 356 975
rect 536 971 540 975
rect 720 971 724 975
rect 904 971 908 975
rect 1080 971 1084 975
rect 1264 971 1268 975
rect 1448 971 1452 975
rect 1632 971 1636 975
rect 2368 971 2372 975
rect 2520 971 2524 975
rect 2680 971 2684 975
rect 2848 971 2852 975
rect 3016 971 3020 975
rect 3176 971 3180 975
rect 3328 971 3332 975
rect 3480 971 3484 975
rect 3624 971 3628 975
rect 3776 971 3780 975
rect 3904 971 3908 975
rect 200 955 204 959
rect 360 955 364 959
rect 400 955 404 959
rect 536 955 540 959
rect 704 955 708 959
rect 728 955 732 959
rect 864 955 868 959
rect 1016 955 1020 959
rect 1152 955 1156 959
rect 1288 955 1292 959
rect 1424 955 1428 959
rect 1560 955 1564 959
rect 400 927 404 931
rect 728 927 732 931
rect 2624 827 2628 831
rect 2744 827 2748 831
rect 2872 827 2876 831
rect 3008 827 3012 831
rect 3144 827 3148 831
rect 3272 827 3276 831
rect 3400 827 3404 831
rect 3528 827 3532 831
rect 3656 827 3660 831
rect 3792 827 3796 831
rect 3904 827 3908 831
rect 224 815 228 819
rect 384 815 388 819
rect 536 815 540 819
rect 680 815 684 819
rect 816 815 820 819
rect 944 815 948 819
rect 1064 815 1068 819
rect 1176 815 1180 819
rect 1296 815 1300 819
rect 1416 815 1420 819
rect 2400 811 2404 815
rect 2536 811 2540 815
rect 2680 811 2684 815
rect 2832 811 2836 815
rect 2984 811 2988 815
rect 3144 811 3148 815
rect 3208 811 3212 815
rect 3304 811 3308 815
rect 3456 811 3460 815
rect 3608 811 3612 815
rect 3768 811 3772 815
rect 3904 811 3908 815
rect 288 803 292 807
rect 448 803 452 807
rect 600 803 604 807
rect 744 803 748 807
rect 880 803 884 807
rect 1016 803 1020 807
rect 1144 803 1148 807
rect 1264 803 1268 807
rect 1392 803 1396 807
rect 1520 803 1524 807
rect 3208 783 3212 787
rect 2136 667 2140 671
rect 2248 667 2252 671
rect 2400 667 2404 671
rect 2552 667 2556 671
rect 2704 667 2708 671
rect 2872 667 2876 671
rect 3048 667 3052 671
rect 3232 667 3236 671
rect 3432 667 3436 671
rect 3640 667 3644 671
rect 3848 667 3852 671
rect 376 659 380 663
rect 536 659 540 663
rect 704 659 708 663
rect 872 659 876 663
rect 1040 659 1044 663
rect 1200 659 1204 663
rect 1360 659 1364 663
rect 1520 659 1524 663
rect 1672 659 1676 663
rect 1832 659 1836 663
rect 1968 659 1972 663
rect 360 647 364 651
rect 512 647 516 651
rect 680 647 684 651
rect 848 647 852 651
rect 1016 647 1020 651
rect 1176 647 1180 651
rect 1328 647 1332 651
rect 1464 647 1468 651
rect 1600 647 1604 651
rect 1728 647 1732 651
rect 1856 647 1860 651
rect 1968 647 1972 651
rect 2136 643 2140 647
rect 2304 643 2308 647
rect 2488 643 2492 647
rect 2688 643 2692 647
rect 2904 643 2908 647
rect 3136 643 3140 647
rect 3384 643 3388 647
rect 3640 643 3644 647
rect 3904 643 3908 647
rect 1520 511 1524 515
rect 304 503 308 507
rect 480 503 484 507
rect 672 503 676 507
rect 864 503 868 507
rect 1056 503 1060 507
rect 1240 503 1244 507
rect 1416 503 1420 507
rect 200 491 204 495
rect 352 491 356 495
rect 528 491 532 495
rect 704 491 708 495
rect 728 491 732 495
rect 872 491 876 495
rect 1032 491 1036 495
rect 1184 491 1188 495
rect 1336 491 1340 495
rect 1480 491 1484 495
rect 728 463 732 467
rect 1584 503 1588 507
rect 1752 503 1756 507
rect 1928 503 1932 507
rect 2256 503 2260 507
rect 2352 503 2356 507
rect 2448 503 2452 507
rect 2544 503 2548 507
rect 2648 503 2652 507
rect 2776 503 2780 507
rect 2936 503 2940 507
rect 3136 503 3140 507
rect 3368 503 3372 507
rect 3616 503 3620 507
rect 3872 503 3876 507
rect 1632 491 1636 495
rect 2496 491 2500 495
rect 2592 491 2596 495
rect 2688 491 2692 495
rect 2792 491 2796 495
rect 2912 491 2916 495
rect 3064 491 3068 495
rect 3240 491 3244 495
rect 3440 491 3444 495
rect 3656 491 3660 495
rect 3872 491 3876 495
rect 1520 463 1524 467
rect 2496 351 2500 355
rect 2592 351 2596 355
rect 2688 351 2692 355
rect 2784 351 2788 355
rect 2880 351 2884 355
rect 2992 351 2996 355
rect 3128 351 3132 355
rect 3288 351 3292 355
rect 3464 351 3468 355
rect 3656 351 3660 355
rect 3848 351 3852 355
rect 200 347 204 351
rect 344 347 348 351
rect 504 347 508 351
rect 648 347 652 351
rect 784 347 788 351
rect 912 347 916 351
rect 1032 347 1036 351
rect 1152 347 1156 351
rect 1272 347 1276 351
rect 1392 347 1396 351
rect 208 335 212 339
rect 232 335 236 339
rect 384 335 388 339
rect 544 335 548 339
rect 696 335 700 339
rect 840 335 844 339
rect 968 335 972 339
rect 1096 335 1100 339
rect 1216 335 1220 339
rect 1336 335 1340 339
rect 1456 335 1460 339
rect 2256 335 2260 339
rect 2392 335 2396 339
rect 2536 335 2540 339
rect 2688 335 2692 339
rect 2848 335 2852 339
rect 3016 335 3020 339
rect 3184 335 3188 339
rect 3360 335 3364 339
rect 3536 335 3540 339
rect 3720 335 3724 339
rect 3904 335 3908 339
rect 232 307 236 311
rect 896 223 900 227
rect 288 191 292 195
rect 456 191 460 195
rect 624 191 628 195
rect 800 191 804 195
rect 2136 195 2140 199
rect 2280 195 2284 199
rect 2464 195 2468 199
rect 2656 195 2660 199
rect 2856 195 2860 199
rect 3048 195 3052 199
rect 3232 195 3236 199
rect 3408 195 3412 199
rect 3576 195 3580 199
rect 3752 195 3756 199
rect 3904 195 3908 199
rect 968 191 972 195
rect 1128 191 1132 195
rect 1280 191 1284 195
rect 1424 191 1428 195
rect 1576 191 1580 195
rect 1728 191 1732 195
rect 2136 159 2140 163
rect 2160 159 2164 163
rect 2256 159 2260 163
rect 2408 159 2412 163
rect 2560 159 2564 163
rect 2712 159 2716 163
rect 2864 159 2868 163
rect 3008 159 3012 163
rect 3136 159 3140 163
rect 3256 159 3260 163
rect 3376 159 3380 163
rect 3488 159 3492 163
rect 3592 159 3596 163
rect 3704 159 3708 163
rect 3808 159 3812 163
rect 3904 159 3908 163
rect 216 147 220 151
rect 240 147 244 151
rect 312 147 316 151
rect 336 147 340 151
rect 408 147 412 151
rect 504 147 508 151
rect 600 147 604 151
rect 696 147 700 151
rect 792 147 796 151
rect 888 147 892 151
rect 896 147 900 151
rect 984 147 988 151
rect 1080 147 1084 151
rect 1176 147 1180 151
rect 1272 147 1276 151
rect 1368 147 1372 151
rect 1400 147 1404 151
rect 1472 147 1476 151
rect 1504 147 1508 151
rect 1576 147 1580 151
rect 1608 147 1612 151
rect 1680 147 1684 151
rect 1776 147 1780 151
rect 1872 147 1876 151
rect 1968 147 1972 151
rect 240 119 244 123
rect 336 119 340 123
rect 1400 119 1404 123
rect 1504 119 1508 123
rect 2160 131 2164 135
rect 1608 119 1612 123
<< m2 >>
rect 2070 3992 2076 3993
rect 2046 3989 2052 3990
rect 2046 3985 2047 3989
rect 2051 3985 2052 3989
rect 2070 3988 2071 3992
rect 2075 3988 2076 3992
rect 2070 3987 2076 3988
rect 2326 3992 2332 3993
rect 2326 3988 2327 3992
rect 2331 3988 2332 3992
rect 2326 3987 2332 3988
rect 2590 3992 2596 3993
rect 2590 3988 2591 3992
rect 2595 3988 2596 3992
rect 2590 3987 2596 3988
rect 2838 3992 2844 3993
rect 2838 3988 2839 3992
rect 2843 3988 2844 3992
rect 2838 3987 2844 3988
rect 3086 3992 3092 3993
rect 3086 3988 3087 3992
rect 3091 3988 3092 3992
rect 3086 3987 3092 3988
rect 3342 3992 3348 3993
rect 3342 3988 3343 3992
rect 3347 3988 3348 3992
rect 3342 3987 3348 3988
rect 3942 3989 3948 3990
rect 2046 3984 2052 3985
rect 3942 3985 3943 3989
rect 3947 3985 3948 3989
rect 3942 3984 3948 3985
rect 2146 3983 2152 3984
rect 2146 3979 2147 3983
rect 2151 3979 2152 3983
rect 2146 3978 2152 3979
rect 2194 3983 2200 3984
rect 2194 3979 2195 3983
rect 2199 3982 2200 3983
rect 2666 3983 2672 3984
rect 2199 3980 2369 3982
rect 2199 3979 2200 3980
rect 2194 3978 2200 3979
rect 2666 3979 2667 3983
rect 2671 3979 2672 3983
rect 2666 3978 2672 3979
rect 2914 3983 2920 3984
rect 2914 3979 2915 3983
rect 2919 3979 2920 3983
rect 2914 3978 2920 3979
rect 3162 3983 3168 3984
rect 3162 3979 3163 3983
rect 3167 3979 3168 3983
rect 3162 3978 3168 3979
rect 3242 3983 3248 3984
rect 3242 3979 3243 3983
rect 3247 3982 3248 3983
rect 3247 3980 3385 3982
rect 3247 3979 3248 3980
rect 3242 3978 3248 3979
rect 2070 3973 2076 3974
rect 310 3972 316 3973
rect 110 3969 116 3970
rect 110 3965 111 3969
rect 115 3965 116 3969
rect 310 3968 311 3972
rect 315 3968 316 3972
rect 310 3967 316 3968
rect 510 3972 516 3973
rect 510 3968 511 3972
rect 515 3968 516 3972
rect 510 3967 516 3968
rect 702 3972 708 3973
rect 702 3968 703 3972
rect 707 3968 708 3972
rect 702 3967 708 3968
rect 886 3972 892 3973
rect 886 3968 887 3972
rect 891 3968 892 3972
rect 886 3967 892 3968
rect 1062 3972 1068 3973
rect 1062 3968 1063 3972
rect 1067 3968 1068 3972
rect 1062 3967 1068 3968
rect 1230 3972 1236 3973
rect 1230 3968 1231 3972
rect 1235 3968 1236 3972
rect 1230 3967 1236 3968
rect 1382 3972 1388 3973
rect 1382 3968 1383 3972
rect 1387 3968 1388 3972
rect 1382 3967 1388 3968
rect 1518 3972 1524 3973
rect 1518 3968 1519 3972
rect 1523 3968 1524 3972
rect 1518 3967 1524 3968
rect 1654 3972 1660 3973
rect 1654 3968 1655 3972
rect 1659 3968 1660 3972
rect 1654 3967 1660 3968
rect 1790 3972 1796 3973
rect 1790 3968 1791 3972
rect 1795 3968 1796 3972
rect 1790 3967 1796 3968
rect 1902 3972 1908 3973
rect 1902 3968 1903 3972
rect 1907 3968 1908 3972
rect 2046 3972 2052 3973
rect 1902 3967 1908 3968
rect 2006 3969 2012 3970
rect 110 3964 116 3965
rect 2006 3965 2007 3969
rect 2011 3965 2012 3969
rect 2046 3968 2047 3972
rect 2051 3968 2052 3972
rect 2070 3969 2071 3973
rect 2075 3969 2076 3973
rect 2070 3968 2076 3969
rect 2326 3973 2332 3974
rect 2326 3969 2327 3973
rect 2331 3969 2332 3973
rect 2326 3968 2332 3969
rect 2590 3973 2596 3974
rect 2590 3969 2591 3973
rect 2595 3969 2596 3973
rect 2590 3968 2596 3969
rect 2838 3973 2844 3974
rect 2838 3969 2839 3973
rect 2843 3969 2844 3973
rect 2838 3968 2844 3969
rect 3086 3973 3092 3974
rect 3086 3969 3087 3973
rect 3091 3969 3092 3973
rect 3086 3968 3092 3969
rect 3342 3973 3348 3974
rect 3342 3969 3343 3973
rect 3347 3969 3348 3973
rect 3342 3968 3348 3969
rect 3942 3972 3948 3973
rect 3942 3968 3943 3972
rect 3947 3968 3948 3972
rect 2046 3967 2052 3968
rect 3942 3967 3948 3968
rect 2006 3964 2012 3965
rect 462 3963 468 3964
rect 462 3962 463 3963
rect 389 3960 463 3962
rect 462 3959 463 3960
rect 467 3959 468 3963
rect 462 3958 468 3959
rect 586 3963 592 3964
rect 586 3959 587 3963
rect 591 3959 592 3963
rect 586 3958 592 3959
rect 778 3963 784 3964
rect 778 3959 779 3963
rect 783 3959 784 3963
rect 1138 3963 1144 3964
rect 778 3958 784 3959
rect 788 3960 929 3962
rect 310 3953 316 3954
rect 110 3952 116 3953
rect 110 3948 111 3952
rect 115 3948 116 3952
rect 310 3949 311 3953
rect 315 3949 316 3953
rect 310 3948 316 3949
rect 510 3953 516 3954
rect 510 3949 511 3953
rect 515 3949 516 3953
rect 510 3948 516 3949
rect 702 3953 708 3954
rect 702 3949 703 3953
rect 707 3949 708 3953
rect 702 3948 708 3949
rect 110 3947 116 3948
rect 634 3947 640 3948
rect 634 3943 635 3947
rect 639 3946 640 3947
rect 788 3946 790 3960
rect 1138 3959 1139 3963
rect 1143 3959 1144 3963
rect 1138 3958 1144 3959
rect 1306 3963 1312 3964
rect 1306 3959 1307 3963
rect 1311 3959 1312 3963
rect 1306 3958 1312 3959
rect 1458 3963 1464 3964
rect 1458 3959 1459 3963
rect 1463 3959 1464 3963
rect 1458 3958 1464 3959
rect 1594 3963 1600 3964
rect 1594 3959 1595 3963
rect 1599 3959 1600 3963
rect 1594 3958 1600 3959
rect 1730 3963 1736 3964
rect 1730 3959 1731 3963
rect 1735 3959 1736 3963
rect 1730 3958 1736 3959
rect 1866 3963 1872 3964
rect 1866 3959 1867 3963
rect 1871 3959 1872 3963
rect 1981 3960 2001 3962
rect 1866 3958 1872 3959
rect 1999 3958 2001 3960
rect 1999 3956 2070 3958
rect 886 3953 892 3954
rect 886 3949 887 3953
rect 891 3949 892 3953
rect 886 3948 892 3949
rect 1062 3953 1068 3954
rect 1062 3949 1063 3953
rect 1067 3949 1068 3953
rect 1062 3948 1068 3949
rect 1230 3953 1236 3954
rect 1230 3949 1231 3953
rect 1235 3949 1236 3953
rect 1230 3948 1236 3949
rect 1382 3953 1388 3954
rect 1382 3949 1383 3953
rect 1387 3949 1388 3953
rect 1382 3948 1388 3949
rect 1518 3953 1524 3954
rect 1518 3949 1519 3953
rect 1523 3949 1524 3953
rect 1518 3948 1524 3949
rect 1654 3953 1660 3954
rect 1654 3949 1655 3953
rect 1659 3949 1660 3953
rect 1654 3948 1660 3949
rect 1790 3953 1796 3954
rect 1790 3949 1791 3953
rect 1795 3949 1796 3953
rect 1790 3948 1796 3949
rect 1902 3953 1908 3954
rect 1902 3949 1903 3953
rect 1907 3949 1908 3953
rect 1902 3948 1908 3949
rect 2006 3952 2012 3953
rect 2006 3948 2007 3952
rect 2011 3948 2012 3952
rect 2068 3950 2070 3956
rect 2135 3951 2141 3952
rect 2135 3950 2136 3951
rect 2068 3948 2136 3950
rect 2006 3947 2012 3948
rect 2135 3947 2136 3948
rect 2140 3947 2141 3951
rect 2135 3946 2141 3947
rect 2146 3951 2152 3952
rect 2146 3947 2147 3951
rect 2151 3950 2152 3951
rect 2391 3951 2397 3952
rect 2391 3950 2392 3951
rect 2151 3948 2392 3950
rect 2151 3947 2152 3948
rect 2146 3946 2152 3947
rect 2391 3947 2392 3948
rect 2396 3947 2397 3951
rect 2391 3946 2397 3947
rect 2655 3951 2664 3952
rect 2655 3947 2656 3951
rect 2663 3947 2664 3951
rect 2655 3946 2664 3947
rect 2666 3951 2672 3952
rect 2666 3947 2667 3951
rect 2671 3950 2672 3951
rect 2903 3951 2909 3952
rect 2903 3950 2904 3951
rect 2671 3948 2904 3950
rect 2671 3947 2672 3948
rect 2666 3946 2672 3947
rect 2903 3947 2904 3948
rect 2908 3947 2909 3951
rect 2903 3946 2909 3947
rect 2914 3951 2920 3952
rect 2914 3947 2915 3951
rect 2919 3950 2920 3951
rect 3151 3951 3157 3952
rect 3151 3950 3152 3951
rect 2919 3948 3152 3950
rect 2919 3947 2920 3948
rect 2914 3946 2920 3947
rect 3151 3947 3152 3948
rect 3156 3947 3157 3951
rect 3151 3946 3157 3947
rect 3162 3951 3168 3952
rect 3162 3947 3163 3951
rect 3167 3950 3168 3951
rect 3407 3951 3413 3952
rect 3407 3950 3408 3951
rect 3167 3948 3408 3950
rect 3167 3947 3168 3948
rect 3162 3946 3168 3947
rect 3407 3947 3408 3948
rect 3412 3947 3413 3951
rect 3407 3946 3413 3947
rect 639 3944 790 3946
rect 639 3943 640 3944
rect 634 3942 640 3943
rect 2191 3939 2200 3940
rect 2191 3935 2192 3939
rect 2199 3935 2200 3939
rect 2191 3934 2200 3935
rect 2202 3939 2208 3940
rect 2202 3935 2203 3939
rect 2207 3938 2208 3939
rect 2335 3939 2341 3940
rect 2335 3938 2336 3939
rect 2207 3936 2336 3938
rect 2207 3935 2208 3936
rect 2202 3934 2208 3935
rect 2335 3935 2336 3936
rect 2340 3935 2341 3939
rect 2335 3934 2341 3935
rect 2346 3939 2352 3940
rect 2346 3935 2347 3939
rect 2351 3938 2352 3939
rect 2503 3939 2509 3940
rect 2503 3938 2504 3939
rect 2351 3936 2504 3938
rect 2351 3935 2352 3936
rect 2346 3934 2352 3935
rect 2503 3935 2504 3936
rect 2508 3935 2509 3939
rect 2503 3934 2509 3935
rect 2514 3939 2520 3940
rect 2514 3935 2515 3939
rect 2519 3938 2520 3939
rect 2679 3939 2685 3940
rect 2679 3938 2680 3939
rect 2519 3936 2680 3938
rect 2519 3935 2520 3936
rect 2514 3934 2520 3935
rect 2679 3935 2680 3936
rect 2684 3935 2685 3939
rect 2679 3934 2685 3935
rect 2690 3939 2696 3940
rect 2690 3935 2691 3939
rect 2695 3938 2696 3939
rect 2863 3939 2869 3940
rect 2863 3938 2864 3939
rect 2695 3936 2864 3938
rect 2695 3935 2696 3936
rect 2690 3934 2696 3935
rect 2863 3935 2864 3936
rect 2868 3935 2869 3939
rect 2863 3934 2869 3935
rect 3047 3939 3056 3940
rect 3047 3935 3048 3939
rect 3055 3935 3056 3939
rect 3047 3934 3056 3935
rect 3239 3939 3248 3940
rect 3239 3935 3240 3939
rect 3247 3935 3248 3939
rect 3239 3934 3248 3935
rect 3250 3939 3256 3940
rect 3250 3935 3251 3939
rect 3255 3938 3256 3939
rect 3431 3939 3437 3940
rect 3431 3938 3432 3939
rect 3255 3936 3432 3938
rect 3255 3935 3256 3936
rect 3250 3934 3256 3935
rect 3431 3935 3432 3936
rect 3436 3935 3437 3939
rect 3431 3934 3437 3935
rect 3442 3939 3448 3940
rect 3442 3935 3443 3939
rect 3447 3938 3448 3939
rect 3623 3939 3629 3940
rect 3623 3938 3624 3939
rect 3447 3936 3624 3938
rect 3447 3935 3448 3936
rect 3442 3934 3448 3935
rect 3623 3935 3624 3936
rect 3628 3935 3629 3939
rect 3623 3934 3629 3935
rect 375 3931 381 3932
rect 375 3927 376 3931
rect 380 3930 381 3931
rect 402 3931 408 3932
rect 402 3930 403 3931
rect 380 3928 403 3930
rect 380 3927 381 3928
rect 375 3926 381 3927
rect 402 3927 403 3928
rect 407 3927 408 3931
rect 402 3926 408 3927
rect 462 3931 468 3932
rect 462 3927 463 3931
rect 467 3930 468 3931
rect 575 3931 581 3932
rect 575 3930 576 3931
rect 467 3928 576 3930
rect 467 3927 468 3928
rect 462 3926 468 3927
rect 575 3927 576 3928
rect 580 3927 581 3931
rect 575 3926 581 3927
rect 586 3931 592 3932
rect 586 3927 587 3931
rect 591 3930 592 3931
rect 767 3931 773 3932
rect 767 3930 768 3931
rect 591 3928 768 3930
rect 591 3927 592 3928
rect 586 3926 592 3927
rect 767 3927 768 3928
rect 772 3927 773 3931
rect 767 3926 773 3927
rect 778 3931 784 3932
rect 778 3927 779 3931
rect 783 3930 784 3931
rect 951 3931 957 3932
rect 951 3930 952 3931
rect 783 3928 952 3930
rect 783 3927 784 3928
rect 778 3926 784 3927
rect 951 3927 952 3928
rect 956 3927 957 3931
rect 951 3926 957 3927
rect 1127 3931 1136 3932
rect 1127 3927 1128 3931
rect 1135 3927 1136 3931
rect 1127 3926 1136 3927
rect 1138 3931 1144 3932
rect 1138 3927 1139 3931
rect 1143 3930 1144 3931
rect 1295 3931 1301 3932
rect 1295 3930 1296 3931
rect 1143 3928 1296 3930
rect 1143 3927 1144 3928
rect 1138 3926 1144 3927
rect 1295 3927 1296 3928
rect 1300 3927 1301 3931
rect 1295 3926 1301 3927
rect 1306 3931 1312 3932
rect 1306 3927 1307 3931
rect 1311 3930 1312 3931
rect 1447 3931 1453 3932
rect 1447 3930 1448 3931
rect 1311 3928 1448 3930
rect 1311 3927 1312 3928
rect 1306 3926 1312 3927
rect 1447 3927 1448 3928
rect 1452 3927 1453 3931
rect 1447 3926 1453 3927
rect 1458 3931 1464 3932
rect 1458 3927 1459 3931
rect 1463 3930 1464 3931
rect 1583 3931 1589 3932
rect 1583 3930 1584 3931
rect 1463 3928 1584 3930
rect 1463 3927 1464 3928
rect 1458 3926 1464 3927
rect 1583 3927 1584 3928
rect 1588 3927 1589 3931
rect 1583 3926 1589 3927
rect 1594 3931 1600 3932
rect 1594 3927 1595 3931
rect 1599 3930 1600 3931
rect 1719 3931 1725 3932
rect 1719 3930 1720 3931
rect 1599 3928 1720 3930
rect 1599 3927 1600 3928
rect 1594 3926 1600 3927
rect 1719 3927 1720 3928
rect 1724 3927 1725 3931
rect 1719 3926 1725 3927
rect 1730 3931 1736 3932
rect 1730 3927 1731 3931
rect 1735 3930 1736 3931
rect 1855 3931 1861 3932
rect 1855 3930 1856 3931
rect 1735 3928 1856 3930
rect 1735 3927 1736 3928
rect 1730 3926 1736 3927
rect 1855 3927 1856 3928
rect 1860 3927 1861 3931
rect 1855 3926 1861 3927
rect 1866 3931 1872 3932
rect 1866 3927 1867 3931
rect 1871 3930 1872 3931
rect 1967 3931 1973 3932
rect 1967 3930 1968 3931
rect 1871 3928 1968 3930
rect 1871 3927 1872 3928
rect 1866 3926 1872 3927
rect 1967 3927 1968 3928
rect 1972 3927 1973 3931
rect 1967 3926 1973 3927
rect 2658 3927 2664 3928
rect 2658 3923 2659 3927
rect 2663 3926 2664 3927
rect 2663 3924 2938 3926
rect 2663 3923 2664 3924
rect 2658 3922 2664 3923
rect 2046 3920 2052 3921
rect 302 3919 308 3920
rect 302 3915 303 3919
rect 307 3918 308 3919
rect 343 3919 349 3920
rect 343 3918 344 3919
rect 307 3916 344 3918
rect 307 3915 308 3916
rect 302 3914 308 3915
rect 343 3915 344 3916
rect 348 3915 349 3919
rect 343 3914 349 3915
rect 354 3919 360 3920
rect 354 3915 355 3919
rect 359 3918 360 3919
rect 479 3919 485 3920
rect 479 3918 480 3919
rect 359 3916 480 3918
rect 359 3915 360 3916
rect 354 3914 360 3915
rect 479 3915 480 3916
rect 484 3915 485 3919
rect 479 3914 485 3915
rect 631 3919 640 3920
rect 631 3915 632 3919
rect 639 3915 640 3919
rect 631 3914 640 3915
rect 642 3919 648 3920
rect 642 3915 643 3919
rect 647 3918 648 3919
rect 799 3919 805 3920
rect 799 3918 800 3919
rect 647 3916 800 3918
rect 647 3915 648 3916
rect 642 3914 648 3915
rect 799 3915 800 3916
rect 804 3915 805 3919
rect 799 3914 805 3915
rect 810 3919 816 3920
rect 810 3915 811 3919
rect 815 3918 816 3919
rect 975 3919 981 3920
rect 975 3918 976 3919
rect 815 3916 976 3918
rect 815 3915 816 3916
rect 810 3914 816 3915
rect 975 3915 976 3916
rect 980 3915 981 3919
rect 975 3914 981 3915
rect 986 3919 992 3920
rect 986 3915 987 3919
rect 991 3918 992 3919
rect 1159 3919 1165 3920
rect 1159 3918 1160 3919
rect 991 3916 1160 3918
rect 991 3915 992 3916
rect 986 3914 992 3915
rect 1159 3915 1160 3916
rect 1164 3915 1165 3919
rect 1159 3914 1165 3915
rect 1351 3919 1357 3920
rect 1351 3915 1352 3919
rect 1356 3918 1357 3919
rect 1370 3919 1376 3920
rect 1370 3918 1371 3919
rect 1356 3916 1371 3918
rect 1356 3915 1357 3916
rect 1351 3914 1357 3915
rect 1370 3915 1371 3916
rect 1375 3915 1376 3919
rect 1370 3914 1376 3915
rect 1543 3919 1549 3920
rect 1543 3915 1544 3919
rect 1548 3918 1549 3919
rect 1567 3919 1573 3920
rect 1567 3918 1568 3919
rect 1548 3916 1568 3918
rect 1548 3915 1549 3916
rect 1543 3914 1549 3915
rect 1567 3915 1568 3916
rect 1572 3915 1573 3919
rect 1567 3914 1573 3915
rect 1706 3919 1712 3920
rect 1706 3915 1707 3919
rect 1711 3918 1712 3919
rect 1743 3919 1749 3920
rect 1743 3918 1744 3919
rect 1711 3916 1744 3918
rect 1711 3915 1712 3916
rect 1706 3914 1712 3915
rect 1743 3915 1744 3916
rect 1748 3915 1749 3919
rect 2046 3916 2047 3920
rect 2051 3916 2052 3920
rect 2046 3915 2052 3916
rect 2126 3919 2132 3920
rect 2126 3915 2127 3919
rect 2131 3915 2132 3919
rect 1743 3914 1749 3915
rect 2126 3914 2132 3915
rect 2270 3919 2276 3920
rect 2270 3915 2271 3919
rect 2275 3915 2276 3919
rect 2270 3914 2276 3915
rect 2438 3919 2444 3920
rect 2438 3915 2439 3919
rect 2443 3915 2444 3919
rect 2438 3914 2444 3915
rect 2614 3919 2620 3920
rect 2614 3915 2615 3919
rect 2619 3915 2620 3919
rect 2614 3914 2620 3915
rect 2798 3919 2804 3920
rect 2798 3915 2799 3919
rect 2803 3915 2804 3919
rect 2798 3914 2804 3915
rect 2202 3911 2208 3912
rect 1130 3907 1136 3908
rect 1130 3903 1131 3907
rect 1135 3906 1136 3907
rect 2202 3907 2203 3911
rect 2207 3907 2208 3911
rect 2202 3906 2208 3907
rect 2346 3911 2352 3912
rect 2346 3907 2347 3911
rect 2351 3907 2352 3911
rect 2346 3906 2352 3907
rect 2514 3911 2520 3912
rect 2514 3907 2515 3911
rect 2519 3907 2520 3911
rect 2514 3906 2520 3907
rect 2690 3911 2696 3912
rect 2690 3907 2691 3911
rect 2695 3907 2696 3911
rect 2936 3910 2938 3924
rect 3942 3920 3948 3921
rect 2982 3919 2988 3920
rect 2982 3915 2983 3919
rect 2987 3915 2988 3919
rect 2982 3914 2988 3915
rect 3174 3919 3180 3920
rect 3174 3915 3175 3919
rect 3179 3915 3180 3919
rect 3174 3914 3180 3915
rect 3366 3919 3372 3920
rect 3366 3915 3367 3919
rect 3371 3915 3372 3919
rect 3366 3914 3372 3915
rect 3558 3919 3564 3920
rect 3558 3915 3559 3919
rect 3563 3915 3564 3919
rect 3942 3916 3943 3920
rect 3947 3916 3948 3920
rect 3942 3915 3948 3916
rect 3558 3914 3564 3915
rect 3250 3911 3256 3912
rect 2936 3908 3025 3910
rect 2690 3906 2696 3907
rect 2874 3907 2880 3908
rect 1135 3904 1246 3906
rect 1135 3903 1136 3904
rect 1130 3902 1136 3903
rect 110 3900 116 3901
rect 110 3896 111 3900
rect 115 3896 116 3900
rect 110 3895 116 3896
rect 278 3899 284 3900
rect 278 3895 279 3899
rect 283 3895 284 3899
rect 278 3894 284 3895
rect 414 3899 420 3900
rect 414 3895 415 3899
rect 419 3895 420 3899
rect 414 3894 420 3895
rect 566 3899 572 3900
rect 566 3895 567 3899
rect 571 3895 572 3899
rect 566 3894 572 3895
rect 734 3899 740 3900
rect 734 3895 735 3899
rect 739 3895 740 3899
rect 734 3894 740 3895
rect 910 3899 916 3900
rect 910 3895 911 3899
rect 915 3895 916 3899
rect 910 3894 916 3895
rect 1094 3899 1100 3900
rect 1094 3895 1095 3899
rect 1099 3895 1100 3899
rect 1094 3894 1100 3895
rect 354 3891 360 3892
rect 354 3887 355 3891
rect 359 3887 360 3891
rect 354 3886 360 3887
rect 402 3891 408 3892
rect 402 3887 403 3891
rect 407 3890 408 3891
rect 642 3891 648 3892
rect 407 3888 457 3890
rect 407 3887 408 3888
rect 402 3886 408 3887
rect 642 3887 643 3891
rect 647 3887 648 3891
rect 642 3886 648 3887
rect 810 3891 816 3892
rect 810 3887 811 3891
rect 815 3887 816 3891
rect 810 3886 816 3887
rect 986 3891 992 3892
rect 986 3887 987 3891
rect 991 3887 992 3891
rect 986 3886 992 3887
rect 1046 3891 1052 3892
rect 1046 3887 1047 3891
rect 1051 3890 1052 3891
rect 1244 3890 1246 3904
rect 2046 3903 2052 3904
rect 2006 3900 2012 3901
rect 1286 3899 1292 3900
rect 1286 3895 1287 3899
rect 1291 3895 1292 3899
rect 1286 3894 1292 3895
rect 1478 3899 1484 3900
rect 1478 3895 1479 3899
rect 1483 3895 1484 3899
rect 1478 3894 1484 3895
rect 1678 3899 1684 3900
rect 1678 3895 1679 3899
rect 1683 3895 1684 3899
rect 2006 3896 2007 3900
rect 2011 3896 2012 3900
rect 2046 3899 2047 3903
rect 2051 3899 2052 3903
rect 2874 3903 2875 3907
rect 2879 3903 2880 3907
rect 3250 3907 3251 3911
rect 3255 3907 3256 3911
rect 3250 3906 3256 3907
rect 3442 3911 3448 3912
rect 3442 3907 3443 3911
rect 3447 3907 3448 3911
rect 3442 3906 3448 3907
rect 3538 3911 3544 3912
rect 3538 3907 3539 3911
rect 3543 3910 3544 3911
rect 3543 3908 3601 3910
rect 3543 3907 3544 3908
rect 3538 3906 3544 3907
rect 2874 3902 2880 3903
rect 3942 3903 3948 3904
rect 2046 3898 2052 3899
rect 2126 3900 2132 3901
rect 2006 3895 2012 3896
rect 2126 3896 2127 3900
rect 2131 3896 2132 3900
rect 2126 3895 2132 3896
rect 2270 3900 2276 3901
rect 2270 3896 2271 3900
rect 2275 3896 2276 3900
rect 2270 3895 2276 3896
rect 2438 3900 2444 3901
rect 2438 3896 2439 3900
rect 2443 3896 2444 3900
rect 2438 3895 2444 3896
rect 2614 3900 2620 3901
rect 2614 3896 2615 3900
rect 2619 3896 2620 3900
rect 2614 3895 2620 3896
rect 2798 3900 2804 3901
rect 2798 3896 2799 3900
rect 2803 3896 2804 3900
rect 2798 3895 2804 3896
rect 2982 3900 2988 3901
rect 2982 3896 2983 3900
rect 2987 3896 2988 3900
rect 2982 3895 2988 3896
rect 3174 3900 3180 3901
rect 3174 3896 3175 3900
rect 3179 3896 3180 3900
rect 3174 3895 3180 3896
rect 3366 3900 3372 3901
rect 3366 3896 3367 3900
rect 3371 3896 3372 3900
rect 3366 3895 3372 3896
rect 3558 3900 3564 3901
rect 3558 3896 3559 3900
rect 3563 3896 3564 3900
rect 3942 3899 3943 3903
rect 3947 3899 3948 3903
rect 3942 3898 3948 3899
rect 3558 3895 3564 3896
rect 1678 3894 1684 3895
rect 1370 3891 1376 3892
rect 1051 3888 1137 3890
rect 1244 3888 1329 3890
rect 1051 3887 1052 3888
rect 1046 3886 1052 3887
rect 1370 3887 1371 3891
rect 1375 3890 1376 3891
rect 1567 3891 1573 3892
rect 1375 3888 1521 3890
rect 1375 3887 1376 3888
rect 1370 3886 1376 3887
rect 1567 3887 1568 3891
rect 1572 3890 1573 3891
rect 1572 3888 1721 3890
rect 1572 3887 1573 3888
rect 1567 3886 1573 3887
rect 110 3883 116 3884
rect 110 3879 111 3883
rect 115 3879 116 3883
rect 2006 3883 2012 3884
rect 110 3878 116 3879
rect 278 3880 284 3881
rect 278 3876 279 3880
rect 283 3876 284 3880
rect 278 3875 284 3876
rect 414 3880 420 3881
rect 414 3876 415 3880
rect 419 3876 420 3880
rect 414 3875 420 3876
rect 566 3880 572 3881
rect 566 3876 567 3880
rect 571 3876 572 3880
rect 566 3875 572 3876
rect 734 3880 740 3881
rect 734 3876 735 3880
rect 739 3876 740 3880
rect 734 3875 740 3876
rect 910 3880 916 3881
rect 910 3876 911 3880
rect 915 3876 916 3880
rect 910 3875 916 3876
rect 1094 3880 1100 3881
rect 1094 3876 1095 3880
rect 1099 3876 1100 3880
rect 1094 3875 1100 3876
rect 1286 3880 1292 3881
rect 1286 3876 1287 3880
rect 1291 3876 1292 3880
rect 1286 3875 1292 3876
rect 1478 3880 1484 3881
rect 1478 3876 1479 3880
rect 1483 3876 1484 3880
rect 1478 3875 1484 3876
rect 1678 3880 1684 3881
rect 1678 3876 1679 3880
rect 1683 3876 1684 3880
rect 2006 3879 2007 3883
rect 2011 3879 2012 3883
rect 2006 3878 2012 3879
rect 1678 3875 1684 3876
rect 2262 3840 2268 3841
rect 2046 3837 2052 3838
rect 2046 3833 2047 3837
rect 2051 3833 2052 3837
rect 2262 3836 2263 3840
rect 2267 3836 2268 3840
rect 2262 3835 2268 3836
rect 2374 3840 2380 3841
rect 2374 3836 2375 3840
rect 2379 3836 2380 3840
rect 2374 3835 2380 3836
rect 2494 3840 2500 3841
rect 2494 3836 2495 3840
rect 2499 3836 2500 3840
rect 2494 3835 2500 3836
rect 2630 3840 2636 3841
rect 2630 3836 2631 3840
rect 2635 3836 2636 3840
rect 2630 3835 2636 3836
rect 2774 3840 2780 3841
rect 2774 3836 2775 3840
rect 2779 3836 2780 3840
rect 2774 3835 2780 3836
rect 2918 3840 2924 3841
rect 2918 3836 2919 3840
rect 2923 3836 2924 3840
rect 2918 3835 2924 3836
rect 3062 3840 3068 3841
rect 3062 3836 3063 3840
rect 3067 3836 3068 3840
rect 3062 3835 3068 3836
rect 3206 3840 3212 3841
rect 3206 3836 3207 3840
rect 3211 3836 3212 3840
rect 3206 3835 3212 3836
rect 3342 3840 3348 3841
rect 3342 3836 3343 3840
rect 3347 3836 3348 3840
rect 3342 3835 3348 3836
rect 3470 3840 3476 3841
rect 3470 3836 3471 3840
rect 3475 3836 3476 3840
rect 3470 3835 3476 3836
rect 3598 3840 3604 3841
rect 3598 3836 3599 3840
rect 3603 3836 3604 3840
rect 3598 3835 3604 3836
rect 3726 3840 3732 3841
rect 3726 3836 3727 3840
rect 3731 3836 3732 3840
rect 3726 3835 3732 3836
rect 3838 3840 3844 3841
rect 3838 3836 3839 3840
rect 3843 3836 3844 3840
rect 3838 3835 3844 3836
rect 3942 3837 3948 3838
rect 2046 3832 2052 3833
rect 3942 3833 3943 3837
rect 3947 3833 3948 3837
rect 3942 3832 3948 3833
rect 2338 3831 2344 3832
rect 2338 3827 2339 3831
rect 2343 3827 2344 3831
rect 2338 3826 2344 3827
rect 2450 3831 2456 3832
rect 2450 3827 2451 3831
rect 2455 3827 2456 3831
rect 2450 3826 2456 3827
rect 2458 3831 2464 3832
rect 2458 3827 2459 3831
rect 2463 3830 2464 3831
rect 2578 3831 2584 3832
rect 2463 3828 2537 3830
rect 2463 3827 2464 3828
rect 2458 3826 2464 3827
rect 2578 3827 2579 3831
rect 2583 3830 2584 3831
rect 2714 3831 2720 3832
rect 2583 3828 2673 3830
rect 2583 3827 2584 3828
rect 2578 3826 2584 3827
rect 2714 3827 2715 3831
rect 2719 3830 2720 3831
rect 2994 3831 3000 3832
rect 2719 3828 2817 3830
rect 2719 3827 2720 3828
rect 2714 3826 2720 3827
rect 2994 3827 2995 3831
rect 2999 3827 3000 3831
rect 2994 3826 3000 3827
rect 3050 3831 3056 3832
rect 3050 3827 3051 3831
rect 3055 3830 3056 3831
rect 3274 3831 3280 3832
rect 3055 3828 3105 3830
rect 3055 3827 3056 3828
rect 3050 3826 3056 3827
rect 3274 3827 3275 3831
rect 3279 3827 3280 3831
rect 3274 3826 3280 3827
rect 3290 3831 3296 3832
rect 3290 3827 3291 3831
rect 3295 3830 3296 3831
rect 3426 3831 3432 3832
rect 3295 3828 3385 3830
rect 3295 3827 3296 3828
rect 3290 3826 3296 3827
rect 3426 3827 3427 3831
rect 3431 3830 3432 3831
rect 3674 3831 3680 3832
rect 3431 3828 3513 3830
rect 3431 3827 3432 3828
rect 3426 3826 3432 3827
rect 3674 3827 3675 3831
rect 3679 3827 3680 3831
rect 3674 3826 3680 3827
rect 3802 3831 3808 3832
rect 3802 3827 3803 3831
rect 3807 3827 3808 3831
rect 3802 3826 3808 3827
rect 3906 3831 3912 3832
rect 3906 3827 3907 3831
rect 3911 3827 3912 3831
rect 3906 3826 3912 3827
rect 2262 3821 2268 3822
rect 2046 3820 2052 3821
rect 2046 3816 2047 3820
rect 2051 3816 2052 3820
rect 2262 3817 2263 3821
rect 2267 3817 2268 3821
rect 2262 3816 2268 3817
rect 2374 3821 2380 3822
rect 2374 3817 2375 3821
rect 2379 3817 2380 3821
rect 2374 3816 2380 3817
rect 2494 3821 2500 3822
rect 2494 3817 2495 3821
rect 2499 3817 2500 3821
rect 2494 3816 2500 3817
rect 2630 3821 2636 3822
rect 2630 3817 2631 3821
rect 2635 3817 2636 3821
rect 2630 3816 2636 3817
rect 2774 3821 2780 3822
rect 2774 3817 2775 3821
rect 2779 3817 2780 3821
rect 2774 3816 2780 3817
rect 2918 3821 2924 3822
rect 2918 3817 2919 3821
rect 2923 3817 2924 3821
rect 2918 3816 2924 3817
rect 3062 3821 3068 3822
rect 3062 3817 3063 3821
rect 3067 3817 3068 3821
rect 3062 3816 3068 3817
rect 3206 3821 3212 3822
rect 3206 3817 3207 3821
rect 3211 3817 3212 3821
rect 3206 3816 3212 3817
rect 3342 3821 3348 3822
rect 3342 3817 3343 3821
rect 3347 3817 3348 3821
rect 3342 3816 3348 3817
rect 3470 3821 3476 3822
rect 3470 3817 3471 3821
rect 3475 3817 3476 3821
rect 3470 3816 3476 3817
rect 3598 3821 3604 3822
rect 3598 3817 3599 3821
rect 3603 3817 3604 3821
rect 3598 3816 3604 3817
rect 3726 3821 3732 3822
rect 3726 3817 3727 3821
rect 3731 3817 3732 3821
rect 3726 3816 3732 3817
rect 3838 3821 3844 3822
rect 3838 3817 3839 3821
rect 3843 3817 3844 3821
rect 3838 3816 3844 3817
rect 3942 3820 3948 3821
rect 3942 3816 3943 3820
rect 3947 3816 3948 3820
rect 2046 3815 2052 3816
rect 3942 3815 3948 3816
rect 230 3812 236 3813
rect 110 3809 116 3810
rect 110 3805 111 3809
rect 115 3805 116 3809
rect 230 3808 231 3812
rect 235 3808 236 3812
rect 230 3807 236 3808
rect 334 3812 340 3813
rect 334 3808 335 3812
rect 339 3808 340 3812
rect 334 3807 340 3808
rect 438 3812 444 3813
rect 438 3808 439 3812
rect 443 3808 444 3812
rect 438 3807 444 3808
rect 534 3812 540 3813
rect 534 3808 535 3812
rect 539 3808 540 3812
rect 534 3807 540 3808
rect 630 3812 636 3813
rect 630 3808 631 3812
rect 635 3808 636 3812
rect 630 3807 636 3808
rect 726 3812 732 3813
rect 726 3808 727 3812
rect 731 3808 732 3812
rect 726 3807 732 3808
rect 830 3812 836 3813
rect 830 3808 831 3812
rect 835 3808 836 3812
rect 830 3807 836 3808
rect 934 3812 940 3813
rect 934 3808 935 3812
rect 939 3808 940 3812
rect 934 3807 940 3808
rect 1038 3812 1044 3813
rect 1038 3808 1039 3812
rect 1043 3808 1044 3812
rect 1038 3807 1044 3808
rect 1150 3812 1156 3813
rect 1150 3808 1151 3812
rect 1155 3808 1156 3812
rect 1150 3807 1156 3808
rect 1262 3812 1268 3813
rect 1262 3808 1263 3812
rect 1267 3808 1268 3812
rect 1262 3807 1268 3808
rect 1382 3812 1388 3813
rect 1382 3808 1383 3812
rect 1387 3808 1388 3812
rect 1382 3807 1388 3808
rect 1502 3812 1508 3813
rect 1502 3808 1503 3812
rect 1507 3808 1508 3812
rect 1502 3807 1508 3808
rect 1630 3812 1636 3813
rect 1630 3808 1631 3812
rect 1635 3808 1636 3812
rect 1630 3807 1636 3808
rect 2006 3809 2012 3810
rect 110 3804 116 3805
rect 2006 3805 2007 3809
rect 2011 3805 2012 3809
rect 2458 3807 2464 3808
rect 2458 3806 2459 3807
rect 2006 3804 2012 3805
rect 2332 3804 2459 3806
rect 302 3803 308 3804
rect 302 3799 303 3803
rect 307 3799 308 3803
rect 302 3798 308 3799
rect 314 3803 320 3804
rect 314 3799 315 3803
rect 319 3802 320 3803
rect 514 3803 520 3804
rect 319 3800 377 3802
rect 319 3799 320 3800
rect 314 3798 320 3799
rect 514 3799 515 3803
rect 519 3799 520 3803
rect 514 3798 520 3799
rect 610 3803 616 3804
rect 610 3799 611 3803
rect 615 3799 616 3803
rect 610 3798 616 3799
rect 706 3803 712 3804
rect 706 3799 707 3803
rect 711 3799 712 3803
rect 706 3798 712 3799
rect 802 3803 808 3804
rect 802 3799 803 3803
rect 807 3799 808 3803
rect 802 3798 808 3799
rect 906 3803 912 3804
rect 906 3799 907 3803
rect 911 3799 912 3803
rect 906 3798 912 3799
rect 1010 3803 1016 3804
rect 1010 3799 1011 3803
rect 1015 3799 1016 3803
rect 1010 3798 1016 3799
rect 1114 3803 1120 3804
rect 1114 3799 1115 3803
rect 1119 3799 1120 3803
rect 1114 3798 1120 3799
rect 1226 3803 1232 3804
rect 1226 3799 1227 3803
rect 1231 3799 1232 3803
rect 1226 3798 1232 3799
rect 1338 3803 1344 3804
rect 1338 3799 1339 3803
rect 1343 3799 1344 3803
rect 1618 3803 1624 3804
rect 1618 3802 1619 3803
rect 1338 3798 1344 3799
rect 1348 3800 1425 3802
rect 1581 3800 1619 3802
rect 230 3793 236 3794
rect 110 3792 116 3793
rect 110 3788 111 3792
rect 115 3788 116 3792
rect 230 3789 231 3793
rect 235 3789 236 3793
rect 230 3788 236 3789
rect 334 3793 340 3794
rect 334 3789 335 3793
rect 339 3789 340 3793
rect 334 3788 340 3789
rect 438 3793 444 3794
rect 438 3789 439 3793
rect 443 3789 444 3793
rect 438 3788 444 3789
rect 534 3793 540 3794
rect 534 3789 535 3793
rect 539 3789 540 3793
rect 534 3788 540 3789
rect 630 3793 636 3794
rect 630 3789 631 3793
rect 635 3789 636 3793
rect 630 3788 636 3789
rect 726 3793 732 3794
rect 726 3789 727 3793
rect 731 3789 732 3793
rect 726 3788 732 3789
rect 830 3793 836 3794
rect 830 3789 831 3793
rect 835 3789 836 3793
rect 830 3788 836 3789
rect 934 3793 940 3794
rect 934 3789 935 3793
rect 939 3789 940 3793
rect 934 3788 940 3789
rect 1038 3793 1044 3794
rect 1038 3789 1039 3793
rect 1043 3789 1044 3793
rect 1038 3788 1044 3789
rect 1150 3793 1156 3794
rect 1150 3789 1151 3793
rect 1155 3789 1156 3793
rect 1150 3788 1156 3789
rect 1262 3793 1268 3794
rect 1262 3789 1263 3793
rect 1267 3789 1268 3793
rect 1262 3788 1268 3789
rect 110 3787 116 3788
rect 818 3787 824 3788
rect 818 3783 819 3787
rect 823 3786 824 3787
rect 1348 3786 1350 3800
rect 1618 3799 1619 3800
rect 1623 3799 1624 3803
rect 1618 3798 1624 3799
rect 1706 3803 1712 3804
rect 1706 3799 1707 3803
rect 1711 3799 1712 3803
rect 2332 3800 2334 3804
rect 2458 3803 2459 3804
rect 2463 3803 2464 3807
rect 2458 3802 2464 3803
rect 3674 3807 3680 3808
rect 3674 3803 3675 3807
rect 3679 3806 3680 3807
rect 3679 3803 3681 3806
rect 3674 3802 3681 3803
rect 1706 3798 1712 3799
rect 2327 3799 2334 3800
rect 2327 3795 2328 3799
rect 2332 3796 2334 3799
rect 2338 3799 2344 3800
rect 2332 3795 2333 3796
rect 2327 3794 2333 3795
rect 2338 3795 2339 3799
rect 2343 3798 2344 3799
rect 2439 3799 2445 3800
rect 2439 3798 2440 3799
rect 2343 3796 2440 3798
rect 2343 3795 2344 3796
rect 2338 3794 2344 3795
rect 2439 3795 2440 3796
rect 2444 3795 2445 3799
rect 2439 3794 2445 3795
rect 2559 3799 2565 3800
rect 2559 3795 2560 3799
rect 2564 3798 2565 3799
rect 2578 3799 2584 3800
rect 2578 3798 2579 3799
rect 2564 3796 2579 3798
rect 2564 3795 2565 3796
rect 2559 3794 2565 3795
rect 2578 3795 2579 3796
rect 2583 3795 2584 3799
rect 2578 3794 2584 3795
rect 2695 3799 2701 3800
rect 2695 3795 2696 3799
rect 2700 3798 2701 3799
rect 2714 3799 2720 3800
rect 2714 3798 2715 3799
rect 2700 3796 2715 3798
rect 2700 3795 2701 3796
rect 2695 3794 2701 3795
rect 2714 3795 2715 3796
rect 2719 3795 2720 3799
rect 2714 3794 2720 3795
rect 2839 3799 2845 3800
rect 2839 3795 2840 3799
rect 2844 3798 2845 3799
rect 2874 3799 2880 3800
rect 2874 3798 2875 3799
rect 2844 3796 2875 3798
rect 2844 3795 2845 3796
rect 2839 3794 2845 3795
rect 2874 3795 2875 3796
rect 2879 3795 2880 3799
rect 2874 3794 2880 3795
rect 2882 3799 2888 3800
rect 2882 3795 2883 3799
rect 2887 3798 2888 3799
rect 2983 3799 2989 3800
rect 2983 3798 2984 3799
rect 2887 3796 2984 3798
rect 2887 3795 2888 3796
rect 2882 3794 2888 3795
rect 2983 3795 2984 3796
rect 2988 3795 2989 3799
rect 2983 3794 2989 3795
rect 2994 3799 3000 3800
rect 2994 3795 2995 3799
rect 2999 3798 3000 3799
rect 3127 3799 3133 3800
rect 3127 3798 3128 3799
rect 2999 3796 3128 3798
rect 2999 3795 3000 3796
rect 2994 3794 3000 3795
rect 3127 3795 3128 3796
rect 3132 3795 3133 3799
rect 3127 3794 3133 3795
rect 3271 3799 3277 3800
rect 3271 3795 3272 3799
rect 3276 3798 3277 3799
rect 3290 3799 3296 3800
rect 3290 3798 3291 3799
rect 3276 3796 3291 3798
rect 3276 3795 3277 3796
rect 3271 3794 3277 3795
rect 3290 3795 3291 3796
rect 3295 3795 3296 3799
rect 3290 3794 3296 3795
rect 3407 3799 3413 3800
rect 3407 3795 3408 3799
rect 3412 3798 3413 3799
rect 3426 3799 3432 3800
rect 3426 3798 3427 3799
rect 3412 3796 3427 3798
rect 3412 3795 3413 3796
rect 3407 3794 3413 3795
rect 3426 3795 3427 3796
rect 3431 3795 3432 3799
rect 3426 3794 3432 3795
rect 3535 3799 3544 3800
rect 3535 3795 3536 3799
rect 3543 3795 3544 3799
rect 3535 3794 3544 3795
rect 3663 3799 3669 3800
rect 3663 3795 3664 3799
rect 3668 3798 3669 3799
rect 3671 3799 3677 3800
rect 3671 3798 3672 3799
rect 3668 3796 3672 3798
rect 3668 3795 3669 3796
rect 3663 3794 3669 3795
rect 3671 3795 3672 3796
rect 3676 3795 3677 3799
rect 3679 3798 3681 3802
rect 3791 3799 3797 3800
rect 3791 3798 3792 3799
rect 3679 3796 3792 3798
rect 3671 3794 3677 3795
rect 3791 3795 3792 3796
rect 3796 3795 3797 3799
rect 3791 3794 3797 3795
rect 3802 3799 3808 3800
rect 3802 3795 3803 3799
rect 3807 3798 3808 3799
rect 3903 3799 3909 3800
rect 3903 3798 3904 3799
rect 3807 3796 3904 3798
rect 3807 3795 3808 3796
rect 3802 3794 3808 3795
rect 3903 3795 3904 3796
rect 3908 3795 3909 3799
rect 3903 3794 3909 3795
rect 1382 3793 1388 3794
rect 1382 3789 1383 3793
rect 1387 3789 1388 3793
rect 1382 3788 1388 3789
rect 1502 3793 1508 3794
rect 1502 3789 1503 3793
rect 1507 3789 1508 3793
rect 1502 3788 1508 3789
rect 1630 3793 1636 3794
rect 1630 3789 1631 3793
rect 1635 3789 1636 3793
rect 1630 3788 1636 3789
rect 2006 3792 2012 3793
rect 2006 3788 2007 3792
rect 2011 3788 2012 3792
rect 2006 3787 2012 3788
rect 823 3784 1350 3786
rect 823 3783 824 3784
rect 818 3782 824 3783
rect 1046 3779 1052 3780
rect 1046 3778 1047 3779
rect 508 3776 1047 3778
rect 508 3772 510 3776
rect 1046 3775 1047 3776
rect 1051 3775 1052 3779
rect 1046 3774 1052 3775
rect 295 3771 301 3772
rect 295 3767 296 3771
rect 300 3770 301 3771
rect 314 3771 320 3772
rect 314 3770 315 3771
rect 300 3768 315 3770
rect 300 3767 301 3768
rect 295 3766 301 3767
rect 314 3767 315 3768
rect 319 3767 320 3771
rect 314 3766 320 3767
rect 399 3771 405 3772
rect 399 3767 400 3771
rect 404 3770 405 3771
rect 447 3771 453 3772
rect 447 3770 448 3771
rect 404 3768 448 3770
rect 404 3767 405 3768
rect 399 3766 405 3767
rect 447 3767 448 3768
rect 452 3767 453 3771
rect 447 3766 453 3767
rect 503 3771 510 3772
rect 503 3767 504 3771
rect 508 3768 510 3771
rect 514 3771 520 3772
rect 508 3767 509 3768
rect 503 3766 509 3767
rect 514 3767 515 3771
rect 519 3770 520 3771
rect 599 3771 605 3772
rect 599 3770 600 3771
rect 519 3768 600 3770
rect 519 3767 520 3768
rect 514 3766 520 3767
rect 599 3767 600 3768
rect 604 3767 605 3771
rect 599 3766 605 3767
rect 610 3771 616 3772
rect 610 3767 611 3771
rect 615 3770 616 3771
rect 695 3771 701 3772
rect 695 3770 696 3771
rect 615 3768 696 3770
rect 615 3767 616 3768
rect 610 3766 616 3767
rect 695 3767 696 3768
rect 700 3767 701 3771
rect 695 3766 701 3767
rect 706 3771 712 3772
rect 706 3767 707 3771
rect 711 3770 712 3771
rect 791 3771 797 3772
rect 791 3770 792 3771
rect 711 3768 792 3770
rect 711 3767 712 3768
rect 706 3766 712 3767
rect 791 3767 792 3768
rect 796 3767 797 3771
rect 791 3766 797 3767
rect 802 3771 808 3772
rect 802 3767 803 3771
rect 807 3770 808 3771
rect 895 3771 901 3772
rect 895 3770 896 3771
rect 807 3768 896 3770
rect 807 3767 808 3768
rect 802 3766 808 3767
rect 895 3767 896 3768
rect 900 3767 901 3771
rect 895 3766 901 3767
rect 906 3771 912 3772
rect 906 3767 907 3771
rect 911 3770 912 3771
rect 999 3771 1005 3772
rect 999 3770 1000 3771
rect 911 3768 1000 3770
rect 911 3767 912 3768
rect 906 3766 912 3767
rect 999 3767 1000 3768
rect 1004 3767 1005 3771
rect 999 3766 1005 3767
rect 1010 3771 1016 3772
rect 1010 3767 1011 3771
rect 1015 3770 1016 3771
rect 1103 3771 1109 3772
rect 1103 3770 1104 3771
rect 1015 3768 1104 3770
rect 1015 3767 1016 3768
rect 1010 3766 1016 3767
rect 1103 3767 1104 3768
rect 1108 3767 1109 3771
rect 1103 3766 1109 3767
rect 1114 3771 1120 3772
rect 1114 3767 1115 3771
rect 1119 3770 1120 3771
rect 1215 3771 1221 3772
rect 1215 3770 1216 3771
rect 1119 3768 1216 3770
rect 1119 3767 1120 3768
rect 1114 3766 1120 3767
rect 1215 3767 1216 3768
rect 1220 3767 1221 3771
rect 1215 3766 1221 3767
rect 1226 3771 1232 3772
rect 1226 3767 1227 3771
rect 1231 3770 1232 3771
rect 1327 3771 1333 3772
rect 1327 3770 1328 3771
rect 1231 3768 1328 3770
rect 1231 3767 1232 3768
rect 1226 3766 1232 3767
rect 1327 3767 1328 3768
rect 1332 3767 1333 3771
rect 1327 3766 1333 3767
rect 1338 3771 1344 3772
rect 1338 3767 1339 3771
rect 1343 3770 1344 3771
rect 1447 3771 1453 3772
rect 1447 3770 1448 3771
rect 1343 3768 1448 3770
rect 1343 3767 1344 3768
rect 1338 3766 1344 3767
rect 1447 3767 1448 3768
rect 1452 3767 1453 3771
rect 1447 3766 1453 3767
rect 1567 3771 1573 3772
rect 1567 3767 1568 3771
rect 1572 3770 1573 3771
rect 1599 3771 1605 3772
rect 1599 3770 1600 3771
rect 1572 3768 1600 3770
rect 1572 3767 1573 3768
rect 1567 3766 1573 3767
rect 1599 3767 1600 3768
rect 1604 3767 1605 3771
rect 1599 3766 1605 3767
rect 1618 3771 1624 3772
rect 1618 3767 1619 3771
rect 1623 3770 1624 3771
rect 1695 3771 1701 3772
rect 1695 3770 1696 3771
rect 1623 3768 1696 3770
rect 1623 3767 1624 3768
rect 1618 3766 1624 3767
rect 1695 3767 1696 3768
rect 1700 3767 1701 3771
rect 1695 3766 1701 3767
rect 2135 3771 2141 3772
rect 2135 3767 2136 3771
rect 2140 3770 2141 3771
rect 2154 3771 2160 3772
rect 2154 3770 2155 3771
rect 2140 3768 2155 3770
rect 2140 3767 2141 3768
rect 2135 3766 2141 3767
rect 2154 3767 2155 3768
rect 2159 3767 2160 3771
rect 2154 3766 2160 3767
rect 2247 3771 2253 3772
rect 2247 3767 2248 3771
rect 2252 3770 2253 3771
rect 2271 3771 2277 3772
rect 2271 3770 2272 3771
rect 2252 3768 2272 3770
rect 2252 3767 2253 3768
rect 2247 3766 2253 3767
rect 2271 3767 2272 3768
rect 2276 3767 2277 3771
rect 2271 3766 2277 3767
rect 2391 3771 2397 3772
rect 2391 3767 2392 3771
rect 2396 3770 2397 3771
rect 2450 3771 2456 3772
rect 2396 3768 2446 3770
rect 2396 3767 2397 3768
rect 2391 3766 2397 3767
rect 2444 3762 2446 3768
rect 2450 3767 2451 3771
rect 2455 3770 2456 3771
rect 2543 3771 2549 3772
rect 2543 3770 2544 3771
rect 2455 3768 2544 3770
rect 2455 3767 2456 3768
rect 2450 3766 2456 3767
rect 2543 3767 2544 3768
rect 2548 3767 2549 3771
rect 2543 3766 2549 3767
rect 2554 3771 2560 3772
rect 2554 3767 2555 3771
rect 2559 3770 2560 3771
rect 2703 3771 2709 3772
rect 2703 3770 2704 3771
rect 2559 3768 2704 3770
rect 2559 3767 2560 3768
rect 2554 3766 2560 3767
rect 2703 3767 2704 3768
rect 2708 3767 2709 3771
rect 2703 3766 2709 3767
rect 2871 3771 2877 3772
rect 2871 3767 2872 3771
rect 2876 3770 2877 3771
rect 2890 3771 2896 3772
rect 2890 3770 2891 3771
rect 2876 3768 2891 3770
rect 2876 3767 2877 3768
rect 2871 3766 2877 3767
rect 2890 3767 2891 3768
rect 2895 3767 2896 3771
rect 2890 3766 2896 3767
rect 3002 3771 3008 3772
rect 3002 3767 3003 3771
rect 3007 3770 3008 3771
rect 3047 3771 3053 3772
rect 3047 3770 3048 3771
rect 3007 3768 3048 3770
rect 3007 3767 3008 3768
rect 3002 3766 3008 3767
rect 3047 3767 3048 3768
rect 3052 3767 3053 3771
rect 3047 3766 3053 3767
rect 3223 3771 3229 3772
rect 3223 3767 3224 3771
rect 3228 3770 3229 3771
rect 3274 3771 3280 3772
rect 3274 3770 3275 3771
rect 3228 3768 3275 3770
rect 3228 3767 3229 3768
rect 3223 3766 3229 3767
rect 3274 3767 3275 3768
rect 3279 3767 3280 3771
rect 3274 3766 3280 3767
rect 3298 3771 3304 3772
rect 3298 3767 3299 3771
rect 3303 3770 3304 3771
rect 3399 3771 3405 3772
rect 3399 3770 3400 3771
rect 3303 3768 3400 3770
rect 3303 3767 3304 3768
rect 3298 3766 3304 3767
rect 3399 3767 3400 3768
rect 3404 3767 3405 3771
rect 3399 3766 3405 3767
rect 3410 3771 3416 3772
rect 3410 3767 3411 3771
rect 3415 3770 3416 3771
rect 3575 3771 3581 3772
rect 3575 3770 3576 3771
rect 3415 3768 3576 3770
rect 3415 3767 3416 3768
rect 3410 3766 3416 3767
rect 3575 3767 3576 3768
rect 3580 3767 3581 3771
rect 3575 3766 3581 3767
rect 3746 3771 3757 3772
rect 3746 3767 3747 3771
rect 3751 3767 3752 3771
rect 3756 3767 3757 3771
rect 3746 3766 3757 3767
rect 3903 3771 3912 3772
rect 3903 3767 3904 3771
rect 3911 3767 3912 3771
rect 3903 3766 3912 3767
rect 2598 3763 2604 3764
rect 2598 3762 2599 3763
rect 2444 3760 2599 3762
rect 222 3759 229 3760
rect 222 3755 223 3759
rect 228 3755 229 3759
rect 222 3754 229 3755
rect 258 3759 264 3760
rect 258 3755 259 3759
rect 263 3758 264 3759
rect 415 3759 421 3760
rect 415 3758 416 3759
rect 263 3756 416 3758
rect 263 3755 264 3756
rect 258 3754 264 3755
rect 415 3755 416 3756
rect 420 3755 421 3759
rect 415 3754 421 3755
rect 426 3759 432 3760
rect 426 3755 427 3759
rect 431 3758 432 3759
rect 615 3759 621 3760
rect 615 3758 616 3759
rect 431 3756 616 3758
rect 431 3755 432 3756
rect 426 3754 432 3755
rect 615 3755 616 3756
rect 620 3755 621 3759
rect 615 3754 621 3755
rect 815 3759 824 3760
rect 815 3755 816 3759
rect 823 3755 824 3759
rect 815 3754 824 3755
rect 906 3759 912 3760
rect 906 3755 907 3759
rect 911 3758 912 3759
rect 1023 3759 1029 3760
rect 1023 3758 1024 3759
rect 911 3756 1024 3758
rect 911 3755 912 3756
rect 906 3754 912 3755
rect 1023 3755 1024 3756
rect 1028 3755 1029 3759
rect 1023 3754 1029 3755
rect 1078 3759 1084 3760
rect 1078 3755 1079 3759
rect 1083 3758 1084 3759
rect 1231 3759 1237 3760
rect 1231 3758 1232 3759
rect 1083 3756 1232 3758
rect 1083 3755 1084 3756
rect 1078 3754 1084 3755
rect 1231 3755 1232 3756
rect 1236 3755 1237 3759
rect 1231 3754 1237 3755
rect 1242 3759 1248 3760
rect 1242 3755 1243 3759
rect 1247 3758 1248 3759
rect 1447 3759 1453 3760
rect 1447 3758 1448 3759
rect 1247 3756 1448 3758
rect 1247 3755 1248 3756
rect 1242 3754 1248 3755
rect 1447 3755 1448 3756
rect 1452 3755 1453 3759
rect 1447 3754 1453 3755
rect 1554 3759 1560 3760
rect 1554 3755 1555 3759
rect 1559 3758 1560 3759
rect 1671 3759 1677 3760
rect 1671 3758 1672 3759
rect 1559 3756 1672 3758
rect 1559 3755 1560 3756
rect 1554 3754 1560 3755
rect 1671 3755 1672 3756
rect 1676 3755 1677 3759
rect 2598 3759 2599 3760
rect 2603 3759 2604 3763
rect 2598 3758 2604 3759
rect 1671 3754 1677 3755
rect 2046 3752 2052 3753
rect 3942 3752 3948 3753
rect 2046 3748 2047 3752
rect 2051 3748 2052 3752
rect 2046 3747 2052 3748
rect 2070 3751 2076 3752
rect 2070 3747 2071 3751
rect 2075 3747 2076 3751
rect 2070 3746 2076 3747
rect 2182 3751 2188 3752
rect 2182 3747 2183 3751
rect 2187 3747 2188 3751
rect 2182 3746 2188 3747
rect 2326 3751 2332 3752
rect 2326 3747 2327 3751
rect 2331 3747 2332 3751
rect 2326 3746 2332 3747
rect 2478 3751 2484 3752
rect 2478 3747 2479 3751
rect 2483 3747 2484 3751
rect 2478 3746 2484 3747
rect 2638 3751 2644 3752
rect 2638 3747 2639 3751
rect 2643 3747 2644 3751
rect 2638 3746 2644 3747
rect 2806 3751 2812 3752
rect 2806 3747 2807 3751
rect 2811 3747 2812 3751
rect 2806 3746 2812 3747
rect 2982 3751 2988 3752
rect 2982 3747 2983 3751
rect 2987 3747 2988 3751
rect 2982 3746 2988 3747
rect 3158 3751 3164 3752
rect 3158 3747 3159 3751
rect 3163 3747 3164 3751
rect 3158 3746 3164 3747
rect 3334 3751 3340 3752
rect 3334 3747 3335 3751
rect 3339 3747 3340 3751
rect 3334 3746 3340 3747
rect 3510 3751 3516 3752
rect 3510 3747 3511 3751
rect 3515 3747 3516 3751
rect 3510 3746 3516 3747
rect 3686 3751 3692 3752
rect 3686 3747 3687 3751
rect 3691 3747 3692 3751
rect 3686 3746 3692 3747
rect 3838 3751 3844 3752
rect 3838 3747 3839 3751
rect 3843 3747 3844 3751
rect 3942 3748 3943 3752
rect 3947 3748 3948 3752
rect 3942 3747 3948 3748
rect 3838 3746 3844 3747
rect 2154 3743 2160 3744
rect 110 3740 116 3741
rect 2006 3740 2012 3741
rect 110 3736 111 3740
rect 115 3736 116 3740
rect 110 3735 116 3736
rect 158 3739 164 3740
rect 158 3735 159 3739
rect 163 3735 164 3739
rect 158 3734 164 3735
rect 350 3739 356 3740
rect 350 3735 351 3739
rect 355 3735 356 3739
rect 350 3734 356 3735
rect 550 3739 556 3740
rect 550 3735 551 3739
rect 555 3735 556 3739
rect 550 3734 556 3735
rect 750 3739 756 3740
rect 750 3735 751 3739
rect 755 3735 756 3739
rect 750 3734 756 3735
rect 958 3739 964 3740
rect 958 3735 959 3739
rect 963 3735 964 3739
rect 958 3734 964 3735
rect 1166 3739 1172 3740
rect 1166 3735 1167 3739
rect 1171 3735 1172 3739
rect 1166 3734 1172 3735
rect 1382 3739 1388 3740
rect 1382 3735 1383 3739
rect 1387 3735 1388 3739
rect 1382 3734 1388 3735
rect 1606 3739 1612 3740
rect 1606 3735 1607 3739
rect 1611 3735 1612 3739
rect 2006 3736 2007 3740
rect 2011 3736 2012 3740
rect 2154 3739 2155 3743
rect 2159 3742 2160 3743
rect 2271 3743 2277 3744
rect 2159 3740 2225 3742
rect 2159 3739 2160 3740
rect 2154 3738 2160 3739
rect 2271 3739 2272 3743
rect 2276 3742 2277 3743
rect 2554 3743 2560 3744
rect 2276 3740 2369 3742
rect 2276 3739 2277 3740
rect 2271 3738 2277 3739
rect 2554 3739 2555 3743
rect 2559 3739 2560 3743
rect 2554 3738 2560 3739
rect 2598 3743 2604 3744
rect 2598 3739 2599 3743
rect 2603 3742 2604 3743
rect 2882 3743 2888 3744
rect 2603 3740 2681 3742
rect 2603 3739 2604 3740
rect 2598 3738 2604 3739
rect 2882 3739 2883 3743
rect 2887 3739 2888 3743
rect 2882 3738 2888 3739
rect 2890 3743 2896 3744
rect 2890 3739 2891 3743
rect 2895 3742 2896 3743
rect 3298 3743 3304 3744
rect 3298 3742 3299 3743
rect 2895 3740 3025 3742
rect 3237 3740 3299 3742
rect 2895 3739 2896 3740
rect 2890 3738 2896 3739
rect 3298 3739 3299 3740
rect 3303 3739 3304 3743
rect 3298 3738 3304 3739
rect 3410 3743 3416 3744
rect 3410 3739 3411 3743
rect 3415 3739 3416 3743
rect 3671 3743 3677 3744
rect 3410 3738 3416 3739
rect 3586 3739 3592 3740
rect 2140 3736 2149 3738
rect 2006 3735 2012 3736
rect 2046 3735 2052 3736
rect 1606 3734 1612 3735
rect 258 3731 264 3732
rect 258 3730 259 3731
rect 237 3728 259 3730
rect 258 3727 259 3728
rect 263 3727 264 3731
rect 258 3726 264 3727
rect 426 3731 432 3732
rect 426 3727 427 3731
rect 431 3727 432 3731
rect 426 3726 432 3727
rect 447 3731 453 3732
rect 447 3727 448 3731
rect 452 3730 453 3731
rect 906 3731 912 3732
rect 906 3730 907 3731
rect 452 3728 593 3730
rect 829 3728 907 3730
rect 452 3727 453 3728
rect 447 3726 453 3727
rect 906 3727 907 3728
rect 911 3727 912 3731
rect 1078 3731 1084 3732
rect 1078 3730 1079 3731
rect 1037 3728 1079 3730
rect 906 3726 912 3727
rect 1078 3727 1079 3728
rect 1083 3727 1084 3731
rect 1078 3726 1084 3727
rect 1242 3731 1248 3732
rect 1242 3727 1243 3731
rect 1247 3727 1248 3731
rect 1242 3726 1248 3727
rect 1346 3731 1352 3732
rect 1346 3727 1347 3731
rect 1351 3730 1352 3731
rect 1599 3731 1605 3732
rect 1351 3728 1425 3730
rect 1351 3727 1352 3728
rect 1346 3726 1352 3727
rect 1599 3727 1600 3731
rect 1604 3730 1605 3731
rect 2046 3731 2047 3735
rect 2051 3731 2052 3735
rect 2138 3735 2144 3736
rect 2046 3730 2052 3731
rect 2070 3732 2076 3733
rect 1604 3728 1649 3730
rect 2070 3728 2071 3732
rect 2075 3728 2076 3732
rect 2138 3731 2139 3735
rect 2143 3731 2144 3735
rect 3586 3735 3587 3739
rect 3591 3735 3592 3739
rect 3671 3739 3672 3743
rect 3676 3742 3677 3743
rect 3676 3740 3729 3742
rect 3676 3739 3677 3740
rect 3671 3738 3677 3739
rect 3908 3736 3917 3738
rect 3586 3734 3592 3735
rect 3906 3735 3912 3736
rect 2138 3730 2144 3731
rect 2182 3732 2188 3733
rect 1604 3727 1605 3728
rect 2070 3727 2076 3728
rect 2182 3728 2183 3732
rect 2187 3728 2188 3732
rect 2182 3727 2188 3728
rect 2326 3732 2332 3733
rect 2326 3728 2327 3732
rect 2331 3728 2332 3732
rect 2326 3727 2332 3728
rect 2478 3732 2484 3733
rect 2478 3728 2479 3732
rect 2483 3728 2484 3732
rect 2478 3727 2484 3728
rect 2638 3732 2644 3733
rect 2638 3728 2639 3732
rect 2643 3728 2644 3732
rect 2638 3727 2644 3728
rect 2806 3732 2812 3733
rect 2806 3728 2807 3732
rect 2811 3728 2812 3732
rect 2806 3727 2812 3728
rect 2982 3732 2988 3733
rect 2982 3728 2983 3732
rect 2987 3728 2988 3732
rect 2982 3727 2988 3728
rect 3158 3732 3164 3733
rect 3158 3728 3159 3732
rect 3163 3728 3164 3732
rect 3158 3727 3164 3728
rect 3334 3732 3340 3733
rect 3334 3728 3335 3732
rect 3339 3728 3340 3732
rect 3334 3727 3340 3728
rect 3510 3732 3516 3733
rect 3510 3728 3511 3732
rect 3515 3728 3516 3732
rect 3510 3727 3516 3728
rect 3686 3732 3692 3733
rect 3686 3728 3687 3732
rect 3691 3728 3692 3732
rect 3686 3727 3692 3728
rect 3838 3732 3844 3733
rect 3838 3728 3839 3732
rect 3843 3728 3844 3732
rect 3906 3731 3907 3735
rect 3911 3731 3912 3735
rect 3906 3730 3912 3731
rect 3942 3735 3948 3736
rect 3942 3731 3943 3735
rect 3947 3731 3948 3735
rect 3942 3730 3948 3731
rect 3838 3727 3844 3728
rect 1599 3726 1605 3727
rect 110 3723 116 3724
rect 110 3719 111 3723
rect 115 3719 116 3723
rect 2006 3723 2012 3724
rect 110 3718 116 3719
rect 158 3720 164 3721
rect 158 3716 159 3720
rect 163 3716 164 3720
rect 158 3715 164 3716
rect 350 3720 356 3721
rect 350 3716 351 3720
rect 355 3716 356 3720
rect 350 3715 356 3716
rect 550 3720 556 3721
rect 550 3716 551 3720
rect 555 3716 556 3720
rect 550 3715 556 3716
rect 750 3720 756 3721
rect 750 3716 751 3720
rect 755 3716 756 3720
rect 750 3715 756 3716
rect 958 3720 964 3721
rect 958 3716 959 3720
rect 963 3716 964 3720
rect 958 3715 964 3716
rect 1166 3720 1172 3721
rect 1166 3716 1167 3720
rect 1171 3716 1172 3720
rect 1166 3715 1172 3716
rect 1382 3720 1388 3721
rect 1382 3716 1383 3720
rect 1387 3716 1388 3720
rect 1382 3715 1388 3716
rect 1606 3720 1612 3721
rect 1606 3716 1607 3720
rect 1611 3716 1612 3720
rect 2006 3719 2007 3723
rect 2011 3719 2012 3723
rect 2006 3718 2012 3719
rect 1606 3715 1612 3716
rect 2070 3660 2076 3661
rect 2046 3657 2052 3658
rect 2046 3653 2047 3657
rect 2051 3653 2052 3657
rect 2070 3656 2071 3660
rect 2075 3656 2076 3660
rect 2070 3655 2076 3656
rect 2198 3660 2204 3661
rect 2198 3656 2199 3660
rect 2203 3656 2204 3660
rect 2198 3655 2204 3656
rect 2366 3660 2372 3661
rect 2366 3656 2367 3660
rect 2371 3656 2372 3660
rect 2366 3655 2372 3656
rect 2550 3660 2556 3661
rect 2550 3656 2551 3660
rect 2555 3656 2556 3660
rect 2550 3655 2556 3656
rect 2734 3660 2740 3661
rect 2734 3656 2735 3660
rect 2739 3656 2740 3660
rect 2734 3655 2740 3656
rect 2926 3660 2932 3661
rect 2926 3656 2927 3660
rect 2931 3656 2932 3660
rect 2926 3655 2932 3656
rect 3110 3660 3116 3661
rect 3110 3656 3111 3660
rect 3115 3656 3116 3660
rect 3110 3655 3116 3656
rect 3294 3660 3300 3661
rect 3294 3656 3295 3660
rect 3299 3656 3300 3660
rect 3294 3655 3300 3656
rect 3478 3660 3484 3661
rect 3478 3656 3479 3660
rect 3483 3656 3484 3660
rect 3478 3655 3484 3656
rect 3670 3660 3676 3661
rect 3670 3656 3671 3660
rect 3675 3656 3676 3660
rect 3670 3655 3676 3656
rect 3838 3660 3844 3661
rect 3838 3656 3839 3660
rect 3843 3656 3844 3660
rect 3838 3655 3844 3656
rect 3942 3657 3948 3658
rect 150 3652 156 3653
rect 110 3649 116 3650
rect 110 3645 111 3649
rect 115 3645 116 3649
rect 150 3648 151 3652
rect 155 3648 156 3652
rect 150 3647 156 3648
rect 382 3652 388 3653
rect 382 3648 383 3652
rect 387 3648 388 3652
rect 382 3647 388 3648
rect 614 3652 620 3653
rect 614 3648 615 3652
rect 619 3648 620 3652
rect 614 3647 620 3648
rect 838 3652 844 3653
rect 838 3648 839 3652
rect 843 3648 844 3652
rect 838 3647 844 3648
rect 1054 3652 1060 3653
rect 1054 3648 1055 3652
rect 1059 3648 1060 3652
rect 1054 3647 1060 3648
rect 1262 3652 1268 3653
rect 1262 3648 1263 3652
rect 1267 3648 1268 3652
rect 1262 3647 1268 3648
rect 1478 3652 1484 3653
rect 1478 3648 1479 3652
rect 1483 3648 1484 3652
rect 1478 3647 1484 3648
rect 1694 3652 1700 3653
rect 2046 3652 2052 3653
rect 3942 3653 3943 3657
rect 3947 3653 3948 3657
rect 3942 3652 3948 3653
rect 1694 3648 1695 3652
rect 1699 3648 1700 3652
rect 2146 3651 2152 3652
rect 1694 3647 1700 3648
rect 2006 3649 2012 3650
rect 110 3644 116 3645
rect 2006 3645 2007 3649
rect 2011 3645 2012 3649
rect 2146 3647 2147 3651
rect 2151 3647 2152 3651
rect 2146 3646 2152 3647
rect 2274 3651 2280 3652
rect 2274 3647 2275 3651
rect 2279 3647 2280 3651
rect 2274 3646 2280 3647
rect 2442 3651 2448 3652
rect 2442 3647 2443 3651
rect 2447 3647 2448 3651
rect 2442 3646 2448 3647
rect 2626 3651 2632 3652
rect 2626 3647 2627 3651
rect 2631 3647 2632 3651
rect 3002 3651 3008 3652
rect 2626 3646 2632 3647
rect 2636 3648 2777 3650
rect 2006 3644 2012 3645
rect 222 3643 228 3644
rect 222 3639 223 3643
rect 227 3639 228 3643
rect 222 3638 228 3639
rect 234 3643 240 3644
rect 234 3639 235 3643
rect 239 3642 240 3643
rect 466 3643 472 3644
rect 239 3640 425 3642
rect 239 3639 240 3640
rect 234 3638 240 3639
rect 466 3639 467 3643
rect 471 3642 472 3643
rect 1038 3643 1044 3644
rect 1038 3642 1039 3643
rect 471 3640 657 3642
rect 917 3640 1039 3642
rect 471 3639 472 3640
rect 466 3638 472 3639
rect 1038 3639 1039 3640
rect 1043 3639 1044 3643
rect 1038 3638 1044 3639
rect 1130 3643 1136 3644
rect 1130 3639 1131 3643
rect 1135 3639 1136 3643
rect 1130 3638 1136 3639
rect 1338 3643 1344 3644
rect 1338 3639 1339 3643
rect 1343 3639 1344 3643
rect 1338 3638 1344 3639
rect 1554 3643 1560 3644
rect 1554 3639 1555 3643
rect 1559 3639 1560 3643
rect 1554 3638 1560 3639
rect 1562 3643 1568 3644
rect 1562 3639 1563 3643
rect 1567 3642 1568 3643
rect 1567 3640 1737 3642
rect 2070 3641 2076 3642
rect 2046 3640 2052 3641
rect 1567 3639 1568 3640
rect 1562 3638 1568 3639
rect 2046 3636 2047 3640
rect 2051 3636 2052 3640
rect 2070 3637 2071 3641
rect 2075 3637 2076 3641
rect 2070 3636 2076 3637
rect 2198 3641 2204 3642
rect 2198 3637 2199 3641
rect 2203 3637 2204 3641
rect 2198 3636 2204 3637
rect 2366 3641 2372 3642
rect 2366 3637 2367 3641
rect 2371 3637 2372 3641
rect 2366 3636 2372 3637
rect 2550 3641 2556 3642
rect 2550 3637 2551 3641
rect 2555 3637 2556 3641
rect 2550 3636 2556 3637
rect 2046 3635 2052 3636
rect 2170 3635 2176 3636
rect 150 3633 156 3634
rect 110 3632 116 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 150 3629 151 3633
rect 155 3629 156 3633
rect 150 3628 156 3629
rect 382 3633 388 3634
rect 382 3629 383 3633
rect 387 3629 388 3633
rect 382 3628 388 3629
rect 614 3633 620 3634
rect 614 3629 615 3633
rect 619 3629 620 3633
rect 614 3628 620 3629
rect 838 3633 844 3634
rect 838 3629 839 3633
rect 843 3629 844 3633
rect 838 3628 844 3629
rect 1054 3633 1060 3634
rect 1054 3629 1055 3633
rect 1059 3629 1060 3633
rect 1054 3628 1060 3629
rect 1262 3633 1268 3634
rect 1262 3629 1263 3633
rect 1267 3629 1268 3633
rect 1262 3628 1268 3629
rect 1478 3633 1484 3634
rect 1478 3629 1479 3633
rect 1483 3629 1484 3633
rect 1478 3628 1484 3629
rect 1694 3633 1700 3634
rect 1694 3629 1695 3633
rect 1699 3629 1700 3633
rect 1694 3628 1700 3629
rect 2006 3632 2012 3633
rect 2006 3628 2007 3632
rect 2011 3628 2012 3632
rect 2170 3631 2171 3635
rect 2175 3634 2176 3635
rect 2636 3634 2638 3648
rect 3002 3647 3003 3651
rect 3007 3647 3008 3651
rect 3002 3646 3008 3647
rect 3186 3651 3192 3652
rect 3186 3647 3187 3651
rect 3191 3647 3192 3651
rect 3186 3646 3192 3647
rect 3194 3651 3200 3652
rect 3194 3647 3195 3651
rect 3199 3650 3200 3651
rect 3378 3651 3384 3652
rect 3199 3648 3337 3650
rect 3199 3647 3200 3648
rect 3194 3646 3200 3647
rect 3378 3647 3379 3651
rect 3383 3650 3384 3651
rect 3746 3651 3752 3652
rect 3383 3648 3521 3650
rect 3383 3647 3384 3648
rect 3378 3646 3384 3647
rect 3746 3647 3747 3651
rect 3751 3647 3752 3651
rect 3746 3646 3752 3647
rect 3914 3651 3920 3652
rect 3914 3647 3915 3651
rect 3919 3647 3920 3651
rect 3914 3646 3920 3647
rect 2734 3641 2740 3642
rect 2734 3637 2735 3641
rect 2739 3637 2740 3641
rect 2734 3636 2740 3637
rect 2926 3641 2932 3642
rect 2926 3637 2927 3641
rect 2931 3637 2932 3641
rect 2926 3636 2932 3637
rect 3110 3641 3116 3642
rect 3110 3637 3111 3641
rect 3115 3637 3116 3641
rect 3110 3636 3116 3637
rect 3294 3641 3300 3642
rect 3294 3637 3295 3641
rect 3299 3637 3300 3641
rect 3294 3636 3300 3637
rect 3478 3641 3484 3642
rect 3478 3637 3479 3641
rect 3483 3637 3484 3641
rect 3478 3636 3484 3637
rect 3670 3641 3676 3642
rect 3670 3637 3671 3641
rect 3675 3637 3676 3641
rect 3670 3636 3676 3637
rect 3838 3641 3844 3642
rect 3838 3637 3839 3641
rect 3843 3637 3844 3641
rect 3838 3636 3844 3637
rect 3942 3640 3948 3641
rect 3942 3636 3943 3640
rect 3947 3636 3948 3640
rect 3942 3635 3948 3636
rect 2175 3632 2638 3634
rect 2175 3631 2176 3632
rect 2170 3630 2176 3631
rect 110 3627 116 3628
rect 2006 3627 2012 3628
rect 1346 3619 1352 3620
rect 1346 3618 1347 3619
rect 1032 3616 1347 3618
rect 215 3611 221 3612
rect 215 3607 216 3611
rect 220 3610 221 3611
rect 234 3611 240 3612
rect 234 3610 235 3611
rect 220 3608 235 3610
rect 220 3607 221 3608
rect 215 3606 221 3607
rect 234 3607 235 3608
rect 239 3607 240 3611
rect 234 3606 240 3607
rect 447 3611 453 3612
rect 447 3607 448 3611
rect 452 3610 453 3611
rect 466 3611 472 3612
rect 466 3610 467 3611
rect 452 3608 467 3610
rect 452 3607 453 3608
rect 447 3606 453 3607
rect 466 3607 467 3608
rect 471 3607 472 3611
rect 466 3606 472 3607
rect 679 3611 688 3612
rect 679 3607 680 3611
rect 687 3607 688 3611
rect 679 3606 688 3607
rect 903 3611 909 3612
rect 903 3607 904 3611
rect 908 3610 909 3611
rect 1032 3610 1034 3616
rect 1346 3615 1347 3616
rect 1351 3615 1352 3619
rect 1346 3614 1352 3615
rect 2135 3619 2144 3620
rect 2135 3615 2136 3619
rect 2143 3615 2144 3619
rect 2135 3614 2144 3615
rect 2146 3619 2152 3620
rect 2146 3615 2147 3619
rect 2151 3618 2152 3619
rect 2263 3619 2269 3620
rect 2263 3618 2264 3619
rect 2151 3616 2264 3618
rect 2151 3615 2152 3616
rect 2146 3614 2152 3615
rect 2263 3615 2264 3616
rect 2268 3615 2269 3619
rect 2263 3614 2269 3615
rect 2274 3619 2280 3620
rect 2274 3615 2275 3619
rect 2279 3618 2280 3619
rect 2431 3619 2437 3620
rect 2431 3618 2432 3619
rect 2279 3616 2432 3618
rect 2279 3615 2280 3616
rect 2274 3614 2280 3615
rect 2431 3615 2432 3616
rect 2436 3615 2437 3619
rect 2431 3614 2437 3615
rect 2442 3619 2448 3620
rect 2442 3615 2443 3619
rect 2447 3618 2448 3619
rect 2615 3619 2621 3620
rect 2615 3618 2616 3619
rect 2447 3616 2616 3618
rect 2447 3615 2448 3616
rect 2442 3614 2448 3615
rect 2615 3615 2616 3616
rect 2620 3615 2621 3619
rect 2615 3614 2621 3615
rect 2626 3619 2632 3620
rect 2626 3615 2627 3619
rect 2631 3618 2632 3619
rect 2799 3619 2805 3620
rect 2799 3618 2800 3619
rect 2631 3616 2800 3618
rect 2631 3615 2632 3616
rect 2626 3614 2632 3615
rect 2799 3615 2800 3616
rect 2804 3615 2805 3619
rect 2799 3614 2805 3615
rect 2991 3619 2997 3620
rect 2991 3615 2992 3619
rect 2996 3618 2997 3619
rect 2999 3619 3005 3620
rect 2999 3618 3000 3619
rect 2996 3616 3000 3618
rect 2996 3615 2997 3616
rect 2991 3614 2997 3615
rect 2999 3615 3000 3616
rect 3004 3615 3005 3619
rect 2999 3614 3005 3615
rect 3175 3619 3181 3620
rect 3175 3615 3176 3619
rect 3180 3618 3181 3619
rect 3194 3619 3200 3620
rect 3194 3618 3195 3619
rect 3180 3616 3195 3618
rect 3180 3615 3181 3616
rect 3175 3614 3181 3615
rect 3194 3615 3195 3616
rect 3199 3615 3200 3619
rect 3194 3614 3200 3615
rect 3359 3619 3365 3620
rect 3359 3615 3360 3619
rect 3364 3618 3365 3619
rect 3378 3619 3384 3620
rect 3378 3618 3379 3619
rect 3364 3616 3379 3618
rect 3364 3615 3365 3616
rect 3359 3614 3365 3615
rect 3378 3615 3379 3616
rect 3383 3615 3384 3619
rect 3378 3614 3384 3615
rect 3543 3619 3549 3620
rect 3543 3615 3544 3619
rect 3548 3618 3549 3619
rect 3586 3619 3592 3620
rect 3586 3618 3587 3619
rect 3548 3616 3587 3618
rect 3548 3615 3549 3616
rect 3543 3614 3549 3615
rect 3586 3615 3587 3616
rect 3591 3615 3592 3619
rect 3586 3614 3592 3615
rect 3714 3619 3720 3620
rect 3714 3615 3715 3619
rect 3719 3618 3720 3619
rect 3735 3619 3741 3620
rect 3735 3618 3736 3619
rect 3719 3616 3736 3618
rect 3719 3615 3720 3616
rect 3714 3614 3720 3615
rect 3735 3615 3736 3616
rect 3740 3615 3741 3619
rect 3735 3614 3741 3615
rect 3903 3619 3912 3620
rect 3903 3615 3904 3619
rect 3911 3615 3912 3619
rect 3903 3614 3912 3615
rect 908 3608 1034 3610
rect 1038 3611 1044 3612
rect 908 3607 909 3608
rect 903 3606 909 3607
rect 1038 3607 1039 3611
rect 1043 3610 1044 3611
rect 1119 3611 1125 3612
rect 1119 3610 1120 3611
rect 1043 3608 1120 3610
rect 1043 3607 1044 3608
rect 1038 3606 1044 3607
rect 1119 3607 1120 3608
rect 1124 3607 1125 3611
rect 1119 3606 1125 3607
rect 1130 3611 1136 3612
rect 1130 3607 1131 3611
rect 1135 3610 1136 3611
rect 1327 3611 1333 3612
rect 1327 3610 1328 3611
rect 1135 3608 1328 3610
rect 1135 3607 1136 3608
rect 1130 3606 1136 3607
rect 1327 3607 1328 3608
rect 1332 3607 1333 3611
rect 1327 3606 1333 3607
rect 1543 3611 1549 3612
rect 1543 3607 1544 3611
rect 1548 3610 1549 3611
rect 1562 3611 1568 3612
rect 1562 3610 1563 3611
rect 1548 3608 1563 3610
rect 1548 3607 1549 3608
rect 1543 3606 1549 3607
rect 1562 3607 1563 3608
rect 1567 3607 1568 3611
rect 1562 3606 1568 3607
rect 1759 3611 1768 3612
rect 1759 3607 1760 3611
rect 1767 3607 1768 3611
rect 1759 3606 1768 3607
rect 2167 3603 2176 3604
rect 2167 3599 2168 3603
rect 2175 3599 2176 3603
rect 2167 3598 2176 3599
rect 2178 3603 2184 3604
rect 2178 3599 2179 3603
rect 2183 3602 2184 3603
rect 2343 3603 2349 3604
rect 2343 3602 2344 3603
rect 2183 3600 2344 3602
rect 2183 3599 2184 3600
rect 2178 3598 2184 3599
rect 2343 3599 2344 3600
rect 2348 3599 2349 3603
rect 2343 3598 2349 3599
rect 2354 3603 2360 3604
rect 2354 3599 2355 3603
rect 2359 3602 2360 3603
rect 2535 3603 2541 3604
rect 2535 3602 2536 3603
rect 2359 3600 2536 3602
rect 2359 3599 2360 3600
rect 2354 3598 2360 3599
rect 2535 3599 2536 3600
rect 2540 3599 2541 3603
rect 2535 3598 2541 3599
rect 2582 3603 2588 3604
rect 2582 3599 2583 3603
rect 2587 3602 2588 3603
rect 2735 3603 2741 3604
rect 2735 3602 2736 3603
rect 2587 3600 2736 3602
rect 2587 3599 2588 3600
rect 2582 3598 2588 3599
rect 2735 3599 2736 3600
rect 2740 3599 2741 3603
rect 2735 3598 2741 3599
rect 2935 3603 2941 3604
rect 2935 3599 2936 3603
rect 2940 3602 2941 3603
rect 2978 3603 2984 3604
rect 2978 3602 2979 3603
rect 2940 3600 2979 3602
rect 2940 3599 2941 3600
rect 2935 3598 2941 3599
rect 2978 3599 2979 3600
rect 2983 3599 2984 3603
rect 2978 3598 2984 3599
rect 2991 3603 2997 3604
rect 2991 3599 2992 3603
rect 2996 3602 2997 3603
rect 3127 3603 3133 3604
rect 3127 3602 3128 3603
rect 2996 3600 3128 3602
rect 2996 3599 2997 3600
rect 2991 3598 2997 3599
rect 3127 3599 3128 3600
rect 3132 3599 3133 3603
rect 3127 3598 3133 3599
rect 3186 3603 3192 3604
rect 3186 3599 3187 3603
rect 3191 3602 3192 3603
rect 3319 3603 3325 3604
rect 3319 3602 3320 3603
rect 3191 3600 3320 3602
rect 3191 3599 3192 3600
rect 3186 3598 3192 3599
rect 3319 3599 3320 3600
rect 3324 3599 3325 3603
rect 3319 3598 3325 3599
rect 3330 3603 3336 3604
rect 3330 3599 3331 3603
rect 3335 3602 3336 3603
rect 3511 3603 3517 3604
rect 3511 3602 3512 3603
rect 3335 3600 3512 3602
rect 3335 3599 3336 3600
rect 3330 3598 3336 3599
rect 3511 3599 3512 3600
rect 3516 3599 3517 3603
rect 3511 3598 3517 3599
rect 3522 3603 3528 3604
rect 3522 3599 3523 3603
rect 3527 3602 3528 3603
rect 3703 3603 3709 3604
rect 3703 3602 3704 3603
rect 3527 3600 3704 3602
rect 3527 3599 3528 3600
rect 3522 3598 3528 3599
rect 3703 3599 3704 3600
rect 3708 3599 3709 3603
rect 3703 3598 3709 3599
rect 3903 3603 3909 3604
rect 3903 3599 3904 3603
rect 3908 3602 3909 3603
rect 3914 3603 3920 3604
rect 3914 3602 3915 3603
rect 3908 3600 3915 3602
rect 3908 3599 3909 3600
rect 3903 3598 3909 3599
rect 3914 3599 3915 3600
rect 3919 3599 3920 3603
rect 3914 3598 3920 3599
rect 231 3595 237 3596
rect 231 3591 232 3595
rect 236 3594 237 3595
rect 242 3595 248 3596
rect 236 3591 238 3594
rect 231 3590 238 3591
rect 242 3591 243 3595
rect 247 3594 248 3595
rect 423 3595 429 3596
rect 423 3594 424 3595
rect 247 3592 424 3594
rect 247 3591 248 3592
rect 242 3590 248 3591
rect 423 3591 424 3592
rect 428 3591 429 3595
rect 423 3590 429 3591
rect 434 3595 440 3596
rect 434 3591 435 3595
rect 439 3594 440 3595
rect 623 3595 629 3596
rect 623 3594 624 3595
rect 439 3592 624 3594
rect 439 3591 440 3592
rect 434 3590 440 3591
rect 623 3591 624 3592
rect 628 3591 629 3595
rect 623 3590 629 3591
rect 634 3595 640 3596
rect 634 3591 635 3595
rect 639 3594 640 3595
rect 839 3595 845 3596
rect 839 3594 840 3595
rect 639 3592 840 3594
rect 639 3591 640 3592
rect 634 3590 640 3591
rect 839 3591 840 3592
rect 844 3591 845 3595
rect 839 3590 845 3591
rect 1055 3595 1061 3596
rect 1055 3591 1056 3595
rect 1060 3594 1061 3595
rect 1127 3595 1133 3596
rect 1127 3594 1128 3595
rect 1060 3592 1128 3594
rect 1060 3591 1061 3592
rect 1055 3590 1061 3591
rect 1127 3591 1128 3592
rect 1132 3591 1133 3595
rect 1127 3590 1133 3591
rect 1279 3595 1285 3596
rect 1279 3591 1280 3595
rect 1284 3594 1285 3595
rect 1298 3595 1304 3596
rect 1298 3594 1299 3595
rect 1284 3592 1299 3594
rect 1284 3591 1285 3592
rect 1279 3590 1285 3591
rect 1298 3591 1299 3592
rect 1303 3591 1304 3595
rect 1298 3590 1304 3591
rect 1338 3595 1344 3596
rect 1338 3591 1339 3595
rect 1343 3594 1344 3595
rect 1511 3595 1517 3596
rect 1511 3594 1512 3595
rect 1343 3592 1512 3594
rect 1343 3591 1344 3592
rect 1338 3590 1344 3591
rect 1511 3591 1512 3592
rect 1516 3591 1517 3595
rect 1511 3590 1517 3591
rect 1751 3595 1760 3596
rect 1751 3591 1752 3595
rect 1759 3591 1760 3595
rect 1751 3590 1760 3591
rect 236 3586 238 3590
rect 271 3587 277 3588
rect 271 3586 272 3587
rect 236 3584 272 3586
rect 271 3583 272 3584
rect 276 3583 277 3587
rect 271 3582 277 3583
rect 2046 3584 2052 3585
rect 3942 3584 3948 3585
rect 2046 3580 2047 3584
rect 2051 3580 2052 3584
rect 2046 3579 2052 3580
rect 2102 3583 2108 3584
rect 2102 3579 2103 3583
rect 2107 3579 2108 3583
rect 2102 3578 2108 3579
rect 2278 3583 2284 3584
rect 2278 3579 2279 3583
rect 2283 3579 2284 3583
rect 2278 3578 2284 3579
rect 2470 3583 2476 3584
rect 2470 3579 2471 3583
rect 2475 3579 2476 3583
rect 2470 3578 2476 3579
rect 2670 3583 2676 3584
rect 2670 3579 2671 3583
rect 2675 3579 2676 3583
rect 2670 3578 2676 3579
rect 2870 3583 2876 3584
rect 2870 3579 2871 3583
rect 2875 3579 2876 3583
rect 2870 3578 2876 3579
rect 3062 3583 3068 3584
rect 3062 3579 3063 3583
rect 3067 3579 3068 3583
rect 3062 3578 3068 3579
rect 3254 3583 3260 3584
rect 3254 3579 3255 3583
rect 3259 3579 3260 3583
rect 3254 3578 3260 3579
rect 3446 3583 3452 3584
rect 3446 3579 3447 3583
rect 3451 3579 3452 3583
rect 3446 3578 3452 3579
rect 3638 3583 3644 3584
rect 3638 3579 3639 3583
rect 3643 3579 3644 3583
rect 3638 3578 3644 3579
rect 3838 3583 3844 3584
rect 3838 3579 3839 3583
rect 3843 3579 3844 3583
rect 3942 3580 3943 3584
rect 3947 3580 3948 3584
rect 3942 3579 3948 3580
rect 3838 3578 3844 3579
rect 110 3576 116 3577
rect 2006 3576 2012 3577
rect 110 3572 111 3576
rect 115 3572 116 3576
rect 110 3571 116 3572
rect 166 3575 172 3576
rect 166 3571 167 3575
rect 171 3571 172 3575
rect 166 3570 172 3571
rect 358 3575 364 3576
rect 358 3571 359 3575
rect 363 3571 364 3575
rect 358 3570 364 3571
rect 558 3575 564 3576
rect 558 3571 559 3575
rect 563 3571 564 3575
rect 558 3570 564 3571
rect 774 3575 780 3576
rect 774 3571 775 3575
rect 779 3571 780 3575
rect 774 3570 780 3571
rect 990 3575 996 3576
rect 990 3571 991 3575
rect 995 3571 996 3575
rect 990 3570 996 3571
rect 1214 3575 1220 3576
rect 1214 3571 1215 3575
rect 1219 3571 1220 3575
rect 1214 3570 1220 3571
rect 1446 3575 1452 3576
rect 1446 3571 1447 3575
rect 1451 3571 1452 3575
rect 1446 3570 1452 3571
rect 1686 3575 1692 3576
rect 1686 3571 1687 3575
rect 1691 3571 1692 3575
rect 2006 3572 2007 3576
rect 2011 3572 2012 3576
rect 2006 3571 2012 3572
rect 2178 3575 2184 3576
rect 2178 3571 2179 3575
rect 2183 3571 2184 3575
rect 1686 3570 1692 3571
rect 2178 3570 2184 3571
rect 2354 3575 2360 3576
rect 2354 3571 2355 3575
rect 2359 3571 2360 3575
rect 2582 3575 2588 3576
rect 2582 3574 2583 3575
rect 2549 3572 2583 3574
rect 2354 3570 2360 3571
rect 2582 3571 2583 3572
rect 2587 3571 2588 3575
rect 2582 3570 2588 3571
rect 2598 3575 2604 3576
rect 2598 3571 2599 3575
rect 2603 3574 2604 3575
rect 2991 3575 2997 3576
rect 2991 3574 2992 3575
rect 2603 3572 2713 3574
rect 2949 3572 2992 3574
rect 2603 3571 2604 3572
rect 2598 3570 2604 3571
rect 2991 3571 2992 3572
rect 2996 3571 2997 3575
rect 2991 3570 2997 3571
rect 2999 3575 3005 3576
rect 2999 3571 3000 3575
rect 3004 3574 3005 3575
rect 3330 3575 3336 3576
rect 3004 3572 3105 3574
rect 3004 3571 3005 3572
rect 2999 3570 3005 3571
rect 3330 3571 3331 3575
rect 3335 3571 3336 3575
rect 3330 3570 3336 3571
rect 3522 3575 3528 3576
rect 3522 3571 3523 3575
rect 3527 3571 3528 3575
rect 3522 3570 3528 3571
rect 3714 3575 3720 3576
rect 3714 3571 3715 3575
rect 3719 3571 3720 3575
rect 3714 3570 3720 3571
rect 3914 3571 3920 3572
rect 242 3567 248 3568
rect 242 3563 243 3567
rect 247 3563 248 3567
rect 242 3562 248 3563
rect 434 3567 440 3568
rect 434 3563 435 3567
rect 439 3563 440 3567
rect 434 3562 440 3563
rect 634 3567 640 3568
rect 634 3563 635 3567
rect 639 3563 640 3567
rect 634 3562 640 3563
rect 682 3567 688 3568
rect 682 3563 683 3567
rect 687 3566 688 3567
rect 1127 3567 1133 3568
rect 687 3564 817 3566
rect 687 3563 688 3564
rect 682 3562 688 3563
rect 1066 3563 1072 3564
rect 110 3559 116 3560
rect 110 3555 111 3559
rect 115 3555 116 3559
rect 1066 3559 1067 3563
rect 1071 3559 1072 3563
rect 1127 3563 1128 3567
rect 1132 3566 1133 3567
rect 1298 3567 1304 3568
rect 1132 3564 1257 3566
rect 1132 3563 1133 3564
rect 1127 3562 1133 3563
rect 1298 3563 1299 3567
rect 1303 3566 1304 3567
rect 1762 3567 1768 3568
rect 1303 3564 1489 3566
rect 1303 3563 1304 3564
rect 1298 3562 1304 3563
rect 1762 3563 1763 3567
rect 1767 3563 1768 3567
rect 1762 3562 1768 3563
rect 2046 3567 2052 3568
rect 2046 3563 2047 3567
rect 2051 3563 2052 3567
rect 3914 3567 3915 3571
rect 3919 3567 3920 3571
rect 3914 3566 3920 3567
rect 3942 3567 3948 3568
rect 2046 3562 2052 3563
rect 2102 3564 2108 3565
rect 2102 3560 2103 3564
rect 2107 3560 2108 3564
rect 1066 3558 1072 3559
rect 2006 3559 2012 3560
rect 2102 3559 2108 3560
rect 2278 3564 2284 3565
rect 2278 3560 2279 3564
rect 2283 3560 2284 3564
rect 2278 3559 2284 3560
rect 2470 3564 2476 3565
rect 2470 3560 2471 3564
rect 2475 3560 2476 3564
rect 2470 3559 2476 3560
rect 2670 3564 2676 3565
rect 2670 3560 2671 3564
rect 2675 3560 2676 3564
rect 2670 3559 2676 3560
rect 2870 3564 2876 3565
rect 2870 3560 2871 3564
rect 2875 3560 2876 3564
rect 2870 3559 2876 3560
rect 3062 3564 3068 3565
rect 3062 3560 3063 3564
rect 3067 3560 3068 3564
rect 3062 3559 3068 3560
rect 3254 3564 3260 3565
rect 3254 3560 3255 3564
rect 3259 3560 3260 3564
rect 3254 3559 3260 3560
rect 3446 3564 3452 3565
rect 3446 3560 3447 3564
rect 3451 3560 3452 3564
rect 3446 3559 3452 3560
rect 3638 3564 3644 3565
rect 3638 3560 3639 3564
rect 3643 3560 3644 3564
rect 3638 3559 3644 3560
rect 3838 3564 3844 3565
rect 3838 3560 3839 3564
rect 3843 3560 3844 3564
rect 3942 3563 3943 3567
rect 3947 3563 3948 3567
rect 3942 3562 3948 3563
rect 3838 3559 3844 3560
rect 110 3554 116 3555
rect 166 3556 172 3557
rect 166 3552 167 3556
rect 171 3552 172 3556
rect 166 3551 172 3552
rect 358 3556 364 3557
rect 358 3552 359 3556
rect 363 3552 364 3556
rect 358 3551 364 3552
rect 558 3556 564 3557
rect 558 3552 559 3556
rect 563 3552 564 3556
rect 558 3551 564 3552
rect 774 3556 780 3557
rect 774 3552 775 3556
rect 779 3552 780 3556
rect 774 3551 780 3552
rect 990 3556 996 3557
rect 990 3552 991 3556
rect 995 3552 996 3556
rect 990 3551 996 3552
rect 1214 3556 1220 3557
rect 1214 3552 1215 3556
rect 1219 3552 1220 3556
rect 1214 3551 1220 3552
rect 1446 3556 1452 3557
rect 1446 3552 1447 3556
rect 1451 3552 1452 3556
rect 1446 3551 1452 3552
rect 1686 3556 1692 3557
rect 1686 3552 1687 3556
rect 1691 3552 1692 3556
rect 2006 3555 2007 3559
rect 2011 3555 2012 3559
rect 2006 3554 2012 3555
rect 1686 3551 1692 3552
rect 2326 3500 2332 3501
rect 2046 3497 2052 3498
rect 2046 3493 2047 3497
rect 2051 3493 2052 3497
rect 2326 3496 2327 3500
rect 2331 3496 2332 3500
rect 2326 3495 2332 3496
rect 2446 3500 2452 3501
rect 2446 3496 2447 3500
rect 2451 3496 2452 3500
rect 2446 3495 2452 3496
rect 2582 3500 2588 3501
rect 2582 3496 2583 3500
rect 2587 3496 2588 3500
rect 2582 3495 2588 3496
rect 2734 3500 2740 3501
rect 2734 3496 2735 3500
rect 2739 3496 2740 3500
rect 2734 3495 2740 3496
rect 2910 3500 2916 3501
rect 2910 3496 2911 3500
rect 2915 3496 2916 3500
rect 2910 3495 2916 3496
rect 3110 3500 3116 3501
rect 3110 3496 3111 3500
rect 3115 3496 3116 3500
rect 3110 3495 3116 3496
rect 3334 3500 3340 3501
rect 3334 3496 3335 3500
rect 3339 3496 3340 3500
rect 3334 3495 3340 3496
rect 3566 3500 3572 3501
rect 3566 3496 3567 3500
rect 3571 3496 3572 3500
rect 3566 3495 3572 3496
rect 3806 3500 3812 3501
rect 3806 3496 3807 3500
rect 3811 3496 3812 3500
rect 3806 3495 3812 3496
rect 3942 3497 3948 3498
rect 2046 3492 2052 3493
rect 3942 3493 3943 3497
rect 3947 3493 3948 3497
rect 3942 3492 3948 3493
rect 2402 3491 2408 3492
rect 294 3488 300 3489
rect 110 3485 116 3486
rect 110 3481 111 3485
rect 115 3481 116 3485
rect 294 3484 295 3488
rect 299 3484 300 3488
rect 294 3483 300 3484
rect 430 3488 436 3489
rect 430 3484 431 3488
rect 435 3484 436 3488
rect 430 3483 436 3484
rect 582 3488 588 3489
rect 582 3484 583 3488
rect 587 3484 588 3488
rect 582 3483 588 3484
rect 742 3488 748 3489
rect 742 3484 743 3488
rect 747 3484 748 3488
rect 742 3483 748 3484
rect 910 3488 916 3489
rect 910 3484 911 3488
rect 915 3484 916 3488
rect 910 3483 916 3484
rect 1078 3488 1084 3489
rect 1078 3484 1079 3488
rect 1083 3484 1084 3488
rect 1078 3483 1084 3484
rect 1246 3488 1252 3489
rect 1246 3484 1247 3488
rect 1251 3484 1252 3488
rect 1246 3483 1252 3484
rect 1422 3488 1428 3489
rect 1422 3484 1423 3488
rect 1427 3484 1428 3488
rect 1422 3483 1428 3484
rect 1598 3488 1604 3489
rect 1598 3484 1599 3488
rect 1603 3484 1604 3488
rect 1598 3483 1604 3484
rect 1774 3488 1780 3489
rect 1774 3484 1775 3488
rect 1779 3484 1780 3488
rect 2402 3487 2403 3491
rect 2407 3487 2408 3491
rect 2402 3486 2408 3487
rect 2522 3491 2528 3492
rect 2522 3487 2523 3491
rect 2527 3487 2528 3491
rect 2710 3491 2716 3492
rect 2710 3490 2711 3491
rect 2661 3488 2711 3490
rect 2522 3486 2528 3487
rect 2710 3487 2711 3488
rect 2715 3487 2716 3491
rect 2978 3491 2984 3492
rect 2710 3486 2716 3487
rect 2720 3488 2777 3490
rect 1774 3483 1780 3484
rect 2006 3485 2012 3486
rect 110 3480 116 3481
rect 2006 3481 2007 3485
rect 2011 3481 2012 3485
rect 2326 3481 2332 3482
rect 2006 3480 2012 3481
rect 2046 3480 2052 3481
rect 271 3479 277 3480
rect 271 3475 272 3479
rect 276 3478 277 3479
rect 378 3479 384 3480
rect 276 3476 337 3478
rect 276 3475 277 3476
rect 271 3474 277 3475
rect 378 3475 379 3479
rect 383 3478 384 3479
rect 514 3479 520 3480
rect 383 3476 473 3478
rect 383 3475 384 3476
rect 378 3474 384 3475
rect 514 3475 515 3479
rect 519 3478 520 3479
rect 666 3479 672 3480
rect 519 3476 625 3478
rect 519 3475 520 3476
rect 514 3474 520 3475
rect 666 3475 667 3479
rect 671 3478 672 3479
rect 826 3479 832 3480
rect 671 3476 785 3478
rect 671 3475 672 3476
rect 666 3474 672 3475
rect 826 3475 827 3479
rect 831 3478 832 3479
rect 1154 3479 1160 3480
rect 831 3476 953 3478
rect 831 3475 832 3476
rect 826 3474 832 3475
rect 1154 3475 1155 3479
rect 1159 3475 1160 3479
rect 1154 3474 1160 3475
rect 1322 3479 1328 3480
rect 1322 3475 1323 3479
rect 1327 3475 1328 3479
rect 1322 3474 1328 3475
rect 1498 3479 1504 3480
rect 1498 3475 1499 3479
rect 1503 3475 1504 3479
rect 1738 3479 1744 3480
rect 1738 3478 1739 3479
rect 1677 3476 1739 3478
rect 1498 3474 1504 3475
rect 1738 3475 1739 3476
rect 1743 3475 1744 3479
rect 1738 3474 1744 3475
rect 1754 3479 1760 3480
rect 1754 3475 1755 3479
rect 1759 3478 1760 3479
rect 1759 3476 1817 3478
rect 2046 3476 2047 3480
rect 2051 3476 2052 3480
rect 2326 3477 2327 3481
rect 2331 3477 2332 3481
rect 2326 3476 2332 3477
rect 2446 3481 2452 3482
rect 2446 3477 2447 3481
rect 2451 3477 2452 3481
rect 2446 3476 2452 3477
rect 2582 3481 2588 3482
rect 2582 3477 2583 3481
rect 2587 3477 2588 3481
rect 2582 3476 2588 3477
rect 1759 3475 1760 3476
rect 2046 3475 2052 3476
rect 2514 3475 2520 3476
rect 1754 3474 1760 3475
rect 2514 3471 2515 3475
rect 2519 3474 2520 3475
rect 2720 3474 2722 3488
rect 2978 3487 2979 3491
rect 2983 3487 2984 3491
rect 2978 3486 2984 3487
rect 2994 3491 3000 3492
rect 2994 3487 2995 3491
rect 2999 3490 3000 3491
rect 3194 3491 3200 3492
rect 2999 3488 3153 3490
rect 2999 3487 3000 3488
rect 2994 3486 3000 3487
rect 3194 3487 3195 3491
rect 3199 3490 3200 3491
rect 3418 3491 3424 3492
rect 3199 3488 3377 3490
rect 3199 3487 3200 3488
rect 3194 3486 3200 3487
rect 3418 3487 3419 3491
rect 3423 3490 3424 3491
rect 3874 3491 3880 3492
rect 3423 3488 3609 3490
rect 3423 3487 3424 3488
rect 3418 3486 3424 3487
rect 3874 3487 3875 3491
rect 3879 3487 3880 3491
rect 3874 3486 3880 3487
rect 2734 3481 2740 3482
rect 2734 3477 2735 3481
rect 2739 3477 2740 3481
rect 2734 3476 2740 3477
rect 2910 3481 2916 3482
rect 2910 3477 2911 3481
rect 2915 3477 2916 3481
rect 2910 3476 2916 3477
rect 3110 3481 3116 3482
rect 3110 3477 3111 3481
rect 3115 3477 3116 3481
rect 3110 3476 3116 3477
rect 3334 3481 3340 3482
rect 3334 3477 3335 3481
rect 3339 3477 3340 3481
rect 3334 3476 3340 3477
rect 3566 3481 3572 3482
rect 3566 3477 3567 3481
rect 3571 3477 3572 3481
rect 3566 3476 3572 3477
rect 3806 3481 3812 3482
rect 3806 3477 3807 3481
rect 3811 3477 3812 3481
rect 3806 3476 3812 3477
rect 3942 3480 3948 3481
rect 3942 3476 3943 3480
rect 3947 3476 3948 3480
rect 3942 3475 3948 3476
rect 2519 3472 2722 3474
rect 2519 3471 2520 3472
rect 2514 3470 2520 3471
rect 294 3469 300 3470
rect 110 3468 116 3469
rect 110 3464 111 3468
rect 115 3464 116 3468
rect 294 3465 295 3469
rect 299 3465 300 3469
rect 294 3464 300 3465
rect 430 3469 436 3470
rect 430 3465 431 3469
rect 435 3465 436 3469
rect 430 3464 436 3465
rect 582 3469 588 3470
rect 582 3465 583 3469
rect 587 3465 588 3469
rect 582 3464 588 3465
rect 742 3469 748 3470
rect 742 3465 743 3469
rect 747 3465 748 3469
rect 742 3464 748 3465
rect 910 3469 916 3470
rect 910 3465 911 3469
rect 915 3465 916 3469
rect 910 3464 916 3465
rect 1078 3469 1084 3470
rect 1078 3465 1079 3469
rect 1083 3465 1084 3469
rect 1078 3464 1084 3465
rect 1246 3469 1252 3470
rect 1246 3465 1247 3469
rect 1251 3465 1252 3469
rect 1246 3464 1252 3465
rect 1422 3469 1428 3470
rect 1422 3465 1423 3469
rect 1427 3465 1428 3469
rect 1422 3464 1428 3465
rect 1598 3469 1604 3470
rect 1598 3465 1599 3469
rect 1603 3465 1604 3469
rect 1598 3464 1604 3465
rect 1774 3469 1780 3470
rect 1774 3465 1775 3469
rect 1779 3465 1780 3469
rect 1774 3464 1780 3465
rect 2006 3468 2012 3469
rect 2006 3464 2007 3468
rect 2011 3464 2012 3468
rect 2598 3467 2604 3468
rect 2598 3466 2599 3467
rect 110 3463 116 3464
rect 2006 3463 2012 3464
rect 2396 3464 2599 3466
rect 2396 3460 2398 3464
rect 2598 3463 2599 3464
rect 2603 3463 2604 3467
rect 2598 3462 2604 3463
rect 2391 3459 2398 3460
rect 2391 3455 2392 3459
rect 2396 3456 2398 3459
rect 2402 3459 2408 3460
rect 2396 3455 2397 3456
rect 2391 3454 2397 3455
rect 2402 3455 2403 3459
rect 2407 3458 2408 3459
rect 2511 3459 2517 3460
rect 2511 3458 2512 3459
rect 2407 3456 2512 3458
rect 2407 3455 2408 3456
rect 2402 3454 2408 3455
rect 2511 3455 2512 3456
rect 2516 3455 2517 3459
rect 2511 3454 2517 3455
rect 2522 3459 2528 3460
rect 2522 3455 2523 3459
rect 2527 3458 2528 3459
rect 2647 3459 2653 3460
rect 2647 3458 2648 3459
rect 2527 3456 2648 3458
rect 2527 3455 2528 3456
rect 2522 3454 2528 3455
rect 2647 3455 2648 3456
rect 2652 3455 2653 3459
rect 2647 3454 2653 3455
rect 2710 3459 2716 3460
rect 2710 3455 2711 3459
rect 2715 3458 2716 3459
rect 2799 3459 2805 3460
rect 2799 3458 2800 3459
rect 2715 3456 2800 3458
rect 2715 3455 2716 3456
rect 2710 3454 2716 3455
rect 2799 3455 2800 3456
rect 2804 3455 2805 3459
rect 2799 3454 2805 3455
rect 2975 3459 2981 3460
rect 2975 3455 2976 3459
rect 2980 3458 2981 3459
rect 2994 3459 3000 3460
rect 2994 3458 2995 3459
rect 2980 3456 2995 3458
rect 2980 3455 2981 3456
rect 2975 3454 2981 3455
rect 2994 3455 2995 3456
rect 2999 3455 3000 3459
rect 2994 3454 3000 3455
rect 3175 3459 3181 3460
rect 3175 3455 3176 3459
rect 3180 3458 3181 3459
rect 3194 3459 3200 3460
rect 3194 3458 3195 3459
rect 3180 3456 3195 3458
rect 3180 3455 3181 3456
rect 3175 3454 3181 3455
rect 3194 3455 3195 3456
rect 3199 3455 3200 3459
rect 3194 3454 3200 3455
rect 3399 3459 3405 3460
rect 3399 3455 3400 3459
rect 3404 3458 3405 3459
rect 3418 3459 3424 3460
rect 3418 3458 3419 3459
rect 3404 3456 3419 3458
rect 3404 3455 3405 3456
rect 3399 3454 3405 3455
rect 3418 3455 3419 3456
rect 3423 3455 3424 3459
rect 3418 3454 3424 3455
rect 3631 3459 3637 3460
rect 3631 3455 3632 3459
rect 3636 3458 3637 3459
rect 3642 3459 3648 3460
rect 3642 3458 3643 3459
rect 3636 3456 3643 3458
rect 3636 3455 3637 3456
rect 3631 3454 3637 3455
rect 3642 3455 3643 3456
rect 3647 3455 3648 3459
rect 3642 3454 3648 3455
rect 3871 3459 3877 3460
rect 3871 3455 3872 3459
rect 3876 3458 3877 3459
rect 3914 3459 3920 3460
rect 3914 3458 3915 3459
rect 3876 3456 3915 3458
rect 3876 3455 3877 3456
rect 3871 3454 3877 3455
rect 3914 3455 3915 3456
rect 3919 3455 3920 3459
rect 3914 3454 3920 3455
rect 359 3447 365 3448
rect 359 3443 360 3447
rect 364 3446 365 3447
rect 378 3447 384 3448
rect 378 3446 379 3447
rect 364 3444 379 3446
rect 364 3443 365 3444
rect 359 3442 365 3443
rect 378 3443 379 3444
rect 383 3443 384 3447
rect 378 3442 384 3443
rect 495 3447 501 3448
rect 495 3443 496 3447
rect 500 3446 501 3447
rect 514 3447 520 3448
rect 514 3446 515 3447
rect 500 3444 515 3446
rect 500 3443 501 3444
rect 495 3442 501 3443
rect 514 3443 515 3444
rect 519 3443 520 3447
rect 514 3442 520 3443
rect 647 3447 653 3448
rect 647 3443 648 3447
rect 652 3446 653 3447
rect 666 3447 672 3448
rect 666 3446 667 3447
rect 652 3444 667 3446
rect 652 3443 653 3444
rect 647 3442 653 3443
rect 666 3443 667 3444
rect 671 3443 672 3447
rect 666 3442 672 3443
rect 807 3447 813 3448
rect 807 3443 808 3447
rect 812 3446 813 3447
rect 826 3447 832 3448
rect 826 3446 827 3447
rect 812 3444 827 3446
rect 812 3443 813 3444
rect 807 3442 813 3443
rect 826 3443 827 3444
rect 831 3443 832 3447
rect 826 3442 832 3443
rect 975 3447 981 3448
rect 975 3443 976 3447
rect 980 3446 981 3447
rect 1034 3447 1040 3448
rect 1034 3446 1035 3447
rect 980 3444 1035 3446
rect 980 3443 981 3444
rect 975 3442 981 3443
rect 1034 3443 1035 3444
rect 1039 3443 1040 3447
rect 1034 3442 1040 3443
rect 1066 3447 1072 3448
rect 1066 3443 1067 3447
rect 1071 3446 1072 3447
rect 1143 3447 1149 3448
rect 1143 3446 1144 3447
rect 1071 3444 1144 3446
rect 1071 3443 1072 3444
rect 1066 3442 1072 3443
rect 1143 3443 1144 3444
rect 1148 3443 1149 3447
rect 1143 3442 1149 3443
rect 1154 3447 1160 3448
rect 1154 3443 1155 3447
rect 1159 3446 1160 3447
rect 1311 3447 1317 3448
rect 1311 3446 1312 3447
rect 1159 3444 1312 3446
rect 1159 3443 1160 3444
rect 1154 3442 1160 3443
rect 1311 3443 1312 3444
rect 1316 3443 1317 3447
rect 1311 3442 1317 3443
rect 1322 3447 1328 3448
rect 1322 3443 1323 3447
rect 1327 3446 1328 3447
rect 1487 3447 1493 3448
rect 1487 3446 1488 3447
rect 1327 3444 1488 3446
rect 1327 3443 1328 3444
rect 1322 3442 1328 3443
rect 1487 3443 1488 3444
rect 1492 3443 1493 3447
rect 1487 3442 1493 3443
rect 1663 3447 1669 3448
rect 1663 3443 1664 3447
rect 1668 3446 1669 3447
rect 1714 3447 1720 3448
rect 1714 3446 1715 3447
rect 1668 3444 1715 3446
rect 1668 3443 1669 3444
rect 1663 3442 1669 3443
rect 1714 3443 1715 3444
rect 1719 3443 1720 3447
rect 1714 3442 1720 3443
rect 1738 3447 1744 3448
rect 1738 3443 1739 3447
rect 1743 3446 1744 3447
rect 1839 3447 1845 3448
rect 1839 3446 1840 3447
rect 1743 3444 1840 3446
rect 1743 3443 1744 3444
rect 1738 3442 1744 3443
rect 1839 3443 1840 3444
rect 1844 3443 1845 3447
rect 1839 3442 1845 3443
rect 2511 3447 2520 3448
rect 2511 3443 2512 3447
rect 2519 3443 2520 3447
rect 2511 3442 2520 3443
rect 2522 3447 2528 3448
rect 2522 3443 2523 3447
rect 2527 3446 2528 3447
rect 2615 3447 2621 3448
rect 2615 3446 2616 3447
rect 2527 3444 2616 3446
rect 2527 3443 2528 3444
rect 2522 3442 2528 3443
rect 2615 3443 2616 3444
rect 2620 3443 2621 3447
rect 2615 3442 2621 3443
rect 2626 3447 2632 3448
rect 2626 3443 2627 3447
rect 2631 3446 2632 3447
rect 2727 3447 2733 3448
rect 2727 3446 2728 3447
rect 2631 3444 2728 3446
rect 2631 3443 2632 3444
rect 2626 3442 2632 3443
rect 2727 3443 2728 3444
rect 2732 3443 2733 3447
rect 2727 3442 2733 3443
rect 2750 3447 2756 3448
rect 2750 3443 2751 3447
rect 2755 3446 2756 3447
rect 2839 3447 2845 3448
rect 2839 3446 2840 3447
rect 2755 3444 2840 3446
rect 2755 3443 2756 3444
rect 2750 3442 2756 3443
rect 2839 3443 2840 3444
rect 2844 3443 2845 3447
rect 2839 3442 2845 3443
rect 2850 3447 2856 3448
rect 2850 3443 2851 3447
rect 2855 3446 2856 3447
rect 2967 3447 2973 3448
rect 2967 3446 2968 3447
rect 2855 3444 2968 3446
rect 2855 3443 2856 3444
rect 2850 3442 2856 3443
rect 2967 3443 2968 3444
rect 2972 3443 2973 3447
rect 2967 3442 2973 3443
rect 3111 3447 3117 3448
rect 3111 3443 3112 3447
rect 3116 3446 3117 3447
rect 3122 3447 3128 3448
rect 3116 3443 3118 3446
rect 3111 3442 3118 3443
rect 3122 3443 3123 3447
rect 3127 3446 3128 3447
rect 3271 3447 3277 3448
rect 3271 3446 3272 3447
rect 3127 3444 3272 3446
rect 3127 3443 3128 3444
rect 3122 3442 3128 3443
rect 3271 3443 3272 3444
rect 3276 3443 3277 3447
rect 3271 3442 3277 3443
rect 3282 3447 3288 3448
rect 3282 3443 3283 3447
rect 3287 3446 3288 3447
rect 3447 3447 3453 3448
rect 3447 3446 3448 3447
rect 3287 3444 3448 3446
rect 3287 3443 3288 3444
rect 3282 3442 3288 3443
rect 3447 3443 3448 3444
rect 3452 3443 3453 3447
rect 3447 3442 3453 3443
rect 3458 3447 3464 3448
rect 3458 3443 3459 3447
rect 3463 3446 3464 3447
rect 3631 3447 3637 3448
rect 3631 3446 3632 3447
rect 3463 3444 3632 3446
rect 3463 3443 3464 3444
rect 3458 3442 3464 3443
rect 3631 3443 3632 3444
rect 3636 3443 3637 3447
rect 3631 3442 3637 3443
rect 3815 3447 3821 3448
rect 3815 3443 3816 3447
rect 3820 3446 3821 3447
rect 3874 3447 3880 3448
rect 3874 3446 3875 3447
rect 3820 3444 3875 3446
rect 3820 3443 3821 3444
rect 3815 3442 3821 3443
rect 3874 3443 3875 3444
rect 3879 3443 3880 3447
rect 3874 3442 3880 3443
rect 3116 3438 3118 3442
rect 3258 3439 3264 3440
rect 3258 3438 3259 3439
rect 3116 3436 3259 3438
rect 3258 3435 3259 3436
rect 3263 3435 3264 3439
rect 3258 3434 3264 3435
rect 2046 3428 2052 3429
rect 3942 3428 3948 3429
rect 2046 3424 2047 3428
rect 2051 3424 2052 3428
rect 2046 3423 2052 3424
rect 2446 3427 2452 3428
rect 2446 3423 2447 3427
rect 2451 3423 2452 3427
rect 2446 3422 2452 3423
rect 2550 3427 2556 3428
rect 2550 3423 2551 3427
rect 2555 3423 2556 3427
rect 2550 3422 2556 3423
rect 2662 3427 2668 3428
rect 2662 3423 2663 3427
rect 2667 3423 2668 3427
rect 2662 3422 2668 3423
rect 2774 3427 2780 3428
rect 2774 3423 2775 3427
rect 2779 3423 2780 3427
rect 2774 3422 2780 3423
rect 2902 3427 2908 3428
rect 2902 3423 2903 3427
rect 2907 3423 2908 3427
rect 2902 3422 2908 3423
rect 3046 3427 3052 3428
rect 3046 3423 3047 3427
rect 3051 3423 3052 3427
rect 3046 3422 3052 3423
rect 3206 3427 3212 3428
rect 3206 3423 3207 3427
rect 3211 3423 3212 3427
rect 3206 3422 3212 3423
rect 3382 3427 3388 3428
rect 3382 3423 3383 3427
rect 3387 3423 3388 3427
rect 3382 3422 3388 3423
rect 3566 3427 3572 3428
rect 3566 3423 3567 3427
rect 3571 3423 3572 3427
rect 3566 3422 3572 3423
rect 3750 3427 3756 3428
rect 3750 3423 3751 3427
rect 3755 3423 3756 3427
rect 3942 3424 3943 3428
rect 3947 3424 3948 3428
rect 3942 3423 3948 3424
rect 3750 3422 3756 3423
rect 2522 3419 2528 3420
rect 559 3415 565 3416
rect 559 3411 560 3415
rect 564 3414 565 3415
rect 618 3415 624 3416
rect 618 3414 619 3415
rect 564 3412 619 3414
rect 564 3411 565 3412
rect 559 3410 565 3411
rect 618 3411 619 3412
rect 623 3411 624 3415
rect 618 3410 624 3411
rect 626 3415 632 3416
rect 626 3411 627 3415
rect 631 3414 632 3415
rect 711 3415 717 3416
rect 711 3414 712 3415
rect 631 3412 712 3414
rect 631 3411 632 3412
rect 626 3410 632 3411
rect 711 3411 712 3412
rect 716 3411 717 3415
rect 711 3410 717 3411
rect 722 3415 728 3416
rect 722 3411 723 3415
rect 727 3414 728 3415
rect 863 3415 869 3416
rect 863 3414 864 3415
rect 727 3412 864 3414
rect 727 3411 728 3412
rect 722 3410 728 3411
rect 863 3411 864 3412
rect 868 3411 869 3415
rect 863 3410 869 3411
rect 874 3415 880 3416
rect 874 3411 875 3415
rect 879 3414 880 3415
rect 1023 3415 1029 3416
rect 1023 3414 1024 3415
rect 879 3412 1024 3414
rect 879 3411 880 3412
rect 874 3410 880 3411
rect 1023 3411 1024 3412
rect 1028 3411 1029 3415
rect 1023 3410 1029 3411
rect 1191 3415 1197 3416
rect 1191 3411 1192 3415
rect 1196 3414 1197 3415
rect 1215 3415 1221 3416
rect 1215 3414 1216 3415
rect 1196 3412 1216 3414
rect 1196 3411 1197 3412
rect 1191 3410 1197 3411
rect 1215 3411 1216 3412
rect 1220 3411 1221 3415
rect 1215 3410 1221 3411
rect 1359 3415 1365 3416
rect 1359 3411 1360 3415
rect 1364 3414 1365 3415
rect 1383 3415 1389 3416
rect 1383 3414 1384 3415
rect 1364 3412 1384 3414
rect 1364 3411 1365 3412
rect 1359 3410 1365 3411
rect 1383 3411 1384 3412
rect 1388 3411 1389 3415
rect 1383 3410 1389 3411
rect 1498 3415 1504 3416
rect 1498 3411 1499 3415
rect 1503 3414 1504 3415
rect 1527 3415 1533 3416
rect 1527 3414 1528 3415
rect 1503 3412 1528 3414
rect 1503 3411 1504 3412
rect 1498 3410 1504 3411
rect 1527 3411 1528 3412
rect 1532 3411 1533 3415
rect 1527 3410 1533 3411
rect 1703 3415 1709 3416
rect 1703 3411 1704 3415
rect 1708 3414 1709 3415
rect 1722 3415 1728 3416
rect 1722 3414 1723 3415
rect 1708 3412 1723 3414
rect 1708 3411 1709 3412
rect 1703 3410 1709 3411
rect 1722 3411 1723 3412
rect 1727 3411 1728 3415
rect 1722 3410 1728 3411
rect 1879 3415 1885 3416
rect 1879 3411 1880 3415
rect 1884 3414 1885 3415
rect 1898 3415 1904 3416
rect 1898 3414 1899 3415
rect 1884 3412 1899 3414
rect 1884 3411 1885 3412
rect 1879 3410 1885 3411
rect 1898 3411 1899 3412
rect 1903 3411 1904 3415
rect 2522 3415 2523 3419
rect 2527 3415 2528 3419
rect 2522 3414 2528 3415
rect 2626 3419 2632 3420
rect 2626 3415 2627 3419
rect 2631 3415 2632 3419
rect 2750 3419 2756 3420
rect 2750 3418 2751 3419
rect 2741 3416 2751 3418
rect 2626 3414 2632 3415
rect 2750 3415 2751 3416
rect 2755 3415 2756 3419
rect 2750 3414 2756 3415
rect 2850 3419 2856 3420
rect 2850 3415 2851 3419
rect 2855 3415 2856 3419
rect 3122 3419 3128 3420
rect 2850 3414 2856 3415
rect 2978 3415 2984 3416
rect 1898 3410 1904 3411
rect 2046 3411 2052 3412
rect 2046 3407 2047 3411
rect 2051 3407 2052 3411
rect 2978 3411 2979 3415
rect 2983 3411 2984 3415
rect 3122 3415 3123 3419
rect 3127 3415 3128 3419
rect 3122 3414 3128 3415
rect 3282 3419 3288 3420
rect 3282 3415 3283 3419
rect 3287 3415 3288 3419
rect 3282 3414 3288 3415
rect 3458 3419 3464 3420
rect 3458 3415 3459 3419
rect 3463 3415 3464 3419
rect 3458 3414 3464 3415
rect 3642 3419 3648 3420
rect 3642 3415 3643 3419
rect 3647 3415 3648 3419
rect 3642 3414 3648 3415
rect 3826 3415 3832 3416
rect 2978 3410 2984 3411
rect 3826 3411 3827 3415
rect 3831 3411 3832 3415
rect 3826 3410 3832 3411
rect 3942 3411 3948 3412
rect 2046 3406 2052 3407
rect 2446 3408 2452 3409
rect 2446 3404 2447 3408
rect 2451 3404 2452 3408
rect 2446 3403 2452 3404
rect 2550 3408 2556 3409
rect 2550 3404 2551 3408
rect 2555 3404 2556 3408
rect 2550 3403 2556 3404
rect 2662 3408 2668 3409
rect 2662 3404 2663 3408
rect 2667 3404 2668 3408
rect 2662 3403 2668 3404
rect 2774 3408 2780 3409
rect 2774 3404 2775 3408
rect 2779 3404 2780 3408
rect 2774 3403 2780 3404
rect 2902 3408 2908 3409
rect 2902 3404 2903 3408
rect 2907 3404 2908 3408
rect 2902 3403 2908 3404
rect 3046 3408 3052 3409
rect 3046 3404 3047 3408
rect 3051 3404 3052 3408
rect 3046 3403 3052 3404
rect 3206 3408 3212 3409
rect 3206 3404 3207 3408
rect 3211 3404 3212 3408
rect 3206 3403 3212 3404
rect 3382 3408 3388 3409
rect 3382 3404 3383 3408
rect 3387 3404 3388 3408
rect 3382 3403 3388 3404
rect 3566 3408 3572 3409
rect 3566 3404 3567 3408
rect 3571 3404 3572 3408
rect 3566 3403 3572 3404
rect 3750 3408 3756 3409
rect 3750 3404 3751 3408
rect 3755 3404 3756 3408
rect 3942 3407 3943 3411
rect 3947 3407 3948 3411
rect 3942 3406 3948 3407
rect 3750 3403 3756 3404
rect 110 3396 116 3397
rect 2006 3396 2012 3397
rect 110 3392 111 3396
rect 115 3392 116 3396
rect 110 3391 116 3392
rect 494 3395 500 3396
rect 494 3391 495 3395
rect 499 3391 500 3395
rect 494 3390 500 3391
rect 646 3395 652 3396
rect 646 3391 647 3395
rect 651 3391 652 3395
rect 646 3390 652 3391
rect 798 3395 804 3396
rect 798 3391 799 3395
rect 803 3391 804 3395
rect 798 3390 804 3391
rect 958 3395 964 3396
rect 958 3391 959 3395
rect 963 3391 964 3395
rect 958 3390 964 3391
rect 1126 3395 1132 3396
rect 1126 3391 1127 3395
rect 1131 3391 1132 3395
rect 1126 3390 1132 3391
rect 1294 3395 1300 3396
rect 1294 3391 1295 3395
rect 1299 3391 1300 3395
rect 1294 3390 1300 3391
rect 1462 3395 1468 3396
rect 1462 3391 1463 3395
rect 1467 3391 1468 3395
rect 1462 3390 1468 3391
rect 1638 3395 1644 3396
rect 1638 3391 1639 3395
rect 1643 3391 1644 3395
rect 1638 3390 1644 3391
rect 1814 3395 1820 3396
rect 1814 3391 1815 3395
rect 1819 3391 1820 3395
rect 2006 3392 2007 3396
rect 2011 3392 2012 3396
rect 2006 3391 2012 3392
rect 1814 3390 1820 3391
rect 626 3387 632 3388
rect 626 3386 627 3387
rect 573 3384 627 3386
rect 626 3383 627 3384
rect 631 3383 632 3387
rect 626 3382 632 3383
rect 722 3387 728 3388
rect 722 3383 723 3387
rect 727 3383 728 3387
rect 722 3382 728 3383
rect 874 3387 880 3388
rect 874 3383 875 3387
rect 879 3383 880 3387
rect 874 3382 880 3383
rect 1034 3387 1040 3388
rect 1034 3383 1035 3387
rect 1039 3383 1040 3387
rect 1215 3387 1221 3388
rect 1034 3382 1040 3383
rect 1202 3383 1208 3384
rect 110 3379 116 3380
rect 110 3375 111 3379
rect 115 3375 116 3379
rect 1202 3379 1203 3383
rect 1207 3379 1208 3383
rect 1215 3383 1216 3387
rect 1220 3386 1221 3387
rect 1383 3387 1389 3388
rect 1220 3384 1337 3386
rect 1220 3383 1221 3384
rect 1215 3382 1221 3383
rect 1383 3383 1384 3387
rect 1388 3386 1389 3387
rect 1714 3387 1720 3388
rect 1388 3384 1505 3386
rect 1388 3383 1389 3384
rect 1383 3382 1389 3383
rect 1714 3383 1715 3387
rect 1719 3383 1720 3387
rect 1714 3382 1720 3383
rect 1722 3387 1728 3388
rect 1722 3383 1723 3387
rect 1727 3386 1728 3387
rect 1727 3384 1857 3386
rect 1727 3383 1728 3384
rect 1722 3382 1728 3383
rect 1202 3378 1208 3379
rect 2006 3379 2012 3380
rect 110 3374 116 3375
rect 494 3376 500 3377
rect 494 3372 495 3376
rect 499 3372 500 3376
rect 494 3371 500 3372
rect 646 3376 652 3377
rect 646 3372 647 3376
rect 651 3372 652 3376
rect 646 3371 652 3372
rect 798 3376 804 3377
rect 798 3372 799 3376
rect 803 3372 804 3376
rect 798 3371 804 3372
rect 958 3376 964 3377
rect 958 3372 959 3376
rect 963 3372 964 3376
rect 958 3371 964 3372
rect 1126 3376 1132 3377
rect 1126 3372 1127 3376
rect 1131 3372 1132 3376
rect 1126 3371 1132 3372
rect 1294 3376 1300 3377
rect 1294 3372 1295 3376
rect 1299 3372 1300 3376
rect 1294 3371 1300 3372
rect 1462 3376 1468 3377
rect 1462 3372 1463 3376
rect 1467 3372 1468 3376
rect 1462 3371 1468 3372
rect 1638 3376 1644 3377
rect 1638 3372 1639 3376
rect 1643 3372 1644 3376
rect 1638 3371 1644 3372
rect 1814 3376 1820 3377
rect 1814 3372 1815 3376
rect 1819 3372 1820 3376
rect 2006 3375 2007 3379
rect 2011 3375 2012 3379
rect 2006 3374 2012 3375
rect 1814 3371 1820 3372
rect 2566 3336 2572 3337
rect 2046 3333 2052 3334
rect 2046 3329 2047 3333
rect 2051 3329 2052 3333
rect 2566 3332 2567 3336
rect 2571 3332 2572 3336
rect 2566 3331 2572 3332
rect 2718 3336 2724 3337
rect 2718 3332 2719 3336
rect 2723 3332 2724 3336
rect 2718 3331 2724 3332
rect 2870 3336 2876 3337
rect 2870 3332 2871 3336
rect 2875 3332 2876 3336
rect 2870 3331 2876 3332
rect 3022 3336 3028 3337
rect 3022 3332 3023 3336
rect 3027 3332 3028 3336
rect 3022 3331 3028 3332
rect 3174 3336 3180 3337
rect 3174 3332 3175 3336
rect 3179 3332 3180 3336
rect 3174 3331 3180 3332
rect 3326 3336 3332 3337
rect 3326 3332 3327 3336
rect 3331 3332 3332 3336
rect 3326 3331 3332 3332
rect 3478 3336 3484 3337
rect 3478 3332 3479 3336
rect 3483 3332 3484 3336
rect 3478 3331 3484 3332
rect 3630 3336 3636 3337
rect 3630 3332 3631 3336
rect 3635 3332 3636 3336
rect 3630 3331 3636 3332
rect 3782 3336 3788 3337
rect 3782 3332 3783 3336
rect 3787 3332 3788 3336
rect 3782 3331 3788 3332
rect 3942 3333 3948 3334
rect 2046 3328 2052 3329
rect 3942 3329 3943 3333
rect 3947 3329 3948 3333
rect 3942 3328 3948 3329
rect 2642 3327 2648 3328
rect 2642 3323 2643 3327
rect 2647 3323 2648 3327
rect 2642 3322 2648 3323
rect 2650 3327 2656 3328
rect 2650 3323 2651 3327
rect 2655 3326 2656 3327
rect 2802 3327 2808 3328
rect 2655 3324 2761 3326
rect 2655 3323 2656 3324
rect 2650 3322 2656 3323
rect 2802 3323 2803 3327
rect 2807 3326 2808 3327
rect 2954 3327 2960 3328
rect 2807 3324 2913 3326
rect 2807 3323 2808 3324
rect 2802 3322 2808 3323
rect 2954 3323 2955 3327
rect 2959 3326 2960 3327
rect 3250 3327 3256 3328
rect 2959 3324 3065 3326
rect 2959 3323 2960 3324
rect 2954 3322 2960 3323
rect 3250 3323 3251 3327
rect 3255 3323 3256 3327
rect 3250 3322 3256 3323
rect 3258 3327 3264 3328
rect 3258 3323 3259 3327
rect 3263 3326 3264 3327
rect 3455 3327 3461 3328
rect 3263 3324 3369 3326
rect 3263 3323 3264 3324
rect 3258 3322 3264 3323
rect 3455 3323 3456 3327
rect 3460 3326 3461 3327
rect 3562 3327 3568 3328
rect 3460 3324 3521 3326
rect 3460 3323 3461 3324
rect 3455 3322 3461 3323
rect 3562 3323 3563 3327
rect 3567 3326 3568 3327
rect 3714 3327 3720 3328
rect 3567 3324 3673 3326
rect 3567 3323 3568 3324
rect 3562 3322 3568 3323
rect 3714 3323 3715 3327
rect 3719 3326 3720 3327
rect 3719 3324 3825 3326
rect 3719 3323 3720 3324
rect 3714 3322 3720 3323
rect 2566 3317 2572 3318
rect 2046 3316 2052 3317
rect 2046 3312 2047 3316
rect 2051 3312 2052 3316
rect 2566 3313 2567 3317
rect 2571 3313 2572 3317
rect 2566 3312 2572 3313
rect 2718 3317 2724 3318
rect 2718 3313 2719 3317
rect 2723 3313 2724 3317
rect 2718 3312 2724 3313
rect 2870 3317 2876 3318
rect 2870 3313 2871 3317
rect 2875 3313 2876 3317
rect 2870 3312 2876 3313
rect 3022 3317 3028 3318
rect 3022 3313 3023 3317
rect 3027 3313 3028 3317
rect 3022 3312 3028 3313
rect 3174 3317 3180 3318
rect 3174 3313 3175 3317
rect 3179 3313 3180 3317
rect 3174 3312 3180 3313
rect 3326 3317 3332 3318
rect 3326 3313 3327 3317
rect 3331 3313 3332 3317
rect 3326 3312 3332 3313
rect 3478 3317 3484 3318
rect 3478 3313 3479 3317
rect 3483 3313 3484 3317
rect 3478 3312 3484 3313
rect 3630 3317 3636 3318
rect 3630 3313 3631 3317
rect 3635 3313 3636 3317
rect 3630 3312 3636 3313
rect 3782 3317 3788 3318
rect 3782 3313 3783 3317
rect 3787 3313 3788 3317
rect 3782 3312 3788 3313
rect 3942 3316 3948 3317
rect 3942 3312 3943 3316
rect 3947 3312 3948 3316
rect 2046 3311 2052 3312
rect 3942 3311 3948 3312
rect 134 3304 140 3305
rect 110 3301 116 3302
rect 110 3297 111 3301
rect 115 3297 116 3301
rect 134 3300 135 3304
rect 139 3300 140 3304
rect 134 3299 140 3300
rect 294 3304 300 3305
rect 294 3300 295 3304
rect 299 3300 300 3304
rect 294 3299 300 3300
rect 478 3304 484 3305
rect 478 3300 479 3304
rect 483 3300 484 3304
rect 478 3299 484 3300
rect 670 3304 676 3305
rect 670 3300 671 3304
rect 675 3300 676 3304
rect 670 3299 676 3300
rect 862 3304 868 3305
rect 862 3300 863 3304
rect 867 3300 868 3304
rect 862 3299 868 3300
rect 1054 3304 1060 3305
rect 1054 3300 1055 3304
rect 1059 3300 1060 3304
rect 1054 3299 1060 3300
rect 1246 3304 1252 3305
rect 1246 3300 1247 3304
rect 1251 3300 1252 3304
rect 1246 3299 1252 3300
rect 1438 3304 1444 3305
rect 1438 3300 1439 3304
rect 1443 3300 1444 3304
rect 1438 3299 1444 3300
rect 1630 3304 1636 3305
rect 1630 3300 1631 3304
rect 1635 3300 1636 3304
rect 1630 3299 1636 3300
rect 1822 3304 1828 3305
rect 1822 3300 1823 3304
rect 1827 3300 1828 3304
rect 1822 3299 1828 3300
rect 2006 3301 2012 3302
rect 110 3296 116 3297
rect 2006 3297 2007 3301
rect 2011 3297 2012 3301
rect 2006 3296 2012 3297
rect 210 3295 216 3296
rect 210 3291 211 3295
rect 215 3291 216 3295
rect 210 3290 216 3291
rect 370 3295 376 3296
rect 370 3291 371 3295
rect 375 3291 376 3295
rect 370 3290 376 3291
rect 386 3295 392 3296
rect 386 3291 387 3295
rect 391 3294 392 3295
rect 618 3295 624 3296
rect 391 3292 521 3294
rect 391 3291 392 3292
rect 386 3290 392 3291
rect 618 3291 619 3295
rect 623 3294 624 3295
rect 754 3295 760 3296
rect 623 3292 713 3294
rect 623 3291 624 3292
rect 618 3290 624 3291
rect 754 3291 755 3295
rect 759 3294 760 3295
rect 1130 3295 1136 3296
rect 759 3292 905 3294
rect 759 3291 760 3292
rect 754 3290 760 3291
rect 1130 3291 1131 3295
rect 1135 3291 1136 3295
rect 1130 3290 1136 3291
rect 1322 3295 1328 3296
rect 1322 3291 1323 3295
rect 1327 3291 1328 3295
rect 1322 3290 1328 3291
rect 1338 3295 1344 3296
rect 1338 3291 1339 3295
rect 1343 3294 1344 3295
rect 1778 3295 1784 3296
rect 1778 3294 1779 3295
rect 1343 3292 1481 3294
rect 1709 3292 1779 3294
rect 1343 3291 1344 3292
rect 1338 3290 1344 3291
rect 1778 3291 1779 3292
rect 1783 3291 1784 3295
rect 1778 3290 1784 3291
rect 1898 3295 1904 3296
rect 1898 3291 1899 3295
rect 1903 3291 1904 3295
rect 1898 3290 1904 3291
rect 2631 3295 2637 3296
rect 2631 3291 2632 3295
rect 2636 3294 2637 3295
rect 2650 3295 2656 3296
rect 2650 3294 2651 3295
rect 2636 3292 2651 3294
rect 2636 3291 2637 3292
rect 2631 3290 2637 3291
rect 2650 3291 2651 3292
rect 2655 3291 2656 3295
rect 2650 3290 2656 3291
rect 2783 3295 2789 3296
rect 2783 3291 2784 3295
rect 2788 3294 2789 3295
rect 2802 3295 2808 3296
rect 2802 3294 2803 3295
rect 2788 3292 2803 3294
rect 2788 3291 2789 3292
rect 2783 3290 2789 3291
rect 2802 3291 2803 3292
rect 2807 3291 2808 3295
rect 2802 3290 2808 3291
rect 2935 3295 2941 3296
rect 2935 3291 2936 3295
rect 2940 3294 2941 3295
rect 2954 3295 2960 3296
rect 2954 3294 2955 3295
rect 2940 3292 2955 3294
rect 2940 3291 2941 3292
rect 2935 3290 2941 3291
rect 2954 3291 2955 3292
rect 2959 3291 2960 3295
rect 2954 3290 2960 3291
rect 2978 3295 2984 3296
rect 2978 3291 2979 3295
rect 2983 3294 2984 3295
rect 3087 3295 3093 3296
rect 3087 3294 3088 3295
rect 2983 3292 3088 3294
rect 2983 3291 2984 3292
rect 2978 3290 2984 3291
rect 3087 3291 3088 3292
rect 3092 3291 3093 3295
rect 3087 3290 3093 3291
rect 3194 3295 3200 3296
rect 3194 3291 3195 3295
rect 3199 3294 3200 3295
rect 3239 3295 3245 3296
rect 3239 3294 3240 3295
rect 3199 3292 3240 3294
rect 3199 3291 3200 3292
rect 3194 3290 3200 3291
rect 3239 3291 3240 3292
rect 3244 3291 3245 3295
rect 3239 3290 3245 3291
rect 3250 3295 3256 3296
rect 3250 3291 3251 3295
rect 3255 3294 3256 3295
rect 3391 3295 3397 3296
rect 3391 3294 3392 3295
rect 3255 3292 3392 3294
rect 3255 3291 3256 3292
rect 3250 3290 3256 3291
rect 3391 3291 3392 3292
rect 3396 3291 3397 3295
rect 3391 3290 3397 3291
rect 3543 3295 3549 3296
rect 3543 3291 3544 3295
rect 3548 3294 3549 3295
rect 3562 3295 3568 3296
rect 3562 3294 3563 3295
rect 3548 3292 3563 3294
rect 3548 3291 3549 3292
rect 3543 3290 3549 3291
rect 3562 3291 3563 3292
rect 3567 3291 3568 3295
rect 3562 3290 3568 3291
rect 3695 3295 3701 3296
rect 3695 3291 3696 3295
rect 3700 3294 3701 3295
rect 3714 3295 3720 3296
rect 3714 3294 3715 3295
rect 3700 3292 3715 3294
rect 3700 3291 3701 3292
rect 3695 3290 3701 3291
rect 3714 3291 3715 3292
rect 3719 3291 3720 3295
rect 3714 3290 3720 3291
rect 3826 3295 3832 3296
rect 3826 3291 3827 3295
rect 3831 3294 3832 3295
rect 3847 3295 3853 3296
rect 3847 3294 3848 3295
rect 3831 3292 3848 3294
rect 3831 3291 3832 3292
rect 3826 3290 3832 3291
rect 3847 3291 3848 3292
rect 3852 3291 3853 3295
rect 3847 3290 3853 3291
rect 134 3285 140 3286
rect 110 3284 116 3285
rect 110 3280 111 3284
rect 115 3280 116 3284
rect 134 3281 135 3285
rect 139 3281 140 3285
rect 134 3280 140 3281
rect 294 3285 300 3286
rect 294 3281 295 3285
rect 299 3281 300 3285
rect 294 3280 300 3281
rect 478 3285 484 3286
rect 478 3281 479 3285
rect 483 3281 484 3285
rect 478 3280 484 3281
rect 670 3285 676 3286
rect 670 3281 671 3285
rect 675 3281 676 3285
rect 670 3280 676 3281
rect 862 3285 868 3286
rect 862 3281 863 3285
rect 867 3281 868 3285
rect 862 3280 868 3281
rect 1054 3285 1060 3286
rect 1054 3281 1055 3285
rect 1059 3281 1060 3285
rect 1054 3280 1060 3281
rect 1246 3285 1252 3286
rect 1246 3281 1247 3285
rect 1251 3281 1252 3285
rect 1246 3280 1252 3281
rect 1438 3285 1444 3286
rect 1438 3281 1439 3285
rect 1443 3281 1444 3285
rect 1438 3280 1444 3281
rect 1630 3285 1636 3286
rect 1630 3281 1631 3285
rect 1635 3281 1636 3285
rect 1630 3280 1636 3281
rect 1822 3285 1828 3286
rect 1822 3281 1823 3285
rect 1827 3281 1828 3285
rect 1822 3280 1828 3281
rect 2006 3284 2012 3285
rect 2006 3280 2007 3284
rect 2011 3280 2012 3284
rect 110 3279 116 3280
rect 2006 3279 2012 3280
rect 2479 3279 2485 3280
rect 2479 3275 2480 3279
rect 2484 3278 2485 3279
rect 2490 3279 2496 3280
rect 2484 3275 2486 3278
rect 2479 3274 2486 3275
rect 2490 3275 2491 3279
rect 2495 3278 2496 3279
rect 2615 3279 2621 3280
rect 2615 3278 2616 3279
rect 2495 3276 2616 3278
rect 2495 3275 2496 3276
rect 2490 3274 2496 3275
rect 2615 3275 2616 3276
rect 2620 3275 2621 3279
rect 2615 3274 2621 3275
rect 2642 3279 2648 3280
rect 2642 3275 2643 3279
rect 2647 3278 2648 3279
rect 2751 3279 2757 3280
rect 2751 3278 2752 3279
rect 2647 3276 2752 3278
rect 2647 3275 2648 3276
rect 2642 3274 2648 3275
rect 2751 3275 2752 3276
rect 2756 3275 2757 3279
rect 2751 3274 2757 3275
rect 2762 3279 2768 3280
rect 2762 3275 2763 3279
rect 2767 3278 2768 3279
rect 2895 3279 2901 3280
rect 2895 3278 2896 3279
rect 2767 3276 2896 3278
rect 2767 3275 2768 3276
rect 2762 3274 2768 3275
rect 2895 3275 2896 3276
rect 2900 3275 2901 3279
rect 2895 3274 2901 3275
rect 2906 3279 2912 3280
rect 2906 3275 2907 3279
rect 2911 3278 2912 3279
rect 3039 3279 3045 3280
rect 3039 3278 3040 3279
rect 2911 3276 3040 3278
rect 2911 3275 2912 3276
rect 2906 3274 2912 3275
rect 3039 3275 3040 3276
rect 3044 3275 3045 3279
rect 3039 3274 3045 3275
rect 3183 3279 3189 3280
rect 3183 3275 3184 3279
rect 3188 3278 3189 3279
rect 3207 3279 3213 3280
rect 3207 3278 3208 3279
rect 3188 3276 3208 3278
rect 3188 3275 3189 3276
rect 3183 3274 3189 3275
rect 3207 3275 3208 3276
rect 3212 3275 3213 3279
rect 3207 3274 3213 3275
rect 3319 3279 3325 3280
rect 3319 3275 3320 3279
rect 3324 3278 3325 3279
rect 3374 3279 3380 3280
rect 3374 3278 3375 3279
rect 3324 3276 3375 3278
rect 3324 3275 3325 3276
rect 3319 3274 3325 3275
rect 3374 3275 3375 3276
rect 3379 3275 3380 3279
rect 3374 3274 3380 3275
rect 3447 3279 3453 3280
rect 3447 3275 3448 3279
rect 3452 3278 3453 3279
rect 3455 3279 3461 3280
rect 3455 3278 3456 3279
rect 3452 3276 3456 3278
rect 3452 3275 3453 3276
rect 3447 3274 3453 3275
rect 3455 3275 3456 3276
rect 3460 3275 3461 3279
rect 3455 3274 3461 3275
rect 3494 3279 3500 3280
rect 3494 3275 3495 3279
rect 3499 3278 3500 3279
rect 3567 3279 3573 3280
rect 3567 3278 3568 3279
rect 3499 3276 3568 3278
rect 3499 3275 3500 3276
rect 3494 3274 3500 3275
rect 3567 3275 3568 3276
rect 3572 3275 3573 3279
rect 3567 3274 3573 3275
rect 3578 3279 3584 3280
rect 3578 3275 3579 3279
rect 3583 3278 3584 3279
rect 3687 3279 3693 3280
rect 3687 3278 3688 3279
rect 3583 3276 3688 3278
rect 3583 3275 3584 3276
rect 3578 3274 3584 3275
rect 3687 3275 3688 3276
rect 3692 3275 3693 3279
rect 3687 3274 3693 3275
rect 3698 3279 3704 3280
rect 3698 3275 3699 3279
rect 3703 3278 3704 3279
rect 3807 3279 3813 3280
rect 3807 3278 3808 3279
rect 3703 3276 3808 3278
rect 3703 3275 3704 3276
rect 3698 3274 3704 3275
rect 3807 3275 3808 3276
rect 3812 3275 3813 3279
rect 3807 3274 3813 3275
rect 3818 3279 3824 3280
rect 3818 3275 3819 3279
rect 3823 3278 3824 3279
rect 3903 3279 3909 3280
rect 3903 3278 3904 3279
rect 3823 3276 3904 3278
rect 3823 3275 3824 3276
rect 3818 3274 3824 3275
rect 3903 3275 3904 3276
rect 3908 3275 3909 3279
rect 3903 3274 3909 3275
rect 1338 3271 1344 3272
rect 1338 3270 1339 3271
rect 1159 3268 1339 3270
rect 210 3263 216 3264
rect 210 3259 211 3263
rect 215 3262 216 3263
rect 359 3263 365 3264
rect 359 3262 360 3263
rect 215 3260 360 3262
rect 215 3259 216 3260
rect 210 3258 216 3259
rect 359 3259 360 3260
rect 364 3259 365 3263
rect 359 3258 365 3259
rect 370 3263 376 3264
rect 370 3259 371 3263
rect 375 3262 376 3263
rect 543 3263 549 3264
rect 543 3262 544 3263
rect 375 3260 544 3262
rect 375 3259 376 3260
rect 370 3258 376 3259
rect 543 3259 544 3260
rect 548 3259 549 3263
rect 543 3258 549 3259
rect 735 3263 741 3264
rect 735 3259 736 3263
rect 740 3262 741 3263
rect 754 3263 760 3264
rect 754 3262 755 3263
rect 740 3260 755 3262
rect 740 3259 741 3260
rect 735 3258 741 3259
rect 754 3259 755 3260
rect 759 3259 760 3263
rect 754 3258 760 3259
rect 927 3263 933 3264
rect 927 3259 928 3263
rect 932 3262 933 3263
rect 986 3263 992 3264
rect 986 3262 987 3263
rect 932 3260 987 3262
rect 932 3259 933 3260
rect 927 3258 933 3259
rect 986 3259 987 3260
rect 991 3259 992 3263
rect 986 3258 992 3259
rect 1119 3263 1125 3264
rect 1119 3259 1120 3263
rect 1124 3262 1125 3263
rect 1159 3262 1161 3268
rect 1338 3267 1339 3268
rect 1343 3267 1344 3271
rect 2484 3270 2486 3274
rect 2926 3271 2932 3272
rect 2926 3270 2927 3271
rect 2484 3268 2927 3270
rect 1338 3266 1344 3267
rect 2926 3267 2927 3268
rect 2931 3267 2932 3271
rect 2926 3266 2932 3267
rect 1124 3260 1161 3262
rect 1202 3263 1208 3264
rect 1124 3259 1125 3260
rect 1119 3258 1125 3259
rect 1202 3259 1203 3263
rect 1207 3262 1208 3263
rect 1311 3263 1317 3264
rect 1311 3262 1312 3263
rect 1207 3260 1312 3262
rect 1207 3259 1208 3260
rect 1202 3258 1208 3259
rect 1311 3259 1312 3260
rect 1316 3259 1317 3263
rect 1311 3258 1317 3259
rect 1322 3263 1328 3264
rect 1322 3259 1323 3263
rect 1327 3262 1328 3263
rect 1503 3263 1509 3264
rect 1503 3262 1504 3263
rect 1327 3260 1504 3262
rect 1327 3259 1328 3260
rect 1322 3258 1328 3259
rect 1503 3259 1504 3260
rect 1508 3259 1509 3263
rect 1503 3258 1509 3259
rect 1695 3263 1701 3264
rect 1695 3259 1696 3263
rect 1700 3262 1701 3263
rect 1706 3263 1712 3264
rect 1706 3262 1707 3263
rect 1700 3260 1707 3262
rect 1700 3259 1701 3260
rect 1695 3258 1701 3259
rect 1706 3259 1707 3260
rect 1711 3259 1712 3263
rect 1706 3258 1712 3259
rect 1778 3263 1784 3264
rect 1778 3259 1779 3263
rect 1783 3262 1784 3263
rect 1887 3263 1893 3264
rect 1887 3262 1888 3263
rect 1783 3260 1888 3262
rect 1783 3259 1784 3260
rect 1778 3258 1784 3259
rect 1887 3259 1888 3260
rect 1892 3259 1893 3263
rect 1887 3258 1893 3259
rect 2046 3260 2052 3261
rect 3942 3260 3948 3261
rect 2046 3256 2047 3260
rect 2051 3256 2052 3260
rect 2046 3255 2052 3256
rect 2414 3259 2420 3260
rect 2414 3255 2415 3259
rect 2419 3255 2420 3259
rect 2414 3254 2420 3255
rect 2550 3259 2556 3260
rect 2550 3255 2551 3259
rect 2555 3255 2556 3259
rect 2550 3254 2556 3255
rect 2686 3259 2692 3260
rect 2686 3255 2687 3259
rect 2691 3255 2692 3259
rect 2686 3254 2692 3255
rect 2830 3259 2836 3260
rect 2830 3255 2831 3259
rect 2835 3255 2836 3259
rect 2830 3254 2836 3255
rect 2974 3259 2980 3260
rect 2974 3255 2975 3259
rect 2979 3255 2980 3259
rect 2974 3254 2980 3255
rect 3118 3259 3124 3260
rect 3118 3255 3119 3259
rect 3123 3255 3124 3259
rect 3118 3254 3124 3255
rect 3254 3259 3260 3260
rect 3254 3255 3255 3259
rect 3259 3255 3260 3259
rect 3254 3254 3260 3255
rect 3382 3259 3388 3260
rect 3382 3255 3383 3259
rect 3387 3255 3388 3259
rect 3382 3254 3388 3255
rect 3502 3259 3508 3260
rect 3502 3255 3503 3259
rect 3507 3255 3508 3259
rect 3502 3254 3508 3255
rect 3622 3259 3628 3260
rect 3622 3255 3623 3259
rect 3627 3255 3628 3259
rect 3622 3254 3628 3255
rect 3742 3259 3748 3260
rect 3742 3255 3743 3259
rect 3747 3255 3748 3259
rect 3742 3254 3748 3255
rect 3838 3259 3844 3260
rect 3838 3255 3839 3259
rect 3843 3255 3844 3259
rect 3942 3256 3943 3260
rect 3947 3256 3948 3260
rect 3942 3255 3948 3256
rect 3838 3254 3844 3255
rect 2490 3251 2496 3252
rect 199 3247 205 3248
rect 199 3243 200 3247
rect 204 3246 205 3247
rect 255 3247 261 3248
rect 255 3246 256 3247
rect 204 3244 256 3246
rect 204 3243 205 3244
rect 199 3242 205 3243
rect 255 3243 256 3244
rect 260 3243 261 3247
rect 255 3242 261 3243
rect 383 3247 392 3248
rect 383 3243 384 3247
rect 391 3243 392 3247
rect 383 3242 392 3243
rect 583 3247 589 3248
rect 583 3243 584 3247
rect 588 3246 589 3247
rect 678 3247 684 3248
rect 678 3246 679 3247
rect 588 3244 679 3246
rect 588 3243 589 3244
rect 583 3242 589 3243
rect 678 3243 679 3244
rect 683 3243 684 3247
rect 678 3242 684 3243
rect 686 3247 692 3248
rect 686 3243 687 3247
rect 691 3246 692 3247
rect 783 3247 789 3248
rect 783 3246 784 3247
rect 691 3244 784 3246
rect 691 3243 692 3244
rect 686 3242 692 3243
rect 783 3243 784 3244
rect 788 3243 789 3247
rect 783 3242 789 3243
rect 794 3247 800 3248
rect 794 3243 795 3247
rect 799 3246 800 3247
rect 975 3247 981 3248
rect 975 3246 976 3247
rect 799 3244 976 3246
rect 799 3243 800 3244
rect 794 3242 800 3243
rect 975 3243 976 3244
rect 980 3243 981 3247
rect 975 3242 981 3243
rect 1130 3247 1136 3248
rect 1130 3243 1131 3247
rect 1135 3246 1136 3247
rect 1159 3247 1165 3248
rect 1159 3246 1160 3247
rect 1135 3244 1160 3246
rect 1135 3243 1136 3244
rect 1130 3242 1136 3243
rect 1159 3243 1160 3244
rect 1164 3243 1165 3247
rect 1159 3242 1165 3243
rect 1170 3247 1176 3248
rect 1170 3243 1171 3247
rect 1175 3246 1176 3247
rect 1335 3247 1341 3248
rect 1335 3246 1336 3247
rect 1175 3244 1336 3246
rect 1175 3243 1176 3244
rect 1170 3242 1176 3243
rect 1335 3243 1336 3244
rect 1340 3243 1341 3247
rect 1335 3242 1341 3243
rect 1346 3247 1352 3248
rect 1346 3243 1347 3247
rect 1351 3246 1352 3247
rect 1511 3247 1517 3248
rect 1511 3246 1512 3247
rect 1351 3244 1512 3246
rect 1351 3243 1352 3244
rect 1346 3242 1352 3243
rect 1511 3243 1512 3244
rect 1516 3243 1517 3247
rect 1511 3242 1517 3243
rect 1650 3247 1656 3248
rect 1650 3243 1651 3247
rect 1655 3246 1656 3247
rect 1687 3247 1693 3248
rect 1687 3246 1688 3247
rect 1655 3244 1688 3246
rect 1655 3243 1656 3244
rect 1650 3242 1656 3243
rect 1687 3243 1688 3244
rect 1692 3243 1693 3247
rect 1687 3242 1693 3243
rect 1698 3247 1704 3248
rect 1698 3243 1699 3247
rect 1703 3246 1704 3247
rect 1863 3247 1869 3248
rect 1863 3246 1864 3247
rect 1703 3244 1864 3246
rect 1703 3243 1704 3244
rect 1698 3242 1704 3243
rect 1863 3243 1864 3244
rect 1868 3243 1869 3247
rect 2490 3247 2491 3251
rect 2495 3247 2496 3251
rect 2762 3251 2768 3252
rect 2490 3246 2496 3247
rect 2626 3247 2632 3248
rect 1863 3242 1869 3243
rect 2046 3243 2052 3244
rect 2046 3239 2047 3243
rect 2051 3239 2052 3243
rect 2626 3243 2627 3247
rect 2631 3243 2632 3247
rect 2762 3247 2763 3251
rect 2767 3247 2768 3251
rect 2762 3246 2768 3247
rect 2906 3251 2912 3252
rect 2906 3247 2907 3251
rect 2911 3247 2912 3251
rect 2906 3246 2912 3247
rect 2926 3251 2932 3252
rect 2926 3247 2927 3251
rect 2931 3250 2932 3251
rect 3194 3251 3200 3252
rect 2931 3248 3017 3250
rect 2931 3247 2932 3248
rect 2926 3246 2932 3247
rect 3194 3247 3195 3251
rect 3199 3247 3200 3251
rect 3194 3246 3200 3247
rect 3207 3251 3213 3252
rect 3207 3247 3208 3251
rect 3212 3250 3213 3251
rect 3494 3251 3500 3252
rect 3494 3250 3495 3251
rect 3212 3248 3297 3250
rect 3461 3248 3495 3250
rect 3212 3247 3213 3248
rect 3207 3246 3213 3247
rect 3494 3247 3495 3248
rect 3499 3247 3500 3251
rect 3494 3246 3500 3247
rect 3578 3251 3584 3252
rect 3578 3247 3579 3251
rect 3583 3247 3584 3251
rect 3578 3246 3584 3247
rect 3698 3251 3704 3252
rect 3698 3247 3699 3251
rect 3703 3247 3704 3251
rect 3698 3246 3704 3247
rect 3818 3251 3824 3252
rect 3818 3247 3819 3251
rect 3823 3247 3824 3251
rect 3818 3246 3824 3247
rect 3914 3247 3920 3248
rect 2626 3242 2632 3243
rect 3914 3243 3915 3247
rect 3919 3243 3920 3247
rect 3914 3242 3920 3243
rect 3942 3243 3948 3244
rect 2046 3238 2052 3239
rect 2414 3240 2420 3241
rect 2414 3236 2415 3240
rect 2419 3236 2420 3240
rect 2414 3235 2420 3236
rect 2550 3240 2556 3241
rect 2550 3236 2551 3240
rect 2555 3236 2556 3240
rect 2550 3235 2556 3236
rect 2686 3240 2692 3241
rect 2686 3236 2687 3240
rect 2691 3236 2692 3240
rect 2686 3235 2692 3236
rect 2830 3240 2836 3241
rect 2830 3236 2831 3240
rect 2835 3236 2836 3240
rect 2830 3235 2836 3236
rect 2974 3240 2980 3241
rect 2974 3236 2975 3240
rect 2979 3236 2980 3240
rect 2974 3235 2980 3236
rect 3118 3240 3124 3241
rect 3118 3236 3119 3240
rect 3123 3236 3124 3240
rect 3118 3235 3124 3236
rect 3254 3240 3260 3241
rect 3254 3236 3255 3240
rect 3259 3236 3260 3240
rect 3254 3235 3260 3236
rect 3382 3240 3388 3241
rect 3382 3236 3383 3240
rect 3387 3236 3388 3240
rect 3382 3235 3388 3236
rect 3502 3240 3508 3241
rect 3502 3236 3503 3240
rect 3507 3236 3508 3240
rect 3502 3235 3508 3236
rect 3622 3240 3628 3241
rect 3622 3236 3623 3240
rect 3627 3236 3628 3240
rect 3622 3235 3628 3236
rect 3742 3240 3748 3241
rect 3742 3236 3743 3240
rect 3747 3236 3748 3240
rect 3742 3235 3748 3236
rect 3838 3240 3844 3241
rect 3838 3236 3839 3240
rect 3843 3236 3844 3240
rect 3942 3239 3943 3243
rect 3947 3239 3948 3243
rect 3942 3238 3948 3239
rect 3838 3235 3844 3236
rect 110 3228 116 3229
rect 2006 3228 2012 3229
rect 110 3224 111 3228
rect 115 3224 116 3228
rect 110 3223 116 3224
rect 134 3227 140 3228
rect 134 3223 135 3227
rect 139 3223 140 3227
rect 134 3222 140 3223
rect 318 3227 324 3228
rect 318 3223 319 3227
rect 323 3223 324 3227
rect 318 3222 324 3223
rect 518 3227 524 3228
rect 518 3223 519 3227
rect 523 3223 524 3227
rect 518 3222 524 3223
rect 718 3227 724 3228
rect 718 3223 719 3227
rect 723 3223 724 3227
rect 718 3222 724 3223
rect 910 3227 916 3228
rect 910 3223 911 3227
rect 915 3223 916 3227
rect 910 3222 916 3223
rect 1094 3227 1100 3228
rect 1094 3223 1095 3227
rect 1099 3223 1100 3227
rect 1094 3222 1100 3223
rect 1270 3227 1276 3228
rect 1270 3223 1271 3227
rect 1275 3223 1276 3227
rect 1270 3222 1276 3223
rect 1446 3227 1452 3228
rect 1446 3223 1447 3227
rect 1451 3223 1452 3227
rect 1446 3222 1452 3223
rect 1622 3227 1628 3228
rect 1622 3223 1623 3227
rect 1627 3223 1628 3227
rect 1622 3222 1628 3223
rect 1798 3227 1804 3228
rect 1798 3223 1799 3227
rect 1803 3223 1804 3227
rect 2006 3224 2007 3228
rect 2011 3224 2012 3228
rect 2006 3223 2012 3224
rect 1798 3222 1804 3223
rect 255 3219 261 3220
rect 210 3215 216 3216
rect 110 3211 116 3212
rect 110 3207 111 3211
rect 115 3207 116 3211
rect 210 3211 211 3215
rect 215 3211 216 3215
rect 255 3215 256 3219
rect 260 3218 261 3219
rect 686 3219 692 3220
rect 686 3218 687 3219
rect 260 3216 361 3218
rect 597 3216 687 3218
rect 260 3215 261 3216
rect 255 3214 261 3215
rect 686 3215 687 3216
rect 691 3215 692 3219
rect 686 3214 692 3215
rect 794 3219 800 3220
rect 794 3215 795 3219
rect 799 3215 800 3219
rect 794 3214 800 3215
rect 986 3219 992 3220
rect 986 3215 987 3219
rect 991 3215 992 3219
rect 986 3214 992 3215
rect 1170 3219 1176 3220
rect 1170 3215 1171 3219
rect 1175 3215 1176 3219
rect 1170 3214 1176 3215
rect 1346 3219 1352 3220
rect 1346 3215 1347 3219
rect 1351 3215 1352 3219
rect 1698 3219 1704 3220
rect 1346 3214 1352 3215
rect 1522 3215 1528 3216
rect 210 3210 216 3211
rect 1522 3211 1523 3215
rect 1527 3211 1528 3215
rect 1698 3215 1699 3219
rect 1703 3215 1704 3219
rect 1698 3214 1704 3215
rect 1706 3219 1712 3220
rect 1706 3215 1707 3219
rect 1711 3218 1712 3219
rect 1711 3216 1841 3218
rect 1711 3215 1712 3216
rect 1706 3214 1712 3215
rect 1522 3210 1528 3211
rect 2006 3211 2012 3212
rect 110 3206 116 3207
rect 134 3208 140 3209
rect 134 3204 135 3208
rect 139 3204 140 3208
rect 134 3203 140 3204
rect 318 3208 324 3209
rect 318 3204 319 3208
rect 323 3204 324 3208
rect 318 3203 324 3204
rect 518 3208 524 3209
rect 518 3204 519 3208
rect 523 3204 524 3208
rect 518 3203 524 3204
rect 718 3208 724 3209
rect 718 3204 719 3208
rect 723 3204 724 3208
rect 718 3203 724 3204
rect 910 3208 916 3209
rect 910 3204 911 3208
rect 915 3204 916 3208
rect 910 3203 916 3204
rect 1094 3208 1100 3209
rect 1094 3204 1095 3208
rect 1099 3204 1100 3208
rect 1094 3203 1100 3204
rect 1270 3208 1276 3209
rect 1270 3204 1271 3208
rect 1275 3204 1276 3208
rect 1270 3203 1276 3204
rect 1446 3208 1452 3209
rect 1446 3204 1447 3208
rect 1451 3204 1452 3208
rect 1446 3203 1452 3204
rect 1622 3208 1628 3209
rect 1622 3204 1623 3208
rect 1627 3204 1628 3208
rect 1622 3203 1628 3204
rect 1798 3208 1804 3209
rect 1798 3204 1799 3208
rect 1803 3204 1804 3208
rect 2006 3207 2007 3211
rect 2011 3207 2012 3211
rect 2006 3206 2012 3207
rect 1798 3203 1804 3204
rect 3374 3175 3380 3176
rect 3374 3171 3375 3175
rect 3379 3174 3380 3175
rect 3379 3172 3534 3174
rect 3379 3171 3380 3172
rect 3374 3170 3380 3171
rect 2246 3168 2252 3169
rect 2046 3165 2052 3166
rect 2046 3161 2047 3165
rect 2051 3161 2052 3165
rect 2246 3164 2247 3168
rect 2251 3164 2252 3168
rect 2246 3163 2252 3164
rect 2398 3168 2404 3169
rect 2398 3164 2399 3168
rect 2403 3164 2404 3168
rect 2398 3163 2404 3164
rect 2558 3168 2564 3169
rect 2558 3164 2559 3168
rect 2563 3164 2564 3168
rect 2558 3163 2564 3164
rect 2726 3168 2732 3169
rect 2726 3164 2727 3168
rect 2731 3164 2732 3168
rect 2726 3163 2732 3164
rect 2902 3168 2908 3169
rect 2902 3164 2903 3168
rect 2907 3164 2908 3168
rect 2902 3163 2908 3164
rect 3078 3168 3084 3169
rect 3078 3164 3079 3168
rect 3083 3164 3084 3168
rect 3078 3163 3084 3164
rect 3262 3168 3268 3169
rect 3262 3164 3263 3168
rect 3267 3164 3268 3168
rect 3262 3163 3268 3164
rect 3446 3168 3452 3169
rect 3446 3164 3447 3168
rect 3451 3164 3452 3168
rect 3446 3163 3452 3164
rect 2046 3160 2052 3161
rect 2322 3159 2328 3160
rect 2322 3155 2323 3159
rect 2327 3155 2328 3159
rect 2322 3154 2328 3155
rect 2330 3159 2336 3160
rect 2330 3155 2331 3159
rect 2335 3158 2336 3159
rect 2634 3159 2640 3160
rect 2335 3156 2441 3158
rect 2335 3155 2336 3156
rect 2330 3154 2336 3155
rect 2634 3155 2635 3159
rect 2639 3155 2640 3159
rect 2634 3154 2640 3155
rect 2802 3159 2808 3160
rect 2802 3155 2803 3159
rect 2807 3155 2808 3159
rect 2802 3154 2808 3155
rect 2839 3159 2845 3160
rect 2839 3155 2840 3159
rect 2844 3158 2845 3159
rect 3154 3159 3160 3160
rect 2844 3156 2945 3158
rect 2844 3155 2845 3156
rect 2839 3154 2845 3155
rect 3154 3155 3155 3159
rect 3159 3155 3160 3159
rect 3154 3154 3160 3155
rect 3338 3159 3344 3160
rect 3338 3155 3339 3159
rect 3343 3155 3344 3159
rect 3338 3154 3344 3155
rect 3522 3159 3528 3160
rect 3522 3155 3523 3159
rect 3527 3155 3528 3159
rect 3532 3158 3534 3172
rect 3630 3168 3636 3169
rect 3630 3164 3631 3168
rect 3635 3164 3636 3168
rect 3630 3163 3636 3164
rect 3814 3168 3820 3169
rect 3814 3164 3815 3168
rect 3819 3164 3820 3168
rect 3814 3163 3820 3164
rect 3942 3165 3948 3166
rect 3942 3161 3943 3165
rect 3947 3161 3948 3165
rect 3942 3160 3948 3161
rect 3890 3159 3896 3160
rect 3532 3156 3673 3158
rect 3522 3154 3528 3155
rect 3890 3155 3891 3159
rect 3895 3155 3896 3159
rect 3890 3154 3896 3155
rect 2246 3149 2252 3150
rect 2046 3148 2052 3149
rect 2046 3144 2047 3148
rect 2051 3144 2052 3148
rect 2246 3145 2247 3149
rect 2251 3145 2252 3149
rect 2246 3144 2252 3145
rect 2398 3149 2404 3150
rect 2398 3145 2399 3149
rect 2403 3145 2404 3149
rect 2398 3144 2404 3145
rect 2558 3149 2564 3150
rect 2558 3145 2559 3149
rect 2563 3145 2564 3149
rect 2558 3144 2564 3145
rect 2726 3149 2732 3150
rect 2726 3145 2727 3149
rect 2731 3145 2732 3149
rect 2726 3144 2732 3145
rect 2902 3149 2908 3150
rect 2902 3145 2903 3149
rect 2907 3145 2908 3149
rect 2902 3144 2908 3145
rect 3078 3149 3084 3150
rect 3078 3145 3079 3149
rect 3083 3145 3084 3149
rect 3078 3144 3084 3145
rect 3262 3149 3268 3150
rect 3262 3145 3263 3149
rect 3267 3145 3268 3149
rect 3262 3144 3268 3145
rect 3446 3149 3452 3150
rect 3446 3145 3447 3149
rect 3451 3145 3452 3149
rect 3446 3144 3452 3145
rect 3630 3149 3636 3150
rect 3630 3145 3631 3149
rect 3635 3145 3636 3149
rect 3630 3144 3636 3145
rect 3814 3149 3820 3150
rect 3814 3145 3815 3149
rect 3819 3145 3820 3149
rect 3814 3144 3820 3145
rect 3942 3148 3948 3149
rect 3942 3144 3943 3148
rect 3947 3144 3948 3148
rect 2046 3143 2052 3144
rect 3942 3143 3948 3144
rect 142 3140 148 3141
rect 110 3137 116 3138
rect 110 3133 111 3137
rect 115 3133 116 3137
rect 142 3136 143 3140
rect 147 3136 148 3140
rect 142 3135 148 3136
rect 342 3140 348 3141
rect 342 3136 343 3140
rect 347 3136 348 3140
rect 342 3135 348 3136
rect 542 3140 548 3141
rect 542 3136 543 3140
rect 547 3136 548 3140
rect 542 3135 548 3136
rect 742 3140 748 3141
rect 742 3136 743 3140
rect 747 3136 748 3140
rect 742 3135 748 3136
rect 926 3140 932 3141
rect 926 3136 927 3140
rect 931 3136 932 3140
rect 926 3135 932 3136
rect 1102 3140 1108 3141
rect 1102 3136 1103 3140
rect 1107 3136 1108 3140
rect 1102 3135 1108 3136
rect 1262 3140 1268 3141
rect 1262 3136 1263 3140
rect 1267 3136 1268 3140
rect 1262 3135 1268 3136
rect 1422 3140 1428 3141
rect 1422 3136 1423 3140
rect 1427 3136 1428 3140
rect 1422 3135 1428 3136
rect 1574 3140 1580 3141
rect 1574 3136 1575 3140
rect 1579 3136 1580 3140
rect 1574 3135 1580 3136
rect 1734 3140 1740 3141
rect 1734 3136 1735 3140
rect 1739 3136 1740 3140
rect 1734 3135 1740 3136
rect 2006 3137 2012 3138
rect 110 3132 116 3133
rect 2006 3133 2007 3137
rect 2011 3133 2012 3137
rect 2839 3135 2845 3136
rect 2839 3134 2840 3135
rect 2006 3132 2012 3133
rect 2616 3132 2840 3134
rect 218 3131 224 3132
rect 218 3127 219 3131
rect 223 3127 224 3131
rect 218 3126 224 3127
rect 418 3131 424 3132
rect 418 3127 419 3131
rect 423 3127 424 3131
rect 630 3131 636 3132
rect 630 3130 631 3131
rect 621 3128 631 3130
rect 418 3126 424 3127
rect 630 3127 631 3128
rect 635 3127 636 3131
rect 630 3126 636 3127
rect 678 3131 684 3132
rect 678 3127 679 3131
rect 683 3130 684 3131
rect 826 3131 832 3132
rect 683 3128 785 3130
rect 683 3127 684 3128
rect 678 3126 684 3127
rect 826 3127 827 3131
rect 831 3130 832 3131
rect 1178 3131 1184 3132
rect 831 3128 969 3130
rect 831 3127 832 3128
rect 826 3126 832 3127
rect 1178 3127 1179 3131
rect 1183 3127 1184 3131
rect 1178 3126 1184 3127
rect 1186 3131 1192 3132
rect 1186 3127 1187 3131
rect 1191 3130 1192 3131
rect 1346 3131 1352 3132
rect 1191 3128 1305 3130
rect 1191 3127 1192 3128
rect 1186 3126 1192 3127
rect 1346 3127 1347 3131
rect 1351 3130 1352 3131
rect 1650 3131 1656 3132
rect 1351 3128 1465 3130
rect 1351 3127 1352 3128
rect 1346 3126 1352 3127
rect 1650 3127 1651 3131
rect 1655 3127 1656 3131
rect 1650 3126 1656 3127
rect 1658 3131 1664 3132
rect 1658 3127 1659 3131
rect 1663 3130 1664 3131
rect 1663 3128 1777 3130
rect 1663 3127 1664 3128
rect 1658 3126 1664 3127
rect 2311 3127 2317 3128
rect 2311 3123 2312 3127
rect 2316 3126 2317 3127
rect 2330 3127 2336 3128
rect 2330 3126 2331 3127
rect 2316 3124 2331 3126
rect 2316 3123 2317 3124
rect 2311 3122 2317 3123
rect 2330 3123 2331 3124
rect 2335 3123 2336 3127
rect 2330 3122 2336 3123
rect 2463 3127 2469 3128
rect 2463 3123 2464 3127
rect 2468 3126 2469 3127
rect 2616 3126 2618 3132
rect 2839 3131 2840 3132
rect 2844 3131 2845 3135
rect 2839 3130 2845 3131
rect 2468 3124 2618 3126
rect 2623 3127 2632 3128
rect 2468 3123 2469 3124
rect 2463 3122 2469 3123
rect 2623 3123 2624 3127
rect 2631 3123 2632 3127
rect 2623 3122 2632 3123
rect 2634 3127 2640 3128
rect 2634 3123 2635 3127
rect 2639 3126 2640 3127
rect 2791 3127 2797 3128
rect 2791 3126 2792 3127
rect 2639 3124 2792 3126
rect 2639 3123 2640 3124
rect 2634 3122 2640 3123
rect 2791 3123 2792 3124
rect 2796 3123 2797 3127
rect 2791 3122 2797 3123
rect 2802 3127 2808 3128
rect 2802 3123 2803 3127
rect 2807 3126 2808 3127
rect 2967 3127 2973 3128
rect 2967 3126 2968 3127
rect 2807 3124 2968 3126
rect 2807 3123 2808 3124
rect 2802 3122 2808 3123
rect 2967 3123 2968 3124
rect 2972 3123 2973 3127
rect 2967 3122 2973 3123
rect 3143 3127 3149 3128
rect 3143 3123 3144 3127
rect 3148 3126 3149 3127
rect 3154 3127 3160 3128
rect 3148 3123 3150 3126
rect 3143 3122 3150 3123
rect 3154 3123 3155 3127
rect 3159 3126 3160 3127
rect 3327 3127 3333 3128
rect 3327 3126 3328 3127
rect 3159 3124 3328 3126
rect 3159 3123 3160 3124
rect 3154 3122 3160 3123
rect 3327 3123 3328 3124
rect 3332 3123 3333 3127
rect 3327 3122 3333 3123
rect 3338 3127 3344 3128
rect 3338 3123 3339 3127
rect 3343 3126 3344 3127
rect 3511 3127 3517 3128
rect 3511 3126 3512 3127
rect 3343 3124 3512 3126
rect 3343 3123 3344 3124
rect 3338 3122 3344 3123
rect 3511 3123 3512 3124
rect 3516 3123 3517 3127
rect 3511 3122 3517 3123
rect 3522 3127 3528 3128
rect 3522 3123 3523 3127
rect 3527 3126 3528 3127
rect 3695 3127 3701 3128
rect 3695 3126 3696 3127
rect 3527 3124 3696 3126
rect 3527 3123 3528 3124
rect 3522 3122 3528 3123
rect 3695 3123 3696 3124
rect 3700 3123 3701 3127
rect 3695 3122 3701 3123
rect 3879 3127 3885 3128
rect 3879 3123 3880 3127
rect 3884 3126 3885 3127
rect 3914 3127 3920 3128
rect 3914 3126 3915 3127
rect 3884 3124 3915 3126
rect 3884 3123 3885 3124
rect 3879 3122 3885 3123
rect 3914 3123 3915 3124
rect 3919 3123 3920 3127
rect 3914 3122 3920 3123
rect 142 3121 148 3122
rect 110 3120 116 3121
rect 110 3116 111 3120
rect 115 3116 116 3120
rect 142 3117 143 3121
rect 147 3117 148 3121
rect 142 3116 148 3117
rect 342 3121 348 3122
rect 342 3117 343 3121
rect 347 3117 348 3121
rect 342 3116 348 3117
rect 542 3121 548 3122
rect 542 3117 543 3121
rect 547 3117 548 3121
rect 542 3116 548 3117
rect 742 3121 748 3122
rect 742 3117 743 3121
rect 747 3117 748 3121
rect 742 3116 748 3117
rect 926 3121 932 3122
rect 926 3117 927 3121
rect 931 3117 932 3121
rect 926 3116 932 3117
rect 1102 3121 1108 3122
rect 1102 3117 1103 3121
rect 1107 3117 1108 3121
rect 1102 3116 1108 3117
rect 1262 3121 1268 3122
rect 1262 3117 1263 3121
rect 1267 3117 1268 3121
rect 1262 3116 1268 3117
rect 1422 3121 1428 3122
rect 1422 3117 1423 3121
rect 1427 3117 1428 3121
rect 1422 3116 1428 3117
rect 1574 3121 1580 3122
rect 1574 3117 1575 3121
rect 1579 3117 1580 3121
rect 1574 3116 1580 3117
rect 1734 3121 1740 3122
rect 1734 3117 1735 3121
rect 1739 3117 1740 3121
rect 1734 3116 1740 3117
rect 2006 3120 2012 3121
rect 2006 3116 2007 3120
rect 2011 3116 2012 3120
rect 3148 3118 3150 3122
rect 3602 3119 3608 3120
rect 3602 3118 3603 3119
rect 3148 3116 3603 3118
rect 110 3115 116 3116
rect 2006 3115 2012 3116
rect 3602 3115 3603 3116
rect 3607 3115 3608 3119
rect 3602 3114 3608 3115
rect 2143 3111 2149 3112
rect 2143 3107 2144 3111
rect 2148 3110 2149 3111
rect 2154 3111 2160 3112
rect 2148 3107 2150 3110
rect 2143 3106 2150 3107
rect 2154 3107 2155 3111
rect 2159 3110 2160 3111
rect 2287 3111 2293 3112
rect 2287 3110 2288 3111
rect 2159 3108 2288 3110
rect 2159 3107 2160 3108
rect 2154 3106 2160 3107
rect 2287 3107 2288 3108
rect 2292 3107 2293 3111
rect 2287 3106 2293 3107
rect 2322 3111 2328 3112
rect 2322 3107 2323 3111
rect 2327 3110 2328 3111
rect 2439 3111 2445 3112
rect 2439 3110 2440 3111
rect 2327 3108 2440 3110
rect 2327 3107 2328 3108
rect 2322 3106 2328 3107
rect 2439 3107 2440 3108
rect 2444 3107 2445 3111
rect 2439 3106 2445 3107
rect 2450 3111 2456 3112
rect 2450 3107 2451 3111
rect 2455 3110 2456 3111
rect 2591 3111 2597 3112
rect 2591 3110 2592 3111
rect 2455 3108 2592 3110
rect 2455 3107 2456 3108
rect 2450 3106 2456 3107
rect 2591 3107 2592 3108
rect 2596 3107 2597 3111
rect 2591 3106 2597 3107
rect 2602 3111 2608 3112
rect 2602 3107 2603 3111
rect 2607 3110 2608 3111
rect 2751 3111 2757 3112
rect 2751 3110 2752 3111
rect 2607 3108 2752 3110
rect 2607 3107 2608 3108
rect 2602 3106 2608 3107
rect 2751 3107 2752 3108
rect 2756 3107 2757 3111
rect 2751 3106 2757 3107
rect 2919 3111 2928 3112
rect 2919 3107 2920 3111
rect 2927 3107 2928 3111
rect 2919 3106 2928 3107
rect 2930 3111 2936 3112
rect 2930 3107 2931 3111
rect 2935 3110 2936 3111
rect 3103 3111 3109 3112
rect 3103 3110 3104 3111
rect 2935 3108 3104 3110
rect 2935 3107 2936 3108
rect 2930 3106 2936 3107
rect 3103 3107 3104 3108
rect 3108 3107 3109 3111
rect 3103 3106 3109 3107
rect 3114 3111 3120 3112
rect 3114 3107 3115 3111
rect 3119 3110 3120 3111
rect 3295 3111 3301 3112
rect 3295 3110 3296 3111
rect 3119 3108 3296 3110
rect 3119 3107 3120 3108
rect 3114 3106 3120 3107
rect 3295 3107 3296 3108
rect 3300 3107 3301 3111
rect 3295 3106 3301 3107
rect 3306 3111 3312 3112
rect 3306 3107 3307 3111
rect 3311 3110 3312 3111
rect 3495 3111 3501 3112
rect 3495 3110 3496 3111
rect 3311 3108 3496 3110
rect 3311 3107 3312 3108
rect 3306 3106 3312 3107
rect 3495 3107 3496 3108
rect 3500 3107 3501 3111
rect 3495 3106 3501 3107
rect 3506 3111 3512 3112
rect 3506 3107 3507 3111
rect 3511 3110 3512 3111
rect 3703 3111 3709 3112
rect 3703 3110 3704 3111
rect 3511 3108 3704 3110
rect 3511 3107 3512 3108
rect 3506 3106 3512 3107
rect 3703 3107 3704 3108
rect 3708 3107 3709 3111
rect 3703 3106 3709 3107
rect 3890 3111 3896 3112
rect 3890 3107 3891 3111
rect 3895 3110 3896 3111
rect 3903 3111 3909 3112
rect 3903 3110 3904 3111
rect 3895 3108 3904 3110
rect 3895 3107 3896 3108
rect 3890 3106 3896 3107
rect 3903 3107 3904 3108
rect 3908 3107 3909 3111
rect 3903 3106 3909 3107
rect 2148 3102 2150 3106
rect 2658 3103 2664 3104
rect 2658 3102 2659 3103
rect 2148 3100 2659 3102
rect 207 3099 216 3100
rect 207 3095 208 3099
rect 215 3095 216 3099
rect 207 3094 216 3095
rect 218 3099 224 3100
rect 218 3095 219 3099
rect 223 3098 224 3099
rect 407 3099 413 3100
rect 407 3098 408 3099
rect 223 3096 408 3098
rect 223 3095 224 3096
rect 218 3094 224 3095
rect 407 3095 408 3096
rect 412 3095 413 3099
rect 407 3094 413 3095
rect 418 3099 424 3100
rect 418 3095 419 3099
rect 423 3098 424 3099
rect 607 3099 613 3100
rect 607 3098 608 3099
rect 423 3096 608 3098
rect 423 3095 424 3096
rect 418 3094 424 3095
rect 607 3095 608 3096
rect 612 3095 613 3099
rect 607 3094 613 3095
rect 807 3099 813 3100
rect 807 3095 808 3099
rect 812 3098 813 3099
rect 826 3099 832 3100
rect 826 3098 827 3099
rect 812 3096 827 3098
rect 812 3095 813 3096
rect 807 3094 813 3095
rect 826 3095 827 3096
rect 831 3095 832 3099
rect 826 3094 832 3095
rect 991 3099 997 3100
rect 991 3095 992 3099
rect 996 3098 997 3099
rect 1050 3099 1056 3100
rect 1050 3098 1051 3099
rect 996 3096 1051 3098
rect 996 3095 997 3096
rect 991 3094 997 3095
rect 1050 3095 1051 3096
rect 1055 3095 1056 3099
rect 1050 3094 1056 3095
rect 1167 3099 1173 3100
rect 1167 3095 1168 3099
rect 1172 3098 1173 3099
rect 1186 3099 1192 3100
rect 1186 3098 1187 3099
rect 1172 3096 1187 3098
rect 1172 3095 1173 3096
rect 1167 3094 1173 3095
rect 1186 3095 1187 3096
rect 1191 3095 1192 3099
rect 1186 3094 1192 3095
rect 1327 3099 1333 3100
rect 1327 3095 1328 3099
rect 1332 3098 1333 3099
rect 1346 3099 1352 3100
rect 1346 3098 1347 3099
rect 1332 3096 1347 3098
rect 1332 3095 1333 3096
rect 1327 3094 1333 3095
rect 1346 3095 1347 3096
rect 1351 3095 1352 3099
rect 1346 3094 1352 3095
rect 1487 3099 1493 3100
rect 1487 3095 1488 3099
rect 1492 3098 1493 3099
rect 1522 3099 1528 3100
rect 1522 3098 1523 3099
rect 1492 3096 1523 3098
rect 1492 3095 1493 3096
rect 1487 3094 1493 3095
rect 1522 3095 1523 3096
rect 1527 3095 1528 3099
rect 1522 3094 1528 3095
rect 1639 3099 1645 3100
rect 1639 3095 1640 3099
rect 1644 3098 1645 3099
rect 1658 3099 1664 3100
rect 1658 3098 1659 3099
rect 1644 3096 1659 3098
rect 1644 3095 1645 3096
rect 1639 3094 1645 3095
rect 1658 3095 1659 3096
rect 1663 3095 1664 3099
rect 1658 3094 1664 3095
rect 1799 3099 1805 3100
rect 1799 3095 1800 3099
rect 1804 3098 1805 3099
rect 1842 3099 1848 3100
rect 1842 3098 1843 3099
rect 1804 3096 1843 3098
rect 1804 3095 1805 3096
rect 1799 3094 1805 3095
rect 1842 3095 1843 3096
rect 1847 3095 1848 3099
rect 2658 3099 2659 3100
rect 2663 3099 2664 3103
rect 2658 3098 2664 3099
rect 1842 3094 1848 3095
rect 2046 3092 2052 3093
rect 3942 3092 3948 3093
rect 2046 3088 2047 3092
rect 2051 3088 2052 3092
rect 327 3087 333 3088
rect 327 3083 328 3087
rect 332 3086 333 3087
rect 386 3087 392 3088
rect 332 3084 382 3086
rect 332 3083 333 3084
rect 327 3082 333 3083
rect 380 3078 382 3084
rect 386 3083 387 3087
rect 391 3086 392 3087
rect 503 3087 509 3088
rect 503 3086 504 3087
rect 391 3084 504 3086
rect 391 3083 392 3084
rect 386 3082 392 3083
rect 503 3083 504 3084
rect 508 3083 509 3087
rect 503 3082 509 3083
rect 630 3087 636 3088
rect 630 3083 631 3087
rect 635 3086 636 3087
rect 679 3087 685 3088
rect 679 3086 680 3087
rect 635 3084 680 3086
rect 635 3083 636 3084
rect 630 3082 636 3083
rect 679 3083 680 3084
rect 684 3083 685 3087
rect 679 3082 685 3083
rect 858 3087 869 3088
rect 858 3083 859 3087
rect 863 3083 864 3087
rect 868 3083 869 3087
rect 858 3082 869 3083
rect 874 3087 880 3088
rect 874 3083 875 3087
rect 879 3086 880 3087
rect 1039 3087 1045 3088
rect 1039 3086 1040 3087
rect 879 3084 1040 3086
rect 879 3083 880 3084
rect 874 3082 880 3083
rect 1039 3083 1040 3084
rect 1044 3083 1045 3087
rect 1039 3082 1045 3083
rect 1178 3087 1184 3088
rect 1178 3083 1179 3087
rect 1183 3086 1184 3087
rect 1207 3087 1213 3088
rect 1207 3086 1208 3087
rect 1183 3084 1208 3086
rect 1183 3083 1184 3084
rect 1178 3082 1184 3083
rect 1207 3083 1208 3084
rect 1212 3083 1213 3087
rect 1207 3082 1213 3083
rect 1218 3087 1224 3088
rect 1218 3083 1219 3087
rect 1223 3086 1224 3087
rect 1367 3087 1373 3088
rect 1367 3086 1368 3087
rect 1223 3084 1368 3086
rect 1223 3083 1224 3084
rect 1218 3082 1224 3083
rect 1367 3083 1368 3084
rect 1372 3083 1373 3087
rect 1367 3082 1373 3083
rect 1378 3087 1384 3088
rect 1378 3083 1379 3087
rect 1383 3086 1384 3087
rect 1519 3087 1525 3088
rect 1519 3086 1520 3087
rect 1383 3084 1520 3086
rect 1383 3083 1384 3084
rect 1378 3082 1384 3083
rect 1519 3083 1520 3084
rect 1524 3083 1525 3087
rect 1519 3082 1525 3083
rect 1530 3087 1536 3088
rect 1530 3083 1531 3087
rect 1535 3086 1536 3087
rect 1671 3087 1677 3088
rect 1671 3086 1672 3087
rect 1535 3084 1672 3086
rect 1535 3083 1536 3084
rect 1530 3082 1536 3083
rect 1671 3083 1672 3084
rect 1676 3083 1677 3087
rect 1671 3082 1677 3083
rect 1682 3087 1688 3088
rect 1682 3083 1683 3087
rect 1687 3086 1688 3087
rect 1831 3087 1837 3088
rect 2046 3087 2052 3088
rect 2078 3091 2084 3092
rect 2078 3087 2079 3091
rect 2083 3087 2084 3091
rect 1831 3086 1832 3087
rect 1687 3084 1832 3086
rect 1687 3083 1688 3084
rect 1682 3082 1688 3083
rect 1831 3083 1832 3084
rect 1836 3083 1837 3087
rect 2078 3086 2084 3087
rect 2222 3091 2228 3092
rect 2222 3087 2223 3091
rect 2227 3087 2228 3091
rect 2222 3086 2228 3087
rect 2374 3091 2380 3092
rect 2374 3087 2375 3091
rect 2379 3087 2380 3091
rect 2374 3086 2380 3087
rect 2526 3091 2532 3092
rect 2526 3087 2527 3091
rect 2531 3087 2532 3091
rect 2526 3086 2532 3087
rect 2686 3091 2692 3092
rect 2686 3087 2687 3091
rect 2691 3087 2692 3091
rect 2686 3086 2692 3087
rect 2854 3091 2860 3092
rect 2854 3087 2855 3091
rect 2859 3087 2860 3091
rect 2854 3086 2860 3087
rect 3038 3091 3044 3092
rect 3038 3087 3039 3091
rect 3043 3087 3044 3091
rect 3038 3086 3044 3087
rect 3230 3091 3236 3092
rect 3230 3087 3231 3091
rect 3235 3087 3236 3091
rect 3230 3086 3236 3087
rect 3430 3091 3436 3092
rect 3430 3087 3431 3091
rect 3435 3087 3436 3091
rect 3430 3086 3436 3087
rect 3638 3091 3644 3092
rect 3638 3087 3639 3091
rect 3643 3087 3644 3091
rect 3638 3086 3644 3087
rect 3838 3091 3844 3092
rect 3838 3087 3839 3091
rect 3843 3087 3844 3091
rect 3942 3088 3943 3092
rect 3947 3088 3948 3092
rect 3942 3087 3948 3088
rect 3838 3086 3844 3087
rect 1831 3082 1837 3083
rect 2154 3083 2160 3084
rect 558 3079 564 3080
rect 558 3078 559 3079
rect 380 3076 559 3078
rect 558 3075 559 3076
rect 563 3075 564 3079
rect 2154 3079 2155 3083
rect 2159 3079 2160 3083
rect 2450 3083 2456 3084
rect 2154 3078 2160 3079
rect 2298 3079 2304 3080
rect 558 3074 564 3075
rect 2046 3075 2052 3076
rect 2046 3071 2047 3075
rect 2051 3071 2052 3075
rect 2298 3075 2299 3079
rect 2303 3075 2304 3079
rect 2450 3079 2451 3083
rect 2455 3079 2456 3083
rect 2450 3078 2456 3079
rect 2602 3083 2608 3084
rect 2602 3079 2603 3083
rect 2607 3079 2608 3083
rect 2602 3078 2608 3079
rect 2658 3083 2664 3084
rect 2658 3079 2659 3083
rect 2663 3082 2664 3083
rect 2930 3083 2936 3084
rect 2663 3080 2729 3082
rect 2663 3079 2664 3080
rect 2658 3078 2664 3079
rect 2930 3079 2931 3083
rect 2935 3079 2936 3083
rect 2930 3078 2936 3079
rect 3114 3083 3120 3084
rect 3114 3079 3115 3083
rect 3119 3079 3120 3083
rect 3114 3078 3120 3079
rect 3306 3083 3312 3084
rect 3306 3079 3307 3083
rect 3311 3079 3312 3083
rect 3306 3078 3312 3079
rect 3506 3083 3512 3084
rect 3506 3079 3507 3083
rect 3511 3079 3512 3083
rect 3506 3078 3512 3079
rect 3602 3083 3608 3084
rect 3602 3079 3603 3083
rect 3607 3082 3608 3083
rect 3607 3080 3681 3082
rect 3607 3079 3608 3080
rect 3602 3078 3608 3079
rect 3914 3079 3920 3080
rect 2298 3074 2304 3075
rect 3914 3075 3915 3079
rect 3919 3075 3920 3079
rect 3914 3074 3920 3075
rect 3942 3075 3948 3076
rect 2046 3070 2052 3071
rect 2078 3072 2084 3073
rect 110 3068 116 3069
rect 2006 3068 2012 3069
rect 110 3064 111 3068
rect 115 3064 116 3068
rect 110 3063 116 3064
rect 262 3067 268 3068
rect 262 3063 263 3067
rect 267 3063 268 3067
rect 262 3062 268 3063
rect 438 3067 444 3068
rect 438 3063 439 3067
rect 443 3063 444 3067
rect 438 3062 444 3063
rect 614 3067 620 3068
rect 614 3063 615 3067
rect 619 3063 620 3067
rect 614 3062 620 3063
rect 798 3067 804 3068
rect 798 3063 799 3067
rect 803 3063 804 3067
rect 798 3062 804 3063
rect 974 3067 980 3068
rect 974 3063 975 3067
rect 979 3063 980 3067
rect 974 3062 980 3063
rect 1142 3067 1148 3068
rect 1142 3063 1143 3067
rect 1147 3063 1148 3067
rect 1142 3062 1148 3063
rect 1302 3067 1308 3068
rect 1302 3063 1303 3067
rect 1307 3063 1308 3067
rect 1302 3062 1308 3063
rect 1454 3067 1460 3068
rect 1454 3063 1455 3067
rect 1459 3063 1460 3067
rect 1454 3062 1460 3063
rect 1606 3067 1612 3068
rect 1606 3063 1607 3067
rect 1611 3063 1612 3067
rect 1606 3062 1612 3063
rect 1766 3067 1772 3068
rect 1766 3063 1767 3067
rect 1771 3063 1772 3067
rect 2006 3064 2007 3068
rect 2011 3064 2012 3068
rect 2078 3068 2079 3072
rect 2083 3068 2084 3072
rect 2078 3067 2084 3068
rect 2222 3072 2228 3073
rect 2222 3068 2223 3072
rect 2227 3068 2228 3072
rect 2222 3067 2228 3068
rect 2374 3072 2380 3073
rect 2374 3068 2375 3072
rect 2379 3068 2380 3072
rect 2374 3067 2380 3068
rect 2526 3072 2532 3073
rect 2526 3068 2527 3072
rect 2531 3068 2532 3072
rect 2526 3067 2532 3068
rect 2686 3072 2692 3073
rect 2686 3068 2687 3072
rect 2691 3068 2692 3072
rect 2686 3067 2692 3068
rect 2854 3072 2860 3073
rect 2854 3068 2855 3072
rect 2859 3068 2860 3072
rect 2854 3067 2860 3068
rect 3038 3072 3044 3073
rect 3038 3068 3039 3072
rect 3043 3068 3044 3072
rect 3038 3067 3044 3068
rect 3230 3072 3236 3073
rect 3230 3068 3231 3072
rect 3235 3068 3236 3072
rect 3230 3067 3236 3068
rect 3430 3072 3436 3073
rect 3430 3068 3431 3072
rect 3435 3068 3436 3072
rect 3430 3067 3436 3068
rect 3638 3072 3644 3073
rect 3638 3068 3639 3072
rect 3643 3068 3644 3072
rect 3638 3067 3644 3068
rect 3838 3072 3844 3073
rect 3838 3068 3839 3072
rect 3843 3068 3844 3072
rect 3942 3071 3943 3075
rect 3947 3071 3948 3075
rect 3942 3070 3948 3071
rect 3838 3067 3844 3068
rect 2006 3063 2012 3064
rect 1766 3062 1772 3063
rect 386 3059 392 3060
rect 386 3058 387 3059
rect 341 3056 387 3058
rect 386 3055 387 3056
rect 391 3055 392 3059
rect 558 3059 564 3060
rect 386 3054 392 3055
rect 514 3055 520 3056
rect 110 3051 116 3052
rect 110 3047 111 3051
rect 115 3047 116 3051
rect 514 3051 515 3055
rect 519 3051 520 3055
rect 558 3055 559 3059
rect 563 3058 564 3059
rect 874 3059 880 3060
rect 563 3056 657 3058
rect 563 3055 564 3056
rect 558 3054 564 3055
rect 874 3055 875 3059
rect 879 3055 880 3059
rect 874 3054 880 3055
rect 1050 3059 1056 3060
rect 1050 3055 1051 3059
rect 1055 3055 1056 3059
rect 1050 3054 1056 3055
rect 1218 3059 1224 3060
rect 1218 3055 1219 3059
rect 1223 3055 1224 3059
rect 1218 3054 1224 3055
rect 1378 3059 1384 3060
rect 1378 3055 1379 3059
rect 1383 3055 1384 3059
rect 1378 3054 1384 3055
rect 1530 3059 1536 3060
rect 1530 3055 1531 3059
rect 1535 3055 1536 3059
rect 1530 3054 1536 3055
rect 1682 3059 1688 3060
rect 1682 3055 1683 3059
rect 1687 3055 1688 3059
rect 1682 3054 1688 3055
rect 1842 3059 1848 3060
rect 1842 3055 1843 3059
rect 1847 3055 1848 3059
rect 1842 3054 1848 3055
rect 514 3050 520 3051
rect 2006 3051 2012 3052
rect 110 3046 116 3047
rect 262 3048 268 3049
rect 262 3044 263 3048
rect 267 3044 268 3048
rect 262 3043 268 3044
rect 438 3048 444 3049
rect 438 3044 439 3048
rect 443 3044 444 3048
rect 438 3043 444 3044
rect 614 3048 620 3049
rect 614 3044 615 3048
rect 619 3044 620 3048
rect 614 3043 620 3044
rect 798 3048 804 3049
rect 798 3044 799 3048
rect 803 3044 804 3048
rect 798 3043 804 3044
rect 974 3048 980 3049
rect 974 3044 975 3048
rect 979 3044 980 3048
rect 974 3043 980 3044
rect 1142 3048 1148 3049
rect 1142 3044 1143 3048
rect 1147 3044 1148 3048
rect 1142 3043 1148 3044
rect 1302 3048 1308 3049
rect 1302 3044 1303 3048
rect 1307 3044 1308 3048
rect 1302 3043 1308 3044
rect 1454 3048 1460 3049
rect 1454 3044 1455 3048
rect 1459 3044 1460 3048
rect 1454 3043 1460 3044
rect 1606 3048 1612 3049
rect 1606 3044 1607 3048
rect 1611 3044 1612 3048
rect 1606 3043 1612 3044
rect 1766 3048 1772 3049
rect 1766 3044 1767 3048
rect 1771 3044 1772 3048
rect 2006 3047 2007 3051
rect 2011 3047 2012 3051
rect 2006 3046 2012 3047
rect 1766 3043 1772 3044
rect 2922 3011 2928 3012
rect 2922 3007 2923 3011
rect 2927 3010 2928 3011
rect 2927 3008 3422 3010
rect 2927 3007 2928 3008
rect 2922 3006 2928 3007
rect 2070 3004 2076 3005
rect 2046 3001 2052 3002
rect 2046 2997 2047 3001
rect 2051 2997 2052 3001
rect 2070 3000 2071 3004
rect 2075 3000 2076 3004
rect 2070 2999 2076 3000
rect 2182 3004 2188 3005
rect 2182 3000 2183 3004
rect 2187 3000 2188 3004
rect 2182 2999 2188 3000
rect 2326 3004 2332 3005
rect 2326 3000 2327 3004
rect 2331 3000 2332 3004
rect 2326 2999 2332 3000
rect 2478 3004 2484 3005
rect 2478 3000 2479 3004
rect 2483 3000 2484 3004
rect 2478 2999 2484 3000
rect 2654 3004 2660 3005
rect 2654 3000 2655 3004
rect 2659 3000 2660 3004
rect 2654 2999 2660 3000
rect 2854 3004 2860 3005
rect 2854 3000 2855 3004
rect 2859 3000 2860 3004
rect 2854 2999 2860 3000
rect 3086 3004 3092 3005
rect 3086 3000 3087 3004
rect 3091 3000 3092 3004
rect 3086 2999 3092 3000
rect 3334 3004 3340 3005
rect 3334 3000 3335 3004
rect 3339 3000 3340 3004
rect 3334 2999 3340 3000
rect 2046 2996 2052 2997
rect 2138 2995 2144 2996
rect 2138 2991 2139 2995
rect 2143 2991 2144 2995
rect 2138 2990 2144 2991
rect 2154 2995 2160 2996
rect 2154 2991 2155 2995
rect 2159 2994 2160 2995
rect 2402 2995 2408 2996
rect 2159 2992 2225 2994
rect 2159 2991 2160 2992
rect 2154 2990 2160 2991
rect 2402 2991 2403 2995
rect 2407 2991 2408 2995
rect 2402 2990 2408 2991
rect 2554 2995 2560 2996
rect 2554 2991 2555 2995
rect 2559 2991 2560 2995
rect 2554 2990 2560 2991
rect 2598 2995 2604 2996
rect 2598 2991 2599 2995
rect 2603 2994 2604 2995
rect 2930 2995 2936 2996
rect 2603 2992 2697 2994
rect 2603 2991 2604 2992
rect 2598 2990 2604 2991
rect 2930 2991 2931 2995
rect 2935 2991 2936 2995
rect 2930 2990 2936 2991
rect 3162 2995 3168 2996
rect 3162 2991 3163 2995
rect 3167 2991 3168 2995
rect 3162 2990 3168 2991
rect 3410 2995 3416 2996
rect 3410 2991 3411 2995
rect 3415 2991 3416 2995
rect 3420 2994 3422 3008
rect 3598 3004 3604 3005
rect 3598 3000 3599 3004
rect 3603 3000 3604 3004
rect 3598 2999 3604 3000
rect 3838 3004 3844 3005
rect 3838 3000 3839 3004
rect 3843 3000 3844 3004
rect 3838 2999 3844 3000
rect 3942 3001 3948 3002
rect 3942 2997 3943 3001
rect 3947 2997 3948 3001
rect 3942 2996 3948 2997
rect 3906 2995 3912 2996
rect 3420 2992 3641 2994
rect 3410 2990 3416 2991
rect 3906 2991 3907 2995
rect 3911 2991 3912 2995
rect 3906 2990 3912 2991
rect 2070 2985 2076 2986
rect 2046 2984 2052 2985
rect 2046 2980 2047 2984
rect 2051 2980 2052 2984
rect 2070 2981 2071 2985
rect 2075 2981 2076 2985
rect 2070 2980 2076 2981
rect 2182 2985 2188 2986
rect 2182 2981 2183 2985
rect 2187 2981 2188 2985
rect 2182 2980 2188 2981
rect 2326 2985 2332 2986
rect 2326 2981 2327 2985
rect 2331 2981 2332 2985
rect 2326 2980 2332 2981
rect 2478 2985 2484 2986
rect 2478 2981 2479 2985
rect 2483 2981 2484 2985
rect 2478 2980 2484 2981
rect 2654 2985 2660 2986
rect 2654 2981 2655 2985
rect 2659 2981 2660 2985
rect 2654 2980 2660 2981
rect 2854 2985 2860 2986
rect 2854 2981 2855 2985
rect 2859 2981 2860 2985
rect 2854 2980 2860 2981
rect 3086 2985 3092 2986
rect 3086 2981 3087 2985
rect 3091 2981 3092 2985
rect 3086 2980 3092 2981
rect 3334 2985 3340 2986
rect 3334 2981 3335 2985
rect 3339 2981 3340 2985
rect 3334 2980 3340 2981
rect 3598 2985 3604 2986
rect 3598 2981 3599 2985
rect 3603 2981 3604 2985
rect 3598 2980 3604 2981
rect 3838 2985 3844 2986
rect 3838 2981 3839 2985
rect 3843 2981 3844 2985
rect 3838 2980 3844 2981
rect 3942 2984 3948 2985
rect 3942 2980 3943 2984
rect 3947 2980 3948 2984
rect 2046 2979 2052 2980
rect 3942 2979 3948 2980
rect 2598 2971 2604 2972
rect 2598 2970 2599 2971
rect 2292 2968 2599 2970
rect 342 2964 348 2965
rect 110 2961 116 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 342 2960 343 2964
rect 347 2960 348 2964
rect 342 2959 348 2960
rect 438 2964 444 2965
rect 438 2960 439 2964
rect 443 2960 444 2964
rect 438 2959 444 2960
rect 542 2964 548 2965
rect 542 2960 543 2964
rect 547 2960 548 2964
rect 542 2959 548 2960
rect 654 2964 660 2965
rect 654 2960 655 2964
rect 659 2960 660 2964
rect 654 2959 660 2960
rect 782 2964 788 2965
rect 782 2960 783 2964
rect 787 2960 788 2964
rect 782 2959 788 2960
rect 934 2964 940 2965
rect 934 2960 935 2964
rect 939 2960 940 2964
rect 934 2959 940 2960
rect 1102 2964 1108 2965
rect 1102 2960 1103 2964
rect 1107 2960 1108 2964
rect 1102 2959 1108 2960
rect 1294 2964 1300 2965
rect 1294 2960 1295 2964
rect 1299 2960 1300 2964
rect 1294 2959 1300 2960
rect 1494 2964 1500 2965
rect 1494 2960 1495 2964
rect 1499 2960 1500 2964
rect 1494 2959 1500 2960
rect 1710 2964 1716 2965
rect 1710 2960 1711 2964
rect 1715 2960 1716 2964
rect 1710 2959 1716 2960
rect 1902 2964 1908 2965
rect 1902 2960 1903 2964
rect 1907 2960 1908 2964
rect 2135 2963 2141 2964
rect 1902 2959 1908 2960
rect 2006 2961 2012 2962
rect 110 2956 116 2957
rect 2006 2957 2007 2961
rect 2011 2957 2012 2961
rect 2135 2959 2136 2963
rect 2140 2962 2141 2963
rect 2154 2963 2160 2964
rect 2154 2962 2155 2963
rect 2140 2960 2155 2962
rect 2140 2959 2141 2960
rect 2135 2958 2141 2959
rect 2154 2959 2155 2960
rect 2159 2959 2160 2963
rect 2154 2958 2160 2959
rect 2247 2963 2253 2964
rect 2247 2959 2248 2963
rect 2252 2962 2253 2963
rect 2292 2962 2294 2968
rect 2598 2967 2599 2968
rect 2603 2967 2604 2971
rect 2598 2966 2604 2967
rect 2252 2960 2294 2962
rect 2298 2963 2304 2964
rect 2252 2959 2253 2960
rect 2247 2958 2253 2959
rect 2298 2959 2299 2963
rect 2303 2962 2304 2963
rect 2391 2963 2397 2964
rect 2391 2962 2392 2963
rect 2303 2960 2392 2962
rect 2303 2959 2304 2960
rect 2298 2958 2304 2959
rect 2391 2959 2392 2960
rect 2396 2959 2397 2963
rect 2391 2958 2397 2959
rect 2402 2963 2408 2964
rect 2402 2959 2403 2963
rect 2407 2962 2408 2963
rect 2543 2963 2549 2964
rect 2543 2962 2544 2963
rect 2407 2960 2544 2962
rect 2407 2959 2408 2960
rect 2402 2958 2408 2959
rect 2543 2959 2544 2960
rect 2548 2959 2549 2963
rect 2543 2958 2549 2959
rect 2554 2963 2560 2964
rect 2554 2959 2555 2963
rect 2559 2962 2560 2963
rect 2719 2963 2725 2964
rect 2719 2962 2720 2963
rect 2559 2960 2720 2962
rect 2559 2959 2560 2960
rect 2554 2958 2560 2959
rect 2719 2959 2720 2960
rect 2724 2959 2725 2963
rect 2719 2958 2725 2959
rect 2919 2963 2925 2964
rect 2919 2959 2920 2963
rect 2924 2962 2925 2963
rect 2930 2963 2936 2964
rect 2924 2959 2926 2962
rect 2919 2958 2926 2959
rect 2930 2959 2931 2963
rect 2935 2962 2936 2963
rect 3151 2963 3157 2964
rect 3151 2962 3152 2963
rect 2935 2960 3152 2962
rect 2935 2959 2936 2960
rect 2930 2958 2936 2959
rect 3151 2959 3152 2960
rect 3156 2959 3157 2963
rect 3151 2958 3157 2959
rect 3162 2963 3168 2964
rect 3162 2959 3163 2963
rect 3167 2962 3168 2963
rect 3399 2963 3405 2964
rect 3399 2962 3400 2963
rect 3167 2960 3400 2962
rect 3167 2959 3168 2960
rect 3162 2958 3168 2959
rect 3399 2959 3400 2960
rect 3404 2959 3405 2963
rect 3399 2958 3405 2959
rect 3410 2963 3416 2964
rect 3410 2959 3411 2963
rect 3415 2962 3416 2963
rect 3663 2963 3669 2964
rect 3663 2962 3664 2963
rect 3415 2960 3664 2962
rect 3415 2959 3416 2960
rect 3410 2958 3416 2959
rect 3663 2959 3664 2960
rect 3668 2959 3669 2963
rect 3663 2958 3669 2959
rect 3903 2963 3909 2964
rect 3903 2959 3904 2963
rect 3908 2962 3909 2963
rect 3914 2963 3920 2964
rect 3914 2962 3915 2963
rect 3908 2960 3915 2962
rect 3908 2959 3909 2960
rect 3903 2958 3909 2959
rect 3914 2959 3915 2960
rect 3919 2959 3920 2963
rect 3914 2958 3920 2959
rect 2006 2956 2012 2957
rect 274 2955 280 2956
rect 274 2951 275 2955
rect 279 2954 280 2955
rect 426 2955 432 2956
rect 279 2952 385 2954
rect 279 2951 280 2952
rect 274 2950 280 2951
rect 426 2951 427 2955
rect 431 2954 432 2955
rect 647 2955 653 2956
rect 647 2954 648 2955
rect 431 2952 481 2954
rect 621 2952 648 2954
rect 431 2951 432 2952
rect 426 2950 432 2951
rect 647 2951 648 2952
rect 652 2951 653 2955
rect 647 2950 653 2951
rect 730 2955 736 2956
rect 730 2951 731 2955
rect 735 2951 736 2955
rect 730 2950 736 2951
rect 858 2955 864 2956
rect 858 2951 859 2955
rect 863 2951 864 2955
rect 858 2950 864 2951
rect 1010 2955 1016 2956
rect 1010 2951 1011 2955
rect 1015 2951 1016 2955
rect 1010 2950 1016 2951
rect 1178 2955 1184 2956
rect 1178 2951 1179 2955
rect 1183 2951 1184 2955
rect 1178 2950 1184 2951
rect 1370 2955 1376 2956
rect 1370 2951 1371 2955
rect 1375 2951 1376 2955
rect 1370 2950 1376 2951
rect 1570 2955 1576 2956
rect 1570 2951 1571 2955
rect 1575 2951 1576 2955
rect 1570 2950 1576 2951
rect 1786 2955 1792 2956
rect 1786 2951 1787 2955
rect 1791 2951 1792 2955
rect 1786 2950 1792 2951
rect 1794 2955 1800 2956
rect 1794 2951 1795 2955
rect 1799 2954 1800 2955
rect 2924 2954 2926 2958
rect 3362 2955 3368 2956
rect 3362 2954 3363 2955
rect 1799 2952 1945 2954
rect 2924 2952 3363 2954
rect 1799 2951 1800 2952
rect 1794 2950 1800 2951
rect 3362 2951 3363 2952
rect 3367 2951 3368 2955
rect 3362 2950 3368 2951
rect 2135 2947 2144 2948
rect 342 2945 348 2946
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 342 2941 343 2945
rect 347 2941 348 2945
rect 342 2940 348 2941
rect 438 2945 444 2946
rect 438 2941 439 2945
rect 443 2941 444 2945
rect 438 2940 444 2941
rect 542 2945 548 2946
rect 542 2941 543 2945
rect 547 2941 548 2945
rect 542 2940 548 2941
rect 654 2945 660 2946
rect 654 2941 655 2945
rect 659 2941 660 2945
rect 654 2940 660 2941
rect 782 2945 788 2946
rect 782 2941 783 2945
rect 787 2941 788 2945
rect 782 2940 788 2941
rect 934 2945 940 2946
rect 934 2941 935 2945
rect 939 2941 940 2945
rect 934 2940 940 2941
rect 1102 2945 1108 2946
rect 1102 2941 1103 2945
rect 1107 2941 1108 2945
rect 1102 2940 1108 2941
rect 1294 2945 1300 2946
rect 1294 2941 1295 2945
rect 1299 2941 1300 2945
rect 1294 2940 1300 2941
rect 1494 2945 1500 2946
rect 1494 2941 1495 2945
rect 1499 2941 1500 2945
rect 1494 2940 1500 2941
rect 1710 2945 1716 2946
rect 1710 2941 1711 2945
rect 1715 2941 1716 2945
rect 1710 2940 1716 2941
rect 1902 2945 1908 2946
rect 1902 2941 1903 2945
rect 1907 2941 1908 2945
rect 1902 2940 1908 2941
rect 2006 2944 2012 2945
rect 2006 2940 2007 2944
rect 2011 2940 2012 2944
rect 2135 2943 2136 2947
rect 2143 2943 2144 2947
rect 2135 2942 2144 2943
rect 2327 2947 2333 2948
rect 2327 2943 2328 2947
rect 2332 2946 2333 2947
rect 2338 2947 2344 2948
rect 2332 2944 2334 2946
rect 2332 2943 2336 2944
rect 2327 2942 2331 2943
rect 110 2939 116 2940
rect 2006 2939 2012 2940
rect 2330 2939 2331 2942
rect 2335 2939 2336 2943
rect 2338 2943 2339 2947
rect 2343 2946 2344 2947
rect 2551 2947 2557 2948
rect 2551 2946 2552 2947
rect 2343 2944 2552 2946
rect 2343 2943 2344 2944
rect 2338 2942 2344 2943
rect 2551 2943 2552 2944
rect 2556 2943 2557 2947
rect 2551 2942 2557 2943
rect 2562 2947 2568 2948
rect 2562 2943 2563 2947
rect 2567 2946 2568 2947
rect 2799 2947 2805 2948
rect 2799 2946 2800 2947
rect 2567 2944 2800 2946
rect 2567 2943 2568 2944
rect 2562 2942 2568 2943
rect 2799 2943 2800 2944
rect 2804 2943 2805 2947
rect 2799 2942 2805 2943
rect 2810 2947 2816 2948
rect 2810 2943 2811 2947
rect 2815 2946 2816 2947
rect 3063 2947 3069 2948
rect 3063 2946 3064 2947
rect 2815 2944 3064 2946
rect 2815 2943 2816 2944
rect 2810 2942 2816 2943
rect 3063 2943 3064 2944
rect 3068 2943 3069 2947
rect 3063 2942 3069 2943
rect 3074 2947 3080 2948
rect 3074 2943 3075 2947
rect 3079 2946 3080 2947
rect 3343 2947 3349 2948
rect 3343 2946 3344 2947
rect 3079 2944 3344 2946
rect 3079 2943 3080 2944
rect 3074 2942 3080 2943
rect 3343 2943 3344 2944
rect 3348 2943 3349 2947
rect 3343 2942 3349 2943
rect 3354 2947 3360 2948
rect 3354 2943 3355 2947
rect 3359 2946 3360 2947
rect 3631 2947 3637 2948
rect 3631 2946 3632 2947
rect 3359 2944 3632 2946
rect 3359 2943 3360 2944
rect 3354 2942 3360 2943
rect 3631 2943 3632 2944
rect 3636 2943 3637 2947
rect 3631 2942 3637 2943
rect 3903 2947 3912 2948
rect 3903 2943 3904 2947
rect 3911 2943 3912 2947
rect 3903 2942 3912 2943
rect 2330 2938 2336 2939
rect 2046 2928 2052 2929
rect 3942 2928 3948 2929
rect 2046 2924 2047 2928
rect 2051 2924 2052 2928
rect 407 2923 413 2924
rect 407 2919 408 2923
rect 412 2922 413 2923
rect 426 2923 432 2924
rect 426 2922 427 2923
rect 412 2920 427 2922
rect 412 2919 413 2920
rect 407 2918 413 2919
rect 426 2919 427 2920
rect 431 2919 432 2923
rect 426 2918 432 2919
rect 503 2923 509 2924
rect 503 2919 504 2923
rect 508 2922 509 2923
rect 514 2923 520 2924
rect 514 2922 515 2923
rect 508 2920 515 2922
rect 508 2919 509 2920
rect 503 2918 509 2919
rect 514 2919 515 2920
rect 519 2919 520 2923
rect 514 2918 520 2919
rect 607 2923 613 2924
rect 607 2919 608 2923
rect 612 2922 613 2923
rect 642 2923 648 2924
rect 642 2922 643 2923
rect 612 2920 643 2922
rect 612 2919 613 2920
rect 607 2918 613 2919
rect 642 2919 643 2920
rect 647 2919 648 2923
rect 642 2918 648 2919
rect 655 2923 661 2924
rect 655 2919 656 2923
rect 660 2922 661 2923
rect 719 2923 725 2924
rect 719 2922 720 2923
rect 660 2920 720 2922
rect 660 2919 661 2920
rect 655 2918 661 2919
rect 719 2919 720 2920
rect 724 2919 725 2923
rect 719 2918 725 2919
rect 730 2923 736 2924
rect 730 2919 731 2923
rect 735 2922 736 2923
rect 847 2923 853 2924
rect 847 2922 848 2923
rect 735 2920 848 2922
rect 735 2919 736 2920
rect 730 2918 736 2919
rect 847 2919 848 2920
rect 852 2919 853 2923
rect 847 2918 853 2919
rect 990 2923 996 2924
rect 990 2919 991 2923
rect 995 2922 996 2923
rect 999 2923 1005 2924
rect 999 2922 1000 2923
rect 995 2920 1000 2922
rect 995 2919 996 2920
rect 990 2918 996 2919
rect 999 2919 1000 2920
rect 1004 2919 1005 2923
rect 999 2918 1005 2919
rect 1010 2923 1016 2924
rect 1010 2919 1011 2923
rect 1015 2922 1016 2923
rect 1167 2923 1173 2924
rect 1167 2922 1168 2923
rect 1015 2920 1168 2922
rect 1015 2919 1016 2920
rect 1010 2918 1016 2919
rect 1167 2919 1168 2920
rect 1172 2919 1173 2923
rect 1167 2918 1173 2919
rect 1178 2923 1184 2924
rect 1178 2919 1179 2923
rect 1183 2922 1184 2923
rect 1359 2923 1365 2924
rect 1359 2922 1360 2923
rect 1183 2920 1360 2922
rect 1183 2919 1184 2920
rect 1178 2918 1184 2919
rect 1359 2919 1360 2920
rect 1364 2919 1365 2923
rect 1359 2918 1365 2919
rect 1370 2923 1376 2924
rect 1370 2919 1371 2923
rect 1375 2922 1376 2923
rect 1559 2923 1565 2924
rect 1559 2922 1560 2923
rect 1375 2920 1560 2922
rect 1375 2919 1376 2920
rect 1370 2918 1376 2919
rect 1559 2919 1560 2920
rect 1564 2919 1565 2923
rect 1559 2918 1565 2919
rect 1775 2923 1781 2924
rect 1775 2919 1776 2923
rect 1780 2922 1781 2923
rect 1794 2923 1800 2924
rect 1794 2922 1795 2923
rect 1780 2920 1795 2922
rect 1780 2919 1781 2920
rect 1775 2918 1781 2919
rect 1794 2919 1795 2920
rect 1799 2919 1800 2923
rect 1794 2918 1800 2919
rect 1967 2923 1973 2924
rect 2046 2923 2052 2924
rect 2070 2927 2076 2928
rect 2070 2923 2071 2927
rect 2075 2923 2076 2927
rect 1967 2919 1968 2923
rect 1972 2922 1973 2923
rect 2070 2922 2076 2923
rect 2262 2927 2268 2928
rect 2262 2923 2263 2927
rect 2267 2923 2268 2927
rect 2262 2922 2268 2923
rect 2486 2927 2492 2928
rect 2486 2923 2487 2927
rect 2491 2923 2492 2927
rect 2486 2922 2492 2923
rect 2734 2927 2740 2928
rect 2734 2923 2735 2927
rect 2739 2923 2740 2927
rect 2734 2922 2740 2923
rect 2998 2927 3004 2928
rect 2998 2923 2999 2927
rect 3003 2923 3004 2927
rect 2998 2922 3004 2923
rect 3278 2927 3284 2928
rect 3278 2923 3279 2927
rect 3283 2923 3284 2927
rect 3278 2922 3284 2923
rect 3566 2927 3572 2928
rect 3566 2923 3567 2927
rect 3571 2923 3572 2927
rect 3566 2922 3572 2923
rect 3838 2927 3844 2928
rect 3838 2923 3839 2927
rect 3843 2923 3844 2927
rect 3942 2924 3943 2928
rect 3947 2924 3948 2928
rect 3942 2923 3948 2924
rect 3838 2922 3844 2923
rect 1972 2920 2001 2922
rect 1972 2919 1973 2920
rect 1967 2918 1973 2919
rect 1999 2918 2001 2920
rect 2338 2919 2344 2920
rect 1999 2916 2113 2918
rect 2338 2915 2339 2919
rect 2343 2915 2344 2919
rect 2338 2914 2344 2915
rect 2562 2919 2568 2920
rect 2562 2915 2563 2919
rect 2567 2915 2568 2919
rect 2562 2914 2568 2915
rect 2810 2919 2816 2920
rect 2810 2915 2811 2919
rect 2815 2915 2816 2919
rect 2810 2914 2816 2915
rect 3074 2919 3080 2920
rect 3074 2915 3075 2919
rect 3079 2915 3080 2919
rect 3074 2914 3080 2915
rect 3354 2919 3360 2920
rect 3354 2915 3355 2919
rect 3359 2915 3360 2919
rect 3354 2914 3360 2915
rect 3362 2919 3368 2920
rect 3362 2915 3363 2919
rect 3367 2918 3368 2919
rect 3367 2916 3609 2918
rect 3367 2915 3368 2916
rect 3362 2914 3368 2915
rect 3914 2915 3920 2916
rect 271 2911 280 2912
rect 271 2907 272 2911
rect 279 2907 280 2911
rect 271 2906 280 2907
rect 282 2911 288 2912
rect 282 2907 283 2911
rect 287 2910 288 2911
rect 391 2911 397 2912
rect 391 2910 392 2911
rect 287 2908 392 2910
rect 287 2907 288 2908
rect 282 2906 288 2907
rect 391 2907 392 2908
rect 396 2907 397 2911
rect 391 2906 397 2907
rect 402 2911 408 2912
rect 402 2907 403 2911
rect 407 2910 408 2911
rect 511 2911 517 2912
rect 511 2910 512 2911
rect 407 2908 512 2910
rect 407 2907 408 2908
rect 402 2906 408 2907
rect 511 2907 512 2908
rect 516 2907 517 2911
rect 511 2906 517 2907
rect 639 2911 645 2912
rect 639 2907 640 2911
rect 644 2910 645 2911
rect 663 2911 669 2912
rect 663 2910 664 2911
rect 644 2908 664 2910
rect 644 2907 645 2908
rect 639 2906 645 2907
rect 663 2907 664 2908
rect 668 2907 669 2911
rect 663 2906 669 2907
rect 767 2911 776 2912
rect 767 2907 768 2911
rect 775 2907 776 2911
rect 767 2906 776 2907
rect 911 2911 917 2912
rect 911 2907 912 2911
rect 916 2910 917 2911
rect 946 2911 952 2912
rect 946 2910 947 2911
rect 916 2908 947 2910
rect 916 2907 917 2908
rect 911 2906 917 2907
rect 946 2907 947 2908
rect 951 2907 952 2911
rect 946 2906 952 2907
rect 974 2911 980 2912
rect 974 2907 975 2911
rect 979 2910 980 2911
rect 1063 2911 1069 2912
rect 1063 2910 1064 2911
rect 979 2908 1064 2910
rect 979 2907 980 2908
rect 974 2906 980 2907
rect 1063 2907 1064 2908
rect 1068 2907 1069 2911
rect 1063 2906 1069 2907
rect 1231 2911 1237 2912
rect 1231 2907 1232 2911
rect 1236 2910 1237 2911
rect 1250 2911 1256 2912
rect 1250 2910 1251 2911
rect 1236 2908 1251 2910
rect 1236 2907 1237 2908
rect 1231 2906 1237 2907
rect 1250 2907 1251 2908
rect 1255 2907 1256 2911
rect 1250 2906 1256 2907
rect 1415 2911 1421 2912
rect 1415 2907 1416 2911
rect 1420 2910 1421 2911
rect 1438 2911 1444 2912
rect 1438 2910 1439 2911
rect 1420 2908 1439 2910
rect 1420 2907 1421 2908
rect 1415 2906 1421 2907
rect 1438 2907 1439 2908
rect 1443 2907 1444 2911
rect 1438 2906 1444 2907
rect 1570 2911 1576 2912
rect 1570 2907 1571 2911
rect 1575 2910 1576 2911
rect 1599 2911 1605 2912
rect 1599 2910 1600 2911
rect 1575 2908 1600 2910
rect 1575 2907 1576 2908
rect 1570 2906 1576 2907
rect 1599 2907 1600 2908
rect 1604 2907 1605 2911
rect 1599 2906 1605 2907
rect 1786 2911 1797 2912
rect 1786 2907 1787 2911
rect 1791 2907 1792 2911
rect 1796 2907 1797 2911
rect 1786 2906 1797 2907
rect 1802 2911 1808 2912
rect 1802 2907 1803 2911
rect 1807 2910 1808 2911
rect 1967 2911 1973 2912
rect 1967 2910 1968 2911
rect 1807 2908 1968 2910
rect 1807 2907 1808 2908
rect 1802 2906 1808 2907
rect 1967 2907 1968 2908
rect 1972 2907 1973 2911
rect 1967 2906 1973 2907
rect 2046 2911 2052 2912
rect 2046 2907 2047 2911
rect 2051 2907 2052 2911
rect 3914 2911 3915 2915
rect 3919 2911 3920 2915
rect 3914 2910 3920 2911
rect 3942 2911 3948 2912
rect 2046 2906 2052 2907
rect 2070 2908 2076 2909
rect 2070 2904 2071 2908
rect 2075 2904 2076 2908
rect 2070 2903 2076 2904
rect 2262 2908 2268 2909
rect 2262 2904 2263 2908
rect 2267 2904 2268 2908
rect 2262 2903 2268 2904
rect 2486 2908 2492 2909
rect 2486 2904 2487 2908
rect 2491 2904 2492 2908
rect 2486 2903 2492 2904
rect 2734 2908 2740 2909
rect 2734 2904 2735 2908
rect 2739 2904 2740 2908
rect 2734 2903 2740 2904
rect 2998 2908 3004 2909
rect 2998 2904 2999 2908
rect 3003 2904 3004 2908
rect 2998 2903 3004 2904
rect 3278 2908 3284 2909
rect 3278 2904 3279 2908
rect 3283 2904 3284 2908
rect 3278 2903 3284 2904
rect 3566 2908 3572 2909
rect 3566 2904 3567 2908
rect 3571 2904 3572 2908
rect 3566 2903 3572 2904
rect 3838 2908 3844 2909
rect 3838 2904 3839 2908
rect 3843 2904 3844 2908
rect 3942 2907 3943 2911
rect 3947 2907 3948 2911
rect 3942 2906 3948 2907
rect 3838 2903 3844 2904
rect 110 2892 116 2893
rect 2006 2892 2012 2893
rect 110 2888 111 2892
rect 115 2888 116 2892
rect 110 2887 116 2888
rect 206 2891 212 2892
rect 206 2887 207 2891
rect 211 2887 212 2891
rect 206 2886 212 2887
rect 326 2891 332 2892
rect 326 2887 327 2891
rect 331 2887 332 2891
rect 326 2886 332 2887
rect 446 2891 452 2892
rect 446 2887 447 2891
rect 451 2887 452 2891
rect 446 2886 452 2887
rect 574 2891 580 2892
rect 574 2887 575 2891
rect 579 2887 580 2891
rect 702 2891 708 2892
rect 574 2886 580 2887
rect 642 2887 648 2888
rect 282 2883 288 2884
rect 282 2879 283 2883
rect 287 2879 288 2883
rect 282 2878 288 2879
rect 402 2883 408 2884
rect 402 2879 403 2883
rect 407 2879 408 2883
rect 642 2883 643 2887
rect 647 2886 648 2887
rect 702 2887 703 2891
rect 707 2887 708 2891
rect 702 2886 708 2887
rect 846 2891 852 2892
rect 846 2887 847 2891
rect 851 2887 852 2891
rect 846 2886 852 2887
rect 998 2891 1004 2892
rect 998 2887 999 2891
rect 1003 2887 1004 2891
rect 998 2886 1004 2887
rect 1166 2891 1172 2892
rect 1166 2887 1167 2891
rect 1171 2887 1172 2891
rect 1166 2886 1172 2887
rect 1350 2891 1356 2892
rect 1350 2887 1351 2891
rect 1355 2887 1356 2891
rect 1350 2886 1356 2887
rect 1534 2891 1540 2892
rect 1534 2887 1535 2891
rect 1539 2887 1540 2891
rect 1534 2886 1540 2887
rect 1726 2891 1732 2892
rect 1726 2887 1727 2891
rect 1731 2887 1732 2891
rect 1726 2886 1732 2887
rect 1902 2891 1908 2892
rect 1902 2887 1903 2891
rect 1907 2887 1908 2891
rect 2006 2888 2007 2892
rect 2011 2888 2012 2892
rect 2006 2887 2012 2888
rect 1902 2886 1908 2887
rect 647 2884 654 2886
rect 647 2883 648 2884
rect 642 2882 648 2883
rect 652 2881 654 2884
rect 663 2883 669 2884
rect 402 2878 408 2879
rect 522 2879 528 2880
rect 110 2875 116 2876
rect 110 2871 111 2875
rect 115 2871 116 2875
rect 522 2875 523 2879
rect 527 2875 528 2879
rect 663 2879 664 2883
rect 668 2882 669 2883
rect 974 2883 980 2884
rect 974 2882 975 2883
rect 668 2880 745 2882
rect 925 2880 975 2882
rect 668 2879 669 2880
rect 663 2878 669 2879
rect 974 2879 975 2880
rect 979 2879 980 2883
rect 974 2878 980 2879
rect 990 2883 996 2884
rect 990 2879 991 2883
rect 995 2882 996 2883
rect 1250 2883 1256 2884
rect 995 2880 1041 2882
rect 995 2879 996 2880
rect 990 2878 996 2879
rect 1242 2879 1248 2880
rect 522 2874 528 2875
rect 1242 2875 1243 2879
rect 1247 2875 1248 2879
rect 1250 2879 1251 2883
rect 1255 2882 1256 2883
rect 1438 2883 1444 2884
rect 1255 2880 1393 2882
rect 1255 2879 1256 2880
rect 1250 2878 1256 2879
rect 1438 2879 1439 2883
rect 1443 2882 1444 2883
rect 1802 2883 1808 2884
rect 1443 2880 1577 2882
rect 1443 2879 1444 2880
rect 1438 2878 1444 2879
rect 1802 2879 1803 2883
rect 1807 2879 1808 2883
rect 1802 2878 1808 2879
rect 1818 2883 1824 2884
rect 1818 2879 1819 2883
rect 1823 2882 1824 2883
rect 1823 2880 1945 2882
rect 1823 2879 1824 2880
rect 1818 2878 1824 2879
rect 1242 2874 1248 2875
rect 2006 2875 2012 2876
rect 110 2870 116 2871
rect 206 2872 212 2873
rect 206 2868 207 2872
rect 211 2868 212 2872
rect 206 2867 212 2868
rect 326 2872 332 2873
rect 326 2868 327 2872
rect 331 2868 332 2872
rect 326 2867 332 2868
rect 446 2872 452 2873
rect 446 2868 447 2872
rect 451 2868 452 2872
rect 446 2867 452 2868
rect 574 2872 580 2873
rect 574 2868 575 2872
rect 579 2868 580 2872
rect 574 2867 580 2868
rect 702 2872 708 2873
rect 702 2868 703 2872
rect 707 2868 708 2872
rect 702 2867 708 2868
rect 846 2872 852 2873
rect 846 2868 847 2872
rect 851 2868 852 2872
rect 846 2867 852 2868
rect 998 2872 1004 2873
rect 998 2868 999 2872
rect 1003 2868 1004 2872
rect 998 2867 1004 2868
rect 1166 2872 1172 2873
rect 1166 2868 1167 2872
rect 1171 2868 1172 2872
rect 1166 2867 1172 2868
rect 1350 2872 1356 2873
rect 1350 2868 1351 2872
rect 1355 2868 1356 2872
rect 1350 2867 1356 2868
rect 1534 2872 1540 2873
rect 1534 2868 1535 2872
rect 1539 2868 1540 2872
rect 1534 2867 1540 2868
rect 1726 2872 1732 2873
rect 1726 2868 1727 2872
rect 1731 2868 1732 2872
rect 1726 2867 1732 2868
rect 1902 2872 1908 2873
rect 1902 2868 1903 2872
rect 1907 2868 1908 2872
rect 2006 2871 2007 2875
rect 2011 2871 2012 2875
rect 2006 2870 2012 2871
rect 1902 2867 1908 2868
rect 2359 2844 2974 2846
rect 2046 2837 2052 2838
rect 2046 2833 2047 2837
rect 2051 2833 2052 2837
rect 2046 2832 2052 2833
rect 2330 2831 2336 2832
rect 2330 2827 2331 2831
rect 2335 2830 2336 2831
rect 2359 2830 2361 2844
rect 2670 2840 2676 2841
rect 2670 2836 2671 2840
rect 2675 2836 2676 2840
rect 2670 2835 2676 2836
rect 2886 2840 2892 2841
rect 2886 2836 2887 2840
rect 2891 2836 2892 2840
rect 2886 2835 2892 2836
rect 2335 2828 2361 2830
rect 2746 2831 2752 2832
rect 2335 2827 2336 2828
rect 2330 2826 2336 2827
rect 2746 2827 2747 2831
rect 2751 2827 2752 2831
rect 2746 2826 2752 2827
rect 2962 2831 2968 2832
rect 2962 2827 2963 2831
rect 2967 2827 2968 2831
rect 2972 2830 2974 2844
rect 3094 2840 3100 2841
rect 3094 2836 3095 2840
rect 3099 2836 3100 2840
rect 3094 2835 3100 2836
rect 3286 2840 3292 2841
rect 3286 2836 3287 2840
rect 3291 2836 3292 2840
rect 3286 2835 3292 2836
rect 3478 2840 3484 2841
rect 3478 2836 3479 2840
rect 3483 2836 3484 2840
rect 3478 2835 3484 2836
rect 3670 2840 3676 2841
rect 3670 2836 3671 2840
rect 3675 2836 3676 2840
rect 3670 2835 3676 2836
rect 3838 2840 3844 2841
rect 3838 2836 3839 2840
rect 3843 2836 3844 2840
rect 3838 2835 3844 2836
rect 3942 2837 3948 2838
rect 3942 2833 3943 2837
rect 3947 2833 3948 2837
rect 3942 2832 3948 2833
rect 3354 2831 3360 2832
rect 2972 2828 3137 2830
rect 2962 2826 2968 2827
rect 3354 2827 3355 2831
rect 3359 2827 3360 2831
rect 3354 2826 3360 2827
rect 3370 2831 3376 2832
rect 3370 2827 3371 2831
rect 3375 2830 3376 2831
rect 3754 2831 3760 2832
rect 3375 2828 3521 2830
rect 3375 2827 3376 2828
rect 3370 2826 3376 2827
rect 3748 2822 3750 2829
rect 3754 2827 3755 2831
rect 3759 2830 3760 2831
rect 3759 2828 3881 2830
rect 3759 2827 3760 2828
rect 3754 2826 3760 2827
rect 3759 2823 3765 2824
rect 3759 2822 3760 2823
rect 2670 2821 2676 2822
rect 2046 2820 2052 2821
rect 2046 2816 2047 2820
rect 2051 2816 2052 2820
rect 2670 2817 2671 2821
rect 2675 2817 2676 2821
rect 2670 2816 2676 2817
rect 2886 2821 2892 2822
rect 2886 2817 2887 2821
rect 2891 2817 2892 2821
rect 2886 2816 2892 2817
rect 3094 2821 3100 2822
rect 3094 2817 3095 2821
rect 3099 2817 3100 2821
rect 3094 2816 3100 2817
rect 3286 2821 3292 2822
rect 3286 2817 3287 2821
rect 3291 2817 3292 2821
rect 3286 2816 3292 2817
rect 3478 2821 3484 2822
rect 3478 2817 3479 2821
rect 3483 2817 3484 2821
rect 3478 2816 3484 2817
rect 3670 2821 3676 2822
rect 3670 2817 3671 2821
rect 3675 2817 3676 2821
rect 3748 2820 3760 2822
rect 3759 2819 3760 2820
rect 3764 2819 3765 2823
rect 3759 2818 3765 2819
rect 3838 2821 3844 2822
rect 3670 2816 3676 2817
rect 3838 2817 3839 2821
rect 3843 2817 3844 2821
rect 3838 2816 3844 2817
rect 3942 2820 3948 2821
rect 3942 2816 3943 2820
rect 3947 2816 3948 2820
rect 2046 2815 2052 2816
rect 3942 2815 3948 2816
rect 134 2808 140 2809
rect 110 2805 116 2806
rect 110 2801 111 2805
rect 115 2801 116 2805
rect 134 2804 135 2808
rect 139 2804 140 2808
rect 134 2803 140 2804
rect 246 2808 252 2809
rect 246 2804 247 2808
rect 251 2804 252 2808
rect 246 2803 252 2804
rect 398 2808 404 2809
rect 398 2804 399 2808
rect 403 2804 404 2808
rect 398 2803 404 2804
rect 550 2808 556 2809
rect 550 2804 551 2808
rect 555 2804 556 2808
rect 550 2803 556 2804
rect 710 2808 716 2809
rect 710 2804 711 2808
rect 715 2804 716 2808
rect 710 2803 716 2804
rect 878 2808 884 2809
rect 878 2804 879 2808
rect 883 2804 884 2808
rect 878 2803 884 2804
rect 1046 2808 1052 2809
rect 1046 2804 1047 2808
rect 1051 2804 1052 2808
rect 1046 2803 1052 2804
rect 1222 2808 1228 2809
rect 1222 2804 1223 2808
rect 1227 2804 1228 2808
rect 1222 2803 1228 2804
rect 1398 2808 1404 2809
rect 1398 2804 1399 2808
rect 1403 2804 1404 2808
rect 1398 2803 1404 2804
rect 1574 2808 1580 2809
rect 1574 2804 1575 2808
rect 1579 2804 1580 2808
rect 1574 2803 1580 2804
rect 1750 2808 1756 2809
rect 1750 2804 1751 2808
rect 1755 2804 1756 2808
rect 1750 2803 1756 2804
rect 1902 2808 1908 2809
rect 1902 2804 1903 2808
rect 1907 2804 1908 2808
rect 1902 2803 1908 2804
rect 2006 2805 2012 2806
rect 110 2800 116 2801
rect 2006 2801 2007 2805
rect 2011 2801 2012 2805
rect 2006 2800 2012 2801
rect 202 2799 208 2800
rect 202 2795 203 2799
rect 207 2795 208 2799
rect 202 2794 208 2795
rect 218 2799 224 2800
rect 218 2795 219 2799
rect 223 2798 224 2799
rect 378 2799 384 2800
rect 223 2796 289 2798
rect 223 2795 224 2796
rect 218 2794 224 2795
rect 378 2795 379 2799
rect 383 2798 384 2799
rect 682 2799 688 2800
rect 682 2798 683 2799
rect 383 2796 441 2798
rect 629 2796 683 2798
rect 383 2795 384 2796
rect 378 2794 384 2795
rect 682 2795 683 2796
rect 687 2795 688 2799
rect 682 2794 688 2795
rect 778 2799 784 2800
rect 778 2795 779 2799
rect 783 2795 784 2799
rect 778 2794 784 2795
rect 946 2799 952 2800
rect 946 2795 947 2799
rect 951 2795 952 2799
rect 946 2794 952 2795
rect 962 2799 968 2800
rect 962 2795 963 2799
rect 967 2798 968 2799
rect 1298 2799 1304 2800
rect 967 2796 1089 2798
rect 967 2795 968 2796
rect 962 2794 968 2795
rect 1298 2795 1299 2799
rect 1303 2795 1304 2799
rect 1298 2794 1304 2795
rect 1474 2799 1480 2800
rect 1474 2795 1475 2799
rect 1479 2795 1480 2799
rect 1474 2794 1480 2795
rect 1650 2799 1656 2800
rect 1650 2795 1651 2799
rect 1655 2795 1656 2799
rect 1650 2794 1656 2795
rect 1826 2799 1832 2800
rect 1826 2795 1827 2799
rect 1831 2795 1832 2799
rect 2682 2799 2688 2800
rect 1981 2796 2001 2798
rect 1826 2794 1832 2795
rect 1999 2794 2001 2796
rect 2682 2795 2683 2799
rect 2687 2798 2688 2799
rect 2735 2799 2741 2800
rect 2735 2798 2736 2799
rect 2687 2796 2736 2798
rect 2687 2795 2688 2796
rect 2682 2794 2688 2795
rect 2735 2795 2736 2796
rect 2740 2795 2741 2799
rect 2735 2794 2741 2795
rect 2746 2799 2752 2800
rect 2746 2795 2747 2799
rect 2751 2798 2752 2799
rect 2951 2799 2957 2800
rect 2951 2798 2952 2799
rect 2751 2796 2952 2798
rect 2751 2795 2752 2796
rect 2746 2794 2752 2795
rect 2951 2795 2952 2796
rect 2956 2795 2957 2799
rect 2951 2794 2957 2795
rect 2962 2799 2968 2800
rect 2962 2795 2963 2799
rect 2967 2798 2968 2799
rect 3159 2799 3165 2800
rect 3159 2798 3160 2799
rect 2967 2796 3160 2798
rect 2967 2795 2968 2796
rect 2962 2794 2968 2795
rect 3159 2795 3160 2796
rect 3164 2795 3165 2799
rect 3159 2794 3165 2795
rect 3351 2799 3357 2800
rect 3351 2795 3352 2799
rect 3356 2798 3357 2799
rect 3370 2799 3376 2800
rect 3370 2798 3371 2799
rect 3356 2796 3371 2798
rect 3356 2795 3357 2796
rect 3351 2794 3357 2795
rect 3370 2795 3371 2796
rect 3375 2795 3376 2799
rect 3370 2794 3376 2795
rect 3522 2799 3528 2800
rect 3522 2795 3523 2799
rect 3527 2798 3528 2799
rect 3543 2799 3549 2800
rect 3543 2798 3544 2799
rect 3527 2796 3544 2798
rect 3527 2795 3528 2796
rect 3522 2794 3528 2795
rect 3543 2795 3544 2796
rect 3548 2795 3549 2799
rect 3543 2794 3549 2795
rect 3735 2799 3741 2800
rect 3735 2795 3736 2799
rect 3740 2798 3741 2799
rect 3754 2799 3760 2800
rect 3754 2798 3755 2799
rect 3740 2796 3755 2798
rect 3740 2795 3741 2796
rect 3735 2794 3741 2795
rect 3754 2795 3755 2796
rect 3759 2795 3760 2799
rect 3754 2794 3760 2795
rect 3903 2799 3912 2800
rect 3903 2795 3904 2799
rect 3911 2795 3912 2799
rect 3903 2794 3912 2795
rect 1999 2792 2070 2794
rect 134 2789 140 2790
rect 110 2788 116 2789
rect 110 2784 111 2788
rect 115 2784 116 2788
rect 134 2785 135 2789
rect 139 2785 140 2789
rect 134 2784 140 2785
rect 246 2789 252 2790
rect 246 2785 247 2789
rect 251 2785 252 2789
rect 246 2784 252 2785
rect 398 2789 404 2790
rect 398 2785 399 2789
rect 403 2785 404 2789
rect 398 2784 404 2785
rect 550 2789 556 2790
rect 550 2785 551 2789
rect 555 2785 556 2789
rect 550 2784 556 2785
rect 710 2789 716 2790
rect 710 2785 711 2789
rect 715 2785 716 2789
rect 710 2784 716 2785
rect 878 2789 884 2790
rect 878 2785 879 2789
rect 883 2785 884 2789
rect 878 2784 884 2785
rect 1046 2789 1052 2790
rect 1046 2785 1047 2789
rect 1051 2785 1052 2789
rect 1046 2784 1052 2785
rect 1222 2789 1228 2790
rect 1222 2785 1223 2789
rect 1227 2785 1228 2789
rect 1222 2784 1228 2785
rect 1398 2789 1404 2790
rect 1398 2785 1399 2789
rect 1403 2785 1404 2789
rect 1398 2784 1404 2785
rect 1574 2789 1580 2790
rect 1574 2785 1575 2789
rect 1579 2785 1580 2789
rect 1574 2784 1580 2785
rect 1750 2789 1756 2790
rect 1750 2785 1751 2789
rect 1755 2785 1756 2789
rect 1750 2784 1756 2785
rect 1902 2789 1908 2790
rect 1902 2785 1903 2789
rect 1907 2785 1908 2789
rect 1902 2784 1908 2785
rect 2006 2788 2012 2789
rect 2006 2784 2007 2788
rect 2011 2784 2012 2788
rect 2068 2786 2070 2792
rect 2135 2787 2141 2788
rect 2135 2786 2136 2787
rect 2068 2784 2136 2786
rect 110 2783 116 2784
rect 2006 2783 2012 2784
rect 2135 2783 2136 2784
rect 2140 2783 2141 2787
rect 2135 2782 2141 2783
rect 2146 2787 2152 2788
rect 2146 2783 2147 2787
rect 2151 2786 2152 2787
rect 2263 2787 2269 2788
rect 2263 2786 2264 2787
rect 2151 2784 2264 2786
rect 2151 2783 2152 2784
rect 2146 2782 2152 2783
rect 2263 2783 2264 2784
rect 2268 2783 2269 2787
rect 2263 2782 2269 2783
rect 2407 2787 2416 2788
rect 2407 2783 2408 2787
rect 2415 2783 2416 2787
rect 2407 2782 2416 2783
rect 2418 2787 2424 2788
rect 2418 2783 2419 2787
rect 2423 2786 2424 2787
rect 2543 2787 2549 2788
rect 2543 2786 2544 2787
rect 2423 2784 2544 2786
rect 2423 2783 2424 2784
rect 2418 2782 2424 2783
rect 2543 2783 2544 2784
rect 2548 2783 2549 2787
rect 2543 2782 2549 2783
rect 2554 2787 2560 2788
rect 2554 2783 2555 2787
rect 2559 2786 2560 2787
rect 2671 2787 2677 2788
rect 2671 2786 2672 2787
rect 2559 2784 2672 2786
rect 2559 2783 2560 2784
rect 2554 2782 2560 2783
rect 2671 2783 2672 2784
rect 2676 2783 2677 2787
rect 2671 2782 2677 2783
rect 2791 2787 2797 2788
rect 2791 2783 2792 2787
rect 2796 2786 2797 2787
rect 2822 2787 2828 2788
rect 2796 2784 2818 2786
rect 2796 2783 2797 2784
rect 2791 2782 2797 2783
rect 2816 2778 2818 2784
rect 2822 2783 2823 2787
rect 2827 2786 2828 2787
rect 2903 2787 2909 2788
rect 2903 2786 2904 2787
rect 2827 2784 2904 2786
rect 2827 2783 2828 2784
rect 2822 2782 2828 2783
rect 2903 2783 2904 2784
rect 2908 2783 2909 2787
rect 2903 2782 2909 2783
rect 3007 2787 3013 2788
rect 3007 2783 3008 2787
rect 3012 2786 3013 2787
rect 3039 2787 3045 2788
rect 3039 2786 3040 2787
rect 3012 2784 3040 2786
rect 3012 2783 3013 2784
rect 3007 2782 3013 2783
rect 3039 2783 3040 2784
rect 3044 2783 3045 2787
rect 3039 2782 3045 2783
rect 3111 2787 3117 2788
rect 3111 2783 3112 2787
rect 3116 2786 3117 2787
rect 3130 2787 3136 2788
rect 3130 2786 3131 2787
rect 3116 2784 3131 2786
rect 3116 2783 3117 2784
rect 3111 2782 3117 2783
rect 3130 2783 3131 2784
rect 3135 2783 3136 2787
rect 3130 2782 3136 2783
rect 3207 2787 3213 2788
rect 3207 2783 3208 2787
rect 3212 2786 3213 2787
rect 3231 2787 3237 2788
rect 3231 2786 3232 2787
rect 3212 2784 3232 2786
rect 3212 2783 3213 2784
rect 3207 2782 3213 2783
rect 3231 2783 3232 2784
rect 3236 2783 3237 2787
rect 3231 2782 3237 2783
rect 3303 2787 3309 2788
rect 3303 2783 3304 2787
rect 3308 2786 3309 2787
rect 3354 2787 3360 2788
rect 3354 2786 3355 2787
rect 3308 2784 3355 2786
rect 3308 2783 3309 2784
rect 3303 2782 3309 2783
rect 3354 2783 3355 2784
rect 3359 2783 3360 2787
rect 3354 2782 3360 2783
rect 3407 2787 3413 2788
rect 3407 2783 3408 2787
rect 3412 2786 3413 2787
rect 3418 2787 3424 2788
rect 3412 2783 3414 2786
rect 3407 2782 3414 2783
rect 3418 2783 3419 2787
rect 3423 2786 3424 2787
rect 3511 2787 3517 2788
rect 3511 2786 3512 2787
rect 3423 2784 3512 2786
rect 3423 2783 3424 2784
rect 3418 2782 3424 2783
rect 3511 2783 3512 2784
rect 3516 2783 3517 2787
rect 3511 2782 3517 2783
rect 3615 2787 3621 2788
rect 3615 2783 3616 2787
rect 3620 2786 3621 2787
rect 3639 2787 3645 2788
rect 3639 2786 3640 2787
rect 3620 2784 3640 2786
rect 3620 2783 3621 2784
rect 3615 2782 3621 2783
rect 3639 2783 3640 2784
rect 3644 2783 3645 2787
rect 3639 2782 3645 2783
rect 3711 2787 3717 2788
rect 3711 2783 3712 2787
rect 3716 2786 3717 2787
rect 3759 2787 3765 2788
rect 3716 2784 3754 2786
rect 3716 2783 3717 2784
rect 3711 2782 3717 2783
rect 2922 2779 2928 2780
rect 2922 2778 2923 2779
rect 2816 2776 2923 2778
rect 2922 2775 2923 2776
rect 2927 2775 2928 2779
rect 3412 2778 3414 2782
rect 3530 2779 3536 2780
rect 3530 2778 3531 2779
rect 3412 2776 3531 2778
rect 2922 2774 2928 2775
rect 3530 2775 3531 2776
rect 3535 2775 3536 2779
rect 3752 2778 3754 2784
rect 3759 2783 3760 2787
rect 3764 2786 3765 2787
rect 3807 2787 3813 2788
rect 3807 2786 3808 2787
rect 3764 2784 3808 2786
rect 3764 2783 3765 2784
rect 3759 2782 3765 2783
rect 3807 2783 3808 2784
rect 3812 2783 3813 2787
rect 3807 2782 3813 2783
rect 3818 2787 3824 2788
rect 3818 2783 3819 2787
rect 3823 2786 3824 2787
rect 3903 2787 3909 2788
rect 3903 2786 3904 2787
rect 3823 2784 3904 2786
rect 3823 2783 3824 2784
rect 3818 2782 3824 2783
rect 3903 2783 3904 2784
rect 3908 2783 3909 2787
rect 3903 2782 3909 2783
rect 3826 2779 3832 2780
rect 3826 2778 3827 2779
rect 3752 2776 3827 2778
rect 3530 2774 3536 2775
rect 3826 2775 3827 2776
rect 3831 2775 3832 2779
rect 3826 2774 3832 2775
rect 2046 2768 2052 2769
rect 3942 2768 3948 2769
rect 199 2767 205 2768
rect 199 2763 200 2767
rect 204 2766 205 2767
rect 218 2767 224 2768
rect 218 2766 219 2767
rect 204 2764 219 2766
rect 204 2763 205 2764
rect 199 2762 205 2763
rect 218 2763 219 2764
rect 223 2763 224 2767
rect 218 2762 224 2763
rect 311 2767 317 2768
rect 311 2763 312 2767
rect 316 2766 317 2767
rect 378 2767 384 2768
rect 378 2766 379 2767
rect 316 2764 379 2766
rect 316 2763 317 2764
rect 311 2762 317 2763
rect 378 2763 379 2764
rect 383 2763 384 2767
rect 378 2762 384 2763
rect 463 2767 469 2768
rect 463 2763 464 2767
rect 468 2766 469 2767
rect 522 2767 528 2768
rect 522 2766 523 2767
rect 468 2764 523 2766
rect 468 2763 469 2764
rect 463 2762 469 2763
rect 522 2763 523 2764
rect 527 2763 528 2767
rect 522 2762 528 2763
rect 615 2767 621 2768
rect 615 2763 616 2767
rect 620 2766 621 2767
rect 650 2767 656 2768
rect 650 2766 651 2767
rect 620 2764 651 2766
rect 620 2763 621 2764
rect 615 2762 621 2763
rect 650 2763 651 2764
rect 655 2763 656 2767
rect 650 2762 656 2763
rect 682 2767 688 2768
rect 682 2763 683 2767
rect 687 2766 688 2767
rect 775 2767 781 2768
rect 775 2766 776 2767
rect 687 2764 776 2766
rect 687 2763 688 2764
rect 682 2762 688 2763
rect 775 2763 776 2764
rect 780 2763 781 2767
rect 775 2762 781 2763
rect 943 2767 949 2768
rect 943 2763 944 2767
rect 948 2766 949 2767
rect 962 2767 968 2768
rect 962 2766 963 2767
rect 948 2764 963 2766
rect 948 2763 949 2764
rect 943 2762 949 2763
rect 962 2763 963 2764
rect 967 2763 968 2767
rect 962 2762 968 2763
rect 1111 2767 1117 2768
rect 1111 2763 1112 2767
rect 1116 2766 1117 2767
rect 1162 2767 1168 2768
rect 1162 2766 1163 2767
rect 1116 2764 1163 2766
rect 1116 2763 1117 2764
rect 1111 2762 1117 2763
rect 1162 2763 1163 2764
rect 1167 2763 1168 2767
rect 1162 2762 1168 2763
rect 1242 2767 1248 2768
rect 1242 2763 1243 2767
rect 1247 2766 1248 2767
rect 1287 2767 1293 2768
rect 1287 2766 1288 2767
rect 1247 2764 1288 2766
rect 1247 2763 1248 2764
rect 1242 2762 1248 2763
rect 1287 2763 1288 2764
rect 1292 2763 1293 2767
rect 1287 2762 1293 2763
rect 1298 2767 1304 2768
rect 1298 2763 1299 2767
rect 1303 2766 1304 2767
rect 1463 2767 1469 2768
rect 1463 2766 1464 2767
rect 1303 2764 1464 2766
rect 1303 2763 1304 2764
rect 1298 2762 1304 2763
rect 1463 2763 1464 2764
rect 1468 2763 1469 2767
rect 1463 2762 1469 2763
rect 1474 2767 1480 2768
rect 1474 2763 1475 2767
rect 1479 2766 1480 2767
rect 1639 2767 1645 2768
rect 1639 2766 1640 2767
rect 1479 2764 1640 2766
rect 1479 2763 1480 2764
rect 1474 2762 1480 2763
rect 1639 2763 1640 2764
rect 1644 2763 1645 2767
rect 1639 2762 1645 2763
rect 1815 2767 1824 2768
rect 1815 2763 1816 2767
rect 1823 2763 1824 2767
rect 1815 2762 1824 2763
rect 1826 2767 1832 2768
rect 1826 2763 1827 2767
rect 1831 2766 1832 2767
rect 1967 2767 1973 2768
rect 1967 2766 1968 2767
rect 1831 2764 1968 2766
rect 1831 2763 1832 2764
rect 1826 2762 1832 2763
rect 1967 2763 1968 2764
rect 1972 2763 1973 2767
rect 2046 2764 2047 2768
rect 2051 2764 2052 2768
rect 2046 2763 2052 2764
rect 2070 2767 2076 2768
rect 2070 2763 2071 2767
rect 2075 2763 2076 2767
rect 1967 2762 1973 2763
rect 2070 2762 2076 2763
rect 2198 2767 2204 2768
rect 2198 2763 2199 2767
rect 2203 2763 2204 2767
rect 2198 2762 2204 2763
rect 2342 2767 2348 2768
rect 2342 2763 2343 2767
rect 2347 2763 2348 2767
rect 2342 2762 2348 2763
rect 2478 2767 2484 2768
rect 2478 2763 2479 2767
rect 2483 2763 2484 2767
rect 2478 2762 2484 2763
rect 2606 2767 2612 2768
rect 2606 2763 2607 2767
rect 2611 2763 2612 2767
rect 2606 2762 2612 2763
rect 2726 2767 2732 2768
rect 2726 2763 2727 2767
rect 2731 2763 2732 2767
rect 2726 2762 2732 2763
rect 2838 2767 2844 2768
rect 2838 2763 2839 2767
rect 2843 2763 2844 2767
rect 2838 2762 2844 2763
rect 2942 2767 2948 2768
rect 2942 2763 2943 2767
rect 2947 2763 2948 2767
rect 2942 2762 2948 2763
rect 3046 2767 3052 2768
rect 3046 2763 3047 2767
rect 3051 2763 3052 2767
rect 3046 2762 3052 2763
rect 3142 2767 3148 2768
rect 3142 2763 3143 2767
rect 3147 2763 3148 2767
rect 3142 2762 3148 2763
rect 3238 2767 3244 2768
rect 3238 2763 3239 2767
rect 3243 2763 3244 2767
rect 3238 2762 3244 2763
rect 3342 2767 3348 2768
rect 3342 2763 3343 2767
rect 3347 2763 3348 2767
rect 3342 2762 3348 2763
rect 3446 2767 3452 2768
rect 3446 2763 3447 2767
rect 3451 2763 3452 2767
rect 3446 2762 3452 2763
rect 3550 2767 3556 2768
rect 3550 2763 3551 2767
rect 3555 2763 3556 2767
rect 3550 2762 3556 2763
rect 3646 2767 3652 2768
rect 3646 2763 3647 2767
rect 3651 2763 3652 2767
rect 3646 2762 3652 2763
rect 3742 2767 3748 2768
rect 3742 2763 3743 2767
rect 3747 2763 3748 2767
rect 3742 2762 3748 2763
rect 3838 2767 3844 2768
rect 3838 2763 3839 2767
rect 3843 2763 3844 2767
rect 3942 2764 3943 2768
rect 3947 2764 3948 2768
rect 3942 2763 3948 2764
rect 3838 2762 3844 2763
rect 2146 2759 2152 2760
rect 2146 2755 2147 2759
rect 2151 2755 2152 2759
rect 2146 2754 2152 2755
rect 2162 2759 2168 2760
rect 2162 2755 2163 2759
rect 2167 2758 2168 2759
rect 2418 2759 2424 2760
rect 2167 2756 2241 2758
rect 2167 2755 2168 2756
rect 2162 2754 2168 2755
rect 2418 2755 2419 2759
rect 2423 2755 2424 2759
rect 2418 2754 2424 2755
rect 2554 2759 2560 2760
rect 2554 2755 2555 2759
rect 2559 2755 2560 2759
rect 2554 2754 2560 2755
rect 2682 2759 2688 2760
rect 2682 2755 2683 2759
rect 2687 2755 2688 2759
rect 2822 2759 2828 2760
rect 2822 2758 2823 2759
rect 2805 2756 2823 2758
rect 2682 2754 2688 2755
rect 2822 2755 2823 2756
rect 2827 2755 2828 2759
rect 2922 2759 2928 2760
rect 2822 2754 2828 2755
rect 2914 2755 2920 2756
rect 2046 2751 2052 2752
rect 199 2747 208 2748
rect 199 2743 200 2747
rect 207 2743 208 2747
rect 199 2742 208 2743
rect 210 2747 216 2748
rect 210 2743 211 2747
rect 215 2746 216 2747
rect 319 2747 325 2748
rect 319 2746 320 2747
rect 215 2744 320 2746
rect 215 2743 216 2744
rect 210 2742 216 2743
rect 319 2743 320 2744
rect 324 2743 325 2747
rect 319 2742 325 2743
rect 330 2747 336 2748
rect 330 2743 331 2747
rect 335 2746 336 2747
rect 471 2747 477 2748
rect 471 2746 472 2747
rect 335 2744 472 2746
rect 335 2743 336 2744
rect 330 2742 336 2743
rect 471 2743 472 2744
rect 476 2743 477 2747
rect 471 2742 477 2743
rect 639 2747 645 2748
rect 639 2743 640 2747
rect 644 2746 645 2747
rect 663 2747 669 2748
rect 663 2746 664 2747
rect 644 2744 664 2746
rect 644 2743 645 2744
rect 639 2742 645 2743
rect 663 2743 664 2744
rect 668 2743 669 2747
rect 663 2742 669 2743
rect 807 2747 813 2748
rect 807 2743 808 2747
rect 812 2746 813 2747
rect 826 2747 832 2748
rect 826 2746 827 2747
rect 812 2744 827 2746
rect 812 2743 813 2744
rect 807 2742 813 2743
rect 826 2743 827 2744
rect 831 2743 832 2747
rect 826 2742 832 2743
rect 983 2747 989 2748
rect 983 2743 984 2747
rect 988 2746 989 2747
rect 1018 2747 1024 2748
rect 1018 2746 1019 2747
rect 988 2744 1019 2746
rect 988 2743 989 2744
rect 983 2742 989 2743
rect 1018 2743 1019 2744
rect 1023 2743 1024 2747
rect 1018 2742 1024 2743
rect 1054 2747 1060 2748
rect 1054 2743 1055 2747
rect 1059 2746 1060 2747
rect 1151 2747 1157 2748
rect 1151 2746 1152 2747
rect 1059 2744 1152 2746
rect 1059 2743 1060 2744
rect 1054 2742 1060 2743
rect 1151 2743 1152 2744
rect 1156 2743 1157 2747
rect 1151 2742 1157 2743
rect 1319 2747 1325 2748
rect 1319 2743 1320 2747
rect 1324 2746 1325 2747
rect 1338 2747 1344 2748
rect 1338 2746 1339 2747
rect 1324 2744 1339 2746
rect 1324 2743 1325 2744
rect 1319 2742 1325 2743
rect 1338 2743 1339 2744
rect 1343 2743 1344 2747
rect 1338 2742 1344 2743
rect 1487 2747 1493 2748
rect 1487 2743 1488 2747
rect 1492 2746 1493 2747
rect 1511 2747 1517 2748
rect 1511 2746 1512 2747
rect 1492 2744 1512 2746
rect 1492 2743 1493 2744
rect 1487 2742 1493 2743
rect 1511 2743 1512 2744
rect 1516 2743 1517 2747
rect 1511 2742 1517 2743
rect 1650 2747 1656 2748
rect 1650 2743 1651 2747
rect 1655 2746 1656 2747
rect 1663 2747 1669 2748
rect 1663 2746 1664 2747
rect 1655 2744 1664 2746
rect 1655 2743 1656 2744
rect 1650 2742 1656 2743
rect 1663 2743 1664 2744
rect 1668 2743 1669 2747
rect 2046 2747 2047 2751
rect 2051 2747 2052 2751
rect 2914 2751 2915 2755
rect 2919 2751 2920 2755
rect 2922 2755 2923 2759
rect 2927 2758 2928 2759
rect 3039 2759 3045 2760
rect 2927 2756 2985 2758
rect 2927 2755 2928 2756
rect 2922 2754 2928 2755
rect 3039 2755 3040 2759
rect 3044 2758 3045 2759
rect 3130 2759 3136 2760
rect 3044 2756 3089 2758
rect 3044 2755 3045 2756
rect 3039 2754 3045 2755
rect 3130 2755 3131 2759
rect 3135 2758 3136 2759
rect 3231 2759 3237 2760
rect 3135 2756 3185 2758
rect 3135 2755 3136 2756
rect 3130 2754 3136 2755
rect 3231 2755 3232 2759
rect 3236 2758 3237 2759
rect 3418 2759 3424 2760
rect 3236 2756 3281 2758
rect 3236 2755 3237 2756
rect 3231 2754 3237 2755
rect 3418 2755 3419 2759
rect 3423 2755 3424 2759
rect 3418 2754 3424 2755
rect 3522 2759 3528 2760
rect 3522 2755 3523 2759
rect 3527 2755 3528 2759
rect 3522 2754 3528 2755
rect 3530 2759 3536 2760
rect 3530 2755 3531 2759
rect 3535 2758 3536 2759
rect 3639 2759 3645 2760
rect 3535 2756 3593 2758
rect 3535 2755 3536 2756
rect 3530 2754 3536 2755
rect 3639 2755 3640 2759
rect 3644 2758 3645 2759
rect 3818 2759 3824 2760
rect 3644 2756 3689 2758
rect 3644 2755 3645 2756
rect 3639 2754 3645 2755
rect 3818 2755 3819 2759
rect 3823 2755 3824 2759
rect 3818 2754 3824 2755
rect 3826 2759 3832 2760
rect 3826 2755 3827 2759
rect 3831 2758 3832 2759
rect 3831 2756 3881 2758
rect 3831 2755 3832 2756
rect 3826 2754 3832 2755
rect 2914 2750 2920 2751
rect 3942 2751 3948 2752
rect 2046 2746 2052 2747
rect 2070 2748 2076 2749
rect 2070 2744 2071 2748
rect 2075 2744 2076 2748
rect 2070 2743 2076 2744
rect 2198 2748 2204 2749
rect 2198 2744 2199 2748
rect 2203 2744 2204 2748
rect 2198 2743 2204 2744
rect 2342 2748 2348 2749
rect 2342 2744 2343 2748
rect 2347 2744 2348 2748
rect 2342 2743 2348 2744
rect 2478 2748 2484 2749
rect 2478 2744 2479 2748
rect 2483 2744 2484 2748
rect 2478 2743 2484 2744
rect 2606 2748 2612 2749
rect 2606 2744 2607 2748
rect 2611 2744 2612 2748
rect 2606 2743 2612 2744
rect 2726 2748 2732 2749
rect 2726 2744 2727 2748
rect 2731 2744 2732 2748
rect 2726 2743 2732 2744
rect 2838 2748 2844 2749
rect 2838 2744 2839 2748
rect 2843 2744 2844 2748
rect 2838 2743 2844 2744
rect 2942 2748 2948 2749
rect 2942 2744 2943 2748
rect 2947 2744 2948 2748
rect 2942 2743 2948 2744
rect 3046 2748 3052 2749
rect 3046 2744 3047 2748
rect 3051 2744 3052 2748
rect 3046 2743 3052 2744
rect 3142 2748 3148 2749
rect 3142 2744 3143 2748
rect 3147 2744 3148 2748
rect 3142 2743 3148 2744
rect 3238 2748 3244 2749
rect 3238 2744 3239 2748
rect 3243 2744 3244 2748
rect 3238 2743 3244 2744
rect 3342 2748 3348 2749
rect 3342 2744 3343 2748
rect 3347 2744 3348 2748
rect 3342 2743 3348 2744
rect 3446 2748 3452 2749
rect 3446 2744 3447 2748
rect 3451 2744 3452 2748
rect 3446 2743 3452 2744
rect 3550 2748 3556 2749
rect 3550 2744 3551 2748
rect 3555 2744 3556 2748
rect 3550 2743 3556 2744
rect 3646 2748 3652 2749
rect 3646 2744 3647 2748
rect 3651 2744 3652 2748
rect 3646 2743 3652 2744
rect 3742 2748 3748 2749
rect 3742 2744 3743 2748
rect 3747 2744 3748 2748
rect 3742 2743 3748 2744
rect 3838 2748 3844 2749
rect 3838 2744 3839 2748
rect 3843 2744 3844 2748
rect 3942 2747 3943 2751
rect 3947 2747 3948 2751
rect 3942 2746 3948 2747
rect 3838 2743 3844 2744
rect 1663 2742 1669 2743
rect 110 2728 116 2729
rect 2006 2728 2012 2729
rect 110 2724 111 2728
rect 115 2724 116 2728
rect 110 2723 116 2724
rect 134 2727 140 2728
rect 134 2723 135 2727
rect 139 2723 140 2727
rect 134 2722 140 2723
rect 254 2727 260 2728
rect 254 2723 255 2727
rect 259 2723 260 2727
rect 254 2722 260 2723
rect 406 2727 412 2728
rect 406 2723 407 2727
rect 411 2723 412 2727
rect 406 2722 412 2723
rect 574 2727 580 2728
rect 574 2723 575 2727
rect 579 2723 580 2727
rect 574 2722 580 2723
rect 742 2727 748 2728
rect 742 2723 743 2727
rect 747 2723 748 2727
rect 742 2722 748 2723
rect 918 2727 924 2728
rect 918 2723 919 2727
rect 923 2723 924 2727
rect 918 2722 924 2723
rect 1086 2727 1092 2728
rect 1086 2723 1087 2727
rect 1091 2723 1092 2727
rect 1086 2722 1092 2723
rect 1254 2727 1260 2728
rect 1254 2723 1255 2727
rect 1259 2723 1260 2727
rect 1254 2722 1260 2723
rect 1422 2727 1428 2728
rect 1422 2723 1423 2727
rect 1427 2723 1428 2727
rect 1422 2722 1428 2723
rect 1598 2727 1604 2728
rect 1598 2723 1599 2727
rect 1603 2723 1604 2727
rect 2006 2724 2007 2728
rect 2011 2724 2012 2728
rect 2006 2723 2012 2724
rect 1598 2722 1604 2723
rect 210 2719 216 2720
rect 210 2715 211 2719
rect 215 2715 216 2719
rect 210 2714 216 2715
rect 330 2719 336 2720
rect 330 2715 331 2719
rect 335 2715 336 2719
rect 330 2714 336 2715
rect 342 2719 348 2720
rect 342 2715 343 2719
rect 347 2718 348 2719
rect 650 2719 656 2720
rect 347 2716 449 2718
rect 347 2715 348 2716
rect 342 2714 348 2715
rect 650 2715 651 2719
rect 655 2715 656 2719
rect 650 2714 656 2715
rect 663 2719 669 2720
rect 663 2715 664 2719
rect 668 2718 669 2719
rect 1054 2719 1060 2720
rect 1054 2718 1055 2719
rect 668 2716 785 2718
rect 997 2716 1055 2718
rect 668 2715 669 2716
rect 663 2714 669 2715
rect 1054 2715 1055 2716
rect 1059 2715 1060 2719
rect 1054 2714 1060 2715
rect 1162 2719 1168 2720
rect 1162 2715 1163 2719
rect 1167 2715 1168 2719
rect 1162 2714 1168 2715
rect 1338 2719 1344 2720
rect 1338 2715 1339 2719
rect 1343 2718 1344 2719
rect 1511 2719 1517 2720
rect 1343 2716 1465 2718
rect 1343 2715 1344 2716
rect 1338 2714 1344 2715
rect 1511 2715 1512 2719
rect 1516 2718 1517 2719
rect 1516 2716 1641 2718
rect 1516 2715 1517 2716
rect 1511 2714 1517 2715
rect 110 2711 116 2712
rect 110 2707 111 2711
rect 115 2707 116 2711
rect 1332 2710 1334 2713
rect 1342 2711 1348 2712
rect 1342 2710 1343 2711
rect 110 2706 116 2707
rect 134 2708 140 2709
rect 134 2704 135 2708
rect 139 2704 140 2708
rect 134 2703 140 2704
rect 254 2708 260 2709
rect 254 2704 255 2708
rect 259 2704 260 2708
rect 254 2703 260 2704
rect 406 2708 412 2709
rect 406 2704 407 2708
rect 411 2704 412 2708
rect 406 2703 412 2704
rect 574 2708 580 2709
rect 574 2704 575 2708
rect 579 2704 580 2708
rect 574 2703 580 2704
rect 742 2708 748 2709
rect 742 2704 743 2708
rect 747 2704 748 2708
rect 742 2703 748 2704
rect 918 2708 924 2709
rect 918 2704 919 2708
rect 923 2704 924 2708
rect 918 2703 924 2704
rect 1086 2708 1092 2709
rect 1086 2704 1087 2708
rect 1091 2704 1092 2708
rect 1086 2703 1092 2704
rect 1254 2708 1260 2709
rect 1332 2708 1343 2710
rect 1254 2704 1255 2708
rect 1259 2704 1260 2708
rect 1342 2707 1343 2708
rect 1347 2707 1348 2711
rect 2006 2711 2012 2712
rect 1342 2706 1348 2707
rect 1422 2708 1428 2709
rect 1254 2703 1260 2704
rect 1422 2704 1423 2708
rect 1427 2704 1428 2708
rect 1422 2703 1428 2704
rect 1598 2708 1604 2709
rect 1598 2704 1599 2708
rect 1603 2704 1604 2708
rect 2006 2707 2007 2711
rect 2011 2707 2012 2711
rect 2006 2706 2012 2707
rect 1598 2703 1604 2704
rect 2094 2668 2100 2669
rect 2046 2665 2052 2666
rect 2046 2661 2047 2665
rect 2051 2661 2052 2665
rect 2094 2664 2095 2668
rect 2099 2664 2100 2668
rect 2094 2663 2100 2664
rect 2262 2668 2268 2669
rect 2262 2664 2263 2668
rect 2267 2664 2268 2668
rect 2262 2663 2268 2664
rect 2438 2668 2444 2669
rect 2438 2664 2439 2668
rect 2443 2664 2444 2668
rect 2438 2663 2444 2664
rect 2614 2668 2620 2669
rect 2614 2664 2615 2668
rect 2619 2664 2620 2668
rect 2614 2663 2620 2664
rect 2782 2668 2788 2669
rect 2782 2664 2783 2668
rect 2787 2664 2788 2668
rect 2782 2663 2788 2664
rect 2942 2668 2948 2669
rect 2942 2664 2943 2668
rect 2947 2664 2948 2668
rect 2942 2663 2948 2664
rect 3094 2668 3100 2669
rect 3094 2664 3095 2668
rect 3099 2664 3100 2668
rect 3094 2663 3100 2664
rect 3238 2668 3244 2669
rect 3238 2664 3239 2668
rect 3243 2664 3244 2668
rect 3238 2663 3244 2664
rect 3382 2668 3388 2669
rect 3382 2664 3383 2668
rect 3387 2664 3388 2668
rect 3382 2663 3388 2664
rect 3534 2668 3540 2669
rect 3534 2664 3535 2668
rect 3539 2664 3540 2668
rect 3534 2663 3540 2664
rect 3942 2665 3948 2666
rect 2046 2660 2052 2661
rect 3942 2661 3943 2665
rect 3947 2661 3948 2665
rect 3942 2660 3948 2661
rect 2170 2659 2176 2660
rect 2170 2655 2171 2659
rect 2175 2655 2176 2659
rect 2170 2654 2176 2655
rect 2330 2659 2336 2660
rect 2330 2655 2331 2659
rect 2335 2655 2336 2659
rect 2330 2654 2336 2655
rect 2410 2659 2416 2660
rect 2410 2655 2411 2659
rect 2415 2658 2416 2659
rect 2522 2659 2528 2660
rect 2415 2656 2481 2658
rect 2415 2655 2416 2656
rect 2410 2654 2416 2655
rect 2522 2655 2523 2659
rect 2527 2658 2528 2659
rect 2719 2659 2725 2660
rect 2527 2656 2657 2658
rect 2527 2655 2528 2656
rect 2522 2654 2528 2655
rect 2719 2655 2720 2659
rect 2724 2658 2725 2659
rect 3018 2659 3024 2660
rect 2724 2656 2825 2658
rect 2724 2655 2725 2656
rect 2719 2654 2725 2655
rect 3018 2655 3019 2659
rect 3023 2655 3024 2659
rect 3018 2654 3024 2655
rect 3170 2659 3176 2660
rect 3170 2655 3171 2659
rect 3175 2655 3176 2659
rect 3170 2654 3176 2655
rect 3314 2659 3320 2660
rect 3314 2655 3315 2659
rect 3319 2655 3320 2659
rect 3314 2654 3320 2655
rect 3458 2659 3464 2660
rect 3458 2655 3459 2659
rect 3463 2655 3464 2659
rect 3458 2654 3464 2655
rect 3466 2659 3472 2660
rect 3466 2655 3467 2659
rect 3471 2658 3472 2659
rect 3471 2656 3577 2658
rect 3471 2655 3472 2656
rect 3466 2654 3472 2655
rect 2094 2649 2100 2650
rect 166 2648 172 2649
rect 110 2645 116 2646
rect 110 2641 111 2645
rect 115 2641 116 2645
rect 166 2644 167 2648
rect 171 2644 172 2648
rect 166 2643 172 2644
rect 358 2648 364 2649
rect 358 2644 359 2648
rect 363 2644 364 2648
rect 358 2643 364 2644
rect 558 2648 564 2649
rect 558 2644 559 2648
rect 563 2644 564 2648
rect 558 2643 564 2644
rect 758 2648 764 2649
rect 758 2644 759 2648
rect 763 2644 764 2648
rect 758 2643 764 2644
rect 950 2648 956 2649
rect 950 2644 951 2648
rect 955 2644 956 2648
rect 950 2643 956 2644
rect 1142 2648 1148 2649
rect 1142 2644 1143 2648
rect 1147 2644 1148 2648
rect 1142 2643 1148 2644
rect 1326 2648 1332 2649
rect 1326 2644 1327 2648
rect 1331 2644 1332 2648
rect 1326 2643 1332 2644
rect 1510 2648 1516 2649
rect 1510 2644 1511 2648
rect 1515 2644 1516 2648
rect 1510 2643 1516 2644
rect 1702 2648 1708 2649
rect 1702 2644 1703 2648
rect 1707 2644 1708 2648
rect 2046 2648 2052 2649
rect 1702 2643 1708 2644
rect 2006 2645 2012 2646
rect 110 2640 116 2641
rect 2006 2641 2007 2645
rect 2011 2641 2012 2645
rect 2046 2644 2047 2648
rect 2051 2644 2052 2648
rect 2094 2645 2095 2649
rect 2099 2645 2100 2649
rect 2094 2644 2100 2645
rect 2262 2649 2268 2650
rect 2262 2645 2263 2649
rect 2267 2645 2268 2649
rect 2262 2644 2268 2645
rect 2438 2649 2444 2650
rect 2438 2645 2439 2649
rect 2443 2645 2444 2649
rect 2438 2644 2444 2645
rect 2614 2649 2620 2650
rect 2614 2645 2615 2649
rect 2619 2645 2620 2649
rect 2614 2644 2620 2645
rect 2782 2649 2788 2650
rect 2782 2645 2783 2649
rect 2787 2645 2788 2649
rect 2782 2644 2788 2645
rect 2942 2649 2948 2650
rect 2942 2645 2943 2649
rect 2947 2645 2948 2649
rect 2942 2644 2948 2645
rect 3094 2649 3100 2650
rect 3094 2645 3095 2649
rect 3099 2645 3100 2649
rect 3094 2644 3100 2645
rect 3238 2649 3244 2650
rect 3238 2645 3239 2649
rect 3243 2645 3244 2649
rect 3238 2644 3244 2645
rect 3382 2649 3388 2650
rect 3382 2645 3383 2649
rect 3387 2645 3388 2649
rect 3382 2644 3388 2645
rect 3534 2649 3540 2650
rect 3534 2645 3535 2649
rect 3539 2645 3540 2649
rect 3534 2644 3540 2645
rect 3942 2648 3948 2649
rect 3942 2644 3943 2648
rect 3947 2644 3948 2648
rect 2046 2643 2052 2644
rect 3942 2643 3948 2644
rect 2006 2640 2012 2641
rect 282 2639 288 2640
rect 282 2638 283 2639
rect 245 2636 283 2638
rect 282 2635 283 2636
rect 287 2635 288 2639
rect 282 2634 288 2635
rect 434 2639 440 2640
rect 434 2635 435 2639
rect 439 2635 440 2639
rect 434 2634 440 2635
rect 634 2639 640 2640
rect 634 2635 635 2639
rect 639 2635 640 2639
rect 634 2634 640 2635
rect 826 2639 832 2640
rect 826 2635 827 2639
rect 831 2635 832 2639
rect 826 2634 832 2635
rect 1018 2639 1024 2640
rect 1018 2635 1019 2639
rect 1023 2635 1024 2639
rect 1018 2634 1024 2635
rect 1034 2639 1040 2640
rect 1034 2635 1035 2639
rect 1039 2638 1040 2639
rect 1402 2639 1408 2640
rect 1039 2636 1185 2638
rect 1039 2635 1040 2636
rect 1034 2634 1040 2635
rect 1402 2635 1403 2639
rect 1407 2635 1408 2639
rect 1402 2634 1408 2635
rect 1586 2639 1592 2640
rect 1586 2635 1587 2639
rect 1591 2635 1592 2639
rect 1586 2634 1592 2635
rect 1778 2639 1784 2640
rect 1778 2635 1779 2639
rect 1783 2635 1784 2639
rect 1778 2634 1784 2635
rect 166 2629 172 2630
rect 110 2628 116 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 166 2625 167 2629
rect 171 2625 172 2629
rect 166 2624 172 2625
rect 358 2629 364 2630
rect 358 2625 359 2629
rect 363 2625 364 2629
rect 358 2624 364 2625
rect 558 2629 564 2630
rect 558 2625 559 2629
rect 563 2625 564 2629
rect 558 2624 564 2625
rect 758 2629 764 2630
rect 758 2625 759 2629
rect 763 2625 764 2629
rect 758 2624 764 2625
rect 950 2629 956 2630
rect 950 2625 951 2629
rect 955 2625 956 2629
rect 950 2624 956 2625
rect 1142 2629 1148 2630
rect 1142 2625 1143 2629
rect 1147 2625 1148 2629
rect 1142 2624 1148 2625
rect 1326 2629 1332 2630
rect 1326 2625 1327 2629
rect 1331 2625 1332 2629
rect 1326 2624 1332 2625
rect 1510 2629 1516 2630
rect 1510 2625 1511 2629
rect 1515 2625 1516 2629
rect 1510 2624 1516 2625
rect 1702 2629 1708 2630
rect 1702 2625 1703 2629
rect 1707 2625 1708 2629
rect 1702 2624 1708 2625
rect 2006 2628 2012 2629
rect 2006 2624 2007 2628
rect 2011 2624 2012 2628
rect 110 2623 116 2624
rect 2006 2623 2012 2624
rect 2159 2627 2168 2628
rect 2159 2623 2160 2627
rect 2167 2623 2168 2627
rect 2159 2622 2168 2623
rect 2170 2627 2176 2628
rect 2170 2623 2171 2627
rect 2175 2626 2176 2627
rect 2327 2627 2333 2628
rect 2327 2626 2328 2627
rect 2175 2624 2328 2626
rect 2175 2623 2176 2624
rect 2170 2622 2176 2623
rect 2327 2623 2328 2624
rect 2332 2623 2333 2627
rect 2327 2622 2333 2623
rect 2503 2627 2509 2628
rect 2503 2623 2504 2627
rect 2508 2626 2509 2627
rect 2522 2627 2528 2628
rect 2522 2626 2523 2627
rect 2508 2624 2523 2626
rect 2508 2623 2509 2624
rect 2503 2622 2509 2623
rect 2522 2623 2523 2624
rect 2527 2623 2528 2627
rect 2522 2622 2528 2623
rect 2679 2627 2685 2628
rect 2679 2623 2680 2627
rect 2684 2626 2685 2627
rect 2719 2627 2725 2628
rect 2719 2626 2720 2627
rect 2684 2624 2720 2626
rect 2684 2623 2685 2624
rect 2679 2622 2685 2623
rect 2719 2623 2720 2624
rect 2724 2623 2725 2627
rect 2719 2622 2725 2623
rect 2746 2627 2752 2628
rect 2746 2623 2747 2627
rect 2751 2626 2752 2627
rect 2847 2627 2853 2628
rect 2847 2626 2848 2627
rect 2751 2624 2848 2626
rect 2751 2623 2752 2624
rect 2746 2622 2752 2623
rect 2847 2623 2848 2624
rect 2852 2623 2853 2627
rect 2847 2622 2853 2623
rect 2914 2627 2920 2628
rect 2914 2623 2915 2627
rect 2919 2626 2920 2627
rect 3007 2627 3013 2628
rect 3007 2626 3008 2627
rect 2919 2624 3008 2626
rect 2919 2623 2920 2624
rect 2914 2622 2920 2623
rect 3007 2623 3008 2624
rect 3012 2623 3013 2627
rect 3007 2622 3013 2623
rect 3018 2627 3024 2628
rect 3018 2623 3019 2627
rect 3023 2626 3024 2627
rect 3159 2627 3165 2628
rect 3159 2626 3160 2627
rect 3023 2624 3160 2626
rect 3023 2623 3024 2624
rect 3018 2622 3024 2623
rect 3159 2623 3160 2624
rect 3164 2623 3165 2627
rect 3159 2622 3165 2623
rect 3170 2627 3176 2628
rect 3170 2623 3171 2627
rect 3175 2626 3176 2627
rect 3303 2627 3309 2628
rect 3303 2626 3304 2627
rect 3175 2624 3304 2626
rect 3175 2623 3176 2624
rect 3170 2622 3176 2623
rect 3303 2623 3304 2624
rect 3308 2623 3309 2627
rect 3303 2622 3309 2623
rect 3314 2627 3320 2628
rect 3314 2623 3315 2627
rect 3319 2626 3320 2627
rect 3447 2627 3453 2628
rect 3447 2626 3448 2627
rect 3319 2624 3448 2626
rect 3319 2623 3320 2624
rect 3314 2622 3320 2623
rect 3447 2623 3448 2624
rect 3452 2623 3453 2627
rect 3447 2622 3453 2623
rect 3458 2627 3464 2628
rect 3458 2623 3459 2627
rect 3463 2626 3464 2627
rect 3599 2627 3605 2628
rect 3599 2626 3600 2627
rect 3463 2624 3600 2626
rect 3463 2623 3464 2624
rect 3458 2622 3464 2623
rect 3599 2623 3600 2624
rect 3604 2623 3605 2627
rect 3599 2622 3605 2623
rect 342 2615 348 2616
rect 342 2614 343 2615
rect 319 2612 343 2614
rect 319 2610 321 2612
rect 342 2611 343 2612
rect 347 2611 348 2615
rect 342 2610 348 2611
rect 276 2608 321 2610
rect 231 2607 237 2608
rect 231 2603 232 2607
rect 236 2606 237 2607
rect 276 2606 278 2608
rect 423 2607 429 2608
rect 423 2606 424 2607
rect 236 2604 278 2606
rect 319 2604 424 2606
rect 236 2603 237 2604
rect 231 2602 237 2603
rect 282 2603 288 2604
rect 282 2599 283 2603
rect 287 2602 288 2603
rect 319 2602 321 2604
rect 423 2603 424 2604
rect 428 2603 429 2607
rect 423 2602 429 2603
rect 434 2607 440 2608
rect 434 2603 435 2607
rect 439 2606 440 2607
rect 623 2607 629 2608
rect 623 2606 624 2607
rect 439 2604 624 2606
rect 439 2603 440 2604
rect 434 2602 440 2603
rect 623 2603 624 2604
rect 628 2603 629 2607
rect 623 2602 629 2603
rect 634 2607 640 2608
rect 634 2603 635 2607
rect 639 2606 640 2607
rect 823 2607 829 2608
rect 823 2606 824 2607
rect 639 2604 824 2606
rect 639 2603 640 2604
rect 634 2602 640 2603
rect 823 2603 824 2604
rect 828 2603 829 2607
rect 823 2602 829 2603
rect 1015 2607 1021 2608
rect 1015 2603 1016 2607
rect 1020 2606 1021 2607
rect 1034 2607 1040 2608
rect 1034 2606 1035 2607
rect 1020 2604 1035 2606
rect 1020 2603 1021 2604
rect 1015 2602 1021 2603
rect 1034 2603 1035 2604
rect 1039 2603 1040 2607
rect 1034 2602 1040 2603
rect 1198 2607 1204 2608
rect 1198 2603 1199 2607
rect 1203 2606 1204 2607
rect 1207 2607 1213 2608
rect 1207 2606 1208 2607
rect 1203 2604 1208 2606
rect 1203 2603 1204 2604
rect 1198 2602 1204 2603
rect 1207 2603 1208 2604
rect 1212 2603 1213 2607
rect 1207 2602 1213 2603
rect 1342 2607 1348 2608
rect 1342 2603 1343 2607
rect 1347 2606 1348 2607
rect 1391 2607 1397 2608
rect 1391 2606 1392 2607
rect 1347 2604 1392 2606
rect 1347 2603 1348 2604
rect 1342 2602 1348 2603
rect 1391 2603 1392 2604
rect 1396 2603 1397 2607
rect 1391 2602 1397 2603
rect 1402 2607 1408 2608
rect 1402 2603 1403 2607
rect 1407 2606 1408 2607
rect 1575 2607 1581 2608
rect 1575 2606 1576 2607
rect 1407 2604 1576 2606
rect 1407 2603 1408 2604
rect 1402 2602 1408 2603
rect 1575 2603 1576 2604
rect 1580 2603 1581 2607
rect 1575 2602 1581 2603
rect 1586 2607 1592 2608
rect 1586 2603 1587 2607
rect 1591 2606 1592 2607
rect 1767 2607 1773 2608
rect 1767 2606 1768 2607
rect 1591 2604 1768 2606
rect 1591 2603 1592 2604
rect 1586 2602 1592 2603
rect 1767 2603 1768 2604
rect 1772 2603 1773 2607
rect 1767 2602 1773 2603
rect 2279 2607 2285 2608
rect 2279 2603 2280 2607
rect 2284 2606 2285 2607
rect 2330 2607 2336 2608
rect 2330 2606 2331 2607
rect 2284 2604 2331 2606
rect 2284 2603 2285 2604
rect 2279 2602 2285 2603
rect 2330 2603 2331 2604
rect 2335 2603 2336 2607
rect 2330 2602 2336 2603
rect 2418 2607 2424 2608
rect 2418 2603 2419 2607
rect 2423 2606 2424 2607
rect 2431 2607 2437 2608
rect 2431 2606 2432 2607
rect 2423 2604 2432 2606
rect 2423 2603 2424 2604
rect 2418 2602 2424 2603
rect 2431 2603 2432 2604
rect 2436 2603 2437 2607
rect 2431 2602 2437 2603
rect 2494 2607 2500 2608
rect 2494 2603 2495 2607
rect 2499 2606 2500 2607
rect 2583 2607 2589 2608
rect 2583 2606 2584 2607
rect 2499 2604 2584 2606
rect 2499 2603 2500 2604
rect 2494 2602 2500 2603
rect 2583 2603 2584 2604
rect 2588 2603 2589 2607
rect 2583 2602 2589 2603
rect 2594 2607 2600 2608
rect 2594 2603 2595 2607
rect 2599 2606 2600 2607
rect 2735 2607 2741 2608
rect 2735 2606 2736 2607
rect 2599 2604 2736 2606
rect 2599 2603 2600 2604
rect 2594 2602 2600 2603
rect 2735 2603 2736 2604
rect 2740 2603 2741 2607
rect 2735 2602 2741 2603
rect 2879 2607 2885 2608
rect 2879 2603 2880 2607
rect 2884 2606 2885 2607
rect 2903 2607 2909 2608
rect 2903 2606 2904 2607
rect 2884 2604 2904 2606
rect 2884 2603 2885 2604
rect 2879 2602 2885 2603
rect 2903 2603 2904 2604
rect 2908 2603 2909 2607
rect 2903 2602 2909 2603
rect 3015 2607 3021 2608
rect 3015 2603 3016 2607
rect 3020 2606 3021 2607
rect 3034 2607 3040 2608
rect 3034 2606 3035 2607
rect 3020 2604 3035 2606
rect 3020 2603 3021 2604
rect 3015 2602 3021 2603
rect 3034 2603 3035 2604
rect 3039 2603 3040 2607
rect 3034 2602 3040 2603
rect 3151 2607 3157 2608
rect 3151 2603 3152 2607
rect 3156 2606 3157 2607
rect 3170 2607 3176 2608
rect 3170 2606 3171 2607
rect 3156 2604 3171 2606
rect 3156 2603 3157 2604
rect 3151 2602 3157 2603
rect 3170 2603 3171 2604
rect 3175 2603 3176 2607
rect 3170 2602 3176 2603
rect 3287 2607 3293 2608
rect 3287 2603 3288 2607
rect 3292 2606 3293 2607
rect 3306 2607 3312 2608
rect 3306 2606 3307 2607
rect 3292 2604 3307 2606
rect 3292 2603 3293 2604
rect 3287 2602 3293 2603
rect 3306 2603 3307 2604
rect 3311 2603 3312 2607
rect 3306 2602 3312 2603
rect 3431 2607 3437 2608
rect 3431 2603 3432 2607
rect 3436 2606 3437 2607
rect 3466 2607 3472 2608
rect 3466 2606 3467 2607
rect 3436 2604 3467 2606
rect 3436 2603 3437 2604
rect 3431 2602 3437 2603
rect 3466 2603 3467 2604
rect 3471 2603 3472 2607
rect 3466 2602 3472 2603
rect 287 2600 321 2602
rect 287 2599 288 2600
rect 282 2598 288 2599
rect 2046 2588 2052 2589
rect 3942 2588 3948 2589
rect 2046 2584 2047 2588
rect 2051 2584 2052 2588
rect 2046 2583 2052 2584
rect 2214 2587 2220 2588
rect 2214 2583 2215 2587
rect 2219 2583 2220 2587
rect 2214 2582 2220 2583
rect 2366 2587 2372 2588
rect 2366 2583 2367 2587
rect 2371 2583 2372 2587
rect 2366 2582 2372 2583
rect 2518 2587 2524 2588
rect 2518 2583 2519 2587
rect 2523 2583 2524 2587
rect 2518 2582 2524 2583
rect 2670 2587 2676 2588
rect 2670 2583 2671 2587
rect 2675 2583 2676 2587
rect 2670 2582 2676 2583
rect 2814 2587 2820 2588
rect 2814 2583 2815 2587
rect 2819 2583 2820 2587
rect 2814 2582 2820 2583
rect 2950 2587 2956 2588
rect 2950 2583 2951 2587
rect 2955 2583 2956 2587
rect 2950 2582 2956 2583
rect 3086 2587 3092 2588
rect 3086 2583 3087 2587
rect 3091 2583 3092 2587
rect 3086 2582 3092 2583
rect 3222 2587 3228 2588
rect 3222 2583 3223 2587
rect 3227 2583 3228 2587
rect 3222 2582 3228 2583
rect 3366 2587 3372 2588
rect 3366 2583 3367 2587
rect 3371 2583 3372 2587
rect 3942 2584 3943 2588
rect 3947 2584 3948 2588
rect 3942 2583 3948 2584
rect 3366 2582 3372 2583
rect 639 2579 645 2580
rect 639 2575 640 2579
rect 644 2578 645 2579
rect 650 2579 656 2580
rect 644 2575 646 2578
rect 639 2574 646 2575
rect 650 2575 651 2579
rect 655 2578 656 2579
rect 751 2579 757 2580
rect 751 2578 752 2579
rect 655 2576 752 2578
rect 655 2575 656 2576
rect 650 2574 656 2575
rect 751 2575 752 2576
rect 756 2575 757 2579
rect 751 2574 757 2575
rect 782 2579 788 2580
rect 782 2575 783 2579
rect 787 2578 788 2579
rect 871 2579 877 2580
rect 871 2578 872 2579
rect 787 2576 872 2578
rect 787 2575 788 2576
rect 782 2574 788 2575
rect 871 2575 872 2576
rect 876 2575 877 2579
rect 871 2574 877 2575
rect 882 2579 888 2580
rect 882 2575 883 2579
rect 887 2578 888 2579
rect 999 2579 1005 2580
rect 999 2578 1000 2579
rect 887 2576 1000 2578
rect 887 2575 888 2576
rect 882 2574 888 2575
rect 999 2575 1000 2576
rect 1004 2575 1005 2579
rect 999 2574 1005 2575
rect 1010 2579 1016 2580
rect 1010 2575 1011 2579
rect 1015 2578 1016 2579
rect 1135 2579 1141 2580
rect 1135 2578 1136 2579
rect 1015 2576 1136 2578
rect 1015 2575 1016 2576
rect 1010 2574 1016 2575
rect 1135 2575 1136 2576
rect 1140 2575 1141 2579
rect 1135 2574 1141 2575
rect 1271 2579 1277 2580
rect 1271 2575 1272 2579
rect 1276 2578 1277 2579
rect 1295 2579 1301 2580
rect 1295 2578 1296 2579
rect 1276 2576 1296 2578
rect 1276 2575 1277 2576
rect 1271 2574 1277 2575
rect 1295 2575 1296 2576
rect 1300 2575 1301 2579
rect 1295 2574 1301 2575
rect 1358 2579 1364 2580
rect 1358 2575 1359 2579
rect 1363 2578 1364 2579
rect 1415 2579 1421 2580
rect 1415 2578 1416 2579
rect 1363 2576 1416 2578
rect 1363 2575 1364 2576
rect 1358 2574 1364 2575
rect 1415 2575 1416 2576
rect 1420 2575 1421 2579
rect 1415 2574 1421 2575
rect 1559 2579 1565 2580
rect 1559 2575 1560 2579
rect 1564 2578 1565 2579
rect 1578 2579 1584 2580
rect 1578 2578 1579 2579
rect 1564 2576 1579 2578
rect 1564 2575 1565 2576
rect 1559 2574 1565 2575
rect 1578 2575 1579 2576
rect 1583 2575 1584 2579
rect 1578 2574 1584 2575
rect 1711 2579 1717 2580
rect 1711 2575 1712 2579
rect 1716 2578 1717 2579
rect 1730 2579 1736 2580
rect 1730 2578 1731 2579
rect 1716 2576 1731 2578
rect 1716 2575 1717 2576
rect 1711 2574 1717 2575
rect 1730 2575 1731 2576
rect 1735 2575 1736 2579
rect 1730 2574 1736 2575
rect 1778 2579 1784 2580
rect 1778 2575 1779 2579
rect 1783 2578 1784 2579
rect 1863 2579 1869 2580
rect 1863 2578 1864 2579
rect 1783 2576 1864 2578
rect 1783 2575 1784 2576
rect 1778 2574 1784 2575
rect 1863 2575 1864 2576
rect 1868 2575 1869 2579
rect 2494 2579 2500 2580
rect 2494 2578 2495 2579
rect 2445 2576 2495 2578
rect 1863 2574 1869 2575
rect 2358 2575 2364 2576
rect 2358 2574 2359 2575
rect 644 2570 646 2574
rect 2293 2572 2359 2574
rect 702 2571 708 2572
rect 702 2570 703 2571
rect 644 2568 703 2570
rect 702 2567 703 2568
rect 707 2567 708 2571
rect 702 2566 708 2567
rect 2046 2571 2052 2572
rect 2046 2567 2047 2571
rect 2051 2567 2052 2571
rect 2358 2571 2359 2572
rect 2363 2571 2364 2575
rect 2494 2575 2495 2576
rect 2499 2575 2500 2579
rect 2494 2574 2500 2575
rect 2594 2579 2600 2580
rect 2594 2575 2595 2579
rect 2599 2575 2600 2579
rect 2594 2574 2600 2575
rect 2746 2579 2752 2580
rect 2746 2575 2747 2579
rect 2751 2575 2752 2579
rect 2746 2574 2752 2575
rect 2786 2579 2792 2580
rect 2786 2575 2787 2579
rect 2791 2578 2792 2579
rect 2903 2579 2909 2580
rect 2791 2576 2857 2578
rect 2791 2575 2792 2576
rect 2786 2574 2792 2575
rect 2903 2575 2904 2579
rect 2908 2578 2909 2579
rect 3034 2579 3040 2580
rect 2908 2576 2993 2578
rect 2908 2575 2909 2576
rect 2903 2574 2909 2575
rect 3034 2575 3035 2579
rect 3039 2578 3040 2579
rect 3170 2579 3176 2580
rect 3039 2576 3129 2578
rect 3039 2575 3040 2576
rect 3034 2574 3040 2575
rect 3170 2575 3171 2579
rect 3175 2578 3176 2579
rect 3306 2579 3312 2580
rect 3175 2576 3265 2578
rect 3175 2575 3176 2576
rect 3170 2574 3176 2575
rect 3306 2575 3307 2579
rect 3311 2578 3312 2579
rect 3311 2576 3409 2578
rect 3311 2575 3312 2576
rect 3306 2574 3312 2575
rect 2358 2570 2364 2571
rect 3942 2571 3948 2572
rect 2046 2566 2052 2567
rect 2214 2568 2220 2569
rect 2214 2564 2215 2568
rect 2219 2564 2220 2568
rect 2214 2563 2220 2564
rect 2366 2568 2372 2569
rect 2366 2564 2367 2568
rect 2371 2564 2372 2568
rect 2366 2563 2372 2564
rect 2518 2568 2524 2569
rect 2518 2564 2519 2568
rect 2523 2564 2524 2568
rect 2518 2563 2524 2564
rect 2670 2568 2676 2569
rect 2670 2564 2671 2568
rect 2675 2564 2676 2568
rect 2670 2563 2676 2564
rect 2814 2568 2820 2569
rect 2814 2564 2815 2568
rect 2819 2564 2820 2568
rect 2814 2563 2820 2564
rect 2950 2568 2956 2569
rect 2950 2564 2951 2568
rect 2955 2564 2956 2568
rect 2950 2563 2956 2564
rect 3086 2568 3092 2569
rect 3086 2564 3087 2568
rect 3091 2564 3092 2568
rect 3086 2563 3092 2564
rect 3222 2568 3228 2569
rect 3222 2564 3223 2568
rect 3227 2564 3228 2568
rect 3222 2563 3228 2564
rect 3366 2568 3372 2569
rect 3366 2564 3367 2568
rect 3371 2564 3372 2568
rect 3942 2567 3943 2571
rect 3947 2567 3948 2571
rect 3942 2566 3948 2567
rect 3366 2563 3372 2564
rect 110 2560 116 2561
rect 2006 2560 2012 2561
rect 110 2556 111 2560
rect 115 2556 116 2560
rect 110 2555 116 2556
rect 574 2559 580 2560
rect 574 2555 575 2559
rect 579 2555 580 2559
rect 574 2554 580 2555
rect 686 2559 692 2560
rect 686 2555 687 2559
rect 691 2555 692 2559
rect 686 2554 692 2555
rect 806 2559 812 2560
rect 806 2555 807 2559
rect 811 2555 812 2559
rect 806 2554 812 2555
rect 934 2559 940 2560
rect 934 2555 935 2559
rect 939 2555 940 2559
rect 934 2554 940 2555
rect 1070 2559 1076 2560
rect 1070 2555 1071 2559
rect 1075 2555 1076 2559
rect 1070 2554 1076 2555
rect 1206 2559 1212 2560
rect 1206 2555 1207 2559
rect 1211 2555 1212 2559
rect 1206 2554 1212 2555
rect 1350 2559 1356 2560
rect 1350 2555 1351 2559
rect 1355 2555 1356 2559
rect 1350 2554 1356 2555
rect 1494 2559 1500 2560
rect 1494 2555 1495 2559
rect 1499 2555 1500 2559
rect 1494 2554 1500 2555
rect 1646 2559 1652 2560
rect 1646 2555 1647 2559
rect 1651 2555 1652 2559
rect 1646 2554 1652 2555
rect 1798 2559 1804 2560
rect 1798 2555 1799 2559
rect 1803 2555 1804 2559
rect 2006 2556 2007 2560
rect 2011 2556 2012 2560
rect 2006 2555 2012 2556
rect 1798 2554 1804 2555
rect 650 2551 656 2552
rect 650 2547 651 2551
rect 655 2547 656 2551
rect 782 2551 788 2552
rect 782 2550 783 2551
rect 765 2548 783 2550
rect 650 2546 656 2547
rect 782 2547 783 2548
rect 787 2547 788 2551
rect 782 2546 788 2547
rect 882 2551 888 2552
rect 882 2547 883 2551
rect 887 2547 888 2551
rect 882 2546 888 2547
rect 1010 2551 1016 2552
rect 1010 2547 1011 2551
rect 1015 2547 1016 2551
rect 1198 2551 1204 2552
rect 1010 2546 1016 2547
rect 1146 2547 1152 2548
rect 110 2543 116 2544
rect 110 2539 111 2543
rect 115 2539 116 2543
rect 1146 2543 1147 2547
rect 1151 2543 1152 2547
rect 1198 2547 1199 2551
rect 1203 2550 1204 2551
rect 1295 2551 1301 2552
rect 1203 2548 1249 2550
rect 1203 2547 1204 2548
rect 1198 2546 1204 2547
rect 1295 2547 1296 2551
rect 1300 2550 1301 2551
rect 1578 2551 1584 2552
rect 1300 2548 1393 2550
rect 1300 2547 1301 2548
rect 1295 2546 1301 2547
rect 1570 2547 1576 2548
rect 1146 2542 1152 2543
rect 1570 2543 1571 2547
rect 1575 2543 1576 2547
rect 1578 2547 1579 2551
rect 1583 2550 1584 2551
rect 1730 2551 1736 2552
rect 1583 2548 1689 2550
rect 1583 2547 1584 2548
rect 1578 2546 1584 2547
rect 1730 2547 1731 2551
rect 1735 2550 1736 2551
rect 1735 2548 1841 2550
rect 1735 2547 1736 2548
rect 1730 2546 1736 2547
rect 1570 2542 1576 2543
rect 2006 2543 2012 2544
rect 110 2538 116 2539
rect 574 2540 580 2541
rect 574 2536 575 2540
rect 579 2536 580 2540
rect 574 2535 580 2536
rect 686 2540 692 2541
rect 686 2536 687 2540
rect 691 2536 692 2540
rect 686 2535 692 2536
rect 806 2540 812 2541
rect 806 2536 807 2540
rect 811 2536 812 2540
rect 806 2535 812 2536
rect 934 2540 940 2541
rect 934 2536 935 2540
rect 939 2536 940 2540
rect 934 2535 940 2536
rect 1070 2540 1076 2541
rect 1070 2536 1071 2540
rect 1075 2536 1076 2540
rect 1070 2535 1076 2536
rect 1206 2540 1212 2541
rect 1206 2536 1207 2540
rect 1211 2536 1212 2540
rect 1206 2535 1212 2536
rect 1350 2540 1356 2541
rect 1350 2536 1351 2540
rect 1355 2536 1356 2540
rect 1350 2535 1356 2536
rect 1494 2540 1500 2541
rect 1494 2536 1495 2540
rect 1499 2536 1500 2540
rect 1494 2535 1500 2536
rect 1646 2540 1652 2541
rect 1646 2536 1647 2540
rect 1651 2536 1652 2540
rect 1646 2535 1652 2536
rect 1798 2540 1804 2541
rect 1798 2536 1799 2540
rect 1803 2536 1804 2540
rect 2006 2539 2007 2543
rect 2011 2539 2012 2543
rect 2006 2538 2012 2539
rect 1798 2535 1804 2536
rect 2094 2504 2100 2505
rect 2046 2501 2052 2502
rect 2046 2497 2047 2501
rect 2051 2497 2052 2501
rect 2094 2500 2095 2504
rect 2099 2500 2100 2504
rect 2094 2499 2100 2500
rect 2214 2504 2220 2505
rect 2214 2500 2215 2504
rect 2219 2500 2220 2504
rect 2214 2499 2220 2500
rect 2342 2504 2348 2505
rect 2342 2500 2343 2504
rect 2347 2500 2348 2504
rect 2342 2499 2348 2500
rect 2470 2504 2476 2505
rect 2470 2500 2471 2504
rect 2475 2500 2476 2504
rect 2470 2499 2476 2500
rect 2598 2504 2604 2505
rect 2598 2500 2599 2504
rect 2603 2500 2604 2504
rect 2598 2499 2604 2500
rect 2718 2504 2724 2505
rect 2718 2500 2719 2504
rect 2723 2500 2724 2504
rect 2718 2499 2724 2500
rect 2838 2504 2844 2505
rect 2838 2500 2839 2504
rect 2843 2500 2844 2504
rect 2838 2499 2844 2500
rect 2966 2504 2972 2505
rect 2966 2500 2967 2504
rect 2971 2500 2972 2504
rect 2966 2499 2972 2500
rect 3094 2504 3100 2505
rect 3094 2500 3095 2504
rect 3099 2500 3100 2504
rect 3094 2499 3100 2500
rect 3222 2504 3228 2505
rect 3222 2500 3223 2504
rect 3227 2500 3228 2504
rect 3222 2499 3228 2500
rect 3942 2501 3948 2502
rect 2046 2496 2052 2497
rect 3942 2497 3943 2501
rect 3947 2497 3948 2501
rect 3942 2496 3948 2497
rect 2170 2495 2176 2496
rect 2170 2491 2171 2495
rect 2175 2491 2176 2495
rect 2170 2490 2176 2491
rect 2290 2495 2296 2496
rect 2290 2491 2291 2495
rect 2295 2491 2296 2495
rect 2290 2490 2296 2491
rect 2418 2495 2424 2496
rect 2418 2491 2419 2495
rect 2423 2491 2424 2495
rect 2418 2490 2424 2491
rect 2546 2495 2552 2496
rect 2546 2491 2547 2495
rect 2551 2491 2552 2495
rect 2546 2490 2552 2491
rect 2666 2495 2672 2496
rect 2666 2491 2667 2495
rect 2671 2491 2672 2495
rect 2666 2490 2672 2491
rect 2794 2495 2800 2496
rect 2794 2491 2795 2495
rect 2799 2491 2800 2495
rect 2794 2490 2800 2491
rect 2914 2495 2920 2496
rect 2914 2491 2915 2495
rect 2919 2491 2920 2495
rect 2914 2490 2920 2491
rect 3042 2495 3048 2496
rect 3042 2491 3043 2495
rect 3047 2491 3048 2495
rect 3042 2490 3048 2491
rect 3170 2495 3176 2496
rect 3170 2491 3171 2495
rect 3175 2491 3176 2495
rect 3170 2490 3176 2491
rect 3214 2495 3220 2496
rect 3214 2491 3215 2495
rect 3219 2494 3220 2495
rect 3219 2492 3265 2494
rect 3219 2491 3220 2492
rect 3214 2490 3220 2491
rect 2094 2485 2100 2486
rect 2046 2484 2052 2485
rect 2046 2480 2047 2484
rect 2051 2480 2052 2484
rect 2094 2481 2095 2485
rect 2099 2481 2100 2485
rect 2094 2480 2100 2481
rect 2214 2485 2220 2486
rect 2214 2481 2215 2485
rect 2219 2481 2220 2485
rect 2214 2480 2220 2481
rect 2342 2485 2348 2486
rect 2342 2481 2343 2485
rect 2347 2481 2348 2485
rect 2342 2480 2348 2481
rect 2470 2485 2476 2486
rect 2470 2481 2471 2485
rect 2475 2481 2476 2485
rect 2470 2480 2476 2481
rect 2598 2485 2604 2486
rect 2598 2481 2599 2485
rect 2603 2481 2604 2485
rect 2598 2480 2604 2481
rect 2718 2485 2724 2486
rect 2718 2481 2719 2485
rect 2723 2481 2724 2485
rect 2718 2480 2724 2481
rect 2838 2485 2844 2486
rect 2838 2481 2839 2485
rect 2843 2481 2844 2485
rect 2838 2480 2844 2481
rect 2966 2485 2972 2486
rect 2966 2481 2967 2485
rect 2971 2481 2972 2485
rect 2966 2480 2972 2481
rect 3094 2485 3100 2486
rect 3094 2481 3095 2485
rect 3099 2481 3100 2485
rect 3094 2480 3100 2481
rect 3222 2485 3228 2486
rect 3222 2481 3223 2485
rect 3227 2481 3228 2485
rect 3222 2480 3228 2481
rect 3942 2484 3948 2485
rect 3942 2480 3943 2484
rect 3947 2480 3948 2484
rect 2046 2479 2052 2480
rect 3942 2479 3948 2480
rect 502 2476 508 2477
rect 110 2473 116 2474
rect 110 2469 111 2473
rect 115 2469 116 2473
rect 502 2472 503 2476
rect 507 2472 508 2476
rect 502 2471 508 2472
rect 606 2476 612 2477
rect 606 2472 607 2476
rect 611 2472 612 2476
rect 606 2471 612 2472
rect 718 2476 724 2477
rect 718 2472 719 2476
rect 723 2472 724 2476
rect 718 2471 724 2472
rect 846 2476 852 2477
rect 846 2472 847 2476
rect 851 2472 852 2476
rect 846 2471 852 2472
rect 982 2476 988 2477
rect 982 2472 983 2476
rect 987 2472 988 2476
rect 982 2471 988 2472
rect 1126 2476 1132 2477
rect 1126 2472 1127 2476
rect 1131 2472 1132 2476
rect 1126 2471 1132 2472
rect 1278 2476 1284 2477
rect 1278 2472 1279 2476
rect 1283 2472 1284 2476
rect 1278 2471 1284 2472
rect 1430 2476 1436 2477
rect 1430 2472 1431 2476
rect 1435 2472 1436 2476
rect 1430 2471 1436 2472
rect 1582 2476 1588 2477
rect 1582 2472 1583 2476
rect 1587 2472 1588 2476
rect 1582 2471 1588 2472
rect 1742 2476 1748 2477
rect 1742 2472 1743 2476
rect 1747 2472 1748 2476
rect 1742 2471 1748 2472
rect 1902 2476 1908 2477
rect 1902 2472 1903 2476
rect 1907 2472 1908 2476
rect 2358 2475 2364 2476
rect 1902 2471 1908 2472
rect 2006 2473 2012 2474
rect 110 2468 116 2469
rect 2006 2469 2007 2473
rect 2011 2469 2012 2473
rect 2358 2471 2359 2475
rect 2363 2474 2364 2475
rect 2363 2472 2422 2474
rect 2363 2471 2364 2472
rect 2358 2470 2364 2471
rect 2006 2468 2012 2469
rect 578 2467 584 2468
rect 578 2463 579 2467
rect 583 2463 584 2467
rect 578 2462 584 2463
rect 682 2467 688 2468
rect 682 2463 683 2467
rect 687 2463 688 2467
rect 682 2462 688 2463
rect 702 2467 708 2468
rect 702 2463 703 2467
rect 707 2466 708 2467
rect 922 2467 928 2468
rect 707 2464 761 2466
rect 707 2463 708 2464
rect 702 2462 708 2463
rect 922 2463 923 2467
rect 927 2463 928 2467
rect 922 2462 928 2463
rect 930 2467 936 2468
rect 930 2463 931 2467
rect 935 2466 936 2467
rect 1066 2467 1072 2468
rect 935 2464 1025 2466
rect 935 2463 936 2464
rect 930 2462 936 2463
rect 1066 2463 1067 2467
rect 1071 2466 1072 2467
rect 1354 2467 1360 2468
rect 1071 2464 1169 2466
rect 1071 2463 1072 2464
rect 1066 2462 1072 2463
rect 1354 2463 1355 2467
rect 1359 2463 1360 2467
rect 1354 2462 1360 2463
rect 1362 2467 1368 2468
rect 1362 2463 1363 2467
rect 1367 2466 1368 2467
rect 1658 2467 1664 2468
rect 1367 2464 1473 2466
rect 1367 2463 1368 2464
rect 1362 2462 1368 2463
rect 1658 2463 1659 2467
rect 1663 2463 1664 2467
rect 1658 2462 1664 2463
rect 1818 2467 1824 2468
rect 1818 2463 1819 2467
rect 1823 2463 1824 2467
rect 1818 2462 1824 2463
rect 1970 2467 1976 2468
rect 1970 2463 1971 2467
rect 1975 2463 1976 2467
rect 1970 2462 1976 2463
rect 2146 2463 2152 2464
rect 2146 2459 2147 2463
rect 2151 2462 2152 2463
rect 2159 2463 2165 2464
rect 2159 2462 2160 2463
rect 2151 2460 2160 2462
rect 2151 2459 2152 2460
rect 2146 2458 2152 2459
rect 2159 2459 2160 2460
rect 2164 2459 2165 2463
rect 2159 2458 2165 2459
rect 2170 2463 2176 2464
rect 2170 2459 2171 2463
rect 2175 2462 2176 2463
rect 2279 2463 2285 2464
rect 2279 2462 2280 2463
rect 2175 2460 2280 2462
rect 2175 2459 2176 2460
rect 2170 2458 2176 2459
rect 2279 2459 2280 2460
rect 2284 2459 2285 2463
rect 2279 2458 2285 2459
rect 2290 2463 2296 2464
rect 2290 2459 2291 2463
rect 2295 2462 2296 2463
rect 2407 2463 2413 2464
rect 2407 2462 2408 2463
rect 2295 2460 2408 2462
rect 2295 2459 2296 2460
rect 2290 2458 2296 2459
rect 2407 2459 2408 2460
rect 2412 2459 2413 2463
rect 2420 2462 2422 2472
rect 2535 2463 2541 2464
rect 2535 2462 2536 2463
rect 2420 2460 2536 2462
rect 2407 2458 2413 2459
rect 2535 2459 2536 2460
rect 2540 2459 2541 2463
rect 2535 2458 2541 2459
rect 2546 2463 2552 2464
rect 2546 2459 2547 2463
rect 2551 2462 2552 2463
rect 2663 2463 2669 2464
rect 2663 2462 2664 2463
rect 2551 2460 2664 2462
rect 2551 2459 2552 2460
rect 2546 2458 2552 2459
rect 2663 2459 2664 2460
rect 2668 2459 2669 2463
rect 2663 2458 2669 2459
rect 2783 2463 2792 2464
rect 2783 2459 2784 2463
rect 2791 2459 2792 2463
rect 2783 2458 2792 2459
rect 2794 2463 2800 2464
rect 2794 2459 2795 2463
rect 2799 2462 2800 2463
rect 2903 2463 2909 2464
rect 2903 2462 2904 2463
rect 2799 2460 2904 2462
rect 2799 2459 2800 2460
rect 2794 2458 2800 2459
rect 2903 2459 2904 2460
rect 2908 2459 2909 2463
rect 2903 2458 2909 2459
rect 2914 2463 2920 2464
rect 2914 2459 2915 2463
rect 2919 2462 2920 2463
rect 3031 2463 3037 2464
rect 3031 2462 3032 2463
rect 2919 2460 3032 2462
rect 2919 2459 2920 2460
rect 2914 2458 2920 2459
rect 3031 2459 3032 2460
rect 3036 2459 3037 2463
rect 3031 2458 3037 2459
rect 3042 2463 3048 2464
rect 3042 2459 3043 2463
rect 3047 2462 3048 2463
rect 3159 2463 3165 2464
rect 3159 2462 3160 2463
rect 3047 2460 3160 2462
rect 3047 2459 3048 2460
rect 3042 2458 3048 2459
rect 3159 2459 3160 2460
rect 3164 2459 3165 2463
rect 3159 2458 3165 2459
rect 3170 2463 3176 2464
rect 3170 2459 3171 2463
rect 3175 2462 3176 2463
rect 3287 2463 3293 2464
rect 3287 2462 3288 2463
rect 3175 2460 3288 2462
rect 3175 2459 3176 2460
rect 3170 2458 3176 2459
rect 3287 2459 3288 2460
rect 3292 2459 3293 2463
rect 3287 2458 3293 2459
rect 502 2457 508 2458
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 502 2453 503 2457
rect 507 2453 508 2457
rect 502 2452 508 2453
rect 606 2457 612 2458
rect 606 2453 607 2457
rect 611 2453 612 2457
rect 606 2452 612 2453
rect 718 2457 724 2458
rect 718 2453 719 2457
rect 723 2453 724 2457
rect 718 2452 724 2453
rect 846 2457 852 2458
rect 846 2453 847 2457
rect 851 2453 852 2457
rect 846 2452 852 2453
rect 982 2457 988 2458
rect 982 2453 983 2457
rect 987 2453 988 2457
rect 982 2452 988 2453
rect 1126 2457 1132 2458
rect 1126 2453 1127 2457
rect 1131 2453 1132 2457
rect 1126 2452 1132 2453
rect 1278 2457 1284 2458
rect 1278 2453 1279 2457
rect 1283 2453 1284 2457
rect 1278 2452 1284 2453
rect 1430 2457 1436 2458
rect 1430 2453 1431 2457
rect 1435 2453 1436 2457
rect 1430 2452 1436 2453
rect 1582 2457 1588 2458
rect 1582 2453 1583 2457
rect 1587 2453 1588 2457
rect 1582 2452 1588 2453
rect 1742 2457 1748 2458
rect 1742 2453 1743 2457
rect 1747 2453 1748 2457
rect 1742 2452 1748 2453
rect 1902 2457 1908 2458
rect 1902 2453 1903 2457
rect 1907 2453 1908 2457
rect 1902 2452 1908 2453
rect 2006 2456 2012 2457
rect 2006 2452 2007 2456
rect 2011 2452 2012 2456
rect 110 2451 116 2452
rect 2006 2451 2012 2452
rect 578 2443 584 2444
rect 578 2439 579 2443
rect 583 2442 584 2443
rect 583 2440 630 2442
rect 583 2439 584 2440
rect 578 2438 584 2439
rect 567 2435 573 2436
rect 567 2431 568 2435
rect 572 2434 573 2435
rect 618 2435 624 2436
rect 618 2434 619 2435
rect 572 2432 619 2434
rect 572 2431 573 2432
rect 567 2430 573 2431
rect 618 2431 619 2432
rect 623 2431 624 2435
rect 628 2434 630 2440
rect 2135 2439 2141 2440
rect 671 2435 677 2436
rect 671 2434 672 2435
rect 628 2432 672 2434
rect 618 2430 624 2431
rect 671 2431 672 2432
rect 676 2431 677 2435
rect 671 2430 677 2431
rect 682 2435 688 2436
rect 682 2431 683 2435
rect 687 2434 688 2435
rect 783 2435 789 2436
rect 783 2434 784 2435
rect 687 2432 784 2434
rect 687 2431 688 2432
rect 682 2430 688 2431
rect 783 2431 784 2432
rect 788 2431 789 2435
rect 783 2430 789 2431
rect 911 2435 917 2436
rect 911 2431 912 2435
rect 916 2434 917 2435
rect 930 2435 936 2436
rect 930 2434 931 2435
rect 916 2432 931 2434
rect 916 2431 917 2432
rect 911 2430 917 2431
rect 930 2431 931 2432
rect 935 2431 936 2435
rect 930 2430 936 2431
rect 1047 2435 1053 2436
rect 1047 2431 1048 2435
rect 1052 2434 1053 2435
rect 1066 2435 1072 2436
rect 1066 2434 1067 2435
rect 1052 2432 1067 2434
rect 1052 2431 1053 2432
rect 1047 2430 1053 2431
rect 1066 2431 1067 2432
rect 1071 2431 1072 2435
rect 1066 2430 1072 2431
rect 1146 2435 1152 2436
rect 1146 2431 1147 2435
rect 1151 2434 1152 2435
rect 1191 2435 1197 2436
rect 1191 2434 1192 2435
rect 1151 2432 1192 2434
rect 1151 2431 1152 2432
rect 1146 2430 1152 2431
rect 1191 2431 1192 2432
rect 1196 2431 1197 2435
rect 1191 2430 1197 2431
rect 1343 2435 1349 2436
rect 1343 2431 1344 2435
rect 1348 2434 1349 2435
rect 1362 2435 1368 2436
rect 1362 2434 1363 2435
rect 1348 2432 1363 2434
rect 1348 2431 1349 2432
rect 1343 2430 1349 2431
rect 1362 2431 1363 2432
rect 1367 2431 1368 2435
rect 1362 2430 1368 2431
rect 1495 2435 1501 2436
rect 1495 2431 1496 2435
rect 1500 2434 1501 2435
rect 1519 2435 1525 2436
rect 1519 2434 1520 2435
rect 1500 2432 1520 2434
rect 1500 2431 1501 2432
rect 1495 2430 1501 2431
rect 1519 2431 1520 2432
rect 1524 2431 1525 2435
rect 1519 2430 1525 2431
rect 1570 2435 1576 2436
rect 1570 2431 1571 2435
rect 1575 2434 1576 2435
rect 1647 2435 1653 2436
rect 1647 2434 1648 2435
rect 1575 2432 1648 2434
rect 1575 2431 1576 2432
rect 1570 2430 1576 2431
rect 1647 2431 1648 2432
rect 1652 2431 1653 2435
rect 1647 2430 1653 2431
rect 1658 2435 1664 2436
rect 1658 2431 1659 2435
rect 1663 2434 1664 2435
rect 1807 2435 1813 2436
rect 1807 2434 1808 2435
rect 1663 2432 1808 2434
rect 1663 2431 1664 2432
rect 1658 2430 1664 2431
rect 1807 2431 1808 2432
rect 1812 2431 1813 2435
rect 1807 2430 1813 2431
rect 1818 2435 1824 2436
rect 1818 2431 1819 2435
rect 1823 2434 1824 2435
rect 1967 2435 1973 2436
rect 1967 2434 1968 2435
rect 1823 2432 1968 2434
rect 1823 2431 1824 2432
rect 1818 2430 1824 2431
rect 1967 2431 1968 2432
rect 1972 2431 1973 2435
rect 2135 2435 2136 2439
rect 2140 2438 2141 2439
rect 2242 2439 2248 2440
rect 2140 2436 2238 2438
rect 2140 2435 2141 2436
rect 2135 2434 2141 2435
rect 1967 2430 1973 2431
rect 2236 2430 2238 2436
rect 2242 2435 2243 2439
rect 2247 2438 2248 2439
rect 2255 2439 2261 2440
rect 2255 2438 2256 2439
rect 2247 2436 2256 2438
rect 2247 2435 2248 2436
rect 2242 2434 2248 2435
rect 2255 2435 2256 2436
rect 2260 2435 2261 2439
rect 2255 2434 2261 2435
rect 2266 2439 2272 2440
rect 2266 2435 2267 2439
rect 2271 2438 2272 2439
rect 2383 2439 2389 2440
rect 2383 2438 2384 2439
rect 2271 2436 2384 2438
rect 2271 2435 2272 2436
rect 2266 2434 2272 2435
rect 2383 2435 2384 2436
rect 2388 2435 2389 2439
rect 2383 2434 2389 2435
rect 2503 2439 2509 2440
rect 2503 2435 2504 2439
rect 2508 2438 2509 2439
rect 2522 2439 2528 2440
rect 2522 2438 2523 2439
rect 2508 2436 2523 2438
rect 2508 2435 2509 2436
rect 2503 2434 2509 2435
rect 2522 2435 2523 2436
rect 2527 2435 2528 2439
rect 2522 2434 2528 2435
rect 2623 2439 2629 2440
rect 2623 2435 2624 2439
rect 2628 2438 2629 2439
rect 2666 2439 2672 2440
rect 2666 2438 2667 2439
rect 2628 2436 2667 2438
rect 2628 2435 2629 2436
rect 2623 2434 2629 2435
rect 2666 2435 2667 2436
rect 2671 2435 2672 2439
rect 2666 2434 2672 2435
rect 2743 2439 2749 2440
rect 2743 2435 2744 2439
rect 2748 2438 2749 2439
rect 2762 2439 2768 2440
rect 2762 2438 2763 2439
rect 2748 2436 2763 2438
rect 2748 2435 2749 2436
rect 2743 2434 2749 2435
rect 2762 2435 2763 2436
rect 2767 2435 2768 2439
rect 2762 2434 2768 2435
rect 2855 2439 2861 2440
rect 2855 2435 2856 2439
rect 2860 2438 2861 2439
rect 2874 2439 2880 2440
rect 2874 2438 2875 2439
rect 2860 2436 2875 2438
rect 2860 2435 2861 2436
rect 2855 2434 2861 2435
rect 2874 2435 2875 2436
rect 2879 2435 2880 2439
rect 2874 2434 2880 2435
rect 2975 2439 2981 2440
rect 2975 2435 2976 2439
rect 2980 2438 2981 2439
rect 2994 2439 3000 2440
rect 2994 2438 2995 2439
rect 2980 2436 2995 2438
rect 2980 2435 2981 2436
rect 2975 2434 2981 2435
rect 2994 2435 2995 2436
rect 2999 2435 3000 2439
rect 2994 2434 3000 2435
rect 3095 2439 3101 2440
rect 3095 2435 3096 2439
rect 3100 2438 3101 2439
rect 3114 2439 3120 2440
rect 3114 2438 3115 2439
rect 3100 2436 3115 2438
rect 3100 2435 3101 2436
rect 3095 2434 3101 2435
rect 3114 2435 3115 2436
rect 3119 2435 3120 2439
rect 3114 2434 3120 2435
rect 3214 2439 3221 2440
rect 3214 2435 3215 2439
rect 3220 2435 3221 2439
rect 3214 2434 3221 2435
rect 2274 2431 2280 2432
rect 2274 2430 2275 2431
rect 2236 2428 2275 2430
rect 2274 2427 2275 2428
rect 2279 2427 2280 2431
rect 2274 2426 2280 2427
rect 2046 2420 2052 2421
rect 3942 2420 3948 2421
rect 2046 2416 2047 2420
rect 2051 2416 2052 2420
rect 922 2415 928 2416
rect 2046 2415 2052 2416
rect 2070 2419 2076 2420
rect 2070 2415 2071 2419
rect 2075 2415 2076 2419
rect 922 2411 923 2415
rect 927 2414 928 2415
rect 2070 2414 2076 2415
rect 2190 2419 2196 2420
rect 2190 2415 2191 2419
rect 2195 2415 2196 2419
rect 2190 2414 2196 2415
rect 2318 2419 2324 2420
rect 2318 2415 2319 2419
rect 2323 2415 2324 2419
rect 2318 2414 2324 2415
rect 2438 2419 2444 2420
rect 2438 2415 2439 2419
rect 2443 2415 2444 2419
rect 2438 2414 2444 2415
rect 2558 2419 2564 2420
rect 2558 2415 2559 2419
rect 2563 2415 2564 2419
rect 2558 2414 2564 2415
rect 2678 2419 2684 2420
rect 2678 2415 2679 2419
rect 2683 2415 2684 2419
rect 2678 2414 2684 2415
rect 2790 2419 2796 2420
rect 2790 2415 2791 2419
rect 2795 2415 2796 2419
rect 2790 2414 2796 2415
rect 2910 2419 2916 2420
rect 2910 2415 2911 2419
rect 2915 2415 2916 2419
rect 2910 2414 2916 2415
rect 3030 2419 3036 2420
rect 3030 2415 3031 2419
rect 3035 2415 3036 2419
rect 3030 2414 3036 2415
rect 3150 2419 3156 2420
rect 3150 2415 3151 2419
rect 3155 2415 3156 2419
rect 3942 2416 3943 2420
rect 3947 2416 3948 2420
rect 3942 2415 3948 2416
rect 3150 2414 3156 2415
rect 927 2412 1018 2414
rect 927 2411 928 2412
rect 922 2410 928 2411
rect 599 2407 605 2408
rect 599 2403 600 2407
rect 604 2406 605 2407
rect 655 2407 661 2408
rect 655 2406 656 2407
rect 604 2404 656 2406
rect 604 2403 605 2404
rect 599 2402 605 2403
rect 655 2403 656 2404
rect 660 2403 661 2407
rect 655 2402 661 2403
rect 730 2407 741 2408
rect 730 2403 731 2407
rect 735 2403 736 2407
rect 740 2403 741 2407
rect 730 2402 741 2403
rect 879 2407 885 2408
rect 879 2403 880 2407
rect 884 2406 885 2407
rect 1016 2406 1018 2412
rect 2146 2411 2152 2412
rect 1023 2407 1029 2408
rect 1023 2406 1024 2407
rect 884 2404 1014 2406
rect 1016 2404 1024 2406
rect 884 2403 885 2404
rect 879 2402 885 2403
rect 1012 2398 1014 2404
rect 1023 2403 1024 2404
rect 1028 2403 1029 2407
rect 1023 2402 1029 2403
rect 1034 2407 1040 2408
rect 1034 2403 1035 2407
rect 1039 2406 1040 2407
rect 1167 2407 1173 2408
rect 1167 2406 1168 2407
rect 1039 2404 1168 2406
rect 1039 2403 1040 2404
rect 1034 2402 1040 2403
rect 1167 2403 1168 2404
rect 1172 2403 1173 2407
rect 1167 2402 1173 2403
rect 1311 2407 1317 2408
rect 1311 2403 1312 2407
rect 1316 2406 1317 2407
rect 1322 2407 1328 2408
rect 1316 2403 1318 2406
rect 1311 2402 1318 2403
rect 1322 2403 1323 2407
rect 1327 2406 1328 2407
rect 1455 2407 1461 2408
rect 1455 2406 1456 2407
rect 1327 2404 1456 2406
rect 1327 2403 1328 2404
rect 1322 2402 1328 2403
rect 1455 2403 1456 2404
rect 1460 2403 1461 2407
rect 1455 2402 1461 2403
rect 1466 2407 1472 2408
rect 1466 2403 1467 2407
rect 1471 2406 1472 2407
rect 1591 2407 1597 2408
rect 1591 2406 1592 2407
rect 1471 2404 1592 2406
rect 1471 2403 1472 2404
rect 1466 2402 1472 2403
rect 1591 2403 1592 2404
rect 1596 2403 1597 2407
rect 1591 2402 1597 2403
rect 1719 2407 1725 2408
rect 1719 2403 1720 2407
rect 1724 2406 1725 2407
rect 1730 2407 1736 2408
rect 1724 2403 1726 2406
rect 1719 2402 1726 2403
rect 1730 2403 1731 2407
rect 1735 2406 1736 2407
rect 1855 2407 1861 2408
rect 1855 2406 1856 2407
rect 1735 2404 1856 2406
rect 1735 2403 1736 2404
rect 1730 2402 1736 2403
rect 1855 2403 1856 2404
rect 1860 2403 1861 2407
rect 1855 2402 1861 2403
rect 1967 2407 1976 2408
rect 1967 2403 1968 2407
rect 1975 2403 1976 2407
rect 2146 2407 2147 2411
rect 2151 2407 2152 2411
rect 2146 2406 2152 2407
rect 2266 2411 2272 2412
rect 2266 2407 2267 2411
rect 2271 2407 2272 2411
rect 2266 2406 2272 2407
rect 2274 2411 2280 2412
rect 2274 2407 2275 2411
rect 2279 2410 2280 2411
rect 2422 2411 2428 2412
rect 2279 2408 2361 2410
rect 2279 2407 2280 2408
rect 2274 2406 2280 2407
rect 2422 2407 2423 2411
rect 2427 2410 2428 2411
rect 2522 2411 2528 2412
rect 2427 2408 2481 2410
rect 2427 2407 2428 2408
rect 2422 2406 2428 2407
rect 2522 2407 2523 2411
rect 2527 2410 2528 2411
rect 2642 2411 2648 2412
rect 2527 2408 2601 2410
rect 2527 2407 2528 2408
rect 2522 2406 2528 2407
rect 2642 2407 2643 2411
rect 2647 2410 2648 2411
rect 2762 2411 2768 2412
rect 2647 2408 2721 2410
rect 2647 2407 2648 2408
rect 2642 2406 2648 2407
rect 2762 2407 2763 2411
rect 2767 2410 2768 2411
rect 2874 2411 2880 2412
rect 2767 2408 2833 2410
rect 2767 2407 2768 2408
rect 2762 2406 2768 2407
rect 2874 2407 2875 2411
rect 2879 2410 2880 2411
rect 2994 2411 3000 2412
rect 2879 2408 2953 2410
rect 2879 2407 2880 2408
rect 2874 2406 2880 2407
rect 2994 2407 2995 2411
rect 2999 2410 3000 2411
rect 3114 2411 3120 2412
rect 2999 2408 3073 2410
rect 2999 2407 3000 2408
rect 2994 2406 3000 2407
rect 3114 2407 3115 2411
rect 3119 2410 3120 2411
rect 3119 2408 3193 2410
rect 3119 2407 3120 2408
rect 3114 2406 3120 2407
rect 1967 2402 1976 2403
rect 2046 2403 2052 2404
rect 1042 2399 1048 2400
rect 1042 2398 1043 2399
rect 1012 2396 1043 2398
rect 1042 2395 1043 2396
rect 1047 2395 1048 2399
rect 1316 2398 1318 2402
rect 1378 2399 1384 2400
rect 1378 2398 1379 2399
rect 1316 2396 1379 2398
rect 1042 2394 1048 2395
rect 1378 2395 1379 2396
rect 1383 2395 1384 2399
rect 1724 2398 1726 2402
rect 1874 2399 1880 2400
rect 1874 2398 1875 2399
rect 1724 2396 1875 2398
rect 1378 2394 1384 2395
rect 1874 2395 1875 2396
rect 1879 2395 1880 2399
rect 2046 2399 2047 2403
rect 2051 2399 2052 2403
rect 3942 2403 3948 2404
rect 2046 2398 2052 2399
rect 2070 2400 2076 2401
rect 2070 2396 2071 2400
rect 2075 2396 2076 2400
rect 2070 2395 2076 2396
rect 2190 2400 2196 2401
rect 2190 2396 2191 2400
rect 2195 2396 2196 2400
rect 2190 2395 2196 2396
rect 2318 2400 2324 2401
rect 2318 2396 2319 2400
rect 2323 2396 2324 2400
rect 2318 2395 2324 2396
rect 2438 2400 2444 2401
rect 2438 2396 2439 2400
rect 2443 2396 2444 2400
rect 2438 2395 2444 2396
rect 2558 2400 2564 2401
rect 2558 2396 2559 2400
rect 2563 2396 2564 2400
rect 2558 2395 2564 2396
rect 2678 2400 2684 2401
rect 2678 2396 2679 2400
rect 2683 2396 2684 2400
rect 2678 2395 2684 2396
rect 2790 2400 2796 2401
rect 2790 2396 2791 2400
rect 2795 2396 2796 2400
rect 2790 2395 2796 2396
rect 2910 2400 2916 2401
rect 2910 2396 2911 2400
rect 2915 2396 2916 2400
rect 2910 2395 2916 2396
rect 3030 2400 3036 2401
rect 3030 2396 3031 2400
rect 3035 2396 3036 2400
rect 3030 2395 3036 2396
rect 3150 2400 3156 2401
rect 3150 2396 3151 2400
rect 3155 2396 3156 2400
rect 3942 2399 3943 2403
rect 3947 2399 3948 2403
rect 3942 2398 3948 2399
rect 3150 2395 3156 2396
rect 1874 2394 1880 2395
rect 110 2388 116 2389
rect 2006 2388 2012 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 534 2387 540 2388
rect 534 2383 535 2387
rect 539 2383 540 2387
rect 534 2382 540 2383
rect 670 2387 676 2388
rect 670 2383 671 2387
rect 675 2383 676 2387
rect 670 2382 676 2383
rect 814 2387 820 2388
rect 814 2383 815 2387
rect 819 2383 820 2387
rect 814 2382 820 2383
rect 958 2387 964 2388
rect 958 2383 959 2387
rect 963 2383 964 2387
rect 958 2382 964 2383
rect 1102 2387 1108 2388
rect 1102 2383 1103 2387
rect 1107 2383 1108 2387
rect 1102 2382 1108 2383
rect 1246 2387 1252 2388
rect 1246 2383 1247 2387
rect 1251 2383 1252 2387
rect 1246 2382 1252 2383
rect 1390 2387 1396 2388
rect 1390 2383 1391 2387
rect 1395 2383 1396 2387
rect 1390 2382 1396 2383
rect 1526 2387 1532 2388
rect 1526 2383 1527 2387
rect 1531 2383 1532 2387
rect 1526 2382 1532 2383
rect 1654 2387 1660 2388
rect 1654 2383 1655 2387
rect 1659 2383 1660 2387
rect 1654 2382 1660 2383
rect 1790 2387 1796 2388
rect 1790 2383 1791 2387
rect 1795 2383 1796 2387
rect 1790 2382 1796 2383
rect 1902 2387 1908 2388
rect 1902 2383 1903 2387
rect 1907 2383 1908 2387
rect 2006 2384 2007 2388
rect 2011 2384 2012 2388
rect 2006 2383 2012 2384
rect 1902 2382 1908 2383
rect 618 2379 624 2380
rect 618 2378 619 2379
rect 613 2376 619 2378
rect 618 2375 619 2376
rect 623 2375 624 2379
rect 618 2374 624 2375
rect 655 2379 661 2380
rect 655 2375 656 2379
rect 660 2378 661 2379
rect 1034 2379 1040 2380
rect 660 2376 713 2378
rect 660 2375 661 2376
rect 655 2374 661 2375
rect 1034 2375 1035 2379
rect 1039 2375 1040 2379
rect 1034 2374 1040 2375
rect 1042 2379 1048 2380
rect 1042 2375 1043 2379
rect 1047 2378 1048 2379
rect 1322 2379 1328 2380
rect 1047 2376 1145 2378
rect 1047 2375 1048 2376
rect 1042 2374 1048 2375
rect 1322 2375 1323 2379
rect 1327 2375 1328 2379
rect 1322 2374 1328 2375
rect 1466 2379 1472 2380
rect 1466 2375 1467 2379
rect 1471 2375 1472 2379
rect 1466 2374 1472 2375
rect 1519 2379 1525 2380
rect 1519 2375 1520 2379
rect 1524 2378 1525 2379
rect 1730 2379 1736 2380
rect 1524 2376 1569 2378
rect 1524 2375 1525 2376
rect 1519 2374 1525 2375
rect 1730 2375 1731 2379
rect 1735 2375 1736 2379
rect 1874 2379 1880 2380
rect 1730 2374 1736 2375
rect 1866 2375 1872 2376
rect 110 2371 116 2372
rect 110 2367 111 2371
rect 115 2367 116 2371
rect 882 2371 888 2372
rect 110 2366 116 2367
rect 534 2368 540 2369
rect 534 2364 535 2368
rect 539 2364 540 2368
rect 534 2363 540 2364
rect 670 2368 676 2369
rect 670 2364 671 2368
rect 675 2364 676 2368
rect 670 2363 676 2364
rect 814 2368 820 2369
rect 814 2364 815 2368
rect 819 2364 820 2368
rect 882 2367 883 2371
rect 887 2370 888 2371
rect 892 2370 894 2373
rect 1866 2371 1867 2375
rect 1871 2371 1872 2375
rect 1874 2375 1875 2379
rect 1879 2378 1880 2379
rect 1879 2376 1945 2378
rect 1879 2375 1880 2376
rect 1874 2374 1880 2375
rect 1866 2370 1872 2371
rect 2006 2371 2012 2372
rect 887 2368 894 2370
rect 958 2368 964 2369
rect 887 2367 888 2368
rect 882 2366 888 2367
rect 814 2363 820 2364
rect 958 2364 959 2368
rect 963 2364 964 2368
rect 958 2363 964 2364
rect 1102 2368 1108 2369
rect 1102 2364 1103 2368
rect 1107 2364 1108 2368
rect 1102 2363 1108 2364
rect 1246 2368 1252 2369
rect 1246 2364 1247 2368
rect 1251 2364 1252 2368
rect 1246 2363 1252 2364
rect 1390 2368 1396 2369
rect 1390 2364 1391 2368
rect 1395 2364 1396 2368
rect 1390 2363 1396 2364
rect 1526 2368 1532 2369
rect 1526 2364 1527 2368
rect 1531 2364 1532 2368
rect 1526 2363 1532 2364
rect 1654 2368 1660 2369
rect 1654 2364 1655 2368
rect 1659 2364 1660 2368
rect 1654 2363 1660 2364
rect 1790 2368 1796 2369
rect 1790 2364 1791 2368
rect 1795 2364 1796 2368
rect 1790 2363 1796 2364
rect 1902 2368 1908 2369
rect 1902 2364 1903 2368
rect 1907 2364 1908 2368
rect 2006 2367 2007 2371
rect 2011 2367 2012 2371
rect 2006 2366 2012 2367
rect 1902 2363 1908 2364
rect 2166 2336 2172 2337
rect 2046 2333 2052 2334
rect 2046 2329 2047 2333
rect 2051 2329 2052 2333
rect 2166 2332 2167 2336
rect 2171 2332 2172 2336
rect 2166 2331 2172 2332
rect 2358 2336 2364 2337
rect 2358 2332 2359 2336
rect 2363 2332 2364 2336
rect 2358 2331 2364 2332
rect 2534 2336 2540 2337
rect 2534 2332 2535 2336
rect 2539 2332 2540 2336
rect 2534 2331 2540 2332
rect 2702 2336 2708 2337
rect 2702 2332 2703 2336
rect 2707 2332 2708 2336
rect 2702 2331 2708 2332
rect 2870 2336 2876 2337
rect 2870 2332 2871 2336
rect 2875 2332 2876 2336
rect 2870 2331 2876 2332
rect 3030 2336 3036 2337
rect 3030 2332 3031 2336
rect 3035 2332 3036 2336
rect 3030 2331 3036 2332
rect 3198 2336 3204 2337
rect 3198 2332 3199 2336
rect 3203 2332 3204 2336
rect 3198 2331 3204 2332
rect 3942 2333 3948 2334
rect 2046 2328 2052 2329
rect 3942 2329 3943 2333
rect 3947 2329 3948 2333
rect 3942 2328 3948 2329
rect 2242 2327 2248 2328
rect 2242 2323 2243 2327
rect 2247 2323 2248 2327
rect 2242 2322 2248 2323
rect 2350 2327 2356 2328
rect 2350 2323 2351 2327
rect 2355 2326 2356 2327
rect 2670 2327 2676 2328
rect 2670 2326 2671 2327
rect 2355 2324 2401 2326
rect 2613 2324 2671 2326
rect 2355 2323 2356 2324
rect 2350 2322 2356 2323
rect 2670 2323 2671 2324
rect 2675 2323 2676 2327
rect 2670 2322 2676 2323
rect 2778 2327 2784 2328
rect 2778 2323 2779 2327
rect 2783 2323 2784 2327
rect 2778 2322 2784 2323
rect 2946 2327 2952 2328
rect 2946 2323 2947 2327
rect 2951 2323 2952 2327
rect 2946 2322 2952 2323
rect 3106 2327 3112 2328
rect 3106 2323 3107 2327
rect 3111 2323 3112 2327
rect 3106 2322 3112 2323
rect 3114 2327 3120 2328
rect 3114 2323 3115 2327
rect 3119 2326 3120 2327
rect 3119 2324 3241 2326
rect 3119 2323 3120 2324
rect 3114 2322 3120 2323
rect 2166 2317 2172 2318
rect 2046 2316 2052 2317
rect 2046 2312 2047 2316
rect 2051 2312 2052 2316
rect 2166 2313 2167 2317
rect 2171 2313 2172 2317
rect 2166 2312 2172 2313
rect 2358 2317 2364 2318
rect 2358 2313 2359 2317
rect 2363 2313 2364 2317
rect 2358 2312 2364 2313
rect 2534 2317 2540 2318
rect 2534 2313 2535 2317
rect 2539 2313 2540 2317
rect 2534 2312 2540 2313
rect 2702 2317 2708 2318
rect 2702 2313 2703 2317
rect 2707 2313 2708 2317
rect 2702 2312 2708 2313
rect 2870 2317 2876 2318
rect 2870 2313 2871 2317
rect 2875 2313 2876 2317
rect 2870 2312 2876 2313
rect 3030 2317 3036 2318
rect 3030 2313 3031 2317
rect 3035 2313 3036 2317
rect 3030 2312 3036 2313
rect 3198 2317 3204 2318
rect 3198 2313 3199 2317
rect 3203 2313 3204 2317
rect 3198 2312 3204 2313
rect 3942 2316 3948 2317
rect 3942 2312 3943 2316
rect 3947 2312 3948 2316
rect 2046 2311 2052 2312
rect 3942 2311 3948 2312
rect 534 2304 540 2305
rect 110 2301 116 2302
rect 110 2297 111 2301
rect 115 2297 116 2301
rect 534 2300 535 2304
rect 539 2300 540 2304
rect 534 2299 540 2300
rect 646 2304 652 2305
rect 646 2300 647 2304
rect 651 2300 652 2304
rect 646 2299 652 2300
rect 766 2304 772 2305
rect 766 2300 767 2304
rect 771 2300 772 2304
rect 766 2299 772 2300
rect 894 2304 900 2305
rect 894 2300 895 2304
rect 899 2300 900 2304
rect 894 2299 900 2300
rect 1030 2304 1036 2305
rect 1030 2300 1031 2304
rect 1035 2300 1036 2304
rect 1030 2299 1036 2300
rect 1166 2304 1172 2305
rect 1166 2300 1167 2304
rect 1171 2300 1172 2304
rect 1166 2299 1172 2300
rect 1294 2304 1300 2305
rect 1294 2300 1295 2304
rect 1299 2300 1300 2304
rect 1294 2299 1300 2300
rect 1422 2304 1428 2305
rect 1422 2300 1423 2304
rect 1427 2300 1428 2304
rect 1422 2299 1428 2300
rect 1550 2304 1556 2305
rect 1550 2300 1551 2304
rect 1555 2300 1556 2304
rect 1550 2299 1556 2300
rect 1670 2304 1676 2305
rect 1670 2300 1671 2304
rect 1675 2300 1676 2304
rect 1670 2299 1676 2300
rect 1798 2304 1804 2305
rect 1798 2300 1799 2304
rect 1803 2300 1804 2304
rect 1798 2299 1804 2300
rect 1902 2304 1908 2305
rect 1902 2300 1903 2304
rect 1907 2300 1908 2304
rect 1902 2299 1908 2300
rect 2006 2301 2012 2302
rect 110 2296 116 2297
rect 2006 2297 2007 2301
rect 2011 2297 2012 2301
rect 2006 2296 2012 2297
rect 2422 2299 2428 2300
rect 610 2295 616 2296
rect 610 2291 611 2295
rect 615 2291 616 2295
rect 730 2295 736 2296
rect 730 2294 731 2295
rect 725 2292 731 2294
rect 610 2290 616 2291
rect 730 2291 731 2292
rect 735 2291 736 2295
rect 887 2295 893 2296
rect 887 2294 888 2295
rect 845 2292 888 2294
rect 730 2290 736 2291
rect 887 2291 888 2292
rect 892 2291 893 2295
rect 887 2290 893 2291
rect 970 2295 976 2296
rect 970 2291 971 2295
rect 975 2291 976 2295
rect 970 2290 976 2291
rect 1106 2295 1112 2296
rect 1106 2291 1107 2295
rect 1111 2291 1112 2295
rect 1106 2290 1112 2291
rect 1114 2295 1120 2296
rect 1114 2291 1115 2295
rect 1119 2294 1120 2295
rect 1370 2295 1376 2296
rect 1119 2292 1209 2294
rect 1119 2291 1120 2292
rect 1114 2290 1120 2291
rect 1370 2291 1371 2295
rect 1375 2291 1376 2295
rect 1370 2290 1376 2291
rect 1378 2295 1384 2296
rect 1378 2291 1379 2295
rect 1383 2294 1384 2295
rect 1506 2295 1512 2296
rect 1383 2292 1465 2294
rect 1383 2291 1384 2292
rect 1378 2290 1384 2291
rect 1506 2291 1507 2295
rect 1511 2294 1512 2295
rect 1634 2295 1640 2296
rect 1511 2292 1593 2294
rect 1511 2291 1512 2292
rect 1506 2290 1512 2291
rect 1634 2291 1635 2295
rect 1639 2294 1640 2295
rect 1874 2295 1880 2296
rect 1639 2292 1713 2294
rect 1639 2291 1640 2292
rect 1634 2290 1640 2291
rect 1874 2291 1875 2295
rect 1879 2291 1880 2295
rect 2231 2295 2240 2296
rect 1981 2292 2001 2294
rect 1874 2290 1880 2291
rect 1999 2290 2001 2292
rect 2231 2291 2232 2295
rect 2239 2291 2240 2295
rect 2422 2295 2423 2299
rect 2427 2298 2428 2299
rect 2427 2297 2429 2298
rect 2422 2294 2424 2295
rect 2423 2293 2424 2294
rect 2428 2293 2429 2297
rect 2423 2292 2429 2293
rect 2599 2295 2605 2296
rect 2231 2290 2240 2291
rect 2599 2291 2600 2295
rect 2604 2294 2605 2295
rect 2642 2295 2648 2296
rect 2642 2294 2643 2295
rect 2604 2292 2643 2294
rect 2604 2291 2605 2292
rect 2599 2290 2605 2291
rect 2642 2291 2643 2292
rect 2647 2291 2648 2295
rect 2642 2290 2648 2291
rect 2670 2295 2676 2296
rect 2670 2291 2671 2295
rect 2675 2294 2676 2295
rect 2767 2295 2773 2296
rect 2767 2294 2768 2295
rect 2675 2292 2768 2294
rect 2675 2291 2676 2292
rect 2670 2290 2676 2291
rect 2767 2291 2768 2292
rect 2772 2291 2773 2295
rect 2767 2290 2773 2291
rect 2778 2295 2784 2296
rect 2778 2291 2779 2295
rect 2783 2294 2784 2295
rect 2935 2295 2941 2296
rect 2935 2294 2936 2295
rect 2783 2292 2936 2294
rect 2783 2291 2784 2292
rect 2778 2290 2784 2291
rect 2935 2291 2936 2292
rect 2940 2291 2941 2295
rect 2935 2290 2941 2291
rect 2946 2295 2952 2296
rect 2946 2291 2947 2295
rect 2951 2294 2952 2295
rect 3095 2295 3101 2296
rect 3095 2294 3096 2295
rect 2951 2292 3096 2294
rect 2951 2291 2952 2292
rect 2946 2290 2952 2291
rect 3095 2291 3096 2292
rect 3100 2291 3101 2295
rect 3095 2290 3101 2291
rect 3106 2295 3112 2296
rect 3106 2291 3107 2295
rect 3111 2294 3112 2295
rect 3263 2295 3269 2296
rect 3263 2294 3264 2295
rect 3111 2292 3264 2294
rect 3111 2291 3112 2292
rect 3106 2290 3112 2291
rect 3263 2291 3264 2292
rect 3268 2291 3269 2295
rect 3263 2290 3269 2291
rect 1999 2288 2070 2290
rect 534 2285 540 2286
rect 110 2284 116 2285
rect 110 2280 111 2284
rect 115 2280 116 2284
rect 534 2281 535 2285
rect 539 2281 540 2285
rect 534 2280 540 2281
rect 646 2285 652 2286
rect 646 2281 647 2285
rect 651 2281 652 2285
rect 646 2280 652 2281
rect 766 2285 772 2286
rect 766 2281 767 2285
rect 771 2281 772 2285
rect 766 2280 772 2281
rect 894 2285 900 2286
rect 894 2281 895 2285
rect 899 2281 900 2285
rect 894 2280 900 2281
rect 1030 2285 1036 2286
rect 1030 2281 1031 2285
rect 1035 2281 1036 2285
rect 1030 2280 1036 2281
rect 1166 2285 1172 2286
rect 1166 2281 1167 2285
rect 1171 2281 1172 2285
rect 1166 2280 1172 2281
rect 1294 2285 1300 2286
rect 1294 2281 1295 2285
rect 1299 2281 1300 2285
rect 1294 2280 1300 2281
rect 1422 2285 1428 2286
rect 1422 2281 1423 2285
rect 1427 2281 1428 2285
rect 1422 2280 1428 2281
rect 1550 2285 1556 2286
rect 1550 2281 1551 2285
rect 1555 2281 1556 2285
rect 1550 2280 1556 2281
rect 1670 2285 1676 2286
rect 1670 2281 1671 2285
rect 1675 2281 1676 2285
rect 1670 2280 1676 2281
rect 1798 2285 1804 2286
rect 1798 2281 1799 2285
rect 1803 2281 1804 2285
rect 1798 2280 1804 2281
rect 1902 2285 1908 2286
rect 1902 2281 1903 2285
rect 1907 2281 1908 2285
rect 1902 2280 1908 2281
rect 2006 2284 2012 2285
rect 2006 2280 2007 2284
rect 2011 2280 2012 2284
rect 2068 2282 2070 2288
rect 2135 2283 2141 2284
rect 2135 2282 2136 2283
rect 2068 2280 2136 2282
rect 110 2279 116 2280
rect 2006 2279 2012 2280
rect 2135 2279 2136 2280
rect 2140 2279 2141 2283
rect 2135 2278 2141 2279
rect 2146 2283 2152 2284
rect 2146 2279 2147 2283
rect 2151 2282 2152 2283
rect 2231 2283 2237 2284
rect 2231 2282 2232 2283
rect 2151 2280 2232 2282
rect 2151 2279 2152 2280
rect 2146 2278 2152 2279
rect 2231 2279 2232 2280
rect 2236 2279 2237 2283
rect 2231 2278 2237 2279
rect 2350 2283 2357 2284
rect 2350 2279 2351 2283
rect 2356 2279 2357 2283
rect 2350 2278 2357 2279
rect 2370 2283 2376 2284
rect 2370 2279 2371 2283
rect 2375 2282 2376 2283
rect 2487 2283 2493 2284
rect 2487 2282 2488 2283
rect 2375 2280 2488 2282
rect 2375 2279 2376 2280
rect 2370 2278 2376 2279
rect 2487 2279 2488 2280
rect 2492 2279 2493 2283
rect 2487 2278 2493 2279
rect 2498 2283 2504 2284
rect 2498 2279 2499 2283
rect 2503 2282 2504 2283
rect 2623 2283 2629 2284
rect 2623 2282 2624 2283
rect 2503 2280 2624 2282
rect 2503 2279 2504 2280
rect 2498 2278 2504 2279
rect 2623 2279 2624 2280
rect 2628 2279 2629 2283
rect 2623 2278 2629 2279
rect 2634 2283 2640 2284
rect 2634 2279 2635 2283
rect 2639 2282 2640 2283
rect 2767 2283 2773 2284
rect 2767 2282 2768 2283
rect 2639 2280 2768 2282
rect 2639 2279 2640 2280
rect 2634 2278 2640 2279
rect 2767 2279 2768 2280
rect 2772 2279 2773 2283
rect 2767 2278 2773 2279
rect 2903 2283 2909 2284
rect 2903 2279 2904 2283
rect 2908 2279 2909 2283
rect 2903 2278 2909 2279
rect 2914 2283 2920 2284
rect 2914 2279 2915 2283
rect 2919 2282 2920 2283
rect 3047 2283 3053 2284
rect 3047 2282 3048 2283
rect 2919 2280 3048 2282
rect 2919 2279 2920 2280
rect 2914 2278 2920 2279
rect 3047 2279 3048 2280
rect 3052 2279 3053 2283
rect 3047 2278 3053 2279
rect 3058 2283 3064 2284
rect 3058 2279 3059 2283
rect 3063 2282 3064 2283
rect 3191 2283 3197 2284
rect 3191 2282 3192 2283
rect 3063 2280 3192 2282
rect 3063 2279 3064 2280
rect 3058 2278 3064 2279
rect 3191 2279 3192 2280
rect 3196 2279 3197 2283
rect 3191 2278 3197 2279
rect 3250 2283 3256 2284
rect 3250 2279 3251 2283
rect 3255 2282 3256 2283
rect 3335 2283 3341 2284
rect 3335 2282 3336 2283
rect 3255 2280 3336 2282
rect 3255 2279 3256 2280
rect 3250 2278 3256 2279
rect 3335 2279 3336 2280
rect 3340 2279 3341 2283
rect 3335 2278 3341 2279
rect 2905 2274 2907 2278
rect 3114 2275 3120 2276
rect 3114 2274 3115 2275
rect 2905 2272 3115 2274
rect 1506 2271 1512 2272
rect 1506 2270 1507 2271
rect 1364 2268 1507 2270
rect 1364 2264 1366 2268
rect 1506 2267 1507 2268
rect 1511 2267 1512 2271
rect 1506 2266 1512 2267
rect 2234 2271 2240 2272
rect 2234 2267 2235 2271
rect 2239 2270 2240 2271
rect 3114 2271 3115 2272
rect 3119 2271 3120 2275
rect 3114 2270 3120 2271
rect 2239 2268 2646 2270
rect 2239 2267 2240 2268
rect 2234 2266 2240 2267
rect 2046 2264 2052 2265
rect 490 2263 496 2264
rect 490 2259 491 2263
rect 495 2262 496 2263
rect 599 2263 605 2264
rect 599 2262 600 2263
rect 495 2260 600 2262
rect 495 2259 496 2260
rect 490 2258 496 2259
rect 599 2259 600 2260
rect 604 2259 605 2263
rect 599 2258 605 2259
rect 610 2263 616 2264
rect 610 2259 611 2263
rect 615 2262 616 2263
rect 711 2263 717 2264
rect 711 2262 712 2263
rect 615 2260 712 2262
rect 615 2259 616 2260
rect 610 2258 616 2259
rect 711 2259 712 2260
rect 716 2259 717 2263
rect 711 2258 717 2259
rect 831 2263 837 2264
rect 831 2259 832 2263
rect 836 2262 837 2263
rect 882 2263 888 2264
rect 882 2262 883 2263
rect 836 2260 883 2262
rect 836 2259 837 2260
rect 831 2258 837 2259
rect 882 2259 883 2260
rect 887 2259 888 2263
rect 882 2258 888 2259
rect 895 2263 901 2264
rect 895 2259 896 2263
rect 900 2262 901 2263
rect 959 2263 965 2264
rect 959 2262 960 2263
rect 900 2260 960 2262
rect 900 2259 901 2260
rect 895 2258 901 2259
rect 959 2259 960 2260
rect 964 2259 965 2263
rect 959 2258 965 2259
rect 970 2263 976 2264
rect 970 2259 971 2263
rect 975 2262 976 2263
rect 1095 2263 1101 2264
rect 1095 2262 1096 2263
rect 975 2260 1096 2262
rect 975 2259 976 2260
rect 970 2258 976 2259
rect 1095 2259 1096 2260
rect 1100 2259 1101 2263
rect 1095 2258 1101 2259
rect 1106 2263 1112 2264
rect 1106 2259 1107 2263
rect 1111 2262 1112 2263
rect 1231 2263 1237 2264
rect 1231 2262 1232 2263
rect 1111 2260 1232 2262
rect 1111 2259 1112 2260
rect 1106 2258 1112 2259
rect 1231 2259 1232 2260
rect 1236 2259 1237 2263
rect 1231 2258 1237 2259
rect 1359 2263 1366 2264
rect 1359 2259 1360 2263
rect 1364 2260 1366 2263
rect 1370 2263 1376 2264
rect 1364 2259 1365 2260
rect 1359 2258 1365 2259
rect 1370 2259 1371 2263
rect 1375 2262 1376 2263
rect 1487 2263 1493 2264
rect 1487 2262 1488 2263
rect 1375 2260 1488 2262
rect 1375 2259 1376 2260
rect 1370 2258 1376 2259
rect 1487 2259 1488 2260
rect 1492 2259 1493 2263
rect 1487 2258 1493 2259
rect 1615 2263 1621 2264
rect 1615 2259 1616 2263
rect 1620 2262 1621 2263
rect 1634 2263 1640 2264
rect 1634 2262 1635 2263
rect 1620 2260 1635 2262
rect 1620 2259 1621 2260
rect 1615 2258 1621 2259
rect 1634 2259 1635 2260
rect 1639 2259 1640 2263
rect 1634 2258 1640 2259
rect 1642 2263 1648 2264
rect 1642 2259 1643 2263
rect 1647 2262 1648 2263
rect 1735 2263 1741 2264
rect 1735 2262 1736 2263
rect 1647 2260 1736 2262
rect 1647 2259 1648 2260
rect 1642 2258 1648 2259
rect 1735 2259 1736 2260
rect 1740 2259 1741 2263
rect 1735 2258 1741 2259
rect 1863 2263 1872 2264
rect 1863 2259 1864 2263
rect 1871 2259 1872 2263
rect 1863 2258 1872 2259
rect 1874 2263 1880 2264
rect 1874 2259 1875 2263
rect 1879 2262 1880 2263
rect 1967 2263 1973 2264
rect 1967 2262 1968 2263
rect 1879 2260 1968 2262
rect 1879 2259 1880 2260
rect 1874 2258 1880 2259
rect 1967 2259 1968 2260
rect 1972 2259 1973 2263
rect 2046 2260 2047 2264
rect 2051 2260 2052 2264
rect 2046 2259 2052 2260
rect 2070 2263 2076 2264
rect 2070 2259 2071 2263
rect 2075 2259 2076 2263
rect 1967 2258 1973 2259
rect 2070 2258 2076 2259
rect 2166 2263 2172 2264
rect 2166 2259 2167 2263
rect 2171 2259 2172 2263
rect 2166 2258 2172 2259
rect 2286 2263 2292 2264
rect 2286 2259 2287 2263
rect 2291 2259 2292 2263
rect 2286 2258 2292 2259
rect 2422 2263 2428 2264
rect 2422 2259 2423 2263
rect 2427 2259 2428 2263
rect 2422 2258 2428 2259
rect 2558 2263 2564 2264
rect 2558 2259 2559 2263
rect 2563 2259 2564 2263
rect 2558 2258 2564 2259
rect 1114 2255 1120 2256
rect 1114 2254 1115 2255
rect 936 2252 1115 2254
rect 479 2247 485 2248
rect 479 2243 480 2247
rect 484 2246 485 2247
rect 498 2247 504 2248
rect 498 2246 499 2247
rect 484 2244 499 2246
rect 484 2243 485 2244
rect 479 2242 485 2243
rect 498 2243 499 2244
rect 503 2243 504 2247
rect 498 2242 504 2243
rect 599 2247 605 2248
rect 599 2243 600 2247
rect 604 2246 605 2247
rect 618 2247 624 2248
rect 618 2246 619 2247
rect 604 2244 619 2246
rect 604 2243 605 2244
rect 599 2242 605 2243
rect 618 2243 619 2244
rect 623 2243 624 2247
rect 618 2242 624 2243
rect 735 2247 741 2248
rect 735 2243 736 2247
rect 740 2246 741 2247
rect 778 2247 784 2248
rect 778 2246 779 2247
rect 740 2244 779 2246
rect 740 2243 741 2244
rect 735 2242 741 2243
rect 778 2243 779 2244
rect 783 2243 784 2247
rect 778 2242 784 2243
rect 887 2247 893 2248
rect 887 2243 888 2247
rect 892 2246 893 2247
rect 936 2246 938 2252
rect 1114 2251 1115 2252
rect 1119 2251 1120 2255
rect 1114 2250 1120 2251
rect 2146 2255 2152 2256
rect 2146 2251 2147 2255
rect 2151 2251 2152 2255
rect 2146 2250 2152 2251
rect 2154 2255 2160 2256
rect 2154 2251 2155 2255
rect 2159 2254 2160 2255
rect 2498 2255 2504 2256
rect 2159 2252 2209 2254
rect 2159 2251 2160 2252
rect 2154 2250 2160 2251
rect 2362 2251 2368 2252
rect 892 2244 938 2246
rect 943 2247 949 2248
rect 892 2243 893 2244
rect 887 2242 893 2243
rect 943 2243 944 2247
rect 948 2246 949 2247
rect 1055 2247 1061 2248
rect 1055 2246 1056 2247
rect 948 2244 1056 2246
rect 948 2243 949 2244
rect 943 2242 949 2243
rect 1055 2243 1056 2244
rect 1060 2243 1061 2247
rect 1055 2242 1061 2243
rect 1066 2247 1072 2248
rect 1066 2243 1067 2247
rect 1071 2246 1072 2247
rect 1239 2247 1245 2248
rect 1239 2246 1240 2247
rect 1071 2244 1240 2246
rect 1071 2243 1072 2244
rect 1066 2242 1072 2243
rect 1239 2243 1240 2244
rect 1244 2243 1245 2247
rect 1239 2242 1245 2243
rect 1250 2247 1256 2248
rect 1250 2243 1251 2247
rect 1255 2246 1256 2247
rect 1431 2247 1437 2248
rect 1431 2246 1432 2247
rect 1255 2244 1432 2246
rect 1255 2243 1256 2244
rect 1250 2242 1256 2243
rect 1431 2243 1432 2244
rect 1436 2243 1437 2247
rect 1431 2242 1437 2243
rect 1631 2247 1637 2248
rect 1631 2243 1632 2247
rect 1636 2246 1637 2247
rect 1650 2247 1656 2248
rect 1650 2246 1651 2247
rect 1636 2244 1651 2246
rect 1636 2243 1637 2244
rect 1631 2242 1637 2243
rect 1650 2243 1651 2244
rect 1655 2243 1656 2247
rect 1650 2242 1656 2243
rect 1754 2247 1760 2248
rect 1754 2243 1755 2247
rect 1759 2246 1760 2247
rect 1831 2247 1837 2248
rect 1831 2246 1832 2247
rect 1759 2244 1832 2246
rect 1759 2243 1760 2244
rect 1754 2242 1760 2243
rect 1831 2243 1832 2244
rect 1836 2243 1837 2247
rect 1831 2242 1837 2243
rect 2046 2247 2052 2248
rect 2046 2243 2047 2247
rect 2051 2243 2052 2247
rect 2362 2247 2363 2251
rect 2367 2247 2368 2251
rect 2498 2251 2499 2255
rect 2503 2251 2504 2255
rect 2498 2250 2504 2251
rect 2634 2255 2640 2256
rect 2634 2251 2635 2255
rect 2639 2251 2640 2255
rect 2644 2254 2646 2268
rect 3942 2264 3948 2265
rect 2702 2263 2708 2264
rect 2702 2259 2703 2263
rect 2707 2259 2708 2263
rect 2702 2258 2708 2259
rect 2838 2263 2844 2264
rect 2838 2259 2839 2263
rect 2843 2259 2844 2263
rect 2838 2258 2844 2259
rect 2982 2263 2988 2264
rect 2982 2259 2983 2263
rect 2987 2259 2988 2263
rect 2982 2258 2988 2259
rect 3126 2263 3132 2264
rect 3126 2259 3127 2263
rect 3131 2259 3132 2263
rect 3126 2258 3132 2259
rect 3270 2263 3276 2264
rect 3270 2259 3271 2263
rect 3275 2259 3276 2263
rect 3942 2260 3943 2264
rect 3947 2260 3948 2264
rect 3942 2259 3948 2260
rect 3270 2258 3276 2259
rect 2914 2255 2920 2256
rect 2644 2252 2745 2254
rect 2634 2250 2640 2251
rect 2914 2251 2915 2255
rect 2919 2251 2920 2255
rect 2914 2250 2920 2251
rect 3058 2255 3064 2256
rect 3058 2251 3059 2255
rect 3063 2251 3064 2255
rect 3250 2255 3256 2256
rect 3250 2254 3251 2255
rect 3205 2252 3251 2254
rect 3058 2250 3064 2251
rect 3250 2251 3251 2252
rect 3255 2251 3256 2255
rect 3250 2250 3256 2251
rect 3258 2255 3264 2256
rect 3258 2251 3259 2255
rect 3263 2254 3264 2255
rect 3263 2252 3313 2254
rect 3263 2251 3264 2252
rect 3258 2250 3264 2251
rect 2362 2246 2368 2247
rect 3942 2247 3948 2248
rect 2046 2242 2052 2243
rect 2070 2244 2076 2245
rect 2070 2240 2071 2244
rect 2075 2240 2076 2244
rect 2070 2239 2076 2240
rect 2166 2244 2172 2245
rect 2166 2240 2167 2244
rect 2171 2240 2172 2244
rect 2166 2239 2172 2240
rect 2286 2244 2292 2245
rect 2286 2240 2287 2244
rect 2291 2240 2292 2244
rect 2286 2239 2292 2240
rect 2422 2244 2428 2245
rect 2422 2240 2423 2244
rect 2427 2240 2428 2244
rect 2422 2239 2428 2240
rect 2558 2244 2564 2245
rect 2558 2240 2559 2244
rect 2563 2240 2564 2244
rect 2558 2239 2564 2240
rect 2702 2244 2708 2245
rect 2702 2240 2703 2244
rect 2707 2240 2708 2244
rect 2702 2239 2708 2240
rect 2838 2244 2844 2245
rect 2838 2240 2839 2244
rect 2843 2240 2844 2244
rect 2838 2239 2844 2240
rect 2982 2244 2988 2245
rect 2982 2240 2983 2244
rect 2987 2240 2988 2244
rect 2982 2239 2988 2240
rect 3126 2244 3132 2245
rect 3126 2240 3127 2244
rect 3131 2240 3132 2244
rect 3126 2239 3132 2240
rect 3270 2244 3276 2245
rect 3270 2240 3271 2244
rect 3275 2240 3276 2244
rect 3942 2243 3943 2247
rect 3947 2243 3948 2247
rect 3942 2242 3948 2243
rect 3270 2239 3276 2240
rect 110 2228 116 2229
rect 2006 2228 2012 2229
rect 110 2224 111 2228
rect 115 2224 116 2228
rect 110 2223 116 2224
rect 414 2227 420 2228
rect 414 2223 415 2227
rect 419 2223 420 2227
rect 414 2222 420 2223
rect 534 2227 540 2228
rect 534 2223 535 2227
rect 539 2223 540 2227
rect 534 2222 540 2223
rect 670 2227 676 2228
rect 670 2223 671 2227
rect 675 2223 676 2227
rect 670 2222 676 2223
rect 822 2227 828 2228
rect 822 2223 823 2227
rect 827 2223 828 2227
rect 822 2222 828 2223
rect 990 2227 996 2228
rect 990 2223 991 2227
rect 995 2223 996 2227
rect 990 2222 996 2223
rect 1174 2227 1180 2228
rect 1174 2223 1175 2227
rect 1179 2223 1180 2227
rect 1174 2222 1180 2223
rect 1366 2227 1372 2228
rect 1366 2223 1367 2227
rect 1371 2223 1372 2227
rect 1366 2222 1372 2223
rect 1566 2227 1572 2228
rect 1566 2223 1567 2227
rect 1571 2223 1572 2227
rect 1566 2222 1572 2223
rect 1766 2227 1772 2228
rect 1766 2223 1767 2227
rect 1771 2223 1772 2227
rect 2006 2224 2007 2228
rect 2011 2224 2012 2228
rect 2006 2223 2012 2224
rect 1766 2222 1772 2223
rect 490 2219 496 2220
rect 490 2215 491 2219
rect 495 2215 496 2219
rect 490 2214 496 2215
rect 498 2219 504 2220
rect 498 2215 499 2219
rect 503 2218 504 2219
rect 618 2219 624 2220
rect 503 2216 577 2218
rect 503 2215 504 2216
rect 498 2214 504 2215
rect 618 2215 619 2219
rect 623 2218 624 2219
rect 943 2219 949 2220
rect 943 2218 944 2219
rect 623 2216 713 2218
rect 901 2216 944 2218
rect 623 2215 624 2216
rect 618 2214 624 2215
rect 943 2215 944 2216
rect 948 2215 949 2219
rect 943 2214 949 2215
rect 1066 2219 1072 2220
rect 1066 2215 1067 2219
rect 1071 2215 1072 2219
rect 1066 2214 1072 2215
rect 1250 2219 1256 2220
rect 1250 2215 1251 2219
rect 1255 2215 1256 2219
rect 1250 2214 1256 2215
rect 1258 2219 1264 2220
rect 1258 2215 1259 2219
rect 1263 2218 1264 2219
rect 1642 2219 1648 2220
rect 1263 2216 1409 2218
rect 1263 2215 1264 2216
rect 1258 2214 1264 2215
rect 1642 2215 1643 2219
rect 1647 2215 1648 2219
rect 1642 2214 1648 2215
rect 1650 2219 1656 2220
rect 1650 2215 1651 2219
rect 1655 2218 1656 2219
rect 1655 2216 1809 2218
rect 1655 2215 1656 2216
rect 1650 2214 1656 2215
rect 110 2211 116 2212
rect 110 2207 111 2211
rect 115 2207 116 2211
rect 2006 2211 2012 2212
rect 110 2206 116 2207
rect 414 2208 420 2209
rect 414 2204 415 2208
rect 419 2204 420 2208
rect 414 2203 420 2204
rect 534 2208 540 2209
rect 534 2204 535 2208
rect 539 2204 540 2208
rect 534 2203 540 2204
rect 670 2208 676 2209
rect 670 2204 671 2208
rect 675 2204 676 2208
rect 670 2203 676 2204
rect 822 2208 828 2209
rect 822 2204 823 2208
rect 827 2204 828 2208
rect 822 2203 828 2204
rect 990 2208 996 2209
rect 990 2204 991 2208
rect 995 2204 996 2208
rect 990 2203 996 2204
rect 1174 2208 1180 2209
rect 1174 2204 1175 2208
rect 1179 2204 1180 2208
rect 1174 2203 1180 2204
rect 1366 2208 1372 2209
rect 1366 2204 1367 2208
rect 1371 2204 1372 2208
rect 1366 2203 1372 2204
rect 1566 2208 1572 2209
rect 1566 2204 1567 2208
rect 1571 2204 1572 2208
rect 1566 2203 1572 2204
rect 1766 2208 1772 2209
rect 1766 2204 1767 2208
rect 1771 2204 1772 2208
rect 2006 2207 2007 2211
rect 2011 2207 2012 2211
rect 2006 2206 2012 2207
rect 1766 2203 1772 2204
rect 2370 2191 2376 2192
rect 2370 2190 2371 2191
rect 2288 2188 2371 2190
rect 2070 2184 2076 2185
rect 2046 2181 2052 2182
rect 2046 2177 2047 2181
rect 2051 2177 2052 2181
rect 2070 2180 2071 2184
rect 2075 2180 2076 2184
rect 2070 2179 2076 2180
rect 2046 2176 2052 2177
rect 2288 2174 2290 2188
rect 2370 2187 2371 2188
rect 2375 2187 2376 2191
rect 2370 2186 2376 2187
rect 2294 2184 2300 2185
rect 2294 2180 2295 2184
rect 2299 2180 2300 2184
rect 2294 2179 2300 2180
rect 2502 2184 2508 2185
rect 2502 2180 2503 2184
rect 2507 2180 2508 2184
rect 2502 2179 2508 2180
rect 2686 2184 2692 2185
rect 2686 2180 2687 2184
rect 2691 2180 2692 2184
rect 2686 2179 2692 2180
rect 2862 2184 2868 2185
rect 2862 2180 2863 2184
rect 2867 2180 2868 2184
rect 2862 2179 2868 2180
rect 3022 2184 3028 2185
rect 3022 2180 3023 2184
rect 3027 2180 3028 2184
rect 3022 2179 3028 2180
rect 3174 2184 3180 2185
rect 3174 2180 3175 2184
rect 3179 2180 3180 2184
rect 3174 2179 3180 2180
rect 3318 2184 3324 2185
rect 3318 2180 3319 2184
rect 3323 2180 3324 2184
rect 3318 2179 3324 2180
rect 3470 2184 3476 2185
rect 3470 2180 3471 2184
rect 3475 2180 3476 2184
rect 3470 2179 3476 2180
rect 3942 2181 3948 2182
rect 3942 2177 3943 2181
rect 3947 2177 3948 2181
rect 3942 2176 3948 2177
rect 2149 2172 2290 2174
rect 2370 2175 2376 2176
rect 2370 2171 2371 2175
rect 2375 2171 2376 2175
rect 2370 2170 2376 2171
rect 2578 2175 2584 2176
rect 2578 2171 2579 2175
rect 2583 2171 2584 2175
rect 2578 2170 2584 2171
rect 2754 2175 2760 2176
rect 2754 2171 2755 2175
rect 2759 2171 2760 2175
rect 2754 2170 2760 2171
rect 2938 2175 2944 2176
rect 2938 2171 2939 2175
rect 2943 2171 2944 2175
rect 2938 2170 2944 2171
rect 3098 2175 3104 2176
rect 3098 2171 3099 2175
rect 3103 2171 3104 2175
rect 3098 2170 3104 2171
rect 3250 2175 3256 2176
rect 3250 2171 3251 2175
rect 3255 2171 3256 2175
rect 3250 2170 3256 2171
rect 3394 2175 3400 2176
rect 3394 2171 3395 2175
rect 3399 2171 3400 2175
rect 3394 2170 3400 2171
rect 3438 2175 3444 2176
rect 3438 2171 3439 2175
rect 3443 2174 3444 2175
rect 3443 2172 3513 2174
rect 3443 2171 3444 2172
rect 3438 2170 3444 2171
rect 2070 2165 2076 2166
rect 2046 2164 2052 2165
rect 2046 2160 2047 2164
rect 2051 2160 2052 2164
rect 2070 2161 2071 2165
rect 2075 2161 2076 2165
rect 2070 2160 2076 2161
rect 2294 2165 2300 2166
rect 2294 2161 2295 2165
rect 2299 2161 2300 2165
rect 2294 2160 2300 2161
rect 2502 2165 2508 2166
rect 2502 2161 2503 2165
rect 2507 2161 2508 2165
rect 2502 2160 2508 2161
rect 2686 2165 2692 2166
rect 2686 2161 2687 2165
rect 2691 2161 2692 2165
rect 2686 2160 2692 2161
rect 2862 2165 2868 2166
rect 2862 2161 2863 2165
rect 2867 2161 2868 2165
rect 2862 2160 2868 2161
rect 3022 2165 3028 2166
rect 3022 2161 3023 2165
rect 3027 2161 3028 2165
rect 3022 2160 3028 2161
rect 3174 2165 3180 2166
rect 3174 2161 3175 2165
rect 3179 2161 3180 2165
rect 3174 2160 3180 2161
rect 3318 2165 3324 2166
rect 3318 2161 3319 2165
rect 3323 2161 3324 2165
rect 3318 2160 3324 2161
rect 3470 2165 3476 2166
rect 3470 2161 3471 2165
rect 3475 2161 3476 2165
rect 3470 2160 3476 2161
rect 3942 2164 3948 2165
rect 3942 2160 3943 2164
rect 3947 2160 3948 2164
rect 2046 2159 2052 2160
rect 3942 2159 3948 2160
rect 3258 2151 3264 2152
rect 3258 2150 3259 2151
rect 2932 2148 3259 2150
rect 2932 2144 2934 2148
rect 3258 2147 3259 2148
rect 3263 2147 3264 2151
rect 3258 2146 3264 2147
rect 2135 2143 2141 2144
rect 134 2140 140 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 246 2140 252 2141
rect 246 2136 247 2140
rect 251 2136 252 2140
rect 246 2135 252 2136
rect 390 2140 396 2141
rect 390 2136 391 2140
rect 395 2136 396 2140
rect 390 2135 396 2136
rect 550 2140 556 2141
rect 550 2136 551 2140
rect 555 2136 556 2140
rect 550 2135 556 2136
rect 710 2140 716 2141
rect 710 2136 711 2140
rect 715 2136 716 2140
rect 710 2135 716 2136
rect 870 2140 876 2141
rect 870 2136 871 2140
rect 875 2136 876 2140
rect 870 2135 876 2136
rect 1030 2140 1036 2141
rect 1030 2136 1031 2140
rect 1035 2136 1036 2140
rect 1030 2135 1036 2136
rect 1190 2140 1196 2141
rect 1190 2136 1191 2140
rect 1195 2136 1196 2140
rect 1190 2135 1196 2136
rect 1350 2140 1356 2141
rect 1350 2136 1351 2140
rect 1355 2136 1356 2140
rect 1350 2135 1356 2136
rect 1510 2140 1516 2141
rect 1510 2136 1511 2140
rect 1515 2136 1516 2140
rect 1510 2135 1516 2136
rect 1678 2140 1684 2141
rect 1678 2136 1679 2140
rect 1683 2136 1684 2140
rect 2135 2139 2136 2143
rect 2140 2142 2141 2143
rect 2154 2143 2160 2144
rect 2154 2142 2155 2143
rect 2140 2140 2155 2142
rect 2140 2139 2141 2140
rect 2135 2138 2141 2139
rect 2154 2139 2155 2140
rect 2159 2139 2160 2143
rect 2154 2138 2160 2139
rect 2359 2143 2368 2144
rect 2359 2139 2360 2143
rect 2367 2139 2368 2143
rect 2359 2138 2368 2139
rect 2370 2143 2376 2144
rect 2370 2139 2371 2143
rect 2375 2142 2376 2143
rect 2567 2143 2573 2144
rect 2567 2142 2568 2143
rect 2375 2140 2568 2142
rect 2375 2139 2376 2140
rect 2370 2138 2376 2139
rect 2567 2139 2568 2140
rect 2572 2139 2573 2143
rect 2567 2138 2573 2139
rect 2578 2143 2584 2144
rect 2578 2139 2579 2143
rect 2583 2142 2584 2143
rect 2751 2143 2757 2144
rect 2751 2142 2752 2143
rect 2583 2140 2752 2142
rect 2583 2139 2584 2140
rect 2578 2138 2584 2139
rect 2751 2139 2752 2140
rect 2756 2139 2757 2143
rect 2751 2138 2757 2139
rect 2927 2143 2934 2144
rect 2927 2139 2928 2143
rect 2932 2140 2934 2143
rect 2938 2143 2944 2144
rect 2932 2139 2933 2140
rect 2927 2138 2933 2139
rect 2938 2139 2939 2143
rect 2943 2142 2944 2143
rect 3087 2143 3093 2144
rect 3087 2142 3088 2143
rect 2943 2140 3088 2142
rect 2943 2139 2944 2140
rect 2938 2138 2944 2139
rect 3087 2139 3088 2140
rect 3092 2139 3093 2143
rect 3087 2138 3093 2139
rect 3098 2143 3104 2144
rect 3098 2139 3099 2143
rect 3103 2142 3104 2143
rect 3239 2143 3245 2144
rect 3239 2142 3240 2143
rect 3103 2140 3240 2142
rect 3103 2139 3104 2140
rect 3098 2138 3104 2139
rect 3239 2139 3240 2140
rect 3244 2139 3245 2143
rect 3239 2138 3245 2139
rect 3250 2143 3256 2144
rect 3250 2139 3251 2143
rect 3255 2142 3256 2143
rect 3383 2143 3389 2144
rect 3383 2142 3384 2143
rect 3255 2140 3384 2142
rect 3255 2139 3256 2140
rect 3250 2138 3256 2139
rect 3383 2139 3384 2140
rect 3388 2139 3389 2143
rect 3383 2138 3389 2139
rect 3394 2143 3400 2144
rect 3394 2139 3395 2143
rect 3399 2142 3400 2143
rect 3535 2143 3541 2144
rect 3535 2142 3536 2143
rect 3399 2140 3536 2142
rect 3399 2139 3400 2140
rect 3394 2138 3400 2139
rect 3535 2139 3536 2140
rect 3540 2139 3541 2143
rect 3535 2138 3541 2139
rect 1678 2135 1684 2136
rect 2006 2137 2012 2138
rect 110 2132 116 2133
rect 2006 2133 2007 2137
rect 2011 2133 2012 2137
rect 2006 2132 2012 2133
rect 239 2131 245 2132
rect 239 2130 240 2131
rect 213 2128 240 2130
rect 239 2127 240 2128
rect 244 2127 245 2131
rect 239 2126 245 2127
rect 322 2131 328 2132
rect 322 2127 323 2131
rect 327 2127 328 2131
rect 322 2126 328 2127
rect 466 2131 472 2132
rect 466 2127 467 2131
rect 471 2127 472 2131
rect 466 2126 472 2127
rect 626 2131 632 2132
rect 626 2127 627 2131
rect 631 2127 632 2131
rect 626 2126 632 2127
rect 778 2131 784 2132
rect 778 2127 779 2131
rect 783 2127 784 2131
rect 778 2126 784 2127
rect 938 2131 944 2132
rect 938 2127 939 2131
rect 943 2127 944 2131
rect 938 2126 944 2127
rect 954 2131 960 2132
rect 954 2127 955 2131
rect 959 2130 960 2131
rect 1127 2131 1133 2132
rect 959 2128 1073 2130
rect 959 2127 960 2128
rect 954 2126 960 2127
rect 1127 2127 1128 2131
rect 1132 2130 1133 2131
rect 1426 2131 1432 2132
rect 1132 2128 1233 2130
rect 1132 2127 1133 2128
rect 1127 2126 1133 2127
rect 1426 2127 1427 2131
rect 1431 2127 1432 2131
rect 1426 2126 1432 2127
rect 1586 2131 1592 2132
rect 1586 2127 1587 2131
rect 1591 2127 1592 2131
rect 1586 2126 1592 2127
rect 1754 2131 1760 2132
rect 1754 2127 1755 2131
rect 1759 2127 1760 2131
rect 1754 2126 1760 2127
rect 134 2121 140 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 134 2117 135 2121
rect 139 2117 140 2121
rect 134 2116 140 2117
rect 246 2121 252 2122
rect 246 2117 247 2121
rect 251 2117 252 2121
rect 246 2116 252 2117
rect 390 2121 396 2122
rect 390 2117 391 2121
rect 395 2117 396 2121
rect 390 2116 396 2117
rect 550 2121 556 2122
rect 550 2117 551 2121
rect 555 2117 556 2121
rect 550 2116 556 2117
rect 710 2121 716 2122
rect 710 2117 711 2121
rect 715 2117 716 2121
rect 710 2116 716 2117
rect 870 2121 876 2122
rect 870 2117 871 2121
rect 875 2117 876 2121
rect 870 2116 876 2117
rect 1030 2121 1036 2122
rect 1030 2117 1031 2121
rect 1035 2117 1036 2121
rect 1030 2116 1036 2117
rect 1190 2121 1196 2122
rect 1190 2117 1191 2121
rect 1195 2117 1196 2121
rect 1190 2116 1196 2117
rect 1350 2121 1356 2122
rect 1350 2117 1351 2121
rect 1355 2117 1356 2121
rect 1350 2116 1356 2117
rect 1510 2121 1516 2122
rect 1510 2117 1511 2121
rect 1515 2117 1516 2121
rect 1510 2116 1516 2117
rect 1678 2121 1684 2122
rect 1678 2117 1679 2121
rect 1683 2117 1684 2121
rect 1678 2116 1684 2117
rect 2006 2120 2012 2121
rect 2006 2116 2007 2120
rect 2011 2116 2012 2120
rect 110 2115 116 2116
rect 2006 2115 2012 2116
rect 2463 2107 2469 2108
rect 2463 2103 2464 2107
rect 2468 2103 2469 2107
rect 2463 2102 2469 2103
rect 2474 2107 2480 2108
rect 2474 2103 2475 2107
rect 2479 2106 2480 2107
rect 2559 2107 2565 2108
rect 2559 2106 2560 2107
rect 2479 2104 2560 2106
rect 2479 2103 2480 2104
rect 2474 2102 2480 2103
rect 2559 2103 2560 2104
rect 2564 2103 2565 2107
rect 2559 2102 2565 2103
rect 2570 2107 2576 2108
rect 2570 2103 2571 2107
rect 2575 2106 2576 2107
rect 2655 2107 2661 2108
rect 2655 2106 2656 2107
rect 2575 2104 2656 2106
rect 2575 2103 2576 2104
rect 2570 2102 2576 2103
rect 2655 2103 2656 2104
rect 2660 2103 2661 2107
rect 2655 2102 2661 2103
rect 2751 2107 2760 2108
rect 2751 2103 2752 2107
rect 2759 2103 2760 2107
rect 2847 2107 2853 2108
rect 2847 2106 2848 2107
rect 2751 2102 2760 2103
rect 2839 2104 2848 2106
rect 199 2099 205 2100
rect 199 2095 200 2099
rect 204 2098 205 2099
rect 210 2099 216 2100
rect 210 2098 211 2099
rect 204 2096 211 2098
rect 204 2095 205 2096
rect 199 2094 205 2095
rect 210 2095 211 2096
rect 215 2095 216 2099
rect 210 2094 216 2095
rect 239 2099 245 2100
rect 239 2095 240 2099
rect 244 2098 245 2099
rect 311 2099 317 2100
rect 311 2098 312 2099
rect 244 2096 312 2098
rect 244 2095 245 2096
rect 239 2094 245 2095
rect 311 2095 312 2096
rect 316 2095 317 2099
rect 311 2094 317 2095
rect 322 2099 328 2100
rect 322 2095 323 2099
rect 327 2098 328 2099
rect 455 2099 461 2100
rect 455 2098 456 2099
rect 327 2096 456 2098
rect 327 2095 328 2096
rect 322 2094 328 2095
rect 455 2095 456 2096
rect 460 2095 461 2099
rect 455 2094 461 2095
rect 466 2099 472 2100
rect 466 2095 467 2099
rect 471 2098 472 2099
rect 615 2099 621 2100
rect 615 2098 616 2099
rect 471 2096 616 2098
rect 471 2095 472 2096
rect 466 2094 472 2095
rect 615 2095 616 2096
rect 620 2095 621 2099
rect 615 2094 621 2095
rect 626 2099 632 2100
rect 626 2095 627 2099
rect 631 2098 632 2099
rect 775 2099 781 2100
rect 775 2098 776 2099
rect 631 2096 776 2098
rect 631 2095 632 2096
rect 626 2094 632 2095
rect 775 2095 776 2096
rect 780 2095 781 2099
rect 775 2094 781 2095
rect 935 2099 941 2100
rect 935 2095 936 2099
rect 940 2098 941 2099
rect 954 2099 960 2100
rect 954 2098 955 2099
rect 940 2096 955 2098
rect 940 2095 941 2096
rect 935 2094 941 2095
rect 954 2095 955 2096
rect 959 2095 960 2099
rect 954 2094 960 2095
rect 1095 2099 1101 2100
rect 1095 2095 1096 2099
rect 1100 2098 1101 2099
rect 1127 2099 1133 2100
rect 1127 2098 1128 2099
rect 1100 2096 1128 2098
rect 1100 2095 1101 2096
rect 1095 2094 1101 2095
rect 1127 2095 1128 2096
rect 1132 2095 1133 2099
rect 1127 2094 1133 2095
rect 1255 2099 1264 2100
rect 1255 2095 1256 2099
rect 1263 2095 1264 2099
rect 1255 2094 1264 2095
rect 1415 2099 1421 2100
rect 1415 2095 1416 2099
rect 1420 2098 1421 2099
rect 1426 2099 1432 2100
rect 1420 2095 1422 2098
rect 1415 2094 1422 2095
rect 1426 2095 1427 2099
rect 1431 2098 1432 2099
rect 1575 2099 1581 2100
rect 1575 2098 1576 2099
rect 1431 2096 1576 2098
rect 1431 2095 1432 2096
rect 1426 2094 1432 2095
rect 1575 2095 1576 2096
rect 1580 2095 1581 2099
rect 1575 2094 1581 2095
rect 1586 2099 1592 2100
rect 1586 2095 1587 2099
rect 1591 2098 1592 2099
rect 1743 2099 1749 2100
rect 1743 2098 1744 2099
rect 1591 2096 1744 2098
rect 1591 2095 1592 2096
rect 1586 2094 1592 2095
rect 1743 2095 1744 2096
rect 1748 2095 1749 2099
rect 1743 2094 1749 2095
rect 2465 2094 2467 2102
rect 2666 2099 2672 2100
rect 2666 2095 2667 2099
rect 2671 2098 2672 2099
rect 2839 2098 2841 2104
rect 2847 2103 2848 2104
rect 2852 2103 2853 2107
rect 2847 2102 2853 2103
rect 2943 2107 2952 2108
rect 2943 2103 2944 2107
rect 2951 2103 2952 2107
rect 2943 2102 2952 2103
rect 2954 2107 2960 2108
rect 2954 2103 2955 2107
rect 2959 2106 2960 2107
rect 3039 2107 3045 2108
rect 3039 2106 3040 2107
rect 2959 2104 3040 2106
rect 2959 2103 2960 2104
rect 2954 2102 2960 2103
rect 3039 2103 3040 2104
rect 3044 2103 3045 2107
rect 3039 2102 3045 2103
rect 3050 2107 3056 2108
rect 3050 2103 3051 2107
rect 3055 2106 3056 2107
rect 3135 2107 3141 2108
rect 3135 2106 3136 2107
rect 3055 2104 3136 2106
rect 3055 2103 3056 2104
rect 3050 2102 3056 2103
rect 3135 2103 3136 2104
rect 3140 2103 3141 2107
rect 3135 2102 3141 2103
rect 3146 2107 3152 2108
rect 3146 2103 3147 2107
rect 3151 2106 3152 2107
rect 3231 2107 3237 2108
rect 3231 2106 3232 2107
rect 3151 2104 3232 2106
rect 3151 2103 3152 2104
rect 3146 2102 3152 2103
rect 3231 2103 3232 2104
rect 3236 2103 3237 2107
rect 3231 2102 3237 2103
rect 3242 2107 3248 2108
rect 3242 2103 3243 2107
rect 3247 2106 3248 2107
rect 3327 2107 3333 2108
rect 3327 2106 3328 2107
rect 3247 2104 3328 2106
rect 3247 2103 3248 2104
rect 3242 2102 3248 2103
rect 3327 2103 3328 2104
rect 3332 2103 3333 2107
rect 3327 2102 3333 2103
rect 3338 2107 3344 2108
rect 3338 2103 3339 2107
rect 3343 2106 3344 2107
rect 3423 2107 3429 2108
rect 3423 2106 3424 2107
rect 3343 2104 3424 2106
rect 3343 2103 3344 2104
rect 3338 2102 3344 2103
rect 3423 2103 3424 2104
rect 3428 2103 3429 2107
rect 3423 2102 3429 2103
rect 3434 2107 3440 2108
rect 3434 2103 3435 2107
rect 3439 2106 3440 2107
rect 3519 2107 3525 2108
rect 3519 2106 3520 2107
rect 3439 2104 3520 2106
rect 3439 2103 3440 2104
rect 3434 2102 3440 2103
rect 3519 2103 3520 2104
rect 3524 2103 3525 2107
rect 3519 2102 3525 2103
rect 3530 2107 3536 2108
rect 3530 2103 3531 2107
rect 3535 2106 3536 2107
rect 3615 2107 3621 2108
rect 3615 2106 3616 2107
rect 3535 2104 3616 2106
rect 3535 2103 3536 2104
rect 3530 2102 3536 2103
rect 3615 2103 3616 2104
rect 3620 2103 3621 2107
rect 3615 2102 3621 2103
rect 3626 2107 3632 2108
rect 3626 2103 3627 2107
rect 3631 2106 3632 2107
rect 3711 2107 3717 2108
rect 3711 2106 3712 2107
rect 3631 2104 3712 2106
rect 3631 2103 3632 2104
rect 3626 2102 3632 2103
rect 3711 2103 3712 2104
rect 3716 2103 3717 2107
rect 3711 2102 3717 2103
rect 3722 2107 3728 2108
rect 3722 2103 3723 2107
rect 3727 2106 3728 2107
rect 3807 2107 3813 2108
rect 3807 2106 3808 2107
rect 3727 2104 3808 2106
rect 3727 2103 3728 2104
rect 3722 2102 3728 2103
rect 3807 2103 3808 2104
rect 3812 2103 3813 2107
rect 3807 2102 3813 2103
rect 3818 2107 3824 2108
rect 3818 2103 3819 2107
rect 3823 2106 3824 2107
rect 3903 2107 3909 2108
rect 3903 2106 3904 2107
rect 3823 2104 3904 2106
rect 3823 2103 3824 2104
rect 3818 2102 3824 2103
rect 3903 2103 3904 2104
rect 3908 2103 3909 2107
rect 3903 2102 3909 2103
rect 2671 2096 2841 2098
rect 2671 2095 2672 2096
rect 2666 2094 2672 2095
rect 1420 2090 1422 2094
rect 2465 2092 2602 2094
rect 1487 2091 1493 2092
rect 1487 2090 1488 2091
rect 1420 2088 1488 2090
rect 1487 2087 1488 2088
rect 1492 2087 1493 2091
rect 2600 2090 2602 2092
rect 1487 2086 1493 2087
rect 2046 2088 2052 2089
rect 2600 2088 2678 2090
rect 3942 2088 3948 2089
rect 2046 2084 2047 2088
rect 2051 2084 2052 2088
rect 2046 2083 2052 2084
rect 2398 2087 2404 2088
rect 2398 2083 2399 2087
rect 2403 2083 2404 2087
rect 2398 2082 2404 2083
rect 2494 2087 2500 2088
rect 2494 2083 2495 2087
rect 2499 2083 2500 2087
rect 2494 2082 2500 2083
rect 2590 2087 2596 2088
rect 2590 2083 2591 2087
rect 2595 2083 2596 2087
rect 2590 2082 2596 2083
rect 199 2079 205 2080
rect 199 2075 200 2079
rect 204 2078 205 2079
rect 218 2079 224 2080
rect 218 2078 219 2079
rect 204 2076 219 2078
rect 204 2075 205 2076
rect 199 2074 205 2075
rect 218 2075 219 2076
rect 223 2075 224 2079
rect 218 2074 224 2075
rect 311 2079 317 2080
rect 311 2075 312 2079
rect 316 2078 317 2079
rect 378 2079 384 2080
rect 378 2078 379 2079
rect 316 2076 379 2078
rect 316 2075 317 2076
rect 311 2074 317 2075
rect 378 2075 379 2076
rect 383 2075 384 2079
rect 378 2074 384 2075
rect 463 2079 469 2080
rect 463 2075 464 2079
rect 468 2078 469 2079
rect 482 2079 488 2080
rect 482 2078 483 2079
rect 468 2076 483 2078
rect 468 2075 469 2076
rect 463 2074 469 2075
rect 482 2075 483 2076
rect 487 2075 488 2079
rect 482 2074 488 2075
rect 615 2079 621 2080
rect 615 2075 616 2079
rect 620 2078 621 2079
rect 634 2079 640 2080
rect 634 2078 635 2079
rect 620 2076 635 2078
rect 620 2075 621 2076
rect 615 2074 621 2075
rect 634 2075 635 2076
rect 639 2075 640 2079
rect 634 2074 640 2075
rect 767 2079 773 2080
rect 767 2075 768 2079
rect 772 2078 773 2079
rect 878 2079 884 2080
rect 878 2078 879 2079
rect 772 2076 879 2078
rect 772 2075 773 2076
rect 767 2074 773 2075
rect 878 2075 879 2076
rect 883 2075 884 2079
rect 878 2074 884 2075
rect 911 2079 917 2080
rect 911 2075 912 2079
rect 916 2078 917 2079
rect 938 2079 944 2080
rect 938 2078 939 2079
rect 916 2076 939 2078
rect 916 2075 917 2076
rect 911 2074 917 2075
rect 938 2075 939 2076
rect 943 2075 944 2079
rect 938 2074 944 2075
rect 970 2079 976 2080
rect 970 2075 971 2079
rect 975 2078 976 2079
rect 1055 2079 1061 2080
rect 1055 2078 1056 2079
rect 975 2076 1056 2078
rect 975 2075 976 2076
rect 970 2074 976 2075
rect 1055 2075 1056 2076
rect 1060 2075 1061 2079
rect 1055 2074 1061 2075
rect 1066 2079 1072 2080
rect 1066 2075 1067 2079
rect 1071 2078 1072 2079
rect 1191 2079 1197 2080
rect 1191 2078 1192 2079
rect 1071 2076 1192 2078
rect 1071 2075 1072 2076
rect 1066 2074 1072 2075
rect 1191 2075 1192 2076
rect 1196 2075 1197 2079
rect 1191 2074 1197 2075
rect 1202 2079 1208 2080
rect 1202 2075 1203 2079
rect 1207 2078 1208 2079
rect 1319 2079 1325 2080
rect 1319 2078 1320 2079
rect 1207 2076 1320 2078
rect 1207 2075 1208 2076
rect 1202 2074 1208 2075
rect 1319 2075 1320 2076
rect 1324 2075 1325 2079
rect 1319 2074 1325 2075
rect 1330 2079 1336 2080
rect 1330 2075 1331 2079
rect 1335 2078 1336 2079
rect 1447 2079 1453 2080
rect 1447 2078 1448 2079
rect 1335 2076 1448 2078
rect 1335 2075 1336 2076
rect 1330 2074 1336 2075
rect 1447 2075 1448 2076
rect 1452 2075 1453 2079
rect 1447 2074 1453 2075
rect 1458 2079 1464 2080
rect 1458 2075 1459 2079
rect 1463 2078 1464 2079
rect 1583 2079 1589 2080
rect 1583 2078 1584 2079
rect 1463 2076 1584 2078
rect 1463 2075 1464 2076
rect 1458 2074 1464 2075
rect 1583 2075 1584 2076
rect 1588 2075 1589 2079
rect 1583 2074 1589 2075
rect 2474 2079 2480 2080
rect 2474 2075 2475 2079
rect 2479 2075 2480 2079
rect 2474 2074 2480 2075
rect 2570 2079 2576 2080
rect 2570 2075 2571 2079
rect 2575 2075 2576 2079
rect 2570 2074 2576 2075
rect 2666 2079 2672 2080
rect 2666 2075 2667 2079
rect 2671 2075 2672 2079
rect 2676 2078 2678 2088
rect 2686 2087 2692 2088
rect 2686 2083 2687 2087
rect 2691 2083 2692 2087
rect 2686 2082 2692 2083
rect 2782 2087 2788 2088
rect 2782 2083 2783 2087
rect 2787 2083 2788 2087
rect 2782 2082 2788 2083
rect 2878 2087 2884 2088
rect 2878 2083 2879 2087
rect 2883 2083 2884 2087
rect 2878 2082 2884 2083
rect 2974 2087 2980 2088
rect 2974 2083 2975 2087
rect 2979 2083 2980 2087
rect 2974 2082 2980 2083
rect 3070 2087 3076 2088
rect 3070 2083 3071 2087
rect 3075 2083 3076 2087
rect 3070 2082 3076 2083
rect 3166 2087 3172 2088
rect 3166 2083 3167 2087
rect 3171 2083 3172 2087
rect 3166 2082 3172 2083
rect 3262 2087 3268 2088
rect 3262 2083 3263 2087
rect 3267 2083 3268 2087
rect 3262 2082 3268 2083
rect 3358 2087 3364 2088
rect 3358 2083 3359 2087
rect 3363 2083 3364 2087
rect 3358 2082 3364 2083
rect 3454 2087 3460 2088
rect 3454 2083 3455 2087
rect 3459 2083 3460 2087
rect 3454 2082 3460 2083
rect 3550 2087 3556 2088
rect 3550 2083 3551 2087
rect 3555 2083 3556 2087
rect 3550 2082 3556 2083
rect 3646 2087 3652 2088
rect 3646 2083 3647 2087
rect 3651 2083 3652 2087
rect 3646 2082 3652 2083
rect 3742 2087 3748 2088
rect 3742 2083 3743 2087
rect 3747 2083 3748 2087
rect 3742 2082 3748 2083
rect 3838 2087 3844 2088
rect 3838 2083 3839 2087
rect 3843 2083 3844 2087
rect 3942 2084 3943 2088
rect 3947 2084 3948 2088
rect 3942 2083 3948 2084
rect 3838 2082 3844 2083
rect 2954 2079 2960 2080
rect 2676 2076 2729 2078
rect 2666 2074 2672 2075
rect 2954 2075 2955 2079
rect 2959 2075 2960 2079
rect 2954 2074 2960 2075
rect 3050 2079 3056 2080
rect 3050 2075 3051 2079
rect 3055 2075 3056 2079
rect 3050 2074 3056 2075
rect 3146 2079 3152 2080
rect 3146 2075 3147 2079
rect 3151 2075 3152 2079
rect 3146 2074 3152 2075
rect 3242 2079 3248 2080
rect 3242 2075 3243 2079
rect 3247 2075 3248 2079
rect 3242 2074 3248 2075
rect 3338 2079 3344 2080
rect 3338 2075 3339 2079
rect 3343 2075 3344 2079
rect 3338 2074 3344 2075
rect 3434 2079 3440 2080
rect 3434 2075 3435 2079
rect 3439 2075 3440 2079
rect 3434 2074 3440 2075
rect 3530 2079 3536 2080
rect 3530 2075 3531 2079
rect 3535 2075 3536 2079
rect 3530 2074 3536 2075
rect 3626 2079 3632 2080
rect 3626 2075 3627 2079
rect 3631 2075 3632 2079
rect 3626 2074 3632 2075
rect 3722 2079 3728 2080
rect 3722 2075 3723 2079
rect 3727 2075 3728 2079
rect 3722 2074 3728 2075
rect 3818 2079 3824 2080
rect 3818 2075 3819 2079
rect 3823 2075 3824 2079
rect 3818 2074 3824 2075
rect 3914 2075 3920 2076
rect 2046 2071 2052 2072
rect 2046 2067 2047 2071
rect 2051 2067 2052 2071
rect 2046 2066 2052 2067
rect 2398 2068 2404 2069
rect 2398 2064 2399 2068
rect 2403 2064 2404 2068
rect 2398 2063 2404 2064
rect 2494 2068 2500 2069
rect 2494 2064 2495 2068
rect 2499 2064 2500 2068
rect 2494 2063 2500 2064
rect 2590 2068 2596 2069
rect 2590 2064 2591 2068
rect 2595 2064 2596 2068
rect 2590 2063 2596 2064
rect 2686 2068 2692 2069
rect 2686 2064 2687 2068
rect 2691 2064 2692 2068
rect 2686 2063 2692 2064
rect 2782 2068 2788 2069
rect 2782 2064 2783 2068
rect 2787 2064 2788 2068
rect 2782 2063 2788 2064
rect 110 2060 116 2061
rect 2006 2060 2012 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 134 2059 140 2060
rect 134 2055 135 2059
rect 139 2055 140 2059
rect 134 2054 140 2055
rect 246 2059 252 2060
rect 246 2055 247 2059
rect 251 2055 252 2059
rect 246 2054 252 2055
rect 398 2059 404 2060
rect 398 2055 399 2059
rect 403 2055 404 2059
rect 398 2054 404 2055
rect 550 2059 556 2060
rect 550 2055 551 2059
rect 555 2055 556 2059
rect 550 2054 556 2055
rect 702 2059 708 2060
rect 702 2055 703 2059
rect 707 2055 708 2059
rect 702 2054 708 2055
rect 846 2059 852 2060
rect 846 2055 847 2059
rect 851 2055 852 2059
rect 846 2054 852 2055
rect 990 2059 996 2060
rect 990 2055 991 2059
rect 995 2055 996 2059
rect 990 2054 996 2055
rect 1126 2059 1132 2060
rect 1126 2055 1127 2059
rect 1131 2055 1132 2059
rect 1126 2054 1132 2055
rect 1254 2059 1260 2060
rect 1254 2055 1255 2059
rect 1259 2055 1260 2059
rect 1254 2054 1260 2055
rect 1382 2059 1388 2060
rect 1382 2055 1383 2059
rect 1387 2055 1388 2059
rect 1382 2054 1388 2055
rect 1518 2059 1524 2060
rect 1518 2055 1519 2059
rect 1523 2055 1524 2059
rect 2006 2056 2007 2060
rect 2011 2056 2012 2060
rect 2860 2058 2862 2073
rect 3914 2071 3915 2075
rect 3919 2071 3920 2075
rect 3914 2070 3920 2071
rect 3942 2071 3948 2072
rect 2878 2068 2884 2069
rect 2878 2064 2879 2068
rect 2883 2064 2884 2068
rect 2878 2063 2884 2064
rect 2974 2068 2980 2069
rect 2974 2064 2975 2068
rect 2979 2064 2980 2068
rect 2974 2063 2980 2064
rect 3070 2068 3076 2069
rect 3070 2064 3071 2068
rect 3075 2064 3076 2068
rect 3070 2063 3076 2064
rect 3166 2068 3172 2069
rect 3166 2064 3167 2068
rect 3171 2064 3172 2068
rect 3166 2063 3172 2064
rect 3262 2068 3268 2069
rect 3262 2064 3263 2068
rect 3267 2064 3268 2068
rect 3262 2063 3268 2064
rect 3358 2068 3364 2069
rect 3358 2064 3359 2068
rect 3363 2064 3364 2068
rect 3358 2063 3364 2064
rect 3454 2068 3460 2069
rect 3454 2064 3455 2068
rect 3459 2064 3460 2068
rect 3454 2063 3460 2064
rect 3550 2068 3556 2069
rect 3550 2064 3551 2068
rect 3555 2064 3556 2068
rect 3550 2063 3556 2064
rect 3646 2068 3652 2069
rect 3646 2064 3647 2068
rect 3651 2064 3652 2068
rect 3646 2063 3652 2064
rect 3742 2068 3748 2069
rect 3742 2064 3743 2068
rect 3747 2064 3748 2068
rect 3742 2063 3748 2064
rect 3838 2068 3844 2069
rect 3838 2064 3839 2068
rect 3843 2064 3844 2068
rect 3942 2067 3943 2071
rect 3947 2067 3948 2071
rect 3942 2066 3948 2067
rect 3838 2063 3844 2064
rect 2903 2059 2909 2060
rect 2903 2058 2904 2059
rect 2860 2056 2904 2058
rect 2006 2055 2012 2056
rect 2903 2055 2904 2056
rect 2908 2055 2909 2059
rect 1518 2054 1524 2055
rect 2903 2054 2909 2055
rect 210 2051 216 2052
rect 210 2047 211 2051
rect 215 2047 216 2051
rect 210 2046 216 2047
rect 218 2051 224 2052
rect 218 2047 219 2051
rect 223 2050 224 2051
rect 378 2051 384 2052
rect 223 2048 289 2050
rect 223 2047 224 2048
rect 218 2046 224 2047
rect 378 2047 379 2051
rect 383 2050 384 2051
rect 482 2051 488 2052
rect 383 2048 441 2050
rect 383 2047 384 2048
rect 378 2046 384 2047
rect 482 2047 483 2051
rect 487 2050 488 2051
rect 634 2051 640 2052
rect 487 2048 593 2050
rect 487 2047 488 2048
rect 482 2046 488 2047
rect 634 2047 635 2051
rect 639 2050 640 2051
rect 970 2051 976 2052
rect 970 2050 971 2051
rect 639 2048 745 2050
rect 925 2048 971 2050
rect 639 2047 640 2048
rect 634 2046 640 2047
rect 970 2047 971 2048
rect 975 2047 976 2051
rect 970 2046 976 2047
rect 1066 2051 1072 2052
rect 1066 2047 1067 2051
rect 1071 2047 1072 2051
rect 1066 2046 1072 2047
rect 1202 2051 1208 2052
rect 1202 2047 1203 2051
rect 1207 2047 1208 2051
rect 1202 2046 1208 2047
rect 1330 2051 1336 2052
rect 1330 2047 1331 2051
rect 1335 2047 1336 2051
rect 1330 2046 1336 2047
rect 1458 2051 1464 2052
rect 1458 2047 1459 2051
rect 1463 2047 1464 2051
rect 1458 2046 1464 2047
rect 1487 2051 1493 2052
rect 1487 2047 1488 2051
rect 1492 2050 1493 2051
rect 1492 2048 1561 2050
rect 1492 2047 1493 2048
rect 1487 2046 1493 2047
rect 110 2043 116 2044
rect 110 2039 111 2043
rect 115 2039 116 2043
rect 2006 2043 2012 2044
rect 110 2038 116 2039
rect 134 2040 140 2041
rect 134 2036 135 2040
rect 139 2036 140 2040
rect 134 2035 140 2036
rect 246 2040 252 2041
rect 246 2036 247 2040
rect 251 2036 252 2040
rect 246 2035 252 2036
rect 398 2040 404 2041
rect 398 2036 399 2040
rect 403 2036 404 2040
rect 398 2035 404 2036
rect 550 2040 556 2041
rect 550 2036 551 2040
rect 555 2036 556 2040
rect 550 2035 556 2036
rect 702 2040 708 2041
rect 702 2036 703 2040
rect 707 2036 708 2040
rect 702 2035 708 2036
rect 846 2040 852 2041
rect 846 2036 847 2040
rect 851 2036 852 2040
rect 846 2035 852 2036
rect 990 2040 996 2041
rect 990 2036 991 2040
rect 995 2036 996 2040
rect 990 2035 996 2036
rect 1126 2040 1132 2041
rect 1126 2036 1127 2040
rect 1131 2036 1132 2040
rect 1126 2035 1132 2036
rect 1254 2040 1260 2041
rect 1254 2036 1255 2040
rect 1259 2036 1260 2040
rect 1254 2035 1260 2036
rect 1382 2040 1388 2041
rect 1382 2036 1383 2040
rect 1387 2036 1388 2040
rect 1382 2035 1388 2036
rect 1518 2040 1524 2041
rect 1518 2036 1519 2040
rect 1523 2036 1524 2040
rect 2006 2039 2007 2043
rect 2011 2039 2012 2043
rect 2006 2038 2012 2039
rect 1518 2035 1524 2036
rect 2190 2008 2196 2009
rect 2046 2005 2052 2006
rect 2046 2001 2047 2005
rect 2051 2001 2052 2005
rect 2190 2004 2191 2008
rect 2195 2004 2196 2008
rect 2190 2003 2196 2004
rect 2398 2008 2404 2009
rect 2398 2004 2399 2008
rect 2403 2004 2404 2008
rect 2398 2003 2404 2004
rect 2646 2008 2652 2009
rect 2646 2004 2647 2008
rect 2651 2004 2652 2008
rect 2646 2003 2652 2004
rect 2918 2008 2924 2009
rect 2918 2004 2919 2008
rect 2923 2004 2924 2008
rect 2918 2003 2924 2004
rect 3214 2008 3220 2009
rect 3214 2004 3215 2008
rect 3219 2004 3220 2008
rect 3214 2003 3220 2004
rect 3526 2008 3532 2009
rect 3526 2004 3527 2008
rect 3531 2004 3532 2008
rect 3526 2003 3532 2004
rect 3838 2008 3844 2009
rect 3838 2004 3839 2008
rect 3843 2004 3844 2008
rect 3838 2003 3844 2004
rect 3942 2005 3948 2006
rect 2046 2000 2052 2001
rect 3942 2001 3943 2005
rect 3947 2001 3948 2005
rect 3942 2000 3948 2001
rect 2314 1999 2320 2000
rect 2314 1998 2315 1999
rect 2269 1996 2315 1998
rect 2314 1995 2315 1996
rect 2319 1995 2320 1999
rect 2314 1994 2320 1995
rect 2474 1999 2480 2000
rect 2474 1995 2475 1999
rect 2479 1995 2480 1999
rect 2474 1994 2480 1995
rect 2522 1999 2528 2000
rect 2522 1995 2523 1999
rect 2527 1998 2528 1999
rect 2994 1999 3000 2000
rect 2527 1996 2689 1998
rect 2527 1995 2528 1996
rect 2522 1994 2528 1995
rect 2994 1995 2995 1999
rect 2999 1995 3000 1999
rect 2994 1994 3000 1995
rect 3002 1999 3008 2000
rect 3002 1995 3003 1999
rect 3007 1998 3008 1999
rect 3610 1999 3616 2000
rect 3007 1996 3257 1998
rect 3007 1995 3008 1996
rect 3002 1994 3008 1995
rect 3604 1990 3606 1997
rect 3610 1995 3611 1999
rect 3615 1998 3616 1999
rect 3615 1996 3881 1998
rect 3615 1995 3616 1996
rect 3610 1994 3616 1995
rect 3791 1991 3797 1992
rect 3791 1990 3792 1991
rect 2190 1989 2196 1990
rect 2046 1988 2052 1989
rect 2046 1984 2047 1988
rect 2051 1984 2052 1988
rect 2190 1985 2191 1989
rect 2195 1985 2196 1989
rect 2190 1984 2196 1985
rect 2398 1989 2404 1990
rect 2398 1985 2399 1989
rect 2403 1985 2404 1989
rect 2398 1984 2404 1985
rect 2646 1989 2652 1990
rect 2646 1985 2647 1989
rect 2651 1985 2652 1989
rect 2646 1984 2652 1985
rect 2918 1989 2924 1990
rect 2918 1985 2919 1989
rect 2923 1985 2924 1989
rect 2918 1984 2924 1985
rect 3214 1989 3220 1990
rect 3214 1985 3215 1989
rect 3219 1985 3220 1989
rect 3214 1984 3220 1985
rect 3526 1989 3532 1990
rect 3526 1985 3527 1989
rect 3531 1985 3532 1989
rect 3604 1988 3792 1990
rect 3791 1987 3792 1988
rect 3796 1987 3797 1991
rect 3791 1986 3797 1987
rect 3838 1989 3844 1990
rect 3526 1984 3532 1985
rect 3838 1985 3839 1989
rect 3843 1985 3844 1989
rect 3838 1984 3844 1985
rect 3942 1988 3948 1989
rect 3942 1984 3943 1988
rect 3947 1984 3948 1988
rect 2046 1983 2052 1984
rect 3942 1983 3948 1984
rect 2522 1975 2528 1976
rect 2522 1974 2523 1975
rect 2308 1972 2523 1974
rect 2255 1967 2261 1968
rect 230 1964 236 1965
rect 110 1961 116 1962
rect 110 1957 111 1961
rect 115 1957 116 1961
rect 230 1960 231 1964
rect 235 1960 236 1964
rect 230 1959 236 1960
rect 390 1964 396 1965
rect 390 1960 391 1964
rect 395 1960 396 1964
rect 390 1959 396 1960
rect 566 1964 572 1965
rect 566 1960 567 1964
rect 571 1960 572 1964
rect 566 1959 572 1960
rect 750 1964 756 1965
rect 750 1960 751 1964
rect 755 1960 756 1964
rect 750 1959 756 1960
rect 942 1964 948 1965
rect 942 1960 943 1964
rect 947 1960 948 1964
rect 942 1959 948 1960
rect 1134 1964 1140 1965
rect 1134 1960 1135 1964
rect 1139 1960 1140 1964
rect 1134 1959 1140 1960
rect 1334 1964 1340 1965
rect 1334 1960 1335 1964
rect 1339 1960 1340 1964
rect 1334 1959 1340 1960
rect 1542 1964 1548 1965
rect 1542 1960 1543 1964
rect 1547 1960 1548 1964
rect 2255 1963 2256 1967
rect 2260 1966 2261 1967
rect 2308 1966 2310 1972
rect 2522 1971 2523 1972
rect 2527 1971 2528 1975
rect 3002 1975 3008 1976
rect 3002 1974 3003 1975
rect 2522 1970 2528 1971
rect 2839 1972 3003 1974
rect 2260 1964 2310 1966
rect 2314 1967 2320 1968
rect 2260 1963 2261 1964
rect 2255 1962 2261 1963
rect 2314 1963 2315 1967
rect 2319 1966 2320 1967
rect 2463 1967 2469 1968
rect 2463 1966 2464 1967
rect 2319 1964 2464 1966
rect 2319 1963 2320 1964
rect 2314 1962 2320 1963
rect 2463 1963 2464 1964
rect 2468 1963 2469 1967
rect 2463 1962 2469 1963
rect 2711 1967 2717 1968
rect 2711 1963 2712 1967
rect 2716 1966 2717 1967
rect 2839 1966 2841 1972
rect 3002 1971 3003 1972
rect 3007 1971 3008 1975
rect 3002 1970 3008 1971
rect 2716 1964 2841 1966
rect 2903 1967 2909 1968
rect 2716 1963 2717 1964
rect 2711 1962 2717 1963
rect 2903 1963 2904 1967
rect 2908 1966 2909 1967
rect 2983 1967 2989 1968
rect 2983 1966 2984 1967
rect 2908 1964 2984 1966
rect 2908 1963 2909 1964
rect 2903 1962 2909 1963
rect 2983 1963 2984 1964
rect 2988 1963 2989 1967
rect 2983 1962 2989 1963
rect 2994 1967 3000 1968
rect 2994 1963 2995 1967
rect 2999 1966 3000 1967
rect 3279 1967 3285 1968
rect 3279 1966 3280 1967
rect 2999 1964 3280 1966
rect 2999 1963 3000 1964
rect 2994 1962 3000 1963
rect 3279 1963 3280 1964
rect 3284 1963 3285 1967
rect 3279 1962 3285 1963
rect 3591 1967 3597 1968
rect 3591 1963 3592 1967
rect 3596 1966 3597 1967
rect 3610 1967 3616 1968
rect 3610 1966 3611 1967
rect 3596 1964 3611 1966
rect 3596 1963 3597 1964
rect 3591 1962 3597 1963
rect 3610 1963 3611 1964
rect 3615 1963 3616 1967
rect 3610 1962 3616 1963
rect 3903 1967 3909 1968
rect 3903 1963 3904 1967
rect 3908 1966 3909 1967
rect 3914 1967 3920 1968
rect 3914 1966 3915 1967
rect 3908 1964 3915 1966
rect 3908 1963 3909 1964
rect 3903 1962 3909 1963
rect 3914 1963 3915 1964
rect 3919 1963 3920 1967
rect 3914 1962 3920 1963
rect 1542 1959 1548 1960
rect 2006 1961 2012 1962
rect 110 1956 116 1957
rect 2006 1957 2007 1961
rect 2011 1957 2012 1961
rect 2006 1956 2012 1957
rect 314 1955 320 1956
rect 314 1954 315 1955
rect 309 1952 315 1954
rect 314 1951 315 1952
rect 319 1951 320 1955
rect 314 1950 320 1951
rect 466 1955 472 1956
rect 466 1951 467 1955
rect 471 1951 472 1955
rect 466 1950 472 1951
rect 642 1955 648 1956
rect 642 1951 643 1955
rect 647 1951 648 1955
rect 642 1950 648 1951
rect 826 1955 832 1956
rect 826 1951 827 1955
rect 831 1951 832 1955
rect 826 1950 832 1951
rect 878 1955 884 1956
rect 878 1951 879 1955
rect 883 1954 884 1955
rect 1210 1955 1216 1956
rect 883 1952 985 1954
rect 883 1951 884 1952
rect 878 1950 884 1951
rect 1210 1951 1211 1955
rect 1215 1951 1216 1955
rect 1210 1950 1216 1951
rect 1402 1955 1408 1956
rect 1402 1951 1403 1955
rect 1407 1951 1408 1955
rect 1402 1950 1408 1951
rect 1458 1955 1464 1956
rect 1458 1951 1459 1955
rect 1463 1954 1464 1955
rect 1463 1952 1585 1954
rect 1463 1951 1464 1952
rect 1458 1950 1464 1951
rect 230 1945 236 1946
rect 110 1944 116 1945
rect 110 1940 111 1944
rect 115 1940 116 1944
rect 230 1941 231 1945
rect 235 1941 236 1945
rect 230 1940 236 1941
rect 390 1945 396 1946
rect 390 1941 391 1945
rect 395 1941 396 1945
rect 390 1940 396 1941
rect 566 1945 572 1946
rect 566 1941 567 1945
rect 571 1941 572 1945
rect 566 1940 572 1941
rect 750 1945 756 1946
rect 750 1941 751 1945
rect 755 1941 756 1945
rect 750 1940 756 1941
rect 942 1945 948 1946
rect 942 1941 943 1945
rect 947 1941 948 1945
rect 942 1940 948 1941
rect 1134 1945 1140 1946
rect 1134 1941 1135 1945
rect 1139 1941 1140 1945
rect 1134 1940 1140 1941
rect 1334 1945 1340 1946
rect 1334 1941 1335 1945
rect 1339 1941 1340 1945
rect 1334 1940 1340 1941
rect 1542 1945 1548 1946
rect 1542 1941 1543 1945
rect 1547 1941 1548 1945
rect 1542 1940 1548 1941
rect 2006 1944 2012 1945
rect 2006 1940 2007 1944
rect 2011 1940 2012 1944
rect 110 1939 116 1940
rect 2006 1939 2012 1940
rect 2135 1943 2141 1944
rect 2135 1939 2136 1943
rect 2140 1939 2141 1943
rect 2135 1938 2141 1939
rect 2146 1943 2152 1944
rect 2146 1939 2147 1943
rect 2151 1942 2152 1943
rect 2303 1943 2309 1944
rect 2303 1942 2304 1943
rect 2151 1940 2304 1942
rect 2151 1939 2152 1940
rect 2146 1938 2152 1939
rect 2303 1939 2304 1940
rect 2308 1939 2309 1943
rect 2303 1938 2309 1939
rect 2474 1943 2480 1944
rect 2474 1939 2475 1943
rect 2479 1942 2480 1943
rect 2511 1943 2517 1944
rect 2511 1942 2512 1943
rect 2479 1940 2512 1942
rect 2479 1939 2480 1940
rect 2474 1938 2480 1939
rect 2511 1939 2512 1940
rect 2516 1939 2517 1943
rect 2511 1938 2517 1939
rect 2522 1943 2528 1944
rect 2522 1939 2523 1943
rect 2527 1942 2528 1943
rect 2735 1943 2741 1944
rect 2735 1942 2736 1943
rect 2527 1940 2736 1942
rect 2527 1939 2528 1940
rect 2522 1938 2528 1939
rect 2735 1939 2736 1940
rect 2740 1939 2741 1943
rect 2735 1938 2741 1939
rect 2746 1943 2752 1944
rect 2746 1939 2747 1943
rect 2751 1942 2752 1943
rect 2959 1943 2965 1944
rect 2959 1942 2960 1943
rect 2751 1940 2960 1942
rect 2751 1939 2752 1940
rect 2746 1938 2752 1939
rect 2959 1939 2960 1940
rect 2964 1939 2965 1943
rect 2959 1938 2965 1939
rect 3191 1943 3197 1944
rect 3191 1939 3192 1943
rect 3196 1942 3197 1943
rect 3215 1943 3221 1944
rect 3215 1942 3216 1943
rect 3196 1940 3216 1942
rect 3196 1939 3197 1940
rect 3191 1938 3197 1939
rect 3215 1939 3216 1940
rect 3220 1939 3221 1943
rect 3215 1938 3221 1939
rect 3423 1943 3429 1944
rect 3423 1939 3424 1943
rect 3428 1942 3429 1943
rect 3442 1943 3448 1944
rect 3442 1942 3443 1943
rect 3428 1940 3443 1942
rect 3428 1939 3429 1940
rect 3423 1938 3429 1939
rect 3442 1939 3443 1940
rect 3447 1939 3448 1943
rect 3442 1938 3448 1939
rect 3654 1943 3661 1944
rect 3654 1939 3655 1943
rect 3660 1939 3661 1943
rect 3654 1938 3661 1939
rect 3791 1943 3797 1944
rect 3791 1939 3792 1943
rect 3796 1942 3797 1943
rect 3895 1943 3901 1944
rect 3895 1942 3896 1943
rect 3796 1940 3896 1942
rect 3796 1939 3797 1940
rect 3791 1938 3797 1939
rect 3895 1939 3896 1940
rect 3900 1939 3901 1943
rect 3895 1938 3901 1939
rect 2137 1934 2139 1938
rect 2778 1935 2784 1936
rect 2778 1934 2779 1935
rect 2137 1932 2779 1934
rect 2778 1931 2779 1932
rect 2783 1931 2784 1935
rect 2778 1930 2784 1931
rect 2046 1924 2052 1925
rect 3942 1924 3948 1925
rect 295 1923 301 1924
rect 295 1919 296 1923
rect 300 1922 301 1923
rect 306 1923 312 1924
rect 306 1922 307 1923
rect 300 1920 307 1922
rect 300 1919 301 1920
rect 295 1918 301 1919
rect 306 1919 307 1920
rect 311 1919 312 1923
rect 306 1918 312 1919
rect 314 1923 320 1924
rect 314 1919 315 1923
rect 319 1922 320 1923
rect 455 1923 461 1924
rect 455 1922 456 1923
rect 319 1920 456 1922
rect 319 1919 320 1920
rect 314 1918 320 1919
rect 455 1919 456 1920
rect 460 1919 461 1923
rect 455 1918 461 1919
rect 466 1923 472 1924
rect 466 1919 467 1923
rect 471 1922 472 1923
rect 631 1923 637 1924
rect 631 1922 632 1923
rect 471 1920 632 1922
rect 471 1919 472 1920
rect 466 1918 472 1919
rect 631 1919 632 1920
rect 636 1919 637 1923
rect 631 1918 637 1919
rect 642 1923 648 1924
rect 642 1919 643 1923
rect 647 1922 648 1923
rect 815 1923 821 1924
rect 815 1922 816 1923
rect 647 1920 816 1922
rect 647 1919 648 1920
rect 642 1918 648 1919
rect 815 1919 816 1920
rect 820 1919 821 1923
rect 815 1918 821 1919
rect 826 1923 832 1924
rect 826 1919 827 1923
rect 831 1922 832 1923
rect 1007 1923 1013 1924
rect 1007 1922 1008 1923
rect 831 1920 1008 1922
rect 831 1919 832 1920
rect 826 1918 832 1919
rect 1007 1919 1008 1920
rect 1012 1919 1013 1923
rect 1007 1918 1013 1919
rect 1199 1923 1208 1924
rect 1199 1919 1200 1923
rect 1207 1919 1208 1923
rect 1199 1918 1208 1919
rect 1210 1923 1216 1924
rect 1210 1919 1211 1923
rect 1215 1922 1216 1923
rect 1399 1923 1405 1924
rect 1399 1922 1400 1923
rect 1215 1920 1400 1922
rect 1215 1919 1216 1920
rect 1210 1918 1216 1919
rect 1399 1919 1400 1920
rect 1404 1919 1405 1923
rect 1399 1918 1405 1919
rect 1530 1923 1536 1924
rect 1530 1919 1531 1923
rect 1535 1922 1536 1923
rect 1607 1923 1613 1924
rect 1607 1922 1608 1923
rect 1535 1920 1608 1922
rect 1535 1919 1536 1920
rect 1530 1918 1536 1919
rect 1607 1919 1608 1920
rect 1612 1919 1613 1923
rect 2046 1920 2047 1924
rect 2051 1920 2052 1924
rect 2046 1919 2052 1920
rect 2070 1923 2076 1924
rect 2070 1919 2071 1923
rect 2075 1919 2076 1923
rect 1607 1918 1613 1919
rect 2070 1918 2076 1919
rect 2238 1923 2244 1924
rect 2238 1919 2239 1923
rect 2243 1919 2244 1923
rect 2238 1918 2244 1919
rect 2446 1923 2452 1924
rect 2446 1919 2447 1923
rect 2451 1919 2452 1923
rect 2446 1918 2452 1919
rect 2670 1923 2676 1924
rect 2670 1919 2671 1923
rect 2675 1919 2676 1923
rect 2670 1918 2676 1919
rect 2894 1923 2900 1924
rect 2894 1919 2895 1923
rect 2899 1919 2900 1923
rect 2894 1918 2900 1919
rect 3126 1923 3132 1924
rect 3126 1919 3127 1923
rect 3131 1919 3132 1923
rect 3126 1918 3132 1919
rect 3358 1923 3364 1924
rect 3358 1919 3359 1923
rect 3363 1919 3364 1923
rect 3358 1918 3364 1919
rect 3590 1923 3596 1924
rect 3590 1919 3591 1923
rect 3595 1919 3596 1923
rect 3590 1918 3596 1919
rect 3830 1923 3836 1924
rect 3830 1919 3831 1923
rect 3835 1919 3836 1923
rect 3942 1920 3943 1924
rect 3947 1920 3948 1924
rect 3942 1919 3948 1920
rect 3830 1918 3836 1919
rect 2146 1915 2152 1916
rect 575 1911 581 1912
rect 575 1907 576 1911
rect 580 1910 581 1911
rect 594 1911 600 1912
rect 594 1910 595 1911
rect 580 1908 595 1910
rect 580 1907 581 1908
rect 575 1906 581 1907
rect 594 1907 595 1908
rect 599 1907 600 1911
rect 594 1906 600 1907
rect 687 1911 693 1912
rect 687 1907 688 1911
rect 692 1910 693 1911
rect 711 1911 717 1912
rect 711 1910 712 1911
rect 692 1908 712 1910
rect 692 1907 693 1908
rect 687 1906 693 1907
rect 711 1907 712 1908
rect 716 1907 717 1911
rect 711 1906 717 1907
rect 807 1911 813 1912
rect 807 1907 808 1911
rect 812 1910 813 1911
rect 831 1911 837 1912
rect 831 1910 832 1911
rect 812 1908 832 1910
rect 812 1907 813 1908
rect 807 1906 813 1907
rect 831 1907 832 1908
rect 836 1907 837 1911
rect 831 1906 837 1907
rect 927 1911 933 1912
rect 927 1907 928 1911
rect 932 1910 933 1911
rect 951 1911 957 1912
rect 951 1910 952 1911
rect 932 1908 952 1910
rect 932 1907 933 1908
rect 927 1906 933 1907
rect 951 1907 952 1908
rect 956 1907 957 1911
rect 951 1906 957 1907
rect 1047 1911 1053 1912
rect 1047 1907 1048 1911
rect 1052 1910 1053 1911
rect 1110 1911 1116 1912
rect 1110 1910 1111 1911
rect 1052 1908 1111 1910
rect 1052 1907 1053 1908
rect 1047 1906 1053 1907
rect 1110 1907 1111 1908
rect 1115 1907 1116 1911
rect 1110 1906 1116 1907
rect 1167 1911 1173 1912
rect 1167 1907 1168 1911
rect 1172 1910 1173 1911
rect 1190 1911 1196 1912
rect 1190 1910 1191 1911
rect 1172 1908 1191 1910
rect 1172 1907 1173 1908
rect 1167 1906 1173 1907
rect 1190 1907 1191 1908
rect 1195 1907 1196 1911
rect 1190 1906 1196 1907
rect 1287 1911 1293 1912
rect 1287 1907 1288 1911
rect 1292 1910 1293 1911
rect 1306 1911 1312 1912
rect 1306 1910 1307 1911
rect 1292 1908 1307 1910
rect 1292 1907 1293 1908
rect 1287 1906 1293 1907
rect 1306 1907 1307 1908
rect 1311 1907 1312 1911
rect 1306 1906 1312 1907
rect 1399 1911 1408 1912
rect 1399 1907 1400 1911
rect 1407 1907 1408 1911
rect 1399 1906 1408 1907
rect 1519 1911 1525 1912
rect 1519 1907 1520 1911
rect 1524 1910 1525 1911
rect 1543 1911 1549 1912
rect 1543 1910 1544 1911
rect 1524 1908 1544 1910
rect 1524 1907 1525 1908
rect 1519 1906 1525 1907
rect 1543 1907 1544 1908
rect 1548 1907 1549 1911
rect 1543 1906 1549 1907
rect 1639 1911 1645 1912
rect 1639 1907 1640 1911
rect 1644 1910 1645 1911
rect 1663 1911 1669 1912
rect 1663 1910 1664 1911
rect 1644 1908 1664 1910
rect 1644 1907 1645 1908
rect 1639 1906 1645 1907
rect 1663 1907 1664 1908
rect 1668 1907 1669 1911
rect 1663 1906 1669 1907
rect 1714 1911 1720 1912
rect 1714 1907 1715 1911
rect 1719 1910 1720 1911
rect 1759 1911 1765 1912
rect 1759 1910 1760 1911
rect 1719 1908 1760 1910
rect 1719 1907 1720 1908
rect 1714 1906 1720 1907
rect 1759 1907 1760 1908
rect 1764 1907 1765 1911
rect 2146 1911 2147 1915
rect 2151 1911 2152 1915
rect 2522 1915 2528 1916
rect 2146 1910 2152 1911
rect 2314 1911 2320 1912
rect 1759 1906 1765 1907
rect 2046 1907 2052 1908
rect 2046 1903 2047 1907
rect 2051 1903 2052 1907
rect 2314 1907 2315 1911
rect 2319 1907 2320 1911
rect 2522 1911 2523 1915
rect 2527 1911 2528 1915
rect 2522 1910 2528 1911
rect 2746 1915 2752 1916
rect 2746 1911 2747 1915
rect 2751 1911 2752 1915
rect 2746 1910 2752 1911
rect 2778 1915 2784 1916
rect 2778 1911 2779 1915
rect 2783 1914 2784 1915
rect 3031 1915 3037 1916
rect 2783 1912 2937 1914
rect 2783 1911 2784 1912
rect 2778 1910 2784 1911
rect 3031 1911 3032 1915
rect 3036 1914 3037 1915
rect 3215 1915 3221 1916
rect 3036 1912 3169 1914
rect 3036 1911 3037 1912
rect 3031 1910 3037 1911
rect 3215 1911 3216 1915
rect 3220 1914 3221 1915
rect 3442 1915 3448 1916
rect 3220 1912 3401 1914
rect 3220 1911 3221 1912
rect 3215 1910 3221 1911
rect 3442 1911 3443 1915
rect 3447 1914 3448 1915
rect 3447 1912 3633 1914
rect 3447 1911 3448 1912
rect 3442 1910 3448 1911
rect 3914 1911 3920 1912
rect 3914 1910 3915 1911
rect 3909 1908 3915 1910
rect 2314 1906 2320 1907
rect 3914 1907 3915 1908
rect 3919 1907 3920 1911
rect 3914 1906 3920 1907
rect 3942 1907 3948 1908
rect 2046 1902 2052 1903
rect 2070 1904 2076 1905
rect 2070 1900 2071 1904
rect 2075 1900 2076 1904
rect 2070 1899 2076 1900
rect 2238 1904 2244 1905
rect 2238 1900 2239 1904
rect 2243 1900 2244 1904
rect 2238 1899 2244 1900
rect 2446 1904 2452 1905
rect 2446 1900 2447 1904
rect 2451 1900 2452 1904
rect 2446 1899 2452 1900
rect 2670 1904 2676 1905
rect 2670 1900 2671 1904
rect 2675 1900 2676 1904
rect 2670 1899 2676 1900
rect 2894 1904 2900 1905
rect 2894 1900 2895 1904
rect 2899 1900 2900 1904
rect 2894 1899 2900 1900
rect 3126 1904 3132 1905
rect 3126 1900 3127 1904
rect 3131 1900 3132 1904
rect 3126 1899 3132 1900
rect 3358 1904 3364 1905
rect 3358 1900 3359 1904
rect 3363 1900 3364 1904
rect 3358 1899 3364 1900
rect 3590 1904 3596 1905
rect 3590 1900 3591 1904
rect 3595 1900 3596 1904
rect 3590 1899 3596 1900
rect 3830 1904 3836 1905
rect 3830 1900 3831 1904
rect 3835 1900 3836 1904
rect 3942 1903 3943 1907
rect 3947 1903 3948 1907
rect 3942 1902 3948 1903
rect 3830 1899 3836 1900
rect 110 1892 116 1893
rect 2006 1892 2012 1893
rect 110 1888 111 1892
rect 115 1888 116 1892
rect 110 1887 116 1888
rect 510 1891 516 1892
rect 510 1887 511 1891
rect 515 1887 516 1891
rect 510 1886 516 1887
rect 622 1891 628 1892
rect 622 1887 623 1891
rect 627 1887 628 1891
rect 622 1886 628 1887
rect 742 1891 748 1892
rect 742 1887 743 1891
rect 747 1887 748 1891
rect 742 1886 748 1887
rect 862 1891 868 1892
rect 862 1887 863 1891
rect 867 1887 868 1891
rect 862 1886 868 1887
rect 982 1891 988 1892
rect 982 1887 983 1891
rect 987 1887 988 1891
rect 982 1886 988 1887
rect 1102 1891 1108 1892
rect 1102 1887 1103 1891
rect 1107 1887 1108 1891
rect 1102 1886 1108 1887
rect 1222 1891 1228 1892
rect 1222 1887 1223 1891
rect 1227 1887 1228 1891
rect 1222 1886 1228 1887
rect 1334 1891 1340 1892
rect 1334 1887 1335 1891
rect 1339 1887 1340 1891
rect 1334 1886 1340 1887
rect 1454 1891 1460 1892
rect 1454 1887 1455 1891
rect 1459 1887 1460 1891
rect 1454 1886 1460 1887
rect 1574 1891 1580 1892
rect 1574 1887 1575 1891
rect 1579 1887 1580 1891
rect 1574 1886 1580 1887
rect 1694 1891 1700 1892
rect 1694 1887 1695 1891
rect 1699 1887 1700 1891
rect 2006 1888 2007 1892
rect 2011 1888 2012 1892
rect 2006 1887 2012 1888
rect 1694 1886 1700 1887
rect 306 1883 312 1884
rect 306 1879 307 1883
rect 311 1882 312 1883
rect 594 1883 600 1884
rect 311 1880 553 1882
rect 311 1879 312 1880
rect 306 1878 312 1879
rect 594 1879 595 1883
rect 599 1882 600 1883
rect 711 1883 717 1884
rect 599 1880 665 1882
rect 599 1879 600 1880
rect 594 1878 600 1879
rect 711 1879 712 1883
rect 716 1882 717 1883
rect 831 1883 837 1884
rect 716 1880 785 1882
rect 716 1879 717 1880
rect 711 1878 717 1879
rect 831 1879 832 1883
rect 836 1882 837 1883
rect 951 1883 957 1884
rect 836 1880 905 1882
rect 836 1879 837 1880
rect 831 1878 837 1879
rect 951 1879 952 1883
rect 956 1882 957 1883
rect 1190 1883 1196 1884
rect 956 1880 1025 1882
rect 956 1879 957 1880
rect 951 1878 957 1879
rect 1178 1879 1184 1880
rect 110 1875 116 1876
rect 110 1871 111 1875
rect 115 1871 116 1875
rect 1178 1875 1179 1879
rect 1183 1875 1184 1879
rect 1190 1879 1191 1883
rect 1195 1882 1196 1883
rect 1306 1883 1312 1884
rect 1195 1880 1265 1882
rect 1195 1879 1196 1880
rect 1190 1878 1196 1879
rect 1306 1879 1307 1883
rect 1311 1882 1312 1883
rect 1530 1883 1536 1884
rect 1311 1880 1377 1882
rect 1311 1879 1312 1880
rect 1306 1878 1312 1879
rect 1530 1879 1531 1883
rect 1535 1879 1536 1883
rect 1530 1878 1536 1879
rect 1543 1883 1549 1884
rect 1543 1879 1544 1883
rect 1548 1882 1549 1883
rect 1663 1883 1669 1884
rect 1548 1880 1617 1882
rect 1548 1879 1549 1880
rect 1543 1878 1549 1879
rect 1663 1879 1664 1883
rect 1668 1882 1669 1883
rect 1668 1880 1737 1882
rect 1668 1879 1669 1880
rect 1663 1878 1669 1879
rect 1178 1874 1184 1875
rect 2006 1875 2012 1876
rect 110 1870 116 1871
rect 510 1872 516 1873
rect 510 1868 511 1872
rect 515 1868 516 1872
rect 510 1867 516 1868
rect 622 1872 628 1873
rect 622 1868 623 1872
rect 627 1868 628 1872
rect 622 1867 628 1868
rect 742 1872 748 1873
rect 742 1868 743 1872
rect 747 1868 748 1872
rect 742 1867 748 1868
rect 862 1872 868 1873
rect 862 1868 863 1872
rect 867 1868 868 1872
rect 862 1867 868 1868
rect 982 1872 988 1873
rect 982 1868 983 1872
rect 987 1868 988 1872
rect 982 1867 988 1868
rect 1102 1872 1108 1873
rect 1102 1868 1103 1872
rect 1107 1868 1108 1872
rect 1102 1867 1108 1868
rect 1222 1872 1228 1873
rect 1222 1868 1223 1872
rect 1227 1868 1228 1872
rect 1222 1867 1228 1868
rect 1334 1872 1340 1873
rect 1334 1868 1335 1872
rect 1339 1868 1340 1872
rect 1334 1867 1340 1868
rect 1454 1872 1460 1873
rect 1454 1868 1455 1872
rect 1459 1868 1460 1872
rect 1454 1867 1460 1868
rect 1574 1872 1580 1873
rect 1574 1868 1575 1872
rect 1579 1868 1580 1872
rect 1574 1867 1580 1868
rect 1694 1872 1700 1873
rect 1694 1868 1695 1872
rect 1699 1868 1700 1872
rect 2006 1871 2007 1875
rect 2011 1871 2012 1875
rect 2006 1870 2012 1871
rect 1694 1867 1700 1868
rect 2070 1844 2076 1845
rect 2046 1841 2052 1842
rect 2046 1837 2047 1841
rect 2051 1837 2052 1841
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2070 1839 2076 1840
rect 2198 1844 2204 1845
rect 2198 1840 2199 1844
rect 2203 1840 2204 1844
rect 2198 1839 2204 1840
rect 2366 1844 2372 1845
rect 2366 1840 2367 1844
rect 2371 1840 2372 1844
rect 2366 1839 2372 1840
rect 2542 1844 2548 1845
rect 2542 1840 2543 1844
rect 2547 1840 2548 1844
rect 2542 1839 2548 1840
rect 2718 1844 2724 1845
rect 2718 1840 2719 1844
rect 2723 1840 2724 1844
rect 2718 1839 2724 1840
rect 2886 1844 2892 1845
rect 2886 1840 2887 1844
rect 2891 1840 2892 1844
rect 2886 1839 2892 1840
rect 3038 1844 3044 1845
rect 3038 1840 3039 1844
rect 3043 1840 3044 1844
rect 3038 1839 3044 1840
rect 3182 1844 3188 1845
rect 3182 1840 3183 1844
rect 3187 1840 3188 1844
rect 3182 1839 3188 1840
rect 3318 1844 3324 1845
rect 3318 1840 3319 1844
rect 3323 1840 3324 1844
rect 3318 1839 3324 1840
rect 3454 1844 3460 1845
rect 3454 1840 3455 1844
rect 3459 1840 3460 1844
rect 3454 1839 3460 1840
rect 3582 1844 3588 1845
rect 3582 1840 3583 1844
rect 3587 1840 3588 1844
rect 3582 1839 3588 1840
rect 3710 1844 3716 1845
rect 3710 1840 3711 1844
rect 3715 1840 3716 1844
rect 3710 1839 3716 1840
rect 3838 1844 3844 1845
rect 3838 1840 3839 1844
rect 3843 1840 3844 1844
rect 3838 1839 3844 1840
rect 3942 1841 3948 1842
rect 2046 1836 2052 1837
rect 3942 1837 3943 1841
rect 3947 1837 3948 1841
rect 3942 1836 3948 1837
rect 2138 1835 2144 1836
rect 2138 1831 2139 1835
rect 2143 1831 2144 1835
rect 2138 1830 2144 1831
rect 2154 1835 2160 1836
rect 2154 1831 2155 1835
rect 2159 1834 2160 1835
rect 2442 1835 2448 1836
rect 2159 1832 2241 1834
rect 2159 1831 2160 1832
rect 2154 1830 2160 1831
rect 2442 1831 2443 1835
rect 2447 1831 2448 1835
rect 2442 1830 2448 1831
rect 2618 1835 2624 1836
rect 2618 1831 2619 1835
rect 2623 1831 2624 1835
rect 2618 1830 2624 1831
rect 2658 1835 2664 1836
rect 2658 1831 2659 1835
rect 2663 1834 2664 1835
rect 2962 1835 2968 1836
rect 2663 1832 2761 1834
rect 2663 1831 2664 1832
rect 2658 1830 2664 1831
rect 2962 1831 2963 1835
rect 2967 1831 2968 1835
rect 2962 1830 2968 1831
rect 3114 1835 3120 1836
rect 3114 1831 3115 1835
rect 3119 1831 3120 1835
rect 3114 1830 3120 1831
rect 3258 1835 3264 1836
rect 3258 1831 3259 1835
rect 3263 1831 3264 1835
rect 3258 1830 3264 1831
rect 3394 1835 3400 1836
rect 3394 1831 3395 1835
rect 3399 1831 3400 1835
rect 3394 1830 3400 1831
rect 3522 1835 3528 1836
rect 3522 1831 3523 1835
rect 3527 1831 3528 1835
rect 3522 1830 3528 1831
rect 3654 1835 3660 1836
rect 3654 1831 3655 1835
rect 3659 1831 3660 1835
rect 3654 1830 3660 1831
rect 3666 1835 3672 1836
rect 3666 1831 3667 1835
rect 3671 1834 3672 1835
rect 3906 1835 3912 1836
rect 3671 1832 3753 1834
rect 3671 1831 3672 1832
rect 3666 1830 3672 1831
rect 3906 1831 3907 1835
rect 3911 1831 3912 1835
rect 3906 1830 3912 1831
rect 2070 1825 2076 1826
rect 2046 1824 2052 1825
rect 2046 1820 2047 1824
rect 2051 1820 2052 1824
rect 2070 1821 2071 1825
rect 2075 1821 2076 1825
rect 2070 1820 2076 1821
rect 2198 1825 2204 1826
rect 2198 1821 2199 1825
rect 2203 1821 2204 1825
rect 2198 1820 2204 1821
rect 2366 1825 2372 1826
rect 2366 1821 2367 1825
rect 2371 1821 2372 1825
rect 2366 1820 2372 1821
rect 2542 1825 2548 1826
rect 2542 1821 2543 1825
rect 2547 1821 2548 1825
rect 2542 1820 2548 1821
rect 2718 1825 2724 1826
rect 2718 1821 2719 1825
rect 2723 1821 2724 1825
rect 2718 1820 2724 1821
rect 2886 1825 2892 1826
rect 2886 1821 2887 1825
rect 2891 1821 2892 1825
rect 2886 1820 2892 1821
rect 3038 1825 3044 1826
rect 3038 1821 3039 1825
rect 3043 1821 3044 1825
rect 3038 1820 3044 1821
rect 3182 1825 3188 1826
rect 3182 1821 3183 1825
rect 3187 1821 3188 1825
rect 3182 1820 3188 1821
rect 3318 1825 3324 1826
rect 3318 1821 3319 1825
rect 3323 1821 3324 1825
rect 3318 1820 3324 1821
rect 3454 1825 3460 1826
rect 3454 1821 3455 1825
rect 3459 1821 3460 1825
rect 3454 1820 3460 1821
rect 3582 1825 3588 1826
rect 3582 1821 3583 1825
rect 3587 1821 3588 1825
rect 3582 1820 3588 1821
rect 3710 1825 3716 1826
rect 3710 1821 3711 1825
rect 3715 1821 3716 1825
rect 3710 1820 3716 1821
rect 3838 1825 3844 1826
rect 3838 1821 3839 1825
rect 3843 1821 3844 1825
rect 3838 1820 3844 1821
rect 3942 1824 3948 1825
rect 3942 1820 3943 1824
rect 3947 1820 3948 1824
rect 2046 1819 2052 1820
rect 3942 1819 3948 1820
rect 2658 1811 2664 1812
rect 2658 1810 2659 1811
rect 2265 1808 2659 1810
rect 614 1804 620 1805
rect 110 1801 116 1802
rect 110 1797 111 1801
rect 115 1797 116 1801
rect 614 1800 615 1804
rect 619 1800 620 1804
rect 614 1799 620 1800
rect 710 1804 716 1805
rect 710 1800 711 1804
rect 715 1800 716 1804
rect 710 1799 716 1800
rect 814 1804 820 1805
rect 814 1800 815 1804
rect 819 1800 820 1804
rect 814 1799 820 1800
rect 926 1804 932 1805
rect 926 1800 927 1804
rect 931 1800 932 1804
rect 926 1799 932 1800
rect 1038 1804 1044 1805
rect 1038 1800 1039 1804
rect 1043 1800 1044 1804
rect 1038 1799 1044 1800
rect 1158 1804 1164 1805
rect 1158 1800 1159 1804
rect 1163 1800 1164 1804
rect 1158 1799 1164 1800
rect 1278 1804 1284 1805
rect 1278 1800 1279 1804
rect 1283 1800 1284 1804
rect 1278 1799 1284 1800
rect 1398 1804 1404 1805
rect 1398 1800 1399 1804
rect 1403 1800 1404 1804
rect 1398 1799 1404 1800
rect 1518 1804 1524 1805
rect 1518 1800 1519 1804
rect 1523 1800 1524 1804
rect 1518 1799 1524 1800
rect 1638 1804 1644 1805
rect 2265 1804 2267 1808
rect 2658 1807 2659 1808
rect 2663 1807 2664 1811
rect 3031 1811 3037 1812
rect 3031 1810 3032 1811
rect 2658 1806 2664 1807
rect 2956 1808 3032 1810
rect 2956 1804 2958 1808
rect 3031 1807 3032 1808
rect 3036 1807 3037 1811
rect 3031 1806 3037 1807
rect 1638 1800 1639 1804
rect 1643 1800 1644 1804
rect 2135 1803 2141 1804
rect 1638 1799 1644 1800
rect 2006 1801 2012 1802
rect 110 1796 116 1797
rect 2006 1797 2007 1801
rect 2011 1797 2012 1801
rect 2135 1799 2136 1803
rect 2140 1802 2141 1803
rect 2154 1803 2160 1804
rect 2154 1802 2155 1803
rect 2140 1800 2155 1802
rect 2140 1799 2141 1800
rect 2135 1798 2141 1799
rect 2154 1799 2155 1800
rect 2159 1799 2160 1803
rect 2154 1798 2160 1799
rect 2263 1803 2269 1804
rect 2263 1799 2264 1803
rect 2268 1799 2269 1803
rect 2263 1798 2269 1799
rect 2314 1803 2320 1804
rect 2314 1799 2315 1803
rect 2319 1802 2320 1803
rect 2431 1803 2437 1804
rect 2431 1802 2432 1803
rect 2319 1800 2432 1802
rect 2319 1799 2320 1800
rect 2314 1798 2320 1799
rect 2431 1799 2432 1800
rect 2436 1799 2437 1803
rect 2431 1798 2437 1799
rect 2442 1803 2448 1804
rect 2442 1799 2443 1803
rect 2447 1802 2448 1803
rect 2607 1803 2613 1804
rect 2607 1802 2608 1803
rect 2447 1800 2608 1802
rect 2447 1799 2448 1800
rect 2442 1798 2448 1799
rect 2607 1799 2608 1800
rect 2612 1799 2613 1803
rect 2607 1798 2613 1799
rect 2618 1803 2624 1804
rect 2618 1799 2619 1803
rect 2623 1802 2624 1803
rect 2783 1803 2789 1804
rect 2783 1802 2784 1803
rect 2623 1800 2784 1802
rect 2623 1799 2624 1800
rect 2618 1798 2624 1799
rect 2783 1799 2784 1800
rect 2788 1799 2789 1803
rect 2783 1798 2789 1799
rect 2951 1803 2958 1804
rect 2951 1799 2952 1803
rect 2956 1800 2958 1803
rect 2962 1803 2968 1804
rect 2956 1799 2957 1800
rect 2951 1798 2957 1799
rect 2962 1799 2963 1803
rect 2967 1802 2968 1803
rect 3103 1803 3109 1804
rect 3103 1802 3104 1803
rect 2967 1800 3104 1802
rect 2967 1799 2968 1800
rect 2962 1798 2968 1799
rect 3103 1799 3104 1800
rect 3108 1799 3109 1803
rect 3103 1798 3109 1799
rect 3114 1803 3120 1804
rect 3114 1799 3115 1803
rect 3119 1802 3120 1803
rect 3247 1803 3253 1804
rect 3247 1802 3248 1803
rect 3119 1800 3248 1802
rect 3119 1799 3120 1800
rect 3114 1798 3120 1799
rect 3247 1799 3248 1800
rect 3252 1799 3253 1803
rect 3247 1798 3253 1799
rect 3258 1803 3264 1804
rect 3258 1799 3259 1803
rect 3263 1802 3264 1803
rect 3383 1803 3389 1804
rect 3383 1802 3384 1803
rect 3263 1800 3384 1802
rect 3263 1799 3264 1800
rect 3258 1798 3264 1799
rect 3383 1799 3384 1800
rect 3388 1799 3389 1803
rect 3383 1798 3389 1799
rect 3394 1803 3400 1804
rect 3394 1799 3395 1803
rect 3399 1802 3400 1803
rect 3519 1803 3525 1804
rect 3519 1802 3520 1803
rect 3399 1800 3520 1802
rect 3399 1799 3400 1800
rect 3394 1798 3400 1799
rect 3519 1799 3520 1800
rect 3524 1799 3525 1803
rect 3519 1798 3525 1799
rect 3647 1803 3653 1804
rect 3647 1799 3648 1803
rect 3652 1802 3653 1803
rect 3666 1803 3672 1804
rect 3666 1802 3667 1803
rect 3652 1800 3667 1802
rect 3652 1799 3653 1800
rect 3647 1798 3653 1799
rect 3666 1799 3667 1800
rect 3671 1799 3672 1803
rect 3666 1798 3672 1799
rect 3722 1803 3728 1804
rect 3722 1799 3723 1803
rect 3727 1802 3728 1803
rect 3775 1803 3781 1804
rect 3775 1802 3776 1803
rect 3727 1800 3776 1802
rect 3727 1799 3728 1800
rect 3722 1798 3728 1799
rect 3775 1799 3776 1800
rect 3780 1799 3781 1803
rect 3775 1798 3781 1799
rect 3903 1803 3909 1804
rect 3903 1799 3904 1803
rect 3908 1802 3909 1803
rect 3914 1803 3920 1804
rect 3914 1802 3915 1803
rect 3908 1800 3915 1802
rect 3908 1799 3909 1800
rect 3903 1798 3909 1799
rect 3914 1799 3915 1800
rect 3919 1799 3920 1803
rect 3914 1798 3920 1799
rect 2006 1796 2012 1797
rect 690 1795 696 1796
rect 690 1791 691 1795
rect 695 1791 696 1795
rect 690 1790 696 1791
rect 786 1795 792 1796
rect 786 1791 787 1795
rect 791 1791 792 1795
rect 786 1790 792 1791
rect 890 1795 896 1796
rect 890 1791 891 1795
rect 895 1791 896 1795
rect 890 1790 896 1791
rect 1002 1795 1008 1796
rect 1002 1791 1003 1795
rect 1007 1791 1008 1795
rect 1002 1790 1008 1791
rect 1110 1795 1116 1796
rect 1110 1791 1111 1795
rect 1115 1791 1116 1795
rect 1110 1790 1116 1791
rect 1234 1795 1240 1796
rect 1234 1791 1235 1795
rect 1239 1791 1240 1795
rect 1234 1790 1240 1791
rect 1354 1795 1360 1796
rect 1354 1791 1355 1795
rect 1359 1791 1360 1795
rect 1354 1790 1360 1791
rect 1390 1795 1396 1796
rect 1390 1791 1391 1795
rect 1395 1794 1396 1795
rect 1594 1795 1600 1796
rect 1395 1792 1441 1794
rect 1395 1791 1396 1792
rect 1390 1790 1396 1791
rect 1594 1791 1595 1795
rect 1599 1791 1600 1795
rect 1594 1790 1600 1791
rect 1714 1795 1720 1796
rect 1714 1791 1715 1795
rect 1719 1791 1720 1795
rect 1714 1790 1720 1791
rect 2135 1787 2144 1788
rect 614 1785 620 1786
rect 110 1784 116 1785
rect 110 1780 111 1784
rect 115 1780 116 1784
rect 614 1781 615 1785
rect 619 1781 620 1785
rect 614 1780 620 1781
rect 710 1785 716 1786
rect 710 1781 711 1785
rect 715 1781 716 1785
rect 710 1780 716 1781
rect 814 1785 820 1786
rect 814 1781 815 1785
rect 819 1781 820 1785
rect 814 1780 820 1781
rect 926 1785 932 1786
rect 926 1781 927 1785
rect 931 1781 932 1785
rect 926 1780 932 1781
rect 1038 1785 1044 1786
rect 1038 1781 1039 1785
rect 1043 1781 1044 1785
rect 1038 1780 1044 1781
rect 1158 1785 1164 1786
rect 1158 1781 1159 1785
rect 1163 1781 1164 1785
rect 1158 1780 1164 1781
rect 1278 1785 1284 1786
rect 1278 1781 1279 1785
rect 1283 1781 1284 1785
rect 1278 1780 1284 1781
rect 1398 1785 1404 1786
rect 1398 1781 1399 1785
rect 1403 1781 1404 1785
rect 1398 1780 1404 1781
rect 1518 1785 1524 1786
rect 1518 1781 1519 1785
rect 1523 1781 1524 1785
rect 1518 1780 1524 1781
rect 1638 1785 1644 1786
rect 1638 1781 1639 1785
rect 1643 1781 1644 1785
rect 1638 1780 1644 1781
rect 2006 1784 2012 1785
rect 2006 1780 2007 1784
rect 2011 1780 2012 1784
rect 2135 1783 2136 1787
rect 2143 1783 2144 1787
rect 2135 1782 2144 1783
rect 2146 1787 2152 1788
rect 2146 1783 2147 1787
rect 2151 1786 2152 1787
rect 2247 1787 2253 1788
rect 2247 1786 2248 1787
rect 2151 1784 2248 1786
rect 2151 1783 2152 1784
rect 2146 1782 2152 1783
rect 2247 1783 2248 1784
rect 2252 1783 2253 1787
rect 2247 1782 2253 1783
rect 2258 1787 2264 1788
rect 2258 1783 2259 1787
rect 2263 1786 2264 1787
rect 2391 1787 2397 1788
rect 2391 1786 2392 1787
rect 2263 1784 2392 1786
rect 2263 1783 2264 1784
rect 2258 1782 2264 1783
rect 2391 1783 2392 1784
rect 2396 1783 2397 1787
rect 2391 1782 2397 1783
rect 2402 1787 2408 1788
rect 2402 1783 2403 1787
rect 2407 1786 2408 1787
rect 2551 1787 2557 1788
rect 2551 1786 2552 1787
rect 2407 1784 2552 1786
rect 2407 1783 2408 1784
rect 2402 1782 2408 1783
rect 2551 1783 2552 1784
rect 2556 1783 2557 1787
rect 2551 1782 2557 1783
rect 2562 1787 2568 1788
rect 2562 1783 2563 1787
rect 2567 1786 2568 1787
rect 2719 1787 2725 1788
rect 2719 1786 2720 1787
rect 2567 1784 2720 1786
rect 2567 1783 2568 1784
rect 2562 1782 2568 1783
rect 2719 1783 2720 1784
rect 2724 1783 2725 1787
rect 2719 1782 2725 1783
rect 2895 1787 2901 1788
rect 2895 1783 2896 1787
rect 2900 1786 2901 1787
rect 2943 1787 2949 1788
rect 2943 1786 2944 1787
rect 2900 1784 2944 1786
rect 2900 1783 2901 1784
rect 2895 1782 2901 1783
rect 2943 1783 2944 1784
rect 2948 1783 2949 1787
rect 2943 1782 2949 1783
rect 3087 1787 3093 1788
rect 3087 1783 3088 1787
rect 3092 1786 3093 1787
rect 3106 1787 3112 1788
rect 3106 1786 3107 1787
rect 3092 1784 3107 1786
rect 3092 1783 3093 1784
rect 3087 1782 3093 1783
rect 3106 1783 3107 1784
rect 3111 1783 3112 1787
rect 3106 1782 3112 1783
rect 3287 1787 3293 1788
rect 3287 1783 3288 1787
rect 3292 1786 3293 1787
rect 3306 1787 3312 1788
rect 3306 1786 3307 1787
rect 3292 1784 3307 1786
rect 3292 1783 3293 1784
rect 3287 1782 3293 1783
rect 3306 1783 3307 1784
rect 3311 1783 3312 1787
rect 3306 1782 3312 1783
rect 3495 1787 3501 1788
rect 3495 1783 3496 1787
rect 3500 1786 3501 1787
rect 3522 1787 3528 1788
rect 3522 1786 3523 1787
rect 3500 1784 3523 1786
rect 3500 1783 3501 1784
rect 3495 1782 3501 1783
rect 3522 1783 3523 1784
rect 3527 1783 3528 1787
rect 3522 1782 3528 1783
rect 3711 1787 3717 1788
rect 3711 1783 3712 1787
rect 3716 1786 3717 1787
rect 3738 1787 3744 1788
rect 3738 1786 3739 1787
rect 3716 1784 3739 1786
rect 3716 1783 3717 1784
rect 3711 1782 3717 1783
rect 3738 1783 3739 1784
rect 3743 1783 3744 1787
rect 3738 1782 3744 1783
rect 3903 1787 3912 1788
rect 3903 1783 3904 1787
rect 3911 1783 3912 1787
rect 3903 1782 3912 1783
rect 110 1779 116 1780
rect 2006 1779 2012 1780
rect 2046 1768 2052 1769
rect 3942 1768 3948 1769
rect 2046 1764 2047 1768
rect 2051 1764 2052 1768
rect 679 1763 688 1764
rect 679 1759 680 1763
rect 687 1759 688 1763
rect 679 1758 688 1759
rect 690 1763 696 1764
rect 690 1759 691 1763
rect 695 1762 696 1763
rect 775 1763 781 1764
rect 775 1762 776 1763
rect 695 1760 776 1762
rect 695 1759 696 1760
rect 690 1758 696 1759
rect 775 1759 776 1760
rect 780 1759 781 1763
rect 775 1758 781 1759
rect 786 1763 792 1764
rect 786 1759 787 1763
rect 791 1762 792 1763
rect 879 1763 885 1764
rect 879 1762 880 1763
rect 791 1760 880 1762
rect 791 1759 792 1760
rect 786 1758 792 1759
rect 879 1759 880 1760
rect 884 1759 885 1763
rect 879 1758 885 1759
rect 890 1763 896 1764
rect 890 1759 891 1763
rect 895 1762 896 1763
rect 991 1763 997 1764
rect 991 1762 992 1763
rect 895 1760 992 1762
rect 895 1759 896 1760
rect 890 1758 896 1759
rect 991 1759 992 1760
rect 996 1759 997 1763
rect 991 1758 997 1759
rect 1002 1763 1008 1764
rect 1002 1759 1003 1763
rect 1007 1762 1008 1763
rect 1103 1763 1109 1764
rect 1103 1762 1104 1763
rect 1007 1760 1104 1762
rect 1007 1759 1008 1760
rect 1002 1758 1008 1759
rect 1103 1759 1104 1760
rect 1108 1759 1109 1763
rect 1103 1758 1109 1759
rect 1178 1763 1184 1764
rect 1178 1759 1179 1763
rect 1183 1762 1184 1763
rect 1223 1763 1229 1764
rect 1223 1762 1224 1763
rect 1183 1760 1224 1762
rect 1183 1759 1184 1760
rect 1178 1758 1184 1759
rect 1223 1759 1224 1760
rect 1228 1759 1229 1763
rect 1223 1758 1229 1759
rect 1234 1763 1240 1764
rect 1234 1759 1235 1763
rect 1239 1762 1240 1763
rect 1343 1763 1349 1764
rect 1343 1762 1344 1763
rect 1239 1760 1344 1762
rect 1239 1759 1240 1760
rect 1234 1758 1240 1759
rect 1343 1759 1344 1760
rect 1348 1759 1349 1763
rect 1343 1758 1349 1759
rect 1354 1763 1360 1764
rect 1354 1759 1355 1763
rect 1359 1762 1360 1763
rect 1463 1763 1469 1764
rect 1463 1762 1464 1763
rect 1359 1760 1464 1762
rect 1359 1759 1360 1760
rect 1354 1758 1360 1759
rect 1463 1759 1464 1760
rect 1468 1759 1469 1763
rect 1463 1758 1469 1759
rect 1583 1763 1592 1764
rect 1583 1759 1584 1763
rect 1591 1759 1592 1763
rect 1583 1758 1592 1759
rect 1594 1763 1600 1764
rect 1594 1759 1595 1763
rect 1599 1762 1600 1763
rect 1703 1763 1709 1764
rect 2046 1763 2052 1764
rect 2070 1767 2076 1768
rect 2070 1763 2071 1767
rect 2075 1763 2076 1767
rect 1703 1762 1704 1763
rect 1599 1760 1704 1762
rect 1599 1759 1600 1760
rect 1594 1758 1600 1759
rect 1703 1759 1704 1760
rect 1708 1759 1709 1763
rect 2070 1762 2076 1763
rect 2182 1767 2188 1768
rect 2182 1763 2183 1767
rect 2187 1763 2188 1767
rect 2182 1762 2188 1763
rect 2326 1767 2332 1768
rect 2326 1763 2327 1767
rect 2331 1763 2332 1767
rect 2326 1762 2332 1763
rect 2486 1767 2492 1768
rect 2486 1763 2487 1767
rect 2491 1763 2492 1767
rect 2486 1762 2492 1763
rect 2654 1767 2660 1768
rect 2654 1763 2655 1767
rect 2659 1763 2660 1767
rect 2654 1762 2660 1763
rect 2830 1767 2836 1768
rect 2830 1763 2831 1767
rect 2835 1763 2836 1767
rect 2830 1762 2836 1763
rect 3022 1767 3028 1768
rect 3022 1763 3023 1767
rect 3027 1763 3028 1767
rect 3022 1762 3028 1763
rect 3222 1767 3228 1768
rect 3222 1763 3223 1767
rect 3227 1763 3228 1767
rect 3222 1762 3228 1763
rect 3430 1767 3436 1768
rect 3430 1763 3431 1767
rect 3435 1763 3436 1767
rect 3430 1762 3436 1763
rect 3646 1767 3652 1768
rect 3646 1763 3647 1767
rect 3651 1763 3652 1767
rect 3646 1762 3652 1763
rect 3838 1767 3844 1768
rect 3838 1763 3839 1767
rect 3843 1763 3844 1767
rect 3942 1764 3943 1768
rect 3947 1764 3948 1768
rect 3942 1763 3948 1764
rect 3838 1762 3844 1763
rect 1703 1758 1709 1759
rect 2146 1759 2152 1760
rect 2146 1755 2147 1759
rect 2151 1755 2152 1759
rect 2146 1754 2152 1755
rect 2258 1759 2264 1760
rect 2258 1755 2259 1759
rect 2263 1755 2264 1759
rect 2258 1754 2264 1755
rect 2402 1759 2408 1760
rect 2402 1755 2403 1759
rect 2407 1755 2408 1759
rect 2402 1754 2408 1755
rect 2562 1759 2568 1760
rect 2562 1755 2563 1759
rect 2567 1755 2568 1759
rect 2562 1754 2568 1755
rect 2598 1759 2604 1760
rect 2598 1755 2599 1759
rect 2603 1758 2604 1759
rect 2943 1759 2949 1760
rect 2603 1756 2697 1758
rect 2603 1755 2604 1756
rect 2598 1754 2604 1755
rect 2906 1755 2912 1756
rect 431 1751 440 1752
rect 431 1747 432 1751
rect 439 1747 440 1751
rect 431 1746 440 1747
rect 442 1751 448 1752
rect 442 1747 443 1751
rect 447 1750 448 1751
rect 559 1751 565 1752
rect 559 1750 560 1751
rect 447 1748 560 1750
rect 447 1747 448 1748
rect 442 1746 448 1747
rect 559 1747 560 1748
rect 564 1747 565 1751
rect 559 1746 565 1747
rect 570 1751 576 1752
rect 570 1747 571 1751
rect 575 1750 576 1751
rect 703 1751 709 1752
rect 703 1750 704 1751
rect 575 1748 704 1750
rect 575 1747 576 1748
rect 570 1746 576 1747
rect 703 1747 704 1748
rect 708 1747 709 1751
rect 703 1746 709 1747
rect 770 1751 776 1752
rect 770 1747 771 1751
rect 775 1750 776 1751
rect 863 1751 869 1752
rect 863 1750 864 1751
rect 775 1748 864 1750
rect 775 1747 776 1748
rect 770 1746 776 1747
rect 863 1747 864 1748
rect 868 1747 869 1751
rect 863 1746 869 1747
rect 874 1751 880 1752
rect 874 1747 875 1751
rect 879 1750 880 1751
rect 1031 1751 1037 1752
rect 1031 1750 1032 1751
rect 879 1748 1032 1750
rect 879 1747 880 1748
rect 874 1746 880 1747
rect 1031 1747 1032 1748
rect 1036 1747 1037 1751
rect 1031 1746 1037 1747
rect 1207 1751 1213 1752
rect 1207 1747 1208 1751
rect 1212 1750 1213 1751
rect 1247 1751 1253 1752
rect 1247 1750 1248 1751
rect 1212 1748 1248 1750
rect 1212 1747 1213 1748
rect 1207 1746 1213 1747
rect 1247 1747 1248 1748
rect 1252 1747 1253 1751
rect 1247 1746 1253 1747
rect 1390 1751 1397 1752
rect 1390 1747 1391 1751
rect 1396 1747 1397 1751
rect 1390 1746 1397 1747
rect 1575 1751 1581 1752
rect 1575 1747 1576 1751
rect 1580 1750 1581 1751
rect 1662 1751 1668 1752
rect 1662 1750 1663 1751
rect 1580 1748 1663 1750
rect 1580 1747 1581 1748
rect 1575 1746 1581 1747
rect 1662 1747 1663 1748
rect 1667 1747 1668 1751
rect 1662 1746 1668 1747
rect 1758 1751 1764 1752
rect 1758 1747 1759 1751
rect 1763 1750 1764 1751
rect 1767 1751 1773 1752
rect 1767 1750 1768 1751
rect 1763 1748 1768 1750
rect 1763 1747 1764 1748
rect 1758 1746 1764 1747
rect 1767 1747 1768 1748
rect 1772 1747 1773 1751
rect 1767 1746 1773 1747
rect 2046 1751 2052 1752
rect 2046 1747 2047 1751
rect 2051 1747 2052 1751
rect 2906 1751 2907 1755
rect 2911 1751 2912 1755
rect 2943 1755 2944 1759
rect 2948 1758 2949 1759
rect 3106 1759 3112 1760
rect 2948 1756 3065 1758
rect 2948 1755 2949 1756
rect 2943 1754 2949 1755
rect 3106 1755 3107 1759
rect 3111 1758 3112 1759
rect 3306 1759 3312 1760
rect 3111 1756 3265 1758
rect 3111 1755 3112 1756
rect 3106 1754 3112 1755
rect 3306 1755 3307 1759
rect 3311 1758 3312 1759
rect 3722 1759 3728 1760
rect 3311 1756 3473 1758
rect 3311 1755 3312 1756
rect 3306 1754 3312 1755
rect 3722 1755 3723 1759
rect 3727 1755 3728 1759
rect 3722 1754 3728 1755
rect 2906 1750 2912 1751
rect 3906 1751 3912 1752
rect 2046 1746 2052 1747
rect 2070 1748 2076 1749
rect 2070 1744 2071 1748
rect 2075 1744 2076 1748
rect 2070 1743 2076 1744
rect 2182 1748 2188 1749
rect 2182 1744 2183 1748
rect 2187 1744 2188 1748
rect 2182 1743 2188 1744
rect 2326 1748 2332 1749
rect 2326 1744 2327 1748
rect 2331 1744 2332 1748
rect 2326 1743 2332 1744
rect 2486 1748 2492 1749
rect 2486 1744 2487 1748
rect 2491 1744 2492 1748
rect 2486 1743 2492 1744
rect 2654 1748 2660 1749
rect 2654 1744 2655 1748
rect 2659 1744 2660 1748
rect 2654 1743 2660 1744
rect 2830 1748 2836 1749
rect 2830 1744 2831 1748
rect 2835 1744 2836 1748
rect 2830 1743 2836 1744
rect 3022 1748 3028 1749
rect 3022 1744 3023 1748
rect 3027 1744 3028 1748
rect 3022 1743 3028 1744
rect 3222 1748 3228 1749
rect 3222 1744 3223 1748
rect 3227 1744 3228 1748
rect 3222 1743 3228 1744
rect 3430 1748 3436 1749
rect 3430 1744 3431 1748
rect 3435 1744 3436 1748
rect 3430 1743 3436 1744
rect 3646 1748 3652 1749
rect 3646 1744 3647 1748
rect 3651 1744 3652 1748
rect 3646 1743 3652 1744
rect 3838 1748 3844 1749
rect 3838 1744 3839 1748
rect 3843 1744 3844 1748
rect 3906 1747 3907 1751
rect 3911 1750 3912 1751
rect 3916 1750 3918 1753
rect 3911 1748 3918 1750
rect 3942 1751 3948 1752
rect 3911 1747 3912 1748
rect 3906 1746 3912 1747
rect 3942 1747 3943 1751
rect 3947 1747 3948 1751
rect 3942 1746 3948 1747
rect 3838 1743 3844 1744
rect 110 1732 116 1733
rect 2006 1732 2012 1733
rect 110 1728 111 1732
rect 115 1728 116 1732
rect 110 1727 116 1728
rect 366 1731 372 1732
rect 366 1727 367 1731
rect 371 1727 372 1731
rect 366 1726 372 1727
rect 494 1731 500 1732
rect 494 1727 495 1731
rect 499 1727 500 1731
rect 494 1726 500 1727
rect 638 1731 644 1732
rect 638 1727 639 1731
rect 643 1727 644 1731
rect 638 1726 644 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 966 1731 972 1732
rect 966 1727 967 1731
rect 971 1727 972 1731
rect 966 1726 972 1727
rect 1142 1731 1148 1732
rect 1142 1727 1143 1731
rect 1147 1727 1148 1731
rect 1142 1726 1148 1727
rect 1326 1731 1332 1732
rect 1326 1727 1327 1731
rect 1331 1727 1332 1731
rect 1326 1726 1332 1727
rect 1510 1731 1516 1732
rect 1510 1727 1511 1731
rect 1515 1727 1516 1731
rect 1510 1726 1516 1727
rect 1702 1731 1708 1732
rect 1702 1727 1703 1731
rect 1707 1727 1708 1731
rect 2006 1728 2007 1732
rect 2011 1728 2012 1732
rect 2006 1727 2012 1728
rect 1702 1726 1708 1727
rect 442 1723 448 1724
rect 442 1719 443 1723
rect 447 1719 448 1723
rect 442 1718 448 1719
rect 570 1723 576 1724
rect 570 1719 571 1723
rect 575 1719 576 1723
rect 770 1723 776 1724
rect 770 1722 771 1723
rect 717 1720 771 1722
rect 570 1718 576 1719
rect 770 1719 771 1720
rect 775 1719 776 1723
rect 770 1718 776 1719
rect 874 1723 880 1724
rect 874 1719 875 1723
rect 879 1719 880 1723
rect 874 1718 880 1719
rect 918 1723 924 1724
rect 918 1719 919 1723
rect 923 1722 924 1723
rect 1054 1723 1060 1724
rect 923 1720 1009 1722
rect 923 1719 924 1720
rect 918 1718 924 1719
rect 1054 1719 1055 1723
rect 1059 1722 1060 1723
rect 1247 1723 1253 1724
rect 1059 1720 1185 1722
rect 1059 1719 1060 1720
rect 1054 1718 1060 1719
rect 1247 1719 1248 1723
rect 1252 1722 1253 1723
rect 1586 1723 1592 1724
rect 1252 1720 1369 1722
rect 1252 1719 1253 1720
rect 1247 1718 1253 1719
rect 1586 1719 1587 1723
rect 1591 1719 1592 1723
rect 1586 1718 1592 1719
rect 1662 1723 1668 1724
rect 1662 1719 1663 1723
rect 1667 1722 1668 1723
rect 1667 1720 1745 1722
rect 1667 1719 1668 1720
rect 1662 1718 1668 1719
rect 110 1715 116 1716
rect 110 1711 111 1715
rect 115 1711 116 1715
rect 2006 1715 2012 1716
rect 110 1710 116 1711
rect 366 1712 372 1713
rect 366 1708 367 1712
rect 371 1708 372 1712
rect 366 1707 372 1708
rect 494 1712 500 1713
rect 494 1708 495 1712
rect 499 1708 500 1712
rect 494 1707 500 1708
rect 638 1712 644 1713
rect 638 1708 639 1712
rect 643 1708 644 1712
rect 638 1707 644 1708
rect 798 1712 804 1713
rect 798 1708 799 1712
rect 803 1708 804 1712
rect 798 1707 804 1708
rect 966 1712 972 1713
rect 966 1708 967 1712
rect 971 1708 972 1712
rect 966 1707 972 1708
rect 1142 1712 1148 1713
rect 1142 1708 1143 1712
rect 1147 1708 1148 1712
rect 1142 1707 1148 1708
rect 1326 1712 1332 1713
rect 1326 1708 1327 1712
rect 1331 1708 1332 1712
rect 1326 1707 1332 1708
rect 1510 1712 1516 1713
rect 1510 1708 1511 1712
rect 1515 1708 1516 1712
rect 1510 1707 1516 1708
rect 1702 1712 1708 1713
rect 1702 1708 1703 1712
rect 1707 1708 1708 1712
rect 2006 1711 2007 1715
rect 2011 1711 2012 1715
rect 2006 1710 2012 1711
rect 1702 1707 1708 1708
rect 2222 1680 2228 1681
rect 2046 1677 2052 1678
rect 2046 1673 2047 1677
rect 2051 1673 2052 1677
rect 2222 1676 2223 1680
rect 2227 1676 2228 1680
rect 2222 1675 2228 1676
rect 2326 1680 2332 1681
rect 2326 1676 2327 1680
rect 2331 1676 2332 1680
rect 2326 1675 2332 1676
rect 2438 1680 2444 1681
rect 2438 1676 2439 1680
rect 2443 1676 2444 1680
rect 2438 1675 2444 1676
rect 2558 1680 2564 1681
rect 2558 1676 2559 1680
rect 2563 1676 2564 1680
rect 2558 1675 2564 1676
rect 2686 1680 2692 1681
rect 2686 1676 2687 1680
rect 2691 1676 2692 1680
rect 2686 1675 2692 1676
rect 2822 1680 2828 1681
rect 2822 1676 2823 1680
rect 2827 1676 2828 1680
rect 2822 1675 2828 1676
rect 2966 1680 2972 1681
rect 2966 1676 2967 1680
rect 2971 1676 2972 1680
rect 2966 1675 2972 1676
rect 3126 1680 3132 1681
rect 3126 1676 3127 1680
rect 3131 1676 3132 1680
rect 3126 1675 3132 1676
rect 3302 1680 3308 1681
rect 3302 1676 3303 1680
rect 3307 1676 3308 1680
rect 3302 1675 3308 1676
rect 3486 1680 3492 1681
rect 3486 1676 3487 1680
rect 3491 1676 3492 1680
rect 3486 1675 3492 1676
rect 3670 1680 3676 1681
rect 3670 1676 3671 1680
rect 3675 1676 3676 1680
rect 3670 1675 3676 1676
rect 3838 1680 3844 1681
rect 3838 1676 3839 1680
rect 3843 1676 3844 1680
rect 3838 1675 3844 1676
rect 3942 1677 3948 1678
rect 2046 1672 2052 1673
rect 3942 1673 3943 1677
rect 3947 1673 3948 1677
rect 3942 1672 3948 1673
rect 2298 1671 2304 1672
rect 2298 1667 2299 1671
rect 2303 1667 2304 1671
rect 2298 1666 2304 1667
rect 2402 1671 2408 1672
rect 2402 1667 2403 1671
rect 2407 1667 2408 1671
rect 2402 1666 2408 1667
rect 2514 1671 2520 1672
rect 2514 1667 2515 1671
rect 2519 1667 2520 1671
rect 2514 1666 2520 1667
rect 2634 1671 2640 1672
rect 2634 1667 2635 1671
rect 2639 1667 2640 1671
rect 2634 1666 2640 1667
rect 2658 1671 2664 1672
rect 2658 1667 2659 1671
rect 2663 1670 2664 1671
rect 2946 1671 2952 1672
rect 2946 1670 2947 1671
rect 2663 1668 2729 1670
rect 2901 1668 2947 1670
rect 2663 1667 2664 1668
rect 2658 1666 2664 1667
rect 2946 1667 2947 1668
rect 2951 1667 2952 1671
rect 2946 1666 2952 1667
rect 3042 1671 3048 1672
rect 3042 1667 3043 1671
rect 3047 1667 3048 1671
rect 3042 1666 3048 1667
rect 3202 1671 3208 1672
rect 3202 1667 3203 1671
rect 3207 1667 3208 1671
rect 3202 1666 3208 1667
rect 3378 1671 3384 1672
rect 3378 1667 3379 1671
rect 3383 1667 3384 1671
rect 3378 1666 3384 1667
rect 3438 1671 3444 1672
rect 3438 1667 3439 1671
rect 3443 1670 3444 1671
rect 3738 1671 3744 1672
rect 3443 1668 3529 1670
rect 3443 1667 3444 1668
rect 3438 1666 3444 1667
rect 3738 1667 3739 1671
rect 3743 1667 3744 1671
rect 3738 1666 3744 1667
rect 3914 1671 3920 1672
rect 3914 1667 3915 1671
rect 3919 1667 3920 1671
rect 3914 1666 3920 1667
rect 2222 1661 2228 1662
rect 2046 1660 2052 1661
rect 2046 1656 2047 1660
rect 2051 1656 2052 1660
rect 2222 1657 2223 1661
rect 2227 1657 2228 1661
rect 2222 1656 2228 1657
rect 2326 1661 2332 1662
rect 2326 1657 2327 1661
rect 2331 1657 2332 1661
rect 2326 1656 2332 1657
rect 2438 1661 2444 1662
rect 2438 1657 2439 1661
rect 2443 1657 2444 1661
rect 2438 1656 2444 1657
rect 2558 1661 2564 1662
rect 2558 1657 2559 1661
rect 2563 1657 2564 1661
rect 2558 1656 2564 1657
rect 2686 1661 2692 1662
rect 2686 1657 2687 1661
rect 2691 1657 2692 1661
rect 2686 1656 2692 1657
rect 2822 1661 2828 1662
rect 2822 1657 2823 1661
rect 2827 1657 2828 1661
rect 2822 1656 2828 1657
rect 2966 1661 2972 1662
rect 2966 1657 2967 1661
rect 2971 1657 2972 1661
rect 2966 1656 2972 1657
rect 3126 1661 3132 1662
rect 3126 1657 3127 1661
rect 3131 1657 3132 1661
rect 3126 1656 3132 1657
rect 3302 1661 3308 1662
rect 3302 1657 3303 1661
rect 3307 1657 3308 1661
rect 3302 1656 3308 1657
rect 3486 1661 3492 1662
rect 3486 1657 3487 1661
rect 3491 1657 3492 1661
rect 3486 1656 3492 1657
rect 3670 1661 3676 1662
rect 3670 1657 3671 1661
rect 3675 1657 3676 1661
rect 3670 1656 3676 1657
rect 3838 1661 3844 1662
rect 3838 1657 3839 1661
rect 3843 1657 3844 1661
rect 3838 1656 3844 1657
rect 3942 1660 3948 1661
rect 3942 1656 3943 1660
rect 3947 1656 3948 1660
rect 434 1655 440 1656
rect 2046 1655 2052 1656
rect 3942 1655 3948 1656
rect 434 1651 435 1655
rect 439 1654 440 1655
rect 439 1652 654 1654
rect 439 1651 440 1652
rect 434 1650 440 1651
rect 134 1648 140 1649
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 134 1644 135 1648
rect 139 1644 140 1648
rect 134 1643 140 1644
rect 246 1648 252 1649
rect 246 1644 247 1648
rect 251 1644 252 1648
rect 246 1643 252 1644
rect 398 1648 404 1649
rect 398 1644 399 1648
rect 403 1644 404 1648
rect 398 1643 404 1644
rect 566 1648 572 1649
rect 566 1644 567 1648
rect 571 1644 572 1648
rect 566 1643 572 1644
rect 110 1640 116 1641
rect 239 1639 245 1640
rect 239 1638 240 1639
rect 213 1636 240 1638
rect 239 1635 240 1636
rect 244 1635 245 1639
rect 239 1634 245 1635
rect 322 1639 328 1640
rect 322 1635 323 1639
rect 327 1635 328 1639
rect 322 1634 328 1635
rect 474 1639 480 1640
rect 474 1635 475 1639
rect 479 1635 480 1639
rect 474 1634 480 1635
rect 642 1639 648 1640
rect 642 1635 643 1639
rect 647 1635 648 1639
rect 652 1638 654 1652
rect 742 1648 748 1649
rect 742 1644 743 1648
rect 747 1644 748 1648
rect 742 1643 748 1644
rect 934 1648 940 1649
rect 934 1644 935 1648
rect 939 1644 940 1648
rect 934 1643 940 1644
rect 1134 1648 1140 1649
rect 1134 1644 1135 1648
rect 1139 1644 1140 1648
rect 1134 1643 1140 1644
rect 1342 1648 1348 1649
rect 1342 1644 1343 1648
rect 1347 1644 1348 1648
rect 1342 1643 1348 1644
rect 1550 1648 1556 1649
rect 1550 1644 1551 1648
rect 1555 1644 1556 1648
rect 1550 1643 1556 1644
rect 1766 1648 1772 1649
rect 1766 1644 1767 1648
rect 1771 1644 1772 1648
rect 2598 1647 2604 1648
rect 2598 1646 2599 1647
rect 1766 1643 1772 1644
rect 2006 1645 2012 1646
rect 2006 1641 2007 1645
rect 2011 1641 2012 1645
rect 2006 1640 2012 1641
rect 2292 1644 2599 1646
rect 2292 1640 2294 1644
rect 2598 1643 2599 1644
rect 2603 1643 2604 1647
rect 2598 1642 2604 1643
rect 1010 1639 1016 1640
rect 652 1636 785 1638
rect 642 1634 648 1635
rect 1010 1635 1011 1639
rect 1015 1635 1016 1639
rect 1010 1634 1016 1635
rect 1210 1639 1216 1640
rect 1210 1635 1211 1639
rect 1215 1635 1216 1639
rect 1210 1634 1216 1635
rect 1410 1639 1416 1640
rect 1410 1635 1411 1639
rect 1415 1635 1416 1639
rect 1666 1639 1672 1640
rect 1666 1638 1667 1639
rect 1629 1636 1667 1638
rect 1410 1634 1416 1635
rect 1666 1635 1667 1636
rect 1671 1635 1672 1639
rect 1666 1634 1672 1635
rect 1758 1639 1764 1640
rect 1758 1635 1759 1639
rect 1763 1638 1764 1639
rect 2287 1639 2294 1640
rect 1763 1636 1809 1638
rect 1763 1635 1764 1636
rect 1758 1634 1764 1635
rect 2287 1635 2288 1639
rect 2292 1636 2294 1639
rect 2298 1639 2304 1640
rect 2292 1635 2293 1636
rect 2287 1634 2293 1635
rect 2298 1635 2299 1639
rect 2303 1638 2304 1639
rect 2391 1639 2397 1640
rect 2391 1638 2392 1639
rect 2303 1636 2392 1638
rect 2303 1635 2304 1636
rect 2298 1634 2304 1635
rect 2391 1635 2392 1636
rect 2396 1635 2397 1639
rect 2391 1634 2397 1635
rect 2402 1639 2408 1640
rect 2402 1635 2403 1639
rect 2407 1638 2408 1639
rect 2503 1639 2509 1640
rect 2503 1638 2504 1639
rect 2407 1636 2504 1638
rect 2407 1635 2408 1636
rect 2402 1634 2408 1635
rect 2503 1635 2504 1636
rect 2508 1635 2509 1639
rect 2503 1634 2509 1635
rect 2514 1639 2520 1640
rect 2514 1635 2515 1639
rect 2519 1638 2520 1639
rect 2623 1639 2629 1640
rect 2623 1638 2624 1639
rect 2519 1636 2624 1638
rect 2519 1635 2520 1636
rect 2514 1634 2520 1635
rect 2623 1635 2624 1636
rect 2628 1635 2629 1639
rect 2623 1634 2629 1635
rect 2634 1639 2640 1640
rect 2634 1635 2635 1639
rect 2639 1638 2640 1639
rect 2751 1639 2757 1640
rect 2751 1638 2752 1639
rect 2639 1636 2752 1638
rect 2639 1635 2640 1636
rect 2634 1634 2640 1635
rect 2751 1635 2752 1636
rect 2756 1635 2757 1639
rect 2751 1634 2757 1635
rect 2887 1639 2893 1640
rect 2887 1635 2888 1639
rect 2892 1638 2893 1639
rect 2906 1639 2912 1640
rect 2906 1638 2907 1639
rect 2892 1636 2907 1638
rect 2892 1635 2893 1636
rect 2887 1634 2893 1635
rect 2906 1635 2907 1636
rect 2911 1635 2912 1639
rect 2906 1634 2912 1635
rect 2946 1639 2952 1640
rect 2946 1635 2947 1639
rect 2951 1638 2952 1639
rect 3031 1639 3037 1640
rect 3031 1638 3032 1639
rect 2951 1636 3032 1638
rect 2951 1635 2952 1636
rect 2946 1634 2952 1635
rect 3031 1635 3032 1636
rect 3036 1635 3037 1639
rect 3031 1634 3037 1635
rect 3042 1639 3048 1640
rect 3042 1635 3043 1639
rect 3047 1638 3048 1639
rect 3191 1639 3197 1640
rect 3191 1638 3192 1639
rect 3047 1636 3192 1638
rect 3047 1635 3048 1636
rect 3042 1634 3048 1635
rect 3191 1635 3192 1636
rect 3196 1635 3197 1639
rect 3191 1634 3197 1635
rect 3202 1639 3208 1640
rect 3202 1635 3203 1639
rect 3207 1638 3208 1639
rect 3367 1639 3373 1640
rect 3367 1638 3368 1639
rect 3207 1636 3368 1638
rect 3207 1635 3208 1636
rect 3202 1634 3208 1635
rect 3367 1635 3368 1636
rect 3372 1635 3373 1639
rect 3367 1634 3373 1635
rect 3378 1639 3384 1640
rect 3378 1635 3379 1639
rect 3383 1638 3384 1639
rect 3551 1639 3557 1640
rect 3551 1638 3552 1639
rect 3383 1636 3552 1638
rect 3383 1635 3384 1636
rect 3378 1634 3384 1635
rect 3551 1635 3552 1636
rect 3556 1635 3557 1639
rect 3551 1634 3557 1635
rect 3735 1639 3741 1640
rect 3735 1635 3736 1639
rect 3740 1638 3741 1639
rect 3794 1639 3800 1640
rect 3794 1638 3795 1639
rect 3740 1636 3795 1638
rect 3740 1635 3741 1636
rect 3735 1634 3741 1635
rect 3794 1635 3795 1636
rect 3799 1635 3800 1639
rect 3794 1634 3800 1635
rect 3903 1639 3912 1640
rect 3903 1635 3904 1639
rect 3911 1635 3912 1639
rect 3903 1634 3912 1635
rect 2658 1631 2664 1632
rect 2658 1630 2659 1631
rect 134 1629 140 1630
rect 110 1628 116 1629
rect 110 1624 111 1628
rect 115 1624 116 1628
rect 134 1625 135 1629
rect 139 1625 140 1629
rect 134 1624 140 1625
rect 246 1629 252 1630
rect 246 1625 247 1629
rect 251 1625 252 1629
rect 246 1624 252 1625
rect 398 1629 404 1630
rect 398 1625 399 1629
rect 403 1625 404 1629
rect 398 1624 404 1625
rect 566 1629 572 1630
rect 566 1625 567 1629
rect 571 1625 572 1629
rect 566 1624 572 1625
rect 742 1629 748 1630
rect 742 1625 743 1629
rect 747 1625 748 1629
rect 742 1624 748 1625
rect 934 1629 940 1630
rect 934 1625 935 1629
rect 939 1625 940 1629
rect 934 1624 940 1625
rect 1134 1629 1140 1630
rect 1134 1625 1135 1629
rect 1139 1625 1140 1629
rect 1134 1624 1140 1625
rect 1342 1629 1348 1630
rect 1342 1625 1343 1629
rect 1347 1625 1348 1629
rect 1342 1624 1348 1625
rect 1550 1629 1556 1630
rect 1550 1625 1551 1629
rect 1555 1625 1556 1629
rect 1550 1624 1556 1625
rect 1766 1629 1772 1630
rect 1766 1625 1767 1629
rect 1771 1625 1772 1629
rect 1766 1624 1772 1625
rect 2006 1628 2012 1629
rect 2006 1624 2007 1628
rect 2011 1624 2012 1628
rect 2460 1628 2659 1630
rect 2460 1624 2462 1628
rect 2658 1627 2659 1628
rect 2663 1627 2664 1631
rect 3438 1631 3444 1632
rect 3438 1630 3439 1631
rect 2658 1626 2664 1627
rect 3044 1628 3439 1630
rect 3044 1624 3046 1628
rect 3438 1627 3439 1628
rect 3443 1627 3444 1631
rect 3438 1626 3444 1627
rect 110 1623 116 1624
rect 2006 1623 2012 1624
rect 2455 1623 2462 1624
rect 2455 1619 2456 1623
rect 2460 1620 2462 1623
rect 2466 1623 2472 1624
rect 2460 1619 2461 1620
rect 2455 1618 2461 1619
rect 2466 1619 2467 1623
rect 2471 1622 2472 1623
rect 2567 1623 2573 1624
rect 2567 1622 2568 1623
rect 2471 1620 2568 1622
rect 2471 1619 2472 1620
rect 2466 1618 2472 1619
rect 2567 1619 2568 1620
rect 2572 1619 2573 1623
rect 2567 1618 2573 1619
rect 2578 1623 2584 1624
rect 2578 1619 2579 1623
rect 2583 1622 2584 1623
rect 2679 1623 2685 1624
rect 2679 1622 2680 1623
rect 2583 1620 2680 1622
rect 2583 1619 2584 1620
rect 2578 1618 2584 1619
rect 2679 1619 2680 1620
rect 2684 1619 2685 1623
rect 2679 1618 2685 1619
rect 2726 1623 2732 1624
rect 2726 1619 2727 1623
rect 2731 1622 2732 1623
rect 2799 1623 2805 1624
rect 2799 1622 2800 1623
rect 2731 1620 2800 1622
rect 2731 1619 2732 1620
rect 2726 1618 2732 1619
rect 2799 1619 2800 1620
rect 2804 1619 2805 1623
rect 2799 1618 2805 1619
rect 2810 1623 2816 1624
rect 2810 1619 2811 1623
rect 2815 1622 2816 1623
rect 2919 1623 2925 1624
rect 2919 1622 2920 1623
rect 2815 1620 2920 1622
rect 2815 1619 2816 1620
rect 2810 1618 2816 1619
rect 2919 1619 2920 1620
rect 2924 1619 2925 1623
rect 2919 1618 2925 1619
rect 3039 1623 3046 1624
rect 3039 1619 3040 1623
rect 3044 1620 3046 1623
rect 3050 1623 3056 1624
rect 3044 1619 3045 1620
rect 3039 1618 3045 1619
rect 3050 1619 3051 1623
rect 3055 1622 3056 1623
rect 3159 1623 3165 1624
rect 3159 1622 3160 1623
rect 3055 1620 3160 1622
rect 3055 1619 3056 1620
rect 3050 1618 3056 1619
rect 3159 1619 3160 1620
rect 3164 1619 3165 1623
rect 3159 1618 3165 1619
rect 3170 1623 3176 1624
rect 3170 1619 3171 1623
rect 3175 1622 3176 1623
rect 3279 1623 3285 1624
rect 3279 1622 3280 1623
rect 3175 1620 3280 1622
rect 3175 1619 3176 1620
rect 3170 1618 3176 1619
rect 3279 1619 3280 1620
rect 3284 1619 3285 1623
rect 3279 1618 3285 1619
rect 3290 1623 3296 1624
rect 3290 1619 3291 1623
rect 3295 1622 3296 1623
rect 3399 1623 3405 1624
rect 3399 1622 3400 1623
rect 3295 1620 3400 1622
rect 3295 1619 3296 1620
rect 3290 1618 3296 1619
rect 3399 1619 3400 1620
rect 3404 1619 3405 1623
rect 3399 1618 3405 1619
rect 3410 1623 3416 1624
rect 3410 1619 3411 1623
rect 3415 1622 3416 1623
rect 3519 1623 3525 1624
rect 3519 1622 3520 1623
rect 3415 1620 3520 1622
rect 3415 1619 3416 1620
rect 3410 1618 3416 1619
rect 3519 1619 3520 1620
rect 3524 1619 3525 1623
rect 3519 1618 3525 1619
rect 1054 1615 1060 1616
rect 1054 1614 1055 1615
rect 1004 1612 1055 1614
rect 1004 1608 1006 1612
rect 1054 1611 1055 1612
rect 1059 1611 1060 1615
rect 1054 1610 1060 1611
rect 199 1607 205 1608
rect 199 1603 200 1607
rect 204 1606 205 1607
rect 210 1607 216 1608
rect 210 1606 211 1607
rect 204 1604 211 1606
rect 204 1603 205 1604
rect 199 1602 205 1603
rect 210 1603 211 1604
rect 215 1603 216 1607
rect 210 1602 216 1603
rect 239 1607 245 1608
rect 239 1603 240 1607
rect 244 1606 245 1607
rect 311 1607 317 1608
rect 311 1606 312 1607
rect 244 1604 312 1606
rect 244 1603 245 1604
rect 239 1602 245 1603
rect 311 1603 312 1604
rect 316 1603 317 1607
rect 311 1602 317 1603
rect 322 1607 328 1608
rect 322 1603 323 1607
rect 327 1606 328 1607
rect 463 1607 469 1608
rect 463 1606 464 1607
rect 327 1604 464 1606
rect 327 1603 328 1604
rect 322 1602 328 1603
rect 463 1603 464 1604
rect 468 1603 469 1607
rect 463 1602 469 1603
rect 474 1607 480 1608
rect 474 1603 475 1607
rect 479 1606 480 1607
rect 631 1607 637 1608
rect 631 1606 632 1607
rect 479 1604 632 1606
rect 479 1603 480 1604
rect 474 1602 480 1603
rect 631 1603 632 1604
rect 636 1603 637 1607
rect 631 1602 637 1603
rect 642 1607 648 1608
rect 642 1603 643 1607
rect 647 1606 648 1607
rect 807 1607 813 1608
rect 807 1606 808 1607
rect 647 1604 808 1606
rect 647 1603 648 1604
rect 642 1602 648 1603
rect 807 1603 808 1604
rect 812 1603 813 1607
rect 807 1602 813 1603
rect 999 1607 1006 1608
rect 999 1603 1000 1607
rect 1004 1604 1006 1607
rect 1010 1607 1016 1608
rect 1004 1603 1005 1604
rect 999 1602 1005 1603
rect 1010 1603 1011 1607
rect 1015 1606 1016 1607
rect 1199 1607 1205 1608
rect 1199 1606 1200 1607
rect 1015 1604 1200 1606
rect 1015 1603 1016 1604
rect 1010 1602 1016 1603
rect 1199 1603 1200 1604
rect 1204 1603 1205 1607
rect 1199 1602 1205 1603
rect 1210 1607 1216 1608
rect 1210 1603 1211 1607
rect 1215 1606 1216 1607
rect 1407 1607 1413 1608
rect 1407 1606 1408 1607
rect 1215 1604 1408 1606
rect 1215 1603 1216 1604
rect 1210 1602 1216 1603
rect 1407 1603 1408 1604
rect 1412 1603 1413 1607
rect 1407 1602 1413 1603
rect 1615 1607 1621 1608
rect 1615 1603 1616 1607
rect 1620 1606 1621 1607
rect 1642 1607 1648 1608
rect 1642 1606 1643 1607
rect 1620 1604 1643 1606
rect 1620 1603 1621 1604
rect 1615 1602 1621 1603
rect 1642 1603 1643 1604
rect 1647 1603 1648 1607
rect 1642 1602 1648 1603
rect 1666 1607 1672 1608
rect 1666 1603 1667 1607
rect 1671 1606 1672 1607
rect 1831 1607 1837 1608
rect 1831 1606 1832 1607
rect 1671 1604 1832 1606
rect 1671 1603 1672 1604
rect 1666 1602 1672 1603
rect 1831 1603 1832 1604
rect 1836 1603 1837 1607
rect 1831 1602 1837 1603
rect 2046 1604 2052 1605
rect 3942 1604 3948 1605
rect 2046 1600 2047 1604
rect 2051 1600 2052 1604
rect 2046 1599 2052 1600
rect 2390 1603 2396 1604
rect 2390 1599 2391 1603
rect 2395 1599 2396 1603
rect 2390 1598 2396 1599
rect 2502 1603 2508 1604
rect 2502 1599 2503 1603
rect 2507 1599 2508 1603
rect 2502 1598 2508 1599
rect 2614 1603 2620 1604
rect 2614 1599 2615 1603
rect 2619 1599 2620 1603
rect 2614 1598 2620 1599
rect 2734 1603 2740 1604
rect 2734 1599 2735 1603
rect 2739 1599 2740 1603
rect 2734 1598 2740 1599
rect 2854 1603 2860 1604
rect 2854 1599 2855 1603
rect 2859 1599 2860 1603
rect 2854 1598 2860 1599
rect 2974 1603 2980 1604
rect 2974 1599 2975 1603
rect 2979 1599 2980 1603
rect 2974 1598 2980 1599
rect 3094 1603 3100 1604
rect 3094 1599 3095 1603
rect 3099 1599 3100 1603
rect 3094 1598 3100 1599
rect 3214 1603 3220 1604
rect 3214 1599 3215 1603
rect 3219 1599 3220 1603
rect 3214 1598 3220 1599
rect 3334 1603 3340 1604
rect 3334 1599 3335 1603
rect 3339 1599 3340 1603
rect 3334 1598 3340 1599
rect 3454 1603 3460 1604
rect 3454 1599 3455 1603
rect 3459 1599 3460 1603
rect 3942 1600 3943 1604
rect 3947 1600 3948 1604
rect 3942 1599 3948 1600
rect 3454 1598 3460 1599
rect 2466 1595 2472 1596
rect 199 1591 205 1592
rect 199 1587 200 1591
rect 204 1590 205 1591
rect 218 1591 224 1592
rect 218 1590 219 1591
rect 204 1588 219 1590
rect 204 1587 205 1588
rect 199 1586 205 1587
rect 218 1587 219 1588
rect 223 1587 224 1591
rect 218 1586 224 1587
rect 319 1591 325 1592
rect 319 1587 320 1591
rect 324 1590 325 1591
rect 338 1591 344 1592
rect 338 1590 339 1591
rect 324 1588 339 1590
rect 324 1587 325 1588
rect 319 1586 325 1587
rect 338 1587 339 1588
rect 343 1587 344 1591
rect 338 1586 344 1587
rect 487 1591 493 1592
rect 487 1587 488 1591
rect 492 1590 493 1591
rect 574 1591 580 1592
rect 574 1590 575 1591
rect 492 1588 575 1590
rect 492 1587 493 1588
rect 487 1586 493 1587
rect 574 1587 575 1588
rect 579 1587 580 1591
rect 574 1586 580 1587
rect 679 1591 685 1592
rect 679 1587 680 1591
rect 684 1590 685 1591
rect 703 1591 709 1592
rect 703 1590 704 1591
rect 684 1588 704 1590
rect 684 1587 685 1588
rect 679 1586 685 1587
rect 703 1587 704 1588
rect 708 1587 709 1591
rect 703 1586 709 1587
rect 850 1591 856 1592
rect 850 1587 851 1591
rect 855 1590 856 1591
rect 895 1591 901 1592
rect 895 1590 896 1591
rect 855 1588 896 1590
rect 855 1587 856 1588
rect 850 1586 856 1587
rect 895 1587 896 1588
rect 900 1587 901 1591
rect 895 1586 901 1587
rect 1127 1591 1133 1592
rect 1127 1587 1128 1591
rect 1132 1590 1133 1591
rect 1146 1591 1152 1592
rect 1146 1590 1147 1591
rect 1132 1588 1147 1590
rect 1132 1587 1133 1588
rect 1127 1586 1133 1587
rect 1146 1587 1147 1588
rect 1151 1587 1152 1591
rect 1146 1586 1152 1587
rect 1375 1591 1381 1592
rect 1375 1587 1376 1591
rect 1380 1590 1381 1591
rect 1410 1591 1416 1592
rect 1410 1590 1411 1591
rect 1380 1588 1411 1590
rect 1380 1587 1381 1588
rect 1375 1586 1381 1587
rect 1410 1587 1411 1588
rect 1415 1587 1416 1591
rect 1410 1586 1416 1587
rect 1631 1591 1637 1592
rect 1631 1587 1632 1591
rect 1636 1590 1637 1591
rect 1650 1591 1656 1592
rect 1650 1590 1651 1591
rect 1636 1588 1651 1590
rect 1636 1587 1637 1588
rect 1631 1586 1637 1587
rect 1650 1587 1651 1588
rect 1655 1587 1656 1591
rect 1650 1586 1656 1587
rect 1810 1591 1816 1592
rect 1810 1587 1811 1591
rect 1815 1590 1816 1591
rect 1895 1591 1901 1592
rect 1895 1590 1896 1591
rect 1815 1588 1896 1590
rect 1815 1587 1816 1588
rect 1810 1586 1816 1587
rect 1895 1587 1896 1588
rect 1900 1587 1901 1591
rect 2466 1591 2467 1595
rect 2471 1591 2472 1595
rect 2466 1590 2472 1591
rect 2578 1595 2584 1596
rect 2578 1591 2579 1595
rect 2583 1591 2584 1595
rect 2726 1595 2732 1596
rect 2726 1594 2727 1595
rect 2693 1592 2727 1594
rect 2578 1590 2584 1591
rect 2726 1591 2727 1592
rect 2731 1591 2732 1595
rect 2726 1590 2732 1591
rect 2810 1595 2816 1596
rect 2810 1591 2811 1595
rect 2815 1591 2816 1595
rect 2810 1590 2816 1591
rect 2818 1595 2824 1596
rect 2818 1591 2819 1595
rect 2823 1594 2824 1595
rect 3050 1595 3056 1596
rect 2823 1592 2897 1594
rect 2823 1591 2824 1592
rect 2818 1590 2824 1591
rect 3050 1591 3051 1595
rect 3055 1591 3056 1595
rect 3050 1590 3056 1591
rect 3170 1595 3176 1596
rect 3170 1591 3171 1595
rect 3175 1591 3176 1595
rect 3170 1590 3176 1591
rect 3290 1595 3296 1596
rect 3290 1591 3291 1595
rect 3295 1591 3296 1595
rect 3290 1590 3296 1591
rect 3410 1595 3416 1596
rect 3410 1591 3411 1595
rect 3415 1591 3416 1595
rect 3410 1590 3416 1591
rect 3418 1595 3424 1596
rect 3418 1591 3419 1595
rect 3423 1594 3424 1595
rect 3423 1592 3497 1594
rect 3423 1591 3424 1592
rect 3418 1590 3424 1591
rect 1895 1586 1901 1587
rect 2046 1587 2052 1588
rect 2046 1583 2047 1587
rect 2051 1583 2052 1587
rect 3942 1587 3948 1588
rect 2046 1582 2052 1583
rect 2390 1584 2396 1585
rect 2390 1580 2391 1584
rect 2395 1580 2396 1584
rect 2390 1579 2396 1580
rect 2502 1584 2508 1585
rect 2502 1580 2503 1584
rect 2507 1580 2508 1584
rect 2502 1579 2508 1580
rect 2614 1584 2620 1585
rect 2614 1580 2615 1584
rect 2619 1580 2620 1584
rect 2614 1579 2620 1580
rect 2734 1584 2740 1585
rect 2734 1580 2735 1584
rect 2739 1580 2740 1584
rect 2734 1579 2740 1580
rect 2854 1584 2860 1585
rect 2854 1580 2855 1584
rect 2859 1580 2860 1584
rect 2854 1579 2860 1580
rect 2974 1584 2980 1585
rect 2974 1580 2975 1584
rect 2979 1580 2980 1584
rect 2974 1579 2980 1580
rect 3094 1584 3100 1585
rect 3094 1580 3095 1584
rect 3099 1580 3100 1584
rect 3094 1579 3100 1580
rect 3214 1584 3220 1585
rect 3214 1580 3215 1584
rect 3219 1580 3220 1584
rect 3214 1579 3220 1580
rect 3334 1584 3340 1585
rect 3334 1580 3335 1584
rect 3339 1580 3340 1584
rect 3334 1579 3340 1580
rect 3454 1584 3460 1585
rect 3454 1580 3455 1584
rect 3459 1580 3460 1584
rect 3942 1583 3943 1587
rect 3947 1583 3948 1587
rect 3942 1582 3948 1583
rect 3454 1579 3460 1580
rect 110 1572 116 1573
rect 2006 1572 2012 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 110 1567 116 1568
rect 134 1571 140 1572
rect 134 1567 135 1571
rect 139 1567 140 1571
rect 134 1566 140 1567
rect 254 1571 260 1572
rect 254 1567 255 1571
rect 259 1567 260 1571
rect 254 1566 260 1567
rect 422 1571 428 1572
rect 422 1567 423 1571
rect 427 1567 428 1571
rect 422 1566 428 1567
rect 614 1571 620 1572
rect 614 1567 615 1571
rect 619 1567 620 1571
rect 614 1566 620 1567
rect 830 1571 836 1572
rect 830 1567 831 1571
rect 835 1567 836 1571
rect 830 1566 836 1567
rect 1062 1571 1068 1572
rect 1062 1567 1063 1571
rect 1067 1567 1068 1571
rect 1062 1566 1068 1567
rect 1310 1571 1316 1572
rect 1310 1567 1311 1571
rect 1315 1567 1316 1571
rect 1310 1566 1316 1567
rect 1566 1571 1572 1572
rect 1566 1567 1567 1571
rect 1571 1567 1572 1571
rect 1566 1566 1572 1567
rect 1830 1571 1836 1572
rect 1830 1567 1831 1571
rect 1835 1567 1836 1571
rect 2006 1568 2007 1572
rect 2011 1568 2012 1572
rect 2006 1567 2012 1568
rect 1830 1566 1836 1567
rect 210 1563 216 1564
rect 210 1559 211 1563
rect 215 1559 216 1563
rect 210 1558 216 1559
rect 218 1563 224 1564
rect 218 1559 219 1563
rect 223 1562 224 1563
rect 338 1563 344 1564
rect 223 1560 297 1562
rect 223 1559 224 1560
rect 218 1558 224 1559
rect 338 1559 339 1563
rect 343 1562 344 1563
rect 574 1563 580 1564
rect 343 1560 465 1562
rect 343 1559 344 1560
rect 338 1558 344 1559
rect 574 1559 575 1563
rect 579 1562 580 1563
rect 703 1563 709 1564
rect 579 1560 657 1562
rect 579 1559 580 1560
rect 574 1558 580 1559
rect 703 1559 704 1563
rect 708 1562 709 1563
rect 1034 1563 1040 1564
rect 708 1560 873 1562
rect 708 1559 709 1560
rect 703 1558 709 1559
rect 1034 1559 1035 1563
rect 1039 1562 1040 1563
rect 1146 1563 1152 1564
rect 1039 1560 1105 1562
rect 1039 1559 1040 1560
rect 1034 1558 1040 1559
rect 1146 1559 1147 1563
rect 1151 1562 1152 1563
rect 1642 1563 1648 1564
rect 1151 1560 1353 1562
rect 1151 1559 1152 1560
rect 1146 1558 1152 1559
rect 1642 1559 1643 1563
rect 1647 1559 1648 1563
rect 1642 1558 1648 1559
rect 1650 1563 1656 1564
rect 1650 1559 1651 1563
rect 1655 1562 1656 1563
rect 1655 1560 1873 1562
rect 1655 1559 1656 1560
rect 1650 1558 1656 1559
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 2006 1555 2012 1556
rect 110 1550 116 1551
rect 134 1552 140 1553
rect 134 1548 135 1552
rect 139 1548 140 1552
rect 134 1547 140 1548
rect 254 1552 260 1553
rect 254 1548 255 1552
rect 259 1548 260 1552
rect 254 1547 260 1548
rect 422 1552 428 1553
rect 422 1548 423 1552
rect 427 1548 428 1552
rect 422 1547 428 1548
rect 614 1552 620 1553
rect 614 1548 615 1552
rect 619 1548 620 1552
rect 614 1547 620 1548
rect 830 1552 836 1553
rect 830 1548 831 1552
rect 835 1548 836 1552
rect 830 1547 836 1548
rect 1062 1552 1068 1553
rect 1062 1548 1063 1552
rect 1067 1548 1068 1552
rect 1062 1547 1068 1548
rect 1310 1552 1316 1553
rect 1310 1548 1311 1552
rect 1315 1548 1316 1552
rect 1310 1547 1316 1548
rect 1566 1552 1572 1553
rect 1566 1548 1567 1552
rect 1571 1548 1572 1552
rect 1566 1547 1572 1548
rect 1830 1552 1836 1553
rect 1830 1548 1831 1552
rect 1835 1548 1836 1552
rect 2006 1551 2007 1555
rect 2011 1551 2012 1555
rect 2006 1550 2012 1551
rect 1830 1547 1836 1548
rect 2542 1524 2548 1525
rect 2046 1521 2052 1522
rect 2046 1517 2047 1521
rect 2051 1517 2052 1521
rect 2542 1520 2543 1524
rect 2547 1520 2548 1524
rect 2542 1519 2548 1520
rect 2670 1524 2676 1525
rect 2670 1520 2671 1524
rect 2675 1520 2676 1524
rect 2670 1519 2676 1520
rect 2798 1524 2804 1525
rect 2798 1520 2799 1524
rect 2803 1520 2804 1524
rect 2798 1519 2804 1520
rect 2934 1524 2940 1525
rect 2934 1520 2935 1524
rect 2939 1520 2940 1524
rect 2934 1519 2940 1520
rect 3070 1524 3076 1525
rect 3070 1520 3071 1524
rect 3075 1520 3076 1524
rect 3070 1519 3076 1520
rect 3206 1524 3212 1525
rect 3206 1520 3207 1524
rect 3211 1520 3212 1524
rect 3206 1519 3212 1520
rect 3334 1524 3340 1525
rect 3334 1520 3335 1524
rect 3339 1520 3340 1524
rect 3334 1519 3340 1520
rect 3462 1524 3468 1525
rect 3462 1520 3463 1524
rect 3467 1520 3468 1524
rect 3462 1519 3468 1520
rect 3590 1524 3596 1525
rect 3590 1520 3591 1524
rect 3595 1520 3596 1524
rect 3590 1519 3596 1520
rect 3726 1524 3732 1525
rect 3726 1520 3727 1524
rect 3731 1520 3732 1524
rect 3726 1519 3732 1520
rect 3838 1524 3844 1525
rect 3838 1520 3839 1524
rect 3843 1520 3844 1524
rect 3838 1519 3844 1520
rect 3942 1521 3948 1522
rect 2046 1516 2052 1517
rect 3942 1517 3943 1521
rect 3947 1517 3948 1521
rect 3942 1516 3948 1517
rect 2618 1515 2624 1516
rect 2618 1511 2619 1515
rect 2623 1511 2624 1515
rect 2618 1510 2624 1511
rect 2746 1515 2752 1516
rect 2746 1511 2747 1515
rect 2751 1511 2752 1515
rect 2746 1510 2752 1511
rect 2874 1515 2880 1516
rect 2874 1511 2875 1515
rect 2879 1511 2880 1515
rect 2874 1510 2880 1511
rect 3010 1515 3016 1516
rect 3010 1511 3011 1515
rect 3015 1511 3016 1515
rect 3010 1510 3016 1511
rect 3146 1515 3152 1516
rect 3146 1511 3147 1515
rect 3151 1511 3152 1515
rect 3146 1510 3152 1511
rect 3282 1515 3288 1516
rect 3282 1511 3283 1515
rect 3287 1511 3288 1515
rect 3282 1510 3288 1511
rect 3410 1515 3416 1516
rect 3410 1511 3411 1515
rect 3415 1511 3416 1515
rect 3410 1510 3416 1511
rect 3538 1515 3544 1516
rect 3538 1511 3539 1515
rect 3543 1511 3544 1515
rect 3719 1515 3725 1516
rect 3719 1514 3720 1515
rect 3669 1512 3720 1514
rect 3538 1510 3544 1511
rect 3719 1511 3720 1512
rect 3724 1511 3725 1515
rect 3719 1510 3725 1511
rect 3794 1515 3800 1516
rect 3794 1511 3795 1515
rect 3799 1511 3800 1515
rect 3794 1510 3800 1511
rect 3906 1515 3912 1516
rect 3906 1511 3907 1515
rect 3911 1511 3912 1515
rect 3906 1510 3912 1511
rect 2542 1505 2548 1506
rect 2046 1504 2052 1505
rect 2046 1500 2047 1504
rect 2051 1500 2052 1504
rect 2542 1501 2543 1505
rect 2547 1501 2548 1505
rect 2542 1500 2548 1501
rect 2670 1505 2676 1506
rect 2670 1501 2671 1505
rect 2675 1501 2676 1505
rect 2670 1500 2676 1501
rect 2798 1505 2804 1506
rect 2798 1501 2799 1505
rect 2803 1501 2804 1505
rect 2798 1500 2804 1501
rect 2934 1505 2940 1506
rect 2934 1501 2935 1505
rect 2939 1501 2940 1505
rect 2934 1500 2940 1501
rect 3070 1505 3076 1506
rect 3070 1501 3071 1505
rect 3075 1501 3076 1505
rect 3070 1500 3076 1501
rect 3206 1505 3212 1506
rect 3206 1501 3207 1505
rect 3211 1501 3212 1505
rect 3206 1500 3212 1501
rect 3334 1505 3340 1506
rect 3334 1501 3335 1505
rect 3339 1501 3340 1505
rect 3334 1500 3340 1501
rect 3462 1505 3468 1506
rect 3462 1501 3463 1505
rect 3467 1501 3468 1505
rect 3462 1500 3468 1501
rect 3590 1505 3596 1506
rect 3590 1501 3591 1505
rect 3595 1501 3596 1505
rect 3590 1500 3596 1501
rect 3726 1505 3732 1506
rect 3726 1501 3727 1505
rect 3731 1501 3732 1505
rect 3726 1500 3732 1501
rect 3838 1505 3844 1506
rect 3838 1501 3839 1505
rect 3843 1501 3844 1505
rect 3838 1500 3844 1501
rect 3942 1504 3948 1505
rect 3942 1500 3943 1504
rect 3947 1500 3948 1504
rect 2046 1499 2052 1500
rect 3942 1499 3948 1500
rect 2818 1491 2824 1492
rect 2818 1490 2819 1491
rect 238 1488 244 1489
rect 110 1485 116 1486
rect 110 1481 111 1485
rect 115 1481 116 1485
rect 238 1484 239 1488
rect 243 1484 244 1488
rect 238 1483 244 1484
rect 406 1488 412 1489
rect 406 1484 407 1488
rect 411 1484 412 1488
rect 406 1483 412 1484
rect 582 1488 588 1489
rect 582 1484 583 1488
rect 587 1484 588 1488
rect 582 1483 588 1484
rect 774 1488 780 1489
rect 774 1484 775 1488
rect 779 1484 780 1488
rect 774 1483 780 1484
rect 966 1488 972 1489
rect 966 1484 967 1488
rect 971 1484 972 1488
rect 966 1483 972 1484
rect 1158 1488 1164 1489
rect 1158 1484 1159 1488
rect 1163 1484 1164 1488
rect 1158 1483 1164 1484
rect 1350 1488 1356 1489
rect 1350 1484 1351 1488
rect 1355 1484 1356 1488
rect 1350 1483 1356 1484
rect 1542 1488 1548 1489
rect 1542 1484 1543 1488
rect 1547 1484 1548 1488
rect 1542 1483 1548 1484
rect 1734 1488 1740 1489
rect 1734 1484 1735 1488
rect 1739 1484 1740 1488
rect 1734 1483 1740 1484
rect 1902 1488 1908 1489
rect 1902 1484 1903 1488
rect 1907 1484 1908 1488
rect 2612 1488 2819 1490
rect 1902 1483 1908 1484
rect 2006 1485 2012 1486
rect 110 1480 116 1481
rect 2006 1481 2007 1485
rect 2011 1481 2012 1485
rect 2612 1484 2614 1488
rect 2818 1487 2819 1488
rect 2823 1487 2824 1491
rect 3418 1491 3424 1492
rect 3418 1490 3419 1491
rect 2818 1486 2824 1487
rect 3276 1488 3419 1490
rect 3276 1484 3278 1488
rect 3418 1487 3419 1488
rect 3423 1487 3424 1491
rect 3418 1486 3424 1487
rect 2006 1480 2012 1481
rect 2607 1483 2614 1484
rect 391 1479 397 1480
rect 391 1478 392 1479
rect 317 1476 392 1478
rect 391 1475 392 1476
rect 396 1475 397 1479
rect 391 1474 397 1475
rect 482 1479 488 1480
rect 482 1475 483 1479
rect 487 1475 488 1479
rect 482 1474 488 1475
rect 658 1479 664 1480
rect 658 1475 659 1479
rect 663 1475 664 1479
rect 658 1474 664 1475
rect 850 1479 856 1480
rect 850 1475 851 1479
rect 855 1475 856 1479
rect 850 1474 856 1475
rect 1042 1479 1048 1480
rect 1042 1475 1043 1479
rect 1047 1475 1048 1479
rect 1042 1474 1048 1475
rect 1234 1479 1240 1480
rect 1234 1475 1235 1479
rect 1239 1475 1240 1479
rect 1442 1479 1448 1480
rect 1442 1478 1443 1479
rect 1429 1476 1443 1478
rect 1234 1474 1240 1475
rect 1442 1475 1443 1476
rect 1447 1475 1448 1479
rect 1442 1474 1448 1475
rect 1618 1479 1624 1480
rect 1618 1475 1619 1479
rect 1623 1475 1624 1479
rect 1618 1474 1624 1475
rect 1810 1479 1816 1480
rect 1810 1475 1811 1479
rect 1815 1475 1816 1479
rect 1810 1474 1816 1475
rect 1818 1479 1824 1480
rect 1818 1475 1819 1479
rect 1823 1478 1824 1479
rect 2607 1479 2608 1483
rect 2612 1480 2614 1483
rect 2618 1483 2624 1484
rect 2612 1479 2613 1480
rect 2607 1478 2613 1479
rect 2618 1479 2619 1483
rect 2623 1482 2624 1483
rect 2735 1483 2741 1484
rect 2735 1482 2736 1483
rect 2623 1480 2736 1482
rect 2623 1479 2624 1480
rect 2618 1478 2624 1479
rect 2735 1479 2736 1480
rect 2740 1479 2741 1483
rect 2735 1478 2741 1479
rect 2746 1483 2752 1484
rect 2746 1479 2747 1483
rect 2751 1482 2752 1483
rect 2863 1483 2869 1484
rect 2863 1482 2864 1483
rect 2751 1480 2864 1482
rect 2751 1479 2752 1480
rect 2746 1478 2752 1479
rect 2863 1479 2864 1480
rect 2868 1479 2869 1483
rect 2863 1478 2869 1479
rect 2874 1483 2880 1484
rect 2874 1479 2875 1483
rect 2879 1482 2880 1483
rect 2999 1483 3005 1484
rect 2999 1482 3000 1483
rect 2879 1480 3000 1482
rect 2879 1479 2880 1480
rect 2874 1478 2880 1479
rect 2999 1479 3000 1480
rect 3004 1479 3005 1483
rect 2999 1478 3005 1479
rect 3010 1483 3016 1484
rect 3010 1479 3011 1483
rect 3015 1482 3016 1483
rect 3135 1483 3141 1484
rect 3135 1482 3136 1483
rect 3015 1480 3136 1482
rect 3015 1479 3016 1480
rect 3010 1478 3016 1479
rect 3135 1479 3136 1480
rect 3140 1479 3141 1483
rect 3135 1478 3141 1479
rect 3271 1483 3278 1484
rect 3271 1479 3272 1483
rect 3276 1480 3278 1483
rect 3282 1483 3288 1484
rect 3276 1479 3277 1480
rect 3271 1478 3277 1479
rect 3282 1479 3283 1483
rect 3287 1482 3288 1483
rect 3399 1483 3405 1484
rect 3399 1482 3400 1483
rect 3287 1480 3400 1482
rect 3287 1479 3288 1480
rect 3282 1478 3288 1479
rect 3399 1479 3400 1480
rect 3404 1479 3405 1483
rect 3399 1478 3405 1479
rect 3410 1483 3416 1484
rect 3410 1479 3411 1483
rect 3415 1482 3416 1483
rect 3527 1483 3533 1484
rect 3527 1482 3528 1483
rect 3415 1480 3528 1482
rect 3415 1479 3416 1480
rect 3410 1478 3416 1479
rect 3527 1479 3528 1480
rect 3532 1479 3533 1483
rect 3527 1478 3533 1479
rect 3538 1483 3544 1484
rect 3538 1479 3539 1483
rect 3543 1482 3544 1483
rect 3655 1483 3661 1484
rect 3655 1482 3656 1483
rect 3543 1480 3656 1482
rect 3543 1479 3544 1480
rect 3538 1478 3544 1479
rect 3655 1479 3656 1480
rect 3660 1479 3661 1483
rect 3655 1478 3661 1479
rect 3790 1483 3797 1484
rect 3790 1479 3791 1483
rect 3796 1479 3797 1483
rect 3790 1478 3797 1479
rect 3903 1483 3909 1484
rect 3903 1479 3904 1483
rect 3908 1482 3909 1483
rect 3914 1483 3920 1484
rect 3914 1482 3915 1483
rect 3908 1480 3915 1482
rect 3908 1479 3909 1480
rect 3903 1478 3909 1479
rect 3914 1479 3915 1480
rect 3919 1479 3920 1483
rect 3914 1478 3920 1479
rect 1823 1476 1945 1478
rect 1823 1475 1824 1476
rect 1818 1474 1824 1475
rect 238 1469 244 1470
rect 110 1468 116 1469
rect 110 1464 111 1468
rect 115 1464 116 1468
rect 238 1465 239 1469
rect 243 1465 244 1469
rect 238 1464 244 1465
rect 406 1469 412 1470
rect 406 1465 407 1469
rect 411 1465 412 1469
rect 406 1464 412 1465
rect 582 1469 588 1470
rect 582 1465 583 1469
rect 587 1465 588 1469
rect 582 1464 588 1465
rect 774 1469 780 1470
rect 774 1465 775 1469
rect 779 1465 780 1469
rect 774 1464 780 1465
rect 966 1469 972 1470
rect 966 1465 967 1469
rect 971 1465 972 1469
rect 966 1464 972 1465
rect 1158 1469 1164 1470
rect 1158 1465 1159 1469
rect 1163 1465 1164 1469
rect 1158 1464 1164 1465
rect 1350 1469 1356 1470
rect 1350 1465 1351 1469
rect 1355 1465 1356 1469
rect 1350 1464 1356 1465
rect 1542 1469 1548 1470
rect 1542 1465 1543 1469
rect 1547 1465 1548 1469
rect 1542 1464 1548 1465
rect 1734 1469 1740 1470
rect 1734 1465 1735 1469
rect 1739 1465 1740 1469
rect 1734 1464 1740 1465
rect 1902 1469 1908 1470
rect 1902 1465 1903 1469
rect 1907 1465 1908 1469
rect 1902 1464 1908 1465
rect 2006 1468 2012 1469
rect 2006 1464 2007 1468
rect 2011 1464 2012 1468
rect 110 1463 116 1464
rect 2006 1463 2012 1464
rect 2583 1459 2589 1460
rect 391 1455 397 1456
rect 391 1451 392 1455
rect 396 1454 397 1455
rect 1818 1455 1824 1456
rect 1818 1454 1819 1455
rect 396 1452 418 1454
rect 396 1451 397 1452
rect 391 1450 397 1451
rect 303 1447 309 1448
rect 303 1443 304 1447
rect 308 1446 309 1447
rect 407 1447 413 1448
rect 407 1446 408 1447
rect 308 1444 408 1446
rect 308 1443 309 1444
rect 303 1442 309 1443
rect 407 1443 408 1444
rect 412 1443 413 1447
rect 416 1446 418 1452
rect 1612 1452 1819 1454
rect 1612 1448 1614 1452
rect 1818 1451 1819 1452
rect 1823 1451 1824 1455
rect 2583 1455 2584 1459
rect 2588 1458 2589 1459
rect 2594 1459 2600 1460
rect 2588 1455 2590 1458
rect 2583 1454 2590 1455
rect 2594 1455 2595 1459
rect 2599 1458 2600 1459
rect 2695 1459 2701 1460
rect 2695 1458 2696 1459
rect 2599 1456 2696 1458
rect 2599 1455 2600 1456
rect 2594 1454 2600 1455
rect 2695 1455 2696 1456
rect 2700 1455 2701 1459
rect 2695 1454 2701 1455
rect 2823 1459 2829 1460
rect 2823 1455 2824 1459
rect 2828 1458 2829 1459
rect 2886 1459 2892 1460
rect 2886 1458 2887 1459
rect 2828 1456 2887 1458
rect 2828 1455 2829 1456
rect 2823 1454 2829 1455
rect 2886 1455 2887 1456
rect 2891 1455 2892 1459
rect 2886 1454 2892 1455
rect 2959 1459 2965 1460
rect 2959 1455 2960 1459
rect 2964 1458 2965 1459
rect 2978 1459 2984 1460
rect 2978 1458 2979 1459
rect 2964 1456 2979 1458
rect 2964 1455 2965 1456
rect 2959 1454 2965 1455
rect 2978 1455 2979 1456
rect 2983 1455 2984 1459
rect 2978 1454 2984 1455
rect 3095 1459 3101 1460
rect 3095 1455 3096 1459
rect 3100 1458 3101 1459
rect 3119 1459 3125 1460
rect 3119 1458 3120 1459
rect 3100 1456 3120 1458
rect 3100 1455 3101 1456
rect 3095 1454 3101 1455
rect 3119 1455 3120 1456
rect 3124 1455 3125 1459
rect 3119 1454 3125 1455
rect 3146 1459 3152 1460
rect 3146 1455 3147 1459
rect 3151 1458 3152 1459
rect 3239 1459 3245 1460
rect 3239 1458 3240 1459
rect 3151 1456 3240 1458
rect 3151 1455 3152 1456
rect 3146 1454 3152 1455
rect 3239 1455 3240 1456
rect 3244 1455 3245 1459
rect 3239 1454 3245 1455
rect 3375 1459 3381 1460
rect 3375 1455 3376 1459
rect 3380 1458 3381 1459
rect 3386 1459 3392 1460
rect 3380 1455 3382 1458
rect 3375 1454 3382 1455
rect 3386 1455 3387 1459
rect 3391 1458 3392 1459
rect 3511 1459 3517 1460
rect 3511 1458 3512 1459
rect 3391 1456 3512 1458
rect 3391 1455 3392 1456
rect 3386 1454 3392 1455
rect 3511 1455 3512 1456
rect 3516 1455 3517 1459
rect 3511 1454 3517 1455
rect 3647 1459 3653 1460
rect 3647 1455 3648 1459
rect 3652 1458 3653 1459
rect 3666 1459 3672 1460
rect 3666 1458 3667 1459
rect 3652 1456 3667 1458
rect 3652 1455 3653 1456
rect 3647 1454 3653 1455
rect 3666 1455 3667 1456
rect 3671 1455 3672 1459
rect 3666 1454 3672 1455
rect 3719 1459 3725 1460
rect 3719 1455 3720 1459
rect 3724 1458 3725 1459
rect 3783 1459 3789 1460
rect 3783 1458 3784 1459
rect 3724 1456 3784 1458
rect 3724 1455 3725 1456
rect 3719 1454 3725 1455
rect 3783 1455 3784 1456
rect 3788 1455 3789 1459
rect 3783 1454 3789 1455
rect 3903 1459 3912 1460
rect 3903 1455 3904 1459
rect 3911 1455 3912 1459
rect 3903 1454 3912 1455
rect 1818 1450 1824 1451
rect 2588 1450 2590 1454
rect 2714 1451 2720 1452
rect 2714 1450 2715 1451
rect 2588 1448 2715 1450
rect 471 1447 477 1448
rect 471 1446 472 1447
rect 416 1444 472 1446
rect 407 1442 413 1443
rect 471 1443 472 1444
rect 476 1443 477 1447
rect 471 1442 477 1443
rect 482 1447 488 1448
rect 482 1443 483 1447
rect 487 1446 488 1447
rect 647 1447 653 1448
rect 647 1446 648 1447
rect 487 1444 648 1446
rect 487 1443 488 1444
rect 482 1442 488 1443
rect 647 1443 648 1444
rect 652 1443 653 1447
rect 647 1442 653 1443
rect 658 1447 664 1448
rect 658 1443 659 1447
rect 663 1446 664 1447
rect 839 1447 845 1448
rect 839 1446 840 1447
rect 663 1444 840 1446
rect 663 1443 664 1444
rect 658 1442 664 1443
rect 839 1443 840 1444
rect 844 1443 845 1447
rect 839 1442 845 1443
rect 1031 1447 1040 1448
rect 1031 1443 1032 1447
rect 1039 1443 1040 1447
rect 1031 1442 1040 1443
rect 1042 1447 1048 1448
rect 1042 1443 1043 1447
rect 1047 1446 1048 1447
rect 1223 1447 1229 1448
rect 1223 1446 1224 1447
rect 1047 1444 1224 1446
rect 1047 1443 1048 1444
rect 1042 1442 1048 1443
rect 1223 1443 1224 1444
rect 1228 1443 1229 1447
rect 1223 1442 1229 1443
rect 1234 1447 1240 1448
rect 1234 1443 1235 1447
rect 1239 1446 1240 1447
rect 1415 1447 1421 1448
rect 1415 1446 1416 1447
rect 1239 1444 1416 1446
rect 1239 1443 1240 1444
rect 1234 1442 1240 1443
rect 1415 1443 1416 1444
rect 1420 1443 1421 1447
rect 1415 1442 1421 1443
rect 1607 1447 1614 1448
rect 1607 1443 1608 1447
rect 1612 1444 1614 1447
rect 1618 1447 1624 1448
rect 1612 1443 1613 1444
rect 1607 1442 1613 1443
rect 1618 1443 1619 1447
rect 1623 1446 1624 1447
rect 1799 1447 1805 1448
rect 1799 1446 1800 1447
rect 1623 1444 1800 1446
rect 1623 1443 1624 1444
rect 1618 1442 1624 1443
rect 1799 1443 1800 1444
rect 1804 1443 1805 1447
rect 1799 1442 1805 1443
rect 1946 1447 1952 1448
rect 1946 1443 1947 1447
rect 1951 1446 1952 1447
rect 1967 1447 1973 1448
rect 1967 1446 1968 1447
rect 1951 1444 1968 1446
rect 1951 1443 1952 1444
rect 1946 1442 1952 1443
rect 1967 1443 1968 1444
rect 1972 1443 1973 1447
rect 2714 1447 2715 1448
rect 2719 1447 2720 1451
rect 3380 1450 3382 1454
rect 3530 1451 3536 1452
rect 3530 1450 3531 1451
rect 3380 1448 3531 1450
rect 2714 1446 2720 1447
rect 3530 1447 3531 1448
rect 3535 1447 3536 1451
rect 3530 1446 3536 1447
rect 1967 1442 1973 1443
rect 2046 1440 2052 1441
rect 3942 1440 3948 1441
rect 2046 1436 2047 1440
rect 2051 1436 2052 1440
rect 2046 1435 2052 1436
rect 2518 1439 2524 1440
rect 2518 1435 2519 1439
rect 2523 1435 2524 1439
rect 2518 1434 2524 1435
rect 2630 1439 2636 1440
rect 2630 1435 2631 1439
rect 2635 1435 2636 1439
rect 2630 1434 2636 1435
rect 2758 1439 2764 1440
rect 2758 1435 2759 1439
rect 2763 1435 2764 1439
rect 2758 1434 2764 1435
rect 2894 1439 2900 1440
rect 2894 1435 2895 1439
rect 2899 1435 2900 1439
rect 2894 1434 2900 1435
rect 3030 1439 3036 1440
rect 3030 1435 3031 1439
rect 3035 1435 3036 1439
rect 3030 1434 3036 1435
rect 3174 1439 3180 1440
rect 3174 1435 3175 1439
rect 3179 1435 3180 1439
rect 3174 1434 3180 1435
rect 3310 1439 3316 1440
rect 3310 1435 3311 1439
rect 3315 1435 3316 1439
rect 3310 1434 3316 1435
rect 3446 1439 3452 1440
rect 3446 1435 3447 1439
rect 3451 1435 3452 1439
rect 3446 1434 3452 1435
rect 3582 1439 3588 1440
rect 3582 1435 3583 1439
rect 3587 1435 3588 1439
rect 3582 1434 3588 1435
rect 3718 1439 3724 1440
rect 3718 1435 3719 1439
rect 3723 1435 3724 1439
rect 3718 1434 3724 1435
rect 3838 1439 3844 1440
rect 3838 1435 3839 1439
rect 3843 1435 3844 1439
rect 3942 1436 3943 1440
rect 3947 1436 3948 1440
rect 3942 1435 3948 1436
rect 3838 1434 3844 1435
rect 2594 1431 2600 1432
rect 527 1427 533 1428
rect 527 1423 528 1427
rect 532 1426 533 1427
rect 551 1427 557 1428
rect 551 1426 552 1427
rect 532 1424 552 1426
rect 532 1423 533 1424
rect 527 1422 533 1423
rect 551 1423 552 1424
rect 556 1423 557 1427
rect 551 1422 557 1423
rect 647 1427 653 1428
rect 647 1423 648 1427
rect 652 1426 653 1427
rect 670 1427 676 1428
rect 670 1426 671 1427
rect 652 1424 671 1426
rect 652 1423 653 1424
rect 647 1422 653 1423
rect 670 1423 671 1424
rect 675 1423 676 1427
rect 670 1422 676 1423
rect 775 1427 781 1428
rect 775 1423 776 1427
rect 780 1426 781 1427
rect 799 1427 805 1428
rect 799 1426 800 1427
rect 780 1424 800 1426
rect 780 1423 781 1424
rect 775 1422 781 1423
rect 799 1423 800 1424
rect 804 1423 805 1427
rect 799 1422 805 1423
rect 919 1427 925 1428
rect 919 1423 920 1427
rect 924 1426 925 1427
rect 938 1427 944 1428
rect 938 1426 939 1427
rect 924 1424 939 1426
rect 924 1423 925 1424
rect 919 1422 925 1423
rect 938 1423 939 1424
rect 943 1423 944 1427
rect 938 1422 944 1423
rect 1071 1427 1077 1428
rect 1071 1423 1072 1427
rect 1076 1426 1077 1427
rect 1114 1427 1120 1428
rect 1114 1426 1115 1427
rect 1076 1424 1115 1426
rect 1076 1423 1077 1424
rect 1071 1422 1077 1423
rect 1114 1423 1115 1424
rect 1119 1423 1120 1427
rect 1114 1422 1120 1423
rect 1231 1427 1237 1428
rect 1231 1423 1232 1427
rect 1236 1426 1237 1427
rect 1250 1427 1256 1428
rect 1250 1426 1251 1427
rect 1236 1424 1251 1426
rect 1236 1423 1237 1424
rect 1231 1422 1237 1423
rect 1250 1423 1251 1424
rect 1255 1423 1256 1427
rect 1250 1422 1256 1423
rect 1399 1427 1405 1428
rect 1399 1423 1400 1427
rect 1404 1426 1405 1427
rect 1423 1427 1429 1428
rect 1423 1426 1424 1427
rect 1404 1424 1424 1426
rect 1404 1423 1405 1424
rect 1399 1422 1405 1423
rect 1423 1423 1424 1424
rect 1428 1423 1429 1427
rect 1423 1422 1429 1423
rect 1442 1427 1448 1428
rect 1442 1423 1443 1427
rect 1447 1426 1448 1427
rect 1575 1427 1581 1428
rect 1575 1426 1576 1427
rect 1447 1424 1576 1426
rect 1447 1423 1448 1424
rect 1442 1422 1448 1423
rect 1575 1423 1576 1424
rect 1580 1423 1581 1427
rect 1575 1422 1581 1423
rect 1751 1427 1757 1428
rect 1751 1423 1752 1427
rect 1756 1426 1757 1427
rect 1822 1427 1828 1428
rect 1822 1426 1823 1427
rect 1756 1424 1823 1426
rect 1756 1423 1757 1424
rect 1751 1422 1757 1423
rect 1822 1423 1823 1424
rect 1827 1423 1828 1427
rect 1822 1422 1828 1423
rect 1830 1427 1836 1428
rect 1830 1423 1831 1427
rect 1835 1426 1836 1427
rect 1935 1427 1941 1428
rect 1935 1426 1936 1427
rect 1835 1424 1936 1426
rect 1835 1423 1836 1424
rect 1830 1422 1836 1423
rect 1935 1423 1936 1424
rect 1940 1423 1941 1427
rect 2594 1427 2595 1431
rect 2599 1427 2600 1431
rect 2714 1431 2720 1432
rect 2594 1426 2600 1427
rect 2706 1427 2712 1428
rect 1935 1422 1941 1423
rect 2046 1423 2052 1424
rect 2046 1419 2047 1423
rect 2051 1419 2052 1423
rect 2706 1423 2707 1427
rect 2711 1423 2712 1427
rect 2714 1427 2715 1431
rect 2719 1430 2720 1431
rect 2886 1431 2892 1432
rect 2719 1428 2801 1430
rect 2719 1427 2720 1428
rect 2714 1426 2720 1427
rect 2886 1427 2887 1431
rect 2891 1430 2892 1431
rect 2978 1431 2984 1432
rect 2891 1428 2937 1430
rect 2891 1427 2892 1428
rect 2886 1426 2892 1427
rect 2978 1427 2979 1431
rect 2983 1430 2984 1431
rect 3119 1431 3125 1432
rect 2983 1428 3073 1430
rect 2983 1427 2984 1428
rect 2978 1426 2984 1427
rect 3119 1427 3120 1431
rect 3124 1430 3125 1431
rect 3386 1431 3392 1432
rect 3124 1428 3217 1430
rect 3124 1427 3125 1428
rect 3119 1426 3125 1427
rect 3386 1427 3387 1431
rect 3391 1427 3392 1431
rect 3386 1426 3392 1427
rect 3530 1431 3536 1432
rect 3530 1427 3531 1431
rect 3535 1430 3536 1431
rect 3666 1431 3672 1432
rect 3535 1428 3625 1430
rect 3535 1427 3536 1428
rect 3530 1426 3536 1427
rect 3666 1427 3667 1431
rect 3671 1430 3672 1431
rect 3671 1428 3761 1430
rect 3671 1427 3672 1428
rect 3666 1426 3672 1427
rect 2706 1422 2712 1423
rect 3524 1422 3526 1425
rect 3574 1423 3580 1424
rect 3574 1422 3575 1423
rect 2046 1418 2052 1419
rect 2518 1420 2524 1421
rect 2518 1416 2519 1420
rect 2523 1416 2524 1420
rect 2518 1415 2524 1416
rect 2630 1420 2636 1421
rect 2630 1416 2631 1420
rect 2635 1416 2636 1420
rect 2630 1415 2636 1416
rect 2758 1420 2764 1421
rect 2758 1416 2759 1420
rect 2763 1416 2764 1420
rect 2758 1415 2764 1416
rect 2894 1420 2900 1421
rect 2894 1416 2895 1420
rect 2899 1416 2900 1420
rect 2894 1415 2900 1416
rect 3030 1420 3036 1421
rect 3030 1416 3031 1420
rect 3035 1416 3036 1420
rect 3030 1415 3036 1416
rect 3174 1420 3180 1421
rect 3174 1416 3175 1420
rect 3179 1416 3180 1420
rect 3174 1415 3180 1416
rect 3310 1420 3316 1421
rect 3310 1416 3311 1420
rect 3315 1416 3316 1420
rect 3310 1415 3316 1416
rect 3446 1420 3452 1421
rect 3524 1420 3575 1422
rect 3446 1416 3447 1420
rect 3451 1416 3452 1420
rect 3574 1419 3575 1420
rect 3579 1419 3580 1423
rect 3906 1423 3912 1424
rect 3574 1418 3580 1419
rect 3582 1420 3588 1421
rect 3446 1415 3452 1416
rect 3582 1416 3583 1420
rect 3587 1416 3588 1420
rect 3582 1415 3588 1416
rect 3718 1420 3724 1421
rect 3718 1416 3719 1420
rect 3723 1416 3724 1420
rect 3718 1415 3724 1416
rect 3838 1420 3844 1421
rect 3838 1416 3839 1420
rect 3843 1416 3844 1420
rect 3906 1419 3907 1423
rect 3911 1422 3912 1423
rect 3916 1422 3918 1425
rect 3911 1420 3918 1422
rect 3942 1423 3948 1424
rect 3911 1419 3912 1420
rect 3906 1418 3912 1419
rect 3942 1419 3943 1423
rect 3947 1419 3948 1423
rect 3942 1418 3948 1419
rect 3838 1415 3844 1416
rect 110 1408 116 1409
rect 2006 1408 2012 1409
rect 110 1404 111 1408
rect 115 1404 116 1408
rect 110 1403 116 1404
rect 462 1407 468 1408
rect 462 1403 463 1407
rect 467 1403 468 1407
rect 462 1402 468 1403
rect 582 1407 588 1408
rect 582 1403 583 1407
rect 587 1403 588 1407
rect 582 1402 588 1403
rect 710 1407 716 1408
rect 710 1403 711 1407
rect 715 1403 716 1407
rect 710 1402 716 1403
rect 854 1407 860 1408
rect 854 1403 855 1407
rect 859 1403 860 1407
rect 854 1402 860 1403
rect 1006 1407 1012 1408
rect 1006 1403 1007 1407
rect 1011 1403 1012 1407
rect 1006 1402 1012 1403
rect 1166 1407 1172 1408
rect 1166 1403 1167 1407
rect 1171 1403 1172 1407
rect 1166 1402 1172 1403
rect 1334 1407 1340 1408
rect 1334 1403 1335 1407
rect 1339 1403 1340 1407
rect 1334 1402 1340 1403
rect 1510 1407 1516 1408
rect 1510 1403 1511 1407
rect 1515 1403 1516 1407
rect 1510 1402 1516 1403
rect 1686 1407 1692 1408
rect 1686 1403 1687 1407
rect 1691 1403 1692 1407
rect 1686 1402 1692 1403
rect 1870 1407 1876 1408
rect 1870 1403 1871 1407
rect 1875 1403 1876 1407
rect 2006 1404 2007 1408
rect 2011 1404 2012 1408
rect 2006 1403 2012 1404
rect 1870 1402 1876 1403
rect 407 1399 413 1400
rect 407 1395 408 1399
rect 412 1398 413 1399
rect 551 1399 557 1400
rect 412 1396 505 1398
rect 412 1395 413 1396
rect 407 1394 413 1395
rect 551 1395 552 1399
rect 556 1398 557 1399
rect 670 1399 676 1400
rect 556 1396 625 1398
rect 556 1395 557 1396
rect 551 1394 557 1395
rect 670 1395 671 1399
rect 675 1398 676 1399
rect 799 1399 805 1400
rect 675 1396 753 1398
rect 675 1395 676 1396
rect 670 1394 676 1395
rect 799 1395 800 1399
rect 804 1398 805 1399
rect 938 1399 944 1400
rect 804 1396 897 1398
rect 804 1395 805 1396
rect 799 1394 805 1395
rect 938 1395 939 1399
rect 943 1398 944 1399
rect 1250 1399 1256 1400
rect 943 1396 1049 1398
rect 943 1395 944 1396
rect 938 1394 944 1395
rect 1242 1395 1248 1396
rect 110 1391 116 1392
rect 110 1387 111 1391
rect 115 1387 116 1391
rect 1242 1391 1243 1395
rect 1247 1391 1248 1395
rect 1250 1395 1251 1399
rect 1255 1398 1256 1399
rect 1423 1399 1429 1400
rect 1255 1396 1377 1398
rect 1255 1395 1256 1396
rect 1250 1394 1256 1395
rect 1423 1395 1424 1399
rect 1428 1398 1429 1399
rect 1830 1399 1836 1400
rect 1830 1398 1831 1399
rect 1428 1396 1553 1398
rect 1765 1396 1831 1398
rect 1428 1395 1429 1396
rect 1423 1394 1429 1395
rect 1830 1395 1831 1396
rect 1835 1395 1836 1399
rect 1830 1394 1836 1395
rect 1946 1399 1952 1400
rect 1946 1395 1947 1399
rect 1951 1395 1952 1399
rect 1946 1394 1952 1395
rect 1242 1390 1248 1391
rect 2006 1391 2012 1392
rect 110 1386 116 1387
rect 462 1388 468 1389
rect 462 1384 463 1388
rect 467 1384 468 1388
rect 462 1383 468 1384
rect 582 1388 588 1389
rect 582 1384 583 1388
rect 587 1384 588 1388
rect 582 1383 588 1384
rect 710 1388 716 1389
rect 710 1384 711 1388
rect 715 1384 716 1388
rect 710 1383 716 1384
rect 854 1388 860 1389
rect 854 1384 855 1388
rect 859 1384 860 1388
rect 854 1383 860 1384
rect 1006 1388 1012 1389
rect 1006 1384 1007 1388
rect 1011 1384 1012 1388
rect 1006 1383 1012 1384
rect 1166 1388 1172 1389
rect 1166 1384 1167 1388
rect 1171 1384 1172 1388
rect 1166 1383 1172 1384
rect 1334 1388 1340 1389
rect 1334 1384 1335 1388
rect 1339 1384 1340 1388
rect 1334 1383 1340 1384
rect 1510 1388 1516 1389
rect 1510 1384 1511 1388
rect 1515 1384 1516 1388
rect 1510 1383 1516 1384
rect 1686 1388 1692 1389
rect 1686 1384 1687 1388
rect 1691 1384 1692 1388
rect 1686 1383 1692 1384
rect 1870 1388 1876 1389
rect 1870 1384 1871 1388
rect 1875 1384 1876 1388
rect 2006 1387 2007 1391
rect 2011 1387 2012 1391
rect 2006 1386 2012 1387
rect 1870 1383 1876 1384
rect 2398 1360 2404 1361
rect 2046 1357 2052 1358
rect 2046 1353 2047 1357
rect 2051 1353 2052 1357
rect 2398 1356 2399 1360
rect 2403 1356 2404 1360
rect 2398 1355 2404 1356
rect 2534 1360 2540 1361
rect 2534 1356 2535 1360
rect 2539 1356 2540 1360
rect 2534 1355 2540 1356
rect 2678 1360 2684 1361
rect 2678 1356 2679 1360
rect 2683 1356 2684 1360
rect 2678 1355 2684 1356
rect 2822 1360 2828 1361
rect 2822 1356 2823 1360
rect 2827 1356 2828 1360
rect 2822 1355 2828 1356
rect 2966 1360 2972 1361
rect 2966 1356 2967 1360
rect 2971 1356 2972 1360
rect 2966 1355 2972 1356
rect 3110 1360 3116 1361
rect 3110 1356 3111 1360
rect 3115 1356 3116 1360
rect 3110 1355 3116 1356
rect 3254 1360 3260 1361
rect 3254 1356 3255 1360
rect 3259 1356 3260 1360
rect 3254 1355 3260 1356
rect 3406 1360 3412 1361
rect 3406 1356 3407 1360
rect 3411 1356 3412 1360
rect 3406 1355 3412 1356
rect 3558 1360 3564 1361
rect 3558 1356 3559 1360
rect 3563 1356 3564 1360
rect 3558 1355 3564 1356
rect 3710 1360 3716 1361
rect 3710 1356 3711 1360
rect 3715 1356 3716 1360
rect 3710 1355 3716 1356
rect 3838 1360 3844 1361
rect 3838 1356 3839 1360
rect 3843 1356 3844 1360
rect 3838 1355 3844 1356
rect 3942 1357 3948 1358
rect 2046 1352 2052 1353
rect 3942 1353 3943 1357
rect 3947 1353 3948 1357
rect 3942 1352 3948 1353
rect 2474 1351 2480 1352
rect 2474 1347 2475 1351
rect 2479 1347 2480 1351
rect 2474 1346 2480 1347
rect 2482 1351 2488 1352
rect 2482 1347 2483 1351
rect 2487 1350 2488 1351
rect 2754 1351 2760 1352
rect 2487 1348 2577 1350
rect 2487 1347 2488 1348
rect 2482 1346 2488 1347
rect 2754 1347 2755 1351
rect 2759 1347 2760 1351
rect 2754 1346 2760 1347
rect 2898 1351 2904 1352
rect 2898 1347 2899 1351
rect 2903 1347 2904 1351
rect 2898 1346 2904 1347
rect 2922 1351 2928 1352
rect 2922 1347 2923 1351
rect 2927 1350 2928 1351
rect 3050 1351 3056 1352
rect 2927 1348 3009 1350
rect 2927 1347 2928 1348
rect 2922 1346 2928 1347
rect 3050 1347 3051 1351
rect 3055 1350 3056 1351
rect 3194 1351 3200 1352
rect 3055 1348 3153 1350
rect 3055 1347 3056 1348
rect 3050 1346 3056 1347
rect 3194 1347 3195 1351
rect 3199 1350 3200 1351
rect 3338 1351 3344 1352
rect 3199 1348 3297 1350
rect 3199 1347 3200 1348
rect 3194 1346 3200 1347
rect 3338 1347 3339 1351
rect 3343 1350 3344 1351
rect 3634 1351 3640 1352
rect 3343 1348 3449 1350
rect 3343 1347 3344 1348
rect 3338 1346 3344 1347
rect 3634 1347 3635 1351
rect 3639 1347 3640 1351
rect 3634 1346 3640 1347
rect 3703 1351 3709 1352
rect 3703 1347 3704 1351
rect 3708 1350 3709 1351
rect 3798 1351 3804 1352
rect 3708 1348 3753 1350
rect 3708 1347 3709 1348
rect 3703 1346 3709 1347
rect 3798 1347 3799 1351
rect 3803 1350 3804 1351
rect 3803 1348 3881 1350
rect 3803 1347 3804 1348
rect 3798 1346 3804 1347
rect 2398 1341 2404 1342
rect 2046 1340 2052 1341
rect 2046 1336 2047 1340
rect 2051 1336 2052 1340
rect 2398 1337 2399 1341
rect 2403 1337 2404 1341
rect 2398 1336 2404 1337
rect 2534 1341 2540 1342
rect 2534 1337 2535 1341
rect 2539 1337 2540 1341
rect 2534 1336 2540 1337
rect 2678 1341 2684 1342
rect 2678 1337 2679 1341
rect 2683 1337 2684 1341
rect 2678 1336 2684 1337
rect 2822 1341 2828 1342
rect 2822 1337 2823 1341
rect 2827 1337 2828 1341
rect 2822 1336 2828 1337
rect 2966 1341 2972 1342
rect 2966 1337 2967 1341
rect 2971 1337 2972 1341
rect 2966 1336 2972 1337
rect 3110 1341 3116 1342
rect 3110 1337 3111 1341
rect 3115 1337 3116 1341
rect 3110 1336 3116 1337
rect 3254 1341 3260 1342
rect 3254 1337 3255 1341
rect 3259 1337 3260 1341
rect 3254 1336 3260 1337
rect 3406 1341 3412 1342
rect 3406 1337 3407 1341
rect 3411 1337 3412 1341
rect 3406 1336 3412 1337
rect 3558 1341 3564 1342
rect 3558 1337 3559 1341
rect 3563 1337 3564 1341
rect 3558 1336 3564 1337
rect 3710 1341 3716 1342
rect 3710 1337 3711 1341
rect 3715 1337 3716 1341
rect 3710 1336 3716 1337
rect 3838 1341 3844 1342
rect 3838 1337 3839 1341
rect 3843 1337 3844 1341
rect 3838 1336 3844 1337
rect 3942 1340 3948 1341
rect 3942 1336 3943 1340
rect 3947 1336 3948 1340
rect 2046 1335 2052 1336
rect 3942 1335 3948 1336
rect 654 1328 660 1329
rect 110 1325 116 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 654 1324 655 1328
rect 659 1324 660 1328
rect 654 1323 660 1324
rect 766 1328 772 1329
rect 766 1324 767 1328
rect 771 1324 772 1328
rect 766 1323 772 1324
rect 886 1328 892 1329
rect 886 1324 887 1328
rect 891 1324 892 1328
rect 886 1323 892 1324
rect 1014 1328 1020 1329
rect 1014 1324 1015 1328
rect 1019 1324 1020 1328
rect 1014 1323 1020 1324
rect 1142 1328 1148 1329
rect 1142 1324 1143 1328
rect 1147 1324 1148 1328
rect 1142 1323 1148 1324
rect 1278 1328 1284 1329
rect 1278 1324 1279 1328
rect 1283 1324 1284 1328
rect 1278 1323 1284 1324
rect 1414 1328 1420 1329
rect 1414 1324 1415 1328
rect 1419 1324 1420 1328
rect 1414 1323 1420 1324
rect 1558 1328 1564 1329
rect 1558 1324 1559 1328
rect 1563 1324 1564 1328
rect 1558 1323 1564 1324
rect 1702 1328 1708 1329
rect 1702 1324 1703 1328
rect 1707 1324 1708 1328
rect 1702 1323 1708 1324
rect 1846 1328 1852 1329
rect 1846 1324 1847 1328
rect 1851 1324 1852 1328
rect 2922 1327 2928 1328
rect 2922 1326 2923 1327
rect 1846 1323 1852 1324
rect 2006 1325 2012 1326
rect 110 1320 116 1321
rect 2006 1321 2007 1325
rect 2011 1321 2012 1325
rect 2006 1320 2012 1321
rect 2700 1324 2923 1326
rect 730 1319 736 1320
rect 730 1315 731 1319
rect 735 1315 736 1319
rect 730 1314 736 1315
rect 842 1319 848 1320
rect 842 1315 843 1319
rect 847 1315 848 1319
rect 842 1314 848 1315
rect 962 1319 968 1320
rect 962 1315 963 1319
rect 967 1315 968 1319
rect 962 1314 968 1315
rect 1090 1319 1096 1320
rect 1090 1315 1091 1319
rect 1095 1315 1096 1319
rect 1090 1314 1096 1315
rect 1114 1319 1120 1320
rect 1114 1315 1115 1319
rect 1119 1318 1120 1319
rect 1354 1319 1360 1320
rect 1119 1316 1185 1318
rect 1119 1315 1120 1316
rect 1114 1314 1120 1315
rect 1354 1315 1355 1319
rect 1359 1315 1360 1319
rect 1354 1314 1360 1315
rect 1482 1319 1488 1320
rect 1482 1315 1483 1319
rect 1487 1315 1488 1319
rect 1482 1314 1488 1315
rect 1634 1319 1640 1320
rect 1634 1315 1635 1319
rect 1639 1315 1640 1319
rect 1634 1314 1640 1315
rect 1778 1319 1784 1320
rect 1778 1315 1779 1319
rect 1783 1315 1784 1319
rect 1778 1314 1784 1315
rect 1822 1319 1828 1320
rect 1822 1315 1823 1319
rect 1827 1318 1828 1319
rect 2463 1319 2469 1320
rect 1827 1316 1889 1318
rect 1827 1315 1828 1316
rect 1822 1314 1828 1315
rect 2463 1315 2464 1319
rect 2468 1318 2469 1319
rect 2482 1319 2488 1320
rect 2482 1318 2483 1319
rect 2468 1316 2483 1318
rect 2468 1315 2469 1316
rect 2463 1314 2469 1315
rect 2482 1315 2483 1316
rect 2487 1315 2488 1319
rect 2482 1314 2488 1315
rect 2599 1319 2605 1320
rect 2599 1315 2600 1319
rect 2604 1318 2605 1319
rect 2700 1318 2702 1324
rect 2922 1323 2923 1324
rect 2927 1323 2928 1327
rect 3703 1327 3709 1328
rect 3703 1326 3704 1327
rect 2922 1322 2928 1323
rect 3576 1324 3704 1326
rect 2604 1316 2702 1318
rect 2706 1319 2712 1320
rect 2604 1315 2605 1316
rect 2599 1314 2605 1315
rect 2706 1315 2707 1319
rect 2711 1318 2712 1319
rect 2743 1319 2749 1320
rect 2743 1318 2744 1319
rect 2711 1316 2744 1318
rect 2711 1315 2712 1316
rect 2706 1314 2712 1315
rect 2743 1315 2744 1316
rect 2748 1315 2749 1319
rect 2743 1314 2749 1315
rect 2754 1319 2760 1320
rect 2754 1315 2755 1319
rect 2759 1318 2760 1319
rect 2887 1319 2893 1320
rect 2887 1318 2888 1319
rect 2759 1316 2888 1318
rect 2759 1315 2760 1316
rect 2754 1314 2760 1315
rect 2887 1315 2888 1316
rect 2892 1315 2893 1319
rect 2887 1314 2893 1315
rect 2898 1319 2904 1320
rect 2898 1315 2899 1319
rect 2903 1318 2904 1319
rect 3031 1319 3037 1320
rect 3031 1318 3032 1319
rect 2903 1316 3032 1318
rect 2903 1315 2904 1316
rect 2898 1314 2904 1315
rect 3031 1315 3032 1316
rect 3036 1315 3037 1319
rect 3031 1314 3037 1315
rect 3175 1319 3181 1320
rect 3175 1315 3176 1319
rect 3180 1318 3181 1319
rect 3194 1319 3200 1320
rect 3194 1318 3195 1319
rect 3180 1316 3195 1318
rect 3180 1315 3181 1316
rect 3175 1314 3181 1315
rect 3194 1315 3195 1316
rect 3199 1315 3200 1319
rect 3194 1314 3200 1315
rect 3319 1319 3325 1320
rect 3319 1315 3320 1319
rect 3324 1318 3325 1319
rect 3338 1319 3344 1320
rect 3338 1318 3339 1319
rect 3324 1316 3339 1318
rect 3324 1315 3325 1316
rect 3319 1314 3325 1315
rect 3338 1315 3339 1316
rect 3343 1315 3344 1319
rect 3338 1314 3344 1315
rect 3471 1319 3477 1320
rect 3471 1315 3472 1319
rect 3476 1318 3477 1319
rect 3576 1318 3578 1324
rect 3703 1323 3704 1324
rect 3708 1323 3709 1327
rect 3703 1322 3709 1323
rect 3476 1316 3578 1318
rect 3582 1319 3588 1320
rect 3476 1315 3477 1316
rect 3471 1314 3477 1315
rect 3582 1315 3583 1319
rect 3587 1318 3588 1319
rect 3623 1319 3629 1320
rect 3623 1318 3624 1319
rect 3587 1316 3624 1318
rect 3587 1315 3588 1316
rect 3582 1314 3588 1315
rect 3623 1315 3624 1316
rect 3628 1315 3629 1319
rect 3623 1314 3629 1315
rect 3634 1319 3640 1320
rect 3634 1315 3635 1319
rect 3639 1318 3640 1319
rect 3775 1319 3781 1320
rect 3775 1318 3776 1319
rect 3639 1316 3776 1318
rect 3639 1315 3640 1316
rect 3634 1314 3640 1315
rect 3775 1315 3776 1316
rect 3780 1315 3781 1319
rect 3775 1314 3781 1315
rect 3903 1319 3909 1320
rect 3903 1315 3904 1319
rect 3908 1318 3909 1319
rect 3914 1319 3920 1320
rect 3914 1318 3915 1319
rect 3908 1316 3915 1318
rect 3908 1315 3909 1316
rect 3903 1314 3909 1315
rect 3914 1315 3915 1316
rect 3919 1315 3920 1319
rect 3914 1314 3920 1315
rect 654 1309 660 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 654 1305 655 1309
rect 659 1305 660 1309
rect 654 1304 660 1305
rect 766 1309 772 1310
rect 766 1305 767 1309
rect 771 1305 772 1309
rect 766 1304 772 1305
rect 886 1309 892 1310
rect 886 1305 887 1309
rect 891 1305 892 1309
rect 886 1304 892 1305
rect 1014 1309 1020 1310
rect 1014 1305 1015 1309
rect 1019 1305 1020 1309
rect 1014 1304 1020 1305
rect 1142 1309 1148 1310
rect 1142 1305 1143 1309
rect 1147 1305 1148 1309
rect 1142 1304 1148 1305
rect 1278 1309 1284 1310
rect 1278 1305 1279 1309
rect 1283 1305 1284 1309
rect 1278 1304 1284 1305
rect 1414 1309 1420 1310
rect 1414 1305 1415 1309
rect 1419 1305 1420 1309
rect 1414 1304 1420 1305
rect 1558 1309 1564 1310
rect 1558 1305 1559 1309
rect 1563 1305 1564 1309
rect 1558 1304 1564 1305
rect 1702 1309 1708 1310
rect 1702 1305 1703 1309
rect 1707 1305 1708 1309
rect 1702 1304 1708 1305
rect 1846 1309 1852 1310
rect 1846 1305 1847 1309
rect 1851 1305 1852 1309
rect 1846 1304 1852 1305
rect 2006 1308 2012 1309
rect 2006 1304 2007 1308
rect 2011 1304 2012 1308
rect 110 1303 116 1304
rect 2006 1303 2012 1304
rect 2311 1303 2317 1304
rect 2311 1299 2312 1303
rect 2316 1302 2317 1303
rect 2366 1303 2372 1304
rect 2366 1302 2367 1303
rect 2316 1300 2367 1302
rect 2316 1299 2317 1300
rect 2311 1298 2317 1299
rect 2366 1299 2367 1300
rect 2371 1299 2372 1303
rect 2366 1298 2372 1299
rect 2439 1303 2445 1304
rect 2439 1299 2440 1303
rect 2444 1302 2445 1303
rect 2474 1303 2480 1304
rect 2444 1300 2470 1302
rect 2444 1299 2445 1300
rect 2439 1298 2445 1299
rect 2468 1294 2470 1300
rect 2474 1299 2475 1303
rect 2479 1302 2480 1303
rect 2575 1303 2581 1304
rect 2575 1302 2576 1303
rect 2479 1300 2576 1302
rect 2479 1299 2480 1300
rect 2474 1298 2480 1299
rect 2575 1299 2576 1300
rect 2580 1299 2581 1303
rect 2575 1298 2581 1299
rect 2586 1303 2592 1304
rect 2586 1299 2587 1303
rect 2591 1302 2592 1303
rect 2711 1303 2717 1304
rect 2711 1302 2712 1303
rect 2591 1300 2712 1302
rect 2591 1299 2592 1300
rect 2586 1298 2592 1299
rect 2711 1299 2712 1300
rect 2716 1299 2717 1303
rect 2711 1298 2717 1299
rect 2722 1303 2728 1304
rect 2722 1299 2723 1303
rect 2727 1302 2728 1303
rect 2855 1303 2861 1304
rect 2855 1302 2856 1303
rect 2727 1300 2856 1302
rect 2727 1299 2728 1300
rect 2722 1298 2728 1299
rect 2855 1299 2856 1300
rect 2860 1299 2861 1303
rect 2855 1298 2861 1299
rect 3007 1303 3013 1304
rect 3007 1299 3008 1303
rect 3012 1302 3013 1303
rect 3050 1303 3056 1304
rect 3050 1302 3051 1303
rect 3012 1300 3051 1302
rect 3012 1299 3013 1300
rect 3007 1298 3013 1299
rect 3050 1299 3051 1300
rect 3055 1299 3056 1303
rect 3050 1298 3056 1299
rect 3078 1303 3084 1304
rect 3078 1299 3079 1303
rect 3083 1302 3084 1303
rect 3175 1303 3181 1304
rect 3175 1302 3176 1303
rect 3083 1300 3176 1302
rect 3083 1299 3084 1300
rect 3078 1298 3084 1299
rect 3175 1299 3176 1300
rect 3180 1299 3181 1303
rect 3175 1298 3181 1299
rect 3186 1303 3192 1304
rect 3186 1299 3187 1303
rect 3191 1302 3192 1303
rect 3351 1303 3357 1304
rect 3351 1302 3352 1303
rect 3191 1300 3352 1302
rect 3191 1299 3192 1300
rect 3186 1298 3192 1299
rect 3351 1299 3352 1300
rect 3356 1299 3357 1303
rect 3351 1298 3357 1299
rect 3362 1303 3368 1304
rect 3362 1299 3363 1303
rect 3367 1302 3368 1303
rect 3535 1303 3541 1304
rect 3535 1302 3536 1303
rect 3367 1300 3536 1302
rect 3367 1299 3368 1300
rect 3362 1298 3368 1299
rect 3535 1299 3536 1300
rect 3540 1299 3541 1303
rect 3535 1298 3541 1299
rect 3546 1303 3552 1304
rect 3546 1299 3547 1303
rect 3551 1302 3552 1303
rect 3727 1303 3733 1304
rect 3727 1302 3728 1303
rect 3551 1300 3728 1302
rect 3551 1299 3552 1300
rect 3546 1298 3552 1299
rect 3727 1299 3728 1300
rect 3732 1299 3733 1303
rect 3727 1298 3733 1299
rect 3903 1303 3912 1304
rect 3903 1299 3904 1303
rect 3911 1299 3912 1303
rect 3903 1298 3912 1299
rect 2730 1295 2736 1296
rect 2730 1294 2731 1295
rect 2468 1292 2731 1294
rect 2730 1291 2731 1292
rect 2735 1291 2736 1295
rect 2730 1290 2736 1291
rect 719 1287 725 1288
rect 719 1283 720 1287
rect 724 1286 725 1287
rect 730 1287 736 1288
rect 724 1283 726 1286
rect 719 1282 726 1283
rect 730 1283 731 1287
rect 735 1286 736 1287
rect 831 1287 837 1288
rect 831 1286 832 1287
rect 735 1284 832 1286
rect 735 1283 736 1284
rect 730 1282 736 1283
rect 831 1283 832 1284
rect 836 1283 837 1287
rect 831 1282 837 1283
rect 842 1287 848 1288
rect 842 1283 843 1287
rect 847 1286 848 1287
rect 951 1287 957 1288
rect 951 1286 952 1287
rect 847 1284 952 1286
rect 847 1283 848 1284
rect 842 1282 848 1283
rect 951 1283 952 1284
rect 956 1283 957 1287
rect 951 1282 957 1283
rect 962 1287 968 1288
rect 962 1283 963 1287
rect 967 1286 968 1287
rect 1079 1287 1085 1288
rect 1079 1286 1080 1287
rect 967 1284 1080 1286
rect 967 1283 968 1284
rect 962 1282 968 1283
rect 1079 1283 1080 1284
rect 1084 1283 1085 1287
rect 1079 1282 1085 1283
rect 1090 1287 1096 1288
rect 1090 1283 1091 1287
rect 1095 1286 1096 1287
rect 1207 1287 1213 1288
rect 1207 1286 1208 1287
rect 1095 1284 1208 1286
rect 1095 1283 1096 1284
rect 1090 1282 1096 1283
rect 1207 1283 1208 1284
rect 1212 1283 1213 1287
rect 1207 1282 1213 1283
rect 1242 1287 1248 1288
rect 1242 1283 1243 1287
rect 1247 1286 1248 1287
rect 1343 1287 1349 1288
rect 1343 1286 1344 1287
rect 1247 1284 1344 1286
rect 1247 1283 1248 1284
rect 1242 1282 1248 1283
rect 1343 1283 1344 1284
rect 1348 1283 1349 1287
rect 1343 1282 1349 1283
rect 1354 1287 1360 1288
rect 1354 1283 1355 1287
rect 1359 1286 1360 1287
rect 1479 1287 1485 1288
rect 1479 1286 1480 1287
rect 1359 1284 1480 1286
rect 1359 1283 1360 1284
rect 1354 1282 1360 1283
rect 1479 1283 1480 1284
rect 1484 1283 1485 1287
rect 1479 1282 1485 1283
rect 1623 1287 1632 1288
rect 1623 1283 1624 1287
rect 1631 1283 1632 1287
rect 1623 1282 1632 1283
rect 1634 1287 1640 1288
rect 1634 1283 1635 1287
rect 1639 1286 1640 1287
rect 1767 1287 1773 1288
rect 1767 1286 1768 1287
rect 1639 1284 1768 1286
rect 1639 1283 1640 1284
rect 1634 1282 1640 1283
rect 1767 1283 1768 1284
rect 1772 1283 1773 1287
rect 1767 1282 1773 1283
rect 1778 1287 1784 1288
rect 1778 1283 1779 1287
rect 1783 1286 1784 1287
rect 1911 1287 1917 1288
rect 1911 1286 1912 1287
rect 1783 1284 1912 1286
rect 1783 1283 1784 1284
rect 1778 1282 1784 1283
rect 1911 1283 1912 1284
rect 1916 1283 1917 1287
rect 1911 1282 1917 1283
rect 2046 1284 2052 1285
rect 3942 1284 3948 1285
rect 724 1278 726 1282
rect 2046 1280 2047 1284
rect 2051 1280 2052 1284
rect 887 1279 893 1280
rect 2046 1279 2052 1280
rect 2246 1283 2252 1284
rect 2246 1279 2247 1283
rect 2251 1279 2252 1283
rect 887 1278 888 1279
rect 724 1276 888 1278
rect 887 1275 888 1276
rect 892 1275 893 1279
rect 2246 1278 2252 1279
rect 2374 1283 2380 1284
rect 2374 1279 2375 1283
rect 2379 1279 2380 1283
rect 2374 1278 2380 1279
rect 2510 1283 2516 1284
rect 2510 1279 2511 1283
rect 2515 1279 2516 1283
rect 2510 1278 2516 1279
rect 2646 1283 2652 1284
rect 2646 1279 2647 1283
rect 2651 1279 2652 1283
rect 2646 1278 2652 1279
rect 2790 1283 2796 1284
rect 2790 1279 2791 1283
rect 2795 1279 2796 1283
rect 2790 1278 2796 1279
rect 2942 1283 2948 1284
rect 2942 1279 2943 1283
rect 2947 1279 2948 1283
rect 2942 1278 2948 1279
rect 3110 1283 3116 1284
rect 3110 1279 3111 1283
rect 3115 1279 3116 1283
rect 3110 1278 3116 1279
rect 3286 1283 3292 1284
rect 3286 1279 3287 1283
rect 3291 1279 3292 1283
rect 3286 1278 3292 1279
rect 3470 1283 3476 1284
rect 3470 1279 3471 1283
rect 3475 1279 3476 1283
rect 3470 1278 3476 1279
rect 3662 1283 3668 1284
rect 3662 1279 3663 1283
rect 3667 1279 3668 1283
rect 3662 1278 3668 1279
rect 3838 1283 3844 1284
rect 3838 1279 3839 1283
rect 3843 1279 3844 1283
rect 3942 1280 3943 1284
rect 3947 1280 3948 1284
rect 3942 1279 3948 1280
rect 3838 1278 3844 1279
rect 887 1274 893 1275
rect 2366 1275 2372 1276
rect 503 1271 509 1272
rect 503 1267 504 1271
rect 508 1270 509 1271
rect 514 1271 520 1272
rect 508 1267 510 1270
rect 503 1266 510 1267
rect 514 1267 515 1271
rect 519 1270 520 1271
rect 615 1271 621 1272
rect 615 1270 616 1271
rect 519 1268 616 1270
rect 519 1267 520 1268
rect 514 1266 520 1267
rect 615 1267 616 1268
rect 620 1267 621 1271
rect 615 1266 621 1267
rect 626 1271 632 1272
rect 626 1267 627 1271
rect 631 1270 632 1271
rect 735 1271 741 1272
rect 735 1270 736 1271
rect 631 1268 736 1270
rect 631 1267 632 1268
rect 626 1266 632 1267
rect 735 1267 736 1268
rect 740 1267 741 1271
rect 735 1266 741 1267
rect 746 1271 752 1272
rect 746 1267 747 1271
rect 751 1270 752 1271
rect 863 1271 869 1272
rect 863 1270 864 1271
rect 751 1268 864 1270
rect 751 1267 752 1268
rect 746 1266 752 1267
rect 863 1267 864 1268
rect 868 1267 869 1271
rect 863 1266 869 1267
rect 874 1271 880 1272
rect 874 1267 875 1271
rect 879 1270 880 1271
rect 999 1271 1005 1272
rect 999 1270 1000 1271
rect 879 1268 1000 1270
rect 879 1267 880 1268
rect 874 1266 880 1267
rect 999 1267 1000 1268
rect 1004 1267 1005 1271
rect 999 1266 1005 1267
rect 1143 1271 1149 1272
rect 1143 1267 1144 1271
rect 1148 1270 1149 1271
rect 1214 1271 1220 1272
rect 1214 1270 1215 1271
rect 1148 1268 1215 1270
rect 1148 1267 1149 1268
rect 1143 1266 1149 1267
rect 1214 1267 1215 1268
rect 1219 1267 1220 1271
rect 1214 1266 1220 1267
rect 1295 1271 1301 1272
rect 1295 1267 1296 1271
rect 1300 1270 1301 1271
rect 1314 1271 1320 1272
rect 1314 1270 1315 1271
rect 1300 1268 1315 1270
rect 1300 1267 1301 1268
rect 1295 1266 1301 1267
rect 1314 1267 1315 1268
rect 1319 1267 1320 1271
rect 1314 1266 1320 1267
rect 1455 1271 1461 1272
rect 1455 1267 1456 1271
rect 1460 1270 1461 1271
rect 1482 1271 1488 1272
rect 1482 1270 1483 1271
rect 1460 1268 1483 1270
rect 1460 1267 1461 1268
rect 1455 1266 1461 1267
rect 1482 1267 1483 1268
rect 1487 1267 1488 1271
rect 1482 1266 1488 1267
rect 1615 1271 1621 1272
rect 1615 1267 1616 1271
rect 1620 1270 1621 1271
rect 1639 1271 1645 1272
rect 1639 1270 1640 1271
rect 1620 1268 1640 1270
rect 1620 1267 1621 1268
rect 1615 1266 1621 1267
rect 1639 1267 1640 1268
rect 1644 1267 1645 1271
rect 1639 1266 1645 1267
rect 1770 1271 1776 1272
rect 1770 1267 1771 1271
rect 1775 1270 1776 1271
rect 1783 1271 1789 1272
rect 1783 1270 1784 1271
rect 1775 1268 1784 1270
rect 1775 1267 1776 1268
rect 1770 1266 1776 1267
rect 1783 1267 1784 1268
rect 1788 1267 1789 1271
rect 2322 1271 2328 1272
rect 1783 1266 1789 1267
rect 2046 1267 2052 1268
rect 508 1262 510 1266
rect 738 1263 744 1264
rect 738 1262 739 1263
rect 508 1260 739 1262
rect 738 1259 739 1260
rect 743 1259 744 1263
rect 2046 1263 2047 1267
rect 2051 1263 2052 1267
rect 2322 1267 2323 1271
rect 2327 1267 2328 1271
rect 2366 1271 2367 1275
rect 2371 1274 2372 1275
rect 2586 1275 2592 1276
rect 2371 1272 2417 1274
rect 2371 1271 2372 1272
rect 2366 1270 2372 1271
rect 2586 1271 2587 1275
rect 2591 1271 2592 1275
rect 2586 1270 2592 1271
rect 2722 1275 2728 1276
rect 2722 1271 2723 1275
rect 2727 1271 2728 1275
rect 2722 1270 2728 1271
rect 2730 1275 2736 1276
rect 2730 1271 2731 1275
rect 2735 1274 2736 1275
rect 3078 1275 3084 1276
rect 3078 1274 3079 1275
rect 2735 1272 2833 1274
rect 3021 1272 3079 1274
rect 2735 1271 2736 1272
rect 2730 1270 2736 1271
rect 3078 1271 3079 1272
rect 3083 1271 3084 1275
rect 3078 1270 3084 1271
rect 3186 1275 3192 1276
rect 3186 1271 3187 1275
rect 3191 1271 3192 1275
rect 3186 1270 3192 1271
rect 3362 1275 3368 1276
rect 3362 1271 3363 1275
rect 3367 1271 3368 1275
rect 3362 1270 3368 1271
rect 3546 1275 3552 1276
rect 3546 1271 3547 1275
rect 3551 1271 3552 1275
rect 3546 1270 3552 1271
rect 3610 1275 3616 1276
rect 3610 1271 3611 1275
rect 3615 1274 3616 1275
rect 3914 1275 3920 1276
rect 3615 1272 3705 1274
rect 3615 1271 3616 1272
rect 3610 1270 3616 1271
rect 3914 1271 3915 1275
rect 3919 1271 3920 1275
rect 3914 1270 3920 1271
rect 2322 1266 2328 1267
rect 3942 1267 3948 1268
rect 2046 1262 2052 1263
rect 2246 1264 2252 1265
rect 2246 1260 2247 1264
rect 2251 1260 2252 1264
rect 2246 1259 2252 1260
rect 2374 1264 2380 1265
rect 2374 1260 2375 1264
rect 2379 1260 2380 1264
rect 2374 1259 2380 1260
rect 2510 1264 2516 1265
rect 2510 1260 2511 1264
rect 2515 1260 2516 1264
rect 2510 1259 2516 1260
rect 2646 1264 2652 1265
rect 2646 1260 2647 1264
rect 2651 1260 2652 1264
rect 2646 1259 2652 1260
rect 2790 1264 2796 1265
rect 2790 1260 2791 1264
rect 2795 1260 2796 1264
rect 2790 1259 2796 1260
rect 2942 1264 2948 1265
rect 2942 1260 2943 1264
rect 2947 1260 2948 1264
rect 2942 1259 2948 1260
rect 3110 1264 3116 1265
rect 3110 1260 3111 1264
rect 3115 1260 3116 1264
rect 3110 1259 3116 1260
rect 3286 1264 3292 1265
rect 3286 1260 3287 1264
rect 3291 1260 3292 1264
rect 3286 1259 3292 1260
rect 3470 1264 3476 1265
rect 3470 1260 3471 1264
rect 3475 1260 3476 1264
rect 3470 1259 3476 1260
rect 3662 1264 3668 1265
rect 3662 1260 3663 1264
rect 3667 1260 3668 1264
rect 3662 1259 3668 1260
rect 3838 1264 3844 1265
rect 3838 1260 3839 1264
rect 3843 1260 3844 1264
rect 3942 1263 3943 1267
rect 3947 1263 3948 1267
rect 3942 1262 3948 1263
rect 3838 1259 3844 1260
rect 738 1258 744 1259
rect 110 1252 116 1253
rect 2006 1252 2012 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 438 1251 444 1252
rect 438 1247 439 1251
rect 443 1247 444 1251
rect 438 1246 444 1247
rect 550 1251 556 1252
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 550 1246 556 1247
rect 670 1251 676 1252
rect 670 1247 671 1251
rect 675 1247 676 1251
rect 670 1246 676 1247
rect 798 1251 804 1252
rect 798 1247 799 1251
rect 803 1247 804 1251
rect 798 1246 804 1247
rect 934 1251 940 1252
rect 934 1247 935 1251
rect 939 1247 940 1251
rect 934 1246 940 1247
rect 1078 1251 1084 1252
rect 1078 1247 1079 1251
rect 1083 1247 1084 1251
rect 1078 1246 1084 1247
rect 1230 1251 1236 1252
rect 1230 1247 1231 1251
rect 1235 1247 1236 1251
rect 1230 1246 1236 1247
rect 1390 1251 1396 1252
rect 1390 1247 1391 1251
rect 1395 1247 1396 1251
rect 1390 1246 1396 1247
rect 1550 1251 1556 1252
rect 1550 1247 1551 1251
rect 1555 1247 1556 1251
rect 1550 1246 1556 1247
rect 1718 1251 1724 1252
rect 1718 1247 1719 1251
rect 1723 1247 1724 1251
rect 2006 1248 2007 1252
rect 2011 1248 2012 1252
rect 2006 1247 2012 1248
rect 1718 1246 1724 1247
rect 514 1243 520 1244
rect 514 1239 515 1243
rect 519 1239 520 1243
rect 514 1238 520 1239
rect 626 1243 632 1244
rect 626 1239 627 1243
rect 631 1239 632 1243
rect 626 1238 632 1239
rect 746 1243 752 1244
rect 746 1239 747 1243
rect 751 1239 752 1243
rect 746 1238 752 1239
rect 874 1243 880 1244
rect 874 1239 875 1243
rect 879 1239 880 1243
rect 874 1238 880 1239
rect 887 1243 893 1244
rect 887 1239 888 1243
rect 892 1242 893 1243
rect 1070 1243 1076 1244
rect 892 1240 977 1242
rect 892 1239 893 1240
rect 887 1238 893 1239
rect 1070 1239 1071 1243
rect 1075 1242 1076 1243
rect 1214 1243 1220 1244
rect 1075 1240 1121 1242
rect 1075 1239 1076 1240
rect 1070 1238 1076 1239
rect 1214 1239 1215 1243
rect 1219 1242 1220 1243
rect 1314 1243 1320 1244
rect 1219 1240 1273 1242
rect 1219 1239 1220 1240
rect 1214 1238 1220 1239
rect 1314 1239 1315 1243
rect 1319 1242 1320 1243
rect 1626 1243 1632 1244
rect 1319 1240 1433 1242
rect 1319 1239 1320 1240
rect 1314 1238 1320 1239
rect 1626 1239 1627 1243
rect 1631 1239 1632 1243
rect 1626 1238 1632 1239
rect 1639 1243 1645 1244
rect 1639 1239 1640 1243
rect 1644 1242 1645 1243
rect 1644 1240 1761 1242
rect 1644 1239 1645 1240
rect 1639 1238 1645 1239
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 2006 1235 2012 1236
rect 110 1230 116 1231
rect 438 1232 444 1233
rect 438 1228 439 1232
rect 443 1228 444 1232
rect 438 1227 444 1228
rect 550 1232 556 1233
rect 550 1228 551 1232
rect 555 1228 556 1232
rect 550 1227 556 1228
rect 670 1232 676 1233
rect 670 1228 671 1232
rect 675 1228 676 1232
rect 670 1227 676 1228
rect 798 1232 804 1233
rect 798 1228 799 1232
rect 803 1228 804 1232
rect 798 1227 804 1228
rect 934 1232 940 1233
rect 934 1228 935 1232
rect 939 1228 940 1232
rect 934 1227 940 1228
rect 1078 1232 1084 1233
rect 1078 1228 1079 1232
rect 1083 1228 1084 1232
rect 1078 1227 1084 1228
rect 1230 1232 1236 1233
rect 1230 1228 1231 1232
rect 1235 1228 1236 1232
rect 1230 1227 1236 1228
rect 1390 1232 1396 1233
rect 1390 1228 1391 1232
rect 1395 1228 1396 1232
rect 1390 1227 1396 1228
rect 1550 1232 1556 1233
rect 1550 1228 1551 1232
rect 1555 1228 1556 1232
rect 1550 1227 1556 1228
rect 1718 1232 1724 1233
rect 1718 1228 1719 1232
rect 1723 1228 1724 1232
rect 2006 1231 2007 1235
rect 2011 1231 2012 1235
rect 2006 1230 2012 1231
rect 1718 1227 1724 1228
rect 2070 1200 2076 1201
rect 2046 1197 2052 1198
rect 2046 1193 2047 1197
rect 2051 1193 2052 1197
rect 2070 1196 2071 1200
rect 2075 1196 2076 1200
rect 2070 1195 2076 1196
rect 2182 1200 2188 1201
rect 2182 1196 2183 1200
rect 2187 1196 2188 1200
rect 2182 1195 2188 1196
rect 2302 1200 2308 1201
rect 2302 1196 2303 1200
rect 2307 1196 2308 1200
rect 2302 1195 2308 1196
rect 2430 1200 2436 1201
rect 2430 1196 2431 1200
rect 2435 1196 2436 1200
rect 2430 1195 2436 1196
rect 2558 1200 2564 1201
rect 2558 1196 2559 1200
rect 2563 1196 2564 1200
rect 2558 1195 2564 1196
rect 2710 1200 2716 1201
rect 2710 1196 2711 1200
rect 2715 1196 2716 1200
rect 2710 1195 2716 1196
rect 2886 1200 2892 1201
rect 2886 1196 2887 1200
rect 2891 1196 2892 1200
rect 2886 1195 2892 1196
rect 3086 1200 3092 1201
rect 3086 1196 3087 1200
rect 3091 1196 3092 1200
rect 3086 1195 3092 1196
rect 3310 1200 3316 1201
rect 3310 1196 3311 1200
rect 3315 1196 3316 1200
rect 3310 1195 3316 1196
rect 3542 1200 3548 1201
rect 3542 1196 3543 1200
rect 3547 1196 3548 1200
rect 3542 1195 3548 1196
rect 3782 1200 3788 1201
rect 3782 1196 3783 1200
rect 3787 1196 3788 1200
rect 3782 1195 3788 1196
rect 3942 1197 3948 1198
rect 2046 1192 2052 1193
rect 3942 1193 3943 1197
rect 3947 1193 3948 1197
rect 3942 1192 3948 1193
rect 2146 1191 2152 1192
rect 2146 1187 2147 1191
rect 2151 1187 2152 1191
rect 2146 1186 2152 1187
rect 2258 1191 2264 1192
rect 2258 1187 2259 1191
rect 2263 1187 2264 1191
rect 2258 1186 2264 1187
rect 2378 1191 2384 1192
rect 2378 1187 2379 1191
rect 2383 1187 2384 1191
rect 2378 1186 2384 1187
rect 2506 1191 2512 1192
rect 2506 1187 2507 1191
rect 2511 1187 2512 1191
rect 2506 1186 2512 1187
rect 2514 1191 2520 1192
rect 2514 1187 2515 1191
rect 2519 1190 2520 1191
rect 2778 1191 2784 1192
rect 2519 1188 2601 1190
rect 2519 1187 2520 1188
rect 2514 1186 2520 1187
rect 2778 1187 2779 1191
rect 2783 1187 2784 1191
rect 2778 1186 2784 1187
rect 2794 1191 2800 1192
rect 2794 1187 2795 1191
rect 2799 1190 2800 1191
rect 2970 1191 2976 1192
rect 2799 1188 2929 1190
rect 2799 1187 2800 1188
rect 2794 1186 2800 1187
rect 2970 1187 2971 1191
rect 2975 1190 2976 1191
rect 3170 1191 3176 1192
rect 2975 1188 3129 1190
rect 2975 1187 2976 1188
rect 2970 1186 2976 1187
rect 3170 1187 3171 1191
rect 3175 1190 3176 1191
rect 3394 1191 3400 1192
rect 3175 1188 3353 1190
rect 3175 1187 3176 1188
rect 3170 1186 3176 1187
rect 3394 1187 3395 1191
rect 3399 1190 3400 1191
rect 3858 1191 3864 1192
rect 3399 1188 3585 1190
rect 3399 1187 3400 1188
rect 3394 1186 3400 1187
rect 3858 1187 3859 1191
rect 3863 1187 3864 1191
rect 3858 1186 3864 1187
rect 2070 1181 2076 1182
rect 2046 1180 2052 1181
rect 2046 1176 2047 1180
rect 2051 1176 2052 1180
rect 2070 1177 2071 1181
rect 2075 1177 2076 1181
rect 2070 1176 2076 1177
rect 2182 1181 2188 1182
rect 2182 1177 2183 1181
rect 2187 1177 2188 1181
rect 2182 1176 2188 1177
rect 2302 1181 2308 1182
rect 2302 1177 2303 1181
rect 2307 1177 2308 1181
rect 2302 1176 2308 1177
rect 2430 1181 2436 1182
rect 2430 1177 2431 1181
rect 2435 1177 2436 1181
rect 2430 1176 2436 1177
rect 2558 1181 2564 1182
rect 2558 1177 2559 1181
rect 2563 1177 2564 1181
rect 2558 1176 2564 1177
rect 2710 1181 2716 1182
rect 2710 1177 2711 1181
rect 2715 1177 2716 1181
rect 2710 1176 2716 1177
rect 2886 1181 2892 1182
rect 2886 1177 2887 1181
rect 2891 1177 2892 1181
rect 2886 1176 2892 1177
rect 3086 1181 3092 1182
rect 3086 1177 3087 1181
rect 3091 1177 3092 1181
rect 3086 1176 3092 1177
rect 3310 1181 3316 1182
rect 3310 1177 3311 1181
rect 3315 1177 3316 1181
rect 3310 1176 3316 1177
rect 3542 1181 3548 1182
rect 3542 1177 3543 1181
rect 3547 1177 3548 1181
rect 3542 1176 3548 1177
rect 3782 1181 3788 1182
rect 3782 1177 3783 1181
rect 3787 1177 3788 1181
rect 3782 1176 3788 1177
rect 3942 1180 3948 1181
rect 3942 1176 3943 1180
rect 3947 1176 3948 1180
rect 2046 1175 2052 1176
rect 3942 1175 3948 1176
rect 166 1172 172 1173
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 166 1168 167 1172
rect 171 1168 172 1172
rect 166 1167 172 1168
rect 302 1172 308 1173
rect 302 1168 303 1172
rect 307 1168 308 1172
rect 302 1167 308 1168
rect 462 1172 468 1173
rect 462 1168 463 1172
rect 467 1168 468 1172
rect 462 1167 468 1168
rect 630 1172 636 1173
rect 630 1168 631 1172
rect 635 1168 636 1172
rect 630 1167 636 1168
rect 806 1172 812 1173
rect 806 1168 807 1172
rect 811 1168 812 1172
rect 806 1167 812 1168
rect 982 1172 988 1173
rect 982 1168 983 1172
rect 987 1168 988 1172
rect 982 1167 988 1168
rect 1158 1172 1164 1173
rect 1158 1168 1159 1172
rect 1163 1168 1164 1172
rect 1158 1167 1164 1168
rect 1334 1172 1340 1173
rect 1334 1168 1335 1172
rect 1339 1168 1340 1172
rect 1334 1167 1340 1168
rect 1510 1172 1516 1173
rect 1510 1168 1511 1172
rect 1515 1168 1516 1172
rect 1510 1167 1516 1168
rect 1694 1172 1700 1173
rect 1694 1168 1695 1172
rect 1699 1168 1700 1172
rect 1694 1167 1700 1168
rect 2006 1169 2012 1170
rect 110 1164 116 1165
rect 2006 1165 2007 1169
rect 2011 1165 2012 1169
rect 2514 1167 2520 1168
rect 2514 1166 2515 1167
rect 2006 1164 2012 1165
rect 2137 1164 2515 1166
rect 242 1163 248 1164
rect 242 1159 243 1163
rect 247 1159 248 1163
rect 242 1158 248 1159
rect 378 1163 384 1164
rect 378 1159 379 1163
rect 383 1159 384 1163
rect 378 1158 384 1159
rect 538 1163 544 1164
rect 538 1159 539 1163
rect 543 1159 544 1163
rect 538 1158 544 1159
rect 706 1163 712 1164
rect 706 1159 707 1163
rect 711 1159 712 1163
rect 706 1158 712 1159
rect 738 1163 744 1164
rect 738 1159 739 1163
rect 743 1162 744 1163
rect 1122 1163 1128 1164
rect 1122 1162 1123 1163
rect 743 1160 849 1162
rect 1061 1160 1123 1162
rect 743 1159 744 1160
rect 738 1158 744 1159
rect 1122 1159 1123 1160
rect 1127 1159 1128 1163
rect 1122 1158 1128 1159
rect 1234 1163 1240 1164
rect 1234 1159 1235 1163
rect 1239 1159 1240 1163
rect 1234 1158 1240 1159
rect 1410 1163 1416 1164
rect 1410 1159 1411 1163
rect 1415 1159 1416 1163
rect 1410 1158 1416 1159
rect 1586 1163 1592 1164
rect 1586 1159 1587 1163
rect 1591 1159 1592 1163
rect 1586 1158 1592 1159
rect 1770 1163 1776 1164
rect 1770 1159 1771 1163
rect 1775 1159 1776 1163
rect 2137 1160 2139 1164
rect 2514 1163 2515 1164
rect 2519 1163 2520 1167
rect 2514 1162 2520 1163
rect 1770 1158 1776 1159
rect 2135 1159 2141 1160
rect 2135 1155 2136 1159
rect 2140 1155 2141 1159
rect 2135 1154 2141 1155
rect 2146 1159 2152 1160
rect 2146 1155 2147 1159
rect 2151 1158 2152 1159
rect 2247 1159 2253 1160
rect 2247 1158 2248 1159
rect 2151 1156 2248 1158
rect 2151 1155 2152 1156
rect 2146 1154 2152 1155
rect 2247 1155 2248 1156
rect 2252 1155 2253 1159
rect 2247 1154 2253 1155
rect 2322 1159 2328 1160
rect 2322 1155 2323 1159
rect 2327 1158 2328 1159
rect 2367 1159 2373 1160
rect 2367 1158 2368 1159
rect 2327 1156 2368 1158
rect 2327 1155 2328 1156
rect 2322 1154 2328 1155
rect 2367 1155 2368 1156
rect 2372 1155 2373 1159
rect 2367 1154 2373 1155
rect 2378 1159 2384 1160
rect 2378 1155 2379 1159
rect 2383 1158 2384 1159
rect 2495 1159 2501 1160
rect 2495 1158 2496 1159
rect 2383 1156 2496 1158
rect 2383 1155 2384 1156
rect 2378 1154 2384 1155
rect 2495 1155 2496 1156
rect 2500 1155 2501 1159
rect 2495 1154 2501 1155
rect 2506 1159 2512 1160
rect 2506 1155 2507 1159
rect 2511 1158 2512 1159
rect 2623 1159 2629 1160
rect 2623 1158 2624 1159
rect 2511 1156 2624 1158
rect 2511 1155 2512 1156
rect 2506 1154 2512 1155
rect 2623 1155 2624 1156
rect 2628 1155 2629 1159
rect 2623 1154 2629 1155
rect 2775 1159 2781 1160
rect 2775 1155 2776 1159
rect 2780 1158 2781 1159
rect 2794 1159 2800 1160
rect 2794 1158 2795 1159
rect 2780 1156 2795 1158
rect 2780 1155 2781 1156
rect 2775 1154 2781 1155
rect 2794 1155 2795 1156
rect 2799 1155 2800 1159
rect 2794 1154 2800 1155
rect 2951 1159 2957 1160
rect 2951 1155 2952 1159
rect 2956 1158 2957 1159
rect 2970 1159 2976 1160
rect 2970 1158 2971 1159
rect 2956 1156 2971 1158
rect 2956 1155 2957 1156
rect 2951 1154 2957 1155
rect 2970 1155 2971 1156
rect 2975 1155 2976 1159
rect 2970 1154 2976 1155
rect 3151 1159 3157 1160
rect 3151 1155 3152 1159
rect 3156 1158 3157 1159
rect 3170 1159 3176 1160
rect 3170 1158 3171 1159
rect 3156 1156 3171 1158
rect 3156 1155 3157 1156
rect 3151 1154 3157 1155
rect 3170 1155 3171 1156
rect 3175 1155 3176 1159
rect 3170 1154 3176 1155
rect 3375 1159 3381 1160
rect 3375 1155 3376 1159
rect 3380 1158 3381 1159
rect 3394 1159 3400 1160
rect 3394 1158 3395 1159
rect 3380 1156 3395 1158
rect 3380 1155 3381 1156
rect 3375 1154 3381 1155
rect 3394 1155 3395 1156
rect 3399 1155 3400 1159
rect 3394 1154 3400 1155
rect 3607 1159 3616 1160
rect 3607 1155 3608 1159
rect 3615 1155 3616 1159
rect 3607 1154 3616 1155
rect 3754 1159 3760 1160
rect 3754 1155 3755 1159
rect 3759 1158 3760 1159
rect 3847 1159 3853 1160
rect 3847 1158 3848 1159
rect 3759 1156 3848 1158
rect 3759 1155 3760 1156
rect 3754 1154 3760 1155
rect 3847 1155 3848 1156
rect 3852 1155 3853 1159
rect 3847 1154 3853 1155
rect 166 1153 172 1154
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 166 1149 167 1153
rect 171 1149 172 1153
rect 166 1148 172 1149
rect 302 1153 308 1154
rect 302 1149 303 1153
rect 307 1149 308 1153
rect 302 1148 308 1149
rect 462 1153 468 1154
rect 462 1149 463 1153
rect 467 1149 468 1153
rect 462 1148 468 1149
rect 630 1153 636 1154
rect 630 1149 631 1153
rect 635 1149 636 1153
rect 630 1148 636 1149
rect 806 1153 812 1154
rect 806 1149 807 1153
rect 811 1149 812 1153
rect 806 1148 812 1149
rect 982 1153 988 1154
rect 982 1149 983 1153
rect 987 1149 988 1153
rect 982 1148 988 1149
rect 1158 1153 1164 1154
rect 1158 1149 1159 1153
rect 1163 1149 1164 1153
rect 1158 1148 1164 1149
rect 1334 1153 1340 1154
rect 1334 1149 1335 1153
rect 1339 1149 1340 1153
rect 1334 1148 1340 1149
rect 1510 1153 1516 1154
rect 1510 1149 1511 1153
rect 1515 1149 1516 1153
rect 1510 1148 1516 1149
rect 1694 1153 1700 1154
rect 1694 1149 1695 1153
rect 1699 1149 1700 1153
rect 1694 1148 1700 1149
rect 2006 1152 2012 1153
rect 2006 1148 2007 1152
rect 2011 1148 2012 1152
rect 110 1147 116 1148
rect 2006 1147 2012 1148
rect 2135 1143 2141 1144
rect 2135 1139 2136 1143
rect 2140 1139 2141 1143
rect 2135 1138 2141 1139
rect 2258 1143 2269 1144
rect 2258 1139 2259 1143
rect 2263 1139 2264 1143
rect 2268 1139 2269 1143
rect 2258 1138 2269 1139
rect 2274 1143 2280 1144
rect 2274 1139 2275 1143
rect 2279 1142 2280 1143
rect 2415 1143 2421 1144
rect 2415 1142 2416 1143
rect 2279 1140 2416 1142
rect 2279 1139 2280 1140
rect 2274 1138 2280 1139
rect 2415 1139 2416 1140
rect 2420 1139 2421 1143
rect 2415 1138 2421 1139
rect 2482 1143 2488 1144
rect 2482 1139 2483 1143
rect 2487 1142 2488 1143
rect 2575 1143 2581 1144
rect 2575 1142 2576 1143
rect 2487 1140 2576 1142
rect 2487 1139 2488 1140
rect 2482 1138 2488 1139
rect 2575 1139 2576 1140
rect 2580 1139 2581 1143
rect 2575 1138 2581 1139
rect 2743 1143 2749 1144
rect 2743 1139 2744 1143
rect 2748 1142 2749 1143
rect 2778 1143 2784 1144
rect 2778 1142 2779 1143
rect 2748 1140 2779 1142
rect 2748 1139 2749 1140
rect 2743 1138 2749 1139
rect 2778 1139 2779 1140
rect 2783 1139 2784 1143
rect 2778 1138 2784 1139
rect 2786 1143 2792 1144
rect 2786 1139 2787 1143
rect 2791 1142 2792 1143
rect 2935 1143 2941 1144
rect 2935 1142 2936 1143
rect 2791 1140 2936 1142
rect 2791 1139 2792 1140
rect 2786 1138 2792 1139
rect 2935 1139 2936 1140
rect 2940 1139 2941 1143
rect 2935 1138 2941 1139
rect 2946 1143 2952 1144
rect 2946 1139 2947 1143
rect 2951 1142 2952 1143
rect 3151 1143 3157 1144
rect 3151 1142 3152 1143
rect 2951 1140 3152 1142
rect 2951 1139 2952 1140
rect 2946 1138 2952 1139
rect 3151 1139 3152 1140
rect 3156 1139 3157 1143
rect 3151 1138 3157 1139
rect 3162 1143 3168 1144
rect 3162 1139 3163 1143
rect 3167 1142 3168 1143
rect 3383 1143 3389 1144
rect 3383 1142 3384 1143
rect 3167 1140 3384 1142
rect 3167 1139 3168 1140
rect 3162 1138 3168 1139
rect 3383 1139 3384 1140
rect 3388 1139 3389 1143
rect 3383 1138 3389 1139
rect 3394 1143 3400 1144
rect 3394 1139 3395 1143
rect 3399 1142 3400 1143
rect 3623 1143 3629 1144
rect 3623 1142 3624 1143
rect 3399 1140 3624 1142
rect 3399 1139 3400 1140
rect 3394 1138 3400 1139
rect 3623 1139 3624 1140
rect 3628 1139 3629 1143
rect 3623 1138 3629 1139
rect 3858 1143 3864 1144
rect 3858 1139 3859 1143
rect 3863 1142 3864 1143
rect 3871 1143 3877 1144
rect 3871 1142 3872 1143
rect 3863 1140 3872 1142
rect 3863 1139 3864 1140
rect 3858 1138 3864 1139
rect 3871 1139 3872 1140
rect 3876 1139 3877 1143
rect 3871 1138 3877 1139
rect 2137 1134 2139 1138
rect 2490 1135 2496 1136
rect 2490 1134 2491 1135
rect 2137 1132 2491 1134
rect 231 1131 237 1132
rect 231 1127 232 1131
rect 236 1127 237 1131
rect 231 1126 237 1127
rect 242 1131 248 1132
rect 242 1127 243 1131
rect 247 1130 248 1131
rect 367 1131 373 1132
rect 367 1130 368 1131
rect 247 1128 368 1130
rect 247 1127 248 1128
rect 242 1126 248 1127
rect 367 1127 368 1128
rect 372 1127 373 1131
rect 367 1126 373 1127
rect 378 1131 384 1132
rect 378 1127 379 1131
rect 383 1130 384 1131
rect 527 1131 533 1132
rect 527 1130 528 1131
rect 383 1128 528 1130
rect 383 1127 384 1128
rect 378 1126 384 1127
rect 527 1127 528 1128
rect 532 1127 533 1131
rect 527 1126 533 1127
rect 538 1131 544 1132
rect 538 1127 539 1131
rect 543 1130 544 1131
rect 695 1131 701 1132
rect 695 1130 696 1131
rect 543 1128 696 1130
rect 543 1127 544 1128
rect 538 1126 544 1127
rect 695 1127 696 1128
rect 700 1127 701 1131
rect 695 1126 701 1127
rect 706 1131 712 1132
rect 706 1127 707 1131
rect 711 1130 712 1131
rect 871 1131 877 1132
rect 871 1130 872 1131
rect 711 1128 872 1130
rect 711 1127 712 1128
rect 706 1126 712 1127
rect 871 1127 872 1128
rect 876 1127 877 1131
rect 871 1126 877 1127
rect 1047 1131 1053 1132
rect 1047 1127 1048 1131
rect 1052 1130 1053 1131
rect 1070 1131 1076 1132
rect 1070 1130 1071 1131
rect 1052 1128 1071 1130
rect 1052 1127 1053 1128
rect 1047 1126 1053 1127
rect 1070 1127 1071 1128
rect 1075 1127 1076 1131
rect 1070 1126 1076 1127
rect 1122 1131 1128 1132
rect 1122 1127 1123 1131
rect 1127 1130 1128 1131
rect 1223 1131 1229 1132
rect 1223 1130 1224 1131
rect 1127 1128 1224 1130
rect 1127 1127 1128 1128
rect 1122 1126 1128 1127
rect 1223 1127 1224 1128
rect 1228 1127 1229 1131
rect 1223 1126 1229 1127
rect 1399 1131 1405 1132
rect 1399 1127 1400 1131
rect 1404 1130 1405 1131
rect 1410 1131 1416 1132
rect 1404 1127 1406 1130
rect 1399 1126 1406 1127
rect 1410 1127 1411 1131
rect 1415 1130 1416 1131
rect 1575 1131 1581 1132
rect 1575 1130 1576 1131
rect 1415 1128 1576 1130
rect 1415 1127 1416 1128
rect 1410 1126 1416 1127
rect 1575 1127 1576 1128
rect 1580 1127 1581 1131
rect 1575 1126 1581 1127
rect 1586 1131 1592 1132
rect 1586 1127 1587 1131
rect 1591 1130 1592 1131
rect 1759 1131 1765 1132
rect 1759 1130 1760 1131
rect 1591 1128 1760 1130
rect 1591 1127 1592 1128
rect 1586 1126 1592 1127
rect 1759 1127 1760 1128
rect 1764 1127 1765 1131
rect 2490 1131 2491 1132
rect 2495 1131 2496 1135
rect 2490 1130 2496 1131
rect 1759 1126 1765 1127
rect 233 1122 235 1126
rect 618 1123 624 1124
rect 618 1122 619 1123
rect 233 1120 619 1122
rect 618 1119 619 1120
rect 623 1119 624 1123
rect 1404 1122 1406 1126
rect 2046 1124 2052 1125
rect 3942 1124 3948 1125
rect 1503 1123 1509 1124
rect 1503 1122 1504 1123
rect 1404 1120 1504 1122
rect 618 1118 624 1119
rect 1503 1119 1504 1120
rect 1508 1119 1509 1123
rect 1503 1118 1509 1119
rect 1900 1120 2001 1122
rect 199 1115 208 1116
rect 199 1111 200 1115
rect 207 1111 208 1115
rect 199 1110 208 1111
rect 210 1115 216 1116
rect 210 1111 211 1115
rect 215 1114 216 1115
rect 303 1115 309 1116
rect 303 1114 304 1115
rect 215 1112 304 1114
rect 215 1111 216 1112
rect 210 1110 216 1111
rect 303 1111 304 1112
rect 308 1111 309 1115
rect 303 1110 309 1111
rect 314 1115 320 1116
rect 314 1111 315 1115
rect 319 1114 320 1115
rect 439 1115 445 1116
rect 439 1114 440 1115
rect 319 1112 440 1114
rect 319 1111 320 1112
rect 314 1110 320 1111
rect 439 1111 440 1112
rect 444 1111 445 1115
rect 439 1110 445 1111
rect 450 1115 456 1116
rect 450 1111 451 1115
rect 455 1114 456 1115
rect 591 1115 597 1116
rect 591 1114 592 1115
rect 455 1112 592 1114
rect 455 1111 456 1112
rect 450 1110 456 1111
rect 591 1111 592 1112
rect 596 1111 597 1115
rect 591 1110 597 1111
rect 602 1115 608 1116
rect 602 1111 603 1115
rect 607 1114 608 1115
rect 759 1115 765 1116
rect 759 1114 760 1115
rect 607 1112 760 1114
rect 607 1111 608 1112
rect 602 1110 608 1111
rect 759 1111 760 1112
rect 764 1111 765 1115
rect 759 1110 765 1111
rect 927 1115 933 1116
rect 927 1111 928 1115
rect 932 1114 933 1115
rect 946 1115 952 1116
rect 946 1114 947 1115
rect 932 1112 947 1114
rect 932 1111 933 1112
rect 927 1110 933 1111
rect 946 1111 947 1112
rect 951 1111 952 1115
rect 946 1110 952 1111
rect 1103 1115 1109 1116
rect 1103 1111 1104 1115
rect 1108 1114 1109 1115
rect 1135 1115 1141 1116
rect 1135 1114 1136 1115
rect 1108 1112 1136 1114
rect 1108 1111 1109 1112
rect 1103 1110 1109 1111
rect 1135 1111 1136 1112
rect 1140 1111 1141 1115
rect 1135 1110 1141 1111
rect 1234 1115 1240 1116
rect 1234 1111 1235 1115
rect 1239 1114 1240 1115
rect 1279 1115 1285 1116
rect 1279 1114 1280 1115
rect 1239 1112 1280 1114
rect 1239 1111 1240 1112
rect 1234 1110 1240 1111
rect 1279 1111 1280 1112
rect 1284 1111 1285 1115
rect 1279 1110 1285 1111
rect 1454 1115 1461 1116
rect 1454 1111 1455 1115
rect 1460 1111 1461 1115
rect 1454 1110 1461 1111
rect 1466 1115 1472 1116
rect 1466 1111 1467 1115
rect 1471 1114 1472 1115
rect 1631 1115 1637 1116
rect 1631 1114 1632 1115
rect 1471 1112 1632 1114
rect 1471 1111 1472 1112
rect 1466 1110 1472 1111
rect 1631 1111 1632 1112
rect 1636 1111 1637 1115
rect 1631 1110 1637 1111
rect 1807 1115 1813 1116
rect 1807 1111 1808 1115
rect 1812 1114 1813 1115
rect 1900 1114 1902 1120
rect 1967 1115 1973 1116
rect 1967 1114 1968 1115
rect 1812 1112 1902 1114
rect 1904 1112 1968 1114
rect 1812 1111 1813 1112
rect 1807 1110 1813 1111
rect 1818 1107 1824 1108
rect 1818 1103 1819 1107
rect 1823 1106 1824 1107
rect 1904 1106 1906 1112
rect 1967 1111 1968 1112
rect 1972 1111 1973 1115
rect 1999 1114 2001 1120
rect 2046 1120 2047 1124
rect 2051 1120 2052 1124
rect 2046 1119 2052 1120
rect 2070 1123 2076 1124
rect 2070 1119 2071 1123
rect 2075 1119 2076 1123
rect 2070 1118 2076 1119
rect 2198 1123 2204 1124
rect 2198 1119 2199 1123
rect 2203 1119 2204 1123
rect 2198 1118 2204 1119
rect 2350 1123 2356 1124
rect 2350 1119 2351 1123
rect 2355 1119 2356 1123
rect 2350 1118 2356 1119
rect 2510 1123 2516 1124
rect 2510 1119 2511 1123
rect 2515 1119 2516 1123
rect 2510 1118 2516 1119
rect 2678 1123 2684 1124
rect 2678 1119 2679 1123
rect 2683 1119 2684 1123
rect 2678 1118 2684 1119
rect 2870 1123 2876 1124
rect 2870 1119 2871 1123
rect 2875 1119 2876 1123
rect 2870 1118 2876 1119
rect 3086 1123 3092 1124
rect 3086 1119 3087 1123
rect 3091 1119 3092 1123
rect 3086 1118 3092 1119
rect 3318 1123 3324 1124
rect 3318 1119 3319 1123
rect 3323 1119 3324 1123
rect 3318 1118 3324 1119
rect 3558 1123 3564 1124
rect 3558 1119 3559 1123
rect 3563 1119 3564 1123
rect 3558 1118 3564 1119
rect 3806 1123 3812 1124
rect 3806 1119 3807 1123
rect 3811 1119 3812 1123
rect 3942 1120 3943 1124
rect 3947 1120 3948 1124
rect 3942 1119 3948 1120
rect 3806 1118 3812 1119
rect 2274 1115 2280 1116
rect 1999 1112 2113 1114
rect 1967 1110 1973 1111
rect 2274 1111 2275 1115
rect 2279 1111 2280 1115
rect 2482 1115 2488 1116
rect 2482 1114 2483 1115
rect 2429 1112 2483 1114
rect 2274 1110 2280 1111
rect 2482 1111 2483 1112
rect 2487 1111 2488 1115
rect 2482 1110 2488 1111
rect 2490 1115 2496 1116
rect 2490 1111 2491 1115
rect 2495 1114 2496 1115
rect 2786 1115 2792 1116
rect 2786 1114 2787 1115
rect 2495 1112 2553 1114
rect 2757 1112 2787 1114
rect 2495 1111 2496 1112
rect 2490 1110 2496 1111
rect 2786 1111 2787 1112
rect 2791 1111 2792 1115
rect 2786 1110 2792 1111
rect 2946 1115 2952 1116
rect 2946 1111 2947 1115
rect 2951 1111 2952 1115
rect 2946 1110 2952 1111
rect 3162 1115 3168 1116
rect 3162 1111 3163 1115
rect 3167 1111 3168 1115
rect 3162 1110 3168 1111
rect 3394 1115 3400 1116
rect 3394 1111 3395 1115
rect 3399 1111 3400 1115
rect 3394 1110 3400 1111
rect 3402 1115 3408 1116
rect 3402 1111 3403 1115
rect 3407 1114 3408 1115
rect 3407 1112 3601 1114
rect 3407 1111 3408 1112
rect 3402 1110 3408 1111
rect 3882 1111 3888 1112
rect 1823 1104 1906 1106
rect 2046 1107 2052 1108
rect 1823 1103 1824 1104
rect 1818 1102 1824 1103
rect 2046 1103 2047 1107
rect 2051 1103 2052 1107
rect 3882 1107 3883 1111
rect 3887 1107 3888 1111
rect 3882 1106 3888 1107
rect 3942 1107 3948 1108
rect 2046 1102 2052 1103
rect 2070 1104 2076 1105
rect 2070 1100 2071 1104
rect 2075 1100 2076 1104
rect 2070 1099 2076 1100
rect 2198 1104 2204 1105
rect 2198 1100 2199 1104
rect 2203 1100 2204 1104
rect 2198 1099 2204 1100
rect 2350 1104 2356 1105
rect 2350 1100 2351 1104
rect 2355 1100 2356 1104
rect 2350 1099 2356 1100
rect 2510 1104 2516 1105
rect 2510 1100 2511 1104
rect 2515 1100 2516 1104
rect 2510 1099 2516 1100
rect 2678 1104 2684 1105
rect 2678 1100 2679 1104
rect 2683 1100 2684 1104
rect 2678 1099 2684 1100
rect 2870 1104 2876 1105
rect 2870 1100 2871 1104
rect 2875 1100 2876 1104
rect 2870 1099 2876 1100
rect 3086 1104 3092 1105
rect 3086 1100 3087 1104
rect 3091 1100 3092 1104
rect 3086 1099 3092 1100
rect 3318 1104 3324 1105
rect 3318 1100 3319 1104
rect 3323 1100 3324 1104
rect 3318 1099 3324 1100
rect 3558 1104 3564 1105
rect 3558 1100 3559 1104
rect 3563 1100 3564 1104
rect 3558 1099 3564 1100
rect 3806 1104 3812 1105
rect 3806 1100 3807 1104
rect 3811 1100 3812 1104
rect 3942 1103 3943 1107
rect 3947 1103 3948 1107
rect 3942 1102 3948 1103
rect 3806 1099 3812 1100
rect 110 1096 116 1097
rect 2006 1096 2012 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 134 1095 140 1096
rect 134 1091 135 1095
rect 139 1091 140 1095
rect 134 1090 140 1091
rect 238 1095 244 1096
rect 238 1091 239 1095
rect 243 1091 244 1095
rect 238 1090 244 1091
rect 374 1095 380 1096
rect 374 1091 375 1095
rect 379 1091 380 1095
rect 374 1090 380 1091
rect 526 1095 532 1096
rect 526 1091 527 1095
rect 531 1091 532 1095
rect 526 1090 532 1091
rect 694 1095 700 1096
rect 694 1091 695 1095
rect 699 1091 700 1095
rect 694 1090 700 1091
rect 862 1095 868 1096
rect 862 1091 863 1095
rect 867 1091 868 1095
rect 862 1090 868 1091
rect 1038 1095 1044 1096
rect 1038 1091 1039 1095
rect 1043 1091 1044 1095
rect 1038 1090 1044 1091
rect 1214 1095 1220 1096
rect 1214 1091 1215 1095
rect 1219 1091 1220 1095
rect 1214 1090 1220 1091
rect 1390 1095 1396 1096
rect 1390 1091 1391 1095
rect 1395 1091 1396 1095
rect 1390 1090 1396 1091
rect 1566 1095 1572 1096
rect 1566 1091 1567 1095
rect 1571 1091 1572 1095
rect 1566 1090 1572 1091
rect 1742 1095 1748 1096
rect 1742 1091 1743 1095
rect 1747 1091 1748 1095
rect 1742 1090 1748 1091
rect 1902 1095 1908 1096
rect 1902 1091 1903 1095
rect 1907 1091 1908 1095
rect 2006 1092 2007 1096
rect 2011 1092 2012 1096
rect 2006 1091 2012 1092
rect 1902 1090 1908 1091
rect 210 1087 216 1088
rect 210 1083 211 1087
rect 215 1083 216 1087
rect 210 1082 216 1083
rect 314 1087 320 1088
rect 314 1083 315 1087
rect 319 1083 320 1087
rect 314 1082 320 1083
rect 450 1087 456 1088
rect 450 1083 451 1087
rect 455 1083 456 1087
rect 450 1082 456 1083
rect 602 1087 608 1088
rect 602 1083 603 1087
rect 607 1083 608 1087
rect 602 1082 608 1083
rect 618 1087 624 1088
rect 618 1083 619 1087
rect 623 1086 624 1087
rect 946 1087 952 1088
rect 623 1084 737 1086
rect 623 1083 624 1084
rect 618 1082 624 1083
rect 938 1083 944 1084
rect 110 1079 116 1080
rect 110 1075 111 1079
rect 115 1075 116 1079
rect 938 1079 939 1083
rect 943 1079 944 1083
rect 946 1083 947 1087
rect 951 1086 952 1087
rect 1135 1087 1141 1088
rect 951 1084 1081 1086
rect 951 1083 952 1084
rect 946 1082 952 1083
rect 1135 1083 1136 1087
rect 1140 1086 1141 1087
rect 1466 1087 1472 1088
rect 1140 1084 1257 1086
rect 1140 1083 1141 1084
rect 1135 1082 1141 1083
rect 1466 1083 1467 1087
rect 1471 1083 1472 1087
rect 1466 1082 1472 1083
rect 1503 1087 1509 1088
rect 1503 1083 1504 1087
rect 1508 1086 1509 1087
rect 1818 1087 1824 1088
rect 1508 1084 1609 1086
rect 1508 1083 1509 1084
rect 1503 1082 1509 1083
rect 1818 1083 1819 1087
rect 1823 1083 1824 1087
rect 2134 1087 2140 1088
rect 2134 1086 2135 1087
rect 1981 1084 2135 1086
rect 1818 1082 1824 1083
rect 2134 1083 2135 1084
rect 2139 1083 2140 1087
rect 2134 1082 2140 1083
rect 938 1078 944 1079
rect 2006 1079 2012 1080
rect 110 1074 116 1075
rect 134 1076 140 1077
rect 134 1072 135 1076
rect 139 1072 140 1076
rect 134 1071 140 1072
rect 238 1076 244 1077
rect 238 1072 239 1076
rect 243 1072 244 1076
rect 238 1071 244 1072
rect 374 1076 380 1077
rect 374 1072 375 1076
rect 379 1072 380 1076
rect 374 1071 380 1072
rect 526 1076 532 1077
rect 526 1072 527 1076
rect 531 1072 532 1076
rect 526 1071 532 1072
rect 694 1076 700 1077
rect 694 1072 695 1076
rect 699 1072 700 1076
rect 694 1071 700 1072
rect 862 1076 868 1077
rect 862 1072 863 1076
rect 867 1072 868 1076
rect 862 1071 868 1072
rect 1038 1076 1044 1077
rect 1038 1072 1039 1076
rect 1043 1072 1044 1076
rect 1038 1071 1044 1072
rect 1214 1076 1220 1077
rect 1214 1072 1215 1076
rect 1219 1072 1220 1076
rect 1214 1071 1220 1072
rect 1390 1076 1396 1077
rect 1390 1072 1391 1076
rect 1395 1072 1396 1076
rect 1390 1071 1396 1072
rect 1566 1076 1572 1077
rect 1566 1072 1567 1076
rect 1571 1072 1572 1076
rect 1566 1071 1572 1072
rect 1742 1076 1748 1077
rect 1742 1072 1743 1076
rect 1747 1072 1748 1076
rect 1742 1071 1748 1072
rect 1902 1076 1908 1077
rect 1902 1072 1903 1076
rect 1907 1072 1908 1076
rect 2006 1075 2007 1079
rect 2011 1075 2012 1079
rect 2006 1074 2012 1075
rect 1902 1071 1908 1072
rect 2070 1032 2076 1033
rect 2046 1029 2052 1030
rect 2046 1025 2047 1029
rect 2051 1025 2052 1029
rect 2070 1028 2071 1032
rect 2075 1028 2076 1032
rect 2070 1027 2076 1028
rect 2262 1032 2268 1033
rect 2262 1028 2263 1032
rect 2267 1028 2268 1032
rect 2262 1027 2268 1028
rect 2486 1032 2492 1033
rect 2486 1028 2487 1032
rect 2491 1028 2492 1032
rect 2486 1027 2492 1028
rect 2702 1032 2708 1033
rect 2702 1028 2703 1032
rect 2707 1028 2708 1032
rect 2702 1027 2708 1028
rect 2918 1032 2924 1033
rect 2918 1028 2919 1032
rect 2923 1028 2924 1032
rect 2918 1027 2924 1028
rect 3118 1032 3124 1033
rect 3118 1028 3119 1032
rect 3123 1028 3124 1032
rect 3118 1027 3124 1028
rect 3310 1032 3316 1033
rect 3310 1028 3311 1032
rect 3315 1028 3316 1032
rect 3310 1027 3316 1028
rect 3494 1032 3500 1033
rect 3494 1028 3495 1032
rect 3499 1028 3500 1032
rect 3494 1027 3500 1028
rect 3678 1032 3684 1033
rect 3678 1028 3679 1032
rect 3683 1028 3684 1032
rect 3678 1027 3684 1028
rect 3838 1032 3844 1033
rect 3838 1028 3839 1032
rect 3843 1028 3844 1032
rect 3838 1027 3844 1028
rect 3942 1029 3948 1030
rect 2046 1024 2052 1025
rect 3942 1025 3943 1029
rect 3947 1025 3948 1029
rect 3942 1024 3948 1025
rect 202 1023 208 1024
rect 202 1019 203 1023
rect 207 1022 208 1023
rect 2146 1023 2152 1024
rect 207 1020 558 1022
rect 207 1019 208 1020
rect 202 1018 208 1019
rect 134 1016 140 1017
rect 110 1013 116 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 134 1012 135 1016
rect 139 1012 140 1016
rect 134 1011 140 1012
rect 286 1016 292 1017
rect 286 1012 287 1016
rect 291 1012 292 1016
rect 286 1011 292 1012
rect 470 1016 476 1017
rect 470 1012 471 1016
rect 475 1012 476 1016
rect 470 1011 476 1012
rect 110 1008 116 1009
rect 222 1007 228 1008
rect 222 1006 223 1007
rect 213 1004 223 1006
rect 222 1003 223 1004
rect 227 1003 228 1007
rect 222 1002 228 1003
rect 362 1007 368 1008
rect 362 1003 363 1007
rect 367 1003 368 1007
rect 362 1002 368 1003
rect 546 1007 552 1008
rect 546 1003 547 1007
rect 551 1003 552 1007
rect 556 1006 558 1020
rect 2146 1019 2147 1023
rect 2151 1019 2152 1023
rect 2146 1018 2152 1019
rect 2338 1023 2344 1024
rect 2338 1019 2339 1023
rect 2343 1019 2344 1023
rect 2338 1018 2344 1019
rect 2562 1023 2568 1024
rect 2562 1019 2563 1023
rect 2567 1019 2568 1023
rect 2562 1018 2568 1019
rect 2570 1023 2576 1024
rect 2570 1019 2571 1023
rect 2575 1022 2576 1023
rect 3002 1023 3008 1024
rect 2575 1020 2745 1022
rect 2575 1019 2576 1020
rect 2570 1018 2576 1019
rect 654 1016 660 1017
rect 654 1012 655 1016
rect 659 1012 660 1016
rect 654 1011 660 1012
rect 838 1016 844 1017
rect 838 1012 839 1016
rect 843 1012 844 1016
rect 838 1011 844 1012
rect 1014 1016 1020 1017
rect 1014 1012 1015 1016
rect 1019 1012 1020 1016
rect 1014 1011 1020 1012
rect 1198 1016 1204 1017
rect 1198 1012 1199 1016
rect 1203 1012 1204 1016
rect 1198 1011 1204 1012
rect 1382 1016 1388 1017
rect 1382 1012 1383 1016
rect 1387 1012 1388 1016
rect 1382 1011 1388 1012
rect 1566 1016 1572 1017
rect 1566 1012 1567 1016
rect 1571 1012 1572 1016
rect 2996 1014 2998 1021
rect 3002 1019 3003 1023
rect 3007 1022 3008 1023
rect 3202 1023 3208 1024
rect 3007 1020 3161 1022
rect 3007 1019 3008 1020
rect 3002 1018 3008 1019
rect 3202 1019 3203 1023
rect 3207 1022 3208 1023
rect 3570 1023 3576 1024
rect 3207 1020 3353 1022
rect 3207 1019 3208 1020
rect 3202 1018 3208 1019
rect 3570 1019 3571 1023
rect 3575 1019 3576 1023
rect 3570 1018 3576 1019
rect 3754 1023 3760 1024
rect 3754 1019 3755 1023
rect 3759 1019 3760 1023
rect 3754 1018 3760 1019
rect 3906 1023 3912 1024
rect 3906 1019 3907 1023
rect 3911 1019 3912 1023
rect 3906 1018 3912 1019
rect 3038 1015 3044 1016
rect 3038 1014 3039 1015
rect 1566 1011 1572 1012
rect 2006 1013 2012 1014
rect 2070 1013 2076 1014
rect 2006 1009 2007 1013
rect 2011 1009 2012 1013
rect 2006 1008 2012 1009
rect 2046 1012 2052 1013
rect 2046 1008 2047 1012
rect 2051 1008 2052 1012
rect 2070 1009 2071 1013
rect 2075 1009 2076 1013
rect 2070 1008 2076 1009
rect 2262 1013 2268 1014
rect 2262 1009 2263 1013
rect 2267 1009 2268 1013
rect 2262 1008 2268 1009
rect 2486 1013 2492 1014
rect 2486 1009 2487 1013
rect 2491 1009 2492 1013
rect 2486 1008 2492 1009
rect 2702 1013 2708 1014
rect 2702 1009 2703 1013
rect 2707 1009 2708 1013
rect 2702 1008 2708 1009
rect 2918 1013 2924 1014
rect 2918 1009 2919 1013
rect 2923 1009 2924 1013
rect 2996 1012 3039 1014
rect 3038 1011 3039 1012
rect 3043 1011 3044 1015
rect 3038 1010 3044 1011
rect 3118 1013 3124 1014
rect 2918 1008 2924 1009
rect 3118 1009 3119 1013
rect 3123 1009 3124 1013
rect 3118 1008 3124 1009
rect 3310 1013 3316 1014
rect 3310 1009 3311 1013
rect 3315 1009 3316 1013
rect 3310 1008 3316 1009
rect 3494 1013 3500 1014
rect 3494 1009 3495 1013
rect 3499 1009 3500 1013
rect 3494 1008 3500 1009
rect 3678 1013 3684 1014
rect 3678 1009 3679 1013
rect 3683 1009 3684 1013
rect 3678 1008 3684 1009
rect 3838 1013 3844 1014
rect 3838 1009 3839 1013
rect 3843 1009 3844 1013
rect 3838 1008 3844 1009
rect 3942 1012 3948 1013
rect 3942 1008 3943 1012
rect 3947 1008 3948 1012
rect 978 1007 984 1008
rect 978 1006 979 1007
rect 556 1004 697 1006
rect 917 1004 979 1006
rect 546 1002 552 1003
rect 978 1003 979 1004
rect 983 1003 984 1007
rect 978 1002 984 1003
rect 1006 1007 1012 1008
rect 1006 1003 1007 1007
rect 1011 1006 1012 1007
rect 1274 1007 1280 1008
rect 1011 1004 1057 1006
rect 1011 1003 1012 1004
rect 1006 1002 1012 1003
rect 1274 1003 1275 1007
rect 1279 1003 1280 1007
rect 1274 1002 1280 1003
rect 1454 1007 1460 1008
rect 1454 1003 1455 1007
rect 1459 1003 1460 1007
rect 1454 1002 1460 1003
rect 1466 1007 1472 1008
rect 2046 1007 2052 1008
rect 3942 1007 3948 1008
rect 1466 1003 1467 1007
rect 1471 1006 1472 1007
rect 1471 1004 1609 1006
rect 1471 1003 1472 1004
rect 1466 1002 1472 1003
rect 134 997 140 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 134 993 135 997
rect 139 993 140 997
rect 134 992 140 993
rect 286 997 292 998
rect 286 993 287 997
rect 291 993 292 997
rect 286 992 292 993
rect 470 997 476 998
rect 470 993 471 997
rect 475 993 476 997
rect 470 992 476 993
rect 654 997 660 998
rect 654 993 655 997
rect 659 993 660 997
rect 654 992 660 993
rect 838 997 844 998
rect 838 993 839 997
rect 843 993 844 997
rect 838 992 844 993
rect 1014 997 1020 998
rect 1014 993 1015 997
rect 1019 993 1020 997
rect 1014 992 1020 993
rect 1198 997 1204 998
rect 1198 993 1199 997
rect 1203 993 1204 997
rect 1198 992 1204 993
rect 1382 997 1388 998
rect 1382 993 1383 997
rect 1387 993 1388 997
rect 1382 992 1388 993
rect 1566 997 1572 998
rect 1566 993 1567 997
rect 1571 993 1572 997
rect 1566 992 1572 993
rect 2006 996 2012 997
rect 2006 992 2007 996
rect 2011 992 2012 996
rect 110 991 116 992
rect 2006 991 2012 992
rect 2134 991 2141 992
rect 2134 987 2135 991
rect 2140 987 2141 991
rect 2134 986 2141 987
rect 2146 991 2152 992
rect 2146 987 2147 991
rect 2151 990 2152 991
rect 2327 991 2333 992
rect 2327 990 2328 991
rect 2151 988 2328 990
rect 2151 987 2152 988
rect 2146 986 2152 987
rect 2327 987 2328 988
rect 2332 987 2333 991
rect 2327 986 2333 987
rect 2338 991 2344 992
rect 2338 987 2339 991
rect 2343 990 2344 991
rect 2551 991 2557 992
rect 2551 990 2552 991
rect 2343 988 2552 990
rect 2343 987 2344 988
rect 2338 986 2344 987
rect 2551 987 2552 988
rect 2556 987 2557 991
rect 2551 986 2557 987
rect 2562 991 2568 992
rect 2562 987 2563 991
rect 2567 990 2568 991
rect 2767 991 2773 992
rect 2767 990 2768 991
rect 2567 988 2768 990
rect 2567 987 2568 988
rect 2562 986 2568 987
rect 2767 987 2768 988
rect 2772 987 2773 991
rect 2767 986 2773 987
rect 2983 991 2989 992
rect 2983 987 2984 991
rect 2988 990 2989 991
rect 3002 991 3008 992
rect 3002 990 3003 991
rect 2988 988 3003 990
rect 2988 987 2989 988
rect 2983 986 2989 987
rect 3002 987 3003 988
rect 3007 987 3008 991
rect 3002 986 3008 987
rect 3183 991 3189 992
rect 3183 987 3184 991
rect 3188 990 3189 991
rect 3202 991 3208 992
rect 3202 990 3203 991
rect 3188 988 3203 990
rect 3188 987 3189 988
rect 3183 986 3189 987
rect 3202 987 3203 988
rect 3207 987 3208 991
rect 3202 986 3208 987
rect 3375 991 3381 992
rect 3375 987 3376 991
rect 3380 990 3381 991
rect 3402 991 3408 992
rect 3402 990 3403 991
rect 3380 988 3403 990
rect 3380 987 3381 988
rect 3375 986 3381 987
rect 3402 987 3403 988
rect 3407 987 3408 991
rect 3402 986 3408 987
rect 3550 991 3556 992
rect 3550 987 3551 991
rect 3555 990 3556 991
rect 3559 991 3565 992
rect 3559 990 3560 991
rect 3555 988 3560 990
rect 3555 987 3556 988
rect 3550 986 3556 987
rect 3559 987 3560 988
rect 3564 987 3565 991
rect 3559 986 3565 987
rect 3570 991 3576 992
rect 3570 987 3571 991
rect 3575 990 3576 991
rect 3743 991 3749 992
rect 3743 990 3744 991
rect 3575 988 3744 990
rect 3575 987 3576 988
rect 3570 986 3576 987
rect 3743 987 3744 988
rect 3748 987 3749 991
rect 3743 986 3749 987
rect 3882 991 3888 992
rect 3882 987 3883 991
rect 3887 990 3888 991
rect 3903 991 3909 992
rect 3903 990 3904 991
rect 3887 988 3904 990
rect 3887 987 3888 988
rect 3882 986 3888 987
rect 3903 987 3904 988
rect 3908 987 3909 991
rect 3903 986 3909 987
rect 1466 983 1472 984
rect 1466 982 1467 983
rect 1268 980 1467 982
rect 1268 976 1270 980
rect 1466 979 1467 980
rect 1471 979 1472 983
rect 2570 983 2576 984
rect 2570 982 2571 983
rect 1466 978 1472 979
rect 2369 980 2571 982
rect 2369 976 2371 980
rect 2570 979 2571 980
rect 2575 979 2576 983
rect 2570 978 2576 979
rect 199 975 205 976
rect 199 971 200 975
rect 204 974 205 975
rect 210 975 216 976
rect 210 974 211 975
rect 204 972 211 974
rect 204 971 205 972
rect 199 970 205 971
rect 210 971 211 972
rect 215 971 216 975
rect 210 970 216 971
rect 222 975 228 976
rect 222 971 223 975
rect 227 974 228 975
rect 351 975 357 976
rect 351 974 352 975
rect 227 972 352 974
rect 227 971 228 972
rect 222 970 228 971
rect 351 971 352 972
rect 356 971 357 975
rect 351 970 357 971
rect 362 975 368 976
rect 362 971 363 975
rect 367 974 368 975
rect 535 975 541 976
rect 535 974 536 975
rect 367 972 536 974
rect 367 971 368 972
rect 362 970 368 971
rect 535 971 536 972
rect 540 971 541 975
rect 535 970 541 971
rect 546 975 552 976
rect 546 971 547 975
rect 551 974 552 975
rect 719 975 725 976
rect 719 974 720 975
rect 551 972 720 974
rect 551 971 552 972
rect 546 970 552 971
rect 719 971 720 972
rect 724 971 725 975
rect 719 970 725 971
rect 903 975 909 976
rect 903 971 904 975
rect 908 974 909 975
rect 938 975 944 976
rect 938 974 939 975
rect 908 972 939 974
rect 908 971 909 972
rect 903 970 909 971
rect 938 971 939 972
rect 943 971 944 975
rect 938 970 944 971
rect 978 975 984 976
rect 978 971 979 975
rect 983 974 984 975
rect 1079 975 1085 976
rect 1079 974 1080 975
rect 983 972 1080 974
rect 983 971 984 972
rect 978 970 984 971
rect 1079 971 1080 972
rect 1084 971 1085 975
rect 1079 970 1085 971
rect 1263 975 1270 976
rect 1263 971 1264 975
rect 1268 972 1270 975
rect 1274 975 1280 976
rect 1268 971 1269 972
rect 1263 970 1269 971
rect 1274 971 1275 975
rect 1279 974 1280 975
rect 1447 975 1453 976
rect 1447 974 1448 975
rect 1279 972 1448 974
rect 1279 971 1280 972
rect 1274 970 1280 971
rect 1447 971 1448 972
rect 1452 971 1453 975
rect 1447 970 1453 971
rect 1582 975 1588 976
rect 1582 971 1583 975
rect 1587 974 1588 975
rect 1631 975 1637 976
rect 1631 974 1632 975
rect 1587 972 1632 974
rect 1587 971 1588 972
rect 1582 970 1588 971
rect 1631 971 1632 972
rect 1636 971 1637 975
rect 1631 970 1637 971
rect 2367 975 2373 976
rect 2367 971 2368 975
rect 2372 971 2373 975
rect 2367 970 2373 971
rect 2378 975 2384 976
rect 2378 971 2379 975
rect 2383 974 2384 975
rect 2519 975 2525 976
rect 2519 974 2520 975
rect 2383 972 2520 974
rect 2383 971 2384 972
rect 2378 970 2384 971
rect 2519 971 2520 972
rect 2524 971 2525 975
rect 2519 970 2525 971
rect 2530 975 2536 976
rect 2530 971 2531 975
rect 2535 974 2536 975
rect 2679 975 2685 976
rect 2679 974 2680 975
rect 2535 972 2680 974
rect 2535 971 2536 972
rect 2530 970 2536 971
rect 2679 971 2680 972
rect 2684 971 2685 975
rect 2679 970 2685 971
rect 2690 975 2696 976
rect 2690 971 2691 975
rect 2695 974 2696 975
rect 2847 975 2853 976
rect 2847 974 2848 975
rect 2695 972 2848 974
rect 2695 971 2696 972
rect 2690 970 2696 971
rect 2847 971 2848 972
rect 2852 971 2853 975
rect 2847 970 2853 971
rect 2858 975 2864 976
rect 2858 971 2859 975
rect 2863 974 2864 975
rect 3015 975 3021 976
rect 3015 974 3016 975
rect 2863 972 3016 974
rect 2863 971 2864 972
rect 2858 970 2864 971
rect 3015 971 3016 972
rect 3020 971 3021 975
rect 3015 970 3021 971
rect 3038 975 3044 976
rect 3038 971 3039 975
rect 3043 974 3044 975
rect 3175 975 3181 976
rect 3175 974 3176 975
rect 3043 972 3176 974
rect 3043 971 3044 972
rect 3038 970 3044 971
rect 3175 971 3176 972
rect 3180 971 3181 975
rect 3175 970 3181 971
rect 3186 975 3192 976
rect 3186 971 3187 975
rect 3191 974 3192 975
rect 3327 975 3333 976
rect 3327 974 3328 975
rect 3191 972 3328 974
rect 3191 971 3192 972
rect 3186 970 3192 971
rect 3327 971 3328 972
rect 3332 971 3333 975
rect 3327 970 3333 971
rect 3338 975 3344 976
rect 3338 971 3339 975
rect 3343 974 3344 975
rect 3479 975 3485 976
rect 3479 974 3480 975
rect 3343 972 3480 974
rect 3343 971 3344 972
rect 3338 970 3344 971
rect 3479 971 3480 972
rect 3484 971 3485 975
rect 3479 970 3485 971
rect 3538 975 3544 976
rect 3538 971 3539 975
rect 3543 974 3544 975
rect 3623 975 3629 976
rect 3623 974 3624 975
rect 3543 972 3624 974
rect 3543 971 3544 972
rect 3538 970 3544 971
rect 3623 971 3624 972
rect 3628 971 3629 975
rect 3623 970 3629 971
rect 3775 975 3781 976
rect 3775 971 3776 975
rect 3780 974 3781 975
rect 3794 975 3800 976
rect 3794 974 3795 975
rect 3780 972 3795 974
rect 3780 971 3781 972
rect 3775 970 3781 971
rect 3794 971 3795 972
rect 3799 971 3800 975
rect 3794 970 3800 971
rect 3903 975 3912 976
rect 3903 971 3904 975
rect 3911 971 3912 975
rect 3903 970 3912 971
rect 199 959 205 960
rect 199 955 200 959
rect 204 958 205 959
rect 270 959 276 960
rect 270 958 271 959
rect 204 956 271 958
rect 204 955 205 956
rect 199 954 205 955
rect 270 955 271 956
rect 275 955 276 959
rect 270 954 276 955
rect 359 959 365 960
rect 359 955 360 959
rect 364 958 365 959
rect 399 959 405 960
rect 399 958 400 959
rect 364 956 400 958
rect 364 955 365 956
rect 359 954 365 955
rect 399 955 400 956
rect 404 955 405 959
rect 399 954 405 955
rect 430 959 436 960
rect 430 955 431 959
rect 435 958 436 959
rect 535 959 541 960
rect 535 958 536 959
rect 435 956 536 958
rect 435 955 436 956
rect 430 954 436 955
rect 535 955 536 956
rect 540 955 541 959
rect 535 954 541 955
rect 703 959 709 960
rect 703 955 704 959
rect 708 958 709 959
rect 727 959 733 960
rect 727 958 728 959
rect 708 956 728 958
rect 708 955 709 956
rect 703 954 709 955
rect 727 955 728 956
rect 732 955 733 959
rect 727 954 733 955
rect 863 959 869 960
rect 863 955 864 959
rect 868 958 869 959
rect 882 959 888 960
rect 882 958 883 959
rect 868 956 883 958
rect 868 955 869 956
rect 863 954 869 955
rect 882 955 883 956
rect 887 955 888 959
rect 882 954 888 955
rect 1006 959 1012 960
rect 1006 955 1007 959
rect 1011 958 1012 959
rect 1015 959 1021 960
rect 1015 958 1016 959
rect 1011 956 1016 958
rect 1011 955 1012 956
rect 1006 954 1012 955
rect 1015 955 1016 956
rect 1020 955 1021 959
rect 1015 954 1021 955
rect 1151 959 1157 960
rect 1151 955 1152 959
rect 1156 958 1157 959
rect 1162 959 1168 960
rect 1156 955 1158 958
rect 1151 954 1158 955
rect 1162 955 1163 959
rect 1167 958 1168 959
rect 1287 959 1293 960
rect 1287 958 1288 959
rect 1167 956 1288 958
rect 1167 955 1168 956
rect 1162 954 1168 955
rect 1287 955 1288 956
rect 1292 955 1293 959
rect 1287 954 1293 955
rect 1298 959 1304 960
rect 1298 955 1299 959
rect 1303 958 1304 959
rect 1423 959 1429 960
rect 1423 958 1424 959
rect 1303 956 1424 958
rect 1303 955 1304 956
rect 1298 954 1304 955
rect 1423 955 1424 956
rect 1428 955 1429 959
rect 1423 954 1429 955
rect 1434 959 1440 960
rect 1434 955 1435 959
rect 1439 958 1440 959
rect 1559 959 1565 960
rect 1559 958 1560 959
rect 1439 956 1560 958
rect 1439 955 1440 956
rect 1434 954 1440 955
rect 1559 955 1560 956
rect 1564 955 1565 959
rect 1559 954 1565 955
rect 2046 956 2052 957
rect 3942 956 3948 957
rect 1156 950 1158 954
rect 2046 952 2047 956
rect 2051 952 2052 956
rect 1314 951 1320 952
rect 2046 951 2052 952
rect 2302 955 2308 956
rect 2302 951 2303 955
rect 2307 951 2308 955
rect 1314 950 1315 951
rect 1156 948 1315 950
rect 1314 947 1315 948
rect 1319 947 1320 951
rect 2302 950 2308 951
rect 2454 955 2460 956
rect 2454 951 2455 955
rect 2459 951 2460 955
rect 2454 950 2460 951
rect 2614 955 2620 956
rect 2614 951 2615 955
rect 2619 951 2620 955
rect 2614 950 2620 951
rect 2782 955 2788 956
rect 2782 951 2783 955
rect 2787 951 2788 955
rect 2782 950 2788 951
rect 2950 955 2956 956
rect 2950 951 2951 955
rect 2955 951 2956 955
rect 2950 950 2956 951
rect 3110 955 3116 956
rect 3110 951 3111 955
rect 3115 951 3116 955
rect 3110 950 3116 951
rect 3262 955 3268 956
rect 3262 951 3263 955
rect 3267 951 3268 955
rect 3262 950 3268 951
rect 3414 955 3420 956
rect 3414 951 3415 955
rect 3419 951 3420 955
rect 3414 950 3420 951
rect 3558 955 3564 956
rect 3558 951 3559 955
rect 3563 951 3564 955
rect 3558 950 3564 951
rect 3710 955 3716 956
rect 3710 951 3711 955
rect 3715 951 3716 955
rect 3710 950 3716 951
rect 3838 955 3844 956
rect 3838 951 3839 955
rect 3843 951 3844 955
rect 3942 952 3943 956
rect 3947 952 3948 956
rect 3942 951 3948 952
rect 3838 950 3844 951
rect 1314 946 1320 947
rect 2378 947 2384 948
rect 2378 943 2379 947
rect 2383 943 2384 947
rect 2378 942 2384 943
rect 2530 947 2536 948
rect 2530 943 2531 947
rect 2535 943 2536 947
rect 2530 942 2536 943
rect 2690 947 2696 948
rect 2690 943 2691 947
rect 2695 943 2696 947
rect 2690 942 2696 943
rect 2858 947 2864 948
rect 2858 943 2859 947
rect 2863 943 2864 947
rect 2858 942 2864 943
rect 2906 947 2912 948
rect 2906 943 2907 947
rect 2911 946 2912 947
rect 3186 947 3192 948
rect 2911 944 2993 946
rect 2911 943 2912 944
rect 2906 942 2912 943
rect 3186 943 3187 947
rect 3191 943 3192 947
rect 3186 942 3192 943
rect 3338 947 3344 948
rect 3338 943 3339 947
rect 3343 943 3344 947
rect 3538 947 3544 948
rect 3538 946 3539 947
rect 3493 944 3539 946
rect 3338 942 3344 943
rect 3538 943 3539 944
rect 3543 943 3544 947
rect 3538 942 3544 943
rect 3550 947 3556 948
rect 3550 943 3551 947
rect 3555 946 3556 947
rect 3642 947 3648 948
rect 3555 944 3601 946
rect 3555 943 3556 944
rect 3550 942 3556 943
rect 3642 943 3643 947
rect 3647 946 3648 947
rect 3647 944 3753 946
rect 3647 943 3648 944
rect 3642 942 3648 943
rect 3914 943 3920 944
rect 110 940 116 941
rect 2006 940 2012 941
rect 110 936 111 940
rect 115 936 116 940
rect 110 935 116 936
rect 134 939 140 940
rect 134 935 135 939
rect 139 935 140 939
rect 134 934 140 935
rect 294 939 300 940
rect 294 935 295 939
rect 299 935 300 939
rect 294 934 300 935
rect 470 939 476 940
rect 470 935 471 939
rect 475 935 476 939
rect 470 934 476 935
rect 638 939 644 940
rect 638 935 639 939
rect 643 935 644 939
rect 638 934 644 935
rect 798 939 804 940
rect 798 935 799 939
rect 803 935 804 939
rect 798 934 804 935
rect 950 939 956 940
rect 950 935 951 939
rect 955 935 956 939
rect 950 934 956 935
rect 1086 939 1092 940
rect 1086 935 1087 939
rect 1091 935 1092 939
rect 1086 934 1092 935
rect 1222 939 1228 940
rect 1222 935 1223 939
rect 1227 935 1228 939
rect 1222 934 1228 935
rect 1358 939 1364 940
rect 1358 935 1359 939
rect 1363 935 1364 939
rect 1358 934 1364 935
rect 1494 939 1500 940
rect 1494 935 1495 939
rect 1499 935 1500 939
rect 2006 936 2007 940
rect 2011 936 2012 940
rect 2006 935 2012 936
rect 2046 939 2052 940
rect 2046 935 2047 939
rect 2051 935 2052 939
rect 3914 939 3915 943
rect 3919 939 3920 943
rect 3914 938 3920 939
rect 3942 939 3948 940
rect 1494 934 1500 935
rect 2046 934 2052 935
rect 2302 936 2308 937
rect 2302 932 2303 936
rect 2307 932 2308 936
rect 210 931 216 932
rect 210 927 211 931
rect 215 927 216 931
rect 210 926 216 927
rect 270 931 276 932
rect 270 927 271 931
rect 275 930 276 931
rect 399 931 405 932
rect 275 928 337 930
rect 275 927 276 928
rect 270 926 276 927
rect 399 927 400 931
rect 404 930 405 931
rect 727 931 733 932
rect 404 928 513 930
rect 404 927 405 928
rect 399 926 405 927
rect 714 927 720 928
rect 110 923 116 924
rect 110 919 111 923
rect 115 919 116 923
rect 714 923 715 927
rect 719 923 720 927
rect 727 927 728 931
rect 732 930 733 931
rect 882 931 888 932
rect 732 928 841 930
rect 732 927 733 928
rect 727 926 733 927
rect 882 927 883 931
rect 887 930 888 931
rect 1162 931 1168 932
rect 887 928 993 930
rect 887 927 888 928
rect 882 926 888 927
rect 1162 927 1163 931
rect 1167 927 1168 931
rect 1162 926 1168 927
rect 1298 931 1304 932
rect 1298 927 1299 931
rect 1303 927 1304 931
rect 1298 926 1304 927
rect 1434 931 1440 932
rect 1434 927 1435 931
rect 1439 927 1440 931
rect 1582 931 1588 932
rect 2302 931 2308 932
rect 2454 936 2460 937
rect 2454 932 2455 936
rect 2459 932 2460 936
rect 2454 931 2460 932
rect 2614 936 2620 937
rect 2614 932 2615 936
rect 2619 932 2620 936
rect 2614 931 2620 932
rect 2782 936 2788 937
rect 2782 932 2783 936
rect 2787 932 2788 936
rect 2782 931 2788 932
rect 2950 936 2956 937
rect 2950 932 2951 936
rect 2955 932 2956 936
rect 2950 931 2956 932
rect 3110 936 3116 937
rect 3110 932 3111 936
rect 3115 932 3116 936
rect 3110 931 3116 932
rect 3262 936 3268 937
rect 3262 932 3263 936
rect 3267 932 3268 936
rect 3262 931 3268 932
rect 3414 936 3420 937
rect 3414 932 3415 936
rect 3419 932 3420 936
rect 3414 931 3420 932
rect 3558 936 3564 937
rect 3558 932 3559 936
rect 3563 932 3564 936
rect 3558 931 3564 932
rect 3710 936 3716 937
rect 3710 932 3711 936
rect 3715 932 3716 936
rect 3710 931 3716 932
rect 3838 936 3844 937
rect 3838 932 3839 936
rect 3843 932 3844 936
rect 3942 935 3943 939
rect 3947 935 3948 939
rect 3942 934 3948 935
rect 3838 931 3844 932
rect 1582 930 1583 931
rect 1573 928 1583 930
rect 1434 926 1440 927
rect 1582 927 1583 928
rect 1587 927 1588 931
rect 1582 926 1588 927
rect 714 922 720 923
rect 2006 923 2012 924
rect 110 918 116 919
rect 134 920 140 921
rect 134 916 135 920
rect 139 916 140 920
rect 134 915 140 916
rect 294 920 300 921
rect 294 916 295 920
rect 299 916 300 920
rect 294 915 300 916
rect 470 920 476 921
rect 470 916 471 920
rect 475 916 476 920
rect 470 915 476 916
rect 638 920 644 921
rect 638 916 639 920
rect 643 916 644 920
rect 638 915 644 916
rect 798 920 804 921
rect 798 916 799 920
rect 803 916 804 920
rect 798 915 804 916
rect 950 920 956 921
rect 950 916 951 920
rect 955 916 956 920
rect 950 915 956 916
rect 1086 920 1092 921
rect 1086 916 1087 920
rect 1091 916 1092 920
rect 1086 915 1092 916
rect 1222 920 1228 921
rect 1222 916 1223 920
rect 1227 916 1228 920
rect 1222 915 1228 916
rect 1358 920 1364 921
rect 1358 916 1359 920
rect 1363 916 1364 920
rect 1358 915 1364 916
rect 1494 920 1500 921
rect 1494 916 1495 920
rect 1499 916 1500 920
rect 2006 919 2007 923
rect 2011 919 2012 923
rect 2006 918 2012 919
rect 1494 915 1500 916
rect 2558 872 2564 873
rect 2046 869 2052 870
rect 2046 865 2047 869
rect 2051 865 2052 869
rect 2558 868 2559 872
rect 2563 868 2564 872
rect 2558 867 2564 868
rect 2678 872 2684 873
rect 2678 868 2679 872
rect 2683 868 2684 872
rect 2678 867 2684 868
rect 2806 872 2812 873
rect 2806 868 2807 872
rect 2811 868 2812 872
rect 2806 867 2812 868
rect 2942 872 2948 873
rect 2942 868 2943 872
rect 2947 868 2948 872
rect 2942 867 2948 868
rect 3078 872 3084 873
rect 3078 868 3079 872
rect 3083 868 3084 872
rect 3078 867 3084 868
rect 3206 872 3212 873
rect 3206 868 3207 872
rect 3211 868 3212 872
rect 3206 867 3212 868
rect 3334 872 3340 873
rect 3334 868 3335 872
rect 3339 868 3340 872
rect 3334 867 3340 868
rect 3462 872 3468 873
rect 3462 868 3463 872
rect 3467 868 3468 872
rect 3462 867 3468 868
rect 3590 872 3596 873
rect 3590 868 3591 872
rect 3595 868 3596 872
rect 3590 867 3596 868
rect 3726 872 3732 873
rect 3726 868 3727 872
rect 3731 868 3732 872
rect 3726 867 3732 868
rect 3838 872 3844 873
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 3838 867 3844 868
rect 3942 869 3948 870
rect 2046 864 2052 865
rect 3942 865 3943 869
rect 3947 865 3948 869
rect 3942 864 3948 865
rect 2634 863 2640 864
rect 158 860 164 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 158 856 159 860
rect 163 856 164 860
rect 158 855 164 856
rect 318 860 324 861
rect 318 856 319 860
rect 323 856 324 860
rect 318 855 324 856
rect 470 860 476 861
rect 470 856 471 860
rect 475 856 476 860
rect 470 855 476 856
rect 614 860 620 861
rect 614 856 615 860
rect 619 856 620 860
rect 614 855 620 856
rect 750 860 756 861
rect 750 856 751 860
rect 755 856 756 860
rect 750 855 756 856
rect 878 860 884 861
rect 878 856 879 860
rect 883 856 884 860
rect 878 855 884 856
rect 998 860 1004 861
rect 998 856 999 860
rect 1003 856 1004 860
rect 998 855 1004 856
rect 1110 860 1116 861
rect 1110 856 1111 860
rect 1115 856 1116 860
rect 1110 855 1116 856
rect 1230 860 1236 861
rect 1230 856 1231 860
rect 1235 856 1236 860
rect 1230 855 1236 856
rect 1350 860 1356 861
rect 1350 856 1351 860
rect 1355 856 1356 860
rect 2634 859 2635 863
rect 2639 859 2640 863
rect 2634 858 2640 859
rect 2754 863 2760 864
rect 2754 859 2755 863
rect 2759 859 2760 863
rect 2754 858 2760 859
rect 2882 863 2888 864
rect 2882 859 2883 863
rect 2887 859 2888 863
rect 2882 858 2888 859
rect 3018 863 3024 864
rect 3018 859 3019 863
rect 3023 859 3024 863
rect 3018 858 3024 859
rect 3026 863 3032 864
rect 3026 859 3027 863
rect 3031 862 3032 863
rect 3162 863 3168 864
rect 3031 860 3121 862
rect 3031 859 3032 860
rect 3026 858 3032 859
rect 3162 859 3163 863
rect 3167 862 3168 863
rect 3290 863 3296 864
rect 3167 860 3249 862
rect 3167 859 3168 860
rect 3162 858 3168 859
rect 3290 859 3291 863
rect 3295 862 3296 863
rect 3418 863 3424 864
rect 3295 860 3377 862
rect 3295 859 3296 860
rect 3290 858 3296 859
rect 3418 859 3419 863
rect 3423 862 3424 863
rect 3666 863 3672 864
rect 3423 860 3505 862
rect 3423 859 3424 860
rect 3418 858 3424 859
rect 3666 859 3667 863
rect 3671 859 3672 863
rect 3666 858 3672 859
rect 3794 863 3800 864
rect 3794 859 3795 863
rect 3799 859 3800 863
rect 3794 858 3800 859
rect 3906 863 3912 864
rect 3906 859 3907 863
rect 3911 859 3912 863
rect 3906 858 3912 859
rect 1350 855 1356 856
rect 2006 857 2012 858
rect 110 852 116 853
rect 2006 853 2007 857
rect 2011 853 2012 857
rect 2558 853 2564 854
rect 2006 852 2012 853
rect 2046 852 2052 853
rect 234 851 240 852
rect 234 847 235 851
rect 239 847 240 851
rect 430 851 436 852
rect 430 850 431 851
rect 397 848 431 850
rect 234 846 240 847
rect 430 847 431 848
rect 435 847 436 851
rect 430 846 436 847
rect 546 851 552 852
rect 546 847 547 851
rect 551 847 552 851
rect 546 846 552 847
rect 554 851 560 852
rect 554 847 555 851
rect 559 850 560 851
rect 698 851 704 852
rect 559 848 657 850
rect 559 847 560 848
rect 554 846 560 847
rect 698 847 699 851
rect 703 850 704 851
rect 990 851 996 852
rect 990 850 991 851
rect 703 848 793 850
rect 957 848 991 850
rect 703 847 704 848
rect 698 846 704 847
rect 990 847 991 848
rect 995 847 996 851
rect 1098 851 1104 852
rect 1098 850 1099 851
rect 1077 848 1099 850
rect 990 846 996 847
rect 1098 847 1099 848
rect 1103 847 1104 851
rect 1098 846 1104 847
rect 1186 851 1192 852
rect 1186 847 1187 851
rect 1191 847 1192 851
rect 1186 846 1192 847
rect 1306 851 1312 852
rect 1306 847 1307 851
rect 1311 847 1312 851
rect 1306 846 1312 847
rect 1314 851 1320 852
rect 1314 847 1315 851
rect 1319 850 1320 851
rect 1319 848 1393 850
rect 2046 848 2047 852
rect 2051 848 2052 852
rect 2558 849 2559 853
rect 2563 849 2564 853
rect 2558 848 2564 849
rect 2678 853 2684 854
rect 2678 849 2679 853
rect 2683 849 2684 853
rect 2678 848 2684 849
rect 2806 853 2812 854
rect 2806 849 2807 853
rect 2811 849 2812 853
rect 2806 848 2812 849
rect 2942 853 2948 854
rect 2942 849 2943 853
rect 2947 849 2948 853
rect 2942 848 2948 849
rect 3078 853 3084 854
rect 3078 849 3079 853
rect 3083 849 3084 853
rect 3078 848 3084 849
rect 3206 853 3212 854
rect 3206 849 3207 853
rect 3211 849 3212 853
rect 3206 848 3212 849
rect 3334 853 3340 854
rect 3334 849 3335 853
rect 3339 849 3340 853
rect 3334 848 3340 849
rect 3462 853 3468 854
rect 3462 849 3463 853
rect 3467 849 3468 853
rect 3462 848 3468 849
rect 3590 853 3596 854
rect 3590 849 3591 853
rect 3595 849 3596 853
rect 3590 848 3596 849
rect 3726 853 3732 854
rect 3726 849 3727 853
rect 3731 849 3732 853
rect 3726 848 3732 849
rect 3838 853 3844 854
rect 3838 849 3839 853
rect 3843 849 3844 853
rect 3838 848 3844 849
rect 3942 852 3948 853
rect 3942 848 3943 852
rect 3947 848 3948 852
rect 1319 847 1320 848
rect 2046 847 2052 848
rect 3942 847 3948 848
rect 1314 846 1320 847
rect 158 841 164 842
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 158 837 159 841
rect 163 837 164 841
rect 158 836 164 837
rect 318 841 324 842
rect 318 837 319 841
rect 323 837 324 841
rect 318 836 324 837
rect 470 841 476 842
rect 470 837 471 841
rect 475 837 476 841
rect 470 836 476 837
rect 614 841 620 842
rect 614 837 615 841
rect 619 837 620 841
rect 614 836 620 837
rect 750 841 756 842
rect 750 837 751 841
rect 755 837 756 841
rect 750 836 756 837
rect 878 841 884 842
rect 878 837 879 841
rect 883 837 884 841
rect 878 836 884 837
rect 998 841 1004 842
rect 998 837 999 841
rect 1003 837 1004 841
rect 998 836 1004 837
rect 1110 841 1116 842
rect 1110 837 1111 841
rect 1115 837 1116 841
rect 1110 836 1116 837
rect 1230 841 1236 842
rect 1230 837 1231 841
rect 1235 837 1236 841
rect 1230 836 1236 837
rect 1350 841 1356 842
rect 1350 837 1351 841
rect 1355 837 1356 841
rect 1350 836 1356 837
rect 2006 840 2012 841
rect 2006 836 2007 840
rect 2011 836 2012 840
rect 2906 839 2912 840
rect 2906 838 2907 839
rect 110 835 116 836
rect 2006 835 2012 836
rect 2625 836 2907 838
rect 2625 832 2627 836
rect 2906 835 2907 836
rect 2911 835 2912 839
rect 3642 839 3648 840
rect 3642 838 3643 839
rect 2906 834 2912 835
rect 3604 836 3643 838
rect 2623 831 2629 832
rect 2623 827 2624 831
rect 2628 827 2629 831
rect 2623 826 2629 827
rect 2634 831 2640 832
rect 2634 827 2635 831
rect 2639 830 2640 831
rect 2743 831 2749 832
rect 2743 830 2744 831
rect 2639 828 2744 830
rect 2639 827 2640 828
rect 2634 826 2640 827
rect 2743 827 2744 828
rect 2748 827 2749 831
rect 2743 826 2749 827
rect 2754 831 2760 832
rect 2754 827 2755 831
rect 2759 830 2760 831
rect 2871 831 2877 832
rect 2871 830 2872 831
rect 2759 828 2872 830
rect 2759 827 2760 828
rect 2754 826 2760 827
rect 2871 827 2872 828
rect 2876 827 2877 831
rect 2871 826 2877 827
rect 2882 831 2888 832
rect 2882 827 2883 831
rect 2887 830 2888 831
rect 3007 831 3013 832
rect 3007 830 3008 831
rect 2887 828 3008 830
rect 2887 827 2888 828
rect 2882 826 2888 827
rect 3007 827 3008 828
rect 3012 827 3013 831
rect 3007 826 3013 827
rect 3018 831 3024 832
rect 3018 827 3019 831
rect 3023 830 3024 831
rect 3143 831 3149 832
rect 3143 830 3144 831
rect 3023 828 3144 830
rect 3023 827 3024 828
rect 3018 826 3024 827
rect 3143 827 3144 828
rect 3148 827 3149 831
rect 3143 826 3149 827
rect 3271 831 3277 832
rect 3271 827 3272 831
rect 3276 830 3277 831
rect 3290 831 3296 832
rect 3290 830 3291 831
rect 3276 828 3291 830
rect 3276 827 3277 828
rect 3271 826 3277 827
rect 3290 827 3291 828
rect 3295 827 3296 831
rect 3290 826 3296 827
rect 3399 831 3405 832
rect 3399 827 3400 831
rect 3404 830 3405 831
rect 3418 831 3424 832
rect 3418 830 3419 831
rect 3404 828 3419 830
rect 3404 827 3405 828
rect 3399 826 3405 827
rect 3418 827 3419 828
rect 3423 827 3424 831
rect 3418 826 3424 827
rect 3527 831 3533 832
rect 3527 827 3528 831
rect 3532 830 3533 831
rect 3604 830 3606 836
rect 3642 835 3643 836
rect 3647 835 3648 839
rect 3642 834 3648 835
rect 3532 828 3606 830
rect 3618 831 3624 832
rect 3532 827 3533 828
rect 3527 826 3533 827
rect 3618 827 3619 831
rect 3623 830 3624 831
rect 3655 831 3661 832
rect 3655 830 3656 831
rect 3623 828 3656 830
rect 3623 827 3624 828
rect 3618 826 3624 827
rect 3655 827 3656 828
rect 3660 827 3661 831
rect 3655 826 3661 827
rect 3666 831 3672 832
rect 3666 827 3667 831
rect 3671 830 3672 831
rect 3791 831 3797 832
rect 3791 830 3792 831
rect 3671 828 3792 830
rect 3671 827 3672 828
rect 3666 826 3672 827
rect 3791 827 3792 828
rect 3796 827 3797 831
rect 3791 826 3797 827
rect 3903 831 3909 832
rect 3903 827 3904 831
rect 3908 830 3909 831
rect 3914 831 3920 832
rect 3914 830 3915 831
rect 3908 828 3915 830
rect 3908 827 3909 828
rect 3903 826 3909 827
rect 3914 827 3915 828
rect 3919 827 3920 831
rect 3914 826 3920 827
rect 214 819 220 820
rect 214 815 215 819
rect 219 818 220 819
rect 223 819 229 820
rect 223 818 224 819
rect 219 816 224 818
rect 219 815 220 816
rect 214 814 220 815
rect 223 815 224 816
rect 228 815 229 819
rect 223 814 229 815
rect 234 819 240 820
rect 234 815 235 819
rect 239 818 240 819
rect 383 819 389 820
rect 383 818 384 819
rect 239 816 384 818
rect 239 815 240 816
rect 234 814 240 815
rect 383 815 384 816
rect 388 815 389 819
rect 383 814 389 815
rect 535 819 541 820
rect 535 815 536 819
rect 540 818 541 819
rect 554 819 560 820
rect 554 818 555 819
rect 540 816 555 818
rect 540 815 541 816
rect 535 814 541 815
rect 554 815 555 816
rect 559 815 560 819
rect 554 814 560 815
rect 679 819 685 820
rect 679 815 680 819
rect 684 818 685 819
rect 698 819 704 820
rect 698 818 699 819
rect 684 816 699 818
rect 684 815 685 816
rect 679 814 685 815
rect 698 815 699 816
rect 703 815 704 819
rect 698 814 704 815
rect 714 819 720 820
rect 714 815 715 819
rect 719 818 720 819
rect 815 819 821 820
rect 815 818 816 819
rect 719 816 816 818
rect 719 815 720 816
rect 714 814 720 815
rect 815 815 816 816
rect 820 815 821 819
rect 815 814 821 815
rect 942 819 949 820
rect 942 815 943 819
rect 948 815 949 819
rect 942 814 949 815
rect 990 819 996 820
rect 990 815 991 819
rect 995 818 996 819
rect 1063 819 1069 820
rect 1063 818 1064 819
rect 995 816 1064 818
rect 995 815 996 816
rect 990 814 996 815
rect 1063 815 1064 816
rect 1068 815 1069 819
rect 1063 814 1069 815
rect 1098 819 1104 820
rect 1098 815 1099 819
rect 1103 818 1104 819
rect 1175 819 1181 820
rect 1175 818 1176 819
rect 1103 816 1176 818
rect 1103 815 1104 816
rect 1098 814 1104 815
rect 1175 815 1176 816
rect 1180 815 1181 819
rect 1175 814 1181 815
rect 1186 819 1192 820
rect 1186 815 1187 819
rect 1191 818 1192 819
rect 1295 819 1301 820
rect 1295 818 1296 819
rect 1191 816 1296 818
rect 1191 815 1192 816
rect 1186 814 1192 815
rect 1295 815 1296 816
rect 1300 815 1301 819
rect 1295 814 1301 815
rect 1306 819 1312 820
rect 1306 815 1307 819
rect 1311 818 1312 819
rect 1415 819 1421 820
rect 1415 818 1416 819
rect 1311 816 1416 818
rect 1311 815 1312 816
rect 1306 814 1312 815
rect 1415 815 1416 816
rect 1420 815 1421 819
rect 1415 814 1421 815
rect 2399 815 2405 816
rect 2399 811 2400 815
rect 2404 814 2405 815
rect 2410 815 2416 816
rect 2404 811 2406 814
rect 2399 810 2406 811
rect 2410 811 2411 815
rect 2415 814 2416 815
rect 2535 815 2541 816
rect 2535 814 2536 815
rect 2415 812 2536 814
rect 2415 811 2416 812
rect 2410 810 2416 811
rect 2535 811 2536 812
rect 2540 811 2541 815
rect 2535 810 2541 811
rect 2546 815 2552 816
rect 2546 811 2547 815
rect 2551 814 2552 815
rect 2679 815 2685 816
rect 2679 814 2680 815
rect 2551 812 2680 814
rect 2551 811 2552 812
rect 2546 810 2552 811
rect 2679 811 2680 812
rect 2684 811 2685 815
rect 2679 810 2685 811
rect 2831 815 2837 816
rect 2831 811 2832 815
rect 2836 814 2837 815
rect 2854 815 2860 816
rect 2854 814 2855 815
rect 2836 812 2855 814
rect 2836 811 2837 812
rect 2831 810 2837 811
rect 2854 811 2855 812
rect 2859 811 2860 815
rect 2854 810 2860 811
rect 2983 815 2989 816
rect 2983 811 2984 815
rect 2988 814 2989 815
rect 3026 815 3032 816
rect 3026 814 3027 815
rect 2988 812 3027 814
rect 2988 811 2989 812
rect 2983 810 2989 811
rect 3026 811 3027 812
rect 3031 811 3032 815
rect 3026 810 3032 811
rect 3143 815 3149 816
rect 3143 811 3144 815
rect 3148 814 3149 815
rect 3162 815 3168 816
rect 3162 814 3163 815
rect 3148 812 3163 814
rect 3148 811 3149 812
rect 3143 810 3149 811
rect 3162 811 3163 812
rect 3167 811 3168 815
rect 3162 810 3168 811
rect 3207 815 3213 816
rect 3207 811 3208 815
rect 3212 814 3213 815
rect 3303 815 3309 816
rect 3303 814 3304 815
rect 3212 812 3304 814
rect 3212 811 3213 812
rect 3207 810 3213 811
rect 3303 811 3304 812
rect 3308 811 3309 815
rect 3303 810 3309 811
rect 3314 815 3320 816
rect 3314 811 3315 815
rect 3319 814 3320 815
rect 3455 815 3461 816
rect 3455 814 3456 815
rect 3319 812 3456 814
rect 3319 811 3320 812
rect 3314 810 3320 811
rect 3455 811 3456 812
rect 3460 811 3461 815
rect 3455 810 3461 811
rect 3607 815 3613 816
rect 3607 811 3608 815
rect 3612 814 3613 815
rect 3642 815 3648 816
rect 3642 814 3643 815
rect 3612 812 3643 814
rect 3612 811 3613 812
rect 3607 810 3613 811
rect 3642 811 3643 812
rect 3647 811 3648 815
rect 3642 810 3648 811
rect 3767 815 3776 816
rect 3767 811 3768 815
rect 3775 811 3776 815
rect 3767 810 3776 811
rect 3903 815 3912 816
rect 3903 811 3904 815
rect 3911 811 3912 815
rect 3903 810 3912 811
rect 287 807 293 808
rect 287 803 288 807
rect 292 806 293 807
rect 306 807 312 808
rect 306 806 307 807
rect 292 804 307 806
rect 292 803 293 804
rect 287 802 293 803
rect 306 803 307 804
rect 311 803 312 807
rect 306 802 312 803
rect 402 807 408 808
rect 402 803 403 807
rect 407 806 408 807
rect 447 807 453 808
rect 447 806 448 807
rect 407 804 448 806
rect 407 803 408 804
rect 402 802 408 803
rect 447 803 448 804
rect 452 803 453 807
rect 447 802 453 803
rect 546 807 552 808
rect 546 803 547 807
rect 551 806 552 807
rect 599 807 605 808
rect 599 806 600 807
rect 551 804 600 806
rect 551 803 552 804
rect 546 802 552 803
rect 599 803 600 804
rect 604 803 605 807
rect 599 802 605 803
rect 634 807 640 808
rect 634 803 635 807
rect 639 806 640 807
rect 743 807 749 808
rect 743 806 744 807
rect 639 804 744 806
rect 639 803 640 804
rect 634 802 640 803
rect 743 803 744 804
rect 748 803 749 807
rect 743 802 749 803
rect 798 807 804 808
rect 798 803 799 807
rect 803 806 804 807
rect 879 807 885 808
rect 879 806 880 807
rect 803 804 880 806
rect 803 803 804 804
rect 798 802 804 803
rect 879 803 880 804
rect 884 803 885 807
rect 879 802 885 803
rect 1015 807 1021 808
rect 1015 803 1016 807
rect 1020 806 1021 807
rect 1066 807 1072 808
rect 1066 806 1067 807
rect 1020 804 1067 806
rect 1020 803 1021 804
rect 1015 802 1021 803
rect 1066 803 1067 804
rect 1071 803 1072 807
rect 1066 802 1072 803
rect 1143 807 1149 808
rect 1143 803 1144 807
rect 1148 806 1149 807
rect 1178 807 1184 808
rect 1178 806 1179 807
rect 1148 804 1179 806
rect 1148 803 1149 804
rect 1143 802 1149 803
rect 1178 803 1179 804
rect 1183 803 1184 807
rect 1178 802 1184 803
rect 1263 807 1269 808
rect 1263 803 1264 807
rect 1268 806 1269 807
rect 1370 807 1376 808
rect 1268 804 1366 806
rect 1268 803 1269 804
rect 1263 802 1269 803
rect 1364 798 1366 804
rect 1370 803 1371 807
rect 1375 806 1376 807
rect 1391 807 1397 808
rect 1391 806 1392 807
rect 1375 804 1392 806
rect 1375 803 1376 804
rect 1370 802 1376 803
rect 1391 803 1392 804
rect 1396 803 1397 807
rect 1391 802 1397 803
rect 1402 807 1408 808
rect 1402 803 1403 807
rect 1407 806 1408 807
rect 1519 807 1525 808
rect 1519 806 1520 807
rect 1407 804 1520 806
rect 1407 803 1408 804
rect 1402 802 1408 803
rect 1519 803 1520 804
rect 1524 803 1525 807
rect 2404 806 2406 810
rect 2718 807 2724 808
rect 2718 806 2719 807
rect 2404 804 2719 806
rect 1519 802 1525 803
rect 2718 803 2719 804
rect 2723 803 2724 807
rect 2718 802 2724 803
rect 1410 799 1416 800
rect 1410 798 1411 799
rect 1364 796 1411 798
rect 1410 795 1411 796
rect 1415 795 1416 799
rect 1410 794 1416 795
rect 2046 796 2052 797
rect 3942 796 3948 797
rect 2046 792 2047 796
rect 2051 792 2052 796
rect 2046 791 2052 792
rect 2334 795 2340 796
rect 2334 791 2335 795
rect 2339 791 2340 795
rect 2334 790 2340 791
rect 2470 795 2476 796
rect 2470 791 2471 795
rect 2475 791 2476 795
rect 2470 790 2476 791
rect 2614 795 2620 796
rect 2614 791 2615 795
rect 2619 791 2620 795
rect 2614 790 2620 791
rect 2766 795 2772 796
rect 2766 791 2767 795
rect 2771 791 2772 795
rect 2766 790 2772 791
rect 2918 795 2924 796
rect 2918 791 2919 795
rect 2923 791 2924 795
rect 2918 790 2924 791
rect 3078 795 3084 796
rect 3078 791 3079 795
rect 3083 791 3084 795
rect 3078 790 3084 791
rect 3238 795 3244 796
rect 3238 791 3239 795
rect 3243 791 3244 795
rect 3238 790 3244 791
rect 3390 795 3396 796
rect 3390 791 3391 795
rect 3395 791 3396 795
rect 3390 790 3396 791
rect 3542 795 3548 796
rect 3542 791 3543 795
rect 3547 791 3548 795
rect 3542 790 3548 791
rect 3702 795 3708 796
rect 3702 791 3703 795
rect 3707 791 3708 795
rect 3702 790 3708 791
rect 3838 795 3844 796
rect 3838 791 3839 795
rect 3843 791 3844 795
rect 3942 792 3943 796
rect 3947 792 3948 796
rect 3942 791 3948 792
rect 3838 790 3844 791
rect 110 788 116 789
rect 2006 788 2012 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 222 787 228 788
rect 222 783 223 787
rect 227 783 228 787
rect 222 782 228 783
rect 382 787 388 788
rect 382 783 383 787
rect 387 783 388 787
rect 382 782 388 783
rect 534 787 540 788
rect 534 783 535 787
rect 539 783 540 787
rect 534 782 540 783
rect 678 787 684 788
rect 678 783 679 787
rect 683 783 684 787
rect 678 782 684 783
rect 814 787 820 788
rect 814 783 815 787
rect 819 783 820 787
rect 814 782 820 783
rect 950 787 956 788
rect 950 783 951 787
rect 955 783 956 787
rect 950 782 956 783
rect 1078 787 1084 788
rect 1078 783 1079 787
rect 1083 783 1084 787
rect 1078 782 1084 783
rect 1198 787 1204 788
rect 1198 783 1199 787
rect 1203 783 1204 787
rect 1198 782 1204 783
rect 1326 787 1332 788
rect 1326 783 1327 787
rect 1331 783 1332 787
rect 1326 782 1332 783
rect 1454 787 1460 788
rect 1454 783 1455 787
rect 1459 783 1460 787
rect 2006 784 2007 788
rect 2011 784 2012 788
rect 2006 783 2012 784
rect 2410 787 2416 788
rect 2410 783 2411 787
rect 2415 783 2416 787
rect 1454 782 1460 783
rect 2410 782 2416 783
rect 2546 787 2552 788
rect 2546 783 2547 787
rect 2551 783 2552 787
rect 2718 787 2724 788
rect 2546 782 2552 783
rect 2690 783 2696 784
rect 214 779 220 780
rect 214 775 215 779
rect 219 778 220 779
rect 306 779 312 780
rect 219 776 265 778
rect 219 775 220 776
rect 214 774 220 775
rect 306 775 307 779
rect 311 778 312 779
rect 634 779 640 780
rect 634 778 635 779
rect 311 776 425 778
rect 613 776 635 778
rect 311 775 312 776
rect 306 774 312 775
rect 634 775 635 776
rect 639 775 640 779
rect 798 779 804 780
rect 798 778 799 779
rect 757 776 799 778
rect 634 774 640 775
rect 798 775 799 776
rect 803 775 804 779
rect 942 779 948 780
rect 798 774 804 775
rect 890 775 896 776
rect 110 771 116 772
rect 110 767 111 771
rect 115 767 116 771
rect 890 771 891 775
rect 895 771 896 775
rect 942 775 943 779
rect 947 778 948 779
rect 1066 779 1072 780
rect 947 776 993 778
rect 947 775 948 776
rect 942 774 948 775
rect 1066 775 1067 779
rect 1071 778 1072 779
rect 1178 779 1184 780
rect 1071 776 1121 778
rect 1071 775 1072 776
rect 1066 774 1072 775
rect 1178 775 1179 779
rect 1183 778 1184 779
rect 1402 779 1408 780
rect 1183 776 1241 778
rect 1183 775 1184 776
rect 1178 774 1184 775
rect 1402 775 1403 779
rect 1407 775 1408 779
rect 1402 774 1408 775
rect 1410 779 1416 780
rect 1410 775 1411 779
rect 1415 778 1416 779
rect 2046 779 2052 780
rect 1415 776 1497 778
rect 1415 775 1416 776
rect 1410 774 1416 775
rect 2046 775 2047 779
rect 2051 775 2052 779
rect 2690 779 2691 783
rect 2695 779 2696 783
rect 2718 783 2719 787
rect 2723 786 2724 787
rect 2854 787 2860 788
rect 2723 784 2809 786
rect 2723 783 2724 784
rect 2718 782 2724 783
rect 2854 783 2855 787
rect 2859 786 2860 787
rect 3207 787 3213 788
rect 3207 786 3208 787
rect 2859 784 2961 786
rect 3157 784 3208 786
rect 2859 783 2860 784
rect 2854 782 2860 783
rect 3207 783 3208 784
rect 3212 783 3213 787
rect 3207 782 3213 783
rect 3314 787 3320 788
rect 3314 783 3315 787
rect 3319 783 3320 787
rect 3618 787 3624 788
rect 3314 782 3320 783
rect 3466 783 3472 784
rect 2690 778 2696 779
rect 3466 779 3467 783
rect 3471 779 3472 783
rect 3618 783 3619 787
rect 3623 783 3624 787
rect 3618 782 3624 783
rect 3642 787 3648 788
rect 3642 783 3643 787
rect 3647 786 3648 787
rect 3647 784 3745 786
rect 3647 783 3648 784
rect 3642 782 3648 783
rect 3914 783 3920 784
rect 3466 778 3472 779
rect 3914 779 3915 783
rect 3919 779 3920 783
rect 3914 778 3920 779
rect 3942 779 3948 780
rect 2046 774 2052 775
rect 2334 776 2340 777
rect 2334 772 2335 776
rect 2339 772 2340 776
rect 890 770 896 771
rect 2006 771 2012 772
rect 2334 771 2340 772
rect 2470 776 2476 777
rect 2470 772 2471 776
rect 2475 772 2476 776
rect 2470 771 2476 772
rect 2614 776 2620 777
rect 2614 772 2615 776
rect 2619 772 2620 776
rect 2614 771 2620 772
rect 2766 776 2772 777
rect 2766 772 2767 776
rect 2771 772 2772 776
rect 2766 771 2772 772
rect 2918 776 2924 777
rect 2918 772 2919 776
rect 2923 772 2924 776
rect 2918 771 2924 772
rect 3078 776 3084 777
rect 3078 772 3079 776
rect 3083 772 3084 776
rect 3078 771 3084 772
rect 3238 776 3244 777
rect 3238 772 3239 776
rect 3243 772 3244 776
rect 3238 771 3244 772
rect 3390 776 3396 777
rect 3390 772 3391 776
rect 3395 772 3396 776
rect 3390 771 3396 772
rect 3542 776 3548 777
rect 3542 772 3543 776
rect 3547 772 3548 776
rect 3542 771 3548 772
rect 3702 776 3708 777
rect 3702 772 3703 776
rect 3707 772 3708 776
rect 3702 771 3708 772
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3942 775 3943 779
rect 3947 775 3948 779
rect 3942 774 3948 775
rect 3838 771 3844 772
rect 110 766 116 767
rect 222 768 228 769
rect 222 764 223 768
rect 227 764 228 768
rect 222 763 228 764
rect 382 768 388 769
rect 382 764 383 768
rect 387 764 388 768
rect 382 763 388 764
rect 534 768 540 769
rect 534 764 535 768
rect 539 764 540 768
rect 534 763 540 764
rect 678 768 684 769
rect 678 764 679 768
rect 683 764 684 768
rect 678 763 684 764
rect 814 768 820 769
rect 814 764 815 768
rect 819 764 820 768
rect 814 763 820 764
rect 950 768 956 769
rect 950 764 951 768
rect 955 764 956 768
rect 950 763 956 764
rect 1078 768 1084 769
rect 1078 764 1079 768
rect 1083 764 1084 768
rect 1078 763 1084 764
rect 1198 768 1204 769
rect 1198 764 1199 768
rect 1203 764 1204 768
rect 1198 763 1204 764
rect 1326 768 1332 769
rect 1326 764 1327 768
rect 1331 764 1332 768
rect 1326 763 1332 764
rect 1454 768 1460 769
rect 1454 764 1455 768
rect 1459 764 1460 768
rect 2006 767 2007 771
rect 2011 767 2012 771
rect 2006 766 2012 767
rect 1454 763 1460 764
rect 2070 712 2076 713
rect 2046 709 2052 710
rect 2046 705 2047 709
rect 2051 705 2052 709
rect 2070 708 2071 712
rect 2075 708 2076 712
rect 2070 707 2076 708
rect 2182 712 2188 713
rect 2182 708 2183 712
rect 2187 708 2188 712
rect 2182 707 2188 708
rect 2334 712 2340 713
rect 2334 708 2335 712
rect 2339 708 2340 712
rect 2334 707 2340 708
rect 2486 712 2492 713
rect 2486 708 2487 712
rect 2491 708 2492 712
rect 2486 707 2492 708
rect 2638 712 2644 713
rect 2638 708 2639 712
rect 2643 708 2644 712
rect 2638 707 2644 708
rect 2806 712 2812 713
rect 2806 708 2807 712
rect 2811 708 2812 712
rect 2806 707 2812 708
rect 2982 712 2988 713
rect 2982 708 2983 712
rect 2987 708 2988 712
rect 2982 707 2988 708
rect 3166 712 3172 713
rect 3166 708 3167 712
rect 3171 708 3172 712
rect 3166 707 3172 708
rect 3366 712 3372 713
rect 3366 708 3367 712
rect 3371 708 3372 712
rect 3366 707 3372 708
rect 3574 712 3580 713
rect 3574 708 3575 712
rect 3579 708 3580 712
rect 3574 707 3580 708
rect 3782 712 3788 713
rect 3782 708 3783 712
rect 3787 708 3788 712
rect 3782 707 3788 708
rect 3942 709 3948 710
rect 310 704 316 705
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 310 700 311 704
rect 315 700 316 704
rect 310 699 316 700
rect 470 704 476 705
rect 470 700 471 704
rect 475 700 476 704
rect 470 699 476 700
rect 638 704 644 705
rect 638 700 639 704
rect 643 700 644 704
rect 638 699 644 700
rect 806 704 812 705
rect 806 700 807 704
rect 811 700 812 704
rect 806 699 812 700
rect 974 704 980 705
rect 974 700 975 704
rect 979 700 980 704
rect 974 699 980 700
rect 1134 704 1140 705
rect 1134 700 1135 704
rect 1139 700 1140 704
rect 1134 699 1140 700
rect 1294 704 1300 705
rect 1294 700 1295 704
rect 1299 700 1300 704
rect 1294 699 1300 700
rect 1454 704 1460 705
rect 1454 700 1455 704
rect 1459 700 1460 704
rect 1454 699 1460 700
rect 1606 704 1612 705
rect 1606 700 1607 704
rect 1611 700 1612 704
rect 1606 699 1612 700
rect 1766 704 1772 705
rect 1766 700 1767 704
rect 1771 700 1772 704
rect 1766 699 1772 700
rect 1902 704 1908 705
rect 2046 704 2052 705
rect 3942 705 3943 709
rect 3947 705 3948 709
rect 3942 704 3948 705
rect 1902 700 1903 704
rect 1907 700 1908 704
rect 2054 703 2060 704
rect 1902 699 1908 700
rect 2006 701 2012 702
rect 110 696 116 697
rect 2006 697 2007 701
rect 2011 697 2012 701
rect 2054 699 2055 703
rect 2059 702 2060 703
rect 2154 703 2160 704
rect 2059 700 2113 702
rect 2059 699 2060 700
rect 2054 698 2060 699
rect 2154 699 2155 703
rect 2159 702 2160 703
rect 2266 703 2272 704
rect 2159 700 2225 702
rect 2159 699 2160 700
rect 2154 698 2160 699
rect 2266 699 2267 703
rect 2271 702 2272 703
rect 2418 703 2424 704
rect 2271 700 2377 702
rect 2271 699 2272 700
rect 2266 698 2272 699
rect 2418 699 2419 703
rect 2423 702 2424 703
rect 2570 703 2576 704
rect 2423 700 2529 702
rect 2423 699 2424 700
rect 2418 698 2424 699
rect 2570 699 2571 703
rect 2575 702 2576 703
rect 2882 703 2888 704
rect 2575 700 2681 702
rect 2575 699 2576 700
rect 2570 698 2576 699
rect 2882 699 2883 703
rect 2887 699 2888 703
rect 2882 698 2888 699
rect 3058 703 3064 704
rect 3058 699 3059 703
rect 3063 699 3064 703
rect 3058 698 3064 699
rect 3242 703 3248 704
rect 3242 699 3243 703
rect 3247 699 3248 703
rect 3242 698 3248 699
rect 3318 703 3324 704
rect 3318 699 3319 703
rect 3323 702 3324 703
rect 3450 703 3456 704
rect 3323 700 3409 702
rect 3323 699 3324 700
rect 3318 698 3324 699
rect 3450 699 3451 703
rect 3455 702 3456 703
rect 3770 703 3776 704
rect 3455 700 3617 702
rect 3455 699 3456 700
rect 3450 698 3456 699
rect 3770 699 3771 703
rect 3775 702 3776 703
rect 3775 700 3825 702
rect 3775 699 3776 700
rect 3770 698 3776 699
rect 2006 696 2012 697
rect 402 695 408 696
rect 402 694 403 695
rect 389 692 403 694
rect 402 691 403 692
rect 407 691 408 695
rect 402 690 408 691
rect 546 695 552 696
rect 546 691 547 695
rect 551 691 552 695
rect 546 690 552 691
rect 554 695 560 696
rect 554 691 555 695
rect 559 694 560 695
rect 942 695 948 696
rect 942 694 943 695
rect 559 692 681 694
rect 885 692 943 694
rect 559 691 560 692
rect 554 690 560 691
rect 942 691 943 692
rect 947 691 948 695
rect 942 690 948 691
rect 1042 695 1048 696
rect 1042 691 1043 695
rect 1047 691 1048 695
rect 1042 690 1048 691
rect 1210 695 1216 696
rect 1210 691 1211 695
rect 1215 691 1216 695
rect 1210 690 1216 691
rect 1370 695 1376 696
rect 1370 691 1371 695
rect 1375 691 1376 695
rect 1582 695 1588 696
rect 1582 694 1583 695
rect 1533 692 1583 694
rect 1370 690 1376 691
rect 1582 691 1583 692
rect 1587 691 1588 695
rect 1582 690 1588 691
rect 1682 695 1688 696
rect 1682 691 1683 695
rect 1687 691 1688 695
rect 1682 690 1688 691
rect 1698 695 1704 696
rect 1698 691 1699 695
rect 1703 694 1704 695
rect 1858 695 1864 696
rect 1703 692 1809 694
rect 1703 691 1704 692
rect 1698 690 1704 691
rect 1858 691 1859 695
rect 1863 694 1864 695
rect 1863 692 1945 694
rect 2070 693 2076 694
rect 2046 692 2052 693
rect 1863 691 1864 692
rect 1858 690 1864 691
rect 2046 688 2047 692
rect 2051 688 2052 692
rect 2070 689 2071 693
rect 2075 689 2076 693
rect 2070 688 2076 689
rect 2182 693 2188 694
rect 2182 689 2183 693
rect 2187 689 2188 693
rect 2182 688 2188 689
rect 2334 693 2340 694
rect 2334 689 2335 693
rect 2339 689 2340 693
rect 2334 688 2340 689
rect 2486 693 2492 694
rect 2486 689 2487 693
rect 2491 689 2492 693
rect 2486 688 2492 689
rect 2638 693 2644 694
rect 2638 689 2639 693
rect 2643 689 2644 693
rect 2638 688 2644 689
rect 2806 693 2812 694
rect 2806 689 2807 693
rect 2811 689 2812 693
rect 2806 688 2812 689
rect 2982 693 2988 694
rect 2982 689 2983 693
rect 2987 689 2988 693
rect 2982 688 2988 689
rect 3166 693 3172 694
rect 3166 689 3167 693
rect 3171 689 3172 693
rect 3166 688 3172 689
rect 3366 693 3372 694
rect 3366 689 3367 693
rect 3371 689 3372 693
rect 3366 688 3372 689
rect 3574 693 3580 694
rect 3574 689 3575 693
rect 3579 689 3580 693
rect 3574 688 3580 689
rect 3782 693 3788 694
rect 3782 689 3783 693
rect 3787 689 3788 693
rect 3782 688 3788 689
rect 3942 692 3948 693
rect 3942 688 3943 692
rect 3947 688 3948 692
rect 2046 687 2052 688
rect 3942 687 3948 688
rect 310 685 316 686
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 310 681 311 685
rect 315 681 316 685
rect 310 680 316 681
rect 470 685 476 686
rect 470 681 471 685
rect 475 681 476 685
rect 470 680 476 681
rect 638 685 644 686
rect 638 681 639 685
rect 643 681 644 685
rect 638 680 644 681
rect 806 685 812 686
rect 806 681 807 685
rect 811 681 812 685
rect 806 680 812 681
rect 974 685 980 686
rect 974 681 975 685
rect 979 681 980 685
rect 974 680 980 681
rect 1134 685 1140 686
rect 1134 681 1135 685
rect 1139 681 1140 685
rect 1134 680 1140 681
rect 1294 685 1300 686
rect 1294 681 1295 685
rect 1299 681 1300 685
rect 1294 680 1300 681
rect 1454 685 1460 686
rect 1454 681 1455 685
rect 1459 681 1460 685
rect 1454 680 1460 681
rect 1606 685 1612 686
rect 1606 681 1607 685
rect 1611 681 1612 685
rect 1606 680 1612 681
rect 1766 685 1772 686
rect 1766 681 1767 685
rect 1771 681 1772 685
rect 1766 680 1772 681
rect 1902 685 1908 686
rect 1902 681 1903 685
rect 1907 681 1908 685
rect 1902 680 1908 681
rect 2006 684 2012 685
rect 2006 680 2007 684
rect 2011 680 2012 684
rect 110 679 116 680
rect 2006 679 2012 680
rect 3318 679 3324 680
rect 3318 678 3319 679
rect 2876 676 3319 678
rect 2876 672 2878 676
rect 3318 675 3319 676
rect 3323 675 3324 679
rect 3318 674 3324 675
rect 3466 675 3472 676
rect 554 671 560 672
rect 554 670 555 671
rect 516 668 555 670
rect 375 663 381 664
rect 375 659 376 663
rect 380 662 381 663
rect 516 662 518 668
rect 554 667 555 668
rect 559 667 560 671
rect 554 666 560 667
rect 2135 671 2141 672
rect 2135 667 2136 671
rect 2140 670 2141 671
rect 2154 671 2160 672
rect 2154 670 2155 671
rect 2140 668 2155 670
rect 2140 667 2141 668
rect 2135 666 2141 667
rect 2154 667 2155 668
rect 2159 667 2160 671
rect 2154 666 2160 667
rect 2247 671 2253 672
rect 2247 667 2248 671
rect 2252 670 2253 671
rect 2266 671 2272 672
rect 2266 670 2267 671
rect 2252 668 2267 670
rect 2252 667 2253 668
rect 2247 666 2253 667
rect 2266 667 2267 668
rect 2271 667 2272 671
rect 2266 666 2272 667
rect 2399 671 2405 672
rect 2399 667 2400 671
rect 2404 670 2405 671
rect 2418 671 2424 672
rect 2418 670 2419 671
rect 2404 668 2419 670
rect 2404 667 2405 668
rect 2399 666 2405 667
rect 2418 667 2419 668
rect 2423 667 2424 671
rect 2418 666 2424 667
rect 2551 671 2557 672
rect 2551 667 2552 671
rect 2556 670 2557 671
rect 2570 671 2576 672
rect 2570 670 2571 671
rect 2556 668 2571 670
rect 2556 667 2557 668
rect 2551 666 2557 667
rect 2570 667 2571 668
rect 2575 667 2576 671
rect 2570 666 2576 667
rect 2690 671 2696 672
rect 2690 667 2691 671
rect 2695 670 2696 671
rect 2703 671 2709 672
rect 2703 670 2704 671
rect 2695 668 2704 670
rect 2695 667 2696 668
rect 2690 666 2696 667
rect 2703 667 2704 668
rect 2708 667 2709 671
rect 2703 666 2709 667
rect 2871 671 2878 672
rect 2871 667 2872 671
rect 2876 668 2878 671
rect 2882 671 2888 672
rect 2876 667 2877 668
rect 2871 666 2877 667
rect 2882 667 2883 671
rect 2887 670 2888 671
rect 3047 671 3053 672
rect 3047 670 3048 671
rect 2887 668 3048 670
rect 2887 667 2888 668
rect 2882 666 2888 667
rect 3047 667 3048 668
rect 3052 667 3053 671
rect 3047 666 3053 667
rect 3058 671 3064 672
rect 3058 667 3059 671
rect 3063 670 3064 671
rect 3231 671 3237 672
rect 3231 670 3232 671
rect 3063 668 3232 670
rect 3063 667 3064 668
rect 3058 666 3064 667
rect 3231 667 3232 668
rect 3236 667 3237 671
rect 3231 666 3237 667
rect 3431 671 3437 672
rect 3431 667 3432 671
rect 3436 670 3437 671
rect 3450 671 3456 672
rect 3450 670 3451 671
rect 3436 668 3451 670
rect 3436 667 3437 668
rect 3431 666 3437 667
rect 3450 667 3451 668
rect 3455 667 3456 671
rect 3466 671 3467 675
rect 3471 674 3472 675
rect 3471 672 3562 674
rect 3471 671 3472 672
rect 3466 670 3472 671
rect 3560 670 3562 672
rect 3639 671 3645 672
rect 3639 670 3640 671
rect 3560 668 3640 670
rect 3450 666 3456 667
rect 3639 667 3640 668
rect 3644 667 3645 671
rect 3639 666 3645 667
rect 3847 671 3853 672
rect 3847 667 3848 671
rect 3852 670 3853 671
rect 3874 671 3880 672
rect 3874 670 3875 671
rect 3852 668 3875 670
rect 3852 667 3853 668
rect 3847 666 3853 667
rect 3874 667 3875 668
rect 3879 667 3880 671
rect 3874 666 3880 667
rect 380 660 518 662
rect 522 663 528 664
rect 380 659 381 660
rect 375 658 381 659
rect 522 659 523 663
rect 527 662 528 663
rect 535 663 541 664
rect 535 662 536 663
rect 527 660 536 662
rect 527 659 528 660
rect 522 658 528 659
rect 535 659 536 660
rect 540 659 541 663
rect 535 658 541 659
rect 546 663 552 664
rect 546 659 547 663
rect 551 662 552 663
rect 703 663 709 664
rect 703 662 704 663
rect 551 660 704 662
rect 551 659 552 660
rect 546 658 552 659
rect 703 659 704 660
rect 708 659 709 663
rect 703 658 709 659
rect 871 663 877 664
rect 871 659 872 663
rect 876 662 877 663
rect 890 663 896 664
rect 890 662 891 663
rect 876 660 891 662
rect 876 659 877 660
rect 871 658 877 659
rect 890 659 891 660
rect 895 659 896 663
rect 890 658 896 659
rect 942 663 948 664
rect 942 659 943 663
rect 947 662 948 663
rect 1039 663 1045 664
rect 1039 662 1040 663
rect 947 660 1040 662
rect 947 659 948 660
rect 942 658 948 659
rect 1039 659 1040 660
rect 1044 659 1045 663
rect 1039 658 1045 659
rect 1199 663 1208 664
rect 1199 659 1200 663
rect 1207 659 1208 663
rect 1199 658 1208 659
rect 1210 663 1216 664
rect 1210 659 1211 663
rect 1215 662 1216 663
rect 1359 663 1365 664
rect 1359 662 1360 663
rect 1215 660 1360 662
rect 1215 659 1216 660
rect 1210 658 1216 659
rect 1359 659 1360 660
rect 1364 659 1365 663
rect 1359 658 1365 659
rect 1474 663 1480 664
rect 1474 659 1475 663
rect 1479 662 1480 663
rect 1519 663 1525 664
rect 1519 662 1520 663
rect 1479 660 1520 662
rect 1479 659 1480 660
rect 1474 658 1480 659
rect 1519 659 1520 660
rect 1524 659 1525 663
rect 1519 658 1525 659
rect 1582 663 1588 664
rect 1582 659 1583 663
rect 1587 662 1588 663
rect 1671 663 1677 664
rect 1671 662 1672 663
rect 1587 660 1672 662
rect 1587 659 1588 660
rect 1582 658 1588 659
rect 1671 659 1672 660
rect 1676 659 1677 663
rect 1671 658 1677 659
rect 1682 663 1688 664
rect 1682 659 1683 663
rect 1687 662 1688 663
rect 1831 663 1837 664
rect 1831 662 1832 663
rect 1687 660 1832 662
rect 1687 659 1688 660
rect 1682 658 1688 659
rect 1831 659 1832 660
rect 1836 659 1837 663
rect 1831 658 1837 659
rect 1967 663 1973 664
rect 1967 659 1968 663
rect 1972 662 1973 663
rect 2054 663 2060 664
rect 2054 662 2055 663
rect 1972 660 2055 662
rect 1972 659 1973 660
rect 1967 658 1973 659
rect 2054 659 2055 660
rect 2059 659 2060 663
rect 2054 658 2060 659
rect 359 651 365 652
rect 359 650 360 651
rect 319 648 360 650
rect 314 647 321 648
rect 314 643 315 647
rect 319 644 321 647
rect 359 647 360 648
rect 364 647 365 651
rect 359 646 365 647
rect 370 651 376 652
rect 370 647 371 651
rect 375 650 376 651
rect 511 651 517 652
rect 511 650 512 651
rect 375 648 512 650
rect 375 647 376 648
rect 370 646 376 647
rect 511 647 512 648
rect 516 647 517 651
rect 511 646 517 647
rect 679 651 685 652
rect 679 647 680 651
rect 684 650 685 651
rect 698 651 704 652
rect 698 650 699 651
rect 684 648 699 650
rect 684 647 685 648
rect 679 646 685 647
rect 698 647 699 648
rect 703 647 704 651
rect 698 646 704 647
rect 847 651 853 652
rect 847 647 848 651
rect 852 650 853 651
rect 866 651 872 652
rect 866 650 867 651
rect 852 648 867 650
rect 852 647 853 648
rect 847 646 853 647
rect 866 647 867 648
rect 871 647 872 651
rect 866 646 872 647
rect 1015 651 1021 652
rect 1015 647 1016 651
rect 1020 650 1021 651
rect 1042 651 1048 652
rect 1042 650 1043 651
rect 1020 648 1043 650
rect 1020 647 1021 648
rect 1015 646 1021 647
rect 1042 647 1043 648
rect 1047 647 1048 651
rect 1042 646 1048 647
rect 1175 651 1181 652
rect 1175 647 1176 651
rect 1180 650 1181 651
rect 1186 651 1192 652
rect 1180 647 1182 650
rect 1175 646 1182 647
rect 1186 647 1187 651
rect 1191 650 1192 651
rect 1327 651 1333 652
rect 1327 650 1328 651
rect 1191 648 1328 650
rect 1191 647 1192 648
rect 1186 646 1192 647
rect 1327 647 1328 648
rect 1332 647 1333 651
rect 1327 646 1333 647
rect 1338 651 1344 652
rect 1338 647 1339 651
rect 1343 650 1344 651
rect 1463 651 1469 652
rect 1463 650 1464 651
rect 1343 648 1464 650
rect 1343 647 1344 648
rect 1338 646 1344 647
rect 1463 647 1464 648
rect 1468 647 1469 651
rect 1463 646 1469 647
rect 1599 651 1605 652
rect 1599 647 1600 651
rect 1604 650 1605 651
rect 1618 651 1624 652
rect 1618 650 1619 651
rect 1604 648 1619 650
rect 1604 647 1605 648
rect 1599 646 1605 647
rect 1618 647 1619 648
rect 1623 647 1624 651
rect 1618 646 1624 647
rect 1727 651 1733 652
rect 1727 647 1728 651
rect 1732 650 1733 651
rect 1818 651 1824 652
rect 1818 650 1819 651
rect 1732 648 1819 650
rect 1732 647 1733 648
rect 1727 646 1733 647
rect 1818 647 1819 648
rect 1823 647 1824 651
rect 1818 646 1824 647
rect 1855 651 1864 652
rect 1855 647 1856 651
rect 1863 647 1864 651
rect 1855 646 1864 647
rect 1866 651 1872 652
rect 1866 647 1867 651
rect 1871 650 1872 651
rect 1967 651 1973 652
rect 1967 650 1968 651
rect 1871 648 1968 650
rect 1871 647 1872 648
rect 1866 646 1872 647
rect 1967 647 1968 648
rect 1972 647 1973 651
rect 1967 646 1973 647
rect 1978 647 1984 648
rect 319 643 320 644
rect 314 642 320 643
rect 1180 642 1182 646
rect 1482 643 1488 644
rect 1482 642 1483 643
rect 1180 640 1483 642
rect 1482 639 1483 640
rect 1487 639 1488 643
rect 1978 643 1979 647
rect 1983 646 1984 647
rect 2135 647 2141 648
rect 2135 646 2136 647
rect 1983 644 2136 646
rect 1983 643 1984 644
rect 1978 642 1984 643
rect 2135 643 2136 644
rect 2140 643 2141 647
rect 2135 642 2141 643
rect 2146 647 2152 648
rect 2146 643 2147 647
rect 2151 646 2152 647
rect 2303 647 2309 648
rect 2303 646 2304 647
rect 2151 644 2304 646
rect 2151 643 2152 644
rect 2146 642 2152 643
rect 2303 643 2304 644
rect 2308 643 2309 647
rect 2303 642 2309 643
rect 2314 647 2320 648
rect 2314 643 2315 647
rect 2319 646 2320 647
rect 2487 647 2493 648
rect 2487 646 2488 647
rect 2319 644 2488 646
rect 2319 643 2320 644
rect 2314 642 2320 643
rect 2487 643 2488 644
rect 2492 643 2493 647
rect 2487 642 2493 643
rect 2687 647 2693 648
rect 2687 643 2688 647
rect 2692 646 2693 647
rect 2762 647 2768 648
rect 2762 646 2763 647
rect 2692 644 2763 646
rect 2692 643 2693 644
rect 2687 642 2693 643
rect 2762 643 2763 644
rect 2767 643 2768 647
rect 2762 642 2768 643
rect 2903 647 2909 648
rect 2903 643 2904 647
rect 2908 646 2909 647
rect 2922 647 2928 648
rect 2922 646 2923 647
rect 2908 644 2923 646
rect 2908 643 2909 644
rect 2903 642 2909 643
rect 2922 643 2923 644
rect 2927 643 2928 647
rect 2922 642 2928 643
rect 3135 647 3141 648
rect 3135 643 3136 647
rect 3140 646 3141 647
rect 3242 647 3248 648
rect 3140 644 3238 646
rect 3140 643 3141 644
rect 3135 642 3141 643
rect 1482 638 1488 639
rect 3236 638 3238 644
rect 3242 643 3243 647
rect 3247 646 3248 647
rect 3383 647 3389 648
rect 3383 646 3384 647
rect 3247 644 3384 646
rect 3247 643 3248 644
rect 3242 642 3248 643
rect 3383 643 3384 644
rect 3388 643 3389 647
rect 3383 642 3389 643
rect 3394 647 3400 648
rect 3394 643 3395 647
rect 3399 646 3400 647
rect 3639 647 3645 648
rect 3639 646 3640 647
rect 3399 644 3640 646
rect 3399 643 3400 644
rect 3394 642 3400 643
rect 3639 643 3640 644
rect 3644 643 3645 647
rect 3639 642 3645 643
rect 3903 647 3909 648
rect 3903 643 3904 647
rect 3908 646 3909 647
rect 3914 647 3920 648
rect 3914 646 3915 647
rect 3908 644 3915 646
rect 3908 643 3909 644
rect 3903 642 3909 643
rect 3914 643 3915 644
rect 3919 643 3920 647
rect 3914 642 3920 643
rect 3402 639 3408 640
rect 3402 638 3403 639
rect 3236 636 3403 638
rect 3402 635 3403 636
rect 3407 635 3408 639
rect 3402 634 3408 635
rect 110 632 116 633
rect 2006 632 2012 633
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 294 631 300 632
rect 294 627 295 631
rect 299 627 300 631
rect 294 626 300 627
rect 446 631 452 632
rect 446 627 447 631
rect 451 627 452 631
rect 446 626 452 627
rect 614 631 620 632
rect 614 627 615 631
rect 619 627 620 631
rect 614 626 620 627
rect 782 631 788 632
rect 782 627 783 631
rect 787 627 788 631
rect 782 626 788 627
rect 950 631 956 632
rect 950 627 951 631
rect 955 627 956 631
rect 950 626 956 627
rect 1110 631 1116 632
rect 1110 627 1111 631
rect 1115 627 1116 631
rect 1110 626 1116 627
rect 1262 631 1268 632
rect 1262 627 1263 631
rect 1267 627 1268 631
rect 1262 626 1268 627
rect 1398 631 1404 632
rect 1398 627 1399 631
rect 1403 627 1404 631
rect 1398 626 1404 627
rect 1534 631 1540 632
rect 1534 627 1535 631
rect 1539 627 1540 631
rect 1534 626 1540 627
rect 1662 631 1668 632
rect 1662 627 1663 631
rect 1667 627 1668 631
rect 1662 626 1668 627
rect 1790 631 1796 632
rect 1790 627 1791 631
rect 1795 627 1796 631
rect 1790 626 1796 627
rect 1902 631 1908 632
rect 1902 627 1903 631
rect 1907 627 1908 631
rect 2006 628 2007 632
rect 2011 628 2012 632
rect 2006 627 2012 628
rect 2046 628 2052 629
rect 3942 628 3948 629
rect 1902 626 1908 627
rect 2046 624 2047 628
rect 2051 624 2052 628
rect 370 623 376 624
rect 370 619 371 623
rect 375 619 376 623
rect 370 618 376 619
rect 522 623 528 624
rect 522 619 523 623
rect 527 619 528 623
rect 698 623 704 624
rect 522 618 528 619
rect 690 619 696 620
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 690 615 691 619
rect 695 615 696 619
rect 698 619 699 623
rect 703 622 704 623
rect 866 623 872 624
rect 703 620 825 622
rect 703 619 704 620
rect 698 618 704 619
rect 866 619 867 623
rect 871 622 872 623
rect 1186 623 1192 624
rect 871 620 993 622
rect 871 619 872 620
rect 866 618 872 619
rect 1186 619 1187 623
rect 1191 619 1192 623
rect 1186 618 1192 619
rect 1338 623 1344 624
rect 1338 619 1339 623
rect 1343 619 1344 623
rect 1338 618 1344 619
rect 1474 623 1480 624
rect 1474 619 1475 623
rect 1479 619 1480 623
rect 1474 618 1480 619
rect 1482 623 1488 624
rect 1482 619 1483 623
rect 1487 622 1488 623
rect 1618 623 1624 624
rect 1487 620 1577 622
rect 1487 619 1488 620
rect 1482 618 1488 619
rect 1618 619 1619 623
rect 1623 622 1624 623
rect 1866 623 1872 624
rect 1623 620 1705 622
rect 1623 619 1624 620
rect 1618 618 1624 619
rect 1866 619 1867 623
rect 1871 619 1872 623
rect 1866 618 1872 619
rect 1978 623 1984 624
rect 2046 623 2052 624
rect 2070 627 2076 628
rect 2070 623 2071 627
rect 2075 623 2076 627
rect 1978 619 1979 623
rect 1983 619 1984 623
rect 2070 622 2076 623
rect 2238 627 2244 628
rect 2238 623 2239 627
rect 2243 623 2244 627
rect 2238 622 2244 623
rect 2422 627 2428 628
rect 2422 623 2423 627
rect 2427 623 2428 627
rect 2422 622 2428 623
rect 2622 627 2628 628
rect 2622 623 2623 627
rect 2627 623 2628 627
rect 2622 622 2628 623
rect 2838 627 2844 628
rect 2838 623 2839 627
rect 2843 623 2844 627
rect 2838 622 2844 623
rect 3070 627 3076 628
rect 3070 623 3071 627
rect 3075 623 3076 627
rect 3070 622 3076 623
rect 3318 627 3324 628
rect 3318 623 3319 627
rect 3323 623 3324 627
rect 3318 622 3324 623
rect 3574 627 3580 628
rect 3574 623 3575 627
rect 3579 623 3580 627
rect 3574 622 3580 623
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3942 624 3943 628
rect 3947 624 3948 628
rect 3942 623 3948 624
rect 3838 622 3844 623
rect 1978 618 1984 619
rect 2146 619 2152 620
rect 690 614 696 615
rect 2006 615 2012 616
rect 110 610 116 611
rect 294 612 300 613
rect 294 608 295 612
rect 299 608 300 612
rect 294 607 300 608
rect 446 612 452 613
rect 446 608 447 612
rect 451 608 452 612
rect 446 607 452 608
rect 614 612 620 613
rect 614 608 615 612
rect 619 608 620 612
rect 614 607 620 608
rect 782 612 788 613
rect 782 608 783 612
rect 787 608 788 612
rect 782 607 788 608
rect 950 612 956 613
rect 950 608 951 612
rect 955 608 956 612
rect 950 607 956 608
rect 1110 612 1116 613
rect 1110 608 1111 612
rect 1115 608 1116 612
rect 1110 607 1116 608
rect 1262 612 1268 613
rect 1262 608 1263 612
rect 1267 608 1268 612
rect 1262 607 1268 608
rect 1398 612 1404 613
rect 1398 608 1399 612
rect 1403 608 1404 612
rect 1398 607 1404 608
rect 1534 612 1540 613
rect 1534 608 1535 612
rect 1539 608 1540 612
rect 1534 607 1540 608
rect 1662 612 1668 613
rect 1662 608 1663 612
rect 1667 608 1668 612
rect 1662 607 1668 608
rect 1790 612 1796 613
rect 1790 608 1791 612
rect 1795 608 1796 612
rect 1790 607 1796 608
rect 1902 612 1908 613
rect 1902 608 1903 612
rect 1907 608 1908 612
rect 2006 611 2007 615
rect 2011 611 2012 615
rect 2146 615 2147 619
rect 2151 615 2152 619
rect 2146 614 2152 615
rect 2314 619 2320 620
rect 2314 615 2315 619
rect 2319 615 2320 619
rect 2314 614 2320 615
rect 2322 619 2328 620
rect 2322 615 2323 619
rect 2327 618 2328 619
rect 2762 619 2768 620
rect 2327 616 2465 618
rect 2327 615 2328 616
rect 2322 614 2328 615
rect 2698 615 2704 616
rect 2006 610 2012 611
rect 2046 611 2052 612
rect 1902 607 1908 608
rect 2046 607 2047 611
rect 2051 607 2052 611
rect 2698 611 2699 615
rect 2703 611 2704 615
rect 2762 615 2763 619
rect 2767 618 2768 619
rect 2922 619 2928 620
rect 2767 616 2881 618
rect 2767 615 2768 616
rect 2762 614 2768 615
rect 2922 615 2923 619
rect 2927 618 2928 619
rect 3394 619 3400 620
rect 2927 616 3113 618
rect 2927 615 2928 616
rect 2922 614 2928 615
rect 3394 615 3395 619
rect 3399 615 3400 619
rect 3394 614 3400 615
rect 3402 619 3408 620
rect 3402 615 3403 619
rect 3407 618 3408 619
rect 3407 616 3617 618
rect 3407 615 3408 616
rect 3402 614 3408 615
rect 3914 615 3920 616
rect 2698 610 2704 611
rect 3914 611 3915 615
rect 3919 611 3920 615
rect 3914 610 3920 611
rect 3942 611 3948 612
rect 2046 606 2052 607
rect 2070 608 2076 609
rect 2070 604 2071 608
rect 2075 604 2076 608
rect 2070 603 2076 604
rect 2238 608 2244 609
rect 2238 604 2239 608
rect 2243 604 2244 608
rect 2238 603 2244 604
rect 2422 608 2428 609
rect 2422 604 2423 608
rect 2427 604 2428 608
rect 2422 603 2428 604
rect 2622 608 2628 609
rect 2622 604 2623 608
rect 2627 604 2628 608
rect 2622 603 2628 604
rect 2838 608 2844 609
rect 2838 604 2839 608
rect 2843 604 2844 608
rect 2838 603 2844 604
rect 3070 608 3076 609
rect 3070 604 3071 608
rect 3075 604 3076 608
rect 3070 603 3076 604
rect 3318 608 3324 609
rect 3318 604 3319 608
rect 3323 604 3324 608
rect 3318 603 3324 604
rect 3574 608 3580 609
rect 3574 604 3575 608
rect 3579 604 3580 608
rect 3574 603 3580 604
rect 3838 608 3844 609
rect 3838 604 3839 608
rect 3843 604 3844 608
rect 3942 607 3943 611
rect 3947 607 3948 611
rect 3942 606 3948 607
rect 3838 603 3844 604
rect 238 548 244 549
rect 110 545 116 546
rect 110 541 111 545
rect 115 541 116 545
rect 238 544 239 548
rect 243 544 244 548
rect 238 543 244 544
rect 414 548 420 549
rect 414 544 415 548
rect 419 544 420 548
rect 414 543 420 544
rect 606 548 612 549
rect 606 544 607 548
rect 611 544 612 548
rect 606 543 612 544
rect 798 548 804 549
rect 798 544 799 548
rect 803 544 804 548
rect 798 543 804 544
rect 990 548 996 549
rect 990 544 991 548
rect 995 544 996 548
rect 990 543 996 544
rect 1174 548 1180 549
rect 1174 544 1175 548
rect 1179 544 1180 548
rect 1174 543 1180 544
rect 1350 548 1356 549
rect 1350 544 1351 548
rect 1355 544 1356 548
rect 1350 543 1356 544
rect 1518 548 1524 549
rect 1518 544 1519 548
rect 1523 544 1524 548
rect 1518 543 1524 544
rect 1686 548 1692 549
rect 1686 544 1687 548
rect 1691 544 1692 548
rect 1686 543 1692 544
rect 1862 548 1868 549
rect 1862 544 1863 548
rect 1867 544 1868 548
rect 2190 548 2196 549
rect 1862 543 1868 544
rect 2006 545 2012 546
rect 110 540 116 541
rect 2006 541 2007 545
rect 2011 541 2012 545
rect 2006 540 2012 541
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2190 544 2191 548
rect 2195 544 2196 548
rect 2190 543 2196 544
rect 2286 548 2292 549
rect 2286 544 2287 548
rect 2291 544 2292 548
rect 2286 543 2292 544
rect 2382 548 2388 549
rect 2382 544 2383 548
rect 2387 544 2388 548
rect 2382 543 2388 544
rect 2478 548 2484 549
rect 2478 544 2479 548
rect 2483 544 2484 548
rect 2478 543 2484 544
rect 2582 548 2588 549
rect 2582 544 2583 548
rect 2587 544 2588 548
rect 2582 543 2588 544
rect 2710 548 2716 549
rect 2710 544 2711 548
rect 2715 544 2716 548
rect 2710 543 2716 544
rect 2870 548 2876 549
rect 2870 544 2871 548
rect 2875 544 2876 548
rect 2870 543 2876 544
rect 3070 548 3076 549
rect 3070 544 3071 548
rect 3075 544 3076 548
rect 3070 543 3076 544
rect 3302 548 3308 549
rect 3302 544 3303 548
rect 3307 544 3308 548
rect 3302 543 3308 544
rect 3550 548 3556 549
rect 3550 544 3551 548
rect 3555 544 3556 548
rect 3550 543 3556 544
rect 3806 548 3812 549
rect 3806 544 3807 548
rect 3811 544 3812 548
rect 3806 543 3812 544
rect 3942 545 3948 546
rect 2046 540 2052 541
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 314 539 320 540
rect 314 535 315 539
rect 319 535 320 539
rect 314 534 320 535
rect 370 539 376 540
rect 370 535 371 539
rect 375 538 376 539
rect 754 539 760 540
rect 754 538 755 539
rect 375 536 457 538
rect 685 536 755 538
rect 375 535 376 536
rect 370 534 376 535
rect 754 535 755 536
rect 759 535 760 539
rect 754 534 760 535
rect 874 539 880 540
rect 874 535 875 539
rect 879 535 880 539
rect 874 534 880 535
rect 882 539 888 540
rect 882 535 883 539
rect 887 538 888 539
rect 1250 539 1256 540
rect 887 536 1033 538
rect 887 535 888 536
rect 882 534 888 535
rect 1250 535 1251 539
rect 1255 535 1256 539
rect 1250 534 1256 535
rect 1426 539 1432 540
rect 1426 535 1427 539
rect 1431 535 1432 539
rect 1426 534 1432 535
rect 1594 539 1600 540
rect 1594 535 1595 539
rect 1599 535 1600 539
rect 1594 534 1600 535
rect 1762 539 1768 540
rect 1762 535 1763 539
rect 1767 535 1768 539
rect 1762 534 1768 535
rect 1818 539 1824 540
rect 1818 535 1819 539
rect 1823 538 1824 539
rect 2266 539 2272 540
rect 1823 536 1905 538
rect 1823 535 1824 536
rect 1818 534 1824 535
rect 2266 535 2267 539
rect 2271 535 2272 539
rect 2266 534 2272 535
rect 2362 539 2368 540
rect 2362 535 2363 539
rect 2367 535 2368 539
rect 2362 534 2368 535
rect 2458 539 2464 540
rect 2458 535 2459 539
rect 2463 535 2464 539
rect 2458 534 2464 535
rect 2554 539 2560 540
rect 2554 535 2555 539
rect 2559 535 2560 539
rect 2554 534 2560 535
rect 2562 539 2568 540
rect 2562 535 2563 539
rect 2567 538 2568 539
rect 2786 539 2792 540
rect 2567 536 2625 538
rect 2567 535 2568 536
rect 2562 534 2568 535
rect 2786 535 2787 539
rect 2791 535 2792 539
rect 2786 534 2792 535
rect 2946 539 2952 540
rect 2946 535 2947 539
rect 2951 535 2952 539
rect 2946 534 2952 535
rect 3146 539 3152 540
rect 3146 535 3147 539
rect 3151 535 3152 539
rect 3478 539 3484 540
rect 3478 538 3479 539
rect 3381 536 3479 538
rect 3146 534 3152 535
rect 3478 535 3479 536
rect 3483 535 3484 539
rect 3478 534 3484 535
rect 3626 539 3632 540
rect 3626 535 3627 539
rect 3631 535 3632 539
rect 3626 534 3632 535
rect 3874 539 3880 540
rect 3874 535 3875 539
rect 3879 535 3880 539
rect 3874 534 3880 535
rect 238 529 244 530
rect 110 528 116 529
rect 110 524 111 528
rect 115 524 116 528
rect 238 525 239 529
rect 243 525 244 529
rect 238 524 244 525
rect 414 529 420 530
rect 414 525 415 529
rect 419 525 420 529
rect 414 524 420 525
rect 606 529 612 530
rect 606 525 607 529
rect 611 525 612 529
rect 606 524 612 525
rect 798 529 804 530
rect 798 525 799 529
rect 803 525 804 529
rect 798 524 804 525
rect 990 529 996 530
rect 990 525 991 529
rect 995 525 996 529
rect 990 524 996 525
rect 1174 529 1180 530
rect 1174 525 1175 529
rect 1179 525 1180 529
rect 1174 524 1180 525
rect 1350 529 1356 530
rect 1350 525 1351 529
rect 1355 525 1356 529
rect 1350 524 1356 525
rect 1518 529 1524 530
rect 1518 525 1519 529
rect 1523 525 1524 529
rect 1518 524 1524 525
rect 1686 529 1692 530
rect 1686 525 1687 529
rect 1691 525 1692 529
rect 1686 524 1692 525
rect 1862 529 1868 530
rect 2190 529 2196 530
rect 1862 525 1863 529
rect 1867 525 1868 529
rect 1862 524 1868 525
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 110 523 116 524
rect 2006 523 2012 524
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2190 525 2191 529
rect 2195 525 2196 529
rect 2190 524 2196 525
rect 2286 529 2292 530
rect 2286 525 2287 529
rect 2291 525 2292 529
rect 2286 524 2292 525
rect 2382 529 2388 530
rect 2382 525 2383 529
rect 2387 525 2388 529
rect 2382 524 2388 525
rect 2478 529 2484 530
rect 2478 525 2479 529
rect 2483 525 2484 529
rect 2478 524 2484 525
rect 2582 529 2588 530
rect 2582 525 2583 529
rect 2587 525 2588 529
rect 2582 524 2588 525
rect 2710 529 2716 530
rect 2710 525 2711 529
rect 2715 525 2716 529
rect 2710 524 2716 525
rect 2870 529 2876 530
rect 2870 525 2871 529
rect 2875 525 2876 529
rect 2870 524 2876 525
rect 3070 529 3076 530
rect 3070 525 3071 529
rect 3075 525 3076 529
rect 3070 524 3076 525
rect 3302 529 3308 530
rect 3302 525 3303 529
rect 3307 525 3308 529
rect 3302 524 3308 525
rect 3550 529 3556 530
rect 3550 525 3551 529
rect 3555 525 3556 529
rect 3550 524 3556 525
rect 3806 529 3812 530
rect 3806 525 3807 529
rect 3811 525 3812 529
rect 3806 524 3812 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 3942 523 3948 524
rect 1519 515 1525 516
rect 1519 514 1520 515
rect 1244 512 1520 514
rect 1244 508 1246 512
rect 1519 511 1520 512
rect 1524 511 1525 515
rect 2322 515 2328 516
rect 2322 514 2323 515
rect 1519 510 1525 511
rect 2260 512 2323 514
rect 2260 508 2262 512
rect 2322 511 2323 512
rect 2327 511 2328 515
rect 2322 510 2328 511
rect 303 507 309 508
rect 303 503 304 507
rect 308 506 309 507
rect 370 507 376 508
rect 370 506 371 507
rect 308 504 371 506
rect 308 503 309 504
rect 303 502 309 503
rect 370 503 371 504
rect 375 503 376 507
rect 370 502 376 503
rect 479 507 485 508
rect 479 503 480 507
rect 484 506 485 507
rect 538 507 544 508
rect 538 506 539 507
rect 484 504 539 506
rect 484 503 485 504
rect 479 502 485 503
rect 538 503 539 504
rect 543 503 544 507
rect 538 502 544 503
rect 671 507 677 508
rect 671 503 672 507
rect 676 506 677 507
rect 690 507 696 508
rect 690 506 691 507
rect 676 504 691 506
rect 676 503 677 504
rect 671 502 677 503
rect 690 503 691 504
rect 695 503 696 507
rect 690 502 696 503
rect 754 507 760 508
rect 754 503 755 507
rect 759 506 760 507
rect 863 507 869 508
rect 863 506 864 507
rect 759 504 864 506
rect 759 503 760 504
rect 754 502 760 503
rect 863 503 864 504
rect 868 503 869 507
rect 863 502 869 503
rect 874 507 880 508
rect 874 503 875 507
rect 879 506 880 507
rect 1055 507 1061 508
rect 1055 506 1056 507
rect 879 504 1056 506
rect 879 503 880 504
rect 874 502 880 503
rect 1055 503 1056 504
rect 1060 503 1061 507
rect 1055 502 1061 503
rect 1239 507 1246 508
rect 1239 503 1240 507
rect 1244 504 1246 507
rect 1250 507 1256 508
rect 1244 503 1245 504
rect 1239 502 1245 503
rect 1250 503 1251 507
rect 1255 506 1256 507
rect 1415 507 1421 508
rect 1415 506 1416 507
rect 1255 504 1416 506
rect 1255 503 1256 504
rect 1250 502 1256 503
rect 1415 503 1416 504
rect 1420 503 1421 507
rect 1415 502 1421 503
rect 1426 507 1432 508
rect 1426 503 1427 507
rect 1431 506 1432 507
rect 1583 507 1589 508
rect 1583 506 1584 507
rect 1431 504 1584 506
rect 1431 503 1432 504
rect 1426 502 1432 503
rect 1583 503 1584 504
rect 1588 503 1589 507
rect 1583 502 1589 503
rect 1594 507 1600 508
rect 1594 503 1595 507
rect 1599 506 1600 507
rect 1751 507 1757 508
rect 1751 506 1752 507
rect 1599 504 1752 506
rect 1599 503 1600 504
rect 1594 502 1600 503
rect 1751 503 1752 504
rect 1756 503 1757 507
rect 1751 502 1757 503
rect 1762 507 1768 508
rect 1762 503 1763 507
rect 1767 506 1768 507
rect 1927 507 1933 508
rect 1927 506 1928 507
rect 1767 504 1928 506
rect 1767 503 1768 504
rect 1762 502 1768 503
rect 1927 503 1928 504
rect 1932 503 1933 507
rect 1927 502 1933 503
rect 2255 507 2262 508
rect 2255 503 2256 507
rect 2260 504 2262 507
rect 2266 507 2272 508
rect 2260 503 2261 504
rect 2255 502 2261 503
rect 2266 503 2267 507
rect 2271 506 2272 507
rect 2351 507 2357 508
rect 2351 506 2352 507
rect 2271 504 2352 506
rect 2271 503 2272 504
rect 2266 502 2272 503
rect 2351 503 2352 504
rect 2356 503 2357 507
rect 2351 502 2357 503
rect 2362 507 2368 508
rect 2362 503 2363 507
rect 2367 506 2368 507
rect 2447 507 2453 508
rect 2447 506 2448 507
rect 2367 504 2448 506
rect 2367 503 2368 504
rect 2362 502 2368 503
rect 2447 503 2448 504
rect 2452 503 2453 507
rect 2447 502 2453 503
rect 2458 507 2464 508
rect 2458 503 2459 507
rect 2463 506 2464 507
rect 2543 507 2549 508
rect 2543 506 2544 507
rect 2463 504 2544 506
rect 2463 503 2464 504
rect 2458 502 2464 503
rect 2543 503 2544 504
rect 2548 503 2549 507
rect 2543 502 2549 503
rect 2554 507 2560 508
rect 2554 503 2555 507
rect 2559 506 2560 507
rect 2647 507 2653 508
rect 2647 506 2648 507
rect 2559 504 2648 506
rect 2559 503 2560 504
rect 2554 502 2560 503
rect 2647 503 2648 504
rect 2652 503 2653 507
rect 2647 502 2653 503
rect 2698 507 2704 508
rect 2698 503 2699 507
rect 2703 506 2704 507
rect 2775 507 2781 508
rect 2775 506 2776 507
rect 2703 504 2776 506
rect 2703 503 2704 504
rect 2698 502 2704 503
rect 2775 503 2776 504
rect 2780 503 2781 507
rect 2775 502 2781 503
rect 2786 507 2792 508
rect 2786 503 2787 507
rect 2791 506 2792 507
rect 2935 507 2941 508
rect 2935 506 2936 507
rect 2791 504 2936 506
rect 2791 503 2792 504
rect 2786 502 2792 503
rect 2935 503 2936 504
rect 2940 503 2941 507
rect 2935 502 2941 503
rect 2946 507 2952 508
rect 2946 503 2947 507
rect 2951 506 2952 507
rect 3135 507 3141 508
rect 3135 506 3136 507
rect 2951 504 3136 506
rect 2951 503 2952 504
rect 2946 502 2952 503
rect 3135 503 3136 504
rect 3140 503 3141 507
rect 3135 502 3141 503
rect 3146 507 3152 508
rect 3146 503 3147 507
rect 3151 506 3152 507
rect 3367 507 3373 508
rect 3367 506 3368 507
rect 3151 504 3368 506
rect 3151 503 3152 504
rect 3146 502 3152 503
rect 3367 503 3368 504
rect 3372 503 3373 507
rect 3367 502 3373 503
rect 3478 507 3484 508
rect 3478 503 3479 507
rect 3483 506 3484 507
rect 3615 507 3621 508
rect 3615 506 3616 507
rect 3483 504 3616 506
rect 3483 503 3484 504
rect 3478 502 3484 503
rect 3615 503 3616 504
rect 3620 503 3621 507
rect 3615 502 3621 503
rect 3871 507 3877 508
rect 3871 503 3872 507
rect 3876 506 3877 507
rect 3914 507 3920 508
rect 3914 506 3915 507
rect 3876 504 3915 506
rect 3876 503 3877 504
rect 3871 502 3877 503
rect 3914 503 3915 504
rect 3919 503 3920 507
rect 3914 502 3920 503
rect 199 495 208 496
rect 199 491 200 495
rect 207 491 208 495
rect 199 490 208 491
rect 210 495 216 496
rect 210 491 211 495
rect 215 494 216 495
rect 351 495 357 496
rect 351 494 352 495
rect 215 492 352 494
rect 215 491 216 492
rect 210 490 216 491
rect 351 491 352 492
rect 356 491 357 495
rect 351 490 357 491
rect 362 495 368 496
rect 362 491 363 495
rect 367 494 368 495
rect 527 495 533 496
rect 527 494 528 495
rect 367 492 528 494
rect 367 491 368 492
rect 362 490 368 491
rect 527 491 528 492
rect 532 491 533 495
rect 527 490 533 491
rect 703 495 709 496
rect 703 491 704 495
rect 708 494 709 495
rect 727 495 733 496
rect 727 494 728 495
rect 708 492 728 494
rect 708 491 709 492
rect 703 490 709 491
rect 727 491 728 492
rect 732 491 733 495
rect 727 490 733 491
rect 871 495 877 496
rect 871 491 872 495
rect 876 494 877 495
rect 882 495 888 496
rect 882 494 883 495
rect 876 492 883 494
rect 876 491 877 492
rect 871 490 877 491
rect 882 491 883 492
rect 887 491 888 495
rect 882 490 888 491
rect 1031 495 1037 496
rect 1031 491 1032 495
rect 1036 494 1037 495
rect 1102 495 1108 496
rect 1036 492 1098 494
rect 1036 491 1037 492
rect 1031 490 1037 491
rect 1096 486 1098 492
rect 1102 491 1103 495
rect 1107 494 1108 495
rect 1183 495 1189 496
rect 1183 494 1184 495
rect 1107 492 1184 494
rect 1107 491 1108 492
rect 1102 490 1108 491
rect 1183 491 1184 492
rect 1188 491 1189 495
rect 1183 490 1189 491
rect 1194 495 1200 496
rect 1194 491 1195 495
rect 1199 494 1200 495
rect 1335 495 1341 496
rect 1335 494 1336 495
rect 1199 492 1336 494
rect 1199 491 1200 492
rect 1194 490 1200 491
rect 1335 491 1336 492
rect 1340 491 1341 495
rect 1335 490 1341 491
rect 1394 495 1400 496
rect 1394 491 1395 495
rect 1399 494 1400 495
rect 1479 495 1485 496
rect 1479 494 1480 495
rect 1399 492 1480 494
rect 1399 491 1400 492
rect 1394 490 1400 491
rect 1479 491 1480 492
rect 1484 491 1485 495
rect 1479 490 1485 491
rect 1490 495 1496 496
rect 1490 491 1491 495
rect 1495 494 1496 495
rect 1631 495 1637 496
rect 1631 494 1632 495
rect 1495 492 1632 494
rect 1495 491 1496 492
rect 1490 490 1496 491
rect 1631 491 1632 492
rect 1636 491 1637 495
rect 1631 490 1637 491
rect 2495 495 2501 496
rect 2495 491 2496 495
rect 2500 491 2501 495
rect 2495 490 2501 491
rect 2506 495 2512 496
rect 2506 491 2507 495
rect 2511 494 2512 495
rect 2591 495 2597 496
rect 2591 494 2592 495
rect 2511 492 2592 494
rect 2511 491 2512 492
rect 2506 490 2512 491
rect 2591 491 2592 492
rect 2596 491 2597 495
rect 2591 490 2597 491
rect 2602 495 2608 496
rect 2602 491 2603 495
rect 2607 494 2608 495
rect 2687 495 2693 496
rect 2687 494 2688 495
rect 2607 492 2688 494
rect 2607 491 2608 492
rect 2602 490 2608 491
rect 2687 491 2688 492
rect 2692 491 2693 495
rect 2687 490 2693 491
rect 2698 495 2704 496
rect 2698 491 2699 495
rect 2703 494 2704 495
rect 2791 495 2797 496
rect 2791 494 2792 495
rect 2703 492 2792 494
rect 2703 491 2704 492
rect 2698 490 2704 491
rect 2791 491 2792 492
rect 2796 491 2797 495
rect 2791 490 2797 491
rect 2802 495 2808 496
rect 2802 491 2803 495
rect 2807 494 2808 495
rect 2911 495 2917 496
rect 2911 494 2912 495
rect 2807 492 2912 494
rect 2807 491 2808 492
rect 2802 490 2808 491
rect 2911 491 2912 492
rect 2916 491 2917 495
rect 2911 490 2917 491
rect 2922 495 2928 496
rect 2922 491 2923 495
rect 2927 494 2928 495
rect 3063 495 3069 496
rect 3063 494 3064 495
rect 2927 492 3064 494
rect 2927 491 2928 492
rect 2922 490 2928 491
rect 3063 491 3064 492
rect 3068 491 3069 495
rect 3063 490 3069 491
rect 3239 495 3245 496
rect 3239 491 3240 495
rect 3244 494 3245 495
rect 3258 495 3264 496
rect 3258 494 3259 495
rect 3244 492 3259 494
rect 3244 491 3245 492
rect 3239 490 3245 491
rect 3258 491 3259 492
rect 3263 491 3264 495
rect 3258 490 3264 491
rect 3439 495 3445 496
rect 3439 491 3440 495
rect 3444 494 3445 495
rect 3458 495 3464 496
rect 3458 494 3459 495
rect 3444 492 3459 494
rect 3444 491 3445 492
rect 3439 490 3445 491
rect 3458 491 3459 492
rect 3463 491 3464 495
rect 3458 490 3464 491
rect 3626 495 3632 496
rect 3626 491 3627 495
rect 3631 494 3632 495
rect 3655 495 3661 496
rect 3655 494 3656 495
rect 3631 492 3656 494
rect 3631 491 3632 492
rect 3626 490 3632 491
rect 3655 491 3656 492
rect 3660 491 3661 495
rect 3655 490 3661 491
rect 3858 495 3864 496
rect 3858 491 3859 495
rect 3863 494 3864 495
rect 3871 495 3877 496
rect 3871 494 3872 495
rect 3863 492 3872 494
rect 3863 491 3864 492
rect 3858 490 3864 491
rect 3871 491 3872 492
rect 3876 491 3877 495
rect 3871 490 3877 491
rect 1290 487 1296 488
rect 1290 486 1291 487
rect 1096 484 1291 486
rect 1290 483 1291 484
rect 1295 483 1296 487
rect 2497 486 2499 490
rect 2562 487 2568 488
rect 2562 486 2563 487
rect 2497 484 2563 486
rect 1290 482 1296 483
rect 2562 483 2563 484
rect 2567 483 2568 487
rect 2562 482 2568 483
rect 110 476 116 477
rect 2006 476 2012 477
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 134 475 140 476
rect 134 471 135 475
rect 139 471 140 475
rect 134 470 140 471
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 462 475 468 476
rect 462 471 463 475
rect 467 471 468 475
rect 462 470 468 471
rect 638 475 644 476
rect 638 471 639 475
rect 643 471 644 475
rect 638 470 644 471
rect 806 475 812 476
rect 806 471 807 475
rect 811 471 812 475
rect 806 470 812 471
rect 966 475 972 476
rect 966 471 967 475
rect 971 471 972 475
rect 966 470 972 471
rect 1118 475 1124 476
rect 1118 471 1119 475
rect 1123 471 1124 475
rect 1118 470 1124 471
rect 1270 475 1276 476
rect 1270 471 1271 475
rect 1275 471 1276 475
rect 1270 470 1276 471
rect 1414 475 1420 476
rect 1414 471 1415 475
rect 1419 471 1420 475
rect 1414 470 1420 471
rect 1566 475 1572 476
rect 1566 471 1567 475
rect 1571 471 1572 475
rect 2006 472 2007 476
rect 2011 472 2012 476
rect 2006 471 2012 472
rect 2046 476 2052 477
rect 3942 476 3948 477
rect 2046 472 2047 476
rect 2051 472 2052 476
rect 2046 471 2052 472
rect 2430 475 2436 476
rect 2430 471 2431 475
rect 2435 471 2436 475
rect 1566 470 1572 471
rect 2430 470 2436 471
rect 2526 475 2532 476
rect 2526 471 2527 475
rect 2531 471 2532 475
rect 2526 470 2532 471
rect 2622 475 2628 476
rect 2622 471 2623 475
rect 2627 471 2628 475
rect 2622 470 2628 471
rect 2726 475 2732 476
rect 2726 471 2727 475
rect 2731 471 2732 475
rect 2726 470 2732 471
rect 2846 475 2852 476
rect 2846 471 2847 475
rect 2851 471 2852 475
rect 2846 470 2852 471
rect 2998 475 3004 476
rect 2998 471 2999 475
rect 3003 471 3004 475
rect 2998 470 3004 471
rect 3174 475 3180 476
rect 3174 471 3175 475
rect 3179 471 3180 475
rect 3174 470 3180 471
rect 3374 475 3380 476
rect 3374 471 3375 475
rect 3379 471 3380 475
rect 3374 470 3380 471
rect 3590 475 3596 476
rect 3590 471 3591 475
rect 3595 471 3596 475
rect 3590 470 3596 471
rect 3806 475 3812 476
rect 3806 471 3807 475
rect 3811 471 3812 475
rect 3942 472 3943 476
rect 3947 472 3948 476
rect 3942 471 3948 472
rect 3806 470 3812 471
rect 210 467 216 468
rect 210 463 211 467
rect 215 463 216 467
rect 210 462 216 463
rect 362 467 368 468
rect 362 463 363 467
rect 367 463 368 467
rect 362 462 368 463
rect 538 467 544 468
rect 538 463 539 467
rect 543 463 544 467
rect 538 462 544 463
rect 546 467 552 468
rect 546 463 547 467
rect 551 466 552 467
rect 727 467 733 468
rect 551 464 681 466
rect 551 463 552 464
rect 546 462 552 463
rect 727 463 728 467
rect 732 466 733 467
rect 1102 467 1108 468
rect 1102 466 1103 467
rect 732 464 849 466
rect 1045 464 1103 466
rect 732 463 733 464
rect 727 462 733 463
rect 1102 463 1103 464
rect 1107 463 1108 467
rect 1102 462 1108 463
rect 1194 467 1200 468
rect 1194 463 1195 467
rect 1199 463 1200 467
rect 1394 467 1400 468
rect 1394 466 1395 467
rect 1349 464 1395 466
rect 1194 462 1200 463
rect 1394 463 1395 464
rect 1399 463 1400 467
rect 1394 462 1400 463
rect 1490 467 1496 468
rect 1490 463 1491 467
rect 1495 463 1496 467
rect 1490 462 1496 463
rect 1519 467 1525 468
rect 1519 463 1520 467
rect 1524 466 1525 467
rect 2506 467 2512 468
rect 1524 464 1609 466
rect 1524 463 1525 464
rect 1519 462 1525 463
rect 2506 463 2507 467
rect 2511 463 2512 467
rect 2506 462 2512 463
rect 2602 467 2608 468
rect 2602 463 2603 467
rect 2607 463 2608 467
rect 2602 462 2608 463
rect 2698 467 2704 468
rect 2698 463 2699 467
rect 2703 463 2704 467
rect 2698 462 2704 463
rect 2802 467 2808 468
rect 2802 463 2803 467
rect 2807 463 2808 467
rect 2802 462 2808 463
rect 2922 467 2928 468
rect 2922 463 2923 467
rect 2927 463 2928 467
rect 2922 462 2928 463
rect 2934 467 2940 468
rect 2934 463 2935 467
rect 2939 466 2940 467
rect 3082 467 3088 468
rect 2939 464 3041 466
rect 2939 463 2940 464
rect 2934 462 2940 463
rect 3082 463 3083 467
rect 3087 466 3088 467
rect 3258 467 3264 468
rect 3087 464 3217 466
rect 3087 463 3088 464
rect 3082 462 3088 463
rect 3258 463 3259 467
rect 3263 466 3264 467
rect 3458 467 3464 468
rect 3263 464 3417 466
rect 3263 463 3264 464
rect 3258 462 3264 463
rect 3458 463 3459 467
rect 3463 466 3464 467
rect 3463 464 3633 466
rect 3463 463 3464 464
rect 3458 462 3464 463
rect 3882 463 3888 464
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 2006 459 2012 460
rect 110 454 116 455
rect 134 456 140 457
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 286 456 292 457
rect 286 452 287 456
rect 291 452 292 456
rect 286 451 292 452
rect 462 456 468 457
rect 462 452 463 456
rect 467 452 468 456
rect 462 451 468 452
rect 638 456 644 457
rect 638 452 639 456
rect 643 452 644 456
rect 638 451 644 452
rect 806 456 812 457
rect 806 452 807 456
rect 811 452 812 456
rect 806 451 812 452
rect 966 456 972 457
rect 966 452 967 456
rect 971 452 972 456
rect 966 451 972 452
rect 1118 456 1124 457
rect 1118 452 1119 456
rect 1123 452 1124 456
rect 1118 451 1124 452
rect 1270 456 1276 457
rect 1270 452 1271 456
rect 1275 452 1276 456
rect 1270 451 1276 452
rect 1414 456 1420 457
rect 1414 452 1415 456
rect 1419 452 1420 456
rect 1414 451 1420 452
rect 1566 456 1572 457
rect 1566 452 1567 456
rect 1571 452 1572 456
rect 2006 455 2007 459
rect 2011 455 2012 459
rect 2006 454 2012 455
rect 2046 459 2052 460
rect 2046 455 2047 459
rect 2051 455 2052 459
rect 3882 459 3883 463
rect 3887 459 3888 463
rect 3882 458 3888 459
rect 3942 459 3948 460
rect 2046 454 2052 455
rect 2430 456 2436 457
rect 1566 451 1572 452
rect 2430 452 2431 456
rect 2435 452 2436 456
rect 2430 451 2436 452
rect 2526 456 2532 457
rect 2526 452 2527 456
rect 2531 452 2532 456
rect 2526 451 2532 452
rect 2622 456 2628 457
rect 2622 452 2623 456
rect 2627 452 2628 456
rect 2622 451 2628 452
rect 2726 456 2732 457
rect 2726 452 2727 456
rect 2731 452 2732 456
rect 2726 451 2732 452
rect 2846 456 2852 457
rect 2846 452 2847 456
rect 2851 452 2852 456
rect 2846 451 2852 452
rect 2998 456 3004 457
rect 2998 452 2999 456
rect 3003 452 3004 456
rect 2998 451 3004 452
rect 3174 456 3180 457
rect 3174 452 3175 456
rect 3179 452 3180 456
rect 3174 451 3180 452
rect 3374 456 3380 457
rect 3374 452 3375 456
rect 3379 452 3380 456
rect 3374 451 3380 452
rect 3590 456 3596 457
rect 3590 452 3591 456
rect 3595 452 3596 456
rect 3590 451 3596 452
rect 3806 456 3812 457
rect 3806 452 3807 456
rect 3811 452 3812 456
rect 3942 455 3943 459
rect 3947 455 3948 459
rect 3942 454 3948 455
rect 3806 451 3812 452
rect 2430 396 2436 397
rect 2046 393 2052 394
rect 134 392 140 393
rect 110 389 116 390
rect 110 385 111 389
rect 115 385 116 389
rect 134 388 135 392
rect 139 388 140 392
rect 134 387 140 388
rect 278 392 284 393
rect 278 388 279 392
rect 283 388 284 392
rect 278 387 284 388
rect 438 392 444 393
rect 438 388 439 392
rect 443 388 444 392
rect 438 387 444 388
rect 582 392 588 393
rect 582 388 583 392
rect 587 388 588 392
rect 582 387 588 388
rect 718 392 724 393
rect 718 388 719 392
rect 723 388 724 392
rect 718 387 724 388
rect 846 392 852 393
rect 846 388 847 392
rect 851 388 852 392
rect 846 387 852 388
rect 966 392 972 393
rect 966 388 967 392
rect 971 388 972 392
rect 966 387 972 388
rect 1086 392 1092 393
rect 1086 388 1087 392
rect 1091 388 1092 392
rect 1086 387 1092 388
rect 1206 392 1212 393
rect 1206 388 1207 392
rect 1211 388 1212 392
rect 1206 387 1212 388
rect 1326 392 1332 393
rect 1326 388 1327 392
rect 1331 388 1332 392
rect 1326 387 1332 388
rect 2006 389 2012 390
rect 110 384 116 385
rect 2006 385 2007 389
rect 2011 385 2012 389
rect 2046 389 2047 393
rect 2051 389 2052 393
rect 2430 392 2431 396
rect 2435 392 2436 396
rect 2430 391 2436 392
rect 2526 396 2532 397
rect 2526 392 2527 396
rect 2531 392 2532 396
rect 2526 391 2532 392
rect 2622 396 2628 397
rect 2622 392 2623 396
rect 2627 392 2628 396
rect 2622 391 2628 392
rect 2718 396 2724 397
rect 2718 392 2719 396
rect 2723 392 2724 396
rect 2718 391 2724 392
rect 2814 396 2820 397
rect 2814 392 2815 396
rect 2819 392 2820 396
rect 2814 391 2820 392
rect 2926 396 2932 397
rect 2926 392 2927 396
rect 2931 392 2932 396
rect 2926 391 2932 392
rect 3062 396 3068 397
rect 3062 392 3063 396
rect 3067 392 3068 396
rect 3062 391 3068 392
rect 3222 396 3228 397
rect 3222 392 3223 396
rect 3227 392 3228 396
rect 3222 391 3228 392
rect 3398 396 3404 397
rect 3398 392 3399 396
rect 3403 392 3404 396
rect 3398 391 3404 392
rect 3590 396 3596 397
rect 3590 392 3591 396
rect 3595 392 3596 396
rect 3590 391 3596 392
rect 3782 396 3788 397
rect 3782 392 3783 396
rect 3787 392 3788 396
rect 3782 391 3788 392
rect 3942 393 3948 394
rect 2046 388 2052 389
rect 3942 389 3943 393
rect 3947 389 3948 393
rect 3942 388 3948 389
rect 2006 384 2012 385
rect 2506 387 2512 388
rect 202 383 208 384
rect 202 379 203 383
rect 207 379 208 383
rect 514 383 520 384
rect 202 378 208 379
rect 260 380 321 382
rect 202 375 208 376
rect 134 373 140 374
rect 110 372 116 373
rect 110 368 111 372
rect 115 368 116 372
rect 134 369 135 373
rect 139 369 140 373
rect 202 371 203 375
rect 207 374 208 375
rect 260 374 262 380
rect 514 379 515 383
rect 519 379 520 383
rect 514 378 520 379
rect 658 383 664 384
rect 658 379 659 383
rect 663 379 664 383
rect 658 378 664 379
rect 794 383 800 384
rect 794 379 795 383
rect 799 379 800 383
rect 794 378 800 379
rect 922 383 928 384
rect 922 379 923 383
rect 927 379 928 383
rect 922 378 928 379
rect 1042 383 1048 384
rect 1042 379 1043 383
rect 1047 379 1048 383
rect 1042 378 1048 379
rect 1162 383 1168 384
rect 1162 379 1163 383
rect 1167 379 1168 383
rect 1162 378 1168 379
rect 1282 383 1288 384
rect 1282 379 1283 383
rect 1287 379 1288 383
rect 1282 378 1288 379
rect 1290 383 1296 384
rect 1290 379 1291 383
rect 1295 382 1296 383
rect 2506 383 2507 387
rect 2511 383 2512 387
rect 2506 382 2512 383
rect 2602 387 2608 388
rect 2602 383 2603 387
rect 2607 383 2608 387
rect 2602 382 2608 383
rect 2610 387 2616 388
rect 2610 383 2611 387
rect 2615 386 2616 387
rect 2706 387 2712 388
rect 2615 384 2665 386
rect 2615 383 2616 384
rect 2610 382 2616 383
rect 2706 383 2707 387
rect 2711 386 2712 387
rect 2802 387 2808 388
rect 2711 384 2761 386
rect 2711 383 2712 384
rect 2706 382 2712 383
rect 2802 383 2803 387
rect 2807 386 2808 387
rect 3002 387 3008 388
rect 2807 384 2857 386
rect 2807 383 2808 384
rect 2802 382 2808 383
rect 3002 383 3003 387
rect 3007 383 3008 387
rect 3002 382 3008 383
rect 3138 387 3144 388
rect 3138 383 3139 387
rect 3143 383 3144 387
rect 3138 382 3144 383
rect 3298 387 3304 388
rect 3298 383 3299 387
rect 3303 383 3304 387
rect 3298 382 3304 383
rect 3474 387 3480 388
rect 3474 383 3475 387
rect 3479 383 3480 387
rect 3474 382 3480 383
rect 3498 387 3504 388
rect 3498 383 3499 387
rect 3503 386 3504 387
rect 3858 387 3864 388
rect 3503 384 3633 386
rect 3503 383 3504 384
rect 3498 382 3504 383
rect 3858 383 3859 387
rect 3863 383 3864 387
rect 3858 382 3864 383
rect 1295 380 1369 382
rect 1295 379 1296 380
rect 1290 378 1296 379
rect 2430 377 2436 378
rect 2046 376 2052 377
rect 207 372 262 374
rect 278 373 284 374
rect 207 371 208 372
rect 202 370 208 371
rect 134 368 140 369
rect 278 369 279 373
rect 283 369 284 373
rect 278 368 284 369
rect 438 373 444 374
rect 438 369 439 373
rect 443 369 444 373
rect 438 368 444 369
rect 582 373 588 374
rect 582 369 583 373
rect 587 369 588 373
rect 582 368 588 369
rect 718 373 724 374
rect 718 369 719 373
rect 723 369 724 373
rect 718 368 724 369
rect 846 373 852 374
rect 846 369 847 373
rect 851 369 852 373
rect 846 368 852 369
rect 966 373 972 374
rect 966 369 967 373
rect 971 369 972 373
rect 966 368 972 369
rect 1086 373 1092 374
rect 1086 369 1087 373
rect 1091 369 1092 373
rect 1086 368 1092 369
rect 1206 373 1212 374
rect 1206 369 1207 373
rect 1211 369 1212 373
rect 1206 368 1212 369
rect 1326 373 1332 374
rect 1326 369 1327 373
rect 1331 369 1332 373
rect 1326 368 1332 369
rect 2006 372 2012 373
rect 2006 368 2007 372
rect 2011 368 2012 372
rect 2046 372 2047 376
rect 2051 372 2052 376
rect 2430 373 2431 377
rect 2435 373 2436 377
rect 2430 372 2436 373
rect 2526 377 2532 378
rect 2526 373 2527 377
rect 2531 373 2532 377
rect 2526 372 2532 373
rect 2622 377 2628 378
rect 2622 373 2623 377
rect 2627 373 2628 377
rect 2622 372 2628 373
rect 2718 377 2724 378
rect 2718 373 2719 377
rect 2723 373 2724 377
rect 2718 372 2724 373
rect 2814 377 2820 378
rect 2814 373 2815 377
rect 2819 373 2820 377
rect 2814 372 2820 373
rect 2926 377 2932 378
rect 2926 373 2927 377
rect 2931 373 2932 377
rect 2926 372 2932 373
rect 3062 377 3068 378
rect 3062 373 3063 377
rect 3067 373 3068 377
rect 3062 372 3068 373
rect 3222 377 3228 378
rect 3222 373 3223 377
rect 3227 373 3228 377
rect 3222 372 3228 373
rect 3398 377 3404 378
rect 3398 373 3399 377
rect 3403 373 3404 377
rect 3398 372 3404 373
rect 3590 377 3596 378
rect 3590 373 3591 377
rect 3595 373 3596 377
rect 3590 372 3596 373
rect 3782 377 3788 378
rect 3782 373 3783 377
rect 3787 373 3788 377
rect 3782 372 3788 373
rect 3942 376 3948 377
rect 3942 372 3943 376
rect 3947 372 3948 376
rect 2046 371 2052 372
rect 3942 371 3948 372
rect 110 367 116 368
rect 2006 367 2012 368
rect 2610 363 2616 364
rect 2610 362 2611 363
rect 2497 360 2611 362
rect 546 359 552 360
rect 546 358 547 359
rect 508 356 547 358
rect 508 352 510 356
rect 546 355 547 356
rect 551 355 552 359
rect 2497 356 2499 360
rect 2610 359 2611 360
rect 2615 359 2616 363
rect 3082 363 3088 364
rect 3082 362 3083 363
rect 2610 358 2616 359
rect 2996 360 3083 362
rect 2996 356 2998 360
rect 3082 359 3083 360
rect 3087 359 3088 363
rect 3082 358 3088 359
rect 546 354 552 355
rect 2495 355 2501 356
rect 199 351 208 352
rect 199 347 200 351
rect 207 347 208 351
rect 199 346 208 347
rect 218 351 224 352
rect 218 347 219 351
rect 223 350 224 351
rect 343 351 349 352
rect 343 350 344 351
rect 223 348 344 350
rect 223 347 224 348
rect 218 346 224 347
rect 343 347 344 348
rect 348 347 349 351
rect 343 346 349 347
rect 503 351 510 352
rect 503 347 504 351
rect 508 348 510 351
rect 514 351 520 352
rect 508 347 509 348
rect 503 346 509 347
rect 514 347 515 351
rect 519 350 520 351
rect 647 351 653 352
rect 647 350 648 351
rect 519 348 648 350
rect 519 347 520 348
rect 514 346 520 347
rect 647 347 648 348
rect 652 347 653 351
rect 647 346 653 347
rect 658 351 664 352
rect 658 347 659 351
rect 663 350 664 351
rect 783 351 789 352
rect 783 350 784 351
rect 663 348 784 350
rect 663 347 664 348
rect 658 346 664 347
rect 783 347 784 348
rect 788 347 789 351
rect 783 346 789 347
rect 894 351 900 352
rect 894 347 895 351
rect 899 350 900 351
rect 911 351 917 352
rect 911 350 912 351
rect 899 348 912 350
rect 899 347 900 348
rect 894 346 900 347
rect 911 347 912 348
rect 916 347 917 351
rect 911 346 917 347
rect 922 351 928 352
rect 922 347 923 351
rect 927 350 928 351
rect 1031 351 1037 352
rect 1031 350 1032 351
rect 927 348 1032 350
rect 927 347 928 348
rect 922 346 928 347
rect 1031 347 1032 348
rect 1036 347 1037 351
rect 1031 346 1037 347
rect 1042 351 1048 352
rect 1042 347 1043 351
rect 1047 350 1048 351
rect 1151 351 1157 352
rect 1151 350 1152 351
rect 1047 348 1152 350
rect 1047 347 1048 348
rect 1042 346 1048 347
rect 1151 347 1152 348
rect 1156 347 1157 351
rect 1151 346 1157 347
rect 1162 351 1168 352
rect 1162 347 1163 351
rect 1167 350 1168 351
rect 1271 351 1277 352
rect 1271 350 1272 351
rect 1167 348 1272 350
rect 1167 347 1168 348
rect 1162 346 1168 347
rect 1271 347 1272 348
rect 1276 347 1277 351
rect 1271 346 1277 347
rect 1282 351 1288 352
rect 1282 347 1283 351
rect 1287 350 1288 351
rect 1391 351 1397 352
rect 1391 350 1392 351
rect 1287 348 1392 350
rect 1287 347 1288 348
rect 1282 346 1288 347
rect 1391 347 1392 348
rect 1396 347 1397 351
rect 2495 351 2496 355
rect 2500 351 2501 355
rect 2495 350 2501 351
rect 2506 355 2512 356
rect 2506 351 2507 355
rect 2511 354 2512 355
rect 2591 355 2597 356
rect 2591 354 2592 355
rect 2511 352 2592 354
rect 2511 351 2512 352
rect 2506 350 2512 351
rect 2591 351 2592 352
rect 2596 351 2597 355
rect 2591 350 2597 351
rect 2687 355 2693 356
rect 2687 351 2688 355
rect 2692 354 2693 355
rect 2706 355 2712 356
rect 2706 354 2707 355
rect 2692 352 2707 354
rect 2692 351 2693 352
rect 2687 350 2693 351
rect 2706 351 2707 352
rect 2711 351 2712 355
rect 2706 350 2712 351
rect 2783 355 2789 356
rect 2783 351 2784 355
rect 2788 354 2789 355
rect 2802 355 2808 356
rect 2802 354 2803 355
rect 2788 352 2803 354
rect 2788 351 2789 352
rect 2783 350 2789 351
rect 2802 351 2803 352
rect 2807 351 2808 355
rect 2802 350 2808 351
rect 2879 355 2885 356
rect 2879 351 2880 355
rect 2884 354 2885 355
rect 2934 355 2940 356
rect 2934 354 2935 355
rect 2884 352 2935 354
rect 2884 351 2885 352
rect 2879 350 2885 351
rect 2934 351 2935 352
rect 2939 351 2940 355
rect 2934 350 2940 351
rect 2991 355 2998 356
rect 2991 351 2992 355
rect 2996 352 2998 355
rect 3002 355 3008 356
rect 2996 351 2997 352
rect 2991 350 2997 351
rect 3002 351 3003 355
rect 3007 354 3008 355
rect 3127 355 3133 356
rect 3127 354 3128 355
rect 3007 352 3128 354
rect 3007 351 3008 352
rect 3002 350 3008 351
rect 3127 351 3128 352
rect 3132 351 3133 355
rect 3127 350 3133 351
rect 3138 355 3144 356
rect 3138 351 3139 355
rect 3143 354 3144 355
rect 3287 355 3293 356
rect 3287 354 3288 355
rect 3143 352 3288 354
rect 3143 351 3144 352
rect 3138 350 3144 351
rect 3287 351 3288 352
rect 3292 351 3293 355
rect 3287 350 3293 351
rect 3298 355 3304 356
rect 3298 351 3299 355
rect 3303 354 3304 355
rect 3463 355 3469 356
rect 3463 354 3464 355
rect 3303 352 3464 354
rect 3303 351 3304 352
rect 3298 350 3304 351
rect 3463 351 3464 352
rect 3468 351 3469 355
rect 3463 350 3469 351
rect 3474 355 3480 356
rect 3474 351 3475 355
rect 3479 354 3480 355
rect 3655 355 3661 356
rect 3655 354 3656 355
rect 3479 352 3656 354
rect 3479 351 3480 352
rect 3474 350 3480 351
rect 3655 351 3656 352
rect 3660 351 3661 355
rect 3655 350 3661 351
rect 3730 355 3736 356
rect 3730 351 3731 355
rect 3735 354 3736 355
rect 3847 355 3853 356
rect 3847 354 3848 355
rect 3735 352 3848 354
rect 3735 351 3736 352
rect 3730 350 3736 351
rect 3847 351 3848 352
rect 3852 351 3853 355
rect 3847 350 3853 351
rect 1391 346 1397 347
rect 2602 347 2608 348
rect 2602 343 2603 347
rect 2607 346 2608 347
rect 3498 347 3504 348
rect 3498 346 3499 347
rect 2607 344 2690 346
rect 2607 343 2608 344
rect 2602 342 2608 343
rect 2688 340 2690 344
rect 3020 344 3499 346
rect 3020 340 3022 344
rect 3498 343 3499 344
rect 3503 343 3504 347
rect 3498 342 3504 343
rect 207 339 213 340
rect 207 335 208 339
rect 212 338 213 339
rect 231 339 237 340
rect 231 338 232 339
rect 212 336 232 338
rect 212 335 213 336
rect 207 334 213 335
rect 231 335 232 336
rect 236 335 237 339
rect 231 334 237 335
rect 383 339 389 340
rect 383 335 384 339
rect 388 338 389 339
rect 498 339 504 340
rect 498 338 499 339
rect 388 336 499 338
rect 388 335 389 336
rect 383 334 389 335
rect 498 335 499 336
rect 503 335 504 339
rect 498 334 504 335
rect 543 339 549 340
rect 543 335 544 339
rect 548 338 549 339
rect 618 339 624 340
rect 548 336 614 338
rect 548 335 549 336
rect 543 334 549 335
rect 612 330 614 336
rect 618 335 619 339
rect 623 338 624 339
rect 695 339 701 340
rect 695 338 696 339
rect 623 336 696 338
rect 623 335 624 336
rect 618 334 624 335
rect 695 335 696 336
rect 700 335 701 339
rect 695 334 701 335
rect 794 339 800 340
rect 794 335 795 339
rect 799 338 800 339
rect 839 339 845 340
rect 839 338 840 339
rect 799 336 840 338
rect 799 335 800 336
rect 794 334 800 335
rect 839 335 840 336
rect 844 335 845 339
rect 839 334 845 335
rect 967 339 973 340
rect 967 335 968 339
rect 972 338 973 339
rect 986 339 992 340
rect 986 338 987 339
rect 972 336 987 338
rect 972 335 973 336
rect 967 334 973 335
rect 986 335 987 336
rect 991 335 992 339
rect 986 334 992 335
rect 1095 339 1101 340
rect 1095 335 1096 339
rect 1100 338 1101 339
rect 1114 339 1120 340
rect 1114 338 1115 339
rect 1100 336 1115 338
rect 1100 335 1101 336
rect 1095 334 1101 335
rect 1114 335 1115 336
rect 1119 335 1120 339
rect 1114 334 1120 335
rect 1215 339 1221 340
rect 1215 335 1216 339
rect 1220 338 1221 339
rect 1234 339 1240 340
rect 1234 338 1235 339
rect 1220 336 1235 338
rect 1220 335 1221 336
rect 1215 334 1221 335
rect 1234 335 1235 336
rect 1239 335 1240 339
rect 1234 334 1240 335
rect 1335 339 1341 340
rect 1335 335 1336 339
rect 1340 338 1341 339
rect 1354 339 1360 340
rect 1354 338 1355 339
rect 1340 336 1355 338
rect 1340 335 1341 336
rect 1335 334 1341 335
rect 1354 335 1355 336
rect 1359 335 1360 339
rect 1354 334 1360 335
rect 1455 339 1461 340
rect 1455 335 1456 339
rect 1460 338 1461 339
rect 1602 339 1608 340
rect 1602 338 1603 339
rect 1460 336 1603 338
rect 1460 335 1461 336
rect 1455 334 1461 335
rect 1602 335 1603 336
rect 1607 335 1608 339
rect 1602 334 1608 335
rect 2255 339 2261 340
rect 2255 335 2256 339
rect 2260 338 2261 339
rect 2314 339 2320 340
rect 2260 336 2310 338
rect 2260 335 2261 336
rect 2255 334 2261 335
rect 746 331 752 332
rect 746 330 747 331
rect 612 328 747 330
rect 746 327 747 328
rect 751 327 752 331
rect 2308 330 2310 336
rect 2314 335 2315 339
rect 2319 338 2320 339
rect 2391 339 2397 340
rect 2391 338 2392 339
rect 2319 336 2392 338
rect 2319 335 2320 336
rect 2314 334 2320 335
rect 2391 335 2392 336
rect 2396 335 2397 339
rect 2391 334 2397 335
rect 2535 339 2541 340
rect 2535 335 2536 339
rect 2540 338 2541 339
rect 2687 339 2693 340
rect 2540 336 2682 338
rect 2540 335 2541 336
rect 2535 334 2541 335
rect 2434 331 2440 332
rect 2434 330 2435 331
rect 2308 328 2435 330
rect 746 326 752 327
rect 2434 327 2435 328
rect 2439 327 2440 331
rect 2680 330 2682 336
rect 2687 335 2688 339
rect 2692 335 2693 339
rect 2687 334 2693 335
rect 2698 339 2704 340
rect 2698 335 2699 339
rect 2703 338 2704 339
rect 2847 339 2853 340
rect 2847 338 2848 339
rect 2703 336 2848 338
rect 2703 335 2704 336
rect 2698 334 2704 335
rect 2847 335 2848 336
rect 2852 335 2853 339
rect 2847 334 2853 335
rect 3015 339 3022 340
rect 3015 335 3016 339
rect 3020 336 3022 339
rect 3026 339 3032 340
rect 3020 335 3021 336
rect 3015 334 3021 335
rect 3026 335 3027 339
rect 3031 338 3032 339
rect 3183 339 3189 340
rect 3183 338 3184 339
rect 3031 336 3184 338
rect 3031 335 3032 336
rect 3026 334 3032 335
rect 3183 335 3184 336
rect 3188 335 3189 339
rect 3183 334 3189 335
rect 3194 339 3200 340
rect 3194 335 3195 339
rect 3199 338 3200 339
rect 3359 339 3365 340
rect 3359 338 3360 339
rect 3199 336 3360 338
rect 3199 335 3200 336
rect 3194 334 3200 335
rect 3359 335 3360 336
rect 3364 335 3365 339
rect 3359 334 3365 335
rect 3370 339 3376 340
rect 3370 335 3371 339
rect 3375 338 3376 339
rect 3535 339 3541 340
rect 3535 338 3536 339
rect 3375 336 3536 338
rect 3375 335 3376 336
rect 3370 334 3376 335
rect 3535 335 3536 336
rect 3540 335 3541 339
rect 3535 334 3541 335
rect 3719 339 3725 340
rect 3719 335 3720 339
rect 3724 338 3725 339
rect 3754 339 3760 340
rect 3754 338 3755 339
rect 3724 336 3755 338
rect 3724 335 3725 336
rect 3719 334 3725 335
rect 3754 335 3755 336
rect 3759 335 3760 339
rect 3754 334 3760 335
rect 3882 339 3888 340
rect 3882 335 3883 339
rect 3887 338 3888 339
rect 3903 339 3909 340
rect 3903 338 3904 339
rect 3887 336 3904 338
rect 3887 335 3888 336
rect 3882 334 3888 335
rect 3903 335 3904 336
rect 3908 335 3909 339
rect 3903 334 3909 335
rect 2706 331 2712 332
rect 2706 330 2707 331
rect 2680 328 2707 330
rect 2434 326 2440 327
rect 2706 327 2707 328
rect 2711 327 2712 331
rect 2706 326 2712 327
rect 110 320 116 321
rect 2006 320 2012 321
rect 110 316 111 320
rect 115 316 116 320
rect 110 315 116 316
rect 142 319 148 320
rect 142 315 143 319
rect 147 315 148 319
rect 142 314 148 315
rect 218 319 224 320
rect 218 315 219 319
rect 223 315 224 319
rect 218 314 224 315
rect 318 319 324 320
rect 318 315 319 319
rect 323 315 324 319
rect 318 314 324 315
rect 478 319 484 320
rect 478 315 479 319
rect 483 315 484 319
rect 478 314 484 315
rect 630 319 636 320
rect 630 315 631 319
rect 635 315 636 319
rect 630 314 636 315
rect 774 319 780 320
rect 774 315 775 319
rect 779 315 780 319
rect 774 314 780 315
rect 902 319 908 320
rect 902 315 903 319
rect 907 315 908 319
rect 902 314 908 315
rect 1030 319 1036 320
rect 1030 315 1031 319
rect 1035 315 1036 319
rect 1030 314 1036 315
rect 1150 319 1156 320
rect 1150 315 1151 319
rect 1155 315 1156 319
rect 1150 314 1156 315
rect 1270 319 1276 320
rect 1270 315 1271 319
rect 1275 315 1276 319
rect 1270 314 1276 315
rect 1390 319 1396 320
rect 1390 315 1391 319
rect 1395 315 1396 319
rect 2006 316 2007 320
rect 2011 316 2012 320
rect 2006 315 2012 316
rect 2046 320 2052 321
rect 3942 320 3948 321
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2190 319 2196 320
rect 2190 315 2191 319
rect 2195 315 2196 319
rect 1390 314 1396 315
rect 2190 314 2196 315
rect 2326 319 2332 320
rect 2326 315 2327 319
rect 2331 315 2332 319
rect 2326 314 2332 315
rect 2470 319 2476 320
rect 2470 315 2471 319
rect 2475 315 2476 319
rect 2470 314 2476 315
rect 2622 319 2628 320
rect 2622 315 2623 319
rect 2627 315 2628 319
rect 2622 314 2628 315
rect 2782 319 2788 320
rect 2782 315 2783 319
rect 2787 315 2788 319
rect 2782 314 2788 315
rect 2950 319 2956 320
rect 2950 315 2951 319
rect 2955 315 2956 319
rect 2950 314 2956 315
rect 3118 319 3124 320
rect 3118 315 3119 319
rect 3123 315 3124 319
rect 3118 314 3124 315
rect 3294 319 3300 320
rect 3294 315 3295 319
rect 3299 315 3300 319
rect 3294 314 3300 315
rect 3470 319 3476 320
rect 3470 315 3471 319
rect 3475 315 3476 319
rect 3470 314 3476 315
rect 3654 319 3660 320
rect 3654 315 3655 319
rect 3659 315 3660 319
rect 3654 314 3660 315
rect 3838 319 3844 320
rect 3838 315 3839 319
rect 3843 315 3844 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3838 314 3844 315
rect 220 309 222 314
rect 231 311 237 312
rect 231 307 232 311
rect 236 310 237 311
rect 618 311 624 312
rect 618 310 619 311
rect 236 308 361 310
rect 557 308 619 310
rect 236 307 237 308
rect 231 306 237 307
rect 618 307 619 308
rect 623 307 624 311
rect 746 311 752 312
rect 618 306 624 307
rect 706 307 712 308
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 706 303 707 307
rect 711 303 712 307
rect 746 307 747 311
rect 751 310 752 311
rect 894 311 900 312
rect 751 308 817 310
rect 751 307 752 308
rect 746 306 752 307
rect 894 307 895 311
rect 899 310 900 311
rect 986 311 992 312
rect 899 308 945 310
rect 899 307 900 308
rect 894 306 900 307
rect 986 307 987 311
rect 991 310 992 311
rect 1114 311 1120 312
rect 991 308 1073 310
rect 991 307 992 308
rect 986 306 992 307
rect 1114 307 1115 311
rect 1119 310 1120 311
rect 1234 311 1240 312
rect 1119 308 1193 310
rect 1119 307 1120 308
rect 1114 306 1120 307
rect 1234 307 1235 311
rect 1239 310 1240 311
rect 1354 311 1360 312
rect 1239 308 1313 310
rect 1239 307 1240 308
rect 1234 306 1240 307
rect 1354 307 1355 311
rect 1359 310 1360 311
rect 2314 311 2320 312
rect 2314 310 2315 311
rect 1359 308 1433 310
rect 2269 308 2315 310
rect 1359 307 1360 308
rect 1354 306 1360 307
rect 2314 307 2315 308
rect 2319 307 2320 311
rect 2434 311 2440 312
rect 2314 306 2320 307
rect 2414 307 2420 308
rect 2414 306 2415 307
rect 2405 304 2415 306
rect 706 302 712 303
rect 2006 303 2012 304
rect 110 298 116 299
rect 142 300 148 301
rect 142 296 143 300
rect 147 296 148 300
rect 142 295 148 296
rect 318 300 324 301
rect 318 296 319 300
rect 323 296 324 300
rect 318 295 324 296
rect 478 300 484 301
rect 478 296 479 300
rect 483 296 484 300
rect 478 295 484 296
rect 630 300 636 301
rect 630 296 631 300
rect 635 296 636 300
rect 630 295 636 296
rect 774 300 780 301
rect 774 296 775 300
rect 779 296 780 300
rect 774 295 780 296
rect 902 300 908 301
rect 902 296 903 300
rect 907 296 908 300
rect 902 295 908 296
rect 1030 300 1036 301
rect 1030 296 1031 300
rect 1035 296 1036 300
rect 1030 295 1036 296
rect 1150 300 1156 301
rect 1150 296 1151 300
rect 1155 296 1156 300
rect 1150 295 1156 296
rect 1270 300 1276 301
rect 1270 296 1271 300
rect 1275 296 1276 300
rect 1270 295 1276 296
rect 1390 300 1396 301
rect 1390 296 1391 300
rect 1395 296 1396 300
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 2414 303 2415 304
rect 2419 303 2420 307
rect 2434 307 2435 311
rect 2439 310 2440 311
rect 2698 311 2704 312
rect 2439 308 2513 310
rect 2439 307 2440 308
rect 2434 306 2440 307
rect 2698 307 2699 311
rect 2703 307 2704 311
rect 2698 306 2704 307
rect 2706 311 2712 312
rect 2706 307 2707 311
rect 2711 310 2712 311
rect 3026 311 3032 312
rect 2711 308 2825 310
rect 2711 307 2712 308
rect 2706 306 2712 307
rect 3026 307 3027 311
rect 3031 307 3032 311
rect 3026 306 3032 307
rect 3194 311 3200 312
rect 3194 307 3195 311
rect 3199 307 3200 311
rect 3194 306 3200 307
rect 3370 311 3376 312
rect 3370 307 3371 311
rect 3375 307 3376 311
rect 3370 306 3376 307
rect 3410 311 3416 312
rect 3410 307 3411 311
rect 3415 310 3416 311
rect 3730 311 3736 312
rect 3415 308 3513 310
rect 3415 307 3416 308
rect 3410 306 3416 307
rect 3730 307 3731 311
rect 3735 307 3736 311
rect 3730 306 3736 307
rect 3914 307 3920 308
rect 2414 302 2420 303
rect 3914 303 3915 307
rect 3919 303 3920 307
rect 3914 302 3920 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2190 300 2196 301
rect 1390 295 1396 296
rect 2190 296 2191 300
rect 2195 296 2196 300
rect 2190 295 2196 296
rect 2326 300 2332 301
rect 2326 296 2327 300
rect 2331 296 2332 300
rect 2326 295 2332 296
rect 2470 300 2476 301
rect 2470 296 2471 300
rect 2475 296 2476 300
rect 2470 295 2476 296
rect 2622 300 2628 301
rect 2622 296 2623 300
rect 2627 296 2628 300
rect 2622 295 2628 296
rect 2782 300 2788 301
rect 2782 296 2783 300
rect 2787 296 2788 300
rect 2782 295 2788 296
rect 2950 300 2956 301
rect 2950 296 2951 300
rect 2955 296 2956 300
rect 2950 295 2956 296
rect 3118 300 3124 301
rect 3118 296 3119 300
rect 3123 296 3124 300
rect 3118 295 3124 296
rect 3294 300 3300 301
rect 3294 296 3295 300
rect 3299 296 3300 300
rect 3294 295 3300 296
rect 3470 300 3476 301
rect 3470 296 3471 300
rect 3475 296 3476 300
rect 3470 295 3476 296
rect 3654 300 3660 301
rect 3654 296 3655 300
rect 3659 296 3660 300
rect 3654 295 3660 296
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3838 295 3844 296
rect 2070 240 2076 241
rect 2046 237 2052 238
rect 222 236 228 237
rect 110 233 116 234
rect 110 229 111 233
rect 115 229 116 233
rect 222 232 223 236
rect 227 232 228 236
rect 222 231 228 232
rect 390 236 396 237
rect 390 232 391 236
rect 395 232 396 236
rect 390 231 396 232
rect 558 236 564 237
rect 558 232 559 236
rect 563 232 564 236
rect 558 231 564 232
rect 734 236 740 237
rect 734 232 735 236
rect 739 232 740 236
rect 734 231 740 232
rect 902 236 908 237
rect 902 232 903 236
rect 907 232 908 236
rect 902 231 908 232
rect 1062 236 1068 237
rect 1062 232 1063 236
rect 1067 232 1068 236
rect 1062 231 1068 232
rect 1214 236 1220 237
rect 1214 232 1215 236
rect 1219 232 1220 236
rect 1214 231 1220 232
rect 1358 236 1364 237
rect 1358 232 1359 236
rect 1363 232 1364 236
rect 1358 231 1364 232
rect 1510 236 1516 237
rect 1510 232 1511 236
rect 1515 232 1516 236
rect 1510 231 1516 232
rect 1662 236 1668 237
rect 1662 232 1663 236
rect 1667 232 1668 236
rect 1662 231 1668 232
rect 2006 233 2012 234
rect 110 228 116 229
rect 2006 229 2007 233
rect 2011 229 2012 233
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2214 240 2220 241
rect 2214 236 2215 240
rect 2219 236 2220 240
rect 2214 235 2220 236
rect 2398 240 2404 241
rect 2398 236 2399 240
rect 2403 236 2404 240
rect 2398 235 2404 236
rect 2590 240 2596 241
rect 2590 236 2591 240
rect 2595 236 2596 240
rect 2590 235 2596 236
rect 2790 240 2796 241
rect 2790 236 2791 240
rect 2795 236 2796 240
rect 2790 235 2796 236
rect 2982 240 2988 241
rect 2982 236 2983 240
rect 2987 236 2988 240
rect 2982 235 2988 236
rect 3166 240 3172 241
rect 3166 236 3167 240
rect 3171 236 3172 240
rect 3166 235 3172 236
rect 3342 240 3348 241
rect 3342 236 3343 240
rect 3347 236 3348 240
rect 3342 235 3348 236
rect 3510 240 3516 241
rect 3510 236 3511 240
rect 3515 236 3516 240
rect 3510 235 3516 236
rect 3686 240 3692 241
rect 3686 236 3687 240
rect 3691 236 3692 240
rect 3686 235 3692 236
rect 3838 240 3844 241
rect 3838 236 3839 240
rect 3843 236 3844 240
rect 3838 235 3844 236
rect 3942 237 3948 238
rect 2046 232 2052 233
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 2006 228 2012 229
rect 2146 231 2152 232
rect 298 227 304 228
rect 298 223 299 227
rect 303 223 304 227
rect 298 222 304 223
rect 466 227 472 228
rect 466 223 467 227
rect 471 223 472 227
rect 466 222 472 223
rect 498 227 504 228
rect 498 223 499 227
rect 503 226 504 227
rect 810 227 816 228
rect 503 224 601 226
rect 503 223 504 224
rect 498 222 504 223
rect 810 223 811 227
rect 815 223 816 227
rect 810 222 816 223
rect 895 227 901 228
rect 895 223 896 227
rect 900 226 901 227
rect 1138 227 1144 228
rect 900 224 945 226
rect 900 223 901 224
rect 895 222 901 223
rect 1138 223 1139 227
rect 1143 223 1144 227
rect 1138 222 1144 223
rect 1290 227 1296 228
rect 1290 223 1291 227
rect 1295 223 1296 227
rect 1290 222 1296 223
rect 1434 227 1440 228
rect 1434 223 1435 227
rect 1439 223 1440 227
rect 1434 222 1440 223
rect 1586 227 1592 228
rect 1586 223 1587 227
rect 1591 223 1592 227
rect 1586 222 1592 223
rect 1602 227 1608 228
rect 1602 223 1603 227
rect 1607 226 1608 227
rect 2146 227 2147 231
rect 2151 227 2152 231
rect 2146 226 2152 227
rect 2290 231 2296 232
rect 2290 227 2291 231
rect 2295 227 2296 231
rect 2290 226 2296 227
rect 2474 231 2480 232
rect 2474 227 2475 231
rect 2479 227 2480 231
rect 2474 226 2480 227
rect 2666 231 2672 232
rect 2666 227 2667 231
rect 2671 227 2672 231
rect 2666 226 2672 227
rect 2674 231 2680 232
rect 2674 227 2675 231
rect 2679 230 2680 231
rect 2874 231 2880 232
rect 2679 228 2833 230
rect 2679 227 2680 228
rect 2674 226 2680 227
rect 2874 227 2875 231
rect 2879 230 2880 231
rect 3066 231 3072 232
rect 2879 228 3025 230
rect 2879 227 2880 228
rect 2874 226 2880 227
rect 3066 227 3067 231
rect 3071 230 3072 231
rect 3250 231 3256 232
rect 3071 228 3209 230
rect 3071 227 3072 228
rect 3066 226 3072 227
rect 3250 227 3251 231
rect 3255 230 3256 231
rect 3586 231 3592 232
rect 3255 228 3385 230
rect 3255 227 3256 228
rect 3250 226 3256 227
rect 3586 227 3587 231
rect 3591 227 3592 231
rect 3586 226 3592 227
rect 3754 231 3760 232
rect 3754 227 3755 231
rect 3759 227 3760 231
rect 3754 226 3760 227
rect 3906 231 3912 232
rect 3906 227 3907 231
rect 3911 227 3912 231
rect 3906 226 3912 227
rect 1607 224 1705 226
rect 1607 223 1608 224
rect 1602 222 1608 223
rect 2070 221 2076 222
rect 2046 220 2052 221
rect 222 217 228 218
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 222 213 223 217
rect 227 213 228 217
rect 222 212 228 213
rect 390 217 396 218
rect 390 213 391 217
rect 395 213 396 217
rect 390 212 396 213
rect 558 217 564 218
rect 558 213 559 217
rect 563 213 564 217
rect 558 212 564 213
rect 734 217 740 218
rect 734 213 735 217
rect 739 213 740 217
rect 734 212 740 213
rect 902 217 908 218
rect 902 213 903 217
rect 907 213 908 217
rect 902 212 908 213
rect 1062 217 1068 218
rect 1062 213 1063 217
rect 1067 213 1068 217
rect 1062 212 1068 213
rect 1214 217 1220 218
rect 1214 213 1215 217
rect 1219 213 1220 217
rect 1214 212 1220 213
rect 1358 217 1364 218
rect 1358 213 1359 217
rect 1363 213 1364 217
rect 1358 212 1364 213
rect 1510 217 1516 218
rect 1510 213 1511 217
rect 1515 213 1516 217
rect 1510 212 1516 213
rect 1662 217 1668 218
rect 1662 213 1663 217
rect 1667 213 1668 217
rect 1662 212 1668 213
rect 2006 216 2012 217
rect 2006 212 2007 216
rect 2011 212 2012 216
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2070 217 2071 221
rect 2075 217 2076 221
rect 2070 216 2076 217
rect 2214 221 2220 222
rect 2214 217 2215 221
rect 2219 217 2220 221
rect 2214 216 2220 217
rect 2398 221 2404 222
rect 2398 217 2399 221
rect 2403 217 2404 221
rect 2398 216 2404 217
rect 2590 221 2596 222
rect 2590 217 2591 221
rect 2595 217 2596 221
rect 2590 216 2596 217
rect 2790 221 2796 222
rect 2790 217 2791 221
rect 2795 217 2796 221
rect 2790 216 2796 217
rect 2982 221 2988 222
rect 2982 217 2983 221
rect 2987 217 2988 221
rect 2982 216 2988 217
rect 3166 221 3172 222
rect 3166 217 3167 221
rect 3171 217 3172 221
rect 3166 216 3172 217
rect 3342 221 3348 222
rect 3342 217 3343 221
rect 3347 217 3348 221
rect 3342 216 3348 217
rect 3510 221 3516 222
rect 3510 217 3511 221
rect 3515 217 3516 221
rect 3510 216 3516 217
rect 3686 221 3692 222
rect 3686 217 3687 221
rect 3691 217 3692 221
rect 3686 216 3692 217
rect 3838 221 3844 222
rect 3838 217 3839 221
rect 3843 217 3844 221
rect 3838 216 3844 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 3942 215 3948 216
rect 110 211 116 212
rect 2006 211 2012 212
rect 2674 207 2680 208
rect 2674 206 2675 207
rect 2140 204 2675 206
rect 2140 200 2142 204
rect 2674 203 2675 204
rect 2679 203 2680 207
rect 2674 202 2680 203
rect 2135 199 2142 200
rect 230 195 236 196
rect 230 191 231 195
rect 235 194 236 195
rect 287 195 293 196
rect 287 194 288 195
rect 235 192 288 194
rect 235 191 236 192
rect 230 190 236 191
rect 287 191 288 192
rect 292 191 293 195
rect 287 190 293 191
rect 298 195 304 196
rect 298 191 299 195
rect 303 194 304 195
rect 455 195 461 196
rect 455 194 456 195
rect 303 192 456 194
rect 303 191 304 192
rect 298 190 304 191
rect 455 191 456 192
rect 460 191 461 195
rect 455 190 461 191
rect 466 195 472 196
rect 466 191 467 195
rect 471 194 472 195
rect 623 195 629 196
rect 623 194 624 195
rect 471 192 624 194
rect 471 191 472 192
rect 466 190 472 191
rect 623 191 624 192
rect 628 191 629 195
rect 623 190 629 191
rect 706 195 712 196
rect 706 191 707 195
rect 711 194 712 195
rect 799 195 805 196
rect 799 194 800 195
rect 711 192 800 194
rect 711 191 712 192
rect 706 190 712 191
rect 799 191 800 192
rect 804 191 805 195
rect 799 190 805 191
rect 810 195 816 196
rect 810 191 811 195
rect 815 194 816 195
rect 967 195 973 196
rect 967 194 968 195
rect 815 192 968 194
rect 815 191 816 192
rect 810 190 816 191
rect 967 191 968 192
rect 972 191 973 195
rect 967 190 973 191
rect 1090 195 1096 196
rect 1090 191 1091 195
rect 1095 194 1096 195
rect 1127 195 1133 196
rect 1127 194 1128 195
rect 1095 192 1128 194
rect 1095 191 1096 192
rect 1090 190 1096 191
rect 1127 191 1128 192
rect 1132 191 1133 195
rect 1127 190 1133 191
rect 1138 195 1144 196
rect 1138 191 1139 195
rect 1143 194 1144 195
rect 1279 195 1285 196
rect 1279 194 1280 195
rect 1143 192 1280 194
rect 1143 191 1144 192
rect 1138 190 1144 191
rect 1279 191 1280 192
rect 1284 191 1285 195
rect 1279 190 1285 191
rect 1290 195 1296 196
rect 1290 191 1291 195
rect 1295 194 1296 195
rect 1423 195 1429 196
rect 1423 194 1424 195
rect 1295 192 1424 194
rect 1295 191 1296 192
rect 1290 190 1296 191
rect 1423 191 1424 192
rect 1428 191 1429 195
rect 1423 190 1429 191
rect 1434 195 1440 196
rect 1434 191 1435 195
rect 1439 194 1440 195
rect 1575 195 1581 196
rect 1575 194 1576 195
rect 1439 192 1576 194
rect 1439 191 1440 192
rect 1434 190 1440 191
rect 1575 191 1576 192
rect 1580 191 1581 195
rect 1575 190 1581 191
rect 1586 195 1592 196
rect 1586 191 1587 195
rect 1591 194 1592 195
rect 1727 195 1733 196
rect 1727 194 1728 195
rect 1591 192 1728 194
rect 1591 191 1592 192
rect 1586 190 1592 191
rect 1727 191 1728 192
rect 1732 191 1733 195
rect 2135 195 2136 199
rect 2140 196 2142 199
rect 2146 199 2152 200
rect 2140 195 2141 196
rect 2135 194 2141 195
rect 2146 195 2147 199
rect 2151 198 2152 199
rect 2279 199 2285 200
rect 2279 198 2280 199
rect 2151 196 2280 198
rect 2151 195 2152 196
rect 2146 194 2152 195
rect 2279 195 2280 196
rect 2284 195 2285 199
rect 2279 194 2285 195
rect 2414 199 2420 200
rect 2414 195 2415 199
rect 2419 198 2420 199
rect 2463 199 2469 200
rect 2463 198 2464 199
rect 2419 196 2464 198
rect 2419 195 2420 196
rect 2414 194 2420 195
rect 2463 195 2464 196
rect 2468 195 2469 199
rect 2463 194 2469 195
rect 2474 199 2480 200
rect 2474 195 2475 199
rect 2479 198 2480 199
rect 2655 199 2661 200
rect 2655 198 2656 199
rect 2479 196 2656 198
rect 2479 195 2480 196
rect 2474 194 2480 195
rect 2655 195 2656 196
rect 2660 195 2661 199
rect 2655 194 2661 195
rect 2666 199 2672 200
rect 2666 195 2667 199
rect 2671 198 2672 199
rect 2855 199 2861 200
rect 2855 198 2856 199
rect 2671 196 2856 198
rect 2671 195 2672 196
rect 2666 194 2672 195
rect 2855 195 2856 196
rect 2860 195 2861 199
rect 2855 194 2861 195
rect 3047 199 3053 200
rect 3047 195 3048 199
rect 3052 198 3053 199
rect 3066 199 3072 200
rect 3066 198 3067 199
rect 3052 196 3067 198
rect 3052 195 3053 196
rect 3047 194 3053 195
rect 3066 195 3067 196
rect 3071 195 3072 199
rect 3066 194 3072 195
rect 3231 199 3237 200
rect 3231 195 3232 199
rect 3236 198 3237 199
rect 3250 199 3256 200
rect 3250 198 3251 199
rect 3236 196 3251 198
rect 3236 195 3237 196
rect 3231 194 3237 195
rect 3250 195 3251 196
rect 3255 195 3256 199
rect 3250 194 3256 195
rect 3407 199 3416 200
rect 3407 195 3408 199
rect 3415 195 3416 199
rect 3407 194 3416 195
rect 3575 199 3581 200
rect 3575 195 3576 199
rect 3580 198 3581 199
rect 3586 199 3592 200
rect 3580 195 3582 198
rect 3575 194 3582 195
rect 3586 195 3587 199
rect 3591 198 3592 199
rect 3751 199 3757 200
rect 3751 198 3752 199
rect 3591 196 3752 198
rect 3591 195 3592 196
rect 3586 194 3592 195
rect 3751 195 3752 196
rect 3756 195 3757 199
rect 3751 194 3757 195
rect 3903 199 3909 200
rect 3903 195 3904 199
rect 3908 198 3909 199
rect 3914 199 3920 200
rect 3914 198 3915 199
rect 3908 196 3915 198
rect 3908 195 3909 196
rect 3903 194 3909 195
rect 3914 195 3915 196
rect 3919 195 3920 199
rect 3914 194 3920 195
rect 1727 190 1733 191
rect 3580 190 3582 194
rect 3630 191 3636 192
rect 3630 190 3631 191
rect 3580 188 3631 190
rect 3630 187 3631 188
rect 3635 187 3636 191
rect 3630 186 3636 187
rect 2135 163 2141 164
rect 2135 159 2136 163
rect 2140 162 2141 163
rect 2159 163 2165 164
rect 2159 162 2160 163
rect 2140 160 2160 162
rect 2140 159 2141 160
rect 2135 158 2141 159
rect 2159 159 2160 160
rect 2164 159 2165 163
rect 2159 158 2165 159
rect 2255 163 2261 164
rect 2255 159 2256 163
rect 2260 159 2261 163
rect 2255 158 2261 159
rect 2290 163 2296 164
rect 2290 159 2291 163
rect 2295 162 2296 163
rect 2407 163 2413 164
rect 2407 162 2408 163
rect 2295 160 2408 162
rect 2295 159 2296 160
rect 2290 158 2296 159
rect 2407 159 2408 160
rect 2412 159 2413 163
rect 2407 158 2413 159
rect 2418 163 2424 164
rect 2418 159 2419 163
rect 2423 162 2424 163
rect 2559 163 2565 164
rect 2559 162 2560 163
rect 2423 160 2560 162
rect 2423 159 2424 160
rect 2418 158 2424 159
rect 2559 159 2560 160
rect 2564 159 2565 163
rect 2559 158 2565 159
rect 2570 163 2576 164
rect 2570 159 2571 163
rect 2575 162 2576 163
rect 2711 163 2717 164
rect 2711 162 2712 163
rect 2575 160 2712 162
rect 2575 159 2576 160
rect 2570 158 2576 159
rect 2711 159 2712 160
rect 2716 159 2717 163
rect 2711 158 2717 159
rect 2863 163 2869 164
rect 2863 159 2864 163
rect 2868 162 2869 163
rect 2874 163 2880 164
rect 2874 162 2875 163
rect 2868 160 2875 162
rect 2868 159 2869 160
rect 2863 158 2869 159
rect 2874 159 2875 160
rect 2879 159 2880 163
rect 2874 158 2880 159
rect 2918 163 2924 164
rect 2918 159 2919 163
rect 2923 162 2924 163
rect 3007 163 3013 164
rect 3007 162 3008 163
rect 2923 160 3008 162
rect 2923 159 2924 160
rect 2918 158 2924 159
rect 3007 159 3008 160
rect 3012 159 3013 163
rect 3007 158 3013 159
rect 3018 163 3024 164
rect 3018 159 3019 163
rect 3023 162 3024 163
rect 3135 163 3141 164
rect 3135 162 3136 163
rect 3023 160 3136 162
rect 3023 159 3024 160
rect 3018 158 3024 159
rect 3135 159 3136 160
rect 3140 159 3141 163
rect 3135 158 3141 159
rect 3146 163 3152 164
rect 3146 159 3147 163
rect 3151 162 3152 163
rect 3255 163 3261 164
rect 3255 162 3256 163
rect 3151 160 3256 162
rect 3151 159 3152 160
rect 3146 158 3152 159
rect 3255 159 3256 160
rect 3260 159 3261 163
rect 3255 158 3261 159
rect 3266 163 3272 164
rect 3266 159 3267 163
rect 3271 162 3272 163
rect 3375 163 3381 164
rect 3375 162 3376 163
rect 3271 160 3376 162
rect 3271 159 3272 160
rect 3266 158 3272 159
rect 3375 159 3376 160
rect 3380 159 3381 163
rect 3375 158 3381 159
rect 3386 163 3392 164
rect 3386 159 3387 163
rect 3391 162 3392 163
rect 3487 163 3493 164
rect 3487 162 3488 163
rect 3391 160 3488 162
rect 3391 159 3392 160
rect 3386 158 3392 159
rect 3487 159 3488 160
rect 3492 159 3493 163
rect 3487 158 3493 159
rect 3498 163 3504 164
rect 3498 159 3499 163
rect 3503 162 3504 163
rect 3591 163 3597 164
rect 3591 162 3592 163
rect 3503 160 3592 162
rect 3503 159 3504 160
rect 3498 158 3504 159
rect 3591 159 3592 160
rect 3596 159 3597 163
rect 3591 158 3597 159
rect 3602 163 3608 164
rect 3602 159 3603 163
rect 3607 162 3608 163
rect 3703 163 3709 164
rect 3703 162 3704 163
rect 3607 160 3704 162
rect 3607 159 3608 160
rect 3602 158 3608 159
rect 3703 159 3704 160
rect 3708 159 3709 163
rect 3703 158 3709 159
rect 3807 163 3813 164
rect 3807 159 3808 163
rect 3812 162 3813 163
rect 3826 163 3832 164
rect 3826 162 3827 163
rect 3812 160 3827 162
rect 3812 159 3813 160
rect 3807 158 3813 159
rect 3826 159 3827 160
rect 3831 159 3832 163
rect 3826 158 3832 159
rect 3903 163 3912 164
rect 3903 159 3904 163
rect 3911 159 3912 163
rect 3903 158 3912 159
rect 2257 154 2259 158
rect 2578 155 2584 156
rect 2578 154 2579 155
rect 2257 152 2579 154
rect 215 151 221 152
rect 215 147 216 151
rect 220 150 221 151
rect 239 151 245 152
rect 239 150 240 151
rect 220 148 240 150
rect 220 147 221 148
rect 215 146 221 147
rect 239 147 240 148
rect 244 147 245 151
rect 239 146 245 147
rect 311 151 317 152
rect 311 147 312 151
rect 316 150 317 151
rect 335 151 341 152
rect 335 150 336 151
rect 316 148 336 150
rect 316 147 317 148
rect 311 146 317 147
rect 335 147 336 148
rect 340 147 341 151
rect 335 146 341 147
rect 407 151 413 152
rect 407 147 408 151
rect 412 150 413 151
rect 426 151 432 152
rect 426 150 427 151
rect 412 148 427 150
rect 412 147 413 148
rect 407 146 413 147
rect 426 147 427 148
rect 431 147 432 151
rect 426 146 432 147
rect 503 151 509 152
rect 503 147 504 151
rect 508 150 509 151
rect 522 151 528 152
rect 522 150 523 151
rect 508 148 523 150
rect 508 147 509 148
rect 503 146 509 147
rect 522 147 523 148
rect 527 147 528 151
rect 522 146 528 147
rect 599 151 605 152
rect 599 147 600 151
rect 604 150 605 151
rect 618 151 624 152
rect 618 150 619 151
rect 604 148 619 150
rect 604 147 605 148
rect 599 146 605 147
rect 618 147 619 148
rect 623 147 624 151
rect 618 146 624 147
rect 695 151 701 152
rect 695 147 696 151
rect 700 150 701 151
rect 714 151 720 152
rect 714 150 715 151
rect 700 148 715 150
rect 700 147 701 148
rect 695 146 701 147
rect 714 147 715 148
rect 719 147 720 151
rect 714 146 720 147
rect 791 151 797 152
rect 791 147 792 151
rect 796 150 797 151
rect 810 151 816 152
rect 810 150 811 151
rect 796 148 811 150
rect 796 147 797 148
rect 791 146 797 147
rect 810 147 811 148
rect 815 147 816 151
rect 810 146 816 147
rect 887 151 893 152
rect 887 147 888 151
rect 892 150 893 151
rect 895 151 901 152
rect 895 150 896 151
rect 892 148 896 150
rect 892 147 893 148
rect 887 146 893 147
rect 895 147 896 148
rect 900 147 901 151
rect 895 146 901 147
rect 983 151 989 152
rect 983 147 984 151
rect 988 150 989 151
rect 994 151 1000 152
rect 988 147 990 150
rect 983 146 990 147
rect 994 147 995 151
rect 999 150 1000 151
rect 1079 151 1085 152
rect 1079 150 1080 151
rect 999 148 1080 150
rect 999 147 1000 148
rect 994 146 1000 147
rect 1079 147 1080 148
rect 1084 147 1085 151
rect 1079 146 1085 147
rect 1175 151 1181 152
rect 1175 147 1176 151
rect 1180 150 1181 151
rect 1194 151 1200 152
rect 1194 150 1195 151
rect 1180 148 1195 150
rect 1180 147 1181 148
rect 1175 146 1181 147
rect 1194 147 1195 148
rect 1199 147 1200 151
rect 1194 146 1200 147
rect 1271 151 1277 152
rect 1271 147 1272 151
rect 1276 150 1277 151
rect 1290 151 1296 152
rect 1290 150 1291 151
rect 1276 148 1291 150
rect 1276 147 1277 148
rect 1271 146 1277 147
rect 1290 147 1291 148
rect 1295 147 1296 151
rect 1290 146 1296 147
rect 1367 151 1373 152
rect 1367 147 1368 151
rect 1372 150 1373 151
rect 1399 151 1405 152
rect 1399 150 1400 151
rect 1372 148 1400 150
rect 1372 147 1373 148
rect 1367 146 1373 147
rect 1399 147 1400 148
rect 1404 147 1405 151
rect 1399 146 1405 147
rect 1471 151 1477 152
rect 1471 147 1472 151
rect 1476 150 1477 151
rect 1503 151 1509 152
rect 1503 150 1504 151
rect 1476 148 1504 150
rect 1476 147 1477 148
rect 1471 146 1477 147
rect 1503 147 1504 148
rect 1508 147 1509 151
rect 1503 146 1509 147
rect 1575 151 1581 152
rect 1575 147 1576 151
rect 1580 150 1581 151
rect 1607 151 1613 152
rect 1607 150 1608 151
rect 1580 148 1608 150
rect 1580 147 1581 148
rect 1575 146 1581 147
rect 1607 147 1608 148
rect 1612 147 1613 151
rect 1607 146 1613 147
rect 1679 151 1685 152
rect 1679 147 1680 151
rect 1684 150 1685 151
rect 1698 151 1704 152
rect 1698 150 1699 151
rect 1684 148 1699 150
rect 1684 147 1685 148
rect 1679 146 1685 147
rect 1698 147 1699 148
rect 1703 147 1704 151
rect 1698 146 1704 147
rect 1775 151 1781 152
rect 1775 147 1776 151
rect 1780 150 1781 151
rect 1794 151 1800 152
rect 1794 150 1795 151
rect 1780 148 1795 150
rect 1780 147 1781 148
rect 1775 146 1781 147
rect 1794 147 1795 148
rect 1799 147 1800 151
rect 1794 146 1800 147
rect 1871 151 1877 152
rect 1871 147 1872 151
rect 1876 150 1877 151
rect 1890 151 1896 152
rect 1890 150 1891 151
rect 1876 148 1891 150
rect 1876 147 1877 148
rect 1871 146 1877 147
rect 1890 147 1891 148
rect 1895 147 1896 151
rect 1890 146 1896 147
rect 1967 151 1973 152
rect 1967 147 1968 151
rect 1972 150 1973 151
rect 2578 151 2579 152
rect 2583 151 2584 155
rect 2578 150 2584 151
rect 1972 148 2058 150
rect 1972 147 1973 148
rect 1967 146 1973 147
rect 988 142 990 146
rect 2046 144 2052 145
rect 1098 143 1104 144
rect 1098 142 1099 143
rect 988 140 1099 142
rect 1098 139 1099 140
rect 1103 139 1104 143
rect 2046 140 2047 144
rect 2051 140 2052 144
rect 2046 139 2052 140
rect 1098 138 1104 139
rect 2056 134 2058 148
rect 3942 144 3948 145
rect 2070 143 2076 144
rect 2070 139 2071 143
rect 2075 139 2076 143
rect 2070 138 2076 139
rect 2190 143 2196 144
rect 2190 139 2191 143
rect 2195 139 2196 143
rect 2190 138 2196 139
rect 2342 143 2348 144
rect 2342 139 2343 143
rect 2347 139 2348 143
rect 2342 138 2348 139
rect 2494 143 2500 144
rect 2494 139 2495 143
rect 2499 139 2500 143
rect 2494 138 2500 139
rect 2646 143 2652 144
rect 2646 139 2647 143
rect 2651 139 2652 143
rect 2646 138 2652 139
rect 2798 143 2804 144
rect 2798 139 2799 143
rect 2803 139 2804 143
rect 2798 138 2804 139
rect 2942 143 2948 144
rect 2942 139 2943 143
rect 2947 139 2948 143
rect 2942 138 2948 139
rect 3070 143 3076 144
rect 3070 139 3071 143
rect 3075 139 3076 143
rect 3070 138 3076 139
rect 3190 143 3196 144
rect 3190 139 3191 143
rect 3195 139 3196 143
rect 3190 138 3196 139
rect 3310 143 3316 144
rect 3310 139 3311 143
rect 3315 139 3316 143
rect 3310 138 3316 139
rect 3422 143 3428 144
rect 3422 139 3423 143
rect 3427 139 3428 143
rect 3422 138 3428 139
rect 3526 143 3532 144
rect 3526 139 3527 143
rect 3531 139 3532 143
rect 3526 138 3532 139
rect 3638 143 3644 144
rect 3638 139 3639 143
rect 3643 139 3644 143
rect 3638 138 3644 139
rect 3742 143 3748 144
rect 3742 139 3743 143
rect 3747 139 3748 143
rect 3742 138 3748 139
rect 3838 143 3844 144
rect 3838 139 3839 143
rect 3843 139 3844 143
rect 3942 140 3943 144
rect 3947 140 3948 144
rect 3942 139 3948 140
rect 3838 138 3844 139
rect 2159 135 2165 136
rect 110 132 116 133
rect 2006 132 2012 133
rect 2056 132 2113 134
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 150 131 156 132
rect 150 127 151 131
rect 155 127 156 131
rect 150 126 156 127
rect 246 131 252 132
rect 246 127 247 131
rect 251 127 252 131
rect 246 126 252 127
rect 342 131 348 132
rect 342 127 343 131
rect 347 127 348 131
rect 342 126 348 127
rect 438 131 444 132
rect 438 127 439 131
rect 443 127 444 131
rect 438 126 444 127
rect 534 131 540 132
rect 534 127 535 131
rect 539 127 540 131
rect 534 126 540 127
rect 630 131 636 132
rect 630 127 631 131
rect 635 127 636 131
rect 630 126 636 127
rect 726 131 732 132
rect 726 127 727 131
rect 731 127 732 131
rect 726 126 732 127
rect 822 131 828 132
rect 822 127 823 131
rect 827 127 828 131
rect 822 126 828 127
rect 918 131 924 132
rect 918 127 919 131
rect 923 127 924 131
rect 918 126 924 127
rect 1014 131 1020 132
rect 1014 127 1015 131
rect 1019 127 1020 131
rect 1014 126 1020 127
rect 1110 131 1116 132
rect 1110 127 1111 131
rect 1115 127 1116 131
rect 1110 126 1116 127
rect 1206 131 1212 132
rect 1206 127 1207 131
rect 1211 127 1212 131
rect 1206 126 1212 127
rect 1302 131 1308 132
rect 1302 127 1303 131
rect 1307 127 1308 131
rect 1302 126 1308 127
rect 1406 131 1412 132
rect 1406 127 1407 131
rect 1411 127 1412 131
rect 1406 126 1412 127
rect 1510 131 1516 132
rect 1510 127 1511 131
rect 1515 127 1516 131
rect 1510 126 1516 127
rect 1614 131 1620 132
rect 1614 127 1615 131
rect 1619 127 1620 131
rect 1614 126 1620 127
rect 1710 131 1716 132
rect 1710 127 1711 131
rect 1715 127 1716 131
rect 1710 126 1716 127
rect 1806 131 1812 132
rect 1806 127 1807 131
rect 1811 127 1812 131
rect 1806 126 1812 127
rect 1902 131 1908 132
rect 1902 127 1903 131
rect 1907 127 1908 131
rect 2006 128 2007 132
rect 2011 128 2012 132
rect 2159 131 2160 135
rect 2164 134 2165 135
rect 2418 135 2424 136
rect 2164 132 2233 134
rect 2164 131 2165 132
rect 2159 130 2165 131
rect 2418 131 2419 135
rect 2423 131 2424 135
rect 2418 130 2424 131
rect 2570 135 2576 136
rect 2570 131 2571 135
rect 2575 131 2576 135
rect 2570 130 2576 131
rect 2578 135 2584 136
rect 2578 131 2579 135
rect 2583 134 2584 135
rect 2918 135 2924 136
rect 2918 134 2919 135
rect 2583 132 2689 134
rect 2877 132 2919 134
rect 2583 131 2584 132
rect 2578 130 2584 131
rect 2918 131 2919 132
rect 2923 131 2924 135
rect 2918 130 2924 131
rect 3018 135 3024 136
rect 3018 131 3019 135
rect 3023 131 3024 135
rect 3018 130 3024 131
rect 3146 135 3152 136
rect 3146 131 3147 135
rect 3151 131 3152 135
rect 3146 130 3152 131
rect 3266 135 3272 136
rect 3266 131 3267 135
rect 3271 131 3272 135
rect 3266 130 3272 131
rect 3386 135 3392 136
rect 3386 131 3387 135
rect 3391 131 3392 135
rect 3386 130 3392 131
rect 3498 135 3504 136
rect 3498 131 3499 135
rect 3503 131 3504 135
rect 3498 130 3504 131
rect 3602 135 3608 136
rect 3602 131 3603 135
rect 3607 131 3608 135
rect 3602 130 3608 131
rect 3630 135 3636 136
rect 3630 131 3631 135
rect 3635 134 3636 135
rect 3826 135 3832 136
rect 3635 132 3681 134
rect 3635 131 3636 132
rect 3630 130 3636 131
rect 3826 131 3827 135
rect 3831 134 3832 135
rect 3831 132 3881 134
rect 3831 131 3832 132
rect 3826 130 3832 131
rect 2006 127 2012 128
rect 2046 127 2052 128
rect 1902 126 1908 127
rect 226 123 232 124
rect 226 119 227 123
rect 231 119 232 123
rect 226 118 232 119
rect 239 123 245 124
rect 239 119 240 123
rect 244 122 245 123
rect 335 123 341 124
rect 244 120 289 122
rect 244 119 245 120
rect 239 118 245 119
rect 335 119 336 123
rect 340 122 341 123
rect 426 123 432 124
rect 340 120 385 122
rect 340 119 341 120
rect 335 118 341 119
rect 426 119 427 123
rect 431 122 432 123
rect 522 123 528 124
rect 431 120 481 122
rect 431 119 432 120
rect 426 118 432 119
rect 522 119 523 123
rect 527 122 528 123
rect 618 123 624 124
rect 527 120 577 122
rect 527 119 528 120
rect 522 118 528 119
rect 618 119 619 123
rect 623 122 624 123
rect 714 123 720 124
rect 623 120 673 122
rect 623 119 624 120
rect 618 118 624 119
rect 714 119 715 123
rect 719 122 720 123
rect 810 123 816 124
rect 719 120 769 122
rect 719 119 720 120
rect 714 118 720 119
rect 810 119 811 123
rect 815 122 816 123
rect 994 123 1000 124
rect 815 120 865 122
rect 815 119 816 120
rect 810 118 816 119
rect 994 119 995 123
rect 999 119 1000 123
rect 994 118 1000 119
rect 1090 123 1096 124
rect 1090 119 1091 123
rect 1095 119 1096 123
rect 1090 118 1096 119
rect 1098 123 1104 124
rect 1098 119 1099 123
rect 1103 122 1104 123
rect 1194 123 1200 124
rect 1103 120 1153 122
rect 1103 119 1104 120
rect 1098 118 1104 119
rect 1194 119 1195 123
rect 1199 122 1200 123
rect 1290 123 1296 124
rect 1199 120 1249 122
rect 1199 119 1200 120
rect 1194 118 1200 119
rect 1290 119 1291 123
rect 1295 122 1296 123
rect 1399 123 1405 124
rect 1295 120 1345 122
rect 1295 119 1296 120
rect 1290 118 1296 119
rect 1399 119 1400 123
rect 1404 122 1405 123
rect 1503 123 1509 124
rect 1404 120 1449 122
rect 1404 119 1405 120
rect 1399 118 1405 119
rect 1503 119 1504 123
rect 1508 122 1509 123
rect 1607 123 1613 124
rect 1508 120 1553 122
rect 1508 119 1509 120
rect 1503 118 1509 119
rect 1607 119 1608 123
rect 1612 122 1613 123
rect 1698 123 1704 124
rect 1612 120 1657 122
rect 1612 119 1613 120
rect 1607 118 1613 119
rect 1698 119 1699 123
rect 1703 122 1704 123
rect 1794 123 1800 124
rect 1703 120 1753 122
rect 1703 119 1704 120
rect 1698 118 1704 119
rect 1794 119 1795 123
rect 1799 122 1800 123
rect 1890 123 1896 124
rect 1799 120 1849 122
rect 1799 119 1800 120
rect 1794 118 1800 119
rect 1890 119 1891 123
rect 1895 122 1896 123
rect 2046 123 2047 127
rect 2051 123 2052 127
rect 3942 127 3948 128
rect 2046 122 2052 123
rect 2070 124 2076 125
rect 1895 120 1945 122
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 1895 119 1896 120
rect 2070 119 2076 120
rect 2190 124 2196 125
rect 2190 120 2191 124
rect 2195 120 2196 124
rect 2190 119 2196 120
rect 2342 124 2348 125
rect 2342 120 2343 124
rect 2347 120 2348 124
rect 2342 119 2348 120
rect 2494 124 2500 125
rect 2494 120 2495 124
rect 2499 120 2500 124
rect 2494 119 2500 120
rect 2646 124 2652 125
rect 2646 120 2647 124
rect 2651 120 2652 124
rect 2646 119 2652 120
rect 2798 124 2804 125
rect 2798 120 2799 124
rect 2803 120 2804 124
rect 2798 119 2804 120
rect 2942 124 2948 125
rect 2942 120 2943 124
rect 2947 120 2948 124
rect 2942 119 2948 120
rect 3070 124 3076 125
rect 3070 120 3071 124
rect 3075 120 3076 124
rect 3070 119 3076 120
rect 3190 124 3196 125
rect 3190 120 3191 124
rect 3195 120 3196 124
rect 3190 119 3196 120
rect 3310 124 3316 125
rect 3310 120 3311 124
rect 3315 120 3316 124
rect 3310 119 3316 120
rect 3422 124 3428 125
rect 3422 120 3423 124
rect 3427 120 3428 124
rect 3422 119 3428 120
rect 3526 124 3532 125
rect 3526 120 3527 124
rect 3531 120 3532 124
rect 3526 119 3532 120
rect 3638 124 3644 125
rect 3638 120 3639 124
rect 3643 120 3644 124
rect 3638 119 3644 120
rect 3742 124 3748 125
rect 3742 120 3743 124
rect 3747 120 3748 124
rect 3742 119 3748 120
rect 3838 124 3844 125
rect 3838 120 3839 124
rect 3843 120 3844 124
rect 3942 123 3943 127
rect 3947 123 3948 127
rect 3942 122 3948 123
rect 3838 119 3844 120
rect 1890 118 1896 119
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 2006 115 2012 116
rect 110 110 116 111
rect 150 112 156 113
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 246 112 252 113
rect 246 108 247 112
rect 251 108 252 112
rect 246 107 252 108
rect 342 112 348 113
rect 342 108 343 112
rect 347 108 348 112
rect 342 107 348 108
rect 438 112 444 113
rect 438 108 439 112
rect 443 108 444 112
rect 438 107 444 108
rect 534 112 540 113
rect 534 108 535 112
rect 539 108 540 112
rect 534 107 540 108
rect 630 112 636 113
rect 630 108 631 112
rect 635 108 636 112
rect 630 107 636 108
rect 726 112 732 113
rect 726 108 727 112
rect 731 108 732 112
rect 726 107 732 108
rect 822 112 828 113
rect 822 108 823 112
rect 827 108 828 112
rect 822 107 828 108
rect 918 112 924 113
rect 918 108 919 112
rect 923 108 924 112
rect 918 107 924 108
rect 1014 112 1020 113
rect 1014 108 1015 112
rect 1019 108 1020 112
rect 1014 107 1020 108
rect 1110 112 1116 113
rect 1110 108 1111 112
rect 1115 108 1116 112
rect 1110 107 1116 108
rect 1206 112 1212 113
rect 1206 108 1207 112
rect 1211 108 1212 112
rect 1206 107 1212 108
rect 1302 112 1308 113
rect 1302 108 1303 112
rect 1307 108 1308 112
rect 1302 107 1308 108
rect 1406 112 1412 113
rect 1406 108 1407 112
rect 1411 108 1412 112
rect 1406 107 1412 108
rect 1510 112 1516 113
rect 1510 108 1511 112
rect 1515 108 1516 112
rect 1510 107 1516 108
rect 1614 112 1620 113
rect 1614 108 1615 112
rect 1619 108 1620 112
rect 1614 107 1620 108
rect 1710 112 1716 113
rect 1710 108 1711 112
rect 1715 108 1716 112
rect 1710 107 1716 108
rect 1806 112 1812 113
rect 1806 108 1807 112
rect 1811 108 1812 112
rect 1806 107 1812 108
rect 1902 112 1908 113
rect 1902 108 1903 112
rect 1907 108 1908 112
rect 2006 111 2007 115
rect 2011 111 2012 115
rect 2006 110 2012 111
rect 1902 107 1908 108
<< m3c >>
rect 2047 3985 2051 3989
rect 2071 3988 2075 3992
rect 2327 3988 2331 3992
rect 2591 3988 2595 3992
rect 2839 3988 2843 3992
rect 3087 3988 3091 3992
rect 3343 3988 3347 3992
rect 3943 3985 3947 3989
rect 2147 3979 2151 3983
rect 2195 3979 2199 3983
rect 2667 3979 2671 3983
rect 2915 3979 2919 3983
rect 3163 3979 3167 3983
rect 3243 3979 3247 3983
rect 111 3965 115 3969
rect 311 3968 315 3972
rect 511 3968 515 3972
rect 703 3968 707 3972
rect 887 3968 891 3972
rect 1063 3968 1067 3972
rect 1231 3968 1235 3972
rect 1383 3968 1387 3972
rect 1519 3968 1523 3972
rect 1655 3968 1659 3972
rect 1791 3968 1795 3972
rect 1903 3968 1907 3972
rect 2007 3965 2011 3969
rect 2047 3968 2051 3972
rect 2071 3969 2075 3973
rect 2327 3969 2331 3973
rect 2591 3969 2595 3973
rect 2839 3969 2843 3973
rect 3087 3969 3091 3973
rect 3343 3969 3347 3973
rect 3943 3968 3947 3972
rect 463 3959 467 3963
rect 587 3959 591 3963
rect 779 3959 783 3963
rect 111 3948 115 3952
rect 311 3949 315 3953
rect 511 3949 515 3953
rect 703 3949 707 3953
rect 635 3943 639 3947
rect 1139 3959 1143 3963
rect 1307 3959 1311 3963
rect 1459 3959 1463 3963
rect 1595 3959 1599 3963
rect 1731 3959 1735 3963
rect 1867 3959 1871 3963
rect 887 3949 891 3953
rect 1063 3949 1067 3953
rect 1231 3949 1235 3953
rect 1383 3949 1387 3953
rect 1519 3949 1523 3953
rect 1655 3949 1659 3953
rect 1791 3949 1795 3953
rect 1903 3949 1907 3953
rect 2007 3948 2011 3952
rect 2147 3947 2151 3951
rect 2659 3947 2660 3951
rect 2660 3947 2663 3951
rect 2667 3947 2671 3951
rect 2915 3947 2919 3951
rect 3163 3947 3167 3951
rect 2195 3935 2196 3939
rect 2196 3935 2199 3939
rect 2203 3935 2207 3939
rect 2347 3935 2351 3939
rect 2515 3935 2519 3939
rect 2691 3935 2695 3939
rect 3051 3935 3052 3939
rect 3052 3935 3055 3939
rect 3243 3935 3244 3939
rect 3244 3935 3247 3939
rect 3251 3935 3255 3939
rect 3443 3935 3447 3939
rect 403 3927 407 3931
rect 463 3927 467 3931
rect 587 3927 591 3931
rect 779 3927 783 3931
rect 1131 3927 1132 3931
rect 1132 3927 1135 3931
rect 1139 3927 1143 3931
rect 1307 3927 1311 3931
rect 1459 3927 1463 3931
rect 1595 3927 1599 3931
rect 1731 3927 1735 3931
rect 1867 3927 1871 3931
rect 2659 3923 2663 3927
rect 303 3915 307 3919
rect 355 3915 359 3919
rect 635 3915 636 3919
rect 636 3915 639 3919
rect 643 3915 647 3919
rect 811 3915 815 3919
rect 987 3915 991 3919
rect 1371 3915 1375 3919
rect 1707 3915 1711 3919
rect 2047 3916 2051 3920
rect 2127 3915 2131 3919
rect 2271 3915 2275 3919
rect 2439 3915 2443 3919
rect 2615 3915 2619 3919
rect 2799 3915 2803 3919
rect 1131 3903 1135 3907
rect 2203 3907 2207 3911
rect 2347 3907 2351 3911
rect 2515 3907 2519 3911
rect 2691 3907 2695 3911
rect 2983 3915 2987 3919
rect 3175 3915 3179 3919
rect 3367 3915 3371 3919
rect 3559 3915 3563 3919
rect 3943 3916 3947 3920
rect 111 3896 115 3900
rect 279 3895 283 3899
rect 415 3895 419 3899
rect 567 3895 571 3899
rect 735 3895 739 3899
rect 911 3895 915 3899
rect 1095 3895 1099 3899
rect 355 3887 359 3891
rect 403 3887 407 3891
rect 643 3887 647 3891
rect 811 3887 815 3891
rect 987 3887 991 3891
rect 1047 3887 1051 3891
rect 1287 3895 1291 3899
rect 1479 3895 1483 3899
rect 1679 3895 1683 3899
rect 2007 3896 2011 3900
rect 2047 3899 2051 3903
rect 2875 3903 2879 3907
rect 3251 3907 3255 3911
rect 3443 3907 3447 3911
rect 3539 3907 3543 3911
rect 2127 3896 2131 3900
rect 2271 3896 2275 3900
rect 2439 3896 2443 3900
rect 2615 3896 2619 3900
rect 2799 3896 2803 3900
rect 2983 3896 2987 3900
rect 3175 3896 3179 3900
rect 3367 3896 3371 3900
rect 3559 3896 3563 3900
rect 3943 3899 3947 3903
rect 1371 3887 1375 3891
rect 111 3879 115 3883
rect 279 3876 283 3880
rect 415 3876 419 3880
rect 567 3876 571 3880
rect 735 3876 739 3880
rect 911 3876 915 3880
rect 1095 3876 1099 3880
rect 1287 3876 1291 3880
rect 1479 3876 1483 3880
rect 1679 3876 1683 3880
rect 2007 3879 2011 3883
rect 2047 3833 2051 3837
rect 2263 3836 2267 3840
rect 2375 3836 2379 3840
rect 2495 3836 2499 3840
rect 2631 3836 2635 3840
rect 2775 3836 2779 3840
rect 2919 3836 2923 3840
rect 3063 3836 3067 3840
rect 3207 3836 3211 3840
rect 3343 3836 3347 3840
rect 3471 3836 3475 3840
rect 3599 3836 3603 3840
rect 3727 3836 3731 3840
rect 3839 3836 3843 3840
rect 3943 3833 3947 3837
rect 2339 3827 2343 3831
rect 2451 3827 2455 3831
rect 2459 3827 2463 3831
rect 2579 3827 2583 3831
rect 2715 3827 2719 3831
rect 2995 3827 2999 3831
rect 3051 3827 3055 3831
rect 3275 3827 3279 3831
rect 3291 3827 3295 3831
rect 3427 3827 3431 3831
rect 3675 3827 3679 3831
rect 3803 3827 3807 3831
rect 3907 3827 3911 3831
rect 2047 3816 2051 3820
rect 2263 3817 2267 3821
rect 2375 3817 2379 3821
rect 2495 3817 2499 3821
rect 2631 3817 2635 3821
rect 2775 3817 2779 3821
rect 2919 3817 2923 3821
rect 3063 3817 3067 3821
rect 3207 3817 3211 3821
rect 3343 3817 3347 3821
rect 3471 3817 3475 3821
rect 3599 3817 3603 3821
rect 3727 3817 3731 3821
rect 3839 3817 3843 3821
rect 3943 3816 3947 3820
rect 111 3805 115 3809
rect 231 3808 235 3812
rect 335 3808 339 3812
rect 439 3808 443 3812
rect 535 3808 539 3812
rect 631 3808 635 3812
rect 727 3808 731 3812
rect 831 3808 835 3812
rect 935 3808 939 3812
rect 1039 3808 1043 3812
rect 1151 3808 1155 3812
rect 1263 3808 1267 3812
rect 1383 3808 1387 3812
rect 1503 3808 1507 3812
rect 1631 3808 1635 3812
rect 2007 3805 2011 3809
rect 303 3799 307 3803
rect 315 3799 319 3803
rect 515 3799 519 3803
rect 611 3799 615 3803
rect 707 3799 711 3803
rect 803 3799 807 3803
rect 907 3799 911 3803
rect 1011 3799 1015 3803
rect 1115 3799 1119 3803
rect 1227 3799 1231 3803
rect 1339 3799 1343 3803
rect 111 3788 115 3792
rect 231 3789 235 3793
rect 335 3789 339 3793
rect 439 3789 443 3793
rect 535 3789 539 3793
rect 631 3789 635 3793
rect 727 3789 731 3793
rect 831 3789 835 3793
rect 935 3789 939 3793
rect 1039 3789 1043 3793
rect 1151 3789 1155 3793
rect 1263 3789 1267 3793
rect 819 3783 823 3787
rect 1619 3799 1623 3803
rect 1707 3799 1711 3803
rect 2459 3803 2463 3807
rect 3675 3803 3679 3807
rect 2339 3795 2343 3799
rect 2579 3795 2583 3799
rect 2715 3795 2719 3799
rect 2875 3795 2879 3799
rect 2883 3795 2887 3799
rect 2995 3795 2999 3799
rect 3291 3795 3295 3799
rect 3427 3795 3431 3799
rect 3539 3795 3540 3799
rect 3540 3795 3543 3799
rect 3803 3795 3807 3799
rect 1383 3789 1387 3793
rect 1503 3789 1507 3793
rect 1631 3789 1635 3793
rect 2007 3788 2011 3792
rect 1047 3775 1051 3779
rect 315 3767 319 3771
rect 515 3767 519 3771
rect 611 3767 615 3771
rect 707 3767 711 3771
rect 803 3767 807 3771
rect 907 3767 911 3771
rect 1011 3767 1015 3771
rect 1115 3767 1119 3771
rect 1227 3767 1231 3771
rect 1339 3767 1343 3771
rect 1619 3767 1623 3771
rect 2155 3767 2159 3771
rect 2451 3767 2455 3771
rect 2555 3767 2559 3771
rect 2891 3767 2895 3771
rect 3003 3767 3007 3771
rect 3275 3767 3279 3771
rect 3299 3767 3303 3771
rect 3411 3767 3415 3771
rect 3747 3767 3751 3771
rect 3907 3767 3908 3771
rect 3908 3767 3911 3771
rect 223 3755 224 3759
rect 224 3755 227 3759
rect 259 3755 263 3759
rect 427 3755 431 3759
rect 819 3755 820 3759
rect 820 3755 823 3759
rect 907 3755 911 3759
rect 1079 3755 1083 3759
rect 1243 3755 1247 3759
rect 1555 3755 1559 3759
rect 2599 3759 2603 3763
rect 2047 3748 2051 3752
rect 2071 3747 2075 3751
rect 2183 3747 2187 3751
rect 2327 3747 2331 3751
rect 2479 3747 2483 3751
rect 2639 3747 2643 3751
rect 2807 3747 2811 3751
rect 2983 3747 2987 3751
rect 3159 3747 3163 3751
rect 3335 3747 3339 3751
rect 3511 3747 3515 3751
rect 3687 3747 3691 3751
rect 3839 3747 3843 3751
rect 3943 3748 3947 3752
rect 111 3736 115 3740
rect 159 3735 163 3739
rect 351 3735 355 3739
rect 551 3735 555 3739
rect 751 3735 755 3739
rect 959 3735 963 3739
rect 1167 3735 1171 3739
rect 1383 3735 1387 3739
rect 1607 3735 1611 3739
rect 2007 3736 2011 3740
rect 2155 3739 2159 3743
rect 2555 3739 2559 3743
rect 2599 3739 2603 3743
rect 2883 3739 2887 3743
rect 2891 3739 2895 3743
rect 3299 3739 3303 3743
rect 3411 3739 3415 3743
rect 259 3727 263 3731
rect 427 3727 431 3731
rect 907 3727 911 3731
rect 1079 3727 1083 3731
rect 1243 3727 1247 3731
rect 1347 3727 1351 3731
rect 2047 3731 2051 3735
rect 2071 3728 2075 3732
rect 2139 3731 2143 3735
rect 3587 3735 3591 3739
rect 2183 3728 2187 3732
rect 2327 3728 2331 3732
rect 2479 3728 2483 3732
rect 2639 3728 2643 3732
rect 2807 3728 2811 3732
rect 2983 3728 2987 3732
rect 3159 3728 3163 3732
rect 3335 3728 3339 3732
rect 3511 3728 3515 3732
rect 3687 3728 3691 3732
rect 3839 3728 3843 3732
rect 3907 3731 3911 3735
rect 3943 3731 3947 3735
rect 111 3719 115 3723
rect 159 3716 163 3720
rect 351 3716 355 3720
rect 551 3716 555 3720
rect 751 3716 755 3720
rect 959 3716 963 3720
rect 1167 3716 1171 3720
rect 1383 3716 1387 3720
rect 1607 3716 1611 3720
rect 2007 3719 2011 3723
rect 2047 3653 2051 3657
rect 2071 3656 2075 3660
rect 2199 3656 2203 3660
rect 2367 3656 2371 3660
rect 2551 3656 2555 3660
rect 2735 3656 2739 3660
rect 2927 3656 2931 3660
rect 3111 3656 3115 3660
rect 3295 3656 3299 3660
rect 3479 3656 3483 3660
rect 3671 3656 3675 3660
rect 3839 3656 3843 3660
rect 111 3645 115 3649
rect 151 3648 155 3652
rect 383 3648 387 3652
rect 615 3648 619 3652
rect 839 3648 843 3652
rect 1055 3648 1059 3652
rect 1263 3648 1267 3652
rect 1479 3648 1483 3652
rect 3943 3653 3947 3657
rect 1695 3648 1699 3652
rect 2007 3645 2011 3649
rect 2147 3647 2151 3651
rect 2275 3647 2279 3651
rect 2443 3647 2447 3651
rect 2627 3647 2631 3651
rect 223 3639 227 3643
rect 235 3639 239 3643
rect 467 3639 471 3643
rect 1039 3639 1043 3643
rect 1131 3639 1135 3643
rect 1339 3639 1343 3643
rect 1555 3639 1559 3643
rect 1563 3639 1567 3643
rect 2047 3636 2051 3640
rect 2071 3637 2075 3641
rect 2199 3637 2203 3641
rect 2367 3637 2371 3641
rect 2551 3637 2555 3641
rect 111 3628 115 3632
rect 151 3629 155 3633
rect 383 3629 387 3633
rect 615 3629 619 3633
rect 839 3629 843 3633
rect 1055 3629 1059 3633
rect 1263 3629 1267 3633
rect 1479 3629 1483 3633
rect 1695 3629 1699 3633
rect 2007 3628 2011 3632
rect 2171 3631 2175 3635
rect 3003 3647 3007 3651
rect 3187 3647 3191 3651
rect 3195 3647 3199 3651
rect 3379 3647 3383 3651
rect 3747 3647 3751 3651
rect 3915 3647 3919 3651
rect 2735 3637 2739 3641
rect 2927 3637 2931 3641
rect 3111 3637 3115 3641
rect 3295 3637 3299 3641
rect 3479 3637 3483 3641
rect 3671 3637 3675 3641
rect 3839 3637 3843 3641
rect 3943 3636 3947 3640
rect 235 3607 239 3611
rect 467 3607 471 3611
rect 683 3607 684 3611
rect 684 3607 687 3611
rect 1347 3615 1351 3619
rect 2139 3615 2140 3619
rect 2140 3615 2143 3619
rect 2147 3615 2151 3619
rect 2275 3615 2279 3619
rect 2443 3615 2447 3619
rect 2627 3615 2631 3619
rect 3195 3615 3199 3619
rect 3379 3615 3383 3619
rect 3587 3615 3591 3619
rect 3715 3615 3719 3619
rect 3907 3615 3908 3619
rect 3908 3615 3911 3619
rect 1039 3607 1043 3611
rect 1131 3607 1135 3611
rect 1563 3607 1567 3611
rect 1763 3607 1764 3611
rect 1764 3607 1767 3611
rect 2171 3599 2172 3603
rect 2172 3599 2175 3603
rect 2179 3599 2183 3603
rect 2355 3599 2359 3603
rect 2583 3599 2587 3603
rect 2979 3599 2983 3603
rect 3187 3599 3191 3603
rect 3331 3599 3335 3603
rect 3523 3599 3527 3603
rect 3915 3599 3919 3603
rect 243 3591 247 3595
rect 435 3591 439 3595
rect 635 3591 639 3595
rect 1299 3591 1303 3595
rect 1339 3591 1343 3595
rect 1755 3591 1756 3595
rect 1756 3591 1759 3595
rect 2047 3580 2051 3584
rect 2103 3579 2107 3583
rect 2279 3579 2283 3583
rect 2471 3579 2475 3583
rect 2671 3579 2675 3583
rect 2871 3579 2875 3583
rect 3063 3579 3067 3583
rect 3255 3579 3259 3583
rect 3447 3579 3451 3583
rect 3639 3579 3643 3583
rect 3839 3579 3843 3583
rect 3943 3580 3947 3584
rect 111 3572 115 3576
rect 167 3571 171 3575
rect 359 3571 363 3575
rect 559 3571 563 3575
rect 775 3571 779 3575
rect 991 3571 995 3575
rect 1215 3571 1219 3575
rect 1447 3571 1451 3575
rect 1687 3571 1691 3575
rect 2007 3572 2011 3576
rect 2179 3571 2183 3575
rect 2355 3571 2359 3575
rect 2583 3571 2587 3575
rect 2599 3571 2603 3575
rect 3331 3571 3335 3575
rect 3523 3571 3527 3575
rect 3715 3571 3719 3575
rect 243 3563 247 3567
rect 435 3563 439 3567
rect 635 3563 639 3567
rect 683 3563 687 3567
rect 111 3555 115 3559
rect 1067 3559 1071 3563
rect 1299 3563 1303 3567
rect 1763 3563 1767 3567
rect 2047 3563 2051 3567
rect 3915 3567 3919 3571
rect 2103 3560 2107 3564
rect 2279 3560 2283 3564
rect 2471 3560 2475 3564
rect 2671 3560 2675 3564
rect 2871 3560 2875 3564
rect 3063 3560 3067 3564
rect 3255 3560 3259 3564
rect 3447 3560 3451 3564
rect 3639 3560 3643 3564
rect 3839 3560 3843 3564
rect 3943 3563 3947 3567
rect 167 3552 171 3556
rect 359 3552 363 3556
rect 559 3552 563 3556
rect 775 3552 779 3556
rect 991 3552 995 3556
rect 1215 3552 1219 3556
rect 1447 3552 1451 3556
rect 1687 3552 1691 3556
rect 2007 3555 2011 3559
rect 2047 3493 2051 3497
rect 2327 3496 2331 3500
rect 2447 3496 2451 3500
rect 2583 3496 2587 3500
rect 2735 3496 2739 3500
rect 2911 3496 2915 3500
rect 3111 3496 3115 3500
rect 3335 3496 3339 3500
rect 3567 3496 3571 3500
rect 3807 3496 3811 3500
rect 3943 3493 3947 3497
rect 111 3481 115 3485
rect 295 3484 299 3488
rect 431 3484 435 3488
rect 583 3484 587 3488
rect 743 3484 747 3488
rect 911 3484 915 3488
rect 1079 3484 1083 3488
rect 1247 3484 1251 3488
rect 1423 3484 1427 3488
rect 1599 3484 1603 3488
rect 1775 3484 1779 3488
rect 2403 3487 2407 3491
rect 2523 3487 2527 3491
rect 2711 3487 2715 3491
rect 2007 3481 2011 3485
rect 379 3475 383 3479
rect 515 3475 519 3479
rect 667 3475 671 3479
rect 827 3475 831 3479
rect 1155 3475 1159 3479
rect 1323 3475 1327 3479
rect 1499 3475 1503 3479
rect 1739 3475 1743 3479
rect 1755 3475 1759 3479
rect 2047 3476 2051 3480
rect 2327 3477 2331 3481
rect 2447 3477 2451 3481
rect 2583 3477 2587 3481
rect 2515 3471 2519 3475
rect 2979 3487 2983 3491
rect 2995 3487 2999 3491
rect 3195 3487 3199 3491
rect 3419 3487 3423 3491
rect 3875 3487 3879 3491
rect 2735 3477 2739 3481
rect 2911 3477 2915 3481
rect 3111 3477 3115 3481
rect 3335 3477 3339 3481
rect 3567 3477 3571 3481
rect 3807 3477 3811 3481
rect 3943 3476 3947 3480
rect 111 3464 115 3468
rect 295 3465 299 3469
rect 431 3465 435 3469
rect 583 3465 587 3469
rect 743 3465 747 3469
rect 911 3465 915 3469
rect 1079 3465 1083 3469
rect 1247 3465 1251 3469
rect 1423 3465 1427 3469
rect 1599 3465 1603 3469
rect 1775 3465 1779 3469
rect 2007 3464 2011 3468
rect 2599 3463 2603 3467
rect 2403 3455 2407 3459
rect 2523 3455 2527 3459
rect 2711 3455 2715 3459
rect 2995 3455 2999 3459
rect 3195 3455 3199 3459
rect 3419 3455 3423 3459
rect 3643 3455 3647 3459
rect 3915 3455 3919 3459
rect 379 3443 383 3447
rect 515 3443 519 3447
rect 667 3443 671 3447
rect 827 3443 831 3447
rect 1035 3443 1039 3447
rect 1067 3443 1071 3447
rect 1155 3443 1159 3447
rect 1323 3443 1327 3447
rect 1715 3443 1719 3447
rect 1739 3443 1743 3447
rect 2515 3443 2516 3447
rect 2516 3443 2519 3447
rect 2523 3443 2527 3447
rect 2627 3443 2631 3447
rect 2751 3443 2755 3447
rect 2851 3443 2855 3447
rect 3123 3443 3127 3447
rect 3283 3443 3287 3447
rect 3459 3443 3463 3447
rect 3875 3443 3879 3447
rect 3259 3435 3263 3439
rect 2047 3424 2051 3428
rect 2447 3423 2451 3427
rect 2551 3423 2555 3427
rect 2663 3423 2667 3427
rect 2775 3423 2779 3427
rect 2903 3423 2907 3427
rect 3047 3423 3051 3427
rect 3207 3423 3211 3427
rect 3383 3423 3387 3427
rect 3567 3423 3571 3427
rect 3751 3423 3755 3427
rect 3943 3424 3947 3428
rect 619 3411 623 3415
rect 627 3411 631 3415
rect 723 3411 727 3415
rect 875 3411 879 3415
rect 1499 3411 1503 3415
rect 1723 3411 1727 3415
rect 1899 3411 1903 3415
rect 2523 3415 2527 3419
rect 2627 3415 2631 3419
rect 2751 3415 2755 3419
rect 2851 3415 2855 3419
rect 2047 3407 2051 3411
rect 2979 3411 2983 3415
rect 3123 3415 3127 3419
rect 3283 3415 3287 3419
rect 3459 3415 3463 3419
rect 3643 3415 3647 3419
rect 3827 3411 3831 3415
rect 2447 3404 2451 3408
rect 2551 3404 2555 3408
rect 2663 3404 2667 3408
rect 2775 3404 2779 3408
rect 2903 3404 2907 3408
rect 3047 3404 3051 3408
rect 3207 3404 3211 3408
rect 3383 3404 3387 3408
rect 3567 3404 3571 3408
rect 3751 3404 3755 3408
rect 3943 3407 3947 3411
rect 111 3392 115 3396
rect 495 3391 499 3395
rect 647 3391 651 3395
rect 799 3391 803 3395
rect 959 3391 963 3395
rect 1127 3391 1131 3395
rect 1295 3391 1299 3395
rect 1463 3391 1467 3395
rect 1639 3391 1643 3395
rect 1815 3391 1819 3395
rect 2007 3392 2011 3396
rect 627 3383 631 3387
rect 723 3383 727 3387
rect 875 3383 879 3387
rect 1035 3383 1039 3387
rect 111 3375 115 3379
rect 1203 3379 1207 3383
rect 1715 3383 1719 3387
rect 1723 3383 1727 3387
rect 495 3372 499 3376
rect 647 3372 651 3376
rect 799 3372 803 3376
rect 959 3372 963 3376
rect 1127 3372 1131 3376
rect 1295 3372 1299 3376
rect 1463 3372 1467 3376
rect 1639 3372 1643 3376
rect 1815 3372 1819 3376
rect 2007 3375 2011 3379
rect 2047 3329 2051 3333
rect 2567 3332 2571 3336
rect 2719 3332 2723 3336
rect 2871 3332 2875 3336
rect 3023 3332 3027 3336
rect 3175 3332 3179 3336
rect 3327 3332 3331 3336
rect 3479 3332 3483 3336
rect 3631 3332 3635 3336
rect 3783 3332 3787 3336
rect 3943 3329 3947 3333
rect 2643 3323 2647 3327
rect 2651 3323 2655 3327
rect 2803 3323 2807 3327
rect 2955 3323 2959 3327
rect 3251 3323 3255 3327
rect 3259 3323 3263 3327
rect 3563 3323 3567 3327
rect 3715 3323 3719 3327
rect 2047 3312 2051 3316
rect 2567 3313 2571 3317
rect 2719 3313 2723 3317
rect 2871 3313 2875 3317
rect 3023 3313 3027 3317
rect 3175 3313 3179 3317
rect 3327 3313 3331 3317
rect 3479 3313 3483 3317
rect 3631 3313 3635 3317
rect 3783 3313 3787 3317
rect 3943 3312 3947 3316
rect 111 3297 115 3301
rect 135 3300 139 3304
rect 295 3300 299 3304
rect 479 3300 483 3304
rect 671 3300 675 3304
rect 863 3300 867 3304
rect 1055 3300 1059 3304
rect 1247 3300 1251 3304
rect 1439 3300 1443 3304
rect 1631 3300 1635 3304
rect 1823 3300 1827 3304
rect 2007 3297 2011 3301
rect 211 3291 215 3295
rect 371 3291 375 3295
rect 387 3291 391 3295
rect 619 3291 623 3295
rect 755 3291 759 3295
rect 1131 3291 1135 3295
rect 1323 3291 1327 3295
rect 1339 3291 1343 3295
rect 1779 3291 1783 3295
rect 1899 3291 1903 3295
rect 2651 3291 2655 3295
rect 2803 3291 2807 3295
rect 2955 3291 2959 3295
rect 2979 3291 2983 3295
rect 3195 3291 3199 3295
rect 3251 3291 3255 3295
rect 3563 3291 3567 3295
rect 3715 3291 3719 3295
rect 3827 3291 3831 3295
rect 111 3280 115 3284
rect 135 3281 139 3285
rect 295 3281 299 3285
rect 479 3281 483 3285
rect 671 3281 675 3285
rect 863 3281 867 3285
rect 1055 3281 1059 3285
rect 1247 3281 1251 3285
rect 1439 3281 1443 3285
rect 1631 3281 1635 3285
rect 1823 3281 1827 3285
rect 2007 3280 2011 3284
rect 2491 3275 2495 3279
rect 2643 3275 2647 3279
rect 2763 3275 2767 3279
rect 2907 3275 2911 3279
rect 3375 3275 3379 3279
rect 3495 3275 3499 3279
rect 3579 3275 3583 3279
rect 3699 3275 3703 3279
rect 3819 3275 3823 3279
rect 211 3259 215 3263
rect 371 3259 375 3263
rect 755 3259 759 3263
rect 987 3259 991 3263
rect 1339 3267 1343 3271
rect 2927 3267 2931 3271
rect 1203 3259 1207 3263
rect 1323 3259 1327 3263
rect 1707 3259 1711 3263
rect 1779 3259 1783 3263
rect 2047 3256 2051 3260
rect 2415 3255 2419 3259
rect 2551 3255 2555 3259
rect 2687 3255 2691 3259
rect 2831 3255 2835 3259
rect 2975 3255 2979 3259
rect 3119 3255 3123 3259
rect 3255 3255 3259 3259
rect 3383 3255 3387 3259
rect 3503 3255 3507 3259
rect 3623 3255 3627 3259
rect 3743 3255 3747 3259
rect 3839 3255 3843 3259
rect 3943 3256 3947 3260
rect 387 3243 388 3247
rect 388 3243 391 3247
rect 679 3243 683 3247
rect 687 3243 691 3247
rect 795 3243 799 3247
rect 1131 3243 1135 3247
rect 1171 3243 1175 3247
rect 1347 3243 1351 3247
rect 1651 3243 1655 3247
rect 1699 3243 1703 3247
rect 2491 3247 2495 3251
rect 2047 3239 2051 3243
rect 2627 3243 2631 3247
rect 2763 3247 2767 3251
rect 2907 3247 2911 3251
rect 2927 3247 2931 3251
rect 3195 3247 3199 3251
rect 3495 3247 3499 3251
rect 3579 3247 3583 3251
rect 3699 3247 3703 3251
rect 3819 3247 3823 3251
rect 3915 3243 3919 3247
rect 2415 3236 2419 3240
rect 2551 3236 2555 3240
rect 2687 3236 2691 3240
rect 2831 3236 2835 3240
rect 2975 3236 2979 3240
rect 3119 3236 3123 3240
rect 3255 3236 3259 3240
rect 3383 3236 3387 3240
rect 3503 3236 3507 3240
rect 3623 3236 3627 3240
rect 3743 3236 3747 3240
rect 3839 3236 3843 3240
rect 3943 3239 3947 3243
rect 111 3224 115 3228
rect 135 3223 139 3227
rect 319 3223 323 3227
rect 519 3223 523 3227
rect 719 3223 723 3227
rect 911 3223 915 3227
rect 1095 3223 1099 3227
rect 1271 3223 1275 3227
rect 1447 3223 1451 3227
rect 1623 3223 1627 3227
rect 1799 3223 1803 3227
rect 2007 3224 2011 3228
rect 111 3207 115 3211
rect 211 3211 215 3215
rect 687 3215 691 3219
rect 795 3215 799 3219
rect 987 3215 991 3219
rect 1171 3215 1175 3219
rect 1347 3215 1351 3219
rect 1523 3211 1527 3215
rect 1699 3215 1703 3219
rect 1707 3215 1711 3219
rect 135 3204 139 3208
rect 319 3204 323 3208
rect 519 3204 523 3208
rect 719 3204 723 3208
rect 911 3204 915 3208
rect 1095 3204 1099 3208
rect 1271 3204 1275 3208
rect 1447 3204 1451 3208
rect 1623 3204 1627 3208
rect 1799 3204 1803 3208
rect 2007 3207 2011 3211
rect 3375 3171 3379 3175
rect 2047 3161 2051 3165
rect 2247 3164 2251 3168
rect 2399 3164 2403 3168
rect 2559 3164 2563 3168
rect 2727 3164 2731 3168
rect 2903 3164 2907 3168
rect 3079 3164 3083 3168
rect 3263 3164 3267 3168
rect 3447 3164 3451 3168
rect 2323 3155 2327 3159
rect 2331 3155 2335 3159
rect 2635 3155 2639 3159
rect 2803 3155 2807 3159
rect 3155 3155 3159 3159
rect 3339 3155 3343 3159
rect 3523 3155 3527 3159
rect 3631 3164 3635 3168
rect 3815 3164 3819 3168
rect 3943 3161 3947 3165
rect 3891 3155 3895 3159
rect 2047 3144 2051 3148
rect 2247 3145 2251 3149
rect 2399 3145 2403 3149
rect 2559 3145 2563 3149
rect 2727 3145 2731 3149
rect 2903 3145 2907 3149
rect 3079 3145 3083 3149
rect 3263 3145 3267 3149
rect 3447 3145 3451 3149
rect 3631 3145 3635 3149
rect 3815 3145 3819 3149
rect 3943 3144 3947 3148
rect 111 3133 115 3137
rect 143 3136 147 3140
rect 343 3136 347 3140
rect 543 3136 547 3140
rect 743 3136 747 3140
rect 927 3136 931 3140
rect 1103 3136 1107 3140
rect 1263 3136 1267 3140
rect 1423 3136 1427 3140
rect 1575 3136 1579 3140
rect 1735 3136 1739 3140
rect 2007 3133 2011 3137
rect 219 3127 223 3131
rect 419 3127 423 3131
rect 631 3127 635 3131
rect 679 3127 683 3131
rect 827 3127 831 3131
rect 1179 3127 1183 3131
rect 1187 3127 1191 3131
rect 1347 3127 1351 3131
rect 1651 3127 1655 3131
rect 1659 3127 1663 3131
rect 2331 3123 2335 3127
rect 2627 3123 2628 3127
rect 2628 3123 2631 3127
rect 2635 3123 2639 3127
rect 2803 3123 2807 3127
rect 3155 3123 3159 3127
rect 3339 3123 3343 3127
rect 3523 3123 3527 3127
rect 3915 3123 3919 3127
rect 111 3116 115 3120
rect 143 3117 147 3121
rect 343 3117 347 3121
rect 543 3117 547 3121
rect 743 3117 747 3121
rect 927 3117 931 3121
rect 1103 3117 1107 3121
rect 1263 3117 1267 3121
rect 1423 3117 1427 3121
rect 1575 3117 1579 3121
rect 1735 3117 1739 3121
rect 2007 3116 2011 3120
rect 3603 3115 3607 3119
rect 2155 3107 2159 3111
rect 2323 3107 2327 3111
rect 2451 3107 2455 3111
rect 2603 3107 2607 3111
rect 2923 3107 2924 3111
rect 2924 3107 2927 3111
rect 2931 3107 2935 3111
rect 3115 3107 3119 3111
rect 3307 3107 3311 3111
rect 3507 3107 3511 3111
rect 3891 3107 3895 3111
rect 211 3095 212 3099
rect 212 3095 215 3099
rect 219 3095 223 3099
rect 419 3095 423 3099
rect 827 3095 831 3099
rect 1051 3095 1055 3099
rect 1187 3095 1191 3099
rect 1347 3095 1351 3099
rect 1523 3095 1527 3099
rect 1659 3095 1663 3099
rect 1843 3095 1847 3099
rect 2659 3099 2663 3103
rect 2047 3088 2051 3092
rect 387 3083 391 3087
rect 631 3083 635 3087
rect 859 3083 863 3087
rect 875 3083 879 3087
rect 1179 3083 1183 3087
rect 1219 3083 1223 3087
rect 1379 3083 1383 3087
rect 1531 3083 1535 3087
rect 1683 3083 1687 3087
rect 2079 3087 2083 3091
rect 2223 3087 2227 3091
rect 2375 3087 2379 3091
rect 2527 3087 2531 3091
rect 2687 3087 2691 3091
rect 2855 3087 2859 3091
rect 3039 3087 3043 3091
rect 3231 3087 3235 3091
rect 3431 3087 3435 3091
rect 3639 3087 3643 3091
rect 3839 3087 3843 3091
rect 3943 3088 3947 3092
rect 559 3075 563 3079
rect 2155 3079 2159 3083
rect 2047 3071 2051 3075
rect 2299 3075 2303 3079
rect 2451 3079 2455 3083
rect 2603 3079 2607 3083
rect 2659 3079 2663 3083
rect 2931 3079 2935 3083
rect 3115 3079 3119 3083
rect 3307 3079 3311 3083
rect 3507 3079 3511 3083
rect 3603 3079 3607 3083
rect 3915 3075 3919 3079
rect 111 3064 115 3068
rect 263 3063 267 3067
rect 439 3063 443 3067
rect 615 3063 619 3067
rect 799 3063 803 3067
rect 975 3063 979 3067
rect 1143 3063 1147 3067
rect 1303 3063 1307 3067
rect 1455 3063 1459 3067
rect 1607 3063 1611 3067
rect 1767 3063 1771 3067
rect 2007 3064 2011 3068
rect 2079 3068 2083 3072
rect 2223 3068 2227 3072
rect 2375 3068 2379 3072
rect 2527 3068 2531 3072
rect 2687 3068 2691 3072
rect 2855 3068 2859 3072
rect 3039 3068 3043 3072
rect 3231 3068 3235 3072
rect 3431 3068 3435 3072
rect 3639 3068 3643 3072
rect 3839 3068 3843 3072
rect 3943 3071 3947 3075
rect 387 3055 391 3059
rect 111 3047 115 3051
rect 515 3051 519 3055
rect 559 3055 563 3059
rect 875 3055 879 3059
rect 1051 3055 1055 3059
rect 1219 3055 1223 3059
rect 1379 3055 1383 3059
rect 1531 3055 1535 3059
rect 1683 3055 1687 3059
rect 1843 3055 1847 3059
rect 263 3044 267 3048
rect 439 3044 443 3048
rect 615 3044 619 3048
rect 799 3044 803 3048
rect 975 3044 979 3048
rect 1143 3044 1147 3048
rect 1303 3044 1307 3048
rect 1455 3044 1459 3048
rect 1607 3044 1611 3048
rect 1767 3044 1771 3048
rect 2007 3047 2011 3051
rect 2923 3007 2927 3011
rect 2047 2997 2051 3001
rect 2071 3000 2075 3004
rect 2183 3000 2187 3004
rect 2327 3000 2331 3004
rect 2479 3000 2483 3004
rect 2655 3000 2659 3004
rect 2855 3000 2859 3004
rect 3087 3000 3091 3004
rect 3335 3000 3339 3004
rect 2139 2991 2143 2995
rect 2155 2991 2159 2995
rect 2403 2991 2407 2995
rect 2555 2991 2559 2995
rect 2599 2991 2603 2995
rect 2931 2991 2935 2995
rect 3163 2991 3167 2995
rect 3411 2991 3415 2995
rect 3599 3000 3603 3004
rect 3839 3000 3843 3004
rect 3943 2997 3947 3001
rect 3907 2991 3911 2995
rect 2047 2980 2051 2984
rect 2071 2981 2075 2985
rect 2183 2981 2187 2985
rect 2327 2981 2331 2985
rect 2479 2981 2483 2985
rect 2655 2981 2659 2985
rect 2855 2981 2859 2985
rect 3087 2981 3091 2985
rect 3335 2981 3339 2985
rect 3599 2981 3603 2985
rect 3839 2981 3843 2985
rect 3943 2980 3947 2984
rect 111 2957 115 2961
rect 343 2960 347 2964
rect 439 2960 443 2964
rect 543 2960 547 2964
rect 655 2960 659 2964
rect 783 2960 787 2964
rect 935 2960 939 2964
rect 1103 2960 1107 2964
rect 1295 2960 1299 2964
rect 1495 2960 1499 2964
rect 1711 2960 1715 2964
rect 1903 2960 1907 2964
rect 2007 2957 2011 2961
rect 2155 2959 2159 2963
rect 2599 2967 2603 2971
rect 2299 2959 2303 2963
rect 2403 2959 2407 2963
rect 2555 2959 2559 2963
rect 2931 2959 2935 2963
rect 3163 2959 3167 2963
rect 3411 2959 3415 2963
rect 3915 2959 3919 2963
rect 275 2951 279 2955
rect 427 2951 431 2955
rect 731 2951 735 2955
rect 859 2951 863 2955
rect 1011 2951 1015 2955
rect 1179 2951 1183 2955
rect 1371 2951 1375 2955
rect 1571 2951 1575 2955
rect 1787 2951 1791 2955
rect 1795 2951 1799 2955
rect 3363 2951 3367 2955
rect 111 2940 115 2944
rect 343 2941 347 2945
rect 439 2941 443 2945
rect 543 2941 547 2945
rect 655 2941 659 2945
rect 783 2941 787 2945
rect 935 2941 939 2945
rect 1103 2941 1107 2945
rect 1295 2941 1299 2945
rect 1495 2941 1499 2945
rect 1711 2941 1715 2945
rect 1903 2941 1907 2945
rect 2007 2940 2011 2944
rect 2139 2943 2140 2947
rect 2140 2943 2143 2947
rect 2331 2939 2335 2943
rect 2339 2943 2343 2947
rect 2563 2943 2567 2947
rect 2811 2943 2815 2947
rect 3075 2943 3079 2947
rect 3355 2943 3359 2947
rect 3907 2943 3908 2947
rect 3908 2943 3911 2947
rect 2047 2924 2051 2928
rect 427 2919 431 2923
rect 515 2919 519 2923
rect 643 2919 647 2923
rect 731 2919 735 2923
rect 991 2919 995 2923
rect 1011 2919 1015 2923
rect 1179 2919 1183 2923
rect 1371 2919 1375 2923
rect 1795 2919 1799 2923
rect 2071 2923 2075 2927
rect 2263 2923 2267 2927
rect 2487 2923 2491 2927
rect 2735 2923 2739 2927
rect 2999 2923 3003 2927
rect 3279 2923 3283 2927
rect 3567 2923 3571 2927
rect 3839 2923 3843 2927
rect 3943 2924 3947 2928
rect 2339 2915 2343 2919
rect 2563 2915 2567 2919
rect 2811 2915 2815 2919
rect 3075 2915 3079 2919
rect 3355 2915 3359 2919
rect 3363 2915 3367 2919
rect 275 2907 276 2911
rect 276 2907 279 2911
rect 283 2907 287 2911
rect 403 2907 407 2911
rect 771 2907 772 2911
rect 772 2907 775 2911
rect 947 2907 951 2911
rect 975 2907 979 2911
rect 1251 2907 1255 2911
rect 1439 2907 1443 2911
rect 1571 2907 1575 2911
rect 1787 2907 1791 2911
rect 1803 2907 1807 2911
rect 2047 2907 2051 2911
rect 3915 2911 3919 2915
rect 2071 2904 2075 2908
rect 2263 2904 2267 2908
rect 2487 2904 2491 2908
rect 2735 2904 2739 2908
rect 2999 2904 3003 2908
rect 3279 2904 3283 2908
rect 3567 2904 3571 2908
rect 3839 2904 3843 2908
rect 3943 2907 3947 2911
rect 111 2888 115 2892
rect 207 2887 211 2891
rect 327 2887 331 2891
rect 447 2887 451 2891
rect 575 2887 579 2891
rect 283 2879 287 2883
rect 403 2879 407 2883
rect 643 2883 647 2887
rect 703 2887 707 2891
rect 847 2887 851 2891
rect 999 2887 1003 2891
rect 1167 2887 1171 2891
rect 1351 2887 1355 2891
rect 1535 2887 1539 2891
rect 1727 2887 1731 2891
rect 1903 2887 1907 2891
rect 2007 2888 2011 2892
rect 111 2871 115 2875
rect 523 2875 527 2879
rect 975 2879 979 2883
rect 991 2879 995 2883
rect 1243 2875 1247 2879
rect 1251 2879 1255 2883
rect 1439 2879 1443 2883
rect 1803 2879 1807 2883
rect 1819 2879 1823 2883
rect 207 2868 211 2872
rect 327 2868 331 2872
rect 447 2868 451 2872
rect 575 2868 579 2872
rect 703 2868 707 2872
rect 847 2868 851 2872
rect 999 2868 1003 2872
rect 1167 2868 1171 2872
rect 1351 2868 1355 2872
rect 1535 2868 1539 2872
rect 1727 2868 1731 2872
rect 1903 2868 1907 2872
rect 2007 2871 2011 2875
rect 2047 2833 2051 2837
rect 2331 2827 2335 2831
rect 2671 2836 2675 2840
rect 2887 2836 2891 2840
rect 2747 2827 2751 2831
rect 2963 2827 2967 2831
rect 3095 2836 3099 2840
rect 3287 2836 3291 2840
rect 3479 2836 3483 2840
rect 3671 2836 3675 2840
rect 3839 2836 3843 2840
rect 3943 2833 3947 2837
rect 3355 2827 3359 2831
rect 3371 2827 3375 2831
rect 3755 2827 3759 2831
rect 2047 2816 2051 2820
rect 2671 2817 2675 2821
rect 2887 2817 2891 2821
rect 3095 2817 3099 2821
rect 3287 2817 3291 2821
rect 3479 2817 3483 2821
rect 3671 2817 3675 2821
rect 3839 2817 3843 2821
rect 3943 2816 3947 2820
rect 111 2801 115 2805
rect 135 2804 139 2808
rect 247 2804 251 2808
rect 399 2804 403 2808
rect 551 2804 555 2808
rect 711 2804 715 2808
rect 879 2804 883 2808
rect 1047 2804 1051 2808
rect 1223 2804 1227 2808
rect 1399 2804 1403 2808
rect 1575 2804 1579 2808
rect 1751 2804 1755 2808
rect 1903 2804 1907 2808
rect 2007 2801 2011 2805
rect 203 2795 207 2799
rect 219 2795 223 2799
rect 379 2795 383 2799
rect 683 2795 687 2799
rect 779 2795 783 2799
rect 947 2795 951 2799
rect 963 2795 967 2799
rect 1299 2795 1303 2799
rect 1475 2795 1479 2799
rect 1651 2795 1655 2799
rect 1827 2795 1831 2799
rect 2683 2795 2687 2799
rect 2747 2795 2751 2799
rect 2963 2795 2967 2799
rect 3371 2795 3375 2799
rect 3523 2795 3527 2799
rect 3755 2795 3759 2799
rect 3907 2795 3908 2799
rect 3908 2795 3911 2799
rect 111 2784 115 2788
rect 135 2785 139 2789
rect 247 2785 251 2789
rect 399 2785 403 2789
rect 551 2785 555 2789
rect 711 2785 715 2789
rect 879 2785 883 2789
rect 1047 2785 1051 2789
rect 1223 2785 1227 2789
rect 1399 2785 1403 2789
rect 1575 2785 1579 2789
rect 1751 2785 1755 2789
rect 1903 2785 1907 2789
rect 2007 2784 2011 2788
rect 2147 2783 2151 2787
rect 2411 2783 2412 2787
rect 2412 2783 2415 2787
rect 2419 2783 2423 2787
rect 2555 2783 2559 2787
rect 2823 2783 2827 2787
rect 3131 2783 3135 2787
rect 3355 2783 3359 2787
rect 3419 2783 3423 2787
rect 2923 2775 2927 2779
rect 3531 2775 3535 2779
rect 3819 2783 3823 2787
rect 3827 2775 3831 2779
rect 219 2763 223 2767
rect 379 2763 383 2767
rect 523 2763 527 2767
rect 651 2763 655 2767
rect 683 2763 687 2767
rect 963 2763 967 2767
rect 1163 2763 1167 2767
rect 1243 2763 1247 2767
rect 1299 2763 1303 2767
rect 1475 2763 1479 2767
rect 1819 2763 1820 2767
rect 1820 2763 1823 2767
rect 1827 2763 1831 2767
rect 2047 2764 2051 2768
rect 2071 2763 2075 2767
rect 2199 2763 2203 2767
rect 2343 2763 2347 2767
rect 2479 2763 2483 2767
rect 2607 2763 2611 2767
rect 2727 2763 2731 2767
rect 2839 2763 2843 2767
rect 2943 2763 2947 2767
rect 3047 2763 3051 2767
rect 3143 2763 3147 2767
rect 3239 2763 3243 2767
rect 3343 2763 3347 2767
rect 3447 2763 3451 2767
rect 3551 2763 3555 2767
rect 3647 2763 3651 2767
rect 3743 2763 3747 2767
rect 3839 2763 3843 2767
rect 3943 2764 3947 2768
rect 2147 2755 2151 2759
rect 2163 2755 2167 2759
rect 2419 2755 2423 2759
rect 2555 2755 2559 2759
rect 2683 2755 2687 2759
rect 2823 2755 2827 2759
rect 203 2743 204 2747
rect 204 2743 207 2747
rect 211 2743 215 2747
rect 331 2743 335 2747
rect 827 2743 831 2747
rect 1019 2743 1023 2747
rect 1055 2743 1059 2747
rect 1339 2743 1343 2747
rect 1651 2743 1655 2747
rect 2047 2747 2051 2751
rect 2915 2751 2919 2755
rect 2923 2755 2927 2759
rect 3131 2755 3135 2759
rect 3419 2755 3423 2759
rect 3523 2755 3527 2759
rect 3531 2755 3535 2759
rect 3819 2755 3823 2759
rect 3827 2755 3831 2759
rect 2071 2744 2075 2748
rect 2199 2744 2203 2748
rect 2343 2744 2347 2748
rect 2479 2744 2483 2748
rect 2607 2744 2611 2748
rect 2727 2744 2731 2748
rect 2839 2744 2843 2748
rect 2943 2744 2947 2748
rect 3047 2744 3051 2748
rect 3143 2744 3147 2748
rect 3239 2744 3243 2748
rect 3343 2744 3347 2748
rect 3447 2744 3451 2748
rect 3551 2744 3555 2748
rect 3647 2744 3651 2748
rect 3743 2744 3747 2748
rect 3839 2744 3843 2748
rect 3943 2747 3947 2751
rect 111 2724 115 2728
rect 135 2723 139 2727
rect 255 2723 259 2727
rect 407 2723 411 2727
rect 575 2723 579 2727
rect 743 2723 747 2727
rect 919 2723 923 2727
rect 1087 2723 1091 2727
rect 1255 2723 1259 2727
rect 1423 2723 1427 2727
rect 1599 2723 1603 2727
rect 2007 2724 2011 2728
rect 211 2715 215 2719
rect 331 2715 335 2719
rect 343 2715 347 2719
rect 651 2715 655 2719
rect 1055 2715 1059 2719
rect 1163 2715 1167 2719
rect 1339 2715 1343 2719
rect 111 2707 115 2711
rect 135 2704 139 2708
rect 255 2704 259 2708
rect 407 2704 411 2708
rect 575 2704 579 2708
rect 743 2704 747 2708
rect 919 2704 923 2708
rect 1087 2704 1091 2708
rect 1255 2704 1259 2708
rect 1343 2707 1347 2711
rect 1423 2704 1427 2708
rect 1599 2704 1603 2708
rect 2007 2707 2011 2711
rect 2047 2661 2051 2665
rect 2095 2664 2099 2668
rect 2263 2664 2267 2668
rect 2439 2664 2443 2668
rect 2615 2664 2619 2668
rect 2783 2664 2787 2668
rect 2943 2664 2947 2668
rect 3095 2664 3099 2668
rect 3239 2664 3243 2668
rect 3383 2664 3387 2668
rect 3535 2664 3539 2668
rect 3943 2661 3947 2665
rect 2171 2655 2175 2659
rect 2331 2655 2335 2659
rect 2411 2655 2415 2659
rect 2523 2655 2527 2659
rect 3019 2655 3023 2659
rect 3171 2655 3175 2659
rect 3315 2655 3319 2659
rect 3459 2655 3463 2659
rect 3467 2655 3471 2659
rect 111 2641 115 2645
rect 167 2644 171 2648
rect 359 2644 363 2648
rect 559 2644 563 2648
rect 759 2644 763 2648
rect 951 2644 955 2648
rect 1143 2644 1147 2648
rect 1327 2644 1331 2648
rect 1511 2644 1515 2648
rect 1703 2644 1707 2648
rect 2007 2641 2011 2645
rect 2047 2644 2051 2648
rect 2095 2645 2099 2649
rect 2263 2645 2267 2649
rect 2439 2645 2443 2649
rect 2615 2645 2619 2649
rect 2783 2645 2787 2649
rect 2943 2645 2947 2649
rect 3095 2645 3099 2649
rect 3239 2645 3243 2649
rect 3383 2645 3387 2649
rect 3535 2645 3539 2649
rect 3943 2644 3947 2648
rect 283 2635 287 2639
rect 435 2635 439 2639
rect 635 2635 639 2639
rect 827 2635 831 2639
rect 1019 2635 1023 2639
rect 1035 2635 1039 2639
rect 1403 2635 1407 2639
rect 1587 2635 1591 2639
rect 1779 2635 1783 2639
rect 111 2624 115 2628
rect 167 2625 171 2629
rect 359 2625 363 2629
rect 559 2625 563 2629
rect 759 2625 763 2629
rect 951 2625 955 2629
rect 1143 2625 1147 2629
rect 1327 2625 1331 2629
rect 1511 2625 1515 2629
rect 1703 2625 1707 2629
rect 2007 2624 2011 2628
rect 2163 2623 2164 2627
rect 2164 2623 2167 2627
rect 2171 2623 2175 2627
rect 2523 2623 2527 2627
rect 2747 2623 2751 2627
rect 2915 2623 2919 2627
rect 3019 2623 3023 2627
rect 3171 2623 3175 2627
rect 3315 2623 3319 2627
rect 3459 2623 3463 2627
rect 343 2611 347 2615
rect 283 2599 287 2603
rect 435 2603 439 2607
rect 635 2603 639 2607
rect 1035 2603 1039 2607
rect 1199 2603 1203 2607
rect 1343 2603 1347 2607
rect 1403 2603 1407 2607
rect 1587 2603 1591 2607
rect 2331 2603 2335 2607
rect 2419 2603 2423 2607
rect 2495 2603 2499 2607
rect 2595 2603 2599 2607
rect 3035 2603 3039 2607
rect 3171 2603 3175 2607
rect 3307 2603 3311 2607
rect 3467 2603 3471 2607
rect 2047 2584 2051 2588
rect 2215 2583 2219 2587
rect 2367 2583 2371 2587
rect 2519 2583 2523 2587
rect 2671 2583 2675 2587
rect 2815 2583 2819 2587
rect 2951 2583 2955 2587
rect 3087 2583 3091 2587
rect 3223 2583 3227 2587
rect 3367 2583 3371 2587
rect 3943 2584 3947 2588
rect 651 2575 655 2579
rect 783 2575 787 2579
rect 883 2575 887 2579
rect 1011 2575 1015 2579
rect 1359 2575 1363 2579
rect 1579 2575 1583 2579
rect 1731 2575 1735 2579
rect 1779 2575 1783 2579
rect 703 2567 707 2571
rect 2047 2567 2051 2571
rect 2359 2571 2363 2575
rect 2495 2575 2499 2579
rect 2595 2575 2599 2579
rect 2747 2575 2751 2579
rect 2787 2575 2791 2579
rect 3035 2575 3039 2579
rect 3171 2575 3175 2579
rect 3307 2575 3311 2579
rect 2215 2564 2219 2568
rect 2367 2564 2371 2568
rect 2519 2564 2523 2568
rect 2671 2564 2675 2568
rect 2815 2564 2819 2568
rect 2951 2564 2955 2568
rect 3087 2564 3091 2568
rect 3223 2564 3227 2568
rect 3367 2564 3371 2568
rect 3943 2567 3947 2571
rect 111 2556 115 2560
rect 575 2555 579 2559
rect 687 2555 691 2559
rect 807 2555 811 2559
rect 935 2555 939 2559
rect 1071 2555 1075 2559
rect 1207 2555 1211 2559
rect 1351 2555 1355 2559
rect 1495 2555 1499 2559
rect 1647 2555 1651 2559
rect 1799 2555 1803 2559
rect 2007 2556 2011 2560
rect 651 2547 655 2551
rect 783 2547 787 2551
rect 883 2547 887 2551
rect 1011 2547 1015 2551
rect 111 2539 115 2543
rect 1147 2543 1151 2547
rect 1199 2547 1203 2551
rect 1571 2543 1575 2547
rect 1579 2547 1583 2551
rect 1731 2547 1735 2551
rect 575 2536 579 2540
rect 687 2536 691 2540
rect 807 2536 811 2540
rect 935 2536 939 2540
rect 1071 2536 1075 2540
rect 1207 2536 1211 2540
rect 1351 2536 1355 2540
rect 1495 2536 1499 2540
rect 1647 2536 1651 2540
rect 1799 2536 1803 2540
rect 2007 2539 2011 2543
rect 2047 2497 2051 2501
rect 2095 2500 2099 2504
rect 2215 2500 2219 2504
rect 2343 2500 2347 2504
rect 2471 2500 2475 2504
rect 2599 2500 2603 2504
rect 2719 2500 2723 2504
rect 2839 2500 2843 2504
rect 2967 2500 2971 2504
rect 3095 2500 3099 2504
rect 3223 2500 3227 2504
rect 3943 2497 3947 2501
rect 2171 2491 2175 2495
rect 2291 2491 2295 2495
rect 2419 2491 2423 2495
rect 2547 2491 2551 2495
rect 2667 2491 2671 2495
rect 2795 2491 2799 2495
rect 2915 2491 2919 2495
rect 3043 2491 3047 2495
rect 3171 2491 3175 2495
rect 3215 2491 3219 2495
rect 2047 2480 2051 2484
rect 2095 2481 2099 2485
rect 2215 2481 2219 2485
rect 2343 2481 2347 2485
rect 2471 2481 2475 2485
rect 2599 2481 2603 2485
rect 2719 2481 2723 2485
rect 2839 2481 2843 2485
rect 2967 2481 2971 2485
rect 3095 2481 3099 2485
rect 3223 2481 3227 2485
rect 3943 2480 3947 2484
rect 111 2469 115 2473
rect 503 2472 507 2476
rect 607 2472 611 2476
rect 719 2472 723 2476
rect 847 2472 851 2476
rect 983 2472 987 2476
rect 1127 2472 1131 2476
rect 1279 2472 1283 2476
rect 1431 2472 1435 2476
rect 1583 2472 1587 2476
rect 1743 2472 1747 2476
rect 1903 2472 1907 2476
rect 2007 2469 2011 2473
rect 2359 2471 2363 2475
rect 579 2463 583 2467
rect 683 2463 687 2467
rect 703 2463 707 2467
rect 923 2463 927 2467
rect 931 2463 935 2467
rect 1067 2463 1071 2467
rect 1355 2463 1359 2467
rect 1363 2463 1367 2467
rect 1659 2463 1663 2467
rect 1819 2463 1823 2467
rect 1971 2463 1975 2467
rect 2147 2459 2151 2463
rect 2171 2459 2175 2463
rect 2291 2459 2295 2463
rect 2547 2459 2551 2463
rect 2787 2459 2788 2463
rect 2788 2459 2791 2463
rect 2795 2459 2799 2463
rect 2915 2459 2919 2463
rect 3043 2459 3047 2463
rect 3171 2459 3175 2463
rect 111 2452 115 2456
rect 503 2453 507 2457
rect 607 2453 611 2457
rect 719 2453 723 2457
rect 847 2453 851 2457
rect 983 2453 987 2457
rect 1127 2453 1131 2457
rect 1279 2453 1283 2457
rect 1431 2453 1435 2457
rect 1583 2453 1587 2457
rect 1743 2453 1747 2457
rect 1903 2453 1907 2457
rect 2007 2452 2011 2456
rect 579 2439 583 2443
rect 619 2431 623 2435
rect 683 2431 687 2435
rect 931 2431 935 2435
rect 1067 2431 1071 2435
rect 1147 2431 1151 2435
rect 1363 2431 1367 2435
rect 1571 2431 1575 2435
rect 1659 2431 1663 2435
rect 1819 2431 1823 2435
rect 2243 2435 2247 2439
rect 2267 2435 2271 2439
rect 2523 2435 2527 2439
rect 2667 2435 2671 2439
rect 2763 2435 2767 2439
rect 2875 2435 2879 2439
rect 2995 2435 2999 2439
rect 3115 2435 3119 2439
rect 3215 2435 3216 2439
rect 3216 2435 3219 2439
rect 2275 2427 2279 2431
rect 2047 2416 2051 2420
rect 2071 2415 2075 2419
rect 923 2411 927 2415
rect 2191 2415 2195 2419
rect 2319 2415 2323 2419
rect 2439 2415 2443 2419
rect 2559 2415 2563 2419
rect 2679 2415 2683 2419
rect 2791 2415 2795 2419
rect 2911 2415 2915 2419
rect 3031 2415 3035 2419
rect 3151 2415 3155 2419
rect 3943 2416 3947 2420
rect 731 2403 735 2407
rect 1035 2403 1039 2407
rect 1323 2403 1327 2407
rect 1467 2403 1471 2407
rect 1731 2403 1735 2407
rect 1971 2403 1972 2407
rect 1972 2403 1975 2407
rect 2147 2407 2151 2411
rect 2267 2407 2271 2411
rect 2275 2407 2279 2411
rect 2423 2407 2427 2411
rect 2523 2407 2527 2411
rect 2643 2407 2647 2411
rect 2763 2407 2767 2411
rect 2875 2407 2879 2411
rect 2995 2407 2999 2411
rect 3115 2407 3119 2411
rect 1043 2395 1047 2399
rect 1379 2395 1383 2399
rect 1875 2395 1879 2399
rect 2047 2399 2051 2403
rect 2071 2396 2075 2400
rect 2191 2396 2195 2400
rect 2319 2396 2323 2400
rect 2439 2396 2443 2400
rect 2559 2396 2563 2400
rect 2679 2396 2683 2400
rect 2791 2396 2795 2400
rect 2911 2396 2915 2400
rect 3031 2396 3035 2400
rect 3151 2396 3155 2400
rect 3943 2399 3947 2403
rect 111 2384 115 2388
rect 535 2383 539 2387
rect 671 2383 675 2387
rect 815 2383 819 2387
rect 959 2383 963 2387
rect 1103 2383 1107 2387
rect 1247 2383 1251 2387
rect 1391 2383 1395 2387
rect 1527 2383 1531 2387
rect 1655 2383 1659 2387
rect 1791 2383 1795 2387
rect 1903 2383 1907 2387
rect 2007 2384 2011 2388
rect 619 2375 623 2379
rect 1035 2375 1039 2379
rect 1043 2375 1047 2379
rect 1323 2375 1327 2379
rect 1467 2375 1471 2379
rect 1731 2375 1735 2379
rect 111 2367 115 2371
rect 535 2364 539 2368
rect 671 2364 675 2368
rect 815 2364 819 2368
rect 883 2367 887 2371
rect 1867 2371 1871 2375
rect 1875 2375 1879 2379
rect 959 2364 963 2368
rect 1103 2364 1107 2368
rect 1247 2364 1251 2368
rect 1391 2364 1395 2368
rect 1527 2364 1531 2368
rect 1655 2364 1659 2368
rect 1791 2364 1795 2368
rect 1903 2364 1907 2368
rect 2007 2367 2011 2371
rect 2047 2329 2051 2333
rect 2167 2332 2171 2336
rect 2359 2332 2363 2336
rect 2535 2332 2539 2336
rect 2703 2332 2707 2336
rect 2871 2332 2875 2336
rect 3031 2332 3035 2336
rect 3199 2332 3203 2336
rect 3943 2329 3947 2333
rect 2243 2323 2247 2327
rect 2351 2323 2355 2327
rect 2671 2323 2675 2327
rect 2779 2323 2783 2327
rect 2947 2323 2951 2327
rect 3107 2323 3111 2327
rect 3115 2323 3119 2327
rect 2047 2312 2051 2316
rect 2167 2313 2171 2317
rect 2359 2313 2363 2317
rect 2535 2313 2539 2317
rect 2703 2313 2707 2317
rect 2871 2313 2875 2317
rect 3031 2313 3035 2317
rect 3199 2313 3203 2317
rect 3943 2312 3947 2316
rect 111 2297 115 2301
rect 535 2300 539 2304
rect 647 2300 651 2304
rect 767 2300 771 2304
rect 895 2300 899 2304
rect 1031 2300 1035 2304
rect 1167 2300 1171 2304
rect 1295 2300 1299 2304
rect 1423 2300 1427 2304
rect 1551 2300 1555 2304
rect 1671 2300 1675 2304
rect 1799 2300 1803 2304
rect 1903 2300 1907 2304
rect 2007 2297 2011 2301
rect 611 2291 615 2295
rect 731 2291 735 2295
rect 971 2291 975 2295
rect 1107 2291 1111 2295
rect 1115 2291 1119 2295
rect 1371 2291 1375 2295
rect 1379 2291 1383 2295
rect 1507 2291 1511 2295
rect 1635 2291 1639 2295
rect 1875 2291 1879 2295
rect 2235 2291 2236 2295
rect 2236 2291 2239 2295
rect 2423 2297 2427 2299
rect 2423 2295 2424 2297
rect 2424 2295 2427 2297
rect 2643 2291 2647 2295
rect 2671 2291 2675 2295
rect 2779 2291 2783 2295
rect 2947 2291 2951 2295
rect 3107 2291 3111 2295
rect 111 2280 115 2284
rect 535 2281 539 2285
rect 647 2281 651 2285
rect 767 2281 771 2285
rect 895 2281 899 2285
rect 1031 2281 1035 2285
rect 1167 2281 1171 2285
rect 1295 2281 1299 2285
rect 1423 2281 1427 2285
rect 1551 2281 1555 2285
rect 1671 2281 1675 2285
rect 1799 2281 1803 2285
rect 1903 2281 1907 2285
rect 2007 2280 2011 2284
rect 2147 2279 2151 2283
rect 2351 2279 2352 2283
rect 2352 2279 2355 2283
rect 2371 2279 2375 2283
rect 2499 2279 2503 2283
rect 2635 2279 2639 2283
rect 2915 2279 2919 2283
rect 3059 2279 3063 2283
rect 3251 2279 3255 2283
rect 1507 2267 1511 2271
rect 2235 2267 2239 2271
rect 3115 2271 3119 2275
rect 491 2259 495 2263
rect 611 2259 615 2263
rect 883 2259 887 2263
rect 971 2259 975 2263
rect 1107 2259 1111 2263
rect 1371 2259 1375 2263
rect 1635 2259 1639 2263
rect 1643 2259 1647 2263
rect 1867 2259 1868 2263
rect 1868 2259 1871 2263
rect 1875 2259 1879 2263
rect 2047 2260 2051 2264
rect 2071 2259 2075 2263
rect 2167 2259 2171 2263
rect 2287 2259 2291 2263
rect 2423 2259 2427 2263
rect 2559 2259 2563 2263
rect 499 2243 503 2247
rect 619 2243 623 2247
rect 779 2243 783 2247
rect 1115 2251 1119 2255
rect 2147 2251 2151 2255
rect 2155 2251 2159 2255
rect 1067 2243 1071 2247
rect 1251 2243 1255 2247
rect 1651 2243 1655 2247
rect 1755 2243 1759 2247
rect 2047 2243 2051 2247
rect 2363 2247 2367 2251
rect 2499 2251 2503 2255
rect 2635 2251 2639 2255
rect 2703 2259 2707 2263
rect 2839 2259 2843 2263
rect 2983 2259 2987 2263
rect 3127 2259 3131 2263
rect 3271 2259 3275 2263
rect 3943 2260 3947 2264
rect 2915 2251 2919 2255
rect 3059 2251 3063 2255
rect 3251 2251 3255 2255
rect 3259 2251 3263 2255
rect 2071 2240 2075 2244
rect 2167 2240 2171 2244
rect 2287 2240 2291 2244
rect 2423 2240 2427 2244
rect 2559 2240 2563 2244
rect 2703 2240 2707 2244
rect 2839 2240 2843 2244
rect 2983 2240 2987 2244
rect 3127 2240 3131 2244
rect 3271 2240 3275 2244
rect 3943 2243 3947 2247
rect 111 2224 115 2228
rect 415 2223 419 2227
rect 535 2223 539 2227
rect 671 2223 675 2227
rect 823 2223 827 2227
rect 991 2223 995 2227
rect 1175 2223 1179 2227
rect 1367 2223 1371 2227
rect 1567 2223 1571 2227
rect 1767 2223 1771 2227
rect 2007 2224 2011 2228
rect 491 2215 495 2219
rect 499 2215 503 2219
rect 619 2215 623 2219
rect 1067 2215 1071 2219
rect 1251 2215 1255 2219
rect 1259 2215 1263 2219
rect 1643 2215 1647 2219
rect 1651 2215 1655 2219
rect 111 2207 115 2211
rect 415 2204 419 2208
rect 535 2204 539 2208
rect 671 2204 675 2208
rect 823 2204 827 2208
rect 991 2204 995 2208
rect 1175 2204 1179 2208
rect 1367 2204 1371 2208
rect 1567 2204 1571 2208
rect 1767 2204 1771 2208
rect 2007 2207 2011 2211
rect 2047 2177 2051 2181
rect 2071 2180 2075 2184
rect 2371 2187 2375 2191
rect 2295 2180 2299 2184
rect 2503 2180 2507 2184
rect 2687 2180 2691 2184
rect 2863 2180 2867 2184
rect 3023 2180 3027 2184
rect 3175 2180 3179 2184
rect 3319 2180 3323 2184
rect 3471 2180 3475 2184
rect 3943 2177 3947 2181
rect 2371 2171 2375 2175
rect 2579 2171 2583 2175
rect 2755 2171 2759 2175
rect 2939 2171 2943 2175
rect 3099 2171 3103 2175
rect 3251 2171 3255 2175
rect 3395 2171 3399 2175
rect 3439 2171 3443 2175
rect 2047 2160 2051 2164
rect 2071 2161 2075 2165
rect 2295 2161 2299 2165
rect 2503 2161 2507 2165
rect 2687 2161 2691 2165
rect 2863 2161 2867 2165
rect 3023 2161 3027 2165
rect 3175 2161 3179 2165
rect 3319 2161 3323 2165
rect 3471 2161 3475 2165
rect 3943 2160 3947 2164
rect 3259 2147 3263 2151
rect 111 2133 115 2137
rect 135 2136 139 2140
rect 247 2136 251 2140
rect 391 2136 395 2140
rect 551 2136 555 2140
rect 711 2136 715 2140
rect 871 2136 875 2140
rect 1031 2136 1035 2140
rect 1191 2136 1195 2140
rect 1351 2136 1355 2140
rect 1511 2136 1515 2140
rect 1679 2136 1683 2140
rect 2155 2139 2159 2143
rect 2363 2139 2364 2143
rect 2364 2139 2367 2143
rect 2371 2139 2375 2143
rect 2579 2139 2583 2143
rect 2939 2139 2943 2143
rect 3099 2139 3103 2143
rect 3251 2139 3255 2143
rect 3395 2139 3399 2143
rect 2007 2133 2011 2137
rect 323 2127 327 2131
rect 467 2127 471 2131
rect 627 2127 631 2131
rect 779 2127 783 2131
rect 939 2127 943 2131
rect 955 2127 959 2131
rect 1427 2127 1431 2131
rect 1587 2127 1591 2131
rect 1755 2127 1759 2131
rect 111 2116 115 2120
rect 135 2117 139 2121
rect 247 2117 251 2121
rect 391 2117 395 2121
rect 551 2117 555 2121
rect 711 2117 715 2121
rect 871 2117 875 2121
rect 1031 2117 1035 2121
rect 1191 2117 1195 2121
rect 1351 2117 1355 2121
rect 1511 2117 1515 2121
rect 1679 2117 1683 2121
rect 2007 2116 2011 2120
rect 2475 2103 2479 2107
rect 2571 2103 2575 2107
rect 2755 2103 2756 2107
rect 2756 2103 2759 2107
rect 211 2095 215 2099
rect 323 2095 327 2099
rect 467 2095 471 2099
rect 627 2095 631 2099
rect 955 2095 959 2099
rect 1259 2095 1260 2099
rect 1260 2095 1263 2099
rect 1427 2095 1431 2099
rect 1587 2095 1591 2099
rect 2667 2095 2671 2099
rect 2947 2103 2948 2107
rect 2948 2103 2951 2107
rect 2955 2103 2959 2107
rect 3051 2103 3055 2107
rect 3147 2103 3151 2107
rect 3243 2103 3247 2107
rect 3339 2103 3343 2107
rect 3435 2103 3439 2107
rect 3531 2103 3535 2107
rect 3627 2103 3631 2107
rect 3723 2103 3727 2107
rect 3819 2103 3823 2107
rect 2047 2084 2051 2088
rect 2399 2083 2403 2087
rect 2495 2083 2499 2087
rect 2591 2083 2595 2087
rect 219 2075 223 2079
rect 379 2075 383 2079
rect 483 2075 487 2079
rect 635 2075 639 2079
rect 879 2075 883 2079
rect 939 2075 943 2079
rect 971 2075 975 2079
rect 1067 2075 1071 2079
rect 1203 2075 1207 2079
rect 1331 2075 1335 2079
rect 1459 2075 1463 2079
rect 2475 2075 2479 2079
rect 2571 2075 2575 2079
rect 2667 2075 2671 2079
rect 2687 2083 2691 2087
rect 2783 2083 2787 2087
rect 2879 2083 2883 2087
rect 2975 2083 2979 2087
rect 3071 2083 3075 2087
rect 3167 2083 3171 2087
rect 3263 2083 3267 2087
rect 3359 2083 3363 2087
rect 3455 2083 3459 2087
rect 3551 2083 3555 2087
rect 3647 2083 3651 2087
rect 3743 2083 3747 2087
rect 3839 2083 3843 2087
rect 3943 2084 3947 2088
rect 2955 2075 2959 2079
rect 3051 2075 3055 2079
rect 3147 2075 3151 2079
rect 3243 2075 3247 2079
rect 3339 2075 3343 2079
rect 3435 2075 3439 2079
rect 3531 2075 3535 2079
rect 3627 2075 3631 2079
rect 3723 2075 3727 2079
rect 3819 2075 3823 2079
rect 2047 2067 2051 2071
rect 2399 2064 2403 2068
rect 2495 2064 2499 2068
rect 2591 2064 2595 2068
rect 2687 2064 2691 2068
rect 2783 2064 2787 2068
rect 111 2056 115 2060
rect 135 2055 139 2059
rect 247 2055 251 2059
rect 399 2055 403 2059
rect 551 2055 555 2059
rect 703 2055 707 2059
rect 847 2055 851 2059
rect 991 2055 995 2059
rect 1127 2055 1131 2059
rect 1255 2055 1259 2059
rect 1383 2055 1387 2059
rect 1519 2055 1523 2059
rect 2007 2056 2011 2060
rect 3915 2071 3919 2075
rect 2879 2064 2883 2068
rect 2975 2064 2979 2068
rect 3071 2064 3075 2068
rect 3167 2064 3171 2068
rect 3263 2064 3267 2068
rect 3359 2064 3363 2068
rect 3455 2064 3459 2068
rect 3551 2064 3555 2068
rect 3647 2064 3651 2068
rect 3743 2064 3747 2068
rect 3839 2064 3843 2068
rect 3943 2067 3947 2071
rect 211 2047 215 2051
rect 219 2047 223 2051
rect 379 2047 383 2051
rect 483 2047 487 2051
rect 635 2047 639 2051
rect 971 2047 975 2051
rect 1067 2047 1071 2051
rect 1203 2047 1207 2051
rect 1331 2047 1335 2051
rect 1459 2047 1463 2051
rect 111 2039 115 2043
rect 135 2036 139 2040
rect 247 2036 251 2040
rect 399 2036 403 2040
rect 551 2036 555 2040
rect 703 2036 707 2040
rect 847 2036 851 2040
rect 991 2036 995 2040
rect 1127 2036 1131 2040
rect 1255 2036 1259 2040
rect 1383 2036 1387 2040
rect 1519 2036 1523 2040
rect 2007 2039 2011 2043
rect 2047 2001 2051 2005
rect 2191 2004 2195 2008
rect 2399 2004 2403 2008
rect 2647 2004 2651 2008
rect 2919 2004 2923 2008
rect 3215 2004 3219 2008
rect 3527 2004 3531 2008
rect 3839 2004 3843 2008
rect 3943 2001 3947 2005
rect 2315 1995 2319 1999
rect 2475 1995 2479 1999
rect 2523 1995 2527 1999
rect 2995 1995 2999 1999
rect 3003 1995 3007 1999
rect 3611 1995 3615 1999
rect 2047 1984 2051 1988
rect 2191 1985 2195 1989
rect 2399 1985 2403 1989
rect 2647 1985 2651 1989
rect 2919 1985 2923 1989
rect 3215 1985 3219 1989
rect 3527 1985 3531 1989
rect 3839 1985 3843 1989
rect 3943 1984 3947 1988
rect 111 1957 115 1961
rect 231 1960 235 1964
rect 391 1960 395 1964
rect 567 1960 571 1964
rect 751 1960 755 1964
rect 943 1960 947 1964
rect 1135 1960 1139 1964
rect 1335 1960 1339 1964
rect 1543 1960 1547 1964
rect 2523 1971 2527 1975
rect 2315 1963 2319 1967
rect 3003 1971 3007 1975
rect 2995 1963 2999 1967
rect 3611 1963 3615 1967
rect 3915 1963 3919 1967
rect 2007 1957 2011 1961
rect 315 1951 319 1955
rect 467 1951 471 1955
rect 643 1951 647 1955
rect 827 1951 831 1955
rect 879 1951 883 1955
rect 1211 1951 1215 1955
rect 1403 1951 1407 1955
rect 1459 1951 1463 1955
rect 111 1940 115 1944
rect 231 1941 235 1945
rect 391 1941 395 1945
rect 567 1941 571 1945
rect 751 1941 755 1945
rect 943 1941 947 1945
rect 1135 1941 1139 1945
rect 1335 1941 1339 1945
rect 1543 1941 1547 1945
rect 2007 1940 2011 1944
rect 2147 1939 2151 1943
rect 2475 1939 2479 1943
rect 2523 1939 2527 1943
rect 2747 1939 2751 1943
rect 3443 1939 3447 1943
rect 3655 1939 3656 1943
rect 3656 1939 3659 1943
rect 2779 1931 2783 1935
rect 307 1919 311 1923
rect 315 1919 319 1923
rect 467 1919 471 1923
rect 643 1919 647 1923
rect 827 1919 831 1923
rect 1203 1919 1204 1923
rect 1204 1919 1207 1923
rect 1211 1919 1215 1923
rect 1531 1919 1535 1923
rect 2047 1920 2051 1924
rect 2071 1919 2075 1923
rect 2239 1919 2243 1923
rect 2447 1919 2451 1923
rect 2671 1919 2675 1923
rect 2895 1919 2899 1923
rect 3127 1919 3131 1923
rect 3359 1919 3363 1923
rect 3591 1919 3595 1923
rect 3831 1919 3835 1923
rect 3943 1920 3947 1924
rect 595 1907 599 1911
rect 1111 1907 1115 1911
rect 1191 1907 1195 1911
rect 1307 1907 1311 1911
rect 1403 1907 1404 1911
rect 1404 1907 1407 1911
rect 1715 1907 1719 1911
rect 2147 1911 2151 1915
rect 2047 1903 2051 1907
rect 2315 1907 2319 1911
rect 2523 1911 2527 1915
rect 2747 1911 2751 1915
rect 2779 1911 2783 1915
rect 3443 1911 3447 1915
rect 3915 1907 3919 1911
rect 2071 1900 2075 1904
rect 2239 1900 2243 1904
rect 2447 1900 2451 1904
rect 2671 1900 2675 1904
rect 2895 1900 2899 1904
rect 3127 1900 3131 1904
rect 3359 1900 3363 1904
rect 3591 1900 3595 1904
rect 3831 1900 3835 1904
rect 3943 1903 3947 1907
rect 111 1888 115 1892
rect 511 1887 515 1891
rect 623 1887 627 1891
rect 743 1887 747 1891
rect 863 1887 867 1891
rect 983 1887 987 1891
rect 1103 1887 1107 1891
rect 1223 1887 1227 1891
rect 1335 1887 1339 1891
rect 1455 1887 1459 1891
rect 1575 1887 1579 1891
rect 1695 1887 1699 1891
rect 2007 1888 2011 1892
rect 307 1879 311 1883
rect 595 1879 599 1883
rect 111 1871 115 1875
rect 1179 1875 1183 1879
rect 1191 1879 1195 1883
rect 1307 1879 1311 1883
rect 1531 1879 1535 1883
rect 511 1868 515 1872
rect 623 1868 627 1872
rect 743 1868 747 1872
rect 863 1868 867 1872
rect 983 1868 987 1872
rect 1103 1868 1107 1872
rect 1223 1868 1227 1872
rect 1335 1868 1339 1872
rect 1455 1868 1459 1872
rect 1575 1868 1579 1872
rect 1695 1868 1699 1872
rect 2007 1871 2011 1875
rect 2047 1837 2051 1841
rect 2071 1840 2075 1844
rect 2199 1840 2203 1844
rect 2367 1840 2371 1844
rect 2543 1840 2547 1844
rect 2719 1840 2723 1844
rect 2887 1840 2891 1844
rect 3039 1840 3043 1844
rect 3183 1840 3187 1844
rect 3319 1840 3323 1844
rect 3455 1840 3459 1844
rect 3583 1840 3587 1844
rect 3711 1840 3715 1844
rect 3839 1840 3843 1844
rect 3943 1837 3947 1841
rect 2139 1831 2143 1835
rect 2155 1831 2159 1835
rect 2443 1831 2447 1835
rect 2619 1831 2623 1835
rect 2659 1831 2663 1835
rect 2963 1831 2967 1835
rect 3115 1831 3119 1835
rect 3259 1831 3263 1835
rect 3395 1831 3399 1835
rect 3523 1831 3527 1835
rect 3655 1831 3659 1835
rect 3667 1831 3671 1835
rect 3907 1831 3911 1835
rect 2047 1820 2051 1824
rect 2071 1821 2075 1825
rect 2199 1821 2203 1825
rect 2367 1821 2371 1825
rect 2543 1821 2547 1825
rect 2719 1821 2723 1825
rect 2887 1821 2891 1825
rect 3039 1821 3043 1825
rect 3183 1821 3187 1825
rect 3319 1821 3323 1825
rect 3455 1821 3459 1825
rect 3583 1821 3587 1825
rect 3711 1821 3715 1825
rect 3839 1821 3843 1825
rect 3943 1820 3947 1824
rect 111 1797 115 1801
rect 615 1800 619 1804
rect 711 1800 715 1804
rect 815 1800 819 1804
rect 927 1800 931 1804
rect 1039 1800 1043 1804
rect 1159 1800 1163 1804
rect 1279 1800 1283 1804
rect 1399 1800 1403 1804
rect 1519 1800 1523 1804
rect 2659 1807 2663 1811
rect 1639 1800 1643 1804
rect 2007 1797 2011 1801
rect 2155 1799 2159 1803
rect 2315 1799 2319 1803
rect 2443 1799 2447 1803
rect 2619 1799 2623 1803
rect 2963 1799 2967 1803
rect 3115 1799 3119 1803
rect 3259 1799 3263 1803
rect 3395 1799 3399 1803
rect 3667 1799 3671 1803
rect 3723 1799 3727 1803
rect 3915 1799 3919 1803
rect 691 1791 695 1795
rect 787 1791 791 1795
rect 891 1791 895 1795
rect 1003 1791 1007 1795
rect 1111 1791 1115 1795
rect 1235 1791 1239 1795
rect 1355 1791 1359 1795
rect 1391 1791 1395 1795
rect 1595 1791 1599 1795
rect 1715 1791 1719 1795
rect 111 1780 115 1784
rect 615 1781 619 1785
rect 711 1781 715 1785
rect 815 1781 819 1785
rect 927 1781 931 1785
rect 1039 1781 1043 1785
rect 1159 1781 1163 1785
rect 1279 1781 1283 1785
rect 1399 1781 1403 1785
rect 1519 1781 1523 1785
rect 1639 1781 1643 1785
rect 2007 1780 2011 1784
rect 2139 1783 2140 1787
rect 2140 1783 2143 1787
rect 2147 1783 2151 1787
rect 2259 1783 2263 1787
rect 2403 1783 2407 1787
rect 2563 1783 2567 1787
rect 3107 1783 3111 1787
rect 3307 1783 3311 1787
rect 3523 1783 3527 1787
rect 3739 1783 3743 1787
rect 3907 1783 3908 1787
rect 3908 1783 3911 1787
rect 2047 1764 2051 1768
rect 683 1759 684 1763
rect 684 1759 687 1763
rect 691 1759 695 1763
rect 787 1759 791 1763
rect 891 1759 895 1763
rect 1003 1759 1007 1763
rect 1179 1759 1183 1763
rect 1235 1759 1239 1763
rect 1355 1759 1359 1763
rect 1587 1759 1588 1763
rect 1588 1759 1591 1763
rect 1595 1759 1599 1763
rect 2071 1763 2075 1767
rect 2183 1763 2187 1767
rect 2327 1763 2331 1767
rect 2487 1763 2491 1767
rect 2655 1763 2659 1767
rect 2831 1763 2835 1767
rect 3023 1763 3027 1767
rect 3223 1763 3227 1767
rect 3431 1763 3435 1767
rect 3647 1763 3651 1767
rect 3839 1763 3843 1767
rect 3943 1764 3947 1768
rect 2147 1755 2151 1759
rect 2259 1755 2263 1759
rect 2403 1755 2407 1759
rect 2563 1755 2567 1759
rect 2599 1755 2603 1759
rect 435 1747 436 1751
rect 436 1747 439 1751
rect 443 1747 447 1751
rect 571 1747 575 1751
rect 771 1747 775 1751
rect 875 1747 879 1751
rect 1391 1747 1392 1751
rect 1392 1747 1395 1751
rect 1663 1747 1667 1751
rect 1759 1747 1763 1751
rect 2047 1747 2051 1751
rect 2907 1751 2911 1755
rect 3107 1755 3111 1759
rect 3307 1755 3311 1759
rect 3723 1755 3727 1759
rect 2071 1744 2075 1748
rect 2183 1744 2187 1748
rect 2327 1744 2331 1748
rect 2487 1744 2491 1748
rect 2655 1744 2659 1748
rect 2831 1744 2835 1748
rect 3023 1744 3027 1748
rect 3223 1744 3227 1748
rect 3431 1744 3435 1748
rect 3647 1744 3651 1748
rect 3839 1744 3843 1748
rect 3907 1747 3911 1751
rect 3943 1747 3947 1751
rect 111 1728 115 1732
rect 367 1727 371 1731
rect 495 1727 499 1731
rect 639 1727 643 1731
rect 799 1727 803 1731
rect 967 1727 971 1731
rect 1143 1727 1147 1731
rect 1327 1727 1331 1731
rect 1511 1727 1515 1731
rect 1703 1727 1707 1731
rect 2007 1728 2011 1732
rect 443 1719 447 1723
rect 571 1719 575 1723
rect 771 1719 775 1723
rect 875 1719 879 1723
rect 919 1719 923 1723
rect 1055 1719 1059 1723
rect 1587 1719 1591 1723
rect 1663 1719 1667 1723
rect 111 1711 115 1715
rect 367 1708 371 1712
rect 495 1708 499 1712
rect 639 1708 643 1712
rect 799 1708 803 1712
rect 967 1708 971 1712
rect 1143 1708 1147 1712
rect 1327 1708 1331 1712
rect 1511 1708 1515 1712
rect 1703 1708 1707 1712
rect 2007 1711 2011 1715
rect 2047 1673 2051 1677
rect 2223 1676 2227 1680
rect 2327 1676 2331 1680
rect 2439 1676 2443 1680
rect 2559 1676 2563 1680
rect 2687 1676 2691 1680
rect 2823 1676 2827 1680
rect 2967 1676 2971 1680
rect 3127 1676 3131 1680
rect 3303 1676 3307 1680
rect 3487 1676 3491 1680
rect 3671 1676 3675 1680
rect 3839 1676 3843 1680
rect 3943 1673 3947 1677
rect 2299 1667 2303 1671
rect 2403 1667 2407 1671
rect 2515 1667 2519 1671
rect 2635 1667 2639 1671
rect 2659 1667 2663 1671
rect 2947 1667 2951 1671
rect 3043 1667 3047 1671
rect 3203 1667 3207 1671
rect 3379 1667 3383 1671
rect 3439 1667 3443 1671
rect 3739 1667 3743 1671
rect 3915 1667 3919 1671
rect 2047 1656 2051 1660
rect 2223 1657 2227 1661
rect 2327 1657 2331 1661
rect 2439 1657 2443 1661
rect 2559 1657 2563 1661
rect 2687 1657 2691 1661
rect 2823 1657 2827 1661
rect 2967 1657 2971 1661
rect 3127 1657 3131 1661
rect 3303 1657 3307 1661
rect 3487 1657 3491 1661
rect 3671 1657 3675 1661
rect 3839 1657 3843 1661
rect 3943 1656 3947 1660
rect 435 1651 439 1655
rect 111 1641 115 1645
rect 135 1644 139 1648
rect 247 1644 251 1648
rect 399 1644 403 1648
rect 567 1644 571 1648
rect 323 1635 327 1639
rect 475 1635 479 1639
rect 643 1635 647 1639
rect 743 1644 747 1648
rect 935 1644 939 1648
rect 1135 1644 1139 1648
rect 1343 1644 1347 1648
rect 1551 1644 1555 1648
rect 1767 1644 1771 1648
rect 2007 1641 2011 1645
rect 2599 1643 2603 1647
rect 1011 1635 1015 1639
rect 1211 1635 1215 1639
rect 1411 1635 1415 1639
rect 1667 1635 1671 1639
rect 1759 1635 1763 1639
rect 2299 1635 2303 1639
rect 2403 1635 2407 1639
rect 2515 1635 2519 1639
rect 2635 1635 2639 1639
rect 2907 1635 2911 1639
rect 2947 1635 2951 1639
rect 3043 1635 3047 1639
rect 3203 1635 3207 1639
rect 3379 1635 3383 1639
rect 3795 1635 3799 1639
rect 3907 1635 3908 1639
rect 3908 1635 3911 1639
rect 111 1624 115 1628
rect 135 1625 139 1629
rect 247 1625 251 1629
rect 399 1625 403 1629
rect 567 1625 571 1629
rect 743 1625 747 1629
rect 935 1625 939 1629
rect 1135 1625 1139 1629
rect 1343 1625 1347 1629
rect 1551 1625 1555 1629
rect 1767 1625 1771 1629
rect 2007 1624 2011 1628
rect 2659 1627 2663 1631
rect 3439 1627 3443 1631
rect 2467 1619 2471 1623
rect 2579 1619 2583 1623
rect 2727 1619 2731 1623
rect 2811 1619 2815 1623
rect 3051 1619 3055 1623
rect 3171 1619 3175 1623
rect 3291 1619 3295 1623
rect 3411 1619 3415 1623
rect 1055 1611 1059 1615
rect 211 1603 215 1607
rect 323 1603 327 1607
rect 475 1603 479 1607
rect 643 1603 647 1607
rect 1011 1603 1015 1607
rect 1211 1603 1215 1607
rect 1643 1603 1647 1607
rect 1667 1603 1671 1607
rect 2047 1600 2051 1604
rect 2391 1599 2395 1603
rect 2503 1599 2507 1603
rect 2615 1599 2619 1603
rect 2735 1599 2739 1603
rect 2855 1599 2859 1603
rect 2975 1599 2979 1603
rect 3095 1599 3099 1603
rect 3215 1599 3219 1603
rect 3335 1599 3339 1603
rect 3455 1599 3459 1603
rect 3943 1600 3947 1604
rect 219 1587 223 1591
rect 339 1587 343 1591
rect 575 1587 579 1591
rect 851 1587 855 1591
rect 1147 1587 1151 1591
rect 1411 1587 1415 1591
rect 1651 1587 1655 1591
rect 1811 1587 1815 1591
rect 2467 1591 2471 1595
rect 2579 1591 2583 1595
rect 2727 1591 2731 1595
rect 2811 1591 2815 1595
rect 2819 1591 2823 1595
rect 3051 1591 3055 1595
rect 3171 1591 3175 1595
rect 3291 1591 3295 1595
rect 3411 1591 3415 1595
rect 3419 1591 3423 1595
rect 2047 1583 2051 1587
rect 2391 1580 2395 1584
rect 2503 1580 2507 1584
rect 2615 1580 2619 1584
rect 2735 1580 2739 1584
rect 2855 1580 2859 1584
rect 2975 1580 2979 1584
rect 3095 1580 3099 1584
rect 3215 1580 3219 1584
rect 3335 1580 3339 1584
rect 3455 1580 3459 1584
rect 3943 1583 3947 1587
rect 111 1568 115 1572
rect 135 1567 139 1571
rect 255 1567 259 1571
rect 423 1567 427 1571
rect 615 1567 619 1571
rect 831 1567 835 1571
rect 1063 1567 1067 1571
rect 1311 1567 1315 1571
rect 1567 1567 1571 1571
rect 1831 1567 1835 1571
rect 2007 1568 2011 1572
rect 211 1559 215 1563
rect 219 1559 223 1563
rect 339 1559 343 1563
rect 575 1559 579 1563
rect 1035 1559 1039 1563
rect 1147 1559 1151 1563
rect 1643 1559 1647 1563
rect 1651 1559 1655 1563
rect 111 1551 115 1555
rect 135 1548 139 1552
rect 255 1548 259 1552
rect 423 1548 427 1552
rect 615 1548 619 1552
rect 831 1548 835 1552
rect 1063 1548 1067 1552
rect 1311 1548 1315 1552
rect 1567 1548 1571 1552
rect 1831 1548 1835 1552
rect 2007 1551 2011 1555
rect 2047 1517 2051 1521
rect 2543 1520 2547 1524
rect 2671 1520 2675 1524
rect 2799 1520 2803 1524
rect 2935 1520 2939 1524
rect 3071 1520 3075 1524
rect 3207 1520 3211 1524
rect 3335 1520 3339 1524
rect 3463 1520 3467 1524
rect 3591 1520 3595 1524
rect 3727 1520 3731 1524
rect 3839 1520 3843 1524
rect 3943 1517 3947 1521
rect 2619 1511 2623 1515
rect 2747 1511 2751 1515
rect 2875 1511 2879 1515
rect 3011 1511 3015 1515
rect 3147 1511 3151 1515
rect 3283 1511 3287 1515
rect 3411 1511 3415 1515
rect 3539 1511 3543 1515
rect 3795 1511 3799 1515
rect 3907 1511 3911 1515
rect 2047 1500 2051 1504
rect 2543 1501 2547 1505
rect 2671 1501 2675 1505
rect 2799 1501 2803 1505
rect 2935 1501 2939 1505
rect 3071 1501 3075 1505
rect 3207 1501 3211 1505
rect 3335 1501 3339 1505
rect 3463 1501 3467 1505
rect 3591 1501 3595 1505
rect 3727 1501 3731 1505
rect 3839 1501 3843 1505
rect 3943 1500 3947 1504
rect 111 1481 115 1485
rect 239 1484 243 1488
rect 407 1484 411 1488
rect 583 1484 587 1488
rect 775 1484 779 1488
rect 967 1484 971 1488
rect 1159 1484 1163 1488
rect 1351 1484 1355 1488
rect 1543 1484 1547 1488
rect 1735 1484 1739 1488
rect 1903 1484 1907 1488
rect 2007 1481 2011 1485
rect 2819 1487 2823 1491
rect 3419 1487 3423 1491
rect 483 1475 487 1479
rect 659 1475 663 1479
rect 851 1475 855 1479
rect 1043 1475 1047 1479
rect 1235 1475 1239 1479
rect 1443 1475 1447 1479
rect 1619 1475 1623 1479
rect 1811 1475 1815 1479
rect 1819 1475 1823 1479
rect 2619 1479 2623 1483
rect 2747 1479 2751 1483
rect 2875 1479 2879 1483
rect 3011 1479 3015 1483
rect 3283 1479 3287 1483
rect 3411 1479 3415 1483
rect 3539 1479 3543 1483
rect 3791 1479 3792 1483
rect 3792 1479 3795 1483
rect 3915 1479 3919 1483
rect 111 1464 115 1468
rect 239 1465 243 1469
rect 407 1465 411 1469
rect 583 1465 587 1469
rect 775 1465 779 1469
rect 967 1465 971 1469
rect 1159 1465 1163 1469
rect 1351 1465 1355 1469
rect 1543 1465 1547 1469
rect 1735 1465 1739 1469
rect 1903 1465 1907 1469
rect 2007 1464 2011 1468
rect 1819 1451 1823 1455
rect 2595 1455 2599 1459
rect 2887 1455 2891 1459
rect 2979 1455 2983 1459
rect 3147 1455 3151 1459
rect 3387 1455 3391 1459
rect 3667 1455 3671 1459
rect 3907 1455 3908 1459
rect 3908 1455 3911 1459
rect 483 1443 487 1447
rect 659 1443 663 1447
rect 1035 1443 1036 1447
rect 1036 1443 1039 1447
rect 1043 1443 1047 1447
rect 1235 1443 1239 1447
rect 1619 1443 1623 1447
rect 1947 1443 1951 1447
rect 2715 1447 2719 1451
rect 3531 1447 3535 1451
rect 2047 1436 2051 1440
rect 2519 1435 2523 1439
rect 2631 1435 2635 1439
rect 2759 1435 2763 1439
rect 2895 1435 2899 1439
rect 3031 1435 3035 1439
rect 3175 1435 3179 1439
rect 3311 1435 3315 1439
rect 3447 1435 3451 1439
rect 3583 1435 3587 1439
rect 3719 1435 3723 1439
rect 3839 1435 3843 1439
rect 3943 1436 3947 1440
rect 671 1423 675 1427
rect 939 1423 943 1427
rect 1115 1423 1119 1427
rect 1251 1423 1255 1427
rect 1443 1423 1447 1427
rect 1823 1423 1827 1427
rect 1831 1423 1835 1427
rect 2595 1427 2599 1431
rect 2047 1419 2051 1423
rect 2707 1423 2711 1427
rect 2715 1427 2719 1431
rect 2887 1427 2891 1431
rect 2979 1427 2983 1431
rect 3387 1427 3391 1431
rect 3531 1427 3535 1431
rect 3667 1427 3671 1431
rect 2519 1416 2523 1420
rect 2631 1416 2635 1420
rect 2759 1416 2763 1420
rect 2895 1416 2899 1420
rect 3031 1416 3035 1420
rect 3175 1416 3179 1420
rect 3311 1416 3315 1420
rect 3447 1416 3451 1420
rect 3575 1419 3579 1423
rect 3583 1416 3587 1420
rect 3719 1416 3723 1420
rect 3839 1416 3843 1420
rect 3907 1419 3911 1423
rect 3943 1419 3947 1423
rect 111 1404 115 1408
rect 463 1403 467 1407
rect 583 1403 587 1407
rect 711 1403 715 1407
rect 855 1403 859 1407
rect 1007 1403 1011 1407
rect 1167 1403 1171 1407
rect 1335 1403 1339 1407
rect 1511 1403 1515 1407
rect 1687 1403 1691 1407
rect 1871 1403 1875 1407
rect 2007 1404 2011 1408
rect 671 1395 675 1399
rect 939 1395 943 1399
rect 111 1387 115 1391
rect 1243 1391 1247 1395
rect 1251 1395 1255 1399
rect 1831 1395 1835 1399
rect 1947 1395 1951 1399
rect 463 1384 467 1388
rect 583 1384 587 1388
rect 711 1384 715 1388
rect 855 1384 859 1388
rect 1007 1384 1011 1388
rect 1167 1384 1171 1388
rect 1335 1384 1339 1388
rect 1511 1384 1515 1388
rect 1687 1384 1691 1388
rect 1871 1384 1875 1388
rect 2007 1387 2011 1391
rect 2047 1353 2051 1357
rect 2399 1356 2403 1360
rect 2535 1356 2539 1360
rect 2679 1356 2683 1360
rect 2823 1356 2827 1360
rect 2967 1356 2971 1360
rect 3111 1356 3115 1360
rect 3255 1356 3259 1360
rect 3407 1356 3411 1360
rect 3559 1356 3563 1360
rect 3711 1356 3715 1360
rect 3839 1356 3843 1360
rect 3943 1353 3947 1357
rect 2475 1347 2479 1351
rect 2483 1347 2487 1351
rect 2755 1347 2759 1351
rect 2899 1347 2903 1351
rect 2923 1347 2927 1351
rect 3051 1347 3055 1351
rect 3195 1347 3199 1351
rect 3339 1347 3343 1351
rect 3635 1347 3639 1351
rect 3799 1347 3803 1351
rect 2047 1336 2051 1340
rect 2399 1337 2403 1341
rect 2535 1337 2539 1341
rect 2679 1337 2683 1341
rect 2823 1337 2827 1341
rect 2967 1337 2971 1341
rect 3111 1337 3115 1341
rect 3255 1337 3259 1341
rect 3407 1337 3411 1341
rect 3559 1337 3563 1341
rect 3711 1337 3715 1341
rect 3839 1337 3843 1341
rect 3943 1336 3947 1340
rect 111 1321 115 1325
rect 655 1324 659 1328
rect 767 1324 771 1328
rect 887 1324 891 1328
rect 1015 1324 1019 1328
rect 1143 1324 1147 1328
rect 1279 1324 1283 1328
rect 1415 1324 1419 1328
rect 1559 1324 1563 1328
rect 1703 1324 1707 1328
rect 1847 1324 1851 1328
rect 2007 1321 2011 1325
rect 731 1315 735 1319
rect 843 1315 847 1319
rect 963 1315 967 1319
rect 1091 1315 1095 1319
rect 1115 1315 1119 1319
rect 1355 1315 1359 1319
rect 1483 1315 1487 1319
rect 1635 1315 1639 1319
rect 1779 1315 1783 1319
rect 1823 1315 1827 1319
rect 2483 1315 2487 1319
rect 2923 1323 2927 1327
rect 2707 1315 2711 1319
rect 2755 1315 2759 1319
rect 2899 1315 2903 1319
rect 3195 1315 3199 1319
rect 3339 1315 3343 1319
rect 3583 1315 3587 1319
rect 3635 1315 3639 1319
rect 3915 1315 3919 1319
rect 111 1304 115 1308
rect 655 1305 659 1309
rect 767 1305 771 1309
rect 887 1305 891 1309
rect 1015 1305 1019 1309
rect 1143 1305 1147 1309
rect 1279 1305 1283 1309
rect 1415 1305 1419 1309
rect 1559 1305 1563 1309
rect 1703 1305 1707 1309
rect 1847 1305 1851 1309
rect 2007 1304 2011 1308
rect 2367 1299 2371 1303
rect 2475 1299 2479 1303
rect 2587 1299 2591 1303
rect 2723 1299 2727 1303
rect 3051 1299 3055 1303
rect 3079 1299 3083 1303
rect 3187 1299 3191 1303
rect 3363 1299 3367 1303
rect 3547 1299 3551 1303
rect 3907 1299 3908 1303
rect 3908 1299 3911 1303
rect 2731 1291 2735 1295
rect 731 1283 735 1287
rect 843 1283 847 1287
rect 963 1283 967 1287
rect 1091 1283 1095 1287
rect 1243 1283 1247 1287
rect 1355 1283 1359 1287
rect 1627 1283 1628 1287
rect 1628 1283 1631 1287
rect 1635 1283 1639 1287
rect 1779 1283 1783 1287
rect 2047 1280 2051 1284
rect 2247 1279 2251 1283
rect 2375 1279 2379 1283
rect 2511 1279 2515 1283
rect 2647 1279 2651 1283
rect 2791 1279 2795 1283
rect 2943 1279 2947 1283
rect 3111 1279 3115 1283
rect 3287 1279 3291 1283
rect 3471 1279 3475 1283
rect 3663 1279 3667 1283
rect 3839 1279 3843 1283
rect 3943 1280 3947 1284
rect 515 1267 519 1271
rect 627 1267 631 1271
rect 747 1267 751 1271
rect 875 1267 879 1271
rect 1215 1267 1219 1271
rect 1315 1267 1319 1271
rect 1483 1267 1487 1271
rect 1771 1267 1775 1271
rect 739 1259 743 1263
rect 2047 1263 2051 1267
rect 2323 1267 2327 1271
rect 2367 1271 2371 1275
rect 2587 1271 2591 1275
rect 2723 1271 2727 1275
rect 2731 1271 2735 1275
rect 3079 1271 3083 1275
rect 3187 1271 3191 1275
rect 3363 1271 3367 1275
rect 3547 1271 3551 1275
rect 3611 1271 3615 1275
rect 3915 1271 3919 1275
rect 2247 1260 2251 1264
rect 2375 1260 2379 1264
rect 2511 1260 2515 1264
rect 2647 1260 2651 1264
rect 2791 1260 2795 1264
rect 2943 1260 2947 1264
rect 3111 1260 3115 1264
rect 3287 1260 3291 1264
rect 3471 1260 3475 1264
rect 3663 1260 3667 1264
rect 3839 1260 3843 1264
rect 3943 1263 3947 1267
rect 111 1248 115 1252
rect 439 1247 443 1251
rect 551 1247 555 1251
rect 671 1247 675 1251
rect 799 1247 803 1251
rect 935 1247 939 1251
rect 1079 1247 1083 1251
rect 1231 1247 1235 1251
rect 1391 1247 1395 1251
rect 1551 1247 1555 1251
rect 1719 1247 1723 1251
rect 2007 1248 2011 1252
rect 515 1239 519 1243
rect 627 1239 631 1243
rect 747 1239 751 1243
rect 875 1239 879 1243
rect 1071 1239 1075 1243
rect 1215 1239 1219 1243
rect 1315 1239 1319 1243
rect 1627 1239 1631 1243
rect 111 1231 115 1235
rect 439 1228 443 1232
rect 551 1228 555 1232
rect 671 1228 675 1232
rect 799 1228 803 1232
rect 935 1228 939 1232
rect 1079 1228 1083 1232
rect 1231 1228 1235 1232
rect 1391 1228 1395 1232
rect 1551 1228 1555 1232
rect 1719 1228 1723 1232
rect 2007 1231 2011 1235
rect 2047 1193 2051 1197
rect 2071 1196 2075 1200
rect 2183 1196 2187 1200
rect 2303 1196 2307 1200
rect 2431 1196 2435 1200
rect 2559 1196 2563 1200
rect 2711 1196 2715 1200
rect 2887 1196 2891 1200
rect 3087 1196 3091 1200
rect 3311 1196 3315 1200
rect 3543 1196 3547 1200
rect 3783 1196 3787 1200
rect 3943 1193 3947 1197
rect 2147 1187 2151 1191
rect 2259 1187 2263 1191
rect 2379 1187 2383 1191
rect 2507 1187 2511 1191
rect 2515 1187 2519 1191
rect 2779 1187 2783 1191
rect 2795 1187 2799 1191
rect 2971 1187 2975 1191
rect 3171 1187 3175 1191
rect 3395 1187 3399 1191
rect 3859 1187 3863 1191
rect 2047 1176 2051 1180
rect 2071 1177 2075 1181
rect 2183 1177 2187 1181
rect 2303 1177 2307 1181
rect 2431 1177 2435 1181
rect 2559 1177 2563 1181
rect 2711 1177 2715 1181
rect 2887 1177 2891 1181
rect 3087 1177 3091 1181
rect 3311 1177 3315 1181
rect 3543 1177 3547 1181
rect 3783 1177 3787 1181
rect 3943 1176 3947 1180
rect 111 1165 115 1169
rect 167 1168 171 1172
rect 303 1168 307 1172
rect 463 1168 467 1172
rect 631 1168 635 1172
rect 807 1168 811 1172
rect 983 1168 987 1172
rect 1159 1168 1163 1172
rect 1335 1168 1339 1172
rect 1511 1168 1515 1172
rect 1695 1168 1699 1172
rect 2007 1165 2011 1169
rect 243 1159 247 1163
rect 379 1159 383 1163
rect 539 1159 543 1163
rect 707 1159 711 1163
rect 739 1159 743 1163
rect 1123 1159 1127 1163
rect 1235 1159 1239 1163
rect 1411 1159 1415 1163
rect 1587 1159 1591 1163
rect 1771 1159 1775 1163
rect 2515 1163 2519 1167
rect 2147 1155 2151 1159
rect 2323 1155 2327 1159
rect 2379 1155 2383 1159
rect 2507 1155 2511 1159
rect 2795 1155 2799 1159
rect 2971 1155 2975 1159
rect 3171 1155 3175 1159
rect 3395 1155 3399 1159
rect 3611 1155 3612 1159
rect 3612 1155 3615 1159
rect 3755 1155 3759 1159
rect 111 1148 115 1152
rect 167 1149 171 1153
rect 303 1149 307 1153
rect 463 1149 467 1153
rect 631 1149 635 1153
rect 807 1149 811 1153
rect 983 1149 987 1153
rect 1159 1149 1163 1153
rect 1335 1149 1339 1153
rect 1511 1149 1515 1153
rect 1695 1149 1699 1153
rect 2007 1148 2011 1152
rect 2259 1139 2263 1143
rect 2275 1139 2279 1143
rect 2483 1139 2487 1143
rect 2779 1139 2783 1143
rect 2787 1139 2791 1143
rect 2947 1139 2951 1143
rect 3163 1139 3167 1143
rect 3395 1139 3399 1143
rect 3859 1139 3863 1143
rect 243 1127 247 1131
rect 379 1127 383 1131
rect 539 1127 543 1131
rect 707 1127 711 1131
rect 1071 1127 1075 1131
rect 1123 1127 1127 1131
rect 1411 1127 1415 1131
rect 1587 1127 1591 1131
rect 2491 1131 2495 1135
rect 619 1119 623 1123
rect 203 1111 204 1115
rect 204 1111 207 1115
rect 211 1111 215 1115
rect 315 1111 319 1115
rect 451 1111 455 1115
rect 603 1111 607 1115
rect 947 1111 951 1115
rect 1235 1111 1239 1115
rect 1455 1111 1456 1115
rect 1456 1111 1459 1115
rect 1467 1111 1471 1115
rect 1819 1103 1823 1107
rect 2047 1120 2051 1124
rect 2071 1119 2075 1123
rect 2199 1119 2203 1123
rect 2351 1119 2355 1123
rect 2511 1119 2515 1123
rect 2679 1119 2683 1123
rect 2871 1119 2875 1123
rect 3087 1119 3091 1123
rect 3319 1119 3323 1123
rect 3559 1119 3563 1123
rect 3807 1119 3811 1123
rect 3943 1120 3947 1124
rect 2275 1111 2279 1115
rect 2483 1111 2487 1115
rect 2491 1111 2495 1115
rect 2787 1111 2791 1115
rect 2947 1111 2951 1115
rect 3163 1111 3167 1115
rect 3395 1111 3399 1115
rect 3403 1111 3407 1115
rect 2047 1103 2051 1107
rect 3883 1107 3887 1111
rect 2071 1100 2075 1104
rect 2199 1100 2203 1104
rect 2351 1100 2355 1104
rect 2511 1100 2515 1104
rect 2679 1100 2683 1104
rect 2871 1100 2875 1104
rect 3087 1100 3091 1104
rect 3319 1100 3323 1104
rect 3559 1100 3563 1104
rect 3807 1100 3811 1104
rect 3943 1103 3947 1107
rect 111 1092 115 1096
rect 135 1091 139 1095
rect 239 1091 243 1095
rect 375 1091 379 1095
rect 527 1091 531 1095
rect 695 1091 699 1095
rect 863 1091 867 1095
rect 1039 1091 1043 1095
rect 1215 1091 1219 1095
rect 1391 1091 1395 1095
rect 1567 1091 1571 1095
rect 1743 1091 1747 1095
rect 1903 1091 1907 1095
rect 2007 1092 2011 1096
rect 211 1083 215 1087
rect 315 1083 319 1087
rect 451 1083 455 1087
rect 603 1083 607 1087
rect 619 1083 623 1087
rect 111 1075 115 1079
rect 939 1079 943 1083
rect 947 1083 951 1087
rect 1467 1083 1471 1087
rect 1819 1083 1823 1087
rect 2135 1083 2139 1087
rect 135 1072 139 1076
rect 239 1072 243 1076
rect 375 1072 379 1076
rect 527 1072 531 1076
rect 695 1072 699 1076
rect 863 1072 867 1076
rect 1039 1072 1043 1076
rect 1215 1072 1219 1076
rect 1391 1072 1395 1076
rect 1567 1072 1571 1076
rect 1743 1072 1747 1076
rect 1903 1072 1907 1076
rect 2007 1075 2011 1079
rect 2047 1025 2051 1029
rect 2071 1028 2075 1032
rect 2263 1028 2267 1032
rect 2487 1028 2491 1032
rect 2703 1028 2707 1032
rect 2919 1028 2923 1032
rect 3119 1028 3123 1032
rect 3311 1028 3315 1032
rect 3495 1028 3499 1032
rect 3679 1028 3683 1032
rect 3839 1028 3843 1032
rect 3943 1025 3947 1029
rect 203 1019 207 1023
rect 111 1009 115 1013
rect 135 1012 139 1016
rect 287 1012 291 1016
rect 471 1012 475 1016
rect 223 1003 227 1007
rect 363 1003 367 1007
rect 547 1003 551 1007
rect 2147 1019 2151 1023
rect 2339 1019 2343 1023
rect 2563 1019 2567 1023
rect 2571 1019 2575 1023
rect 655 1012 659 1016
rect 839 1012 843 1016
rect 1015 1012 1019 1016
rect 1199 1012 1203 1016
rect 1383 1012 1387 1016
rect 1567 1012 1571 1016
rect 3003 1019 3007 1023
rect 3203 1019 3207 1023
rect 3571 1019 3575 1023
rect 3755 1019 3759 1023
rect 3907 1019 3911 1023
rect 2007 1009 2011 1013
rect 2047 1008 2051 1012
rect 2071 1009 2075 1013
rect 2263 1009 2267 1013
rect 2487 1009 2491 1013
rect 2703 1009 2707 1013
rect 2919 1009 2923 1013
rect 3039 1011 3043 1015
rect 3119 1009 3123 1013
rect 3311 1009 3315 1013
rect 3495 1009 3499 1013
rect 3679 1009 3683 1013
rect 3839 1009 3843 1013
rect 3943 1008 3947 1012
rect 979 1003 983 1007
rect 1007 1003 1011 1007
rect 1275 1003 1279 1007
rect 1455 1003 1459 1007
rect 1467 1003 1471 1007
rect 111 992 115 996
rect 135 993 139 997
rect 287 993 291 997
rect 471 993 475 997
rect 655 993 659 997
rect 839 993 843 997
rect 1015 993 1019 997
rect 1199 993 1203 997
rect 1383 993 1387 997
rect 1567 993 1571 997
rect 2007 992 2011 996
rect 2135 987 2136 991
rect 2136 987 2139 991
rect 2147 987 2151 991
rect 2339 987 2343 991
rect 2563 987 2567 991
rect 3003 987 3007 991
rect 3203 987 3207 991
rect 3403 987 3407 991
rect 3551 987 3555 991
rect 3571 987 3575 991
rect 3883 987 3887 991
rect 1467 979 1471 983
rect 2571 979 2575 983
rect 211 971 215 975
rect 223 971 227 975
rect 363 971 367 975
rect 547 971 551 975
rect 939 971 943 975
rect 979 971 983 975
rect 1275 971 1279 975
rect 1583 971 1587 975
rect 2379 971 2383 975
rect 2531 971 2535 975
rect 2691 971 2695 975
rect 2859 971 2863 975
rect 3039 971 3043 975
rect 3187 971 3191 975
rect 3339 971 3343 975
rect 3539 971 3543 975
rect 3795 971 3799 975
rect 3907 971 3908 975
rect 3908 971 3911 975
rect 271 955 275 959
rect 431 955 435 959
rect 883 955 887 959
rect 1007 955 1011 959
rect 1163 955 1167 959
rect 1299 955 1303 959
rect 1435 955 1439 959
rect 2047 952 2051 956
rect 2303 951 2307 955
rect 1315 947 1319 951
rect 2455 951 2459 955
rect 2615 951 2619 955
rect 2783 951 2787 955
rect 2951 951 2955 955
rect 3111 951 3115 955
rect 3263 951 3267 955
rect 3415 951 3419 955
rect 3559 951 3563 955
rect 3711 951 3715 955
rect 3839 951 3843 955
rect 3943 952 3947 956
rect 2379 943 2383 947
rect 2531 943 2535 947
rect 2691 943 2695 947
rect 2859 943 2863 947
rect 2907 943 2911 947
rect 3187 943 3191 947
rect 3339 943 3343 947
rect 3539 943 3543 947
rect 3551 943 3555 947
rect 3643 943 3647 947
rect 111 936 115 940
rect 135 935 139 939
rect 295 935 299 939
rect 471 935 475 939
rect 639 935 643 939
rect 799 935 803 939
rect 951 935 955 939
rect 1087 935 1091 939
rect 1223 935 1227 939
rect 1359 935 1363 939
rect 1495 935 1499 939
rect 2007 936 2011 940
rect 2047 935 2051 939
rect 3915 939 3919 943
rect 2303 932 2307 936
rect 211 927 215 931
rect 271 927 275 931
rect 111 919 115 923
rect 715 923 719 927
rect 883 927 887 931
rect 1163 927 1167 931
rect 1299 927 1303 931
rect 1435 927 1439 931
rect 2455 932 2459 936
rect 2615 932 2619 936
rect 2783 932 2787 936
rect 2951 932 2955 936
rect 3111 932 3115 936
rect 3263 932 3267 936
rect 3415 932 3419 936
rect 3559 932 3563 936
rect 3711 932 3715 936
rect 3839 932 3843 936
rect 3943 935 3947 939
rect 1583 927 1587 931
rect 135 916 139 920
rect 295 916 299 920
rect 471 916 475 920
rect 639 916 643 920
rect 799 916 803 920
rect 951 916 955 920
rect 1087 916 1091 920
rect 1223 916 1227 920
rect 1359 916 1363 920
rect 1495 916 1499 920
rect 2007 919 2011 923
rect 2047 865 2051 869
rect 2559 868 2563 872
rect 2679 868 2683 872
rect 2807 868 2811 872
rect 2943 868 2947 872
rect 3079 868 3083 872
rect 3207 868 3211 872
rect 3335 868 3339 872
rect 3463 868 3467 872
rect 3591 868 3595 872
rect 3727 868 3731 872
rect 3839 868 3843 872
rect 3943 865 3947 869
rect 111 853 115 857
rect 159 856 163 860
rect 319 856 323 860
rect 471 856 475 860
rect 615 856 619 860
rect 751 856 755 860
rect 879 856 883 860
rect 999 856 1003 860
rect 1111 856 1115 860
rect 1231 856 1235 860
rect 1351 856 1355 860
rect 2635 859 2639 863
rect 2755 859 2759 863
rect 2883 859 2887 863
rect 3019 859 3023 863
rect 3027 859 3031 863
rect 3163 859 3167 863
rect 3291 859 3295 863
rect 3419 859 3423 863
rect 3667 859 3671 863
rect 3795 859 3799 863
rect 3907 859 3911 863
rect 2007 853 2011 857
rect 235 847 239 851
rect 431 847 435 851
rect 547 847 551 851
rect 555 847 559 851
rect 699 847 703 851
rect 991 847 995 851
rect 1099 847 1103 851
rect 1187 847 1191 851
rect 1307 847 1311 851
rect 1315 847 1319 851
rect 2047 848 2051 852
rect 2559 849 2563 853
rect 2679 849 2683 853
rect 2807 849 2811 853
rect 2943 849 2947 853
rect 3079 849 3083 853
rect 3207 849 3211 853
rect 3335 849 3339 853
rect 3463 849 3467 853
rect 3591 849 3595 853
rect 3727 849 3731 853
rect 3839 849 3843 853
rect 3943 848 3947 852
rect 111 836 115 840
rect 159 837 163 841
rect 319 837 323 841
rect 471 837 475 841
rect 615 837 619 841
rect 751 837 755 841
rect 879 837 883 841
rect 999 837 1003 841
rect 1111 837 1115 841
rect 1231 837 1235 841
rect 1351 837 1355 841
rect 2007 836 2011 840
rect 2907 835 2911 839
rect 2635 827 2639 831
rect 2755 827 2759 831
rect 2883 827 2887 831
rect 3019 827 3023 831
rect 3291 827 3295 831
rect 3419 827 3423 831
rect 3643 835 3647 839
rect 3619 827 3623 831
rect 3667 827 3671 831
rect 3915 827 3919 831
rect 215 815 219 819
rect 235 815 239 819
rect 555 815 559 819
rect 699 815 703 819
rect 715 815 719 819
rect 943 815 944 819
rect 944 815 947 819
rect 991 815 995 819
rect 1099 815 1103 819
rect 1187 815 1191 819
rect 1307 815 1311 819
rect 2411 811 2415 815
rect 2547 811 2551 815
rect 2855 811 2859 815
rect 3027 811 3031 815
rect 3163 811 3167 815
rect 3315 811 3319 815
rect 3643 811 3647 815
rect 3771 811 3772 815
rect 3772 811 3775 815
rect 3907 811 3908 815
rect 3908 811 3911 815
rect 307 803 311 807
rect 403 803 407 807
rect 547 803 551 807
rect 635 803 639 807
rect 799 803 803 807
rect 1067 803 1071 807
rect 1179 803 1183 807
rect 1371 803 1375 807
rect 1403 803 1407 807
rect 2719 803 2723 807
rect 1411 795 1415 799
rect 2047 792 2051 796
rect 2335 791 2339 795
rect 2471 791 2475 795
rect 2615 791 2619 795
rect 2767 791 2771 795
rect 2919 791 2923 795
rect 3079 791 3083 795
rect 3239 791 3243 795
rect 3391 791 3395 795
rect 3543 791 3547 795
rect 3703 791 3707 795
rect 3839 791 3843 795
rect 3943 792 3947 796
rect 111 784 115 788
rect 223 783 227 787
rect 383 783 387 787
rect 535 783 539 787
rect 679 783 683 787
rect 815 783 819 787
rect 951 783 955 787
rect 1079 783 1083 787
rect 1199 783 1203 787
rect 1327 783 1331 787
rect 1455 783 1459 787
rect 2007 784 2011 788
rect 2411 783 2415 787
rect 2547 783 2551 787
rect 215 775 219 779
rect 307 775 311 779
rect 635 775 639 779
rect 799 775 803 779
rect 111 767 115 771
rect 891 771 895 775
rect 943 775 947 779
rect 1067 775 1071 779
rect 1179 775 1183 779
rect 1403 775 1407 779
rect 1411 775 1415 779
rect 2047 775 2051 779
rect 2691 779 2695 783
rect 2719 783 2723 787
rect 2855 783 2859 787
rect 3315 783 3319 787
rect 3467 779 3471 783
rect 3619 783 3623 787
rect 3643 783 3647 787
rect 3915 779 3919 783
rect 2335 772 2339 776
rect 2471 772 2475 776
rect 2615 772 2619 776
rect 2767 772 2771 776
rect 2919 772 2923 776
rect 3079 772 3083 776
rect 3239 772 3243 776
rect 3391 772 3395 776
rect 3543 772 3547 776
rect 3703 772 3707 776
rect 3839 772 3843 776
rect 3943 775 3947 779
rect 223 764 227 768
rect 383 764 387 768
rect 535 764 539 768
rect 679 764 683 768
rect 815 764 819 768
rect 951 764 955 768
rect 1079 764 1083 768
rect 1199 764 1203 768
rect 1327 764 1331 768
rect 1455 764 1459 768
rect 2007 767 2011 771
rect 2047 705 2051 709
rect 2071 708 2075 712
rect 2183 708 2187 712
rect 2335 708 2339 712
rect 2487 708 2491 712
rect 2639 708 2643 712
rect 2807 708 2811 712
rect 2983 708 2987 712
rect 3167 708 3171 712
rect 3367 708 3371 712
rect 3575 708 3579 712
rect 3783 708 3787 712
rect 111 697 115 701
rect 311 700 315 704
rect 471 700 475 704
rect 639 700 643 704
rect 807 700 811 704
rect 975 700 979 704
rect 1135 700 1139 704
rect 1295 700 1299 704
rect 1455 700 1459 704
rect 1607 700 1611 704
rect 1767 700 1771 704
rect 3943 705 3947 709
rect 1903 700 1907 704
rect 2007 697 2011 701
rect 2055 699 2059 703
rect 2155 699 2159 703
rect 2267 699 2271 703
rect 2419 699 2423 703
rect 2571 699 2575 703
rect 2883 699 2887 703
rect 3059 699 3063 703
rect 3243 699 3247 703
rect 3319 699 3323 703
rect 3451 699 3455 703
rect 3771 699 3775 703
rect 403 691 407 695
rect 547 691 551 695
rect 555 691 559 695
rect 943 691 947 695
rect 1043 691 1047 695
rect 1211 691 1215 695
rect 1371 691 1375 695
rect 1583 691 1587 695
rect 1683 691 1687 695
rect 1699 691 1703 695
rect 1859 691 1863 695
rect 2047 688 2051 692
rect 2071 689 2075 693
rect 2183 689 2187 693
rect 2335 689 2339 693
rect 2487 689 2491 693
rect 2639 689 2643 693
rect 2807 689 2811 693
rect 2983 689 2987 693
rect 3167 689 3171 693
rect 3367 689 3371 693
rect 3575 689 3579 693
rect 3783 689 3787 693
rect 3943 688 3947 692
rect 111 680 115 684
rect 311 681 315 685
rect 471 681 475 685
rect 639 681 643 685
rect 807 681 811 685
rect 975 681 979 685
rect 1135 681 1139 685
rect 1295 681 1299 685
rect 1455 681 1459 685
rect 1607 681 1611 685
rect 1767 681 1771 685
rect 1903 681 1907 685
rect 2007 680 2011 684
rect 3319 675 3323 679
rect 555 667 559 671
rect 2155 667 2159 671
rect 2267 667 2271 671
rect 2419 667 2423 671
rect 2571 667 2575 671
rect 2691 667 2695 671
rect 2883 667 2887 671
rect 3059 667 3063 671
rect 3451 667 3455 671
rect 3467 671 3471 675
rect 3875 667 3879 671
rect 523 659 527 663
rect 547 659 551 663
rect 891 659 895 663
rect 943 659 947 663
rect 1203 659 1204 663
rect 1204 659 1207 663
rect 1211 659 1215 663
rect 1475 659 1479 663
rect 1583 659 1587 663
rect 1683 659 1687 663
rect 2055 659 2059 663
rect 315 643 319 647
rect 371 647 375 651
rect 699 647 703 651
rect 867 647 871 651
rect 1043 647 1047 651
rect 1187 647 1191 651
rect 1339 647 1343 651
rect 1619 647 1623 651
rect 1819 647 1823 651
rect 1859 647 1860 651
rect 1860 647 1863 651
rect 1867 647 1871 651
rect 1483 639 1487 643
rect 1979 643 1983 647
rect 2147 643 2151 647
rect 2315 643 2319 647
rect 2763 643 2767 647
rect 2923 643 2927 647
rect 3243 643 3247 647
rect 3395 643 3399 647
rect 3915 643 3919 647
rect 3403 635 3407 639
rect 111 628 115 632
rect 295 627 299 631
rect 447 627 451 631
rect 615 627 619 631
rect 783 627 787 631
rect 951 627 955 631
rect 1111 627 1115 631
rect 1263 627 1267 631
rect 1399 627 1403 631
rect 1535 627 1539 631
rect 1663 627 1667 631
rect 1791 627 1795 631
rect 1903 627 1907 631
rect 2007 628 2011 632
rect 2047 624 2051 628
rect 371 619 375 623
rect 523 619 527 623
rect 111 611 115 615
rect 691 615 695 619
rect 699 619 703 623
rect 867 619 871 623
rect 1187 619 1191 623
rect 1339 619 1343 623
rect 1475 619 1479 623
rect 1483 619 1487 623
rect 1619 619 1623 623
rect 1867 619 1871 623
rect 2071 623 2075 627
rect 1979 619 1983 623
rect 2239 623 2243 627
rect 2423 623 2427 627
rect 2623 623 2627 627
rect 2839 623 2843 627
rect 3071 623 3075 627
rect 3319 623 3323 627
rect 3575 623 3579 627
rect 3839 623 3843 627
rect 3943 624 3947 628
rect 295 608 299 612
rect 447 608 451 612
rect 615 608 619 612
rect 783 608 787 612
rect 951 608 955 612
rect 1111 608 1115 612
rect 1263 608 1267 612
rect 1399 608 1403 612
rect 1535 608 1539 612
rect 1663 608 1667 612
rect 1791 608 1795 612
rect 1903 608 1907 612
rect 2007 611 2011 615
rect 2147 615 2151 619
rect 2315 615 2319 619
rect 2323 615 2327 619
rect 2047 607 2051 611
rect 2699 611 2703 615
rect 2763 615 2767 619
rect 2923 615 2927 619
rect 3395 615 3399 619
rect 3403 615 3407 619
rect 3915 611 3919 615
rect 2071 604 2075 608
rect 2239 604 2243 608
rect 2423 604 2427 608
rect 2623 604 2627 608
rect 2839 604 2843 608
rect 3071 604 3075 608
rect 3319 604 3323 608
rect 3575 604 3579 608
rect 3839 604 3843 608
rect 3943 607 3947 611
rect 111 541 115 545
rect 239 544 243 548
rect 415 544 419 548
rect 607 544 611 548
rect 799 544 803 548
rect 991 544 995 548
rect 1175 544 1179 548
rect 1351 544 1355 548
rect 1519 544 1523 548
rect 1687 544 1691 548
rect 1863 544 1867 548
rect 2007 541 2011 545
rect 2047 541 2051 545
rect 2191 544 2195 548
rect 2287 544 2291 548
rect 2383 544 2387 548
rect 2479 544 2483 548
rect 2583 544 2587 548
rect 2711 544 2715 548
rect 2871 544 2875 548
rect 3071 544 3075 548
rect 3303 544 3307 548
rect 3551 544 3555 548
rect 3807 544 3811 548
rect 3943 541 3947 545
rect 315 535 319 539
rect 371 535 375 539
rect 755 535 759 539
rect 875 535 879 539
rect 883 535 887 539
rect 1251 535 1255 539
rect 1427 535 1431 539
rect 1595 535 1599 539
rect 1763 535 1767 539
rect 1819 535 1823 539
rect 2267 535 2271 539
rect 2363 535 2367 539
rect 2459 535 2463 539
rect 2555 535 2559 539
rect 2563 535 2567 539
rect 2787 535 2791 539
rect 2947 535 2951 539
rect 3147 535 3151 539
rect 3479 535 3483 539
rect 3627 535 3631 539
rect 3875 535 3879 539
rect 111 524 115 528
rect 239 525 243 529
rect 415 525 419 529
rect 607 525 611 529
rect 799 525 803 529
rect 991 525 995 529
rect 1175 525 1179 529
rect 1351 525 1355 529
rect 1519 525 1523 529
rect 1687 525 1691 529
rect 1863 525 1867 529
rect 2007 524 2011 528
rect 2047 524 2051 528
rect 2191 525 2195 529
rect 2287 525 2291 529
rect 2383 525 2387 529
rect 2479 525 2483 529
rect 2583 525 2587 529
rect 2711 525 2715 529
rect 2871 525 2875 529
rect 3071 525 3075 529
rect 3303 525 3307 529
rect 3551 525 3555 529
rect 3807 525 3811 529
rect 3943 524 3947 528
rect 2323 511 2327 515
rect 371 503 375 507
rect 539 503 543 507
rect 691 503 695 507
rect 755 503 759 507
rect 875 503 879 507
rect 1251 503 1255 507
rect 1427 503 1431 507
rect 1595 503 1599 507
rect 1763 503 1767 507
rect 2267 503 2271 507
rect 2363 503 2367 507
rect 2459 503 2463 507
rect 2555 503 2559 507
rect 2699 503 2703 507
rect 2787 503 2791 507
rect 2947 503 2951 507
rect 3147 503 3151 507
rect 3479 503 3483 507
rect 3915 503 3919 507
rect 203 491 204 495
rect 204 491 207 495
rect 211 491 215 495
rect 363 491 367 495
rect 883 491 887 495
rect 1103 491 1107 495
rect 1195 491 1199 495
rect 1395 491 1399 495
rect 1491 491 1495 495
rect 2507 491 2511 495
rect 2603 491 2607 495
rect 2699 491 2703 495
rect 2803 491 2807 495
rect 2923 491 2927 495
rect 3259 491 3263 495
rect 3459 491 3463 495
rect 3627 491 3631 495
rect 3859 491 3863 495
rect 1291 483 1295 487
rect 2563 483 2567 487
rect 111 472 115 476
rect 135 471 139 475
rect 287 471 291 475
rect 463 471 467 475
rect 639 471 643 475
rect 807 471 811 475
rect 967 471 971 475
rect 1119 471 1123 475
rect 1271 471 1275 475
rect 1415 471 1419 475
rect 1567 471 1571 475
rect 2007 472 2011 476
rect 2047 472 2051 476
rect 2431 471 2435 475
rect 2527 471 2531 475
rect 2623 471 2627 475
rect 2727 471 2731 475
rect 2847 471 2851 475
rect 2999 471 3003 475
rect 3175 471 3179 475
rect 3375 471 3379 475
rect 3591 471 3595 475
rect 3807 471 3811 475
rect 3943 472 3947 476
rect 211 463 215 467
rect 363 463 367 467
rect 539 463 543 467
rect 547 463 551 467
rect 1103 463 1107 467
rect 1195 463 1199 467
rect 1395 463 1399 467
rect 1491 463 1495 467
rect 2507 463 2511 467
rect 2603 463 2607 467
rect 2699 463 2703 467
rect 2803 463 2807 467
rect 2923 463 2927 467
rect 2935 463 2939 467
rect 3083 463 3087 467
rect 3259 463 3263 467
rect 3459 463 3463 467
rect 111 455 115 459
rect 135 452 139 456
rect 287 452 291 456
rect 463 452 467 456
rect 639 452 643 456
rect 807 452 811 456
rect 967 452 971 456
rect 1119 452 1123 456
rect 1271 452 1275 456
rect 1415 452 1419 456
rect 1567 452 1571 456
rect 2007 455 2011 459
rect 2047 455 2051 459
rect 3883 459 3887 463
rect 2431 452 2435 456
rect 2527 452 2531 456
rect 2623 452 2627 456
rect 2727 452 2731 456
rect 2847 452 2851 456
rect 2999 452 3003 456
rect 3175 452 3179 456
rect 3375 452 3379 456
rect 3591 452 3595 456
rect 3807 452 3811 456
rect 3943 455 3947 459
rect 111 385 115 389
rect 135 388 139 392
rect 279 388 283 392
rect 439 388 443 392
rect 583 388 587 392
rect 719 388 723 392
rect 847 388 851 392
rect 967 388 971 392
rect 1087 388 1091 392
rect 1207 388 1211 392
rect 1327 388 1331 392
rect 2007 385 2011 389
rect 2047 389 2051 393
rect 2431 392 2435 396
rect 2527 392 2531 396
rect 2623 392 2627 396
rect 2719 392 2723 396
rect 2815 392 2819 396
rect 2927 392 2931 396
rect 3063 392 3067 396
rect 3223 392 3227 396
rect 3399 392 3403 396
rect 3591 392 3595 396
rect 3783 392 3787 396
rect 3943 389 3947 393
rect 203 379 207 383
rect 111 368 115 372
rect 135 369 139 373
rect 203 371 207 375
rect 515 379 519 383
rect 659 379 663 383
rect 795 379 799 383
rect 923 379 927 383
rect 1043 379 1047 383
rect 1163 379 1167 383
rect 1283 379 1287 383
rect 1291 379 1295 383
rect 2507 383 2511 387
rect 2603 383 2607 387
rect 2611 383 2615 387
rect 2707 383 2711 387
rect 2803 383 2807 387
rect 3003 383 3007 387
rect 3139 383 3143 387
rect 3299 383 3303 387
rect 3475 383 3479 387
rect 3499 383 3503 387
rect 3859 383 3863 387
rect 279 369 283 373
rect 439 369 443 373
rect 583 369 587 373
rect 719 369 723 373
rect 847 369 851 373
rect 967 369 971 373
rect 1087 369 1091 373
rect 1207 369 1211 373
rect 1327 369 1331 373
rect 2007 368 2011 372
rect 2047 372 2051 376
rect 2431 373 2435 377
rect 2527 373 2531 377
rect 2623 373 2627 377
rect 2719 373 2723 377
rect 2815 373 2819 377
rect 2927 373 2931 377
rect 3063 373 3067 377
rect 3223 373 3227 377
rect 3399 373 3403 377
rect 3591 373 3595 377
rect 3783 373 3787 377
rect 3943 372 3947 376
rect 547 355 551 359
rect 2611 359 2615 363
rect 3083 359 3087 363
rect 203 347 204 351
rect 204 347 207 351
rect 219 347 223 351
rect 515 347 519 351
rect 659 347 663 351
rect 895 347 899 351
rect 923 347 927 351
rect 1043 347 1047 351
rect 1163 347 1167 351
rect 1283 347 1287 351
rect 2507 351 2511 355
rect 2707 351 2711 355
rect 2803 351 2807 355
rect 2935 351 2939 355
rect 3003 351 3007 355
rect 3139 351 3143 355
rect 3299 351 3303 355
rect 3475 351 3479 355
rect 3731 351 3735 355
rect 2603 343 2607 347
rect 3499 343 3503 347
rect 499 335 503 339
rect 619 335 623 339
rect 795 335 799 339
rect 987 335 991 339
rect 1115 335 1119 339
rect 1235 335 1239 339
rect 1355 335 1359 339
rect 1603 335 1607 339
rect 747 327 751 331
rect 2315 335 2319 339
rect 2435 327 2439 331
rect 2699 335 2703 339
rect 3027 335 3031 339
rect 3195 335 3199 339
rect 3371 335 3375 339
rect 3755 335 3759 339
rect 3883 335 3887 339
rect 2707 327 2711 331
rect 111 316 115 320
rect 143 315 147 319
rect 219 315 223 319
rect 319 315 323 319
rect 479 315 483 319
rect 631 315 635 319
rect 775 315 779 319
rect 903 315 907 319
rect 1031 315 1035 319
rect 1151 315 1155 319
rect 1271 315 1275 319
rect 1391 315 1395 319
rect 2007 316 2011 320
rect 2047 316 2051 320
rect 2191 315 2195 319
rect 2327 315 2331 319
rect 2471 315 2475 319
rect 2623 315 2627 319
rect 2783 315 2787 319
rect 2951 315 2955 319
rect 3119 315 3123 319
rect 3295 315 3299 319
rect 3471 315 3475 319
rect 3655 315 3659 319
rect 3839 315 3843 319
rect 3943 316 3947 320
rect 619 307 623 311
rect 111 299 115 303
rect 707 303 711 307
rect 747 307 751 311
rect 895 307 899 311
rect 987 307 991 311
rect 1115 307 1119 311
rect 1235 307 1239 311
rect 1355 307 1359 311
rect 2315 307 2319 311
rect 143 296 147 300
rect 319 296 323 300
rect 479 296 483 300
rect 631 296 635 300
rect 775 296 779 300
rect 903 296 907 300
rect 1031 296 1035 300
rect 1151 296 1155 300
rect 1271 296 1275 300
rect 1391 296 1395 300
rect 2007 299 2011 303
rect 2047 299 2051 303
rect 2415 303 2419 307
rect 2435 307 2439 311
rect 2699 307 2703 311
rect 2707 307 2711 311
rect 3027 307 3031 311
rect 3195 307 3199 311
rect 3371 307 3375 311
rect 3411 307 3415 311
rect 3731 307 3735 311
rect 3915 303 3919 307
rect 2191 296 2195 300
rect 2327 296 2331 300
rect 2471 296 2475 300
rect 2623 296 2627 300
rect 2783 296 2787 300
rect 2951 296 2955 300
rect 3119 296 3123 300
rect 3295 296 3299 300
rect 3471 296 3475 300
rect 3655 296 3659 300
rect 3839 296 3843 300
rect 3943 299 3947 303
rect 111 229 115 233
rect 223 232 227 236
rect 391 232 395 236
rect 559 232 563 236
rect 735 232 739 236
rect 903 232 907 236
rect 1063 232 1067 236
rect 1215 232 1219 236
rect 1359 232 1363 236
rect 1511 232 1515 236
rect 1663 232 1667 236
rect 2007 229 2011 233
rect 2047 233 2051 237
rect 2071 236 2075 240
rect 2215 236 2219 240
rect 2399 236 2403 240
rect 2591 236 2595 240
rect 2791 236 2795 240
rect 2983 236 2987 240
rect 3167 236 3171 240
rect 3343 236 3347 240
rect 3511 236 3515 240
rect 3687 236 3691 240
rect 3839 236 3843 240
rect 3943 233 3947 237
rect 299 223 303 227
rect 467 223 471 227
rect 499 223 503 227
rect 811 223 815 227
rect 1139 223 1143 227
rect 1291 223 1295 227
rect 1435 223 1439 227
rect 1587 223 1591 227
rect 1603 223 1607 227
rect 2147 227 2151 231
rect 2291 227 2295 231
rect 2475 227 2479 231
rect 2667 227 2671 231
rect 2675 227 2679 231
rect 2875 227 2879 231
rect 3067 227 3071 231
rect 3251 227 3255 231
rect 3587 227 3591 231
rect 3755 227 3759 231
rect 3907 227 3911 231
rect 111 212 115 216
rect 223 213 227 217
rect 391 213 395 217
rect 559 213 563 217
rect 735 213 739 217
rect 903 213 907 217
rect 1063 213 1067 217
rect 1215 213 1219 217
rect 1359 213 1363 217
rect 1511 213 1515 217
rect 1663 213 1667 217
rect 2007 212 2011 216
rect 2047 216 2051 220
rect 2071 217 2075 221
rect 2215 217 2219 221
rect 2399 217 2403 221
rect 2591 217 2595 221
rect 2791 217 2795 221
rect 2983 217 2987 221
rect 3167 217 3171 221
rect 3343 217 3347 221
rect 3511 217 3515 221
rect 3687 217 3691 221
rect 3839 217 3843 221
rect 3943 216 3947 220
rect 2675 203 2679 207
rect 231 191 235 195
rect 299 191 303 195
rect 467 191 471 195
rect 707 191 711 195
rect 811 191 815 195
rect 1091 191 1095 195
rect 1139 191 1143 195
rect 1291 191 1295 195
rect 1435 191 1439 195
rect 1587 191 1591 195
rect 2147 195 2151 199
rect 2415 195 2419 199
rect 2475 195 2479 199
rect 2667 195 2671 199
rect 3067 195 3071 199
rect 3251 195 3255 199
rect 3411 195 3412 199
rect 3412 195 3415 199
rect 3587 195 3591 199
rect 3915 195 3919 199
rect 3631 187 3635 191
rect 2291 159 2295 163
rect 2419 159 2423 163
rect 2571 159 2575 163
rect 2875 159 2879 163
rect 2919 159 2923 163
rect 3019 159 3023 163
rect 3147 159 3151 163
rect 3267 159 3271 163
rect 3387 159 3391 163
rect 3499 159 3503 163
rect 3603 159 3607 163
rect 3827 159 3831 163
rect 3907 159 3908 163
rect 3908 159 3911 163
rect 427 147 431 151
rect 523 147 527 151
rect 619 147 623 151
rect 715 147 719 151
rect 811 147 815 151
rect 995 147 999 151
rect 1195 147 1199 151
rect 1291 147 1295 151
rect 1699 147 1703 151
rect 1795 147 1799 151
rect 1891 147 1895 151
rect 2579 151 2583 155
rect 1099 139 1103 143
rect 2047 140 2051 144
rect 2071 139 2075 143
rect 2191 139 2195 143
rect 2343 139 2347 143
rect 2495 139 2499 143
rect 2647 139 2651 143
rect 2799 139 2803 143
rect 2943 139 2947 143
rect 3071 139 3075 143
rect 3191 139 3195 143
rect 3311 139 3315 143
rect 3423 139 3427 143
rect 3527 139 3531 143
rect 3639 139 3643 143
rect 3743 139 3747 143
rect 3839 139 3843 143
rect 3943 140 3947 144
rect 111 128 115 132
rect 151 127 155 131
rect 247 127 251 131
rect 343 127 347 131
rect 439 127 443 131
rect 535 127 539 131
rect 631 127 635 131
rect 727 127 731 131
rect 823 127 827 131
rect 919 127 923 131
rect 1015 127 1019 131
rect 1111 127 1115 131
rect 1207 127 1211 131
rect 1303 127 1307 131
rect 1407 127 1411 131
rect 1511 127 1515 131
rect 1615 127 1619 131
rect 1711 127 1715 131
rect 1807 127 1811 131
rect 1903 127 1907 131
rect 2007 128 2011 132
rect 2419 131 2423 135
rect 2571 131 2575 135
rect 2579 131 2583 135
rect 2919 131 2923 135
rect 3019 131 3023 135
rect 3147 131 3151 135
rect 3267 131 3271 135
rect 3387 131 3391 135
rect 3499 131 3503 135
rect 3603 131 3607 135
rect 3631 131 3635 135
rect 3827 131 3831 135
rect 227 119 231 123
rect 427 119 431 123
rect 523 119 527 123
rect 619 119 623 123
rect 715 119 719 123
rect 811 119 815 123
rect 995 119 999 123
rect 1091 119 1095 123
rect 1099 119 1103 123
rect 1195 119 1199 123
rect 1291 119 1295 123
rect 1699 119 1703 123
rect 1795 119 1799 123
rect 1891 119 1895 123
rect 2047 123 2051 127
rect 2071 120 2075 124
rect 2191 120 2195 124
rect 2343 120 2347 124
rect 2495 120 2499 124
rect 2647 120 2651 124
rect 2799 120 2803 124
rect 2943 120 2947 124
rect 3071 120 3075 124
rect 3191 120 3195 124
rect 3311 120 3315 124
rect 3423 120 3427 124
rect 3527 120 3531 124
rect 3639 120 3643 124
rect 3743 120 3747 124
rect 3839 120 3843 124
rect 3943 123 3947 127
rect 111 111 115 115
rect 151 108 155 112
rect 247 108 251 112
rect 343 108 347 112
rect 439 108 443 112
rect 535 108 539 112
rect 631 108 635 112
rect 727 108 731 112
rect 823 108 827 112
rect 919 108 923 112
rect 1015 108 1019 112
rect 1111 108 1115 112
rect 1207 108 1211 112
rect 1303 108 1307 112
rect 1407 108 1411 112
rect 1511 108 1515 112
rect 1615 108 1619 112
rect 1711 108 1715 112
rect 1807 108 1811 112
rect 1903 108 1907 112
rect 2007 111 2011 115
<< m3 >>
rect 2047 4022 2051 4023
rect 2047 4017 2051 4018
rect 2071 4022 2075 4023
rect 2071 4017 2075 4018
rect 2327 4022 2331 4023
rect 2327 4017 2331 4018
rect 2591 4022 2595 4023
rect 2591 4017 2595 4018
rect 2839 4022 2843 4023
rect 2839 4017 2843 4018
rect 3087 4022 3091 4023
rect 3087 4017 3091 4018
rect 3343 4022 3347 4023
rect 3343 4017 3347 4018
rect 3943 4022 3947 4023
rect 3943 4017 3947 4018
rect 111 4002 115 4003
rect 111 3997 115 3998
rect 311 4002 315 4003
rect 311 3997 315 3998
rect 511 4002 515 4003
rect 511 3997 515 3998
rect 703 4002 707 4003
rect 703 3997 707 3998
rect 887 4002 891 4003
rect 887 3997 891 3998
rect 1063 4002 1067 4003
rect 1063 3997 1067 3998
rect 1231 4002 1235 4003
rect 1231 3997 1235 3998
rect 1383 4002 1387 4003
rect 1383 3997 1387 3998
rect 1519 4002 1523 4003
rect 1519 3997 1523 3998
rect 1655 4002 1659 4003
rect 1655 3997 1659 3998
rect 1791 4002 1795 4003
rect 1791 3997 1795 3998
rect 1903 4002 1907 4003
rect 1903 3997 1907 3998
rect 2007 4002 2011 4003
rect 2007 3997 2011 3998
rect 112 3970 114 3997
rect 312 3973 314 3997
rect 512 3973 514 3997
rect 704 3973 706 3997
rect 888 3973 890 3997
rect 1064 3973 1066 3997
rect 1232 3973 1234 3997
rect 1384 3973 1386 3997
rect 1520 3973 1522 3997
rect 1656 3973 1658 3997
rect 1792 3973 1794 3997
rect 1904 3973 1906 3997
rect 310 3972 316 3973
rect 110 3969 116 3970
rect 110 3965 111 3969
rect 115 3965 116 3969
rect 310 3968 311 3972
rect 315 3968 316 3972
rect 310 3967 316 3968
rect 510 3972 516 3973
rect 510 3968 511 3972
rect 515 3968 516 3972
rect 510 3967 516 3968
rect 702 3972 708 3973
rect 702 3968 703 3972
rect 707 3968 708 3972
rect 702 3967 708 3968
rect 886 3972 892 3973
rect 886 3968 887 3972
rect 891 3968 892 3972
rect 886 3967 892 3968
rect 1062 3972 1068 3973
rect 1062 3968 1063 3972
rect 1067 3968 1068 3972
rect 1062 3967 1068 3968
rect 1230 3972 1236 3973
rect 1230 3968 1231 3972
rect 1235 3968 1236 3972
rect 1230 3967 1236 3968
rect 1382 3972 1388 3973
rect 1382 3968 1383 3972
rect 1387 3968 1388 3972
rect 1382 3967 1388 3968
rect 1518 3972 1524 3973
rect 1518 3968 1519 3972
rect 1523 3968 1524 3972
rect 1518 3967 1524 3968
rect 1654 3972 1660 3973
rect 1654 3968 1655 3972
rect 1659 3968 1660 3972
rect 1654 3967 1660 3968
rect 1790 3972 1796 3973
rect 1790 3968 1791 3972
rect 1795 3968 1796 3972
rect 1790 3967 1796 3968
rect 1902 3972 1908 3973
rect 1902 3968 1903 3972
rect 1907 3968 1908 3972
rect 2008 3970 2010 3997
rect 2048 3990 2050 4017
rect 2072 3993 2074 4017
rect 2328 3993 2330 4017
rect 2592 3993 2594 4017
rect 2840 3993 2842 4017
rect 3088 3993 3090 4017
rect 3344 3993 3346 4017
rect 2070 3992 2076 3993
rect 2046 3989 2052 3990
rect 2046 3985 2047 3989
rect 2051 3985 2052 3989
rect 2070 3988 2071 3992
rect 2075 3988 2076 3992
rect 2070 3987 2076 3988
rect 2326 3992 2332 3993
rect 2326 3988 2327 3992
rect 2331 3988 2332 3992
rect 2326 3987 2332 3988
rect 2590 3992 2596 3993
rect 2590 3988 2591 3992
rect 2595 3988 2596 3992
rect 2590 3987 2596 3988
rect 2838 3992 2844 3993
rect 2838 3988 2839 3992
rect 2843 3988 2844 3992
rect 2838 3987 2844 3988
rect 3086 3992 3092 3993
rect 3086 3988 3087 3992
rect 3091 3988 3092 3992
rect 3086 3987 3092 3988
rect 3342 3992 3348 3993
rect 3342 3988 3343 3992
rect 3347 3988 3348 3992
rect 3944 3990 3946 4017
rect 3342 3987 3348 3988
rect 3942 3989 3948 3990
rect 2046 3984 2052 3985
rect 3942 3985 3943 3989
rect 3947 3985 3948 3989
rect 3942 3984 3948 3985
rect 2146 3983 2152 3984
rect 2146 3979 2147 3983
rect 2151 3979 2152 3983
rect 2146 3978 2152 3979
rect 2194 3983 2200 3984
rect 2194 3979 2195 3983
rect 2199 3979 2200 3983
rect 2194 3978 2200 3979
rect 2666 3983 2672 3984
rect 2666 3979 2667 3983
rect 2671 3979 2672 3983
rect 2666 3978 2672 3979
rect 2914 3983 2920 3984
rect 2914 3979 2915 3983
rect 2919 3979 2920 3983
rect 2914 3978 2920 3979
rect 3162 3983 3168 3984
rect 3162 3979 3163 3983
rect 3167 3979 3168 3983
rect 3162 3978 3168 3979
rect 3242 3983 3248 3984
rect 3242 3979 3243 3983
rect 3247 3979 3248 3983
rect 3242 3978 3248 3979
rect 2070 3973 2076 3974
rect 2046 3972 2052 3973
rect 1902 3967 1908 3968
rect 2006 3969 2012 3970
rect 110 3964 116 3965
rect 2006 3965 2007 3969
rect 2011 3965 2012 3969
rect 2046 3968 2047 3972
rect 2051 3968 2052 3972
rect 2070 3969 2071 3973
rect 2075 3969 2076 3973
rect 2070 3968 2076 3969
rect 2046 3967 2052 3968
rect 2006 3964 2012 3965
rect 462 3963 468 3964
rect 462 3959 463 3963
rect 467 3959 468 3963
rect 462 3958 468 3959
rect 586 3963 592 3964
rect 586 3959 587 3963
rect 591 3959 592 3963
rect 586 3958 592 3959
rect 778 3963 784 3964
rect 778 3959 779 3963
rect 783 3959 784 3963
rect 778 3958 784 3959
rect 1138 3963 1144 3964
rect 1138 3959 1139 3963
rect 1143 3959 1144 3963
rect 1138 3958 1144 3959
rect 1306 3963 1312 3964
rect 1306 3959 1307 3963
rect 1311 3959 1312 3963
rect 1306 3958 1312 3959
rect 1458 3963 1464 3964
rect 1458 3959 1459 3963
rect 1463 3959 1464 3963
rect 1458 3958 1464 3959
rect 1594 3963 1600 3964
rect 1594 3959 1595 3963
rect 1599 3959 1600 3963
rect 1594 3958 1600 3959
rect 1730 3963 1736 3964
rect 1730 3959 1731 3963
rect 1735 3959 1736 3963
rect 1730 3958 1736 3959
rect 1866 3963 1872 3964
rect 1866 3959 1867 3963
rect 1871 3959 1872 3963
rect 1866 3958 1872 3959
rect 310 3953 316 3954
rect 110 3952 116 3953
rect 110 3948 111 3952
rect 115 3948 116 3952
rect 310 3949 311 3953
rect 315 3949 316 3953
rect 310 3948 316 3949
rect 110 3947 116 3948
rect 112 3927 114 3947
rect 312 3927 314 3948
rect 464 3932 466 3958
rect 510 3953 516 3954
rect 510 3949 511 3953
rect 515 3949 516 3953
rect 510 3948 516 3949
rect 402 3931 408 3932
rect 402 3927 403 3931
rect 407 3927 408 3931
rect 462 3931 468 3932
rect 462 3927 463 3931
rect 467 3927 468 3931
rect 512 3927 514 3948
rect 588 3932 590 3958
rect 702 3953 708 3954
rect 702 3949 703 3953
rect 707 3949 708 3953
rect 702 3948 708 3949
rect 634 3947 640 3948
rect 634 3943 635 3947
rect 639 3943 640 3947
rect 634 3942 640 3943
rect 586 3931 592 3932
rect 586 3927 587 3931
rect 591 3927 592 3931
rect 111 3926 115 3927
rect 111 3921 115 3922
rect 279 3926 283 3927
rect 279 3921 283 3922
rect 311 3926 315 3927
rect 402 3926 408 3927
rect 415 3926 419 3927
rect 462 3926 468 3927
rect 511 3926 515 3927
rect 311 3921 315 3922
rect 112 3901 114 3921
rect 110 3900 116 3901
rect 280 3900 282 3921
rect 302 3919 308 3920
rect 302 3915 303 3919
rect 307 3915 308 3919
rect 302 3914 308 3915
rect 354 3919 360 3920
rect 354 3915 355 3919
rect 359 3915 360 3919
rect 354 3914 360 3915
rect 110 3896 111 3900
rect 115 3896 116 3900
rect 110 3895 116 3896
rect 278 3899 284 3900
rect 278 3895 279 3899
rect 283 3895 284 3899
rect 278 3894 284 3895
rect 110 3883 116 3884
rect 110 3879 111 3883
rect 115 3879 116 3883
rect 110 3878 116 3879
rect 278 3880 284 3881
rect 112 3843 114 3878
rect 278 3876 279 3880
rect 283 3876 284 3880
rect 278 3875 284 3876
rect 280 3843 282 3875
rect 111 3842 115 3843
rect 111 3837 115 3838
rect 231 3842 235 3843
rect 231 3837 235 3838
rect 279 3842 283 3843
rect 279 3837 283 3838
rect 112 3810 114 3837
rect 232 3813 234 3837
rect 230 3812 236 3813
rect 110 3809 116 3810
rect 110 3805 111 3809
rect 115 3805 116 3809
rect 230 3808 231 3812
rect 235 3808 236 3812
rect 230 3807 236 3808
rect 110 3804 116 3805
rect 304 3804 306 3914
rect 356 3892 358 3914
rect 404 3892 406 3926
rect 415 3921 419 3922
rect 511 3921 515 3922
rect 567 3926 571 3927
rect 586 3926 592 3927
rect 567 3921 571 3922
rect 416 3900 418 3921
rect 568 3900 570 3921
rect 636 3920 638 3942
rect 704 3927 706 3948
rect 780 3932 782 3958
rect 886 3953 892 3954
rect 886 3949 887 3953
rect 891 3949 892 3953
rect 886 3948 892 3949
rect 1062 3953 1068 3954
rect 1062 3949 1063 3953
rect 1067 3949 1068 3953
rect 1062 3948 1068 3949
rect 778 3931 784 3932
rect 778 3927 779 3931
rect 783 3927 784 3931
rect 888 3927 890 3948
rect 1064 3927 1066 3948
rect 1140 3932 1142 3958
rect 1230 3953 1236 3954
rect 1230 3949 1231 3953
rect 1235 3949 1236 3953
rect 1230 3948 1236 3949
rect 1130 3931 1136 3932
rect 1130 3927 1131 3931
rect 1135 3927 1136 3931
rect 703 3926 707 3927
rect 703 3921 707 3922
rect 735 3926 739 3927
rect 778 3926 784 3927
rect 887 3926 891 3927
rect 735 3921 739 3922
rect 887 3921 891 3922
rect 911 3926 915 3927
rect 911 3921 915 3922
rect 1063 3926 1067 3927
rect 1063 3921 1067 3922
rect 1095 3926 1099 3927
rect 1130 3926 1136 3927
rect 1138 3931 1144 3932
rect 1138 3927 1139 3931
rect 1143 3927 1144 3931
rect 1232 3927 1234 3948
rect 1308 3932 1310 3958
rect 1382 3953 1388 3954
rect 1382 3949 1383 3953
rect 1387 3949 1388 3953
rect 1382 3948 1388 3949
rect 1306 3931 1312 3932
rect 1306 3927 1307 3931
rect 1311 3927 1312 3931
rect 1384 3927 1386 3948
rect 1460 3932 1462 3958
rect 1518 3953 1524 3954
rect 1518 3949 1519 3953
rect 1523 3949 1524 3953
rect 1518 3948 1524 3949
rect 1458 3931 1464 3932
rect 1458 3927 1459 3931
rect 1463 3927 1464 3931
rect 1520 3927 1522 3948
rect 1596 3932 1598 3958
rect 1654 3953 1660 3954
rect 1654 3949 1655 3953
rect 1659 3949 1660 3953
rect 1654 3948 1660 3949
rect 1594 3931 1600 3932
rect 1594 3927 1595 3931
rect 1599 3927 1600 3931
rect 1656 3927 1658 3948
rect 1732 3932 1734 3958
rect 1790 3953 1796 3954
rect 1790 3949 1791 3953
rect 1795 3949 1796 3953
rect 1790 3948 1796 3949
rect 1730 3931 1736 3932
rect 1730 3927 1731 3931
rect 1735 3927 1736 3931
rect 1792 3927 1794 3948
rect 1868 3932 1870 3958
rect 1902 3953 1908 3954
rect 1902 3949 1903 3953
rect 1907 3949 1908 3953
rect 1902 3948 1908 3949
rect 2006 3952 2012 3953
rect 2006 3948 2007 3952
rect 2011 3948 2012 3952
rect 1866 3931 1872 3932
rect 1866 3927 1867 3931
rect 1871 3927 1872 3931
rect 1904 3927 1906 3948
rect 2006 3947 2012 3948
rect 2048 3947 2050 3967
rect 2072 3947 2074 3968
rect 2148 3952 2150 3978
rect 2146 3951 2152 3952
rect 2146 3947 2147 3951
rect 2151 3947 2152 3951
rect 2008 3927 2010 3947
rect 2047 3946 2051 3947
rect 2047 3941 2051 3942
rect 2071 3946 2075 3947
rect 2071 3941 2075 3942
rect 2127 3946 2131 3947
rect 2146 3946 2152 3947
rect 2127 3941 2131 3942
rect 1138 3926 1144 3927
rect 1231 3926 1235 3927
rect 1095 3921 1099 3922
rect 634 3919 640 3920
rect 634 3915 635 3919
rect 639 3915 640 3919
rect 634 3914 640 3915
rect 642 3919 648 3920
rect 642 3915 643 3919
rect 647 3915 648 3919
rect 642 3914 648 3915
rect 414 3899 420 3900
rect 414 3895 415 3899
rect 419 3895 420 3899
rect 414 3894 420 3895
rect 566 3899 572 3900
rect 566 3895 567 3899
rect 571 3895 572 3899
rect 566 3894 572 3895
rect 644 3892 646 3914
rect 736 3900 738 3921
rect 810 3919 816 3920
rect 810 3915 811 3919
rect 815 3915 816 3919
rect 810 3914 816 3915
rect 734 3899 740 3900
rect 734 3895 735 3899
rect 739 3895 740 3899
rect 734 3894 740 3895
rect 812 3892 814 3914
rect 912 3900 914 3921
rect 986 3919 992 3920
rect 986 3915 987 3919
rect 991 3915 992 3919
rect 986 3914 992 3915
rect 910 3899 916 3900
rect 910 3895 911 3899
rect 915 3895 916 3899
rect 910 3894 916 3895
rect 988 3892 990 3914
rect 1096 3900 1098 3921
rect 1132 3908 1134 3926
rect 1231 3921 1235 3922
rect 1287 3926 1291 3927
rect 1306 3926 1312 3927
rect 1383 3926 1387 3927
rect 1458 3926 1464 3927
rect 1479 3926 1483 3927
rect 1287 3921 1291 3922
rect 1383 3921 1387 3922
rect 1479 3921 1483 3922
rect 1519 3926 1523 3927
rect 1594 3926 1600 3927
rect 1655 3926 1659 3927
rect 1519 3921 1523 3922
rect 1655 3921 1659 3922
rect 1679 3926 1683 3927
rect 1730 3926 1736 3927
rect 1791 3926 1795 3927
rect 1866 3926 1872 3927
rect 1903 3926 1907 3927
rect 1679 3921 1683 3922
rect 1791 3921 1795 3922
rect 1903 3921 1907 3922
rect 2007 3926 2011 3927
rect 2007 3921 2011 3922
rect 2048 3921 2050 3941
rect 1130 3907 1136 3908
rect 1130 3903 1131 3907
rect 1135 3903 1136 3907
rect 1130 3902 1136 3903
rect 1288 3900 1290 3921
rect 1370 3919 1376 3920
rect 1370 3915 1371 3919
rect 1375 3915 1376 3919
rect 1370 3914 1376 3915
rect 1094 3899 1100 3900
rect 1094 3895 1095 3899
rect 1099 3895 1100 3899
rect 1094 3894 1100 3895
rect 1286 3899 1292 3900
rect 1286 3895 1287 3899
rect 1291 3895 1292 3899
rect 1286 3894 1292 3895
rect 1372 3892 1374 3914
rect 1480 3900 1482 3921
rect 1680 3900 1682 3921
rect 1706 3919 1712 3920
rect 1706 3915 1707 3919
rect 1711 3915 1712 3919
rect 1706 3914 1712 3915
rect 1478 3899 1484 3900
rect 1478 3895 1479 3899
rect 1483 3895 1484 3899
rect 1478 3894 1484 3895
rect 1678 3899 1684 3900
rect 1678 3895 1679 3899
rect 1683 3895 1684 3899
rect 1678 3894 1684 3895
rect 354 3891 360 3892
rect 354 3887 355 3891
rect 359 3887 360 3891
rect 354 3886 360 3887
rect 402 3891 408 3892
rect 402 3887 403 3891
rect 407 3887 408 3891
rect 402 3886 408 3887
rect 642 3891 648 3892
rect 642 3887 643 3891
rect 647 3887 648 3891
rect 642 3886 648 3887
rect 810 3891 816 3892
rect 810 3887 811 3891
rect 815 3887 816 3891
rect 810 3886 816 3887
rect 986 3891 992 3892
rect 986 3887 987 3891
rect 991 3887 992 3891
rect 986 3886 992 3887
rect 1046 3891 1052 3892
rect 1046 3887 1047 3891
rect 1051 3887 1052 3891
rect 1046 3886 1052 3887
rect 1370 3891 1376 3892
rect 1370 3887 1371 3891
rect 1375 3887 1376 3891
rect 1370 3886 1376 3887
rect 414 3880 420 3881
rect 414 3876 415 3880
rect 419 3876 420 3880
rect 414 3875 420 3876
rect 566 3880 572 3881
rect 566 3876 567 3880
rect 571 3876 572 3880
rect 566 3875 572 3876
rect 734 3880 740 3881
rect 734 3876 735 3880
rect 739 3876 740 3880
rect 734 3875 740 3876
rect 910 3880 916 3881
rect 910 3876 911 3880
rect 915 3876 916 3880
rect 910 3875 916 3876
rect 416 3843 418 3875
rect 568 3843 570 3875
rect 736 3843 738 3875
rect 912 3843 914 3875
rect 335 3842 339 3843
rect 335 3837 339 3838
rect 415 3842 419 3843
rect 415 3837 419 3838
rect 439 3842 443 3843
rect 439 3837 443 3838
rect 535 3842 539 3843
rect 535 3837 539 3838
rect 567 3842 571 3843
rect 567 3837 571 3838
rect 631 3842 635 3843
rect 631 3837 635 3838
rect 727 3842 731 3843
rect 727 3837 731 3838
rect 735 3842 739 3843
rect 735 3837 739 3838
rect 831 3842 835 3843
rect 831 3837 835 3838
rect 911 3842 915 3843
rect 911 3837 915 3838
rect 935 3842 939 3843
rect 935 3837 939 3838
rect 1039 3842 1043 3843
rect 1039 3837 1043 3838
rect 336 3813 338 3837
rect 440 3813 442 3837
rect 536 3813 538 3837
rect 632 3813 634 3837
rect 728 3813 730 3837
rect 832 3813 834 3837
rect 936 3813 938 3837
rect 1040 3813 1042 3837
rect 334 3812 340 3813
rect 334 3808 335 3812
rect 339 3808 340 3812
rect 334 3807 340 3808
rect 438 3812 444 3813
rect 438 3808 439 3812
rect 443 3808 444 3812
rect 438 3807 444 3808
rect 534 3812 540 3813
rect 534 3808 535 3812
rect 539 3808 540 3812
rect 534 3807 540 3808
rect 630 3812 636 3813
rect 630 3808 631 3812
rect 635 3808 636 3812
rect 630 3807 636 3808
rect 726 3812 732 3813
rect 726 3808 727 3812
rect 731 3808 732 3812
rect 726 3807 732 3808
rect 830 3812 836 3813
rect 830 3808 831 3812
rect 835 3808 836 3812
rect 830 3807 836 3808
rect 934 3812 940 3813
rect 934 3808 935 3812
rect 939 3808 940 3812
rect 934 3807 940 3808
rect 1038 3812 1044 3813
rect 1038 3808 1039 3812
rect 1043 3808 1044 3812
rect 1038 3807 1044 3808
rect 302 3803 308 3804
rect 302 3799 303 3803
rect 307 3799 308 3803
rect 302 3798 308 3799
rect 314 3803 320 3804
rect 314 3799 315 3803
rect 319 3799 320 3803
rect 314 3798 320 3799
rect 514 3803 520 3804
rect 514 3799 515 3803
rect 519 3799 520 3803
rect 514 3798 520 3799
rect 610 3803 616 3804
rect 610 3799 611 3803
rect 615 3799 616 3803
rect 610 3798 616 3799
rect 706 3803 712 3804
rect 706 3799 707 3803
rect 711 3799 712 3803
rect 706 3798 712 3799
rect 802 3803 808 3804
rect 802 3799 803 3803
rect 807 3799 808 3803
rect 802 3798 808 3799
rect 906 3803 912 3804
rect 906 3799 907 3803
rect 911 3799 912 3803
rect 906 3798 912 3799
rect 1010 3803 1016 3804
rect 1010 3799 1011 3803
rect 1015 3799 1016 3803
rect 1010 3798 1016 3799
rect 230 3793 236 3794
rect 110 3792 116 3793
rect 110 3788 111 3792
rect 115 3788 116 3792
rect 230 3789 231 3793
rect 235 3789 236 3793
rect 230 3788 236 3789
rect 110 3787 116 3788
rect 112 3767 114 3787
rect 232 3767 234 3788
rect 316 3772 318 3798
rect 334 3793 340 3794
rect 334 3789 335 3793
rect 339 3789 340 3793
rect 334 3788 340 3789
rect 438 3793 444 3794
rect 438 3789 439 3793
rect 443 3789 444 3793
rect 438 3788 444 3789
rect 314 3771 320 3772
rect 314 3767 315 3771
rect 319 3767 320 3771
rect 336 3767 338 3788
rect 440 3767 442 3788
rect 516 3772 518 3798
rect 534 3793 540 3794
rect 534 3789 535 3793
rect 539 3789 540 3793
rect 534 3788 540 3789
rect 514 3771 520 3772
rect 514 3767 515 3771
rect 519 3767 520 3771
rect 536 3767 538 3788
rect 612 3772 614 3798
rect 630 3793 636 3794
rect 630 3789 631 3793
rect 635 3789 636 3793
rect 630 3788 636 3789
rect 610 3771 616 3772
rect 610 3767 611 3771
rect 615 3767 616 3771
rect 632 3767 634 3788
rect 708 3772 710 3798
rect 726 3793 732 3794
rect 726 3789 727 3793
rect 731 3789 732 3793
rect 726 3788 732 3789
rect 706 3771 712 3772
rect 706 3767 707 3771
rect 711 3767 712 3771
rect 728 3767 730 3788
rect 804 3772 806 3798
rect 830 3793 836 3794
rect 830 3789 831 3793
rect 835 3789 836 3793
rect 830 3788 836 3789
rect 818 3787 824 3788
rect 818 3783 819 3787
rect 823 3783 824 3787
rect 818 3782 824 3783
rect 802 3771 808 3772
rect 802 3767 803 3771
rect 807 3767 808 3771
rect 111 3766 115 3767
rect 111 3761 115 3762
rect 159 3766 163 3767
rect 159 3761 163 3762
rect 231 3766 235 3767
rect 314 3766 320 3767
rect 335 3766 339 3767
rect 231 3761 235 3762
rect 335 3761 339 3762
rect 351 3766 355 3767
rect 351 3761 355 3762
rect 439 3766 443 3767
rect 514 3766 520 3767
rect 535 3766 539 3767
rect 439 3761 443 3762
rect 535 3761 539 3762
rect 551 3766 555 3767
rect 610 3766 616 3767
rect 631 3766 635 3767
rect 706 3766 712 3767
rect 727 3766 731 3767
rect 551 3761 555 3762
rect 631 3761 635 3762
rect 727 3761 731 3762
rect 751 3766 755 3767
rect 802 3766 808 3767
rect 751 3761 755 3762
rect 112 3741 114 3761
rect 110 3740 116 3741
rect 160 3740 162 3761
rect 222 3759 228 3760
rect 222 3755 223 3759
rect 227 3755 228 3759
rect 222 3754 228 3755
rect 258 3759 264 3760
rect 258 3755 259 3759
rect 263 3755 264 3759
rect 258 3754 264 3755
rect 110 3736 111 3740
rect 115 3736 116 3740
rect 110 3735 116 3736
rect 158 3739 164 3740
rect 158 3735 159 3739
rect 163 3735 164 3739
rect 158 3734 164 3735
rect 110 3723 116 3724
rect 110 3719 111 3723
rect 115 3719 116 3723
rect 110 3718 116 3719
rect 158 3720 164 3721
rect 112 3683 114 3718
rect 158 3716 159 3720
rect 163 3716 164 3720
rect 158 3715 164 3716
rect 160 3683 162 3715
rect 111 3682 115 3683
rect 111 3677 115 3678
rect 151 3682 155 3683
rect 151 3677 155 3678
rect 159 3682 163 3683
rect 159 3677 163 3678
rect 112 3650 114 3677
rect 152 3653 154 3677
rect 150 3652 156 3653
rect 110 3649 116 3650
rect 110 3645 111 3649
rect 115 3645 116 3649
rect 150 3648 151 3652
rect 155 3648 156 3652
rect 150 3647 156 3648
rect 110 3644 116 3645
rect 224 3644 226 3754
rect 260 3732 262 3754
rect 352 3740 354 3761
rect 426 3759 432 3760
rect 426 3755 427 3759
rect 431 3755 432 3759
rect 426 3754 432 3755
rect 350 3739 356 3740
rect 350 3735 351 3739
rect 355 3735 356 3739
rect 350 3734 356 3735
rect 428 3732 430 3754
rect 552 3740 554 3761
rect 752 3740 754 3761
rect 820 3760 822 3782
rect 832 3767 834 3788
rect 908 3772 910 3798
rect 934 3793 940 3794
rect 934 3789 935 3793
rect 939 3789 940 3793
rect 934 3788 940 3789
rect 906 3771 912 3772
rect 906 3767 907 3771
rect 911 3767 912 3771
rect 936 3767 938 3788
rect 1012 3772 1014 3798
rect 1038 3793 1044 3794
rect 1038 3789 1039 3793
rect 1043 3789 1044 3793
rect 1038 3788 1044 3789
rect 1010 3771 1016 3772
rect 1010 3767 1011 3771
rect 1015 3767 1016 3771
rect 1040 3767 1042 3788
rect 1048 3780 1050 3886
rect 1094 3880 1100 3881
rect 1094 3876 1095 3880
rect 1099 3876 1100 3880
rect 1094 3875 1100 3876
rect 1286 3880 1292 3881
rect 1286 3876 1287 3880
rect 1291 3876 1292 3880
rect 1286 3875 1292 3876
rect 1478 3880 1484 3881
rect 1478 3876 1479 3880
rect 1483 3876 1484 3880
rect 1478 3875 1484 3876
rect 1678 3880 1684 3881
rect 1678 3876 1679 3880
rect 1683 3876 1684 3880
rect 1678 3875 1684 3876
rect 1096 3843 1098 3875
rect 1288 3843 1290 3875
rect 1480 3843 1482 3875
rect 1680 3843 1682 3875
rect 1095 3842 1099 3843
rect 1095 3837 1099 3838
rect 1151 3842 1155 3843
rect 1151 3837 1155 3838
rect 1263 3842 1267 3843
rect 1263 3837 1267 3838
rect 1287 3842 1291 3843
rect 1287 3837 1291 3838
rect 1383 3842 1387 3843
rect 1383 3837 1387 3838
rect 1479 3842 1483 3843
rect 1479 3837 1483 3838
rect 1503 3842 1507 3843
rect 1503 3837 1507 3838
rect 1631 3842 1635 3843
rect 1631 3837 1635 3838
rect 1679 3842 1683 3843
rect 1679 3837 1683 3838
rect 1152 3813 1154 3837
rect 1264 3813 1266 3837
rect 1384 3813 1386 3837
rect 1504 3813 1506 3837
rect 1632 3813 1634 3837
rect 1150 3812 1156 3813
rect 1150 3808 1151 3812
rect 1155 3808 1156 3812
rect 1150 3807 1156 3808
rect 1262 3812 1268 3813
rect 1262 3808 1263 3812
rect 1267 3808 1268 3812
rect 1262 3807 1268 3808
rect 1382 3812 1388 3813
rect 1382 3808 1383 3812
rect 1387 3808 1388 3812
rect 1382 3807 1388 3808
rect 1502 3812 1508 3813
rect 1502 3808 1503 3812
rect 1507 3808 1508 3812
rect 1502 3807 1508 3808
rect 1630 3812 1636 3813
rect 1630 3808 1631 3812
rect 1635 3808 1636 3812
rect 1630 3807 1636 3808
rect 1708 3804 1710 3914
rect 2008 3901 2010 3921
rect 2046 3920 2052 3921
rect 2128 3920 2130 3941
rect 2196 3940 2198 3978
rect 2326 3973 2332 3974
rect 2326 3969 2327 3973
rect 2331 3969 2332 3973
rect 2326 3968 2332 3969
rect 2590 3973 2596 3974
rect 2590 3969 2591 3973
rect 2595 3969 2596 3973
rect 2590 3968 2596 3969
rect 2328 3947 2330 3968
rect 2592 3947 2594 3968
rect 2668 3952 2670 3978
rect 2838 3973 2844 3974
rect 2838 3969 2839 3973
rect 2843 3969 2844 3973
rect 2838 3968 2844 3969
rect 2658 3951 2664 3952
rect 2658 3947 2659 3951
rect 2663 3947 2664 3951
rect 2271 3946 2275 3947
rect 2271 3941 2275 3942
rect 2327 3946 2331 3947
rect 2327 3941 2331 3942
rect 2439 3946 2443 3947
rect 2439 3941 2443 3942
rect 2591 3946 2595 3947
rect 2591 3941 2595 3942
rect 2615 3946 2619 3947
rect 2658 3946 2664 3947
rect 2666 3951 2672 3952
rect 2666 3947 2667 3951
rect 2671 3947 2672 3951
rect 2840 3947 2842 3968
rect 2916 3952 2918 3978
rect 3086 3973 3092 3974
rect 3086 3969 3087 3973
rect 3091 3969 3092 3973
rect 3086 3968 3092 3969
rect 2914 3951 2920 3952
rect 2914 3947 2915 3951
rect 2919 3947 2920 3951
rect 3088 3947 3090 3968
rect 3164 3952 3166 3978
rect 3162 3951 3168 3952
rect 3162 3947 3163 3951
rect 3167 3947 3168 3951
rect 2666 3946 2672 3947
rect 2799 3946 2803 3947
rect 2615 3941 2619 3942
rect 2194 3939 2200 3940
rect 2194 3935 2195 3939
rect 2199 3935 2200 3939
rect 2194 3934 2200 3935
rect 2202 3939 2208 3940
rect 2202 3935 2203 3939
rect 2207 3935 2208 3939
rect 2202 3934 2208 3935
rect 2046 3916 2047 3920
rect 2051 3916 2052 3920
rect 2046 3915 2052 3916
rect 2126 3919 2132 3920
rect 2126 3915 2127 3919
rect 2131 3915 2132 3919
rect 2126 3914 2132 3915
rect 2204 3912 2206 3934
rect 2272 3920 2274 3941
rect 2346 3939 2352 3940
rect 2346 3935 2347 3939
rect 2351 3935 2352 3939
rect 2346 3934 2352 3935
rect 2270 3919 2276 3920
rect 2270 3915 2271 3919
rect 2275 3915 2276 3919
rect 2270 3914 2276 3915
rect 2348 3912 2350 3934
rect 2440 3920 2442 3941
rect 2514 3939 2520 3940
rect 2514 3935 2515 3939
rect 2519 3935 2520 3939
rect 2514 3934 2520 3935
rect 2438 3919 2444 3920
rect 2438 3915 2439 3919
rect 2443 3915 2444 3919
rect 2438 3914 2444 3915
rect 2516 3912 2518 3934
rect 2616 3920 2618 3941
rect 2660 3928 2662 3946
rect 2799 3941 2803 3942
rect 2839 3946 2843 3947
rect 2914 3946 2920 3947
rect 2983 3946 2987 3947
rect 2839 3941 2843 3942
rect 2983 3941 2987 3942
rect 3087 3946 3091 3947
rect 3162 3946 3168 3947
rect 3175 3946 3179 3947
rect 3087 3941 3091 3942
rect 3175 3941 3179 3942
rect 2690 3939 2696 3940
rect 2690 3935 2691 3939
rect 2695 3935 2696 3939
rect 2690 3934 2696 3935
rect 2658 3927 2664 3928
rect 2658 3923 2659 3927
rect 2663 3923 2664 3927
rect 2658 3922 2664 3923
rect 2614 3919 2620 3920
rect 2614 3915 2615 3919
rect 2619 3915 2620 3919
rect 2614 3914 2620 3915
rect 2692 3912 2694 3934
rect 2800 3920 2802 3941
rect 2984 3920 2986 3941
rect 3050 3939 3056 3940
rect 3050 3935 3051 3939
rect 3055 3935 3056 3939
rect 3050 3934 3056 3935
rect 2798 3919 2804 3920
rect 2798 3915 2799 3919
rect 2803 3915 2804 3919
rect 2798 3914 2804 3915
rect 2982 3919 2988 3920
rect 2982 3915 2983 3919
rect 2987 3915 2988 3919
rect 2982 3914 2988 3915
rect 2202 3911 2208 3912
rect 2202 3907 2203 3911
rect 2207 3907 2208 3911
rect 2202 3906 2208 3907
rect 2346 3911 2352 3912
rect 2346 3907 2347 3911
rect 2351 3907 2352 3911
rect 2346 3906 2352 3907
rect 2514 3911 2520 3912
rect 2514 3907 2515 3911
rect 2519 3907 2520 3911
rect 2514 3906 2520 3907
rect 2690 3911 2696 3912
rect 2690 3907 2691 3911
rect 2695 3907 2696 3911
rect 2690 3906 2696 3907
rect 2874 3907 2880 3908
rect 2046 3903 2052 3904
rect 2006 3900 2012 3901
rect 2006 3896 2007 3900
rect 2011 3896 2012 3900
rect 2046 3899 2047 3903
rect 2051 3899 2052 3903
rect 2874 3903 2875 3907
rect 2879 3903 2880 3907
rect 2874 3902 2880 3903
rect 2046 3898 2052 3899
rect 2126 3900 2132 3901
rect 2006 3895 2012 3896
rect 2006 3883 2012 3884
rect 2006 3879 2007 3883
rect 2011 3879 2012 3883
rect 2006 3878 2012 3879
rect 2008 3843 2010 3878
rect 2048 3871 2050 3898
rect 2126 3896 2127 3900
rect 2131 3896 2132 3900
rect 2126 3895 2132 3896
rect 2270 3900 2276 3901
rect 2270 3896 2271 3900
rect 2275 3896 2276 3900
rect 2270 3895 2276 3896
rect 2438 3900 2444 3901
rect 2438 3896 2439 3900
rect 2443 3896 2444 3900
rect 2438 3895 2444 3896
rect 2614 3900 2620 3901
rect 2614 3896 2615 3900
rect 2619 3896 2620 3900
rect 2614 3895 2620 3896
rect 2798 3900 2804 3901
rect 2798 3896 2799 3900
rect 2803 3896 2804 3900
rect 2798 3895 2804 3896
rect 2128 3871 2130 3895
rect 2272 3871 2274 3895
rect 2440 3871 2442 3895
rect 2616 3871 2618 3895
rect 2800 3871 2802 3895
rect 2047 3870 2051 3871
rect 2047 3865 2051 3866
rect 2127 3870 2131 3871
rect 2127 3865 2131 3866
rect 2263 3870 2267 3871
rect 2263 3865 2267 3866
rect 2271 3870 2275 3871
rect 2271 3865 2275 3866
rect 2375 3870 2379 3871
rect 2375 3865 2379 3866
rect 2439 3870 2443 3871
rect 2439 3865 2443 3866
rect 2495 3870 2499 3871
rect 2495 3865 2499 3866
rect 2615 3870 2619 3871
rect 2615 3865 2619 3866
rect 2631 3870 2635 3871
rect 2631 3865 2635 3866
rect 2775 3870 2779 3871
rect 2775 3865 2779 3866
rect 2799 3870 2803 3871
rect 2799 3865 2803 3866
rect 2007 3842 2011 3843
rect 2048 3838 2050 3865
rect 2264 3841 2266 3865
rect 2376 3841 2378 3865
rect 2496 3841 2498 3865
rect 2632 3841 2634 3865
rect 2776 3841 2778 3865
rect 2262 3840 2268 3841
rect 2007 3837 2011 3838
rect 2046 3837 2052 3838
rect 2008 3810 2010 3837
rect 2046 3833 2047 3837
rect 2051 3833 2052 3837
rect 2262 3836 2263 3840
rect 2267 3836 2268 3840
rect 2262 3835 2268 3836
rect 2374 3840 2380 3841
rect 2374 3836 2375 3840
rect 2379 3836 2380 3840
rect 2374 3835 2380 3836
rect 2494 3840 2500 3841
rect 2494 3836 2495 3840
rect 2499 3836 2500 3840
rect 2494 3835 2500 3836
rect 2630 3840 2636 3841
rect 2630 3836 2631 3840
rect 2635 3836 2636 3840
rect 2630 3835 2636 3836
rect 2774 3840 2780 3841
rect 2774 3836 2775 3840
rect 2779 3836 2780 3840
rect 2774 3835 2780 3836
rect 2046 3832 2052 3833
rect 2338 3831 2344 3832
rect 2338 3827 2339 3831
rect 2343 3827 2344 3831
rect 2338 3826 2344 3827
rect 2450 3831 2456 3832
rect 2450 3827 2451 3831
rect 2455 3827 2456 3831
rect 2450 3826 2456 3827
rect 2458 3831 2464 3832
rect 2458 3827 2459 3831
rect 2463 3827 2464 3831
rect 2458 3826 2464 3827
rect 2578 3831 2584 3832
rect 2578 3827 2579 3831
rect 2583 3827 2584 3831
rect 2578 3826 2584 3827
rect 2714 3831 2720 3832
rect 2714 3827 2715 3831
rect 2719 3827 2720 3831
rect 2714 3826 2720 3827
rect 2262 3821 2268 3822
rect 2046 3820 2052 3821
rect 2046 3816 2047 3820
rect 2051 3816 2052 3820
rect 2262 3817 2263 3821
rect 2267 3817 2268 3821
rect 2262 3816 2268 3817
rect 2046 3815 2052 3816
rect 2006 3809 2012 3810
rect 2006 3805 2007 3809
rect 2011 3805 2012 3809
rect 2006 3804 2012 3805
rect 1114 3803 1120 3804
rect 1114 3799 1115 3803
rect 1119 3799 1120 3803
rect 1114 3798 1120 3799
rect 1226 3803 1232 3804
rect 1226 3799 1227 3803
rect 1231 3799 1232 3803
rect 1226 3798 1232 3799
rect 1338 3803 1344 3804
rect 1338 3799 1339 3803
rect 1343 3799 1344 3803
rect 1338 3798 1344 3799
rect 1618 3803 1624 3804
rect 1618 3799 1619 3803
rect 1623 3799 1624 3803
rect 1618 3798 1624 3799
rect 1706 3803 1712 3804
rect 1706 3799 1707 3803
rect 1711 3799 1712 3803
rect 1706 3798 1712 3799
rect 1046 3779 1052 3780
rect 1046 3775 1047 3779
rect 1051 3775 1052 3779
rect 1046 3774 1052 3775
rect 1116 3772 1118 3798
rect 1150 3793 1156 3794
rect 1150 3789 1151 3793
rect 1155 3789 1156 3793
rect 1150 3788 1156 3789
rect 1114 3771 1120 3772
rect 1114 3767 1115 3771
rect 1119 3767 1120 3771
rect 1152 3767 1154 3788
rect 1228 3772 1230 3798
rect 1262 3793 1268 3794
rect 1262 3789 1263 3793
rect 1267 3789 1268 3793
rect 1262 3788 1268 3789
rect 1226 3771 1232 3772
rect 1226 3767 1227 3771
rect 1231 3767 1232 3771
rect 1264 3767 1266 3788
rect 1340 3772 1342 3798
rect 1382 3793 1388 3794
rect 1382 3789 1383 3793
rect 1387 3789 1388 3793
rect 1382 3788 1388 3789
rect 1502 3793 1508 3794
rect 1502 3789 1503 3793
rect 1507 3789 1508 3793
rect 1502 3788 1508 3789
rect 1338 3771 1344 3772
rect 1338 3767 1339 3771
rect 1343 3767 1344 3771
rect 1384 3767 1386 3788
rect 1504 3767 1506 3788
rect 1620 3772 1622 3798
rect 1630 3793 1636 3794
rect 1630 3789 1631 3793
rect 1635 3789 1636 3793
rect 1630 3788 1636 3789
rect 2006 3792 2012 3793
rect 2006 3788 2007 3792
rect 2011 3788 2012 3792
rect 1618 3771 1624 3772
rect 1618 3767 1619 3771
rect 1623 3767 1624 3771
rect 1632 3767 1634 3788
rect 2006 3787 2012 3788
rect 2008 3767 2010 3787
rect 2048 3779 2050 3815
rect 2264 3779 2266 3816
rect 2340 3800 2342 3826
rect 2374 3821 2380 3822
rect 2374 3817 2375 3821
rect 2379 3817 2380 3821
rect 2374 3816 2380 3817
rect 2338 3799 2344 3800
rect 2338 3795 2339 3799
rect 2343 3795 2344 3799
rect 2338 3794 2344 3795
rect 2376 3779 2378 3816
rect 2047 3778 2051 3779
rect 2047 3773 2051 3774
rect 2071 3778 2075 3779
rect 2071 3773 2075 3774
rect 2183 3778 2187 3779
rect 2183 3773 2187 3774
rect 2263 3778 2267 3779
rect 2263 3773 2267 3774
rect 2327 3778 2331 3779
rect 2327 3773 2331 3774
rect 2375 3778 2379 3779
rect 2375 3773 2379 3774
rect 831 3766 835 3767
rect 906 3766 912 3767
rect 935 3766 939 3767
rect 831 3761 835 3762
rect 935 3761 939 3762
rect 959 3766 963 3767
rect 1010 3766 1016 3767
rect 1039 3766 1043 3767
rect 1114 3766 1120 3767
rect 1151 3766 1155 3767
rect 959 3761 963 3762
rect 1039 3761 1043 3762
rect 1151 3761 1155 3762
rect 1167 3766 1171 3767
rect 1226 3766 1232 3767
rect 1263 3766 1267 3767
rect 1338 3766 1344 3767
rect 1383 3766 1387 3767
rect 1167 3761 1171 3762
rect 1263 3761 1267 3762
rect 1383 3761 1387 3762
rect 1503 3766 1507 3767
rect 1503 3761 1507 3762
rect 1607 3766 1611 3767
rect 1618 3766 1624 3767
rect 1631 3766 1635 3767
rect 1607 3761 1611 3762
rect 1631 3761 1635 3762
rect 2007 3766 2011 3767
rect 2007 3761 2011 3762
rect 818 3759 824 3760
rect 818 3755 819 3759
rect 823 3755 824 3759
rect 818 3754 824 3755
rect 906 3759 912 3760
rect 906 3755 907 3759
rect 911 3755 912 3759
rect 906 3754 912 3755
rect 550 3739 556 3740
rect 550 3735 551 3739
rect 555 3735 556 3739
rect 550 3734 556 3735
rect 750 3739 756 3740
rect 750 3735 751 3739
rect 755 3735 756 3739
rect 750 3734 756 3735
rect 908 3732 910 3754
rect 960 3740 962 3761
rect 1078 3759 1084 3760
rect 1078 3755 1079 3759
rect 1083 3755 1084 3759
rect 1078 3754 1084 3755
rect 958 3739 964 3740
rect 958 3735 959 3739
rect 963 3735 964 3739
rect 958 3734 964 3735
rect 1080 3732 1082 3754
rect 1168 3740 1170 3761
rect 1242 3759 1248 3760
rect 1242 3755 1243 3759
rect 1247 3755 1248 3759
rect 1242 3754 1248 3755
rect 1166 3739 1172 3740
rect 1166 3735 1167 3739
rect 1171 3735 1172 3739
rect 1166 3734 1172 3735
rect 1244 3732 1246 3754
rect 1384 3740 1386 3761
rect 1554 3759 1560 3760
rect 1554 3755 1555 3759
rect 1559 3755 1560 3759
rect 1554 3754 1560 3755
rect 1382 3739 1388 3740
rect 1382 3735 1383 3739
rect 1387 3735 1388 3739
rect 1382 3734 1388 3735
rect 258 3731 264 3732
rect 258 3727 259 3731
rect 263 3727 264 3731
rect 258 3726 264 3727
rect 426 3731 432 3732
rect 426 3727 427 3731
rect 431 3727 432 3731
rect 426 3726 432 3727
rect 906 3731 912 3732
rect 906 3727 907 3731
rect 911 3727 912 3731
rect 906 3726 912 3727
rect 1078 3731 1084 3732
rect 1078 3727 1079 3731
rect 1083 3727 1084 3731
rect 1078 3726 1084 3727
rect 1242 3731 1248 3732
rect 1242 3727 1243 3731
rect 1247 3727 1248 3731
rect 1242 3726 1248 3727
rect 1346 3731 1352 3732
rect 1346 3727 1347 3731
rect 1351 3727 1352 3731
rect 1346 3726 1352 3727
rect 350 3720 356 3721
rect 350 3716 351 3720
rect 355 3716 356 3720
rect 350 3715 356 3716
rect 550 3720 556 3721
rect 550 3716 551 3720
rect 555 3716 556 3720
rect 550 3715 556 3716
rect 750 3720 756 3721
rect 750 3716 751 3720
rect 755 3716 756 3720
rect 750 3715 756 3716
rect 958 3720 964 3721
rect 958 3716 959 3720
rect 963 3716 964 3720
rect 958 3715 964 3716
rect 1166 3720 1172 3721
rect 1166 3716 1167 3720
rect 1171 3716 1172 3720
rect 1166 3715 1172 3716
rect 352 3683 354 3715
rect 552 3683 554 3715
rect 752 3683 754 3715
rect 960 3683 962 3715
rect 1168 3683 1170 3715
rect 351 3682 355 3683
rect 351 3677 355 3678
rect 383 3682 387 3683
rect 383 3677 387 3678
rect 551 3682 555 3683
rect 551 3677 555 3678
rect 615 3682 619 3683
rect 615 3677 619 3678
rect 751 3682 755 3683
rect 751 3677 755 3678
rect 839 3682 843 3683
rect 839 3677 843 3678
rect 959 3682 963 3683
rect 959 3677 963 3678
rect 1055 3682 1059 3683
rect 1055 3677 1059 3678
rect 1167 3682 1171 3683
rect 1167 3677 1171 3678
rect 1263 3682 1267 3683
rect 1263 3677 1267 3678
rect 384 3653 386 3677
rect 616 3653 618 3677
rect 840 3653 842 3677
rect 1056 3653 1058 3677
rect 1264 3653 1266 3677
rect 382 3652 388 3653
rect 382 3648 383 3652
rect 387 3648 388 3652
rect 382 3647 388 3648
rect 614 3652 620 3653
rect 614 3648 615 3652
rect 619 3648 620 3652
rect 614 3647 620 3648
rect 838 3652 844 3653
rect 838 3648 839 3652
rect 843 3648 844 3652
rect 838 3647 844 3648
rect 1054 3652 1060 3653
rect 1054 3648 1055 3652
rect 1059 3648 1060 3652
rect 1054 3647 1060 3648
rect 1262 3652 1268 3653
rect 1262 3648 1263 3652
rect 1267 3648 1268 3652
rect 1262 3647 1268 3648
rect 222 3643 228 3644
rect 222 3639 223 3643
rect 227 3639 228 3643
rect 222 3638 228 3639
rect 234 3643 240 3644
rect 234 3639 235 3643
rect 239 3639 240 3643
rect 234 3638 240 3639
rect 466 3643 472 3644
rect 466 3639 467 3643
rect 471 3639 472 3643
rect 466 3638 472 3639
rect 1038 3643 1044 3644
rect 1038 3639 1039 3643
rect 1043 3639 1044 3643
rect 1038 3638 1044 3639
rect 1130 3643 1136 3644
rect 1130 3639 1131 3643
rect 1135 3639 1136 3643
rect 1130 3638 1136 3639
rect 1338 3643 1344 3644
rect 1338 3639 1339 3643
rect 1343 3639 1344 3643
rect 1338 3638 1344 3639
rect 150 3633 156 3634
rect 110 3632 116 3633
rect 110 3628 111 3632
rect 115 3628 116 3632
rect 150 3629 151 3633
rect 155 3629 156 3633
rect 150 3628 156 3629
rect 110 3627 116 3628
rect 112 3603 114 3627
rect 152 3603 154 3628
rect 236 3612 238 3638
rect 382 3633 388 3634
rect 382 3629 383 3633
rect 387 3629 388 3633
rect 382 3628 388 3629
rect 234 3611 240 3612
rect 234 3607 235 3611
rect 239 3607 240 3611
rect 234 3606 240 3607
rect 384 3603 386 3628
rect 468 3612 470 3638
rect 614 3633 620 3634
rect 614 3629 615 3633
rect 619 3629 620 3633
rect 614 3628 620 3629
rect 838 3633 844 3634
rect 838 3629 839 3633
rect 843 3629 844 3633
rect 838 3628 844 3629
rect 466 3611 472 3612
rect 466 3607 467 3611
rect 471 3607 472 3611
rect 466 3606 472 3607
rect 616 3603 618 3628
rect 682 3611 688 3612
rect 682 3607 683 3611
rect 687 3607 688 3611
rect 682 3606 688 3607
rect 111 3602 115 3603
rect 111 3597 115 3598
rect 151 3602 155 3603
rect 151 3597 155 3598
rect 167 3602 171 3603
rect 167 3597 171 3598
rect 359 3602 363 3603
rect 359 3597 363 3598
rect 383 3602 387 3603
rect 383 3597 387 3598
rect 559 3602 563 3603
rect 559 3597 563 3598
rect 615 3602 619 3603
rect 615 3597 619 3598
rect 112 3577 114 3597
rect 110 3576 116 3577
rect 168 3576 170 3597
rect 242 3595 248 3596
rect 242 3591 243 3595
rect 247 3591 248 3595
rect 242 3590 248 3591
rect 110 3572 111 3576
rect 115 3572 116 3576
rect 110 3571 116 3572
rect 166 3575 172 3576
rect 166 3571 167 3575
rect 171 3571 172 3575
rect 166 3570 172 3571
rect 244 3568 246 3590
rect 360 3576 362 3597
rect 434 3595 440 3596
rect 434 3591 435 3595
rect 439 3591 440 3595
rect 434 3590 440 3591
rect 358 3575 364 3576
rect 358 3571 359 3575
rect 363 3571 364 3575
rect 358 3570 364 3571
rect 436 3568 438 3590
rect 560 3576 562 3597
rect 634 3595 640 3596
rect 634 3591 635 3595
rect 639 3591 640 3595
rect 634 3590 640 3591
rect 558 3575 564 3576
rect 558 3571 559 3575
rect 563 3571 564 3575
rect 558 3570 564 3571
rect 636 3568 638 3590
rect 684 3568 686 3606
rect 840 3603 842 3628
rect 1040 3612 1042 3638
rect 1054 3633 1060 3634
rect 1054 3629 1055 3633
rect 1059 3629 1060 3633
rect 1054 3628 1060 3629
rect 1038 3611 1044 3612
rect 1038 3607 1039 3611
rect 1043 3607 1044 3611
rect 1038 3606 1044 3607
rect 1056 3603 1058 3628
rect 1132 3612 1134 3638
rect 1262 3633 1268 3634
rect 1262 3629 1263 3633
rect 1267 3629 1268 3633
rect 1262 3628 1268 3629
rect 1130 3611 1136 3612
rect 1130 3607 1131 3611
rect 1135 3607 1136 3611
rect 1130 3606 1136 3607
rect 1264 3603 1266 3628
rect 775 3602 779 3603
rect 775 3597 779 3598
rect 839 3602 843 3603
rect 839 3597 843 3598
rect 991 3602 995 3603
rect 991 3597 995 3598
rect 1055 3602 1059 3603
rect 1055 3597 1059 3598
rect 1215 3602 1219 3603
rect 1215 3597 1219 3598
rect 1263 3602 1267 3603
rect 1263 3597 1267 3598
rect 776 3576 778 3597
rect 992 3576 994 3597
rect 1216 3576 1218 3597
rect 1340 3596 1342 3638
rect 1348 3620 1350 3726
rect 1382 3720 1388 3721
rect 1382 3716 1383 3720
rect 1387 3716 1388 3720
rect 1382 3715 1388 3716
rect 1384 3683 1386 3715
rect 1383 3682 1387 3683
rect 1383 3677 1387 3678
rect 1479 3682 1483 3683
rect 1479 3677 1483 3678
rect 1480 3653 1482 3677
rect 1478 3652 1484 3653
rect 1478 3648 1479 3652
rect 1483 3648 1484 3652
rect 1478 3647 1484 3648
rect 1556 3644 1558 3754
rect 1608 3740 1610 3761
rect 2008 3741 2010 3761
rect 2048 3753 2050 3773
rect 2046 3752 2052 3753
rect 2072 3752 2074 3773
rect 2154 3771 2160 3772
rect 2154 3767 2155 3771
rect 2159 3767 2160 3771
rect 2154 3766 2160 3767
rect 2046 3748 2047 3752
rect 2051 3748 2052 3752
rect 2046 3747 2052 3748
rect 2070 3751 2076 3752
rect 2070 3747 2071 3751
rect 2075 3747 2076 3751
rect 2070 3746 2076 3747
rect 2156 3744 2158 3766
rect 2184 3752 2186 3773
rect 2328 3752 2330 3773
rect 2452 3772 2454 3826
rect 2460 3808 2462 3826
rect 2494 3821 2500 3822
rect 2494 3817 2495 3821
rect 2499 3817 2500 3821
rect 2494 3816 2500 3817
rect 2458 3807 2464 3808
rect 2458 3803 2459 3807
rect 2463 3803 2464 3807
rect 2458 3802 2464 3803
rect 2496 3779 2498 3816
rect 2580 3800 2582 3826
rect 2630 3821 2636 3822
rect 2630 3817 2631 3821
rect 2635 3817 2636 3821
rect 2630 3816 2636 3817
rect 2578 3799 2584 3800
rect 2578 3795 2579 3799
rect 2583 3795 2584 3799
rect 2578 3794 2584 3795
rect 2632 3779 2634 3816
rect 2716 3800 2718 3826
rect 2774 3821 2780 3822
rect 2774 3817 2775 3821
rect 2779 3817 2780 3821
rect 2774 3816 2780 3817
rect 2714 3799 2720 3800
rect 2714 3795 2715 3799
rect 2719 3795 2720 3799
rect 2714 3794 2720 3795
rect 2776 3779 2778 3816
rect 2876 3800 2878 3902
rect 2982 3900 2988 3901
rect 2982 3896 2983 3900
rect 2987 3896 2988 3900
rect 2982 3895 2988 3896
rect 2984 3871 2986 3895
rect 2919 3870 2923 3871
rect 2919 3865 2923 3866
rect 2983 3870 2987 3871
rect 2983 3865 2987 3866
rect 2920 3841 2922 3865
rect 2918 3840 2924 3841
rect 2918 3836 2919 3840
rect 2923 3836 2924 3840
rect 2918 3835 2924 3836
rect 3052 3832 3054 3934
rect 3176 3920 3178 3941
rect 3244 3940 3246 3978
rect 3342 3973 3348 3974
rect 3342 3969 3343 3973
rect 3347 3969 3348 3973
rect 3342 3968 3348 3969
rect 3942 3972 3948 3973
rect 3942 3968 3943 3972
rect 3947 3968 3948 3972
rect 3344 3947 3346 3968
rect 3942 3967 3948 3968
rect 3944 3947 3946 3967
rect 3343 3946 3347 3947
rect 3343 3941 3347 3942
rect 3367 3946 3371 3947
rect 3367 3941 3371 3942
rect 3559 3946 3563 3947
rect 3559 3941 3563 3942
rect 3943 3946 3947 3947
rect 3943 3941 3947 3942
rect 3242 3939 3248 3940
rect 3242 3935 3243 3939
rect 3247 3935 3248 3939
rect 3242 3934 3248 3935
rect 3250 3939 3256 3940
rect 3250 3935 3251 3939
rect 3255 3935 3256 3939
rect 3250 3934 3256 3935
rect 3174 3919 3180 3920
rect 3174 3915 3175 3919
rect 3179 3915 3180 3919
rect 3174 3914 3180 3915
rect 3252 3912 3254 3934
rect 3368 3920 3370 3941
rect 3442 3939 3448 3940
rect 3442 3935 3443 3939
rect 3447 3935 3448 3939
rect 3442 3934 3448 3935
rect 3366 3919 3372 3920
rect 3366 3915 3367 3919
rect 3371 3915 3372 3919
rect 3366 3914 3372 3915
rect 3444 3912 3446 3934
rect 3560 3920 3562 3941
rect 3944 3921 3946 3941
rect 3942 3920 3948 3921
rect 3558 3919 3564 3920
rect 3558 3915 3559 3919
rect 3563 3915 3564 3919
rect 3942 3916 3943 3920
rect 3947 3916 3948 3920
rect 3942 3915 3948 3916
rect 3558 3914 3564 3915
rect 3250 3911 3256 3912
rect 3250 3907 3251 3911
rect 3255 3907 3256 3911
rect 3250 3906 3256 3907
rect 3442 3911 3448 3912
rect 3442 3907 3443 3911
rect 3447 3907 3448 3911
rect 3442 3906 3448 3907
rect 3538 3911 3544 3912
rect 3538 3907 3539 3911
rect 3543 3907 3544 3911
rect 3538 3906 3544 3907
rect 3174 3900 3180 3901
rect 3174 3896 3175 3900
rect 3179 3896 3180 3900
rect 3174 3895 3180 3896
rect 3366 3900 3372 3901
rect 3366 3896 3367 3900
rect 3371 3896 3372 3900
rect 3366 3895 3372 3896
rect 3176 3871 3178 3895
rect 3368 3871 3370 3895
rect 3063 3870 3067 3871
rect 3063 3865 3067 3866
rect 3175 3870 3179 3871
rect 3175 3865 3179 3866
rect 3207 3870 3211 3871
rect 3207 3865 3211 3866
rect 3343 3870 3347 3871
rect 3343 3865 3347 3866
rect 3367 3870 3371 3871
rect 3367 3865 3371 3866
rect 3471 3870 3475 3871
rect 3471 3865 3475 3866
rect 3064 3841 3066 3865
rect 3208 3841 3210 3865
rect 3344 3841 3346 3865
rect 3472 3841 3474 3865
rect 3062 3840 3068 3841
rect 3062 3836 3063 3840
rect 3067 3836 3068 3840
rect 3062 3835 3068 3836
rect 3206 3840 3212 3841
rect 3206 3836 3207 3840
rect 3211 3836 3212 3840
rect 3206 3835 3212 3836
rect 3342 3840 3348 3841
rect 3342 3836 3343 3840
rect 3347 3836 3348 3840
rect 3342 3835 3348 3836
rect 3470 3840 3476 3841
rect 3470 3836 3471 3840
rect 3475 3836 3476 3840
rect 3470 3835 3476 3836
rect 2994 3831 3000 3832
rect 2994 3827 2995 3831
rect 2999 3827 3000 3831
rect 2994 3826 3000 3827
rect 3050 3831 3056 3832
rect 3050 3827 3051 3831
rect 3055 3827 3056 3831
rect 3050 3826 3056 3827
rect 3274 3831 3280 3832
rect 3274 3827 3275 3831
rect 3279 3827 3280 3831
rect 3274 3826 3280 3827
rect 3290 3831 3296 3832
rect 3290 3827 3291 3831
rect 3295 3827 3296 3831
rect 3290 3826 3296 3827
rect 3426 3831 3432 3832
rect 3426 3827 3427 3831
rect 3431 3827 3432 3831
rect 3426 3826 3432 3827
rect 2918 3821 2924 3822
rect 2918 3817 2919 3821
rect 2923 3817 2924 3821
rect 2918 3816 2924 3817
rect 2874 3799 2880 3800
rect 2874 3795 2875 3799
rect 2879 3795 2880 3799
rect 2874 3794 2880 3795
rect 2882 3799 2888 3800
rect 2882 3795 2883 3799
rect 2887 3795 2888 3799
rect 2882 3794 2888 3795
rect 2479 3778 2483 3779
rect 2479 3773 2483 3774
rect 2495 3778 2499 3779
rect 2495 3773 2499 3774
rect 2631 3778 2635 3779
rect 2631 3773 2635 3774
rect 2639 3778 2643 3779
rect 2639 3773 2643 3774
rect 2775 3778 2779 3779
rect 2775 3773 2779 3774
rect 2807 3778 2811 3779
rect 2807 3773 2811 3774
rect 2450 3771 2456 3772
rect 2450 3767 2451 3771
rect 2455 3767 2456 3771
rect 2450 3766 2456 3767
rect 2480 3752 2482 3773
rect 2554 3771 2560 3772
rect 2554 3767 2555 3771
rect 2559 3767 2560 3771
rect 2554 3766 2560 3767
rect 2182 3751 2188 3752
rect 2182 3747 2183 3751
rect 2187 3747 2188 3751
rect 2182 3746 2188 3747
rect 2326 3751 2332 3752
rect 2326 3747 2327 3751
rect 2331 3747 2332 3751
rect 2326 3746 2332 3747
rect 2478 3751 2484 3752
rect 2478 3747 2479 3751
rect 2483 3747 2484 3751
rect 2478 3746 2484 3747
rect 2556 3744 2558 3766
rect 2598 3763 2604 3764
rect 2598 3759 2599 3763
rect 2603 3759 2604 3763
rect 2598 3758 2604 3759
rect 2600 3744 2602 3758
rect 2640 3752 2642 3773
rect 2808 3752 2810 3773
rect 2638 3751 2644 3752
rect 2638 3747 2639 3751
rect 2643 3747 2644 3751
rect 2638 3746 2644 3747
rect 2806 3751 2812 3752
rect 2806 3747 2807 3751
rect 2811 3747 2812 3751
rect 2806 3746 2812 3747
rect 2884 3744 2886 3794
rect 2920 3779 2922 3816
rect 2996 3800 2998 3826
rect 3062 3821 3068 3822
rect 3062 3817 3063 3821
rect 3067 3817 3068 3821
rect 3062 3816 3068 3817
rect 3206 3821 3212 3822
rect 3206 3817 3207 3821
rect 3211 3817 3212 3821
rect 3206 3816 3212 3817
rect 2994 3799 3000 3800
rect 2994 3795 2995 3799
rect 2999 3795 3000 3799
rect 2994 3794 3000 3795
rect 3064 3779 3066 3816
rect 3208 3779 3210 3816
rect 2919 3778 2923 3779
rect 2919 3773 2923 3774
rect 2983 3778 2987 3779
rect 2983 3773 2987 3774
rect 3063 3778 3067 3779
rect 3063 3773 3067 3774
rect 3159 3778 3163 3779
rect 3159 3773 3163 3774
rect 3207 3778 3211 3779
rect 3207 3773 3211 3774
rect 2890 3771 2896 3772
rect 2890 3767 2891 3771
rect 2895 3767 2896 3771
rect 2890 3766 2896 3767
rect 2892 3744 2894 3766
rect 2984 3752 2986 3773
rect 3002 3771 3008 3772
rect 3002 3767 3003 3771
rect 3007 3767 3008 3771
rect 3002 3766 3008 3767
rect 2982 3751 2988 3752
rect 2982 3747 2983 3751
rect 2987 3747 2988 3751
rect 2982 3746 2988 3747
rect 2154 3743 2160 3744
rect 2006 3740 2012 3741
rect 1606 3739 1612 3740
rect 1606 3735 1607 3739
rect 1611 3735 1612 3739
rect 2006 3736 2007 3740
rect 2011 3736 2012 3740
rect 2154 3739 2155 3743
rect 2159 3739 2160 3743
rect 2154 3738 2160 3739
rect 2554 3743 2560 3744
rect 2554 3739 2555 3743
rect 2559 3739 2560 3743
rect 2554 3738 2560 3739
rect 2598 3743 2604 3744
rect 2598 3739 2599 3743
rect 2603 3739 2604 3743
rect 2598 3738 2604 3739
rect 2882 3743 2888 3744
rect 2882 3739 2883 3743
rect 2887 3739 2888 3743
rect 2882 3738 2888 3739
rect 2890 3743 2896 3744
rect 2890 3739 2891 3743
rect 2895 3739 2896 3743
rect 2890 3738 2896 3739
rect 2006 3735 2012 3736
rect 2046 3735 2052 3736
rect 1606 3734 1612 3735
rect 2046 3731 2047 3735
rect 2051 3731 2052 3735
rect 2138 3735 2144 3736
rect 2046 3730 2052 3731
rect 2070 3732 2076 3733
rect 2006 3723 2012 3724
rect 1606 3720 1612 3721
rect 1606 3716 1607 3720
rect 1611 3716 1612 3720
rect 2006 3719 2007 3723
rect 2011 3719 2012 3723
rect 2006 3718 2012 3719
rect 1606 3715 1612 3716
rect 1608 3683 1610 3715
rect 2008 3683 2010 3718
rect 2048 3691 2050 3730
rect 2070 3728 2071 3732
rect 2075 3728 2076 3732
rect 2138 3731 2139 3735
rect 2143 3731 2144 3735
rect 2138 3730 2144 3731
rect 2182 3732 2188 3733
rect 2070 3727 2076 3728
rect 2072 3691 2074 3727
rect 2047 3690 2051 3691
rect 2047 3685 2051 3686
rect 2071 3690 2075 3691
rect 2071 3685 2075 3686
rect 1607 3682 1611 3683
rect 1607 3677 1611 3678
rect 1695 3682 1699 3683
rect 1695 3677 1699 3678
rect 2007 3682 2011 3683
rect 2007 3677 2011 3678
rect 1696 3653 1698 3677
rect 1694 3652 1700 3653
rect 1694 3648 1695 3652
rect 1699 3648 1700 3652
rect 2008 3650 2010 3677
rect 2048 3658 2050 3685
rect 2072 3661 2074 3685
rect 2070 3660 2076 3661
rect 2046 3657 2052 3658
rect 2046 3653 2047 3657
rect 2051 3653 2052 3657
rect 2070 3656 2071 3660
rect 2075 3656 2076 3660
rect 2070 3655 2076 3656
rect 2046 3652 2052 3653
rect 1694 3647 1700 3648
rect 2006 3649 2012 3650
rect 2006 3645 2007 3649
rect 2011 3645 2012 3649
rect 2006 3644 2012 3645
rect 1554 3643 1560 3644
rect 1554 3639 1555 3643
rect 1559 3639 1560 3643
rect 1554 3638 1560 3639
rect 1562 3643 1568 3644
rect 1562 3639 1563 3643
rect 1567 3639 1568 3643
rect 2070 3641 2076 3642
rect 1562 3638 1568 3639
rect 2046 3640 2052 3641
rect 1478 3633 1484 3634
rect 1478 3629 1479 3633
rect 1483 3629 1484 3633
rect 1478 3628 1484 3629
rect 1346 3619 1352 3620
rect 1346 3615 1347 3619
rect 1351 3615 1352 3619
rect 1346 3614 1352 3615
rect 1480 3603 1482 3628
rect 1564 3612 1566 3638
rect 2046 3636 2047 3640
rect 2051 3636 2052 3640
rect 2070 3637 2071 3641
rect 2075 3637 2076 3641
rect 2070 3636 2076 3637
rect 2046 3635 2052 3636
rect 1694 3633 1700 3634
rect 1694 3629 1695 3633
rect 1699 3629 1700 3633
rect 1694 3628 1700 3629
rect 2006 3632 2012 3633
rect 2006 3628 2007 3632
rect 2011 3628 2012 3632
rect 1562 3611 1568 3612
rect 1562 3607 1563 3611
rect 1567 3607 1568 3611
rect 1562 3606 1568 3607
rect 1696 3603 1698 3628
rect 2006 3627 2012 3628
rect 1762 3611 1768 3612
rect 1762 3607 1763 3611
rect 1767 3607 1768 3611
rect 1762 3606 1768 3607
rect 1447 3602 1451 3603
rect 1447 3597 1451 3598
rect 1479 3602 1483 3603
rect 1479 3597 1483 3598
rect 1687 3602 1691 3603
rect 1687 3597 1691 3598
rect 1695 3602 1699 3603
rect 1695 3597 1699 3598
rect 1298 3595 1304 3596
rect 1298 3591 1299 3595
rect 1303 3591 1304 3595
rect 1298 3590 1304 3591
rect 1338 3595 1344 3596
rect 1338 3591 1339 3595
rect 1343 3591 1344 3595
rect 1338 3590 1344 3591
rect 774 3575 780 3576
rect 774 3571 775 3575
rect 779 3571 780 3575
rect 774 3570 780 3571
rect 990 3575 996 3576
rect 990 3571 991 3575
rect 995 3571 996 3575
rect 990 3570 996 3571
rect 1214 3575 1220 3576
rect 1214 3571 1215 3575
rect 1219 3571 1220 3575
rect 1214 3570 1220 3571
rect 1300 3568 1302 3590
rect 1448 3576 1450 3597
rect 1688 3576 1690 3597
rect 1754 3595 1760 3596
rect 1754 3591 1755 3595
rect 1759 3591 1760 3595
rect 1754 3590 1760 3591
rect 1446 3575 1452 3576
rect 1446 3571 1447 3575
rect 1451 3571 1452 3575
rect 1446 3570 1452 3571
rect 1686 3575 1692 3576
rect 1686 3571 1687 3575
rect 1691 3571 1692 3575
rect 1686 3570 1692 3571
rect 242 3567 248 3568
rect 242 3563 243 3567
rect 247 3563 248 3567
rect 242 3562 248 3563
rect 434 3567 440 3568
rect 434 3563 435 3567
rect 439 3563 440 3567
rect 434 3562 440 3563
rect 634 3567 640 3568
rect 634 3563 635 3567
rect 639 3563 640 3567
rect 634 3562 640 3563
rect 682 3567 688 3568
rect 682 3563 683 3567
rect 687 3563 688 3567
rect 1298 3567 1304 3568
rect 682 3562 688 3563
rect 1066 3563 1072 3564
rect 110 3559 116 3560
rect 110 3555 111 3559
rect 115 3555 116 3559
rect 1066 3559 1067 3563
rect 1071 3559 1072 3563
rect 1298 3563 1299 3567
rect 1303 3563 1304 3567
rect 1298 3562 1304 3563
rect 1066 3558 1072 3559
rect 110 3554 116 3555
rect 166 3556 172 3557
rect 112 3519 114 3554
rect 166 3552 167 3556
rect 171 3552 172 3556
rect 166 3551 172 3552
rect 358 3556 364 3557
rect 358 3552 359 3556
rect 363 3552 364 3556
rect 358 3551 364 3552
rect 558 3556 564 3557
rect 558 3552 559 3556
rect 563 3552 564 3556
rect 558 3551 564 3552
rect 774 3556 780 3557
rect 774 3552 775 3556
rect 779 3552 780 3556
rect 774 3551 780 3552
rect 990 3556 996 3557
rect 990 3552 991 3556
rect 995 3552 996 3556
rect 990 3551 996 3552
rect 168 3519 170 3551
rect 360 3519 362 3551
rect 560 3519 562 3551
rect 776 3519 778 3551
rect 992 3519 994 3551
rect 111 3518 115 3519
rect 111 3513 115 3514
rect 167 3518 171 3519
rect 167 3513 171 3514
rect 295 3518 299 3519
rect 295 3513 299 3514
rect 359 3518 363 3519
rect 359 3513 363 3514
rect 431 3518 435 3519
rect 431 3513 435 3514
rect 559 3518 563 3519
rect 559 3513 563 3514
rect 583 3518 587 3519
rect 583 3513 587 3514
rect 743 3518 747 3519
rect 743 3513 747 3514
rect 775 3518 779 3519
rect 775 3513 779 3514
rect 911 3518 915 3519
rect 911 3513 915 3514
rect 991 3518 995 3519
rect 991 3513 995 3514
rect 112 3486 114 3513
rect 296 3489 298 3513
rect 432 3489 434 3513
rect 584 3489 586 3513
rect 744 3489 746 3513
rect 912 3489 914 3513
rect 294 3488 300 3489
rect 110 3485 116 3486
rect 110 3481 111 3485
rect 115 3481 116 3485
rect 294 3484 295 3488
rect 299 3484 300 3488
rect 294 3483 300 3484
rect 430 3488 436 3489
rect 430 3484 431 3488
rect 435 3484 436 3488
rect 430 3483 436 3484
rect 582 3488 588 3489
rect 582 3484 583 3488
rect 587 3484 588 3488
rect 582 3483 588 3484
rect 742 3488 748 3489
rect 742 3484 743 3488
rect 747 3484 748 3488
rect 742 3483 748 3484
rect 910 3488 916 3489
rect 910 3484 911 3488
rect 915 3484 916 3488
rect 910 3483 916 3484
rect 110 3480 116 3481
rect 378 3479 384 3480
rect 378 3475 379 3479
rect 383 3475 384 3479
rect 378 3474 384 3475
rect 514 3479 520 3480
rect 514 3475 515 3479
rect 519 3475 520 3479
rect 514 3474 520 3475
rect 666 3479 672 3480
rect 666 3475 667 3479
rect 671 3475 672 3479
rect 666 3474 672 3475
rect 826 3479 832 3480
rect 826 3475 827 3479
rect 831 3475 832 3479
rect 826 3474 832 3475
rect 294 3469 300 3470
rect 110 3468 116 3469
rect 110 3464 111 3468
rect 115 3464 116 3468
rect 294 3465 295 3469
rect 299 3465 300 3469
rect 294 3464 300 3465
rect 110 3463 116 3464
rect 112 3423 114 3463
rect 296 3423 298 3464
rect 380 3448 382 3474
rect 430 3469 436 3470
rect 430 3465 431 3469
rect 435 3465 436 3469
rect 430 3464 436 3465
rect 378 3447 384 3448
rect 378 3443 379 3447
rect 383 3443 384 3447
rect 378 3442 384 3443
rect 432 3423 434 3464
rect 516 3448 518 3474
rect 582 3469 588 3470
rect 582 3465 583 3469
rect 587 3465 588 3469
rect 582 3464 588 3465
rect 514 3447 520 3448
rect 514 3443 515 3447
rect 519 3443 520 3447
rect 514 3442 520 3443
rect 584 3423 586 3464
rect 668 3448 670 3474
rect 742 3469 748 3470
rect 742 3465 743 3469
rect 747 3465 748 3469
rect 742 3464 748 3465
rect 666 3447 672 3448
rect 666 3443 667 3447
rect 671 3443 672 3447
rect 666 3442 672 3443
rect 744 3423 746 3464
rect 828 3448 830 3474
rect 910 3469 916 3470
rect 910 3465 911 3469
rect 915 3465 916 3469
rect 910 3464 916 3465
rect 826 3447 832 3448
rect 826 3443 827 3447
rect 831 3443 832 3447
rect 826 3442 832 3443
rect 912 3423 914 3464
rect 1068 3448 1070 3558
rect 1214 3556 1220 3557
rect 1214 3552 1215 3556
rect 1219 3552 1220 3556
rect 1214 3551 1220 3552
rect 1446 3556 1452 3557
rect 1446 3552 1447 3556
rect 1451 3552 1452 3556
rect 1446 3551 1452 3552
rect 1686 3556 1692 3557
rect 1686 3552 1687 3556
rect 1691 3552 1692 3556
rect 1686 3551 1692 3552
rect 1216 3519 1218 3551
rect 1448 3519 1450 3551
rect 1688 3519 1690 3551
rect 1079 3518 1083 3519
rect 1079 3513 1083 3514
rect 1215 3518 1219 3519
rect 1215 3513 1219 3514
rect 1247 3518 1251 3519
rect 1247 3513 1251 3514
rect 1423 3518 1427 3519
rect 1423 3513 1427 3514
rect 1447 3518 1451 3519
rect 1447 3513 1451 3514
rect 1599 3518 1603 3519
rect 1599 3513 1603 3514
rect 1687 3518 1691 3519
rect 1687 3513 1691 3514
rect 1080 3489 1082 3513
rect 1248 3489 1250 3513
rect 1424 3489 1426 3513
rect 1600 3489 1602 3513
rect 1078 3488 1084 3489
rect 1078 3484 1079 3488
rect 1083 3484 1084 3488
rect 1078 3483 1084 3484
rect 1246 3488 1252 3489
rect 1246 3484 1247 3488
rect 1251 3484 1252 3488
rect 1246 3483 1252 3484
rect 1422 3488 1428 3489
rect 1422 3484 1423 3488
rect 1427 3484 1428 3488
rect 1422 3483 1428 3484
rect 1598 3488 1604 3489
rect 1598 3484 1599 3488
rect 1603 3484 1604 3488
rect 1598 3483 1604 3484
rect 1756 3480 1758 3590
rect 1764 3568 1766 3606
rect 2008 3603 2010 3627
rect 2048 3611 2050 3635
rect 2072 3611 2074 3636
rect 2140 3620 2142 3730
rect 2182 3728 2183 3732
rect 2187 3728 2188 3732
rect 2182 3727 2188 3728
rect 2326 3732 2332 3733
rect 2326 3728 2327 3732
rect 2331 3728 2332 3732
rect 2326 3727 2332 3728
rect 2478 3732 2484 3733
rect 2478 3728 2479 3732
rect 2483 3728 2484 3732
rect 2478 3727 2484 3728
rect 2638 3732 2644 3733
rect 2638 3728 2639 3732
rect 2643 3728 2644 3732
rect 2638 3727 2644 3728
rect 2806 3732 2812 3733
rect 2806 3728 2807 3732
rect 2811 3728 2812 3732
rect 2806 3727 2812 3728
rect 2982 3732 2988 3733
rect 2982 3728 2983 3732
rect 2987 3728 2988 3732
rect 2982 3727 2988 3728
rect 2184 3691 2186 3727
rect 2328 3691 2330 3727
rect 2480 3691 2482 3727
rect 2640 3691 2642 3727
rect 2808 3691 2810 3727
rect 2984 3691 2986 3727
rect 2183 3690 2187 3691
rect 2183 3685 2187 3686
rect 2199 3690 2203 3691
rect 2199 3685 2203 3686
rect 2327 3690 2331 3691
rect 2327 3685 2331 3686
rect 2367 3690 2371 3691
rect 2367 3685 2371 3686
rect 2479 3690 2483 3691
rect 2479 3685 2483 3686
rect 2551 3690 2555 3691
rect 2551 3685 2555 3686
rect 2639 3690 2643 3691
rect 2639 3685 2643 3686
rect 2735 3690 2739 3691
rect 2735 3685 2739 3686
rect 2807 3690 2811 3691
rect 2807 3685 2811 3686
rect 2927 3690 2931 3691
rect 2927 3685 2931 3686
rect 2983 3690 2987 3691
rect 2983 3685 2987 3686
rect 2200 3661 2202 3685
rect 2368 3661 2370 3685
rect 2552 3661 2554 3685
rect 2736 3661 2738 3685
rect 2928 3661 2930 3685
rect 2198 3660 2204 3661
rect 2198 3656 2199 3660
rect 2203 3656 2204 3660
rect 2198 3655 2204 3656
rect 2366 3660 2372 3661
rect 2366 3656 2367 3660
rect 2371 3656 2372 3660
rect 2366 3655 2372 3656
rect 2550 3660 2556 3661
rect 2550 3656 2551 3660
rect 2555 3656 2556 3660
rect 2550 3655 2556 3656
rect 2734 3660 2740 3661
rect 2734 3656 2735 3660
rect 2739 3656 2740 3660
rect 2734 3655 2740 3656
rect 2926 3660 2932 3661
rect 2926 3656 2927 3660
rect 2931 3656 2932 3660
rect 2926 3655 2932 3656
rect 3004 3652 3006 3766
rect 3160 3752 3162 3773
rect 3276 3772 3278 3826
rect 3292 3800 3294 3826
rect 3342 3821 3348 3822
rect 3342 3817 3343 3821
rect 3347 3817 3348 3821
rect 3342 3816 3348 3817
rect 3290 3799 3296 3800
rect 3290 3795 3291 3799
rect 3295 3795 3296 3799
rect 3290 3794 3296 3795
rect 3344 3779 3346 3816
rect 3428 3800 3430 3826
rect 3470 3821 3476 3822
rect 3470 3817 3471 3821
rect 3475 3817 3476 3821
rect 3470 3816 3476 3817
rect 3426 3799 3432 3800
rect 3426 3795 3427 3799
rect 3431 3795 3432 3799
rect 3426 3794 3432 3795
rect 3472 3779 3474 3816
rect 3540 3800 3542 3906
rect 3942 3903 3948 3904
rect 3558 3900 3564 3901
rect 3558 3896 3559 3900
rect 3563 3896 3564 3900
rect 3942 3899 3943 3903
rect 3947 3899 3948 3903
rect 3942 3898 3948 3899
rect 3558 3895 3564 3896
rect 3560 3871 3562 3895
rect 3944 3871 3946 3898
rect 3559 3870 3563 3871
rect 3559 3865 3563 3866
rect 3599 3870 3603 3871
rect 3599 3865 3603 3866
rect 3727 3870 3731 3871
rect 3727 3865 3731 3866
rect 3839 3870 3843 3871
rect 3839 3865 3843 3866
rect 3943 3870 3947 3871
rect 3943 3865 3947 3866
rect 3600 3841 3602 3865
rect 3728 3841 3730 3865
rect 3840 3841 3842 3865
rect 3598 3840 3604 3841
rect 3598 3836 3599 3840
rect 3603 3836 3604 3840
rect 3598 3835 3604 3836
rect 3726 3840 3732 3841
rect 3726 3836 3727 3840
rect 3731 3836 3732 3840
rect 3726 3835 3732 3836
rect 3838 3840 3844 3841
rect 3838 3836 3839 3840
rect 3843 3836 3844 3840
rect 3944 3838 3946 3865
rect 3838 3835 3844 3836
rect 3942 3837 3948 3838
rect 3942 3833 3943 3837
rect 3947 3833 3948 3837
rect 3942 3832 3948 3833
rect 3674 3831 3680 3832
rect 3674 3827 3675 3831
rect 3679 3827 3680 3831
rect 3674 3826 3680 3827
rect 3802 3831 3808 3832
rect 3802 3827 3803 3831
rect 3807 3827 3808 3831
rect 3802 3826 3808 3827
rect 3906 3831 3912 3832
rect 3906 3827 3907 3831
rect 3911 3827 3912 3831
rect 3906 3826 3912 3827
rect 3598 3821 3604 3822
rect 3598 3817 3599 3821
rect 3603 3817 3604 3821
rect 3598 3816 3604 3817
rect 3538 3799 3544 3800
rect 3538 3795 3539 3799
rect 3543 3795 3544 3799
rect 3538 3794 3544 3795
rect 3600 3779 3602 3816
rect 3676 3808 3678 3826
rect 3726 3821 3732 3822
rect 3726 3817 3727 3821
rect 3731 3817 3732 3821
rect 3726 3816 3732 3817
rect 3674 3807 3680 3808
rect 3674 3803 3675 3807
rect 3679 3803 3680 3807
rect 3674 3802 3680 3803
rect 3728 3779 3730 3816
rect 3804 3800 3806 3826
rect 3838 3821 3844 3822
rect 3838 3817 3839 3821
rect 3843 3817 3844 3821
rect 3838 3816 3844 3817
rect 3802 3799 3808 3800
rect 3802 3795 3803 3799
rect 3807 3795 3808 3799
rect 3802 3794 3808 3795
rect 3840 3779 3842 3816
rect 3335 3778 3339 3779
rect 3335 3773 3339 3774
rect 3343 3778 3347 3779
rect 3343 3773 3347 3774
rect 3471 3778 3475 3779
rect 3471 3773 3475 3774
rect 3511 3778 3515 3779
rect 3511 3773 3515 3774
rect 3599 3778 3603 3779
rect 3599 3773 3603 3774
rect 3687 3778 3691 3779
rect 3687 3773 3691 3774
rect 3727 3778 3731 3779
rect 3727 3773 3731 3774
rect 3839 3778 3843 3779
rect 3839 3773 3843 3774
rect 3274 3771 3280 3772
rect 3274 3767 3275 3771
rect 3279 3767 3280 3771
rect 3274 3766 3280 3767
rect 3298 3771 3304 3772
rect 3298 3767 3299 3771
rect 3303 3767 3304 3771
rect 3298 3766 3304 3767
rect 3158 3751 3164 3752
rect 3158 3747 3159 3751
rect 3163 3747 3164 3751
rect 3158 3746 3164 3747
rect 3300 3744 3302 3766
rect 3336 3752 3338 3773
rect 3410 3771 3416 3772
rect 3410 3767 3411 3771
rect 3415 3767 3416 3771
rect 3410 3766 3416 3767
rect 3334 3751 3340 3752
rect 3334 3747 3335 3751
rect 3339 3747 3340 3751
rect 3334 3746 3340 3747
rect 3412 3744 3414 3766
rect 3512 3752 3514 3773
rect 3688 3752 3690 3773
rect 3746 3771 3752 3772
rect 3746 3767 3747 3771
rect 3751 3767 3752 3771
rect 3746 3766 3752 3767
rect 3510 3751 3516 3752
rect 3510 3747 3511 3751
rect 3515 3747 3516 3751
rect 3510 3746 3516 3747
rect 3686 3751 3692 3752
rect 3686 3747 3687 3751
rect 3691 3747 3692 3751
rect 3686 3746 3692 3747
rect 3298 3743 3304 3744
rect 3298 3739 3299 3743
rect 3303 3739 3304 3743
rect 3298 3738 3304 3739
rect 3410 3743 3416 3744
rect 3410 3739 3411 3743
rect 3415 3739 3416 3743
rect 3410 3738 3416 3739
rect 3586 3739 3592 3740
rect 3586 3735 3587 3739
rect 3591 3735 3592 3739
rect 3586 3734 3592 3735
rect 3158 3732 3164 3733
rect 3158 3728 3159 3732
rect 3163 3728 3164 3732
rect 3158 3727 3164 3728
rect 3334 3732 3340 3733
rect 3334 3728 3335 3732
rect 3339 3728 3340 3732
rect 3334 3727 3340 3728
rect 3510 3732 3516 3733
rect 3510 3728 3511 3732
rect 3515 3728 3516 3732
rect 3510 3727 3516 3728
rect 3160 3691 3162 3727
rect 3336 3691 3338 3727
rect 3512 3691 3514 3727
rect 3111 3690 3115 3691
rect 3111 3685 3115 3686
rect 3159 3690 3163 3691
rect 3159 3685 3163 3686
rect 3295 3690 3299 3691
rect 3295 3685 3299 3686
rect 3335 3690 3339 3691
rect 3335 3685 3339 3686
rect 3479 3690 3483 3691
rect 3479 3685 3483 3686
rect 3511 3690 3515 3691
rect 3511 3685 3515 3686
rect 3112 3661 3114 3685
rect 3296 3661 3298 3685
rect 3480 3661 3482 3685
rect 3110 3660 3116 3661
rect 3110 3656 3111 3660
rect 3115 3656 3116 3660
rect 3110 3655 3116 3656
rect 3294 3660 3300 3661
rect 3294 3656 3295 3660
rect 3299 3656 3300 3660
rect 3294 3655 3300 3656
rect 3478 3660 3484 3661
rect 3478 3656 3479 3660
rect 3483 3656 3484 3660
rect 3478 3655 3484 3656
rect 2146 3651 2152 3652
rect 2146 3647 2147 3651
rect 2151 3647 2152 3651
rect 2146 3646 2152 3647
rect 2274 3651 2280 3652
rect 2274 3647 2275 3651
rect 2279 3647 2280 3651
rect 2274 3646 2280 3647
rect 2442 3651 2448 3652
rect 2442 3647 2443 3651
rect 2447 3647 2448 3651
rect 2442 3646 2448 3647
rect 2626 3651 2632 3652
rect 2626 3647 2627 3651
rect 2631 3647 2632 3651
rect 2626 3646 2632 3647
rect 3002 3651 3008 3652
rect 3002 3647 3003 3651
rect 3007 3647 3008 3651
rect 3002 3646 3008 3647
rect 3186 3651 3192 3652
rect 3186 3647 3187 3651
rect 3191 3647 3192 3651
rect 3186 3646 3192 3647
rect 3194 3651 3200 3652
rect 3194 3647 3195 3651
rect 3199 3647 3200 3651
rect 3194 3646 3200 3647
rect 3378 3651 3384 3652
rect 3378 3647 3379 3651
rect 3383 3647 3384 3651
rect 3378 3646 3384 3647
rect 2148 3620 2150 3646
rect 2198 3641 2204 3642
rect 2198 3637 2199 3641
rect 2203 3637 2204 3641
rect 2198 3636 2204 3637
rect 2170 3635 2176 3636
rect 2170 3631 2171 3635
rect 2175 3631 2176 3635
rect 2170 3630 2176 3631
rect 2138 3619 2144 3620
rect 2138 3615 2139 3619
rect 2143 3615 2144 3619
rect 2138 3614 2144 3615
rect 2146 3619 2152 3620
rect 2146 3615 2147 3619
rect 2151 3615 2152 3619
rect 2146 3614 2152 3615
rect 2047 3610 2051 3611
rect 2047 3605 2051 3606
rect 2071 3610 2075 3611
rect 2071 3605 2075 3606
rect 2103 3610 2107 3611
rect 2103 3605 2107 3606
rect 2007 3602 2011 3603
rect 2007 3597 2011 3598
rect 2008 3577 2010 3597
rect 2048 3585 2050 3605
rect 2046 3584 2052 3585
rect 2104 3584 2106 3605
rect 2172 3604 2174 3630
rect 2200 3611 2202 3636
rect 2276 3620 2278 3646
rect 2366 3641 2372 3642
rect 2366 3637 2367 3641
rect 2371 3637 2372 3641
rect 2366 3636 2372 3637
rect 2274 3619 2280 3620
rect 2274 3615 2275 3619
rect 2279 3615 2280 3619
rect 2274 3614 2280 3615
rect 2368 3611 2370 3636
rect 2444 3620 2446 3646
rect 2550 3641 2556 3642
rect 2550 3637 2551 3641
rect 2555 3637 2556 3641
rect 2550 3636 2556 3637
rect 2442 3619 2448 3620
rect 2442 3615 2443 3619
rect 2447 3615 2448 3619
rect 2442 3614 2448 3615
rect 2552 3611 2554 3636
rect 2628 3620 2630 3646
rect 2734 3641 2740 3642
rect 2734 3637 2735 3641
rect 2739 3637 2740 3641
rect 2734 3636 2740 3637
rect 2926 3641 2932 3642
rect 2926 3637 2927 3641
rect 2931 3637 2932 3641
rect 2926 3636 2932 3637
rect 3110 3641 3116 3642
rect 3110 3637 3111 3641
rect 3115 3637 3116 3641
rect 3110 3636 3116 3637
rect 2626 3619 2632 3620
rect 2626 3615 2627 3619
rect 2631 3615 2632 3619
rect 2626 3614 2632 3615
rect 2736 3611 2738 3636
rect 2928 3611 2930 3636
rect 3112 3611 3114 3636
rect 2199 3610 2203 3611
rect 2199 3605 2203 3606
rect 2279 3610 2283 3611
rect 2279 3605 2283 3606
rect 2367 3610 2371 3611
rect 2367 3605 2371 3606
rect 2471 3610 2475 3611
rect 2471 3605 2475 3606
rect 2551 3610 2555 3611
rect 2551 3605 2555 3606
rect 2671 3610 2675 3611
rect 2671 3605 2675 3606
rect 2735 3610 2739 3611
rect 2735 3605 2739 3606
rect 2871 3610 2875 3611
rect 2871 3605 2875 3606
rect 2927 3610 2931 3611
rect 2927 3605 2931 3606
rect 3063 3610 3067 3611
rect 3063 3605 3067 3606
rect 3111 3610 3115 3611
rect 3111 3605 3115 3606
rect 2170 3603 2176 3604
rect 2170 3599 2171 3603
rect 2175 3599 2176 3603
rect 2170 3598 2176 3599
rect 2178 3603 2184 3604
rect 2178 3599 2179 3603
rect 2183 3599 2184 3603
rect 2178 3598 2184 3599
rect 2046 3580 2047 3584
rect 2051 3580 2052 3584
rect 2046 3579 2052 3580
rect 2102 3583 2108 3584
rect 2102 3579 2103 3583
rect 2107 3579 2108 3583
rect 2102 3578 2108 3579
rect 2006 3576 2012 3577
rect 2180 3576 2182 3598
rect 2280 3584 2282 3605
rect 2354 3603 2360 3604
rect 2354 3599 2355 3603
rect 2359 3599 2360 3603
rect 2354 3598 2360 3599
rect 2278 3583 2284 3584
rect 2278 3579 2279 3583
rect 2283 3579 2284 3583
rect 2278 3578 2284 3579
rect 2356 3576 2358 3598
rect 2472 3584 2474 3605
rect 2582 3603 2588 3604
rect 2582 3599 2583 3603
rect 2587 3599 2588 3603
rect 2582 3598 2588 3599
rect 2470 3583 2476 3584
rect 2470 3579 2471 3583
rect 2475 3579 2476 3583
rect 2470 3578 2476 3579
rect 2584 3576 2586 3598
rect 2672 3584 2674 3605
rect 2872 3584 2874 3605
rect 2978 3603 2984 3604
rect 2978 3599 2979 3603
rect 2983 3599 2984 3603
rect 2978 3598 2984 3599
rect 2670 3583 2676 3584
rect 2670 3579 2671 3583
rect 2675 3579 2676 3583
rect 2670 3578 2676 3579
rect 2870 3583 2876 3584
rect 2870 3579 2871 3583
rect 2875 3579 2876 3583
rect 2870 3578 2876 3579
rect 2006 3572 2007 3576
rect 2011 3572 2012 3576
rect 2006 3571 2012 3572
rect 2178 3575 2184 3576
rect 2178 3571 2179 3575
rect 2183 3571 2184 3575
rect 2178 3570 2184 3571
rect 2354 3575 2360 3576
rect 2354 3571 2355 3575
rect 2359 3571 2360 3575
rect 2354 3570 2360 3571
rect 2582 3575 2588 3576
rect 2582 3571 2583 3575
rect 2587 3571 2588 3575
rect 2582 3570 2588 3571
rect 2598 3575 2604 3576
rect 2598 3571 2599 3575
rect 2603 3571 2604 3575
rect 2598 3570 2604 3571
rect 1762 3567 1768 3568
rect 1762 3563 1763 3567
rect 1767 3563 1768 3567
rect 1762 3562 1768 3563
rect 2046 3567 2052 3568
rect 2046 3563 2047 3567
rect 2051 3563 2052 3567
rect 2046 3562 2052 3563
rect 2102 3564 2108 3565
rect 2006 3559 2012 3560
rect 2006 3555 2007 3559
rect 2011 3555 2012 3559
rect 2006 3554 2012 3555
rect 2008 3519 2010 3554
rect 2048 3531 2050 3562
rect 2102 3560 2103 3564
rect 2107 3560 2108 3564
rect 2102 3559 2108 3560
rect 2278 3564 2284 3565
rect 2278 3560 2279 3564
rect 2283 3560 2284 3564
rect 2278 3559 2284 3560
rect 2470 3564 2476 3565
rect 2470 3560 2471 3564
rect 2475 3560 2476 3564
rect 2470 3559 2476 3560
rect 2104 3531 2106 3559
rect 2280 3531 2282 3559
rect 2472 3531 2474 3559
rect 2047 3530 2051 3531
rect 2047 3525 2051 3526
rect 2103 3530 2107 3531
rect 2103 3525 2107 3526
rect 2279 3530 2283 3531
rect 2279 3525 2283 3526
rect 2327 3530 2331 3531
rect 2327 3525 2331 3526
rect 2447 3530 2451 3531
rect 2447 3525 2451 3526
rect 2471 3530 2475 3531
rect 2471 3525 2475 3526
rect 2583 3530 2587 3531
rect 2583 3525 2587 3526
rect 1775 3518 1779 3519
rect 1775 3513 1779 3514
rect 2007 3518 2011 3519
rect 2007 3513 2011 3514
rect 1776 3489 1778 3513
rect 1774 3488 1780 3489
rect 1774 3484 1775 3488
rect 1779 3484 1780 3488
rect 2008 3486 2010 3513
rect 2048 3498 2050 3525
rect 2328 3501 2330 3525
rect 2448 3501 2450 3525
rect 2584 3501 2586 3525
rect 2326 3500 2332 3501
rect 2046 3497 2052 3498
rect 2046 3493 2047 3497
rect 2051 3493 2052 3497
rect 2326 3496 2327 3500
rect 2331 3496 2332 3500
rect 2326 3495 2332 3496
rect 2446 3500 2452 3501
rect 2446 3496 2447 3500
rect 2451 3496 2452 3500
rect 2446 3495 2452 3496
rect 2582 3500 2588 3501
rect 2582 3496 2583 3500
rect 2587 3496 2588 3500
rect 2582 3495 2588 3496
rect 2046 3492 2052 3493
rect 2402 3491 2408 3492
rect 2402 3487 2403 3491
rect 2407 3487 2408 3491
rect 2402 3486 2408 3487
rect 2522 3491 2528 3492
rect 2522 3487 2523 3491
rect 2527 3487 2528 3491
rect 2522 3486 2528 3487
rect 1774 3483 1780 3484
rect 2006 3485 2012 3486
rect 2006 3481 2007 3485
rect 2011 3481 2012 3485
rect 2326 3481 2332 3482
rect 2006 3480 2012 3481
rect 2046 3480 2052 3481
rect 1154 3479 1160 3480
rect 1154 3475 1155 3479
rect 1159 3475 1160 3479
rect 1154 3474 1160 3475
rect 1322 3479 1328 3480
rect 1322 3475 1323 3479
rect 1327 3475 1328 3479
rect 1322 3474 1328 3475
rect 1498 3479 1504 3480
rect 1498 3475 1499 3479
rect 1503 3475 1504 3479
rect 1498 3474 1504 3475
rect 1738 3479 1744 3480
rect 1738 3475 1739 3479
rect 1743 3475 1744 3479
rect 1738 3474 1744 3475
rect 1754 3479 1760 3480
rect 1754 3475 1755 3479
rect 1759 3475 1760 3479
rect 2046 3476 2047 3480
rect 2051 3476 2052 3480
rect 2326 3477 2327 3481
rect 2331 3477 2332 3481
rect 2326 3476 2332 3477
rect 2046 3475 2052 3476
rect 1754 3474 1760 3475
rect 1078 3469 1084 3470
rect 1078 3465 1079 3469
rect 1083 3465 1084 3469
rect 1078 3464 1084 3465
rect 1034 3447 1040 3448
rect 1034 3443 1035 3447
rect 1039 3443 1040 3447
rect 1034 3442 1040 3443
rect 1066 3447 1072 3448
rect 1066 3443 1067 3447
rect 1071 3443 1072 3447
rect 1066 3442 1072 3443
rect 111 3422 115 3423
rect 111 3417 115 3418
rect 295 3422 299 3423
rect 295 3417 299 3418
rect 431 3422 435 3423
rect 431 3417 435 3418
rect 495 3422 499 3423
rect 495 3417 499 3418
rect 583 3422 587 3423
rect 583 3417 587 3418
rect 647 3422 651 3423
rect 647 3417 651 3418
rect 743 3422 747 3423
rect 743 3417 747 3418
rect 799 3422 803 3423
rect 799 3417 803 3418
rect 911 3422 915 3423
rect 911 3417 915 3418
rect 959 3422 963 3423
rect 959 3417 963 3418
rect 112 3397 114 3417
rect 110 3396 116 3397
rect 496 3396 498 3417
rect 618 3415 624 3416
rect 618 3411 619 3415
rect 623 3411 624 3415
rect 618 3410 624 3411
rect 626 3415 632 3416
rect 626 3411 627 3415
rect 631 3411 632 3415
rect 626 3410 632 3411
rect 110 3392 111 3396
rect 115 3392 116 3396
rect 110 3391 116 3392
rect 494 3395 500 3396
rect 494 3391 495 3395
rect 499 3391 500 3395
rect 494 3390 500 3391
rect 110 3379 116 3380
rect 110 3375 111 3379
rect 115 3375 116 3379
rect 110 3374 116 3375
rect 494 3376 500 3377
rect 112 3335 114 3374
rect 494 3372 495 3376
rect 499 3372 500 3376
rect 494 3371 500 3372
rect 496 3335 498 3371
rect 111 3334 115 3335
rect 111 3329 115 3330
rect 135 3334 139 3335
rect 135 3329 139 3330
rect 295 3334 299 3335
rect 295 3329 299 3330
rect 479 3334 483 3335
rect 479 3329 483 3330
rect 495 3334 499 3335
rect 495 3329 499 3330
rect 112 3302 114 3329
rect 136 3305 138 3329
rect 296 3305 298 3329
rect 480 3305 482 3329
rect 134 3304 140 3305
rect 110 3301 116 3302
rect 110 3297 111 3301
rect 115 3297 116 3301
rect 134 3300 135 3304
rect 139 3300 140 3304
rect 134 3299 140 3300
rect 294 3304 300 3305
rect 294 3300 295 3304
rect 299 3300 300 3304
rect 294 3299 300 3300
rect 478 3304 484 3305
rect 478 3300 479 3304
rect 483 3300 484 3304
rect 478 3299 484 3300
rect 110 3296 116 3297
rect 620 3296 622 3410
rect 628 3388 630 3410
rect 648 3396 650 3417
rect 722 3415 728 3416
rect 722 3411 723 3415
rect 727 3411 728 3415
rect 722 3410 728 3411
rect 646 3395 652 3396
rect 646 3391 647 3395
rect 651 3391 652 3395
rect 646 3390 652 3391
rect 724 3388 726 3410
rect 800 3396 802 3417
rect 874 3415 880 3416
rect 874 3411 875 3415
rect 879 3411 880 3415
rect 874 3410 880 3411
rect 798 3395 804 3396
rect 798 3391 799 3395
rect 803 3391 804 3395
rect 798 3390 804 3391
rect 876 3388 878 3410
rect 960 3396 962 3417
rect 958 3395 964 3396
rect 958 3391 959 3395
rect 963 3391 964 3395
rect 958 3390 964 3391
rect 1036 3388 1038 3442
rect 1080 3423 1082 3464
rect 1156 3448 1158 3474
rect 1246 3469 1252 3470
rect 1246 3465 1247 3469
rect 1251 3465 1252 3469
rect 1246 3464 1252 3465
rect 1154 3447 1160 3448
rect 1154 3443 1155 3447
rect 1159 3443 1160 3447
rect 1154 3442 1160 3443
rect 1248 3423 1250 3464
rect 1324 3448 1326 3474
rect 1422 3469 1428 3470
rect 1422 3465 1423 3469
rect 1427 3465 1428 3469
rect 1422 3464 1428 3465
rect 1322 3447 1328 3448
rect 1322 3443 1323 3447
rect 1327 3443 1328 3447
rect 1322 3442 1328 3443
rect 1424 3423 1426 3464
rect 1079 3422 1083 3423
rect 1079 3417 1083 3418
rect 1127 3422 1131 3423
rect 1127 3417 1131 3418
rect 1247 3422 1251 3423
rect 1247 3417 1251 3418
rect 1295 3422 1299 3423
rect 1295 3417 1299 3418
rect 1423 3422 1427 3423
rect 1423 3417 1427 3418
rect 1463 3422 1467 3423
rect 1463 3417 1467 3418
rect 1128 3396 1130 3417
rect 1296 3396 1298 3417
rect 1464 3396 1466 3417
rect 1500 3416 1502 3474
rect 1598 3469 1604 3470
rect 1598 3465 1599 3469
rect 1603 3465 1604 3469
rect 1598 3464 1604 3465
rect 1600 3423 1602 3464
rect 1740 3448 1742 3474
rect 1774 3469 1780 3470
rect 1774 3465 1775 3469
rect 1779 3465 1780 3469
rect 1774 3464 1780 3465
rect 2006 3468 2012 3469
rect 2006 3464 2007 3468
rect 2011 3464 2012 3468
rect 1714 3447 1720 3448
rect 1714 3443 1715 3447
rect 1719 3443 1720 3447
rect 1714 3442 1720 3443
rect 1738 3447 1744 3448
rect 1738 3443 1739 3447
rect 1743 3443 1744 3447
rect 1738 3442 1744 3443
rect 1599 3422 1603 3423
rect 1599 3417 1603 3418
rect 1639 3422 1643 3423
rect 1639 3417 1643 3418
rect 1498 3415 1504 3416
rect 1498 3411 1499 3415
rect 1503 3411 1504 3415
rect 1498 3410 1504 3411
rect 1640 3396 1642 3417
rect 1126 3395 1132 3396
rect 1126 3391 1127 3395
rect 1131 3391 1132 3395
rect 1126 3390 1132 3391
rect 1294 3395 1300 3396
rect 1294 3391 1295 3395
rect 1299 3391 1300 3395
rect 1294 3390 1300 3391
rect 1462 3395 1468 3396
rect 1462 3391 1463 3395
rect 1467 3391 1468 3395
rect 1462 3390 1468 3391
rect 1638 3395 1644 3396
rect 1638 3391 1639 3395
rect 1643 3391 1644 3395
rect 1638 3390 1644 3391
rect 1716 3388 1718 3442
rect 1776 3423 1778 3464
rect 2006 3463 2012 3464
rect 2008 3423 2010 3463
rect 2048 3455 2050 3475
rect 2328 3455 2330 3476
rect 2404 3460 2406 3486
rect 2446 3481 2452 3482
rect 2446 3477 2447 3481
rect 2451 3477 2452 3481
rect 2446 3476 2452 3477
rect 2402 3459 2408 3460
rect 2402 3455 2403 3459
rect 2407 3455 2408 3459
rect 2448 3455 2450 3476
rect 2514 3475 2520 3476
rect 2514 3471 2515 3475
rect 2519 3471 2520 3475
rect 2514 3470 2520 3471
rect 2047 3454 2051 3455
rect 2047 3449 2051 3450
rect 2327 3454 2331 3455
rect 2402 3454 2408 3455
rect 2447 3454 2451 3455
rect 2327 3449 2331 3450
rect 2447 3449 2451 3450
rect 2048 3429 2050 3449
rect 2046 3428 2052 3429
rect 2448 3428 2450 3449
rect 2516 3448 2518 3470
rect 2524 3460 2526 3486
rect 2582 3481 2588 3482
rect 2582 3477 2583 3481
rect 2587 3477 2588 3481
rect 2582 3476 2588 3477
rect 2522 3459 2528 3460
rect 2522 3455 2523 3459
rect 2527 3455 2528 3459
rect 2584 3455 2586 3476
rect 2600 3468 2602 3570
rect 2670 3564 2676 3565
rect 2670 3560 2671 3564
rect 2675 3560 2676 3564
rect 2670 3559 2676 3560
rect 2870 3564 2876 3565
rect 2870 3560 2871 3564
rect 2875 3560 2876 3564
rect 2870 3559 2876 3560
rect 2672 3531 2674 3559
rect 2872 3531 2874 3559
rect 2671 3530 2675 3531
rect 2671 3525 2675 3526
rect 2735 3530 2739 3531
rect 2735 3525 2739 3526
rect 2871 3530 2875 3531
rect 2871 3525 2875 3526
rect 2911 3530 2915 3531
rect 2911 3525 2915 3526
rect 2736 3501 2738 3525
rect 2912 3501 2914 3525
rect 2734 3500 2740 3501
rect 2734 3496 2735 3500
rect 2739 3496 2740 3500
rect 2734 3495 2740 3496
rect 2910 3500 2916 3501
rect 2910 3496 2911 3500
rect 2915 3496 2916 3500
rect 2910 3495 2916 3496
rect 2980 3492 2982 3598
rect 3064 3584 3066 3605
rect 3188 3604 3190 3646
rect 3196 3620 3198 3646
rect 3294 3641 3300 3642
rect 3294 3637 3295 3641
rect 3299 3637 3300 3641
rect 3294 3636 3300 3637
rect 3194 3619 3200 3620
rect 3194 3615 3195 3619
rect 3199 3615 3200 3619
rect 3194 3614 3200 3615
rect 3296 3611 3298 3636
rect 3380 3620 3382 3646
rect 3478 3641 3484 3642
rect 3478 3637 3479 3641
rect 3483 3637 3484 3641
rect 3478 3636 3484 3637
rect 3378 3619 3384 3620
rect 3378 3615 3379 3619
rect 3383 3615 3384 3619
rect 3378 3614 3384 3615
rect 3480 3611 3482 3636
rect 3588 3620 3590 3734
rect 3686 3732 3692 3733
rect 3686 3728 3687 3732
rect 3691 3728 3692 3732
rect 3686 3727 3692 3728
rect 3688 3691 3690 3727
rect 3671 3690 3675 3691
rect 3671 3685 3675 3686
rect 3687 3690 3691 3691
rect 3687 3685 3691 3686
rect 3672 3661 3674 3685
rect 3670 3660 3676 3661
rect 3670 3656 3671 3660
rect 3675 3656 3676 3660
rect 3670 3655 3676 3656
rect 3748 3652 3750 3766
rect 3840 3752 3842 3773
rect 3908 3772 3910 3826
rect 3942 3820 3948 3821
rect 3942 3816 3943 3820
rect 3947 3816 3948 3820
rect 3942 3815 3948 3816
rect 3944 3779 3946 3815
rect 3943 3778 3947 3779
rect 3943 3773 3947 3774
rect 3906 3771 3912 3772
rect 3906 3767 3907 3771
rect 3911 3767 3912 3771
rect 3906 3766 3912 3767
rect 3944 3753 3946 3773
rect 3942 3752 3948 3753
rect 3838 3751 3844 3752
rect 3838 3747 3839 3751
rect 3843 3747 3844 3751
rect 3942 3748 3943 3752
rect 3947 3748 3948 3752
rect 3942 3747 3948 3748
rect 3838 3746 3844 3747
rect 3906 3735 3912 3736
rect 3838 3732 3844 3733
rect 3838 3728 3839 3732
rect 3843 3728 3844 3732
rect 3906 3731 3907 3735
rect 3911 3731 3912 3735
rect 3906 3730 3912 3731
rect 3942 3735 3948 3736
rect 3942 3731 3943 3735
rect 3947 3731 3948 3735
rect 3942 3730 3948 3731
rect 3838 3727 3844 3728
rect 3840 3691 3842 3727
rect 3839 3690 3843 3691
rect 3839 3685 3843 3686
rect 3840 3661 3842 3685
rect 3838 3660 3844 3661
rect 3838 3656 3839 3660
rect 3843 3656 3844 3660
rect 3838 3655 3844 3656
rect 3746 3651 3752 3652
rect 3746 3647 3747 3651
rect 3751 3647 3752 3651
rect 3746 3646 3752 3647
rect 3670 3641 3676 3642
rect 3670 3637 3671 3641
rect 3675 3637 3676 3641
rect 3670 3636 3676 3637
rect 3838 3641 3844 3642
rect 3838 3637 3839 3641
rect 3843 3637 3844 3641
rect 3838 3636 3844 3637
rect 3586 3619 3592 3620
rect 3586 3615 3587 3619
rect 3591 3615 3592 3619
rect 3586 3614 3592 3615
rect 3672 3611 3674 3636
rect 3714 3619 3720 3620
rect 3714 3615 3715 3619
rect 3719 3615 3720 3619
rect 3714 3614 3720 3615
rect 3255 3610 3259 3611
rect 3255 3605 3259 3606
rect 3295 3610 3299 3611
rect 3295 3605 3299 3606
rect 3447 3610 3451 3611
rect 3447 3605 3451 3606
rect 3479 3610 3483 3611
rect 3479 3605 3483 3606
rect 3639 3610 3643 3611
rect 3639 3605 3643 3606
rect 3671 3610 3675 3611
rect 3671 3605 3675 3606
rect 3186 3603 3192 3604
rect 3186 3599 3187 3603
rect 3191 3599 3192 3603
rect 3186 3598 3192 3599
rect 3256 3584 3258 3605
rect 3330 3603 3336 3604
rect 3330 3599 3331 3603
rect 3335 3599 3336 3603
rect 3330 3598 3336 3599
rect 3062 3583 3068 3584
rect 3062 3579 3063 3583
rect 3067 3579 3068 3583
rect 3062 3578 3068 3579
rect 3254 3583 3260 3584
rect 3254 3579 3255 3583
rect 3259 3579 3260 3583
rect 3254 3578 3260 3579
rect 3332 3576 3334 3598
rect 3448 3584 3450 3605
rect 3522 3603 3528 3604
rect 3522 3599 3523 3603
rect 3527 3599 3528 3603
rect 3522 3598 3528 3599
rect 3446 3583 3452 3584
rect 3446 3579 3447 3583
rect 3451 3579 3452 3583
rect 3446 3578 3452 3579
rect 3524 3576 3526 3598
rect 3640 3584 3642 3605
rect 3638 3583 3644 3584
rect 3638 3579 3639 3583
rect 3643 3579 3644 3583
rect 3638 3578 3644 3579
rect 3716 3576 3718 3614
rect 3840 3611 3842 3636
rect 3908 3620 3910 3730
rect 3944 3691 3946 3730
rect 3943 3690 3947 3691
rect 3943 3685 3947 3686
rect 3944 3658 3946 3685
rect 3942 3657 3948 3658
rect 3942 3653 3943 3657
rect 3947 3653 3948 3657
rect 3942 3652 3948 3653
rect 3914 3651 3920 3652
rect 3914 3647 3915 3651
rect 3919 3647 3920 3651
rect 3914 3646 3920 3647
rect 3906 3619 3912 3620
rect 3906 3615 3907 3619
rect 3911 3615 3912 3619
rect 3906 3614 3912 3615
rect 3839 3610 3843 3611
rect 3839 3605 3843 3606
rect 3840 3584 3842 3605
rect 3916 3604 3918 3646
rect 3942 3640 3948 3641
rect 3942 3636 3943 3640
rect 3947 3636 3948 3640
rect 3942 3635 3948 3636
rect 3944 3611 3946 3635
rect 3943 3610 3947 3611
rect 3943 3605 3947 3606
rect 3914 3603 3920 3604
rect 3914 3599 3915 3603
rect 3919 3599 3920 3603
rect 3914 3598 3920 3599
rect 3944 3585 3946 3605
rect 3942 3584 3948 3585
rect 3838 3583 3844 3584
rect 3838 3579 3839 3583
rect 3843 3579 3844 3583
rect 3942 3580 3943 3584
rect 3947 3580 3948 3584
rect 3942 3579 3948 3580
rect 3838 3578 3844 3579
rect 3330 3575 3336 3576
rect 3330 3571 3331 3575
rect 3335 3571 3336 3575
rect 3330 3570 3336 3571
rect 3522 3575 3528 3576
rect 3522 3571 3523 3575
rect 3527 3571 3528 3575
rect 3522 3570 3528 3571
rect 3714 3575 3720 3576
rect 3714 3571 3715 3575
rect 3719 3571 3720 3575
rect 3714 3570 3720 3571
rect 3914 3571 3920 3572
rect 3914 3567 3915 3571
rect 3919 3567 3920 3571
rect 3914 3566 3920 3567
rect 3942 3567 3948 3568
rect 3062 3564 3068 3565
rect 3062 3560 3063 3564
rect 3067 3560 3068 3564
rect 3062 3559 3068 3560
rect 3254 3564 3260 3565
rect 3254 3560 3255 3564
rect 3259 3560 3260 3564
rect 3254 3559 3260 3560
rect 3446 3564 3452 3565
rect 3446 3560 3447 3564
rect 3451 3560 3452 3564
rect 3446 3559 3452 3560
rect 3638 3564 3644 3565
rect 3638 3560 3639 3564
rect 3643 3560 3644 3564
rect 3638 3559 3644 3560
rect 3838 3564 3844 3565
rect 3838 3560 3839 3564
rect 3843 3560 3844 3564
rect 3838 3559 3844 3560
rect 3064 3531 3066 3559
rect 3256 3531 3258 3559
rect 3448 3531 3450 3559
rect 3640 3531 3642 3559
rect 3840 3531 3842 3559
rect 3063 3530 3067 3531
rect 3063 3525 3067 3526
rect 3111 3530 3115 3531
rect 3111 3525 3115 3526
rect 3255 3530 3259 3531
rect 3255 3525 3259 3526
rect 3335 3530 3339 3531
rect 3335 3525 3339 3526
rect 3447 3530 3451 3531
rect 3447 3525 3451 3526
rect 3567 3530 3571 3531
rect 3567 3525 3571 3526
rect 3639 3530 3643 3531
rect 3639 3525 3643 3526
rect 3807 3530 3811 3531
rect 3807 3525 3811 3526
rect 3839 3530 3843 3531
rect 3839 3525 3843 3526
rect 3112 3501 3114 3525
rect 3336 3501 3338 3525
rect 3568 3501 3570 3525
rect 3808 3501 3810 3525
rect 3110 3500 3116 3501
rect 3110 3496 3111 3500
rect 3115 3496 3116 3500
rect 3110 3495 3116 3496
rect 3334 3500 3340 3501
rect 3334 3496 3335 3500
rect 3339 3496 3340 3500
rect 3334 3495 3340 3496
rect 3566 3500 3572 3501
rect 3566 3496 3567 3500
rect 3571 3496 3572 3500
rect 3566 3495 3572 3496
rect 3806 3500 3812 3501
rect 3806 3496 3807 3500
rect 3811 3496 3812 3500
rect 3806 3495 3812 3496
rect 2710 3491 2716 3492
rect 2710 3487 2711 3491
rect 2715 3487 2716 3491
rect 2710 3486 2716 3487
rect 2978 3491 2984 3492
rect 2978 3487 2979 3491
rect 2983 3487 2984 3491
rect 2978 3486 2984 3487
rect 2994 3491 3000 3492
rect 2994 3487 2995 3491
rect 2999 3487 3000 3491
rect 2994 3486 3000 3487
rect 3194 3491 3200 3492
rect 3194 3487 3195 3491
rect 3199 3487 3200 3491
rect 3194 3486 3200 3487
rect 3418 3491 3424 3492
rect 3418 3487 3419 3491
rect 3423 3487 3424 3491
rect 3418 3486 3424 3487
rect 3874 3491 3880 3492
rect 3874 3487 3875 3491
rect 3879 3487 3880 3491
rect 3874 3486 3880 3487
rect 2598 3467 2604 3468
rect 2598 3463 2599 3467
rect 2603 3463 2604 3467
rect 2598 3462 2604 3463
rect 2712 3460 2714 3486
rect 2734 3481 2740 3482
rect 2734 3477 2735 3481
rect 2739 3477 2740 3481
rect 2734 3476 2740 3477
rect 2910 3481 2916 3482
rect 2910 3477 2911 3481
rect 2915 3477 2916 3481
rect 2910 3476 2916 3477
rect 2710 3459 2716 3460
rect 2710 3455 2711 3459
rect 2715 3455 2716 3459
rect 2736 3455 2738 3476
rect 2912 3455 2914 3476
rect 2996 3460 2998 3486
rect 3110 3481 3116 3482
rect 3110 3477 3111 3481
rect 3115 3477 3116 3481
rect 3110 3476 3116 3477
rect 2994 3459 3000 3460
rect 2994 3455 2995 3459
rect 2999 3455 3000 3459
rect 3112 3455 3114 3476
rect 3196 3460 3198 3486
rect 3334 3481 3340 3482
rect 3334 3477 3335 3481
rect 3339 3477 3340 3481
rect 3334 3476 3340 3477
rect 3194 3459 3200 3460
rect 3194 3455 3195 3459
rect 3199 3455 3200 3459
rect 3336 3455 3338 3476
rect 3420 3460 3422 3486
rect 3566 3481 3572 3482
rect 3566 3477 3567 3481
rect 3571 3477 3572 3481
rect 3566 3476 3572 3477
rect 3806 3481 3812 3482
rect 3806 3477 3807 3481
rect 3811 3477 3812 3481
rect 3806 3476 3812 3477
rect 3418 3459 3424 3460
rect 3418 3455 3419 3459
rect 3423 3455 3424 3459
rect 3568 3455 3570 3476
rect 3642 3459 3648 3460
rect 3642 3455 3643 3459
rect 3647 3455 3648 3459
rect 3808 3455 3810 3476
rect 2522 3454 2528 3455
rect 2551 3454 2555 3455
rect 2551 3449 2555 3450
rect 2583 3454 2587 3455
rect 2583 3449 2587 3450
rect 2663 3454 2667 3455
rect 2710 3454 2716 3455
rect 2735 3454 2739 3455
rect 2663 3449 2667 3450
rect 2735 3449 2739 3450
rect 2775 3454 2779 3455
rect 2775 3449 2779 3450
rect 2903 3454 2907 3455
rect 2903 3449 2907 3450
rect 2911 3454 2915 3455
rect 2994 3454 3000 3455
rect 3047 3454 3051 3455
rect 2911 3449 2915 3450
rect 3047 3449 3051 3450
rect 3111 3454 3115 3455
rect 3194 3454 3200 3455
rect 3207 3454 3211 3455
rect 3111 3449 3115 3450
rect 3207 3449 3211 3450
rect 3335 3454 3339 3455
rect 3335 3449 3339 3450
rect 3383 3454 3387 3455
rect 3418 3454 3424 3455
rect 3567 3454 3571 3455
rect 3642 3454 3648 3455
rect 3751 3454 3755 3455
rect 3383 3449 3387 3450
rect 3567 3449 3571 3450
rect 2514 3447 2520 3448
rect 2514 3443 2515 3447
rect 2519 3443 2520 3447
rect 2514 3442 2520 3443
rect 2522 3447 2528 3448
rect 2522 3443 2523 3447
rect 2527 3443 2528 3447
rect 2522 3442 2528 3443
rect 2046 3424 2047 3428
rect 2051 3424 2052 3428
rect 2046 3423 2052 3424
rect 2446 3427 2452 3428
rect 2446 3423 2447 3427
rect 2451 3423 2452 3427
rect 1775 3422 1779 3423
rect 1775 3417 1779 3418
rect 1815 3422 1819 3423
rect 1815 3417 1819 3418
rect 2007 3422 2011 3423
rect 2446 3422 2452 3423
rect 2524 3420 2526 3442
rect 2552 3428 2554 3449
rect 2626 3447 2632 3448
rect 2626 3443 2627 3447
rect 2631 3443 2632 3447
rect 2626 3442 2632 3443
rect 2550 3427 2556 3428
rect 2550 3423 2551 3427
rect 2555 3423 2556 3427
rect 2550 3422 2556 3423
rect 2628 3420 2630 3442
rect 2664 3428 2666 3449
rect 2750 3447 2756 3448
rect 2750 3443 2751 3447
rect 2755 3443 2756 3447
rect 2750 3442 2756 3443
rect 2662 3427 2668 3428
rect 2662 3423 2663 3427
rect 2667 3423 2668 3427
rect 2662 3422 2668 3423
rect 2752 3420 2754 3442
rect 2776 3428 2778 3449
rect 2850 3447 2856 3448
rect 2850 3443 2851 3447
rect 2855 3443 2856 3447
rect 2850 3442 2856 3443
rect 2774 3427 2780 3428
rect 2774 3423 2775 3427
rect 2779 3423 2780 3427
rect 2774 3422 2780 3423
rect 2852 3420 2854 3442
rect 2904 3428 2906 3449
rect 3048 3428 3050 3449
rect 3122 3447 3128 3448
rect 3122 3443 3123 3447
rect 3127 3443 3128 3447
rect 3122 3442 3128 3443
rect 2902 3427 2908 3428
rect 2902 3423 2903 3427
rect 2907 3423 2908 3427
rect 2902 3422 2908 3423
rect 3046 3427 3052 3428
rect 3046 3423 3047 3427
rect 3051 3423 3052 3427
rect 3046 3422 3052 3423
rect 3124 3420 3126 3442
rect 3208 3428 3210 3449
rect 3282 3447 3288 3448
rect 3282 3443 3283 3447
rect 3287 3443 3288 3447
rect 3282 3442 3288 3443
rect 3258 3439 3264 3440
rect 3258 3435 3259 3439
rect 3263 3435 3264 3439
rect 3258 3434 3264 3435
rect 3206 3427 3212 3428
rect 3206 3423 3207 3427
rect 3211 3423 3212 3427
rect 3206 3422 3212 3423
rect 2007 3417 2011 3418
rect 2522 3419 2528 3420
rect 1722 3415 1728 3416
rect 1722 3411 1723 3415
rect 1727 3411 1728 3415
rect 1722 3410 1728 3411
rect 1724 3388 1726 3410
rect 1816 3396 1818 3417
rect 1898 3415 1904 3416
rect 1898 3411 1899 3415
rect 1903 3411 1904 3415
rect 1898 3410 1904 3411
rect 1814 3395 1820 3396
rect 1814 3391 1815 3395
rect 1819 3391 1820 3395
rect 1814 3390 1820 3391
rect 626 3387 632 3388
rect 626 3383 627 3387
rect 631 3383 632 3387
rect 626 3382 632 3383
rect 722 3387 728 3388
rect 722 3383 723 3387
rect 727 3383 728 3387
rect 722 3382 728 3383
rect 874 3387 880 3388
rect 874 3383 875 3387
rect 879 3383 880 3387
rect 874 3382 880 3383
rect 1034 3387 1040 3388
rect 1034 3383 1035 3387
rect 1039 3383 1040 3387
rect 1714 3387 1720 3388
rect 1034 3382 1040 3383
rect 1202 3383 1208 3384
rect 1202 3379 1203 3383
rect 1207 3379 1208 3383
rect 1714 3383 1715 3387
rect 1719 3383 1720 3387
rect 1714 3382 1720 3383
rect 1722 3387 1728 3388
rect 1722 3383 1723 3387
rect 1727 3383 1728 3387
rect 1722 3382 1728 3383
rect 1202 3378 1208 3379
rect 646 3376 652 3377
rect 646 3372 647 3376
rect 651 3372 652 3376
rect 646 3371 652 3372
rect 798 3376 804 3377
rect 798 3372 799 3376
rect 803 3372 804 3376
rect 798 3371 804 3372
rect 958 3376 964 3377
rect 958 3372 959 3376
rect 963 3372 964 3376
rect 958 3371 964 3372
rect 1126 3376 1132 3377
rect 1126 3372 1127 3376
rect 1131 3372 1132 3376
rect 1126 3371 1132 3372
rect 648 3335 650 3371
rect 800 3335 802 3371
rect 960 3335 962 3371
rect 1128 3335 1130 3371
rect 647 3334 651 3335
rect 647 3329 651 3330
rect 671 3334 675 3335
rect 671 3329 675 3330
rect 799 3334 803 3335
rect 799 3329 803 3330
rect 863 3334 867 3335
rect 863 3329 867 3330
rect 959 3334 963 3335
rect 959 3329 963 3330
rect 1055 3334 1059 3335
rect 1055 3329 1059 3330
rect 1127 3334 1131 3335
rect 1127 3329 1131 3330
rect 672 3305 674 3329
rect 864 3305 866 3329
rect 1056 3305 1058 3329
rect 670 3304 676 3305
rect 670 3300 671 3304
rect 675 3300 676 3304
rect 670 3299 676 3300
rect 862 3304 868 3305
rect 862 3300 863 3304
rect 867 3300 868 3304
rect 862 3299 868 3300
rect 1054 3304 1060 3305
rect 1054 3300 1055 3304
rect 1059 3300 1060 3304
rect 1054 3299 1060 3300
rect 210 3295 216 3296
rect 210 3291 211 3295
rect 215 3291 216 3295
rect 210 3290 216 3291
rect 370 3295 376 3296
rect 370 3291 371 3295
rect 375 3291 376 3295
rect 370 3290 376 3291
rect 386 3295 392 3296
rect 386 3291 387 3295
rect 391 3291 392 3295
rect 386 3290 392 3291
rect 618 3295 624 3296
rect 618 3291 619 3295
rect 623 3291 624 3295
rect 618 3290 624 3291
rect 754 3295 760 3296
rect 754 3291 755 3295
rect 759 3291 760 3295
rect 754 3290 760 3291
rect 1130 3295 1136 3296
rect 1130 3291 1131 3295
rect 1135 3291 1136 3295
rect 1130 3290 1136 3291
rect 134 3285 140 3286
rect 110 3284 116 3285
rect 110 3280 111 3284
rect 115 3280 116 3284
rect 134 3281 135 3285
rect 139 3281 140 3285
rect 134 3280 140 3281
rect 110 3279 116 3280
rect 112 3255 114 3279
rect 136 3255 138 3280
rect 212 3264 214 3290
rect 294 3285 300 3286
rect 294 3281 295 3285
rect 299 3281 300 3285
rect 294 3280 300 3281
rect 210 3263 216 3264
rect 210 3259 211 3263
rect 215 3259 216 3263
rect 210 3258 216 3259
rect 296 3255 298 3280
rect 372 3264 374 3290
rect 370 3263 376 3264
rect 370 3259 371 3263
rect 375 3259 376 3263
rect 370 3258 376 3259
rect 111 3254 115 3255
rect 111 3249 115 3250
rect 135 3254 139 3255
rect 135 3249 139 3250
rect 295 3254 299 3255
rect 295 3249 299 3250
rect 319 3254 323 3255
rect 319 3249 323 3250
rect 112 3229 114 3249
rect 110 3228 116 3229
rect 136 3228 138 3249
rect 320 3228 322 3249
rect 388 3248 390 3290
rect 478 3285 484 3286
rect 478 3281 479 3285
rect 483 3281 484 3285
rect 478 3280 484 3281
rect 670 3285 676 3286
rect 670 3281 671 3285
rect 675 3281 676 3285
rect 670 3280 676 3281
rect 480 3255 482 3280
rect 672 3255 674 3280
rect 756 3264 758 3290
rect 862 3285 868 3286
rect 862 3281 863 3285
rect 867 3281 868 3285
rect 862 3280 868 3281
rect 1054 3285 1060 3286
rect 1054 3281 1055 3285
rect 1059 3281 1060 3285
rect 1054 3280 1060 3281
rect 754 3263 760 3264
rect 754 3259 755 3263
rect 759 3259 760 3263
rect 754 3258 760 3259
rect 864 3255 866 3280
rect 986 3263 992 3264
rect 986 3259 987 3263
rect 991 3259 992 3263
rect 986 3258 992 3259
rect 479 3254 483 3255
rect 479 3249 483 3250
rect 519 3254 523 3255
rect 519 3249 523 3250
rect 671 3254 675 3255
rect 671 3249 675 3250
rect 719 3254 723 3255
rect 719 3249 723 3250
rect 863 3254 867 3255
rect 863 3249 867 3250
rect 911 3254 915 3255
rect 911 3249 915 3250
rect 386 3247 392 3248
rect 386 3243 387 3247
rect 391 3243 392 3247
rect 386 3242 392 3243
rect 520 3228 522 3249
rect 678 3247 684 3248
rect 678 3243 679 3247
rect 683 3243 684 3247
rect 678 3242 684 3243
rect 686 3247 692 3248
rect 686 3243 687 3247
rect 691 3243 692 3247
rect 686 3242 692 3243
rect 110 3224 111 3228
rect 115 3224 116 3228
rect 110 3223 116 3224
rect 134 3227 140 3228
rect 134 3223 135 3227
rect 139 3223 140 3227
rect 134 3222 140 3223
rect 318 3227 324 3228
rect 318 3223 319 3227
rect 323 3223 324 3227
rect 318 3222 324 3223
rect 518 3227 524 3228
rect 518 3223 519 3227
rect 523 3223 524 3227
rect 518 3222 524 3223
rect 210 3215 216 3216
rect 110 3211 116 3212
rect 110 3207 111 3211
rect 115 3207 116 3211
rect 210 3211 211 3215
rect 215 3211 216 3215
rect 210 3210 216 3211
rect 110 3206 116 3207
rect 134 3208 140 3209
rect 112 3171 114 3206
rect 134 3204 135 3208
rect 139 3204 140 3208
rect 134 3203 140 3204
rect 136 3171 138 3203
rect 111 3170 115 3171
rect 111 3165 115 3166
rect 135 3170 139 3171
rect 135 3165 139 3166
rect 143 3170 147 3171
rect 143 3165 147 3166
rect 112 3138 114 3165
rect 144 3141 146 3165
rect 142 3140 148 3141
rect 110 3137 116 3138
rect 110 3133 111 3137
rect 115 3133 116 3137
rect 142 3136 143 3140
rect 147 3136 148 3140
rect 142 3135 148 3136
rect 110 3132 116 3133
rect 142 3121 148 3122
rect 110 3120 116 3121
rect 110 3116 111 3120
rect 115 3116 116 3120
rect 142 3117 143 3121
rect 147 3117 148 3121
rect 142 3116 148 3117
rect 110 3115 116 3116
rect 112 3095 114 3115
rect 144 3095 146 3116
rect 212 3100 214 3210
rect 318 3208 324 3209
rect 318 3204 319 3208
rect 323 3204 324 3208
rect 318 3203 324 3204
rect 518 3208 524 3209
rect 518 3204 519 3208
rect 523 3204 524 3208
rect 518 3203 524 3204
rect 320 3171 322 3203
rect 520 3171 522 3203
rect 319 3170 323 3171
rect 319 3165 323 3166
rect 343 3170 347 3171
rect 343 3165 347 3166
rect 519 3170 523 3171
rect 519 3165 523 3166
rect 543 3170 547 3171
rect 543 3165 547 3166
rect 344 3141 346 3165
rect 544 3141 546 3165
rect 342 3140 348 3141
rect 342 3136 343 3140
rect 347 3136 348 3140
rect 342 3135 348 3136
rect 542 3140 548 3141
rect 542 3136 543 3140
rect 547 3136 548 3140
rect 542 3135 548 3136
rect 680 3132 682 3242
rect 688 3220 690 3242
rect 720 3228 722 3249
rect 794 3247 800 3248
rect 794 3243 795 3247
rect 799 3243 800 3247
rect 794 3242 800 3243
rect 718 3227 724 3228
rect 718 3223 719 3227
rect 723 3223 724 3227
rect 718 3222 724 3223
rect 796 3220 798 3242
rect 912 3228 914 3249
rect 910 3227 916 3228
rect 910 3223 911 3227
rect 915 3223 916 3227
rect 910 3222 916 3223
rect 988 3220 990 3258
rect 1056 3255 1058 3280
rect 1055 3254 1059 3255
rect 1055 3249 1059 3250
rect 1095 3254 1099 3255
rect 1095 3249 1099 3250
rect 1096 3228 1098 3249
rect 1132 3248 1134 3290
rect 1204 3264 1206 3378
rect 1294 3376 1300 3377
rect 1294 3372 1295 3376
rect 1299 3372 1300 3376
rect 1294 3371 1300 3372
rect 1462 3376 1468 3377
rect 1462 3372 1463 3376
rect 1467 3372 1468 3376
rect 1462 3371 1468 3372
rect 1638 3376 1644 3377
rect 1638 3372 1639 3376
rect 1643 3372 1644 3376
rect 1638 3371 1644 3372
rect 1814 3376 1820 3377
rect 1814 3372 1815 3376
rect 1819 3372 1820 3376
rect 1814 3371 1820 3372
rect 1296 3335 1298 3371
rect 1464 3335 1466 3371
rect 1640 3335 1642 3371
rect 1816 3335 1818 3371
rect 1247 3334 1251 3335
rect 1247 3329 1251 3330
rect 1295 3334 1299 3335
rect 1295 3329 1299 3330
rect 1439 3334 1443 3335
rect 1439 3329 1443 3330
rect 1463 3334 1467 3335
rect 1463 3329 1467 3330
rect 1631 3334 1635 3335
rect 1631 3329 1635 3330
rect 1639 3334 1643 3335
rect 1639 3329 1643 3330
rect 1815 3334 1819 3335
rect 1815 3329 1819 3330
rect 1823 3334 1827 3335
rect 1823 3329 1827 3330
rect 1248 3305 1250 3329
rect 1440 3305 1442 3329
rect 1632 3305 1634 3329
rect 1824 3305 1826 3329
rect 1246 3304 1252 3305
rect 1246 3300 1247 3304
rect 1251 3300 1252 3304
rect 1246 3299 1252 3300
rect 1438 3304 1444 3305
rect 1438 3300 1439 3304
rect 1443 3300 1444 3304
rect 1438 3299 1444 3300
rect 1630 3304 1636 3305
rect 1630 3300 1631 3304
rect 1635 3300 1636 3304
rect 1630 3299 1636 3300
rect 1822 3304 1828 3305
rect 1822 3300 1823 3304
rect 1827 3300 1828 3304
rect 1822 3299 1828 3300
rect 1900 3296 1902 3410
rect 2008 3397 2010 3417
rect 2522 3415 2523 3419
rect 2527 3415 2528 3419
rect 2522 3414 2528 3415
rect 2626 3419 2632 3420
rect 2626 3415 2627 3419
rect 2631 3415 2632 3419
rect 2626 3414 2632 3415
rect 2750 3419 2756 3420
rect 2750 3415 2751 3419
rect 2755 3415 2756 3419
rect 2750 3414 2756 3415
rect 2850 3419 2856 3420
rect 2850 3415 2851 3419
rect 2855 3415 2856 3419
rect 3122 3419 3128 3420
rect 2850 3414 2856 3415
rect 2978 3415 2984 3416
rect 2046 3411 2052 3412
rect 2046 3407 2047 3411
rect 2051 3407 2052 3411
rect 2978 3411 2979 3415
rect 2983 3411 2984 3415
rect 3122 3415 3123 3419
rect 3127 3415 3128 3419
rect 3122 3414 3128 3415
rect 2978 3410 2984 3411
rect 2046 3406 2052 3407
rect 2446 3408 2452 3409
rect 2006 3396 2012 3397
rect 2006 3392 2007 3396
rect 2011 3392 2012 3396
rect 2006 3391 2012 3392
rect 2006 3379 2012 3380
rect 2006 3375 2007 3379
rect 2011 3375 2012 3379
rect 2006 3374 2012 3375
rect 2008 3335 2010 3374
rect 2048 3367 2050 3406
rect 2446 3404 2447 3408
rect 2451 3404 2452 3408
rect 2446 3403 2452 3404
rect 2550 3408 2556 3409
rect 2550 3404 2551 3408
rect 2555 3404 2556 3408
rect 2550 3403 2556 3404
rect 2662 3408 2668 3409
rect 2662 3404 2663 3408
rect 2667 3404 2668 3408
rect 2662 3403 2668 3404
rect 2774 3408 2780 3409
rect 2774 3404 2775 3408
rect 2779 3404 2780 3408
rect 2774 3403 2780 3404
rect 2902 3408 2908 3409
rect 2902 3404 2903 3408
rect 2907 3404 2908 3408
rect 2902 3403 2908 3404
rect 2448 3367 2450 3403
rect 2552 3367 2554 3403
rect 2664 3367 2666 3403
rect 2776 3367 2778 3403
rect 2904 3367 2906 3403
rect 2047 3366 2051 3367
rect 2047 3361 2051 3362
rect 2447 3366 2451 3367
rect 2447 3361 2451 3362
rect 2551 3366 2555 3367
rect 2551 3361 2555 3362
rect 2567 3366 2571 3367
rect 2567 3361 2571 3362
rect 2663 3366 2667 3367
rect 2663 3361 2667 3362
rect 2719 3366 2723 3367
rect 2719 3361 2723 3362
rect 2775 3366 2779 3367
rect 2775 3361 2779 3362
rect 2871 3366 2875 3367
rect 2871 3361 2875 3362
rect 2903 3366 2907 3367
rect 2903 3361 2907 3362
rect 2007 3334 2011 3335
rect 2048 3334 2050 3361
rect 2568 3337 2570 3361
rect 2720 3337 2722 3361
rect 2872 3337 2874 3361
rect 2566 3336 2572 3337
rect 2007 3329 2011 3330
rect 2046 3333 2052 3334
rect 2046 3329 2047 3333
rect 2051 3329 2052 3333
rect 2566 3332 2567 3336
rect 2571 3332 2572 3336
rect 2566 3331 2572 3332
rect 2718 3336 2724 3337
rect 2718 3332 2719 3336
rect 2723 3332 2724 3336
rect 2718 3331 2724 3332
rect 2870 3336 2876 3337
rect 2870 3332 2871 3336
rect 2875 3332 2876 3336
rect 2870 3331 2876 3332
rect 2008 3302 2010 3329
rect 2046 3328 2052 3329
rect 2642 3327 2648 3328
rect 2642 3323 2643 3327
rect 2647 3323 2648 3327
rect 2642 3322 2648 3323
rect 2650 3327 2656 3328
rect 2650 3323 2651 3327
rect 2655 3323 2656 3327
rect 2650 3322 2656 3323
rect 2802 3327 2808 3328
rect 2802 3323 2803 3327
rect 2807 3323 2808 3327
rect 2802 3322 2808 3323
rect 2954 3327 2960 3328
rect 2954 3323 2955 3327
rect 2959 3323 2960 3327
rect 2954 3322 2960 3323
rect 2566 3317 2572 3318
rect 2046 3316 2052 3317
rect 2046 3312 2047 3316
rect 2051 3312 2052 3316
rect 2566 3313 2567 3317
rect 2571 3313 2572 3317
rect 2566 3312 2572 3313
rect 2046 3311 2052 3312
rect 2006 3301 2012 3302
rect 2006 3297 2007 3301
rect 2011 3297 2012 3301
rect 2006 3296 2012 3297
rect 1322 3295 1328 3296
rect 1322 3291 1323 3295
rect 1327 3291 1328 3295
rect 1322 3290 1328 3291
rect 1338 3295 1344 3296
rect 1338 3291 1339 3295
rect 1343 3291 1344 3295
rect 1338 3290 1344 3291
rect 1778 3295 1784 3296
rect 1778 3291 1779 3295
rect 1783 3291 1784 3295
rect 1778 3290 1784 3291
rect 1898 3295 1904 3296
rect 1898 3291 1899 3295
rect 1903 3291 1904 3295
rect 1898 3290 1904 3291
rect 1246 3285 1252 3286
rect 1246 3281 1247 3285
rect 1251 3281 1252 3285
rect 1246 3280 1252 3281
rect 1202 3263 1208 3264
rect 1202 3259 1203 3263
rect 1207 3259 1208 3263
rect 1202 3258 1208 3259
rect 1248 3255 1250 3280
rect 1324 3264 1326 3290
rect 1340 3272 1342 3290
rect 1438 3285 1444 3286
rect 1438 3281 1439 3285
rect 1443 3281 1444 3285
rect 1438 3280 1444 3281
rect 1630 3285 1636 3286
rect 1630 3281 1631 3285
rect 1635 3281 1636 3285
rect 1630 3280 1636 3281
rect 1338 3271 1344 3272
rect 1338 3267 1339 3271
rect 1343 3267 1344 3271
rect 1338 3266 1344 3267
rect 1322 3263 1328 3264
rect 1322 3259 1323 3263
rect 1327 3259 1328 3263
rect 1322 3258 1328 3259
rect 1440 3255 1442 3280
rect 1632 3255 1634 3280
rect 1780 3264 1782 3290
rect 2048 3287 2050 3311
rect 2568 3287 2570 3312
rect 2047 3286 2051 3287
rect 1822 3285 1828 3286
rect 1822 3281 1823 3285
rect 1827 3281 1828 3285
rect 1822 3280 1828 3281
rect 2006 3284 2012 3285
rect 2006 3280 2007 3284
rect 2011 3280 2012 3284
rect 2047 3281 2051 3282
rect 2415 3286 2419 3287
rect 2415 3281 2419 3282
rect 2551 3286 2555 3287
rect 2551 3281 2555 3282
rect 2567 3286 2571 3287
rect 2567 3281 2571 3282
rect 1706 3263 1712 3264
rect 1706 3259 1707 3263
rect 1711 3259 1712 3263
rect 1706 3258 1712 3259
rect 1778 3263 1784 3264
rect 1778 3259 1779 3263
rect 1783 3259 1784 3263
rect 1778 3258 1784 3259
rect 1247 3254 1251 3255
rect 1247 3249 1251 3250
rect 1271 3254 1275 3255
rect 1271 3249 1275 3250
rect 1439 3254 1443 3255
rect 1439 3249 1443 3250
rect 1447 3254 1451 3255
rect 1447 3249 1451 3250
rect 1623 3254 1627 3255
rect 1623 3249 1627 3250
rect 1631 3254 1635 3255
rect 1631 3249 1635 3250
rect 1130 3247 1136 3248
rect 1130 3243 1131 3247
rect 1135 3243 1136 3247
rect 1130 3242 1136 3243
rect 1170 3247 1176 3248
rect 1170 3243 1171 3247
rect 1175 3243 1176 3247
rect 1170 3242 1176 3243
rect 1094 3227 1100 3228
rect 1094 3223 1095 3227
rect 1099 3223 1100 3227
rect 1094 3222 1100 3223
rect 1172 3220 1174 3242
rect 1272 3228 1274 3249
rect 1346 3247 1352 3248
rect 1346 3243 1347 3247
rect 1351 3243 1352 3247
rect 1346 3242 1352 3243
rect 1270 3227 1276 3228
rect 1270 3223 1271 3227
rect 1275 3223 1276 3227
rect 1270 3222 1276 3223
rect 1348 3220 1350 3242
rect 1448 3228 1450 3249
rect 1624 3228 1626 3249
rect 1650 3247 1656 3248
rect 1650 3243 1651 3247
rect 1655 3243 1656 3247
rect 1650 3242 1656 3243
rect 1698 3247 1704 3248
rect 1698 3243 1699 3247
rect 1703 3243 1704 3247
rect 1698 3242 1704 3243
rect 1446 3227 1452 3228
rect 1446 3223 1447 3227
rect 1451 3223 1452 3227
rect 1446 3222 1452 3223
rect 1622 3227 1628 3228
rect 1622 3223 1623 3227
rect 1627 3223 1628 3227
rect 1622 3222 1628 3223
rect 686 3219 692 3220
rect 686 3215 687 3219
rect 691 3215 692 3219
rect 686 3214 692 3215
rect 794 3219 800 3220
rect 794 3215 795 3219
rect 799 3215 800 3219
rect 794 3214 800 3215
rect 986 3219 992 3220
rect 986 3215 987 3219
rect 991 3215 992 3219
rect 986 3214 992 3215
rect 1170 3219 1176 3220
rect 1170 3215 1171 3219
rect 1175 3215 1176 3219
rect 1170 3214 1176 3215
rect 1346 3219 1352 3220
rect 1346 3215 1347 3219
rect 1351 3215 1352 3219
rect 1346 3214 1352 3215
rect 1522 3215 1528 3216
rect 1522 3211 1523 3215
rect 1527 3211 1528 3215
rect 1522 3210 1528 3211
rect 718 3208 724 3209
rect 718 3204 719 3208
rect 723 3204 724 3208
rect 718 3203 724 3204
rect 910 3208 916 3209
rect 910 3204 911 3208
rect 915 3204 916 3208
rect 910 3203 916 3204
rect 1094 3208 1100 3209
rect 1094 3204 1095 3208
rect 1099 3204 1100 3208
rect 1094 3203 1100 3204
rect 1270 3208 1276 3209
rect 1270 3204 1271 3208
rect 1275 3204 1276 3208
rect 1270 3203 1276 3204
rect 1446 3208 1452 3209
rect 1446 3204 1447 3208
rect 1451 3204 1452 3208
rect 1446 3203 1452 3204
rect 720 3171 722 3203
rect 912 3171 914 3203
rect 1096 3171 1098 3203
rect 1272 3171 1274 3203
rect 1448 3171 1450 3203
rect 719 3170 723 3171
rect 719 3165 723 3166
rect 743 3170 747 3171
rect 743 3165 747 3166
rect 911 3170 915 3171
rect 911 3165 915 3166
rect 927 3170 931 3171
rect 927 3165 931 3166
rect 1095 3170 1099 3171
rect 1095 3165 1099 3166
rect 1103 3170 1107 3171
rect 1103 3165 1107 3166
rect 1263 3170 1267 3171
rect 1263 3165 1267 3166
rect 1271 3170 1275 3171
rect 1271 3165 1275 3166
rect 1423 3170 1427 3171
rect 1423 3165 1427 3166
rect 1447 3170 1451 3171
rect 1447 3165 1451 3166
rect 744 3141 746 3165
rect 928 3141 930 3165
rect 1104 3141 1106 3165
rect 1264 3141 1266 3165
rect 1424 3141 1426 3165
rect 742 3140 748 3141
rect 742 3136 743 3140
rect 747 3136 748 3140
rect 742 3135 748 3136
rect 926 3140 932 3141
rect 926 3136 927 3140
rect 931 3136 932 3140
rect 926 3135 932 3136
rect 1102 3140 1108 3141
rect 1102 3136 1103 3140
rect 1107 3136 1108 3140
rect 1102 3135 1108 3136
rect 1262 3140 1268 3141
rect 1262 3136 1263 3140
rect 1267 3136 1268 3140
rect 1262 3135 1268 3136
rect 1422 3140 1428 3141
rect 1422 3136 1423 3140
rect 1427 3136 1428 3140
rect 1422 3135 1428 3136
rect 218 3131 224 3132
rect 218 3127 219 3131
rect 223 3127 224 3131
rect 218 3126 224 3127
rect 418 3131 424 3132
rect 418 3127 419 3131
rect 423 3127 424 3131
rect 418 3126 424 3127
rect 630 3131 636 3132
rect 630 3127 631 3131
rect 635 3127 636 3131
rect 630 3126 636 3127
rect 678 3131 684 3132
rect 678 3127 679 3131
rect 683 3127 684 3131
rect 678 3126 684 3127
rect 826 3131 832 3132
rect 826 3127 827 3131
rect 831 3127 832 3131
rect 826 3126 832 3127
rect 1178 3131 1184 3132
rect 1178 3127 1179 3131
rect 1183 3127 1184 3131
rect 1178 3126 1184 3127
rect 1186 3131 1192 3132
rect 1186 3127 1187 3131
rect 1191 3127 1192 3131
rect 1186 3126 1192 3127
rect 1346 3131 1352 3132
rect 1346 3127 1347 3131
rect 1351 3127 1352 3131
rect 1346 3126 1352 3127
rect 220 3100 222 3126
rect 342 3121 348 3122
rect 342 3117 343 3121
rect 347 3117 348 3121
rect 342 3116 348 3117
rect 210 3099 216 3100
rect 210 3095 211 3099
rect 215 3095 216 3099
rect 111 3094 115 3095
rect 111 3089 115 3090
rect 143 3094 147 3095
rect 210 3094 216 3095
rect 218 3099 224 3100
rect 218 3095 219 3099
rect 223 3095 224 3099
rect 344 3095 346 3116
rect 420 3100 422 3126
rect 542 3121 548 3122
rect 542 3117 543 3121
rect 547 3117 548 3121
rect 542 3116 548 3117
rect 418 3099 424 3100
rect 418 3095 419 3099
rect 423 3095 424 3099
rect 544 3095 546 3116
rect 218 3094 224 3095
rect 263 3094 267 3095
rect 143 3089 147 3090
rect 263 3089 267 3090
rect 343 3094 347 3095
rect 418 3094 424 3095
rect 439 3094 443 3095
rect 343 3089 347 3090
rect 439 3089 443 3090
rect 543 3094 547 3095
rect 543 3089 547 3090
rect 615 3094 619 3095
rect 615 3089 619 3090
rect 112 3069 114 3089
rect 110 3068 116 3069
rect 264 3068 266 3089
rect 386 3087 392 3088
rect 386 3083 387 3087
rect 391 3083 392 3087
rect 386 3082 392 3083
rect 110 3064 111 3068
rect 115 3064 116 3068
rect 110 3063 116 3064
rect 262 3067 268 3068
rect 262 3063 263 3067
rect 267 3063 268 3067
rect 262 3062 268 3063
rect 388 3060 390 3082
rect 440 3068 442 3089
rect 558 3079 564 3080
rect 558 3075 559 3079
rect 563 3075 564 3079
rect 558 3074 564 3075
rect 438 3067 444 3068
rect 438 3063 439 3067
rect 443 3063 444 3067
rect 438 3062 444 3063
rect 560 3060 562 3074
rect 616 3068 618 3089
rect 632 3088 634 3126
rect 742 3121 748 3122
rect 742 3117 743 3121
rect 747 3117 748 3121
rect 742 3116 748 3117
rect 744 3095 746 3116
rect 828 3100 830 3126
rect 926 3121 932 3122
rect 926 3117 927 3121
rect 931 3117 932 3121
rect 926 3116 932 3117
rect 1102 3121 1108 3122
rect 1102 3117 1103 3121
rect 1107 3117 1108 3121
rect 1102 3116 1108 3117
rect 826 3099 832 3100
rect 826 3095 827 3099
rect 831 3095 832 3099
rect 928 3095 930 3116
rect 1050 3099 1056 3100
rect 1050 3095 1051 3099
rect 1055 3095 1056 3099
rect 1104 3095 1106 3116
rect 743 3094 747 3095
rect 743 3089 747 3090
rect 799 3094 803 3095
rect 826 3094 832 3095
rect 927 3094 931 3095
rect 799 3089 803 3090
rect 927 3089 931 3090
rect 975 3094 979 3095
rect 1050 3094 1056 3095
rect 1103 3094 1107 3095
rect 975 3089 979 3090
rect 630 3087 636 3088
rect 630 3083 631 3087
rect 635 3083 636 3087
rect 630 3082 636 3083
rect 800 3068 802 3089
rect 858 3087 864 3088
rect 858 3083 859 3087
rect 863 3083 864 3087
rect 858 3082 864 3083
rect 874 3087 880 3088
rect 874 3083 875 3087
rect 879 3083 880 3087
rect 874 3082 880 3083
rect 614 3067 620 3068
rect 614 3063 615 3067
rect 619 3063 620 3067
rect 614 3062 620 3063
rect 798 3067 804 3068
rect 798 3063 799 3067
rect 803 3063 804 3067
rect 798 3062 804 3063
rect 386 3059 392 3060
rect 386 3055 387 3059
rect 391 3055 392 3059
rect 558 3059 564 3060
rect 386 3054 392 3055
rect 514 3055 520 3056
rect 110 3051 116 3052
rect 110 3047 111 3051
rect 115 3047 116 3051
rect 514 3051 515 3055
rect 519 3051 520 3055
rect 558 3055 559 3059
rect 563 3055 564 3059
rect 558 3054 564 3055
rect 514 3050 520 3051
rect 110 3046 116 3047
rect 262 3048 268 3049
rect 112 2995 114 3046
rect 262 3044 263 3048
rect 267 3044 268 3048
rect 262 3043 268 3044
rect 438 3048 444 3049
rect 438 3044 439 3048
rect 443 3044 444 3048
rect 438 3043 444 3044
rect 264 2995 266 3043
rect 440 2995 442 3043
rect 111 2994 115 2995
rect 111 2989 115 2990
rect 263 2994 267 2995
rect 263 2989 267 2990
rect 343 2994 347 2995
rect 343 2989 347 2990
rect 439 2994 443 2995
rect 439 2989 443 2990
rect 112 2962 114 2989
rect 344 2965 346 2989
rect 440 2965 442 2989
rect 342 2964 348 2965
rect 110 2961 116 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 342 2960 343 2964
rect 347 2960 348 2964
rect 342 2959 348 2960
rect 438 2964 444 2965
rect 438 2960 439 2964
rect 443 2960 444 2964
rect 438 2959 444 2960
rect 110 2956 116 2957
rect 274 2955 280 2956
rect 274 2951 275 2955
rect 279 2951 280 2955
rect 274 2950 280 2951
rect 426 2955 432 2956
rect 426 2951 427 2955
rect 431 2951 432 2955
rect 426 2950 432 2951
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 110 2939 116 2940
rect 112 2919 114 2939
rect 111 2918 115 2919
rect 111 2913 115 2914
rect 207 2918 211 2919
rect 207 2913 211 2914
rect 112 2893 114 2913
rect 110 2892 116 2893
rect 208 2892 210 2913
rect 276 2912 278 2950
rect 342 2945 348 2946
rect 342 2941 343 2945
rect 347 2941 348 2945
rect 342 2940 348 2941
rect 344 2919 346 2940
rect 428 2924 430 2950
rect 438 2945 444 2946
rect 438 2941 439 2945
rect 443 2941 444 2945
rect 438 2940 444 2941
rect 426 2923 432 2924
rect 426 2919 427 2923
rect 431 2919 432 2923
rect 440 2919 442 2940
rect 516 2924 518 3050
rect 614 3048 620 3049
rect 614 3044 615 3048
rect 619 3044 620 3048
rect 614 3043 620 3044
rect 798 3048 804 3049
rect 798 3044 799 3048
rect 803 3044 804 3048
rect 798 3043 804 3044
rect 616 2995 618 3043
rect 800 2995 802 3043
rect 543 2994 547 2995
rect 543 2989 547 2990
rect 615 2994 619 2995
rect 615 2989 619 2990
rect 655 2994 659 2995
rect 655 2989 659 2990
rect 783 2994 787 2995
rect 783 2989 787 2990
rect 799 2994 803 2995
rect 799 2989 803 2990
rect 544 2965 546 2989
rect 656 2965 658 2989
rect 784 2965 786 2989
rect 542 2964 548 2965
rect 542 2960 543 2964
rect 547 2960 548 2964
rect 542 2959 548 2960
rect 654 2964 660 2965
rect 654 2960 655 2964
rect 659 2960 660 2964
rect 654 2959 660 2960
rect 782 2964 788 2965
rect 782 2960 783 2964
rect 787 2960 788 2964
rect 782 2959 788 2960
rect 860 2956 862 3082
rect 876 3060 878 3082
rect 976 3068 978 3089
rect 974 3067 980 3068
rect 974 3063 975 3067
rect 979 3063 980 3067
rect 974 3062 980 3063
rect 1052 3060 1054 3094
rect 1103 3089 1107 3090
rect 1143 3094 1147 3095
rect 1143 3089 1147 3090
rect 1144 3068 1146 3089
rect 1180 3088 1182 3126
rect 1188 3100 1190 3126
rect 1262 3121 1268 3122
rect 1262 3117 1263 3121
rect 1267 3117 1268 3121
rect 1262 3116 1268 3117
rect 1186 3099 1192 3100
rect 1186 3095 1187 3099
rect 1191 3095 1192 3099
rect 1264 3095 1266 3116
rect 1348 3100 1350 3126
rect 1422 3121 1428 3122
rect 1422 3117 1423 3121
rect 1427 3117 1428 3121
rect 1422 3116 1428 3117
rect 1346 3099 1352 3100
rect 1346 3095 1347 3099
rect 1351 3095 1352 3099
rect 1424 3095 1426 3116
rect 1524 3100 1526 3210
rect 1622 3208 1628 3209
rect 1622 3204 1623 3208
rect 1627 3204 1628 3208
rect 1622 3203 1628 3204
rect 1624 3171 1626 3203
rect 1575 3170 1579 3171
rect 1575 3165 1579 3166
rect 1623 3170 1627 3171
rect 1623 3165 1627 3166
rect 1576 3141 1578 3165
rect 1574 3140 1580 3141
rect 1574 3136 1575 3140
rect 1579 3136 1580 3140
rect 1574 3135 1580 3136
rect 1652 3132 1654 3242
rect 1700 3220 1702 3242
rect 1708 3220 1710 3258
rect 1824 3255 1826 3280
rect 2006 3279 2012 3280
rect 2008 3255 2010 3279
rect 2048 3261 2050 3281
rect 2046 3260 2052 3261
rect 2416 3260 2418 3281
rect 2490 3279 2496 3280
rect 2490 3275 2491 3279
rect 2495 3275 2496 3279
rect 2490 3274 2496 3275
rect 2046 3256 2047 3260
rect 2051 3256 2052 3260
rect 2046 3255 2052 3256
rect 2414 3259 2420 3260
rect 2414 3255 2415 3259
rect 2419 3255 2420 3259
rect 1799 3254 1803 3255
rect 1799 3249 1803 3250
rect 1823 3254 1827 3255
rect 1823 3249 1827 3250
rect 2007 3254 2011 3255
rect 2414 3254 2420 3255
rect 2492 3252 2494 3274
rect 2552 3260 2554 3281
rect 2644 3280 2646 3322
rect 2652 3296 2654 3322
rect 2718 3317 2724 3318
rect 2718 3313 2719 3317
rect 2723 3313 2724 3317
rect 2718 3312 2724 3313
rect 2650 3295 2656 3296
rect 2650 3291 2651 3295
rect 2655 3291 2656 3295
rect 2650 3290 2656 3291
rect 2720 3287 2722 3312
rect 2804 3296 2806 3322
rect 2870 3317 2876 3318
rect 2870 3313 2871 3317
rect 2875 3313 2876 3317
rect 2870 3312 2876 3313
rect 2802 3295 2808 3296
rect 2802 3291 2803 3295
rect 2807 3291 2808 3295
rect 2802 3290 2808 3291
rect 2872 3287 2874 3312
rect 2956 3296 2958 3322
rect 2980 3296 2982 3410
rect 3046 3408 3052 3409
rect 3046 3404 3047 3408
rect 3051 3404 3052 3408
rect 3046 3403 3052 3404
rect 3206 3408 3212 3409
rect 3206 3404 3207 3408
rect 3211 3404 3212 3408
rect 3206 3403 3212 3404
rect 3048 3367 3050 3403
rect 3208 3367 3210 3403
rect 3023 3366 3027 3367
rect 3023 3361 3027 3362
rect 3047 3366 3051 3367
rect 3047 3361 3051 3362
rect 3175 3366 3179 3367
rect 3175 3361 3179 3362
rect 3207 3366 3211 3367
rect 3207 3361 3211 3362
rect 3024 3337 3026 3361
rect 3176 3337 3178 3361
rect 3022 3336 3028 3337
rect 3022 3332 3023 3336
rect 3027 3332 3028 3336
rect 3022 3331 3028 3332
rect 3174 3336 3180 3337
rect 3174 3332 3175 3336
rect 3179 3332 3180 3336
rect 3174 3331 3180 3332
rect 3260 3328 3262 3434
rect 3284 3420 3286 3442
rect 3384 3428 3386 3449
rect 3458 3447 3464 3448
rect 3458 3443 3459 3447
rect 3463 3443 3464 3447
rect 3458 3442 3464 3443
rect 3382 3427 3388 3428
rect 3382 3423 3383 3427
rect 3387 3423 3388 3427
rect 3382 3422 3388 3423
rect 3460 3420 3462 3442
rect 3568 3428 3570 3449
rect 3566 3427 3572 3428
rect 3566 3423 3567 3427
rect 3571 3423 3572 3427
rect 3566 3422 3572 3423
rect 3644 3420 3646 3454
rect 3751 3449 3755 3450
rect 3807 3454 3811 3455
rect 3807 3449 3811 3450
rect 3752 3428 3754 3449
rect 3876 3448 3878 3486
rect 3916 3460 3918 3566
rect 3942 3563 3943 3567
rect 3947 3563 3948 3567
rect 3942 3562 3948 3563
rect 3944 3531 3946 3562
rect 3943 3530 3947 3531
rect 3943 3525 3947 3526
rect 3944 3498 3946 3525
rect 3942 3497 3948 3498
rect 3942 3493 3943 3497
rect 3947 3493 3948 3497
rect 3942 3492 3948 3493
rect 3942 3480 3948 3481
rect 3942 3476 3943 3480
rect 3947 3476 3948 3480
rect 3942 3475 3948 3476
rect 3914 3459 3920 3460
rect 3914 3455 3915 3459
rect 3919 3455 3920 3459
rect 3944 3455 3946 3475
rect 3914 3454 3920 3455
rect 3943 3454 3947 3455
rect 3943 3449 3947 3450
rect 3874 3447 3880 3448
rect 3874 3443 3875 3447
rect 3879 3443 3880 3447
rect 3874 3442 3880 3443
rect 3944 3429 3946 3449
rect 3942 3428 3948 3429
rect 3750 3427 3756 3428
rect 3750 3423 3751 3427
rect 3755 3423 3756 3427
rect 3942 3424 3943 3428
rect 3947 3424 3948 3428
rect 3942 3423 3948 3424
rect 3750 3422 3756 3423
rect 3282 3419 3288 3420
rect 3282 3415 3283 3419
rect 3287 3415 3288 3419
rect 3282 3414 3288 3415
rect 3458 3419 3464 3420
rect 3458 3415 3459 3419
rect 3463 3415 3464 3419
rect 3458 3414 3464 3415
rect 3642 3419 3648 3420
rect 3642 3415 3643 3419
rect 3647 3415 3648 3419
rect 3642 3414 3648 3415
rect 3826 3415 3832 3416
rect 3826 3411 3827 3415
rect 3831 3411 3832 3415
rect 3826 3410 3832 3411
rect 3942 3411 3948 3412
rect 3382 3408 3388 3409
rect 3382 3404 3383 3408
rect 3387 3404 3388 3408
rect 3382 3403 3388 3404
rect 3566 3408 3572 3409
rect 3566 3404 3567 3408
rect 3571 3404 3572 3408
rect 3566 3403 3572 3404
rect 3750 3408 3756 3409
rect 3750 3404 3751 3408
rect 3755 3404 3756 3408
rect 3750 3403 3756 3404
rect 3384 3367 3386 3403
rect 3568 3367 3570 3403
rect 3752 3367 3754 3403
rect 3327 3366 3331 3367
rect 3327 3361 3331 3362
rect 3383 3366 3387 3367
rect 3383 3361 3387 3362
rect 3479 3366 3483 3367
rect 3479 3361 3483 3362
rect 3567 3366 3571 3367
rect 3567 3361 3571 3362
rect 3631 3366 3635 3367
rect 3631 3361 3635 3362
rect 3751 3366 3755 3367
rect 3751 3361 3755 3362
rect 3783 3366 3787 3367
rect 3783 3361 3787 3362
rect 3328 3337 3330 3361
rect 3480 3337 3482 3361
rect 3632 3337 3634 3361
rect 3784 3337 3786 3361
rect 3326 3336 3332 3337
rect 3326 3332 3327 3336
rect 3331 3332 3332 3336
rect 3326 3331 3332 3332
rect 3478 3336 3484 3337
rect 3478 3332 3479 3336
rect 3483 3332 3484 3336
rect 3478 3331 3484 3332
rect 3630 3336 3636 3337
rect 3630 3332 3631 3336
rect 3635 3332 3636 3336
rect 3630 3331 3636 3332
rect 3782 3336 3788 3337
rect 3782 3332 3783 3336
rect 3787 3332 3788 3336
rect 3782 3331 3788 3332
rect 3250 3327 3256 3328
rect 3250 3323 3251 3327
rect 3255 3323 3256 3327
rect 3250 3322 3256 3323
rect 3258 3327 3264 3328
rect 3258 3323 3259 3327
rect 3263 3323 3264 3327
rect 3258 3322 3264 3323
rect 3562 3327 3568 3328
rect 3562 3323 3563 3327
rect 3567 3323 3568 3327
rect 3562 3322 3568 3323
rect 3714 3327 3720 3328
rect 3714 3323 3715 3327
rect 3719 3323 3720 3327
rect 3714 3322 3720 3323
rect 3022 3317 3028 3318
rect 3022 3313 3023 3317
rect 3027 3313 3028 3317
rect 3022 3312 3028 3313
rect 3174 3317 3180 3318
rect 3174 3313 3175 3317
rect 3179 3313 3180 3317
rect 3174 3312 3180 3313
rect 2954 3295 2960 3296
rect 2954 3291 2955 3295
rect 2959 3291 2960 3295
rect 2954 3290 2960 3291
rect 2978 3295 2984 3296
rect 2978 3291 2979 3295
rect 2983 3291 2984 3295
rect 2978 3290 2984 3291
rect 3024 3287 3026 3312
rect 3176 3287 3178 3312
rect 3252 3296 3254 3322
rect 3326 3317 3332 3318
rect 3326 3313 3327 3317
rect 3331 3313 3332 3317
rect 3326 3312 3332 3313
rect 3478 3317 3484 3318
rect 3478 3313 3479 3317
rect 3483 3313 3484 3317
rect 3478 3312 3484 3313
rect 3194 3295 3200 3296
rect 3194 3291 3195 3295
rect 3199 3291 3200 3295
rect 3194 3290 3200 3291
rect 3250 3295 3256 3296
rect 3250 3291 3251 3295
rect 3255 3291 3256 3295
rect 3250 3290 3256 3291
rect 2687 3286 2691 3287
rect 2687 3281 2691 3282
rect 2719 3286 2723 3287
rect 2719 3281 2723 3282
rect 2831 3286 2835 3287
rect 2831 3281 2835 3282
rect 2871 3286 2875 3287
rect 2871 3281 2875 3282
rect 2975 3286 2979 3287
rect 2975 3281 2979 3282
rect 3023 3286 3027 3287
rect 3023 3281 3027 3282
rect 3119 3286 3123 3287
rect 3119 3281 3123 3282
rect 3175 3286 3179 3287
rect 3175 3281 3179 3282
rect 2642 3279 2648 3280
rect 2642 3275 2643 3279
rect 2647 3275 2648 3279
rect 2642 3274 2648 3275
rect 2688 3260 2690 3281
rect 2762 3279 2768 3280
rect 2762 3275 2763 3279
rect 2767 3275 2768 3279
rect 2762 3274 2768 3275
rect 2550 3259 2556 3260
rect 2550 3255 2551 3259
rect 2555 3255 2556 3259
rect 2550 3254 2556 3255
rect 2686 3259 2692 3260
rect 2686 3255 2687 3259
rect 2691 3255 2692 3259
rect 2686 3254 2692 3255
rect 2764 3252 2766 3274
rect 2832 3260 2834 3281
rect 2906 3279 2912 3280
rect 2906 3275 2907 3279
rect 2911 3275 2912 3279
rect 2906 3274 2912 3275
rect 2830 3259 2836 3260
rect 2830 3255 2831 3259
rect 2835 3255 2836 3259
rect 2830 3254 2836 3255
rect 2908 3252 2910 3274
rect 2926 3271 2932 3272
rect 2926 3267 2927 3271
rect 2931 3267 2932 3271
rect 2926 3266 2932 3267
rect 2928 3252 2930 3266
rect 2976 3260 2978 3281
rect 3120 3260 3122 3281
rect 2974 3259 2980 3260
rect 2974 3255 2975 3259
rect 2979 3255 2980 3259
rect 2974 3254 2980 3255
rect 3118 3259 3124 3260
rect 3118 3255 3119 3259
rect 3123 3255 3124 3259
rect 3118 3254 3124 3255
rect 3196 3252 3198 3290
rect 3328 3287 3330 3312
rect 3480 3287 3482 3312
rect 3564 3296 3566 3322
rect 3630 3317 3636 3318
rect 3630 3313 3631 3317
rect 3635 3313 3636 3317
rect 3630 3312 3636 3313
rect 3562 3295 3568 3296
rect 3562 3291 3563 3295
rect 3567 3291 3568 3295
rect 3562 3290 3568 3291
rect 3632 3287 3634 3312
rect 3716 3296 3718 3322
rect 3782 3317 3788 3318
rect 3782 3313 3783 3317
rect 3787 3313 3788 3317
rect 3782 3312 3788 3313
rect 3714 3295 3720 3296
rect 3714 3291 3715 3295
rect 3719 3291 3720 3295
rect 3714 3290 3720 3291
rect 3784 3287 3786 3312
rect 3828 3296 3830 3410
rect 3942 3407 3943 3411
rect 3947 3407 3948 3411
rect 3942 3406 3948 3407
rect 3944 3367 3946 3406
rect 3943 3366 3947 3367
rect 3943 3361 3947 3362
rect 3944 3334 3946 3361
rect 3942 3333 3948 3334
rect 3942 3329 3943 3333
rect 3947 3329 3948 3333
rect 3942 3328 3948 3329
rect 3942 3316 3948 3317
rect 3942 3312 3943 3316
rect 3947 3312 3948 3316
rect 3942 3311 3948 3312
rect 3826 3295 3832 3296
rect 3826 3291 3827 3295
rect 3831 3291 3832 3295
rect 3826 3290 3832 3291
rect 3944 3287 3946 3311
rect 3255 3286 3259 3287
rect 3255 3281 3259 3282
rect 3327 3286 3331 3287
rect 3327 3281 3331 3282
rect 3383 3286 3387 3287
rect 3383 3281 3387 3282
rect 3479 3286 3483 3287
rect 3479 3281 3483 3282
rect 3503 3286 3507 3287
rect 3503 3281 3507 3282
rect 3623 3286 3627 3287
rect 3623 3281 3627 3282
rect 3631 3286 3635 3287
rect 3631 3281 3635 3282
rect 3743 3286 3747 3287
rect 3743 3281 3747 3282
rect 3783 3286 3787 3287
rect 3783 3281 3787 3282
rect 3839 3286 3843 3287
rect 3839 3281 3843 3282
rect 3943 3286 3947 3287
rect 3943 3281 3947 3282
rect 3256 3260 3258 3281
rect 3374 3279 3380 3280
rect 3374 3275 3375 3279
rect 3379 3275 3380 3279
rect 3374 3274 3380 3275
rect 3254 3259 3260 3260
rect 3254 3255 3255 3259
rect 3259 3255 3260 3259
rect 3254 3254 3260 3255
rect 2007 3249 2011 3250
rect 2490 3251 2496 3252
rect 1800 3228 1802 3249
rect 2008 3229 2010 3249
rect 2490 3247 2491 3251
rect 2495 3247 2496 3251
rect 2762 3251 2768 3252
rect 2490 3246 2496 3247
rect 2626 3247 2632 3248
rect 2046 3243 2052 3244
rect 2046 3239 2047 3243
rect 2051 3239 2052 3243
rect 2626 3243 2627 3247
rect 2631 3243 2632 3247
rect 2762 3247 2763 3251
rect 2767 3247 2768 3251
rect 2762 3246 2768 3247
rect 2906 3251 2912 3252
rect 2906 3247 2907 3251
rect 2911 3247 2912 3251
rect 2906 3246 2912 3247
rect 2926 3251 2932 3252
rect 2926 3247 2927 3251
rect 2931 3247 2932 3251
rect 2926 3246 2932 3247
rect 3194 3251 3200 3252
rect 3194 3247 3195 3251
rect 3199 3247 3200 3251
rect 3194 3246 3200 3247
rect 2626 3242 2632 3243
rect 2046 3238 2052 3239
rect 2414 3240 2420 3241
rect 2006 3228 2012 3229
rect 1798 3227 1804 3228
rect 1798 3223 1799 3227
rect 1803 3223 1804 3227
rect 2006 3224 2007 3228
rect 2011 3224 2012 3228
rect 2006 3223 2012 3224
rect 1798 3222 1804 3223
rect 1698 3219 1704 3220
rect 1698 3215 1699 3219
rect 1703 3215 1704 3219
rect 1698 3214 1704 3215
rect 1706 3219 1712 3220
rect 1706 3215 1707 3219
rect 1711 3215 1712 3219
rect 1706 3214 1712 3215
rect 2006 3211 2012 3212
rect 1798 3208 1804 3209
rect 1798 3204 1799 3208
rect 1803 3204 1804 3208
rect 2006 3207 2007 3211
rect 2011 3207 2012 3211
rect 2006 3206 2012 3207
rect 1798 3203 1804 3204
rect 1800 3171 1802 3203
rect 2008 3171 2010 3206
rect 2048 3199 2050 3238
rect 2414 3236 2415 3240
rect 2419 3236 2420 3240
rect 2414 3235 2420 3236
rect 2550 3240 2556 3241
rect 2550 3236 2551 3240
rect 2555 3236 2556 3240
rect 2550 3235 2556 3236
rect 2416 3199 2418 3235
rect 2552 3199 2554 3235
rect 2047 3198 2051 3199
rect 2047 3193 2051 3194
rect 2247 3198 2251 3199
rect 2247 3193 2251 3194
rect 2399 3198 2403 3199
rect 2399 3193 2403 3194
rect 2415 3198 2419 3199
rect 2415 3193 2419 3194
rect 2551 3198 2555 3199
rect 2551 3193 2555 3194
rect 2559 3198 2563 3199
rect 2559 3193 2563 3194
rect 1735 3170 1739 3171
rect 1735 3165 1739 3166
rect 1799 3170 1803 3171
rect 1799 3165 1803 3166
rect 2007 3170 2011 3171
rect 2048 3166 2050 3193
rect 2248 3169 2250 3193
rect 2400 3169 2402 3193
rect 2560 3169 2562 3193
rect 2246 3168 2252 3169
rect 2007 3165 2011 3166
rect 2046 3165 2052 3166
rect 1736 3141 1738 3165
rect 1734 3140 1740 3141
rect 1734 3136 1735 3140
rect 1739 3136 1740 3140
rect 2008 3138 2010 3165
rect 2046 3161 2047 3165
rect 2051 3161 2052 3165
rect 2246 3164 2247 3168
rect 2251 3164 2252 3168
rect 2246 3163 2252 3164
rect 2398 3168 2404 3169
rect 2398 3164 2399 3168
rect 2403 3164 2404 3168
rect 2398 3163 2404 3164
rect 2558 3168 2564 3169
rect 2558 3164 2559 3168
rect 2563 3164 2564 3168
rect 2558 3163 2564 3164
rect 2046 3160 2052 3161
rect 2322 3159 2328 3160
rect 2322 3155 2323 3159
rect 2327 3155 2328 3159
rect 2322 3154 2328 3155
rect 2330 3159 2336 3160
rect 2330 3155 2331 3159
rect 2335 3155 2336 3159
rect 2330 3154 2336 3155
rect 2246 3149 2252 3150
rect 2046 3148 2052 3149
rect 2046 3144 2047 3148
rect 2051 3144 2052 3148
rect 2246 3145 2247 3149
rect 2251 3145 2252 3149
rect 2246 3144 2252 3145
rect 2046 3143 2052 3144
rect 1734 3135 1740 3136
rect 2006 3137 2012 3138
rect 2006 3133 2007 3137
rect 2011 3133 2012 3137
rect 2006 3132 2012 3133
rect 1650 3131 1656 3132
rect 1650 3127 1651 3131
rect 1655 3127 1656 3131
rect 1650 3126 1656 3127
rect 1658 3131 1664 3132
rect 1658 3127 1659 3131
rect 1663 3127 1664 3131
rect 1658 3126 1664 3127
rect 1574 3121 1580 3122
rect 1574 3117 1575 3121
rect 1579 3117 1580 3121
rect 1574 3116 1580 3117
rect 1522 3099 1528 3100
rect 1522 3095 1523 3099
rect 1527 3095 1528 3099
rect 1576 3095 1578 3116
rect 1660 3100 1662 3126
rect 1734 3121 1740 3122
rect 1734 3117 1735 3121
rect 1739 3117 1740 3121
rect 1734 3116 1740 3117
rect 2006 3120 2012 3121
rect 2006 3116 2007 3120
rect 2011 3116 2012 3120
rect 2048 3119 2050 3143
rect 2248 3119 2250 3144
rect 1658 3099 1664 3100
rect 1658 3095 1659 3099
rect 1663 3095 1664 3099
rect 1736 3095 1738 3116
rect 2006 3115 2012 3116
rect 2047 3118 2051 3119
rect 1842 3099 1848 3100
rect 1842 3095 1843 3099
rect 1847 3095 1848 3099
rect 2008 3095 2010 3115
rect 2047 3113 2051 3114
rect 2079 3118 2083 3119
rect 2079 3113 2083 3114
rect 2223 3118 2227 3119
rect 2223 3113 2227 3114
rect 2247 3118 2251 3119
rect 2247 3113 2251 3114
rect 1186 3094 1192 3095
rect 1263 3094 1267 3095
rect 1263 3089 1267 3090
rect 1303 3094 1307 3095
rect 1346 3094 1352 3095
rect 1423 3094 1427 3095
rect 1303 3089 1307 3090
rect 1423 3089 1427 3090
rect 1455 3094 1459 3095
rect 1522 3094 1528 3095
rect 1575 3094 1579 3095
rect 1455 3089 1459 3090
rect 1575 3089 1579 3090
rect 1607 3094 1611 3095
rect 1658 3094 1664 3095
rect 1735 3094 1739 3095
rect 1607 3089 1611 3090
rect 1735 3089 1739 3090
rect 1767 3094 1771 3095
rect 1842 3094 1848 3095
rect 2007 3094 2011 3095
rect 1767 3089 1771 3090
rect 1178 3087 1184 3088
rect 1178 3083 1179 3087
rect 1183 3083 1184 3087
rect 1178 3082 1184 3083
rect 1218 3087 1224 3088
rect 1218 3083 1219 3087
rect 1223 3083 1224 3087
rect 1218 3082 1224 3083
rect 1142 3067 1148 3068
rect 1142 3063 1143 3067
rect 1147 3063 1148 3067
rect 1142 3062 1148 3063
rect 1220 3060 1222 3082
rect 1304 3068 1306 3089
rect 1378 3087 1384 3088
rect 1378 3083 1379 3087
rect 1383 3083 1384 3087
rect 1378 3082 1384 3083
rect 1302 3067 1308 3068
rect 1302 3063 1303 3067
rect 1307 3063 1308 3067
rect 1302 3062 1308 3063
rect 1380 3060 1382 3082
rect 1456 3068 1458 3089
rect 1530 3087 1536 3088
rect 1530 3083 1531 3087
rect 1535 3083 1536 3087
rect 1530 3082 1536 3083
rect 1454 3067 1460 3068
rect 1454 3063 1455 3067
rect 1459 3063 1460 3067
rect 1454 3062 1460 3063
rect 1532 3060 1534 3082
rect 1608 3068 1610 3089
rect 1682 3087 1688 3088
rect 1682 3083 1683 3087
rect 1687 3083 1688 3087
rect 1682 3082 1688 3083
rect 1606 3067 1612 3068
rect 1606 3063 1607 3067
rect 1611 3063 1612 3067
rect 1606 3062 1612 3063
rect 1684 3060 1686 3082
rect 1768 3068 1770 3089
rect 1766 3067 1772 3068
rect 1766 3063 1767 3067
rect 1771 3063 1772 3067
rect 1766 3062 1772 3063
rect 1844 3060 1846 3094
rect 2048 3093 2050 3113
rect 2007 3089 2011 3090
rect 2046 3092 2052 3093
rect 2080 3092 2082 3113
rect 2154 3111 2160 3112
rect 2154 3107 2155 3111
rect 2159 3107 2160 3111
rect 2154 3106 2160 3107
rect 2008 3069 2010 3089
rect 2046 3088 2047 3092
rect 2051 3088 2052 3092
rect 2046 3087 2052 3088
rect 2078 3091 2084 3092
rect 2078 3087 2079 3091
rect 2083 3087 2084 3091
rect 2078 3086 2084 3087
rect 2156 3084 2158 3106
rect 2224 3092 2226 3113
rect 2324 3112 2326 3154
rect 2332 3128 2334 3154
rect 2398 3149 2404 3150
rect 2398 3145 2399 3149
rect 2403 3145 2404 3149
rect 2398 3144 2404 3145
rect 2558 3149 2564 3150
rect 2558 3145 2559 3149
rect 2563 3145 2564 3149
rect 2558 3144 2564 3145
rect 2330 3127 2336 3128
rect 2330 3123 2331 3127
rect 2335 3123 2336 3127
rect 2330 3122 2336 3123
rect 2400 3119 2402 3144
rect 2560 3119 2562 3144
rect 2628 3128 2630 3242
rect 2686 3240 2692 3241
rect 2686 3236 2687 3240
rect 2691 3236 2692 3240
rect 2686 3235 2692 3236
rect 2830 3240 2836 3241
rect 2830 3236 2831 3240
rect 2835 3236 2836 3240
rect 2830 3235 2836 3236
rect 2974 3240 2980 3241
rect 2974 3236 2975 3240
rect 2979 3236 2980 3240
rect 2974 3235 2980 3236
rect 3118 3240 3124 3241
rect 3118 3236 3119 3240
rect 3123 3236 3124 3240
rect 3118 3235 3124 3236
rect 3254 3240 3260 3241
rect 3254 3236 3255 3240
rect 3259 3236 3260 3240
rect 3254 3235 3260 3236
rect 2688 3199 2690 3235
rect 2832 3199 2834 3235
rect 2976 3199 2978 3235
rect 3120 3199 3122 3235
rect 3256 3199 3258 3235
rect 2687 3198 2691 3199
rect 2687 3193 2691 3194
rect 2727 3198 2731 3199
rect 2727 3193 2731 3194
rect 2831 3198 2835 3199
rect 2831 3193 2835 3194
rect 2903 3198 2907 3199
rect 2903 3193 2907 3194
rect 2975 3198 2979 3199
rect 2975 3193 2979 3194
rect 3079 3198 3083 3199
rect 3079 3193 3083 3194
rect 3119 3198 3123 3199
rect 3119 3193 3123 3194
rect 3255 3198 3259 3199
rect 3255 3193 3259 3194
rect 3263 3198 3267 3199
rect 3263 3193 3267 3194
rect 2728 3169 2730 3193
rect 2904 3169 2906 3193
rect 3080 3169 3082 3193
rect 3264 3169 3266 3193
rect 3376 3176 3378 3274
rect 3384 3260 3386 3281
rect 3494 3279 3500 3280
rect 3494 3275 3495 3279
rect 3499 3275 3500 3279
rect 3494 3274 3500 3275
rect 3382 3259 3388 3260
rect 3382 3255 3383 3259
rect 3387 3255 3388 3259
rect 3382 3254 3388 3255
rect 3496 3252 3498 3274
rect 3504 3260 3506 3281
rect 3578 3279 3584 3280
rect 3578 3275 3579 3279
rect 3583 3275 3584 3279
rect 3578 3274 3584 3275
rect 3502 3259 3508 3260
rect 3502 3255 3503 3259
rect 3507 3255 3508 3259
rect 3502 3254 3508 3255
rect 3580 3252 3582 3274
rect 3624 3260 3626 3281
rect 3698 3279 3704 3280
rect 3698 3275 3699 3279
rect 3703 3275 3704 3279
rect 3698 3274 3704 3275
rect 3622 3259 3628 3260
rect 3622 3255 3623 3259
rect 3627 3255 3628 3259
rect 3622 3254 3628 3255
rect 3700 3252 3702 3274
rect 3744 3260 3746 3281
rect 3818 3279 3824 3280
rect 3818 3275 3819 3279
rect 3823 3275 3824 3279
rect 3818 3274 3824 3275
rect 3742 3259 3748 3260
rect 3742 3255 3743 3259
rect 3747 3255 3748 3259
rect 3742 3254 3748 3255
rect 3820 3252 3822 3274
rect 3840 3260 3842 3281
rect 3944 3261 3946 3281
rect 3942 3260 3948 3261
rect 3838 3259 3844 3260
rect 3838 3255 3839 3259
rect 3843 3255 3844 3259
rect 3942 3256 3943 3260
rect 3947 3256 3948 3260
rect 3942 3255 3948 3256
rect 3838 3254 3844 3255
rect 3494 3251 3500 3252
rect 3494 3247 3495 3251
rect 3499 3247 3500 3251
rect 3494 3246 3500 3247
rect 3578 3251 3584 3252
rect 3578 3247 3579 3251
rect 3583 3247 3584 3251
rect 3578 3246 3584 3247
rect 3698 3251 3704 3252
rect 3698 3247 3699 3251
rect 3703 3247 3704 3251
rect 3698 3246 3704 3247
rect 3818 3251 3824 3252
rect 3818 3247 3819 3251
rect 3823 3247 3824 3251
rect 3818 3246 3824 3247
rect 3914 3247 3920 3248
rect 3914 3243 3915 3247
rect 3919 3243 3920 3247
rect 3914 3242 3920 3243
rect 3942 3243 3948 3244
rect 3382 3240 3388 3241
rect 3382 3236 3383 3240
rect 3387 3236 3388 3240
rect 3382 3235 3388 3236
rect 3502 3240 3508 3241
rect 3502 3236 3503 3240
rect 3507 3236 3508 3240
rect 3502 3235 3508 3236
rect 3622 3240 3628 3241
rect 3622 3236 3623 3240
rect 3627 3236 3628 3240
rect 3622 3235 3628 3236
rect 3742 3240 3748 3241
rect 3742 3236 3743 3240
rect 3747 3236 3748 3240
rect 3742 3235 3748 3236
rect 3838 3240 3844 3241
rect 3838 3236 3839 3240
rect 3843 3236 3844 3240
rect 3838 3235 3844 3236
rect 3384 3199 3386 3235
rect 3504 3199 3506 3235
rect 3624 3199 3626 3235
rect 3744 3199 3746 3235
rect 3840 3199 3842 3235
rect 3383 3198 3387 3199
rect 3383 3193 3387 3194
rect 3447 3198 3451 3199
rect 3447 3193 3451 3194
rect 3503 3198 3507 3199
rect 3503 3193 3507 3194
rect 3623 3198 3627 3199
rect 3623 3193 3627 3194
rect 3631 3198 3635 3199
rect 3631 3193 3635 3194
rect 3743 3198 3747 3199
rect 3743 3193 3747 3194
rect 3815 3198 3819 3199
rect 3815 3193 3819 3194
rect 3839 3198 3843 3199
rect 3839 3193 3843 3194
rect 3374 3175 3380 3176
rect 3374 3171 3375 3175
rect 3379 3171 3380 3175
rect 3374 3170 3380 3171
rect 3448 3169 3450 3193
rect 3632 3169 3634 3193
rect 3816 3169 3818 3193
rect 2726 3168 2732 3169
rect 2726 3164 2727 3168
rect 2731 3164 2732 3168
rect 2726 3163 2732 3164
rect 2902 3168 2908 3169
rect 2902 3164 2903 3168
rect 2907 3164 2908 3168
rect 2902 3163 2908 3164
rect 3078 3168 3084 3169
rect 3078 3164 3079 3168
rect 3083 3164 3084 3168
rect 3078 3163 3084 3164
rect 3262 3168 3268 3169
rect 3262 3164 3263 3168
rect 3267 3164 3268 3168
rect 3262 3163 3268 3164
rect 3446 3168 3452 3169
rect 3446 3164 3447 3168
rect 3451 3164 3452 3168
rect 3446 3163 3452 3164
rect 3630 3168 3636 3169
rect 3630 3164 3631 3168
rect 3635 3164 3636 3168
rect 3630 3163 3636 3164
rect 3814 3168 3820 3169
rect 3814 3164 3815 3168
rect 3819 3164 3820 3168
rect 3814 3163 3820 3164
rect 2634 3159 2640 3160
rect 2634 3155 2635 3159
rect 2639 3155 2640 3159
rect 2634 3154 2640 3155
rect 2802 3159 2808 3160
rect 2802 3155 2803 3159
rect 2807 3155 2808 3159
rect 2802 3154 2808 3155
rect 3154 3159 3160 3160
rect 3154 3155 3155 3159
rect 3159 3155 3160 3159
rect 3154 3154 3160 3155
rect 3338 3159 3344 3160
rect 3338 3155 3339 3159
rect 3343 3155 3344 3159
rect 3338 3154 3344 3155
rect 3522 3159 3528 3160
rect 3522 3155 3523 3159
rect 3527 3155 3528 3159
rect 3522 3154 3528 3155
rect 3890 3159 3896 3160
rect 3890 3155 3891 3159
rect 3895 3155 3896 3159
rect 3890 3154 3896 3155
rect 2636 3128 2638 3154
rect 2726 3149 2732 3150
rect 2726 3145 2727 3149
rect 2731 3145 2732 3149
rect 2726 3144 2732 3145
rect 2626 3127 2632 3128
rect 2626 3123 2627 3127
rect 2631 3123 2632 3127
rect 2626 3122 2632 3123
rect 2634 3127 2640 3128
rect 2634 3123 2635 3127
rect 2639 3123 2640 3127
rect 2634 3122 2640 3123
rect 2728 3119 2730 3144
rect 2804 3128 2806 3154
rect 2902 3149 2908 3150
rect 2902 3145 2903 3149
rect 2907 3145 2908 3149
rect 2902 3144 2908 3145
rect 3078 3149 3084 3150
rect 3078 3145 3079 3149
rect 3083 3145 3084 3149
rect 3078 3144 3084 3145
rect 2802 3127 2808 3128
rect 2802 3123 2803 3127
rect 2807 3123 2808 3127
rect 2802 3122 2808 3123
rect 2904 3119 2906 3144
rect 3080 3119 3082 3144
rect 3156 3128 3158 3154
rect 3262 3149 3268 3150
rect 3262 3145 3263 3149
rect 3267 3145 3268 3149
rect 3262 3144 3268 3145
rect 3154 3127 3160 3128
rect 3154 3123 3155 3127
rect 3159 3123 3160 3127
rect 3154 3122 3160 3123
rect 3264 3119 3266 3144
rect 3340 3128 3342 3154
rect 3446 3149 3452 3150
rect 3446 3145 3447 3149
rect 3451 3145 3452 3149
rect 3446 3144 3452 3145
rect 3338 3127 3344 3128
rect 3338 3123 3339 3127
rect 3343 3123 3344 3127
rect 3338 3122 3344 3123
rect 3448 3119 3450 3144
rect 3524 3128 3526 3154
rect 3630 3149 3636 3150
rect 3630 3145 3631 3149
rect 3635 3145 3636 3149
rect 3630 3144 3636 3145
rect 3814 3149 3820 3150
rect 3814 3145 3815 3149
rect 3819 3145 3820 3149
rect 3814 3144 3820 3145
rect 3522 3127 3528 3128
rect 3522 3123 3523 3127
rect 3527 3123 3528 3127
rect 3522 3122 3528 3123
rect 3602 3119 3608 3120
rect 3632 3119 3634 3144
rect 3816 3119 3818 3144
rect 2375 3118 2379 3119
rect 2375 3113 2379 3114
rect 2399 3118 2403 3119
rect 2399 3113 2403 3114
rect 2527 3118 2531 3119
rect 2527 3113 2531 3114
rect 2559 3118 2563 3119
rect 2559 3113 2563 3114
rect 2687 3118 2691 3119
rect 2687 3113 2691 3114
rect 2727 3118 2731 3119
rect 2727 3113 2731 3114
rect 2855 3118 2859 3119
rect 2855 3113 2859 3114
rect 2903 3118 2907 3119
rect 2903 3113 2907 3114
rect 3039 3118 3043 3119
rect 3039 3113 3043 3114
rect 3079 3118 3083 3119
rect 3079 3113 3083 3114
rect 3231 3118 3235 3119
rect 3231 3113 3235 3114
rect 3263 3118 3267 3119
rect 3263 3113 3267 3114
rect 3431 3118 3435 3119
rect 3431 3113 3435 3114
rect 3447 3118 3451 3119
rect 3602 3115 3603 3119
rect 3607 3115 3608 3119
rect 3602 3114 3608 3115
rect 3631 3118 3635 3119
rect 3447 3113 3451 3114
rect 2322 3111 2328 3112
rect 2322 3107 2323 3111
rect 2327 3107 2328 3111
rect 2322 3106 2328 3107
rect 2376 3092 2378 3113
rect 2450 3111 2456 3112
rect 2450 3107 2451 3111
rect 2455 3107 2456 3111
rect 2450 3106 2456 3107
rect 2222 3091 2228 3092
rect 2222 3087 2223 3091
rect 2227 3087 2228 3091
rect 2222 3086 2228 3087
rect 2374 3091 2380 3092
rect 2374 3087 2375 3091
rect 2379 3087 2380 3091
rect 2374 3086 2380 3087
rect 2452 3084 2454 3106
rect 2528 3092 2530 3113
rect 2602 3111 2608 3112
rect 2602 3107 2603 3111
rect 2607 3107 2608 3111
rect 2602 3106 2608 3107
rect 2526 3091 2532 3092
rect 2526 3087 2527 3091
rect 2531 3087 2532 3091
rect 2526 3086 2532 3087
rect 2604 3084 2606 3106
rect 2658 3103 2664 3104
rect 2658 3099 2659 3103
rect 2663 3099 2664 3103
rect 2658 3098 2664 3099
rect 2660 3084 2662 3098
rect 2688 3092 2690 3113
rect 2856 3092 2858 3113
rect 2922 3111 2928 3112
rect 2922 3107 2923 3111
rect 2927 3107 2928 3111
rect 2922 3106 2928 3107
rect 2930 3111 2936 3112
rect 2930 3107 2931 3111
rect 2935 3107 2936 3111
rect 2930 3106 2936 3107
rect 2686 3091 2692 3092
rect 2686 3087 2687 3091
rect 2691 3087 2692 3091
rect 2686 3086 2692 3087
rect 2854 3091 2860 3092
rect 2854 3087 2855 3091
rect 2859 3087 2860 3091
rect 2854 3086 2860 3087
rect 2154 3083 2160 3084
rect 2154 3079 2155 3083
rect 2159 3079 2160 3083
rect 2450 3083 2456 3084
rect 2154 3078 2160 3079
rect 2298 3079 2304 3080
rect 2046 3075 2052 3076
rect 2046 3071 2047 3075
rect 2051 3071 2052 3075
rect 2298 3075 2299 3079
rect 2303 3075 2304 3079
rect 2450 3079 2451 3083
rect 2455 3079 2456 3083
rect 2450 3078 2456 3079
rect 2602 3083 2608 3084
rect 2602 3079 2603 3083
rect 2607 3079 2608 3083
rect 2602 3078 2608 3079
rect 2658 3083 2664 3084
rect 2658 3079 2659 3083
rect 2663 3079 2664 3083
rect 2658 3078 2664 3079
rect 2298 3074 2304 3075
rect 2046 3070 2052 3071
rect 2078 3072 2084 3073
rect 2006 3068 2012 3069
rect 2006 3064 2007 3068
rect 2011 3064 2012 3068
rect 2006 3063 2012 3064
rect 874 3059 880 3060
rect 874 3055 875 3059
rect 879 3055 880 3059
rect 874 3054 880 3055
rect 1050 3059 1056 3060
rect 1050 3055 1051 3059
rect 1055 3055 1056 3059
rect 1050 3054 1056 3055
rect 1218 3059 1224 3060
rect 1218 3055 1219 3059
rect 1223 3055 1224 3059
rect 1218 3054 1224 3055
rect 1378 3059 1384 3060
rect 1378 3055 1379 3059
rect 1383 3055 1384 3059
rect 1378 3054 1384 3055
rect 1530 3059 1536 3060
rect 1530 3055 1531 3059
rect 1535 3055 1536 3059
rect 1530 3054 1536 3055
rect 1682 3059 1688 3060
rect 1682 3055 1683 3059
rect 1687 3055 1688 3059
rect 1682 3054 1688 3055
rect 1842 3059 1848 3060
rect 1842 3055 1843 3059
rect 1847 3055 1848 3059
rect 1842 3054 1848 3055
rect 2006 3051 2012 3052
rect 974 3048 980 3049
rect 974 3044 975 3048
rect 979 3044 980 3048
rect 974 3043 980 3044
rect 1142 3048 1148 3049
rect 1142 3044 1143 3048
rect 1147 3044 1148 3048
rect 1142 3043 1148 3044
rect 1302 3048 1308 3049
rect 1302 3044 1303 3048
rect 1307 3044 1308 3048
rect 1302 3043 1308 3044
rect 1454 3048 1460 3049
rect 1454 3044 1455 3048
rect 1459 3044 1460 3048
rect 1454 3043 1460 3044
rect 1606 3048 1612 3049
rect 1606 3044 1607 3048
rect 1611 3044 1612 3048
rect 1606 3043 1612 3044
rect 1766 3048 1772 3049
rect 1766 3044 1767 3048
rect 1771 3044 1772 3048
rect 2006 3047 2007 3051
rect 2011 3047 2012 3051
rect 2006 3046 2012 3047
rect 1766 3043 1772 3044
rect 976 2995 978 3043
rect 1144 2995 1146 3043
rect 1304 2995 1306 3043
rect 1456 2995 1458 3043
rect 1608 2995 1610 3043
rect 1768 2995 1770 3043
rect 2008 2995 2010 3046
rect 2048 3035 2050 3070
rect 2078 3068 2079 3072
rect 2083 3068 2084 3072
rect 2078 3067 2084 3068
rect 2222 3072 2228 3073
rect 2222 3068 2223 3072
rect 2227 3068 2228 3072
rect 2222 3067 2228 3068
rect 2080 3035 2082 3067
rect 2224 3035 2226 3067
rect 2047 3034 2051 3035
rect 2047 3029 2051 3030
rect 2071 3034 2075 3035
rect 2071 3029 2075 3030
rect 2079 3034 2083 3035
rect 2079 3029 2083 3030
rect 2183 3034 2187 3035
rect 2183 3029 2187 3030
rect 2223 3034 2227 3035
rect 2223 3029 2227 3030
rect 2048 3002 2050 3029
rect 2072 3005 2074 3029
rect 2184 3005 2186 3029
rect 2070 3004 2076 3005
rect 2046 3001 2052 3002
rect 2046 2997 2047 3001
rect 2051 2997 2052 3001
rect 2070 3000 2071 3004
rect 2075 3000 2076 3004
rect 2070 2999 2076 3000
rect 2182 3004 2188 3005
rect 2182 3000 2183 3004
rect 2187 3000 2188 3004
rect 2182 2999 2188 3000
rect 2046 2996 2052 2997
rect 2138 2995 2144 2996
rect 935 2994 939 2995
rect 935 2989 939 2990
rect 975 2994 979 2995
rect 975 2989 979 2990
rect 1103 2994 1107 2995
rect 1103 2989 1107 2990
rect 1143 2994 1147 2995
rect 1143 2989 1147 2990
rect 1295 2994 1299 2995
rect 1295 2989 1299 2990
rect 1303 2994 1307 2995
rect 1303 2989 1307 2990
rect 1455 2994 1459 2995
rect 1455 2989 1459 2990
rect 1495 2994 1499 2995
rect 1495 2989 1499 2990
rect 1607 2994 1611 2995
rect 1607 2989 1611 2990
rect 1711 2994 1715 2995
rect 1711 2989 1715 2990
rect 1767 2994 1771 2995
rect 1767 2989 1771 2990
rect 1903 2994 1907 2995
rect 1903 2989 1907 2990
rect 2007 2994 2011 2995
rect 2138 2991 2139 2995
rect 2143 2991 2144 2995
rect 2138 2990 2144 2991
rect 2154 2995 2160 2996
rect 2154 2991 2155 2995
rect 2159 2991 2160 2995
rect 2154 2990 2160 2991
rect 2007 2989 2011 2990
rect 936 2965 938 2989
rect 1104 2965 1106 2989
rect 1296 2965 1298 2989
rect 1496 2965 1498 2989
rect 1712 2965 1714 2989
rect 1904 2965 1906 2989
rect 934 2964 940 2965
rect 934 2960 935 2964
rect 939 2960 940 2964
rect 934 2959 940 2960
rect 1102 2964 1108 2965
rect 1102 2960 1103 2964
rect 1107 2960 1108 2964
rect 1102 2959 1108 2960
rect 1294 2964 1300 2965
rect 1294 2960 1295 2964
rect 1299 2960 1300 2964
rect 1294 2959 1300 2960
rect 1494 2964 1500 2965
rect 1494 2960 1495 2964
rect 1499 2960 1500 2964
rect 1494 2959 1500 2960
rect 1710 2964 1716 2965
rect 1710 2960 1711 2964
rect 1715 2960 1716 2964
rect 1710 2959 1716 2960
rect 1902 2964 1908 2965
rect 1902 2960 1903 2964
rect 1907 2960 1908 2964
rect 2008 2962 2010 2989
rect 2070 2985 2076 2986
rect 2046 2984 2052 2985
rect 2046 2980 2047 2984
rect 2051 2980 2052 2984
rect 2070 2981 2071 2985
rect 2075 2981 2076 2985
rect 2070 2980 2076 2981
rect 2046 2979 2052 2980
rect 1902 2959 1908 2960
rect 2006 2961 2012 2962
rect 2006 2957 2007 2961
rect 2011 2957 2012 2961
rect 2006 2956 2012 2957
rect 730 2955 736 2956
rect 730 2951 731 2955
rect 735 2951 736 2955
rect 730 2950 736 2951
rect 858 2955 864 2956
rect 858 2951 859 2955
rect 863 2951 864 2955
rect 858 2950 864 2951
rect 1010 2955 1016 2956
rect 1010 2951 1011 2955
rect 1015 2951 1016 2955
rect 1010 2950 1016 2951
rect 1178 2955 1184 2956
rect 1178 2951 1179 2955
rect 1183 2951 1184 2955
rect 1178 2950 1184 2951
rect 1370 2955 1376 2956
rect 1370 2951 1371 2955
rect 1375 2951 1376 2955
rect 1370 2950 1376 2951
rect 1570 2955 1576 2956
rect 1570 2951 1571 2955
rect 1575 2951 1576 2955
rect 1570 2950 1576 2951
rect 1786 2955 1792 2956
rect 1786 2951 1787 2955
rect 1791 2951 1792 2955
rect 1786 2950 1792 2951
rect 1794 2955 1800 2956
rect 2048 2955 2050 2979
rect 2072 2955 2074 2980
rect 1794 2951 1795 2955
rect 1799 2951 1800 2955
rect 1794 2950 1800 2951
rect 2047 2954 2051 2955
rect 542 2945 548 2946
rect 542 2941 543 2945
rect 547 2941 548 2945
rect 542 2940 548 2941
rect 654 2945 660 2946
rect 654 2941 655 2945
rect 659 2941 660 2945
rect 654 2940 660 2941
rect 514 2923 520 2924
rect 514 2919 515 2923
rect 519 2919 520 2923
rect 544 2919 546 2940
rect 642 2923 648 2924
rect 642 2919 643 2923
rect 647 2919 648 2923
rect 656 2919 658 2940
rect 732 2924 734 2950
rect 782 2945 788 2946
rect 782 2941 783 2945
rect 787 2941 788 2945
rect 782 2940 788 2941
rect 934 2945 940 2946
rect 934 2941 935 2945
rect 939 2941 940 2945
rect 934 2940 940 2941
rect 730 2923 736 2924
rect 730 2919 731 2923
rect 735 2919 736 2923
rect 784 2919 786 2940
rect 936 2919 938 2940
rect 1012 2924 1014 2950
rect 1102 2945 1108 2946
rect 1102 2941 1103 2945
rect 1107 2941 1108 2945
rect 1102 2940 1108 2941
rect 990 2923 996 2924
rect 990 2919 991 2923
rect 995 2919 996 2923
rect 1010 2923 1016 2924
rect 1010 2919 1011 2923
rect 1015 2919 1016 2923
rect 1104 2919 1106 2940
rect 1180 2924 1182 2950
rect 1294 2945 1300 2946
rect 1294 2941 1295 2945
rect 1299 2941 1300 2945
rect 1294 2940 1300 2941
rect 1178 2923 1184 2924
rect 1178 2919 1179 2923
rect 1183 2919 1184 2923
rect 1296 2919 1298 2940
rect 1372 2924 1374 2950
rect 1494 2945 1500 2946
rect 1494 2941 1495 2945
rect 1499 2941 1500 2945
rect 1494 2940 1500 2941
rect 1370 2923 1376 2924
rect 1370 2919 1371 2923
rect 1375 2919 1376 2923
rect 1496 2919 1498 2940
rect 327 2918 331 2919
rect 327 2913 331 2914
rect 343 2918 347 2919
rect 426 2918 432 2919
rect 439 2918 443 2919
rect 343 2913 347 2914
rect 439 2913 443 2914
rect 447 2918 451 2919
rect 514 2918 520 2919
rect 543 2918 547 2919
rect 447 2913 451 2914
rect 543 2913 547 2914
rect 575 2918 579 2919
rect 642 2918 648 2919
rect 655 2918 659 2919
rect 575 2913 579 2914
rect 274 2911 280 2912
rect 274 2907 275 2911
rect 279 2907 280 2911
rect 274 2906 280 2907
rect 282 2911 288 2912
rect 282 2907 283 2911
rect 287 2907 288 2911
rect 282 2906 288 2907
rect 110 2888 111 2892
rect 115 2888 116 2892
rect 110 2887 116 2888
rect 206 2891 212 2892
rect 206 2887 207 2891
rect 211 2887 212 2891
rect 206 2886 212 2887
rect 284 2884 286 2906
rect 328 2892 330 2913
rect 402 2911 408 2912
rect 402 2907 403 2911
rect 407 2907 408 2911
rect 402 2906 408 2907
rect 326 2891 332 2892
rect 326 2887 327 2891
rect 331 2887 332 2891
rect 326 2886 332 2887
rect 404 2884 406 2906
rect 448 2892 450 2913
rect 576 2892 578 2913
rect 446 2891 452 2892
rect 446 2887 447 2891
rect 451 2887 452 2891
rect 446 2886 452 2887
rect 574 2891 580 2892
rect 574 2887 575 2891
rect 579 2887 580 2891
rect 644 2888 646 2918
rect 655 2913 659 2914
rect 703 2918 707 2919
rect 730 2918 736 2919
rect 783 2918 787 2919
rect 703 2913 707 2914
rect 783 2913 787 2914
rect 847 2918 851 2919
rect 847 2913 851 2914
rect 935 2918 939 2919
rect 990 2918 996 2919
rect 999 2918 1003 2919
rect 1010 2918 1016 2919
rect 1103 2918 1107 2919
rect 935 2913 939 2914
rect 704 2892 706 2913
rect 770 2911 776 2912
rect 770 2907 771 2911
rect 775 2907 776 2911
rect 770 2906 776 2907
rect 702 2891 708 2892
rect 574 2886 580 2887
rect 642 2887 648 2888
rect 282 2883 288 2884
rect 282 2879 283 2883
rect 287 2879 288 2883
rect 282 2878 288 2879
rect 402 2883 408 2884
rect 402 2879 403 2883
rect 407 2879 408 2883
rect 642 2883 643 2887
rect 647 2883 648 2887
rect 702 2887 703 2891
rect 707 2887 708 2891
rect 702 2886 708 2887
rect 642 2882 648 2883
rect 402 2878 408 2879
rect 522 2879 528 2880
rect 110 2875 116 2876
rect 110 2871 111 2875
rect 115 2871 116 2875
rect 522 2875 523 2879
rect 527 2875 528 2879
rect 522 2874 528 2875
rect 110 2870 116 2871
rect 206 2872 212 2873
rect 112 2839 114 2870
rect 206 2868 207 2872
rect 211 2868 212 2872
rect 206 2867 212 2868
rect 326 2872 332 2873
rect 326 2868 327 2872
rect 331 2868 332 2872
rect 326 2867 332 2868
rect 446 2872 452 2873
rect 446 2868 447 2872
rect 451 2868 452 2872
rect 446 2867 452 2868
rect 208 2839 210 2867
rect 328 2839 330 2867
rect 448 2839 450 2867
rect 111 2838 115 2839
rect 111 2833 115 2834
rect 135 2838 139 2839
rect 135 2833 139 2834
rect 207 2838 211 2839
rect 207 2833 211 2834
rect 247 2838 251 2839
rect 247 2833 251 2834
rect 327 2838 331 2839
rect 327 2833 331 2834
rect 399 2838 403 2839
rect 399 2833 403 2834
rect 447 2838 451 2839
rect 447 2833 451 2834
rect 112 2806 114 2833
rect 136 2809 138 2833
rect 248 2809 250 2833
rect 400 2809 402 2833
rect 134 2808 140 2809
rect 110 2805 116 2806
rect 110 2801 111 2805
rect 115 2801 116 2805
rect 134 2804 135 2808
rect 139 2804 140 2808
rect 134 2803 140 2804
rect 246 2808 252 2809
rect 246 2804 247 2808
rect 251 2804 252 2808
rect 246 2803 252 2804
rect 398 2808 404 2809
rect 398 2804 399 2808
rect 403 2804 404 2808
rect 398 2803 404 2804
rect 110 2800 116 2801
rect 202 2799 208 2800
rect 202 2795 203 2799
rect 207 2795 208 2799
rect 202 2794 208 2795
rect 218 2799 224 2800
rect 218 2795 219 2799
rect 223 2795 224 2799
rect 218 2794 224 2795
rect 378 2799 384 2800
rect 378 2795 379 2799
rect 383 2795 384 2799
rect 378 2794 384 2795
rect 134 2789 140 2790
rect 110 2788 116 2789
rect 110 2784 111 2788
rect 115 2784 116 2788
rect 134 2785 135 2789
rect 139 2785 140 2789
rect 134 2784 140 2785
rect 110 2783 116 2784
rect 112 2755 114 2783
rect 136 2755 138 2784
rect 111 2754 115 2755
rect 111 2749 115 2750
rect 135 2754 139 2755
rect 135 2749 139 2750
rect 112 2729 114 2749
rect 110 2728 116 2729
rect 136 2728 138 2749
rect 204 2748 206 2794
rect 220 2768 222 2794
rect 246 2789 252 2790
rect 246 2785 247 2789
rect 251 2785 252 2789
rect 246 2784 252 2785
rect 218 2767 224 2768
rect 218 2763 219 2767
rect 223 2763 224 2767
rect 218 2762 224 2763
rect 248 2755 250 2784
rect 380 2768 382 2794
rect 398 2789 404 2790
rect 398 2785 399 2789
rect 403 2785 404 2789
rect 398 2784 404 2785
rect 378 2767 384 2768
rect 378 2763 379 2767
rect 383 2763 384 2767
rect 378 2762 384 2763
rect 400 2755 402 2784
rect 524 2768 526 2874
rect 574 2872 580 2873
rect 574 2868 575 2872
rect 579 2868 580 2872
rect 574 2867 580 2868
rect 702 2872 708 2873
rect 702 2868 703 2872
rect 707 2868 708 2872
rect 702 2867 708 2868
rect 576 2839 578 2867
rect 704 2839 706 2867
rect 551 2838 555 2839
rect 551 2833 555 2834
rect 575 2838 579 2839
rect 575 2833 579 2834
rect 703 2838 707 2839
rect 703 2833 707 2834
rect 711 2838 715 2839
rect 711 2833 715 2834
rect 772 2833 774 2906
rect 848 2892 850 2913
rect 946 2911 952 2912
rect 946 2907 947 2911
rect 951 2907 952 2911
rect 946 2906 952 2907
rect 974 2911 980 2912
rect 974 2907 975 2911
rect 979 2907 980 2911
rect 974 2906 980 2907
rect 846 2891 852 2892
rect 846 2887 847 2891
rect 851 2887 852 2891
rect 846 2886 852 2887
rect 846 2872 852 2873
rect 846 2868 847 2872
rect 851 2868 852 2872
rect 846 2867 852 2868
rect 848 2839 850 2867
rect 847 2838 851 2839
rect 847 2833 851 2834
rect 879 2838 883 2839
rect 879 2833 883 2834
rect 552 2809 554 2833
rect 712 2809 714 2833
rect 772 2831 782 2833
rect 550 2808 556 2809
rect 550 2804 551 2808
rect 555 2804 556 2808
rect 550 2803 556 2804
rect 710 2808 716 2809
rect 710 2804 711 2808
rect 715 2804 716 2808
rect 710 2803 716 2804
rect 780 2800 782 2831
rect 880 2809 882 2833
rect 878 2808 884 2809
rect 878 2804 879 2808
rect 883 2804 884 2808
rect 878 2803 884 2804
rect 948 2800 950 2906
rect 976 2884 978 2906
rect 992 2884 994 2918
rect 999 2913 1003 2914
rect 1103 2913 1107 2914
rect 1167 2918 1171 2919
rect 1178 2918 1184 2919
rect 1295 2918 1299 2919
rect 1167 2913 1171 2914
rect 1295 2913 1299 2914
rect 1351 2918 1355 2919
rect 1370 2918 1376 2919
rect 1495 2918 1499 2919
rect 1351 2913 1355 2914
rect 1495 2913 1499 2914
rect 1535 2918 1539 2919
rect 1535 2913 1539 2914
rect 1000 2892 1002 2913
rect 1168 2892 1170 2913
rect 1250 2911 1256 2912
rect 1250 2907 1251 2911
rect 1255 2907 1256 2911
rect 1250 2906 1256 2907
rect 998 2891 1004 2892
rect 998 2887 999 2891
rect 1003 2887 1004 2891
rect 998 2886 1004 2887
rect 1166 2891 1172 2892
rect 1166 2887 1167 2891
rect 1171 2887 1172 2891
rect 1166 2886 1172 2887
rect 1252 2884 1254 2906
rect 1352 2892 1354 2913
rect 1438 2911 1444 2912
rect 1438 2907 1439 2911
rect 1443 2907 1444 2911
rect 1438 2906 1444 2907
rect 1350 2891 1356 2892
rect 1350 2887 1351 2891
rect 1355 2887 1356 2891
rect 1350 2886 1356 2887
rect 1440 2884 1442 2906
rect 1536 2892 1538 2913
rect 1572 2912 1574 2950
rect 1710 2945 1716 2946
rect 1710 2941 1711 2945
rect 1715 2941 1716 2945
rect 1710 2940 1716 2941
rect 1712 2919 1714 2940
rect 1711 2918 1715 2919
rect 1711 2913 1715 2914
rect 1727 2918 1731 2919
rect 1727 2913 1731 2914
rect 1570 2911 1576 2912
rect 1570 2907 1571 2911
rect 1575 2907 1576 2911
rect 1570 2906 1576 2907
rect 1728 2892 1730 2913
rect 1788 2912 1790 2950
rect 1796 2924 1798 2950
rect 2047 2949 2051 2950
rect 2071 2954 2075 2955
rect 2071 2949 2075 2950
rect 1902 2945 1908 2946
rect 1902 2941 1903 2945
rect 1907 2941 1908 2945
rect 1902 2940 1908 2941
rect 2006 2944 2012 2945
rect 2006 2940 2007 2944
rect 2011 2940 2012 2944
rect 1794 2923 1800 2924
rect 1794 2919 1795 2923
rect 1799 2919 1800 2923
rect 1904 2919 1906 2940
rect 2006 2939 2012 2940
rect 2008 2919 2010 2939
rect 2048 2929 2050 2949
rect 2046 2928 2052 2929
rect 2072 2928 2074 2949
rect 2140 2948 2142 2990
rect 2156 2964 2158 2990
rect 2182 2985 2188 2986
rect 2182 2981 2183 2985
rect 2187 2981 2188 2985
rect 2182 2980 2188 2981
rect 2154 2963 2160 2964
rect 2154 2959 2155 2963
rect 2159 2959 2160 2963
rect 2154 2958 2160 2959
rect 2184 2955 2186 2980
rect 2300 2964 2302 3074
rect 2374 3072 2380 3073
rect 2374 3068 2375 3072
rect 2379 3068 2380 3072
rect 2374 3067 2380 3068
rect 2526 3072 2532 3073
rect 2526 3068 2527 3072
rect 2531 3068 2532 3072
rect 2526 3067 2532 3068
rect 2686 3072 2692 3073
rect 2686 3068 2687 3072
rect 2691 3068 2692 3072
rect 2686 3067 2692 3068
rect 2854 3072 2860 3073
rect 2854 3068 2855 3072
rect 2859 3068 2860 3072
rect 2854 3067 2860 3068
rect 2376 3035 2378 3067
rect 2528 3035 2530 3067
rect 2688 3035 2690 3067
rect 2856 3035 2858 3067
rect 2327 3034 2331 3035
rect 2327 3029 2331 3030
rect 2375 3034 2379 3035
rect 2375 3029 2379 3030
rect 2479 3034 2483 3035
rect 2479 3029 2483 3030
rect 2527 3034 2531 3035
rect 2527 3029 2531 3030
rect 2655 3034 2659 3035
rect 2655 3029 2659 3030
rect 2687 3034 2691 3035
rect 2687 3029 2691 3030
rect 2855 3034 2859 3035
rect 2855 3029 2859 3030
rect 2328 3005 2330 3029
rect 2480 3005 2482 3029
rect 2656 3005 2658 3029
rect 2856 3005 2858 3029
rect 2924 3012 2926 3106
rect 2932 3084 2934 3106
rect 3040 3092 3042 3113
rect 3114 3111 3120 3112
rect 3114 3107 3115 3111
rect 3119 3107 3120 3111
rect 3114 3106 3120 3107
rect 3038 3091 3044 3092
rect 3038 3087 3039 3091
rect 3043 3087 3044 3091
rect 3038 3086 3044 3087
rect 3116 3084 3118 3106
rect 3232 3092 3234 3113
rect 3306 3111 3312 3112
rect 3306 3107 3307 3111
rect 3311 3107 3312 3111
rect 3306 3106 3312 3107
rect 3230 3091 3236 3092
rect 3230 3087 3231 3091
rect 3235 3087 3236 3091
rect 3230 3086 3236 3087
rect 3308 3084 3310 3106
rect 3432 3092 3434 3113
rect 3506 3111 3512 3112
rect 3506 3107 3507 3111
rect 3511 3107 3512 3111
rect 3506 3106 3512 3107
rect 3430 3091 3436 3092
rect 3430 3087 3431 3091
rect 3435 3087 3436 3091
rect 3430 3086 3436 3087
rect 3508 3084 3510 3106
rect 3604 3084 3606 3114
rect 3631 3113 3635 3114
rect 3639 3118 3643 3119
rect 3639 3113 3643 3114
rect 3815 3118 3819 3119
rect 3815 3113 3819 3114
rect 3839 3118 3843 3119
rect 3839 3113 3843 3114
rect 3640 3092 3642 3113
rect 3840 3092 3842 3113
rect 3892 3112 3894 3154
rect 3916 3128 3918 3242
rect 3942 3239 3943 3243
rect 3947 3239 3948 3243
rect 3942 3238 3948 3239
rect 3944 3199 3946 3238
rect 3943 3198 3947 3199
rect 3943 3193 3947 3194
rect 3944 3166 3946 3193
rect 3942 3165 3948 3166
rect 3942 3161 3943 3165
rect 3947 3161 3948 3165
rect 3942 3160 3948 3161
rect 3942 3148 3948 3149
rect 3942 3144 3943 3148
rect 3947 3144 3948 3148
rect 3942 3143 3948 3144
rect 3914 3127 3920 3128
rect 3914 3123 3915 3127
rect 3919 3123 3920 3127
rect 3914 3122 3920 3123
rect 3944 3119 3946 3143
rect 3943 3118 3947 3119
rect 3943 3113 3947 3114
rect 3890 3111 3896 3112
rect 3890 3107 3891 3111
rect 3895 3107 3896 3111
rect 3890 3106 3896 3107
rect 3944 3093 3946 3113
rect 3942 3092 3948 3093
rect 3638 3091 3644 3092
rect 3638 3087 3639 3091
rect 3643 3087 3644 3091
rect 3638 3086 3644 3087
rect 3838 3091 3844 3092
rect 3838 3087 3839 3091
rect 3843 3087 3844 3091
rect 3942 3088 3943 3092
rect 3947 3088 3948 3092
rect 3942 3087 3948 3088
rect 3838 3086 3844 3087
rect 2930 3083 2936 3084
rect 2930 3079 2931 3083
rect 2935 3079 2936 3083
rect 2930 3078 2936 3079
rect 3114 3083 3120 3084
rect 3114 3079 3115 3083
rect 3119 3079 3120 3083
rect 3114 3078 3120 3079
rect 3306 3083 3312 3084
rect 3306 3079 3307 3083
rect 3311 3079 3312 3083
rect 3306 3078 3312 3079
rect 3506 3083 3512 3084
rect 3506 3079 3507 3083
rect 3511 3079 3512 3083
rect 3506 3078 3512 3079
rect 3602 3083 3608 3084
rect 3602 3079 3603 3083
rect 3607 3079 3608 3083
rect 3602 3078 3608 3079
rect 3914 3079 3920 3080
rect 3914 3075 3915 3079
rect 3919 3075 3920 3079
rect 3914 3074 3920 3075
rect 3942 3075 3948 3076
rect 3038 3072 3044 3073
rect 3038 3068 3039 3072
rect 3043 3068 3044 3072
rect 3038 3067 3044 3068
rect 3230 3072 3236 3073
rect 3230 3068 3231 3072
rect 3235 3068 3236 3072
rect 3230 3067 3236 3068
rect 3430 3072 3436 3073
rect 3430 3068 3431 3072
rect 3435 3068 3436 3072
rect 3430 3067 3436 3068
rect 3638 3072 3644 3073
rect 3638 3068 3639 3072
rect 3643 3068 3644 3072
rect 3638 3067 3644 3068
rect 3838 3072 3844 3073
rect 3838 3068 3839 3072
rect 3843 3068 3844 3072
rect 3838 3067 3844 3068
rect 3040 3035 3042 3067
rect 3232 3035 3234 3067
rect 3432 3035 3434 3067
rect 3640 3035 3642 3067
rect 3840 3035 3842 3067
rect 3039 3034 3043 3035
rect 3039 3029 3043 3030
rect 3087 3034 3091 3035
rect 3087 3029 3091 3030
rect 3231 3034 3235 3035
rect 3231 3029 3235 3030
rect 3335 3034 3339 3035
rect 3335 3029 3339 3030
rect 3431 3034 3435 3035
rect 3431 3029 3435 3030
rect 3599 3034 3603 3035
rect 3599 3029 3603 3030
rect 3639 3034 3643 3035
rect 3639 3029 3643 3030
rect 3839 3034 3843 3035
rect 3839 3029 3843 3030
rect 2922 3011 2928 3012
rect 2922 3007 2923 3011
rect 2927 3007 2928 3011
rect 2922 3006 2928 3007
rect 3088 3005 3090 3029
rect 3336 3005 3338 3029
rect 3600 3005 3602 3029
rect 3840 3005 3842 3029
rect 2326 3004 2332 3005
rect 2326 3000 2327 3004
rect 2331 3000 2332 3004
rect 2326 2999 2332 3000
rect 2478 3004 2484 3005
rect 2478 3000 2479 3004
rect 2483 3000 2484 3004
rect 2478 2999 2484 3000
rect 2654 3004 2660 3005
rect 2654 3000 2655 3004
rect 2659 3000 2660 3004
rect 2654 2999 2660 3000
rect 2854 3004 2860 3005
rect 2854 3000 2855 3004
rect 2859 3000 2860 3004
rect 2854 2999 2860 3000
rect 3086 3004 3092 3005
rect 3086 3000 3087 3004
rect 3091 3000 3092 3004
rect 3086 2999 3092 3000
rect 3334 3004 3340 3005
rect 3334 3000 3335 3004
rect 3339 3000 3340 3004
rect 3334 2999 3340 3000
rect 3598 3004 3604 3005
rect 3598 3000 3599 3004
rect 3603 3000 3604 3004
rect 3598 2999 3604 3000
rect 3838 3004 3844 3005
rect 3838 3000 3839 3004
rect 3843 3000 3844 3004
rect 3838 2999 3844 3000
rect 2402 2995 2408 2996
rect 2402 2991 2403 2995
rect 2407 2991 2408 2995
rect 2402 2990 2408 2991
rect 2554 2995 2560 2996
rect 2554 2991 2555 2995
rect 2559 2991 2560 2995
rect 2554 2990 2560 2991
rect 2598 2995 2604 2996
rect 2598 2991 2599 2995
rect 2603 2991 2604 2995
rect 2598 2990 2604 2991
rect 2930 2995 2936 2996
rect 2930 2991 2931 2995
rect 2935 2991 2936 2995
rect 2930 2990 2936 2991
rect 3162 2995 3168 2996
rect 3162 2991 3163 2995
rect 3167 2991 3168 2995
rect 3162 2990 3168 2991
rect 3410 2995 3416 2996
rect 3410 2991 3411 2995
rect 3415 2991 3416 2995
rect 3410 2990 3416 2991
rect 3906 2995 3912 2996
rect 3906 2991 3907 2995
rect 3911 2991 3912 2995
rect 3906 2990 3912 2991
rect 2326 2985 2332 2986
rect 2326 2981 2327 2985
rect 2331 2981 2332 2985
rect 2326 2980 2332 2981
rect 2298 2963 2304 2964
rect 2298 2959 2299 2963
rect 2303 2959 2304 2963
rect 2298 2958 2304 2959
rect 2328 2955 2330 2980
rect 2404 2964 2406 2990
rect 2478 2985 2484 2986
rect 2478 2981 2479 2985
rect 2483 2981 2484 2985
rect 2478 2980 2484 2981
rect 2402 2963 2408 2964
rect 2402 2959 2403 2963
rect 2407 2959 2408 2963
rect 2402 2958 2408 2959
rect 2480 2955 2482 2980
rect 2556 2964 2558 2990
rect 2600 2972 2602 2990
rect 2654 2985 2660 2986
rect 2654 2981 2655 2985
rect 2659 2981 2660 2985
rect 2654 2980 2660 2981
rect 2854 2985 2860 2986
rect 2854 2981 2855 2985
rect 2859 2981 2860 2985
rect 2854 2980 2860 2981
rect 2598 2971 2604 2972
rect 2598 2967 2599 2971
rect 2603 2967 2604 2971
rect 2598 2966 2604 2967
rect 2554 2963 2560 2964
rect 2554 2959 2555 2963
rect 2559 2959 2560 2963
rect 2554 2958 2560 2959
rect 2656 2955 2658 2980
rect 2856 2955 2858 2980
rect 2932 2964 2934 2990
rect 3086 2985 3092 2986
rect 3086 2981 3087 2985
rect 3091 2981 3092 2985
rect 3086 2980 3092 2981
rect 2930 2963 2936 2964
rect 2930 2959 2931 2963
rect 2935 2959 2936 2963
rect 2930 2958 2936 2959
rect 3088 2955 3090 2980
rect 3164 2964 3166 2990
rect 3334 2985 3340 2986
rect 3334 2981 3335 2985
rect 3339 2981 3340 2985
rect 3334 2980 3340 2981
rect 3162 2963 3168 2964
rect 3162 2959 3163 2963
rect 3167 2959 3168 2963
rect 3162 2958 3168 2959
rect 3336 2955 3338 2980
rect 3412 2964 3414 2990
rect 3598 2985 3604 2986
rect 3598 2981 3599 2985
rect 3603 2981 3604 2985
rect 3598 2980 3604 2981
rect 3838 2985 3844 2986
rect 3838 2981 3839 2985
rect 3843 2981 3844 2985
rect 3838 2980 3844 2981
rect 3410 2963 3416 2964
rect 3410 2959 3411 2963
rect 3415 2959 3416 2963
rect 3410 2958 3416 2959
rect 3362 2955 3368 2956
rect 3600 2955 3602 2980
rect 3840 2955 3842 2980
rect 2183 2954 2187 2955
rect 2183 2949 2187 2950
rect 2263 2954 2267 2955
rect 2263 2949 2267 2950
rect 2327 2954 2331 2955
rect 2327 2949 2331 2950
rect 2479 2954 2483 2955
rect 2479 2949 2483 2950
rect 2487 2954 2491 2955
rect 2487 2949 2491 2950
rect 2655 2954 2659 2955
rect 2655 2949 2659 2950
rect 2735 2954 2739 2955
rect 2735 2949 2739 2950
rect 2855 2954 2859 2955
rect 2855 2949 2859 2950
rect 2999 2954 3003 2955
rect 2999 2949 3003 2950
rect 3087 2954 3091 2955
rect 3087 2949 3091 2950
rect 3279 2954 3283 2955
rect 3279 2949 3283 2950
rect 3335 2954 3339 2955
rect 3362 2951 3363 2955
rect 3367 2951 3368 2955
rect 3362 2950 3368 2951
rect 3567 2954 3571 2955
rect 3335 2949 3339 2950
rect 2138 2947 2144 2948
rect 2138 2943 2139 2947
rect 2143 2943 2144 2947
rect 2138 2942 2144 2943
rect 2264 2928 2266 2949
rect 2338 2947 2344 2948
rect 2330 2943 2336 2944
rect 2330 2939 2331 2943
rect 2335 2939 2336 2943
rect 2338 2943 2339 2947
rect 2343 2943 2344 2947
rect 2338 2942 2344 2943
rect 2330 2938 2336 2939
rect 2046 2924 2047 2928
rect 2051 2924 2052 2928
rect 2046 2923 2052 2924
rect 2070 2927 2076 2928
rect 2070 2923 2071 2927
rect 2075 2923 2076 2927
rect 2070 2922 2076 2923
rect 2262 2927 2268 2928
rect 2262 2923 2263 2927
rect 2267 2923 2268 2927
rect 2262 2922 2268 2923
rect 1794 2918 1800 2919
rect 1903 2918 1907 2919
rect 1903 2913 1907 2914
rect 2007 2918 2011 2919
rect 2007 2913 2011 2914
rect 1786 2911 1792 2912
rect 1786 2907 1787 2911
rect 1791 2907 1792 2911
rect 1786 2906 1792 2907
rect 1802 2911 1808 2912
rect 1802 2907 1803 2911
rect 1807 2907 1808 2911
rect 1802 2906 1808 2907
rect 1534 2891 1540 2892
rect 1534 2887 1535 2891
rect 1539 2887 1540 2891
rect 1534 2886 1540 2887
rect 1726 2891 1732 2892
rect 1726 2887 1727 2891
rect 1731 2887 1732 2891
rect 1726 2886 1732 2887
rect 1804 2884 1806 2906
rect 1904 2892 1906 2913
rect 2008 2893 2010 2913
rect 2046 2911 2052 2912
rect 2046 2907 2047 2911
rect 2051 2907 2052 2911
rect 2046 2906 2052 2907
rect 2070 2908 2076 2909
rect 2006 2892 2012 2893
rect 1902 2891 1908 2892
rect 1902 2887 1903 2891
rect 1907 2887 1908 2891
rect 2006 2888 2007 2892
rect 2011 2888 2012 2892
rect 2006 2887 2012 2888
rect 1902 2886 1908 2887
rect 974 2883 980 2884
rect 974 2879 975 2883
rect 979 2879 980 2883
rect 974 2878 980 2879
rect 990 2883 996 2884
rect 990 2879 991 2883
rect 995 2879 996 2883
rect 1250 2883 1256 2884
rect 990 2878 996 2879
rect 1242 2879 1248 2880
rect 1242 2875 1243 2879
rect 1247 2875 1248 2879
rect 1250 2879 1251 2883
rect 1255 2879 1256 2883
rect 1250 2878 1256 2879
rect 1438 2883 1444 2884
rect 1438 2879 1439 2883
rect 1443 2879 1444 2883
rect 1438 2878 1444 2879
rect 1802 2883 1808 2884
rect 1802 2879 1803 2883
rect 1807 2879 1808 2883
rect 1802 2878 1808 2879
rect 1818 2883 1824 2884
rect 1818 2879 1819 2883
rect 1823 2879 1824 2883
rect 1818 2878 1824 2879
rect 1242 2874 1248 2875
rect 998 2872 1004 2873
rect 998 2868 999 2872
rect 1003 2868 1004 2872
rect 998 2867 1004 2868
rect 1166 2872 1172 2873
rect 1166 2868 1167 2872
rect 1171 2868 1172 2872
rect 1166 2867 1172 2868
rect 1000 2839 1002 2867
rect 1168 2839 1170 2867
rect 999 2838 1003 2839
rect 999 2833 1003 2834
rect 1047 2838 1051 2839
rect 1047 2833 1051 2834
rect 1167 2838 1171 2839
rect 1167 2833 1171 2834
rect 1223 2838 1227 2839
rect 1223 2833 1227 2834
rect 1048 2809 1050 2833
rect 1224 2809 1226 2833
rect 1046 2808 1052 2809
rect 1046 2804 1047 2808
rect 1051 2804 1052 2808
rect 1046 2803 1052 2804
rect 1222 2808 1228 2809
rect 1222 2804 1223 2808
rect 1227 2804 1228 2808
rect 1222 2803 1228 2804
rect 682 2799 688 2800
rect 682 2795 683 2799
rect 687 2795 688 2799
rect 682 2794 688 2795
rect 778 2799 784 2800
rect 778 2795 779 2799
rect 783 2795 784 2799
rect 778 2794 784 2795
rect 946 2799 952 2800
rect 946 2795 947 2799
rect 951 2795 952 2799
rect 946 2794 952 2795
rect 962 2799 968 2800
rect 962 2795 963 2799
rect 967 2795 968 2799
rect 962 2794 968 2795
rect 550 2789 556 2790
rect 550 2785 551 2789
rect 555 2785 556 2789
rect 550 2784 556 2785
rect 522 2767 528 2768
rect 522 2763 523 2767
rect 527 2763 528 2767
rect 522 2762 528 2763
rect 552 2755 554 2784
rect 684 2768 686 2794
rect 710 2789 716 2790
rect 710 2785 711 2789
rect 715 2785 716 2789
rect 710 2784 716 2785
rect 878 2789 884 2790
rect 878 2785 879 2789
rect 883 2785 884 2789
rect 878 2784 884 2785
rect 650 2767 656 2768
rect 650 2763 651 2767
rect 655 2763 656 2767
rect 650 2762 656 2763
rect 682 2767 688 2768
rect 682 2763 683 2767
rect 687 2763 688 2767
rect 682 2762 688 2763
rect 247 2754 251 2755
rect 247 2749 251 2750
rect 255 2754 259 2755
rect 255 2749 259 2750
rect 399 2754 403 2755
rect 399 2749 403 2750
rect 407 2754 411 2755
rect 407 2749 411 2750
rect 551 2754 555 2755
rect 551 2749 555 2750
rect 575 2754 579 2755
rect 575 2749 579 2750
rect 202 2747 208 2748
rect 202 2743 203 2747
rect 207 2743 208 2747
rect 202 2742 208 2743
rect 210 2747 216 2748
rect 210 2743 211 2747
rect 215 2743 216 2747
rect 210 2742 216 2743
rect 110 2724 111 2728
rect 115 2724 116 2728
rect 110 2723 116 2724
rect 134 2727 140 2728
rect 134 2723 135 2727
rect 139 2723 140 2727
rect 134 2722 140 2723
rect 212 2720 214 2742
rect 256 2728 258 2749
rect 330 2747 336 2748
rect 330 2743 331 2747
rect 335 2743 336 2747
rect 330 2742 336 2743
rect 254 2727 260 2728
rect 254 2723 255 2727
rect 259 2723 260 2727
rect 254 2722 260 2723
rect 332 2720 334 2742
rect 408 2728 410 2749
rect 576 2728 578 2749
rect 406 2727 412 2728
rect 406 2723 407 2727
rect 411 2723 412 2727
rect 406 2722 412 2723
rect 574 2727 580 2728
rect 574 2723 575 2727
rect 579 2723 580 2727
rect 574 2722 580 2723
rect 652 2720 654 2762
rect 712 2755 714 2784
rect 880 2755 882 2784
rect 964 2768 966 2794
rect 1046 2789 1052 2790
rect 1046 2785 1047 2789
rect 1051 2785 1052 2789
rect 1046 2784 1052 2785
rect 1222 2789 1228 2790
rect 1222 2785 1223 2789
rect 1227 2785 1228 2789
rect 1222 2784 1228 2785
rect 962 2767 968 2768
rect 962 2763 963 2767
rect 967 2763 968 2767
rect 962 2762 968 2763
rect 1048 2755 1050 2784
rect 1162 2767 1168 2768
rect 1162 2763 1163 2767
rect 1167 2763 1168 2767
rect 1162 2762 1168 2763
rect 711 2754 715 2755
rect 711 2749 715 2750
rect 743 2754 747 2755
rect 743 2749 747 2750
rect 879 2754 883 2755
rect 879 2749 883 2750
rect 919 2754 923 2755
rect 919 2749 923 2750
rect 1047 2754 1051 2755
rect 1047 2749 1051 2750
rect 1087 2754 1091 2755
rect 1087 2749 1091 2750
rect 744 2728 746 2749
rect 826 2747 832 2748
rect 826 2743 827 2747
rect 831 2743 832 2747
rect 826 2742 832 2743
rect 742 2727 748 2728
rect 742 2723 743 2727
rect 747 2723 748 2727
rect 742 2722 748 2723
rect 210 2719 216 2720
rect 210 2715 211 2719
rect 215 2715 216 2719
rect 210 2714 216 2715
rect 330 2719 336 2720
rect 330 2715 331 2719
rect 335 2715 336 2719
rect 330 2714 336 2715
rect 342 2719 348 2720
rect 342 2715 343 2719
rect 347 2715 348 2719
rect 342 2714 348 2715
rect 650 2719 656 2720
rect 650 2715 651 2719
rect 655 2715 656 2719
rect 650 2714 656 2715
rect 110 2711 116 2712
rect 110 2707 111 2711
rect 115 2707 116 2711
rect 110 2706 116 2707
rect 134 2708 140 2709
rect 112 2679 114 2706
rect 134 2704 135 2708
rect 139 2704 140 2708
rect 134 2703 140 2704
rect 254 2708 260 2709
rect 254 2704 255 2708
rect 259 2704 260 2708
rect 254 2703 260 2704
rect 136 2679 138 2703
rect 256 2679 258 2703
rect 111 2678 115 2679
rect 111 2673 115 2674
rect 135 2678 139 2679
rect 135 2673 139 2674
rect 167 2678 171 2679
rect 167 2673 171 2674
rect 255 2678 259 2679
rect 255 2673 259 2674
rect 112 2646 114 2673
rect 168 2649 170 2673
rect 166 2648 172 2649
rect 110 2645 116 2646
rect 110 2641 111 2645
rect 115 2641 116 2645
rect 166 2644 167 2648
rect 171 2644 172 2648
rect 166 2643 172 2644
rect 110 2640 116 2641
rect 282 2639 288 2640
rect 282 2635 283 2639
rect 287 2635 288 2639
rect 282 2634 288 2635
rect 166 2629 172 2630
rect 110 2628 116 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 166 2625 167 2629
rect 171 2625 172 2629
rect 166 2624 172 2625
rect 110 2623 116 2624
rect 112 2587 114 2623
rect 168 2587 170 2624
rect 284 2604 286 2634
rect 344 2616 346 2714
rect 406 2708 412 2709
rect 406 2704 407 2708
rect 411 2704 412 2708
rect 406 2703 412 2704
rect 574 2708 580 2709
rect 574 2704 575 2708
rect 579 2704 580 2708
rect 574 2703 580 2704
rect 742 2708 748 2709
rect 742 2704 743 2708
rect 747 2704 748 2708
rect 742 2703 748 2704
rect 408 2679 410 2703
rect 576 2679 578 2703
rect 744 2679 746 2703
rect 359 2678 363 2679
rect 359 2673 363 2674
rect 407 2678 411 2679
rect 407 2673 411 2674
rect 559 2678 563 2679
rect 559 2673 563 2674
rect 575 2678 579 2679
rect 575 2673 579 2674
rect 743 2678 747 2679
rect 743 2673 747 2674
rect 759 2678 763 2679
rect 759 2673 763 2674
rect 360 2649 362 2673
rect 560 2649 562 2673
rect 760 2649 762 2673
rect 358 2648 364 2649
rect 358 2644 359 2648
rect 363 2644 364 2648
rect 358 2643 364 2644
rect 558 2648 564 2649
rect 558 2644 559 2648
rect 563 2644 564 2648
rect 558 2643 564 2644
rect 758 2648 764 2649
rect 758 2644 759 2648
rect 763 2644 764 2648
rect 758 2643 764 2644
rect 828 2640 830 2742
rect 920 2728 922 2749
rect 1018 2747 1024 2748
rect 1018 2743 1019 2747
rect 1023 2743 1024 2747
rect 1018 2742 1024 2743
rect 1054 2747 1060 2748
rect 1054 2743 1055 2747
rect 1059 2743 1060 2747
rect 1054 2742 1060 2743
rect 918 2727 924 2728
rect 918 2723 919 2727
rect 923 2723 924 2727
rect 918 2722 924 2723
rect 918 2708 924 2709
rect 918 2704 919 2708
rect 923 2704 924 2708
rect 918 2703 924 2704
rect 920 2679 922 2703
rect 919 2678 923 2679
rect 919 2673 923 2674
rect 951 2678 955 2679
rect 951 2673 955 2674
rect 952 2649 954 2673
rect 950 2648 956 2649
rect 950 2644 951 2648
rect 955 2644 956 2648
rect 950 2643 956 2644
rect 1020 2640 1022 2742
rect 1056 2720 1058 2742
rect 1088 2728 1090 2749
rect 1086 2727 1092 2728
rect 1086 2723 1087 2727
rect 1091 2723 1092 2727
rect 1086 2722 1092 2723
rect 1164 2720 1166 2762
rect 1224 2755 1226 2784
rect 1244 2768 1246 2874
rect 1350 2872 1356 2873
rect 1350 2868 1351 2872
rect 1355 2868 1356 2872
rect 1350 2867 1356 2868
rect 1534 2872 1540 2873
rect 1534 2868 1535 2872
rect 1539 2868 1540 2872
rect 1534 2867 1540 2868
rect 1726 2872 1732 2873
rect 1726 2868 1727 2872
rect 1731 2868 1732 2872
rect 1726 2867 1732 2868
rect 1352 2839 1354 2867
rect 1536 2839 1538 2867
rect 1728 2839 1730 2867
rect 1351 2838 1355 2839
rect 1351 2833 1355 2834
rect 1399 2838 1403 2839
rect 1399 2833 1403 2834
rect 1535 2838 1539 2839
rect 1535 2833 1539 2834
rect 1575 2838 1579 2839
rect 1575 2833 1579 2834
rect 1727 2838 1731 2839
rect 1727 2833 1731 2834
rect 1751 2838 1755 2839
rect 1751 2833 1755 2834
rect 1400 2809 1402 2833
rect 1576 2809 1578 2833
rect 1752 2809 1754 2833
rect 1398 2808 1404 2809
rect 1398 2804 1399 2808
rect 1403 2804 1404 2808
rect 1398 2803 1404 2804
rect 1574 2808 1580 2809
rect 1574 2804 1575 2808
rect 1579 2804 1580 2808
rect 1574 2803 1580 2804
rect 1750 2808 1756 2809
rect 1750 2804 1751 2808
rect 1755 2804 1756 2808
rect 1750 2803 1756 2804
rect 1298 2799 1304 2800
rect 1298 2795 1299 2799
rect 1303 2795 1304 2799
rect 1298 2794 1304 2795
rect 1474 2799 1480 2800
rect 1474 2795 1475 2799
rect 1479 2795 1480 2799
rect 1474 2794 1480 2795
rect 1650 2799 1656 2800
rect 1650 2795 1651 2799
rect 1655 2795 1656 2799
rect 1650 2794 1656 2795
rect 1300 2768 1302 2794
rect 1398 2789 1404 2790
rect 1398 2785 1399 2789
rect 1403 2785 1404 2789
rect 1398 2784 1404 2785
rect 1242 2767 1248 2768
rect 1242 2763 1243 2767
rect 1247 2763 1248 2767
rect 1242 2762 1248 2763
rect 1298 2767 1304 2768
rect 1298 2763 1299 2767
rect 1303 2763 1304 2767
rect 1298 2762 1304 2763
rect 1400 2755 1402 2784
rect 1476 2768 1478 2794
rect 1574 2789 1580 2790
rect 1574 2785 1575 2789
rect 1579 2785 1580 2789
rect 1574 2784 1580 2785
rect 1474 2767 1480 2768
rect 1474 2763 1475 2767
rect 1479 2763 1480 2767
rect 1474 2762 1480 2763
rect 1576 2755 1578 2784
rect 1223 2754 1227 2755
rect 1223 2749 1227 2750
rect 1255 2754 1259 2755
rect 1255 2749 1259 2750
rect 1399 2754 1403 2755
rect 1399 2749 1403 2750
rect 1423 2754 1427 2755
rect 1423 2749 1427 2750
rect 1575 2754 1579 2755
rect 1575 2749 1579 2750
rect 1599 2754 1603 2755
rect 1599 2749 1603 2750
rect 1256 2728 1258 2749
rect 1338 2747 1344 2748
rect 1338 2743 1339 2747
rect 1343 2743 1344 2747
rect 1338 2742 1344 2743
rect 1254 2727 1260 2728
rect 1254 2723 1255 2727
rect 1259 2723 1260 2727
rect 1254 2722 1260 2723
rect 1340 2720 1342 2742
rect 1424 2728 1426 2749
rect 1600 2728 1602 2749
rect 1652 2748 1654 2794
rect 1750 2789 1756 2790
rect 1750 2785 1751 2789
rect 1755 2785 1756 2789
rect 1750 2784 1756 2785
rect 1752 2755 1754 2784
rect 1820 2768 1822 2878
rect 2006 2875 2012 2876
rect 1902 2872 1908 2873
rect 1902 2868 1903 2872
rect 1907 2868 1908 2872
rect 2006 2871 2007 2875
rect 2011 2871 2012 2875
rect 2048 2871 2050 2906
rect 2070 2904 2071 2908
rect 2075 2904 2076 2908
rect 2070 2903 2076 2904
rect 2262 2908 2268 2909
rect 2262 2904 2263 2908
rect 2267 2904 2268 2908
rect 2262 2903 2268 2904
rect 2072 2871 2074 2903
rect 2264 2871 2266 2903
rect 2006 2870 2012 2871
rect 2047 2870 2051 2871
rect 1902 2867 1908 2868
rect 1904 2839 1906 2867
rect 2008 2839 2010 2870
rect 2047 2865 2051 2866
rect 2071 2870 2075 2871
rect 2071 2865 2075 2866
rect 2263 2870 2267 2871
rect 2263 2865 2267 2866
rect 1903 2838 1907 2839
rect 1903 2833 1907 2834
rect 2007 2838 2011 2839
rect 2048 2838 2050 2865
rect 2007 2833 2011 2834
rect 2046 2837 2052 2838
rect 2046 2833 2047 2837
rect 2051 2833 2052 2837
rect 1904 2809 1906 2833
rect 1902 2808 1908 2809
rect 1902 2804 1903 2808
rect 1907 2804 1908 2808
rect 2008 2806 2010 2833
rect 2046 2832 2052 2833
rect 2332 2832 2334 2938
rect 2340 2920 2342 2942
rect 2488 2928 2490 2949
rect 2562 2947 2568 2948
rect 2562 2943 2563 2947
rect 2567 2943 2568 2947
rect 2562 2942 2568 2943
rect 2486 2927 2492 2928
rect 2486 2923 2487 2927
rect 2491 2923 2492 2927
rect 2486 2922 2492 2923
rect 2564 2920 2566 2942
rect 2736 2928 2738 2949
rect 2810 2947 2816 2948
rect 2810 2943 2811 2947
rect 2815 2943 2816 2947
rect 2810 2942 2816 2943
rect 2734 2927 2740 2928
rect 2734 2923 2735 2927
rect 2739 2923 2740 2927
rect 2734 2922 2740 2923
rect 2812 2920 2814 2942
rect 3000 2928 3002 2949
rect 3074 2947 3080 2948
rect 3074 2943 3075 2947
rect 3079 2943 3080 2947
rect 3074 2942 3080 2943
rect 2998 2927 3004 2928
rect 2998 2923 2999 2927
rect 3003 2923 3004 2927
rect 2998 2922 3004 2923
rect 3076 2920 3078 2942
rect 3280 2928 3282 2949
rect 3354 2947 3360 2948
rect 3354 2943 3355 2947
rect 3359 2943 3360 2947
rect 3354 2942 3360 2943
rect 3278 2927 3284 2928
rect 3278 2923 3279 2927
rect 3283 2923 3284 2927
rect 3278 2922 3284 2923
rect 3356 2920 3358 2942
rect 3364 2920 3366 2950
rect 3567 2949 3571 2950
rect 3599 2954 3603 2955
rect 3599 2949 3603 2950
rect 3839 2954 3843 2955
rect 3839 2949 3843 2950
rect 3568 2928 3570 2949
rect 3840 2928 3842 2949
rect 3908 2948 3910 2990
rect 3916 2964 3918 3074
rect 3942 3071 3943 3075
rect 3947 3071 3948 3075
rect 3942 3070 3948 3071
rect 3944 3035 3946 3070
rect 3943 3034 3947 3035
rect 3943 3029 3947 3030
rect 3944 3002 3946 3029
rect 3942 3001 3948 3002
rect 3942 2997 3943 3001
rect 3947 2997 3948 3001
rect 3942 2996 3948 2997
rect 3942 2984 3948 2985
rect 3942 2980 3943 2984
rect 3947 2980 3948 2984
rect 3942 2979 3948 2980
rect 3914 2963 3920 2964
rect 3914 2959 3915 2963
rect 3919 2959 3920 2963
rect 3914 2958 3920 2959
rect 3944 2955 3946 2979
rect 3943 2954 3947 2955
rect 3943 2949 3947 2950
rect 3906 2947 3912 2948
rect 3906 2943 3907 2947
rect 3911 2943 3912 2947
rect 3906 2942 3912 2943
rect 3944 2929 3946 2949
rect 3942 2928 3948 2929
rect 3566 2927 3572 2928
rect 3566 2923 3567 2927
rect 3571 2923 3572 2927
rect 3566 2922 3572 2923
rect 3838 2927 3844 2928
rect 3838 2923 3839 2927
rect 3843 2923 3844 2927
rect 3942 2924 3943 2928
rect 3947 2924 3948 2928
rect 3942 2923 3948 2924
rect 3838 2922 3844 2923
rect 2338 2919 2344 2920
rect 2338 2915 2339 2919
rect 2343 2915 2344 2919
rect 2338 2914 2344 2915
rect 2562 2919 2568 2920
rect 2562 2915 2563 2919
rect 2567 2915 2568 2919
rect 2562 2914 2568 2915
rect 2810 2919 2816 2920
rect 2810 2915 2811 2919
rect 2815 2915 2816 2919
rect 2810 2914 2816 2915
rect 3074 2919 3080 2920
rect 3074 2915 3075 2919
rect 3079 2915 3080 2919
rect 3074 2914 3080 2915
rect 3354 2919 3360 2920
rect 3354 2915 3355 2919
rect 3359 2915 3360 2919
rect 3354 2914 3360 2915
rect 3362 2919 3368 2920
rect 3362 2915 3363 2919
rect 3367 2915 3368 2919
rect 3362 2914 3368 2915
rect 3914 2915 3920 2916
rect 3914 2911 3915 2915
rect 3919 2911 3920 2915
rect 3914 2910 3920 2911
rect 3942 2911 3948 2912
rect 2486 2908 2492 2909
rect 2486 2904 2487 2908
rect 2491 2904 2492 2908
rect 2486 2903 2492 2904
rect 2734 2908 2740 2909
rect 2734 2904 2735 2908
rect 2739 2904 2740 2908
rect 2734 2903 2740 2904
rect 2998 2908 3004 2909
rect 2998 2904 2999 2908
rect 3003 2904 3004 2908
rect 2998 2903 3004 2904
rect 3278 2908 3284 2909
rect 3278 2904 3279 2908
rect 3283 2904 3284 2908
rect 3278 2903 3284 2904
rect 3566 2908 3572 2909
rect 3566 2904 3567 2908
rect 3571 2904 3572 2908
rect 3566 2903 3572 2904
rect 3838 2908 3844 2909
rect 3838 2904 3839 2908
rect 3843 2904 3844 2908
rect 3838 2903 3844 2904
rect 2488 2871 2490 2903
rect 2736 2871 2738 2903
rect 3000 2871 3002 2903
rect 3280 2871 3282 2903
rect 3568 2871 3570 2903
rect 3840 2871 3842 2903
rect 2487 2870 2491 2871
rect 2487 2865 2491 2866
rect 2671 2870 2675 2871
rect 2671 2865 2675 2866
rect 2735 2870 2739 2871
rect 2735 2865 2739 2866
rect 2887 2870 2891 2871
rect 2887 2865 2891 2866
rect 2999 2870 3003 2871
rect 2999 2865 3003 2866
rect 3095 2870 3099 2871
rect 3095 2865 3099 2866
rect 3279 2870 3283 2871
rect 3279 2865 3283 2866
rect 3287 2870 3291 2871
rect 3287 2865 3291 2866
rect 3479 2870 3483 2871
rect 3479 2865 3483 2866
rect 3567 2870 3571 2871
rect 3567 2865 3571 2866
rect 3671 2870 3675 2871
rect 3671 2865 3675 2866
rect 3839 2870 3843 2871
rect 3839 2865 3843 2866
rect 2672 2841 2674 2865
rect 2888 2841 2890 2865
rect 3096 2841 3098 2865
rect 3288 2841 3290 2865
rect 3480 2841 3482 2865
rect 3672 2841 3674 2865
rect 3840 2841 3842 2865
rect 2670 2840 2676 2841
rect 2670 2836 2671 2840
rect 2675 2836 2676 2840
rect 2670 2835 2676 2836
rect 2886 2840 2892 2841
rect 2886 2836 2887 2840
rect 2891 2836 2892 2840
rect 2886 2835 2892 2836
rect 3094 2840 3100 2841
rect 3094 2836 3095 2840
rect 3099 2836 3100 2840
rect 3094 2835 3100 2836
rect 3286 2840 3292 2841
rect 3286 2836 3287 2840
rect 3291 2836 3292 2840
rect 3286 2835 3292 2836
rect 3478 2840 3484 2841
rect 3478 2836 3479 2840
rect 3483 2836 3484 2840
rect 3478 2835 3484 2836
rect 3670 2840 3676 2841
rect 3670 2836 3671 2840
rect 3675 2836 3676 2840
rect 3670 2835 3676 2836
rect 3838 2840 3844 2841
rect 3838 2836 3839 2840
rect 3843 2836 3844 2840
rect 3838 2835 3844 2836
rect 3916 2833 3918 2910
rect 3942 2907 3943 2911
rect 3947 2907 3948 2911
rect 3942 2906 3948 2907
rect 3944 2871 3946 2906
rect 3943 2870 3947 2871
rect 3943 2865 3947 2866
rect 3944 2838 3946 2865
rect 2330 2831 2336 2832
rect 2330 2827 2331 2831
rect 2335 2827 2336 2831
rect 2330 2826 2336 2827
rect 2746 2831 2752 2832
rect 2746 2827 2747 2831
rect 2751 2827 2752 2831
rect 2746 2826 2752 2827
rect 2962 2831 2968 2832
rect 2962 2827 2963 2831
rect 2967 2827 2968 2831
rect 2962 2826 2968 2827
rect 3354 2831 3360 2832
rect 3354 2827 3355 2831
rect 3359 2827 3360 2831
rect 3354 2826 3360 2827
rect 3370 2831 3376 2832
rect 3370 2827 3371 2831
rect 3375 2827 3376 2831
rect 3370 2826 3376 2827
rect 3754 2831 3760 2832
rect 3754 2827 3755 2831
rect 3759 2827 3760 2831
rect 3754 2826 3760 2827
rect 3908 2831 3918 2833
rect 3942 2837 3948 2838
rect 3942 2833 3943 2837
rect 3947 2833 3948 2837
rect 3942 2832 3948 2833
rect 2670 2821 2676 2822
rect 2046 2820 2052 2821
rect 2046 2816 2047 2820
rect 2051 2816 2052 2820
rect 2670 2817 2671 2821
rect 2675 2817 2676 2821
rect 2670 2816 2676 2817
rect 2046 2815 2052 2816
rect 1902 2803 1908 2804
rect 2006 2805 2012 2806
rect 2006 2801 2007 2805
rect 2011 2801 2012 2805
rect 2006 2800 2012 2801
rect 1826 2799 1832 2800
rect 1826 2795 1827 2799
rect 1831 2795 1832 2799
rect 2048 2795 2050 2815
rect 2672 2795 2674 2816
rect 2748 2800 2750 2826
rect 2886 2821 2892 2822
rect 2886 2817 2887 2821
rect 2891 2817 2892 2821
rect 2886 2816 2892 2817
rect 2682 2799 2688 2800
rect 2682 2795 2683 2799
rect 2687 2795 2688 2799
rect 2746 2799 2752 2800
rect 2746 2795 2747 2799
rect 2751 2795 2752 2799
rect 2888 2795 2890 2816
rect 2964 2800 2966 2826
rect 3094 2821 3100 2822
rect 3094 2817 3095 2821
rect 3099 2817 3100 2821
rect 3094 2816 3100 2817
rect 3286 2821 3292 2822
rect 3286 2817 3287 2821
rect 3291 2817 3292 2821
rect 3286 2816 3292 2817
rect 2962 2799 2968 2800
rect 2962 2795 2963 2799
rect 2967 2795 2968 2799
rect 3096 2795 3098 2816
rect 3288 2795 3290 2816
rect 1826 2794 1832 2795
rect 2047 2794 2051 2795
rect 1828 2768 1830 2794
rect 1902 2789 1908 2790
rect 2047 2789 2051 2790
rect 2071 2794 2075 2795
rect 2071 2789 2075 2790
rect 2199 2794 2203 2795
rect 2199 2789 2203 2790
rect 2343 2794 2347 2795
rect 2343 2789 2347 2790
rect 2479 2794 2483 2795
rect 2479 2789 2483 2790
rect 2607 2794 2611 2795
rect 2607 2789 2611 2790
rect 2671 2794 2675 2795
rect 2682 2794 2688 2795
rect 2727 2794 2731 2795
rect 2746 2794 2752 2795
rect 2839 2794 2843 2795
rect 2671 2789 2675 2790
rect 1902 2785 1903 2789
rect 1907 2785 1908 2789
rect 1902 2784 1908 2785
rect 2006 2788 2012 2789
rect 2006 2784 2007 2788
rect 2011 2784 2012 2788
rect 1818 2767 1824 2768
rect 1818 2763 1819 2767
rect 1823 2763 1824 2767
rect 1818 2762 1824 2763
rect 1826 2767 1832 2768
rect 1826 2763 1827 2767
rect 1831 2763 1832 2767
rect 1826 2762 1832 2763
rect 1904 2755 1906 2784
rect 2006 2783 2012 2784
rect 2008 2755 2010 2783
rect 2048 2769 2050 2789
rect 2046 2768 2052 2769
rect 2072 2768 2074 2789
rect 2146 2787 2152 2788
rect 2146 2783 2147 2787
rect 2151 2783 2152 2787
rect 2146 2782 2152 2783
rect 2046 2764 2047 2768
rect 2051 2764 2052 2768
rect 2046 2763 2052 2764
rect 2070 2767 2076 2768
rect 2070 2763 2071 2767
rect 2075 2763 2076 2767
rect 2070 2762 2076 2763
rect 2148 2760 2150 2782
rect 2200 2768 2202 2789
rect 2344 2768 2346 2789
rect 2410 2787 2416 2788
rect 2410 2783 2411 2787
rect 2415 2783 2416 2787
rect 2410 2782 2416 2783
rect 2418 2787 2424 2788
rect 2418 2783 2419 2787
rect 2423 2783 2424 2787
rect 2418 2782 2424 2783
rect 2198 2767 2204 2768
rect 2198 2763 2199 2767
rect 2203 2763 2204 2767
rect 2198 2762 2204 2763
rect 2342 2767 2348 2768
rect 2342 2763 2343 2767
rect 2347 2763 2348 2767
rect 2342 2762 2348 2763
rect 2146 2759 2152 2760
rect 2146 2755 2147 2759
rect 2151 2755 2152 2759
rect 1751 2754 1755 2755
rect 1751 2749 1755 2750
rect 1903 2754 1907 2755
rect 1903 2749 1907 2750
rect 2007 2754 2011 2755
rect 2146 2754 2152 2755
rect 2162 2759 2168 2760
rect 2162 2755 2163 2759
rect 2167 2755 2168 2759
rect 2162 2754 2168 2755
rect 2007 2749 2011 2750
rect 2046 2751 2052 2752
rect 1650 2747 1656 2748
rect 1650 2743 1651 2747
rect 1655 2743 1656 2747
rect 1650 2742 1656 2743
rect 2008 2729 2010 2749
rect 2046 2747 2047 2751
rect 2051 2747 2052 2751
rect 2046 2746 2052 2747
rect 2070 2748 2076 2749
rect 2006 2728 2012 2729
rect 1422 2727 1428 2728
rect 1422 2723 1423 2727
rect 1427 2723 1428 2727
rect 1422 2722 1428 2723
rect 1598 2727 1604 2728
rect 1598 2723 1599 2727
rect 1603 2723 1604 2727
rect 2006 2724 2007 2728
rect 2011 2724 2012 2728
rect 2006 2723 2012 2724
rect 1598 2722 1604 2723
rect 1054 2719 1060 2720
rect 1054 2715 1055 2719
rect 1059 2715 1060 2719
rect 1054 2714 1060 2715
rect 1162 2719 1168 2720
rect 1162 2715 1163 2719
rect 1167 2715 1168 2719
rect 1162 2714 1168 2715
rect 1338 2719 1344 2720
rect 1338 2715 1339 2719
rect 1343 2715 1344 2719
rect 1338 2714 1344 2715
rect 1342 2711 1348 2712
rect 1086 2708 1092 2709
rect 1086 2704 1087 2708
rect 1091 2704 1092 2708
rect 1086 2703 1092 2704
rect 1254 2708 1260 2709
rect 1254 2704 1255 2708
rect 1259 2704 1260 2708
rect 1342 2707 1343 2711
rect 1347 2707 1348 2711
rect 2006 2711 2012 2712
rect 1342 2706 1348 2707
rect 1422 2708 1428 2709
rect 1254 2703 1260 2704
rect 1088 2679 1090 2703
rect 1256 2679 1258 2703
rect 1087 2678 1091 2679
rect 1087 2673 1091 2674
rect 1143 2678 1147 2679
rect 1143 2673 1147 2674
rect 1255 2678 1259 2679
rect 1255 2673 1259 2674
rect 1327 2678 1331 2679
rect 1327 2673 1331 2674
rect 1144 2649 1146 2673
rect 1328 2649 1330 2673
rect 1142 2648 1148 2649
rect 1142 2644 1143 2648
rect 1147 2644 1148 2648
rect 1142 2643 1148 2644
rect 1326 2648 1332 2649
rect 1326 2644 1327 2648
rect 1331 2644 1332 2648
rect 1326 2643 1332 2644
rect 434 2639 440 2640
rect 434 2635 435 2639
rect 439 2635 440 2639
rect 434 2634 440 2635
rect 634 2639 640 2640
rect 634 2635 635 2639
rect 639 2635 640 2639
rect 634 2634 640 2635
rect 826 2639 832 2640
rect 826 2635 827 2639
rect 831 2635 832 2639
rect 826 2634 832 2635
rect 1018 2639 1024 2640
rect 1018 2635 1019 2639
rect 1023 2635 1024 2639
rect 1018 2634 1024 2635
rect 1034 2639 1040 2640
rect 1034 2635 1035 2639
rect 1039 2635 1040 2639
rect 1034 2634 1040 2635
rect 358 2629 364 2630
rect 358 2625 359 2629
rect 363 2625 364 2629
rect 358 2624 364 2625
rect 342 2615 348 2616
rect 342 2611 343 2615
rect 347 2611 348 2615
rect 342 2610 348 2611
rect 282 2603 288 2604
rect 282 2599 283 2603
rect 287 2599 288 2603
rect 282 2598 288 2599
rect 360 2587 362 2624
rect 436 2608 438 2634
rect 558 2629 564 2630
rect 558 2625 559 2629
rect 563 2625 564 2629
rect 558 2624 564 2625
rect 434 2607 440 2608
rect 434 2603 435 2607
rect 439 2603 440 2607
rect 434 2602 440 2603
rect 560 2587 562 2624
rect 636 2608 638 2634
rect 758 2629 764 2630
rect 758 2625 759 2629
rect 763 2625 764 2629
rect 758 2624 764 2625
rect 950 2629 956 2630
rect 950 2625 951 2629
rect 955 2625 956 2629
rect 950 2624 956 2625
rect 634 2607 640 2608
rect 634 2603 635 2607
rect 639 2603 640 2607
rect 634 2602 640 2603
rect 760 2587 762 2624
rect 952 2587 954 2624
rect 1036 2608 1038 2634
rect 1142 2629 1148 2630
rect 1142 2625 1143 2629
rect 1147 2625 1148 2629
rect 1142 2624 1148 2625
rect 1326 2629 1332 2630
rect 1326 2625 1327 2629
rect 1331 2625 1332 2629
rect 1326 2624 1332 2625
rect 1034 2607 1040 2608
rect 1034 2603 1035 2607
rect 1039 2603 1040 2607
rect 1034 2602 1040 2603
rect 1144 2587 1146 2624
rect 1198 2607 1204 2608
rect 1198 2603 1199 2607
rect 1203 2603 1204 2607
rect 1198 2602 1204 2603
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 167 2586 171 2587
rect 167 2581 171 2582
rect 359 2586 363 2587
rect 359 2581 363 2582
rect 559 2586 563 2587
rect 559 2581 563 2582
rect 575 2586 579 2587
rect 575 2581 579 2582
rect 687 2586 691 2587
rect 687 2581 691 2582
rect 759 2586 763 2587
rect 759 2581 763 2582
rect 807 2586 811 2587
rect 807 2581 811 2582
rect 935 2586 939 2587
rect 935 2581 939 2582
rect 951 2586 955 2587
rect 951 2581 955 2582
rect 1071 2586 1075 2587
rect 1071 2581 1075 2582
rect 1143 2586 1147 2587
rect 1143 2581 1147 2582
rect 112 2561 114 2581
rect 110 2560 116 2561
rect 576 2560 578 2581
rect 650 2579 656 2580
rect 650 2575 651 2579
rect 655 2575 656 2579
rect 650 2574 656 2575
rect 110 2556 111 2560
rect 115 2556 116 2560
rect 110 2555 116 2556
rect 574 2559 580 2560
rect 574 2555 575 2559
rect 579 2555 580 2559
rect 574 2554 580 2555
rect 652 2552 654 2574
rect 688 2560 690 2581
rect 782 2579 788 2580
rect 782 2575 783 2579
rect 787 2575 788 2579
rect 782 2574 788 2575
rect 702 2571 708 2572
rect 702 2567 703 2571
rect 707 2567 708 2571
rect 702 2566 708 2567
rect 686 2559 692 2560
rect 686 2555 687 2559
rect 691 2555 692 2559
rect 686 2554 692 2555
rect 650 2551 656 2552
rect 650 2547 651 2551
rect 655 2547 656 2551
rect 650 2546 656 2547
rect 110 2543 116 2544
rect 110 2539 111 2543
rect 115 2539 116 2543
rect 110 2538 116 2539
rect 574 2540 580 2541
rect 112 2507 114 2538
rect 574 2536 575 2540
rect 579 2536 580 2540
rect 574 2535 580 2536
rect 686 2540 692 2541
rect 686 2536 687 2540
rect 691 2536 692 2540
rect 686 2535 692 2536
rect 576 2507 578 2535
rect 688 2507 690 2535
rect 111 2506 115 2507
rect 111 2501 115 2502
rect 503 2506 507 2507
rect 503 2501 507 2502
rect 575 2506 579 2507
rect 575 2501 579 2502
rect 607 2506 611 2507
rect 607 2501 611 2502
rect 687 2506 691 2507
rect 687 2501 691 2502
rect 112 2474 114 2501
rect 504 2477 506 2501
rect 608 2477 610 2501
rect 502 2476 508 2477
rect 110 2473 116 2474
rect 110 2469 111 2473
rect 115 2469 116 2473
rect 502 2472 503 2476
rect 507 2472 508 2476
rect 502 2471 508 2472
rect 606 2476 612 2477
rect 606 2472 607 2476
rect 611 2472 612 2476
rect 606 2471 612 2472
rect 110 2468 116 2469
rect 704 2468 706 2566
rect 784 2552 786 2574
rect 808 2560 810 2581
rect 882 2579 888 2580
rect 882 2575 883 2579
rect 887 2575 888 2579
rect 882 2574 888 2575
rect 806 2559 812 2560
rect 806 2555 807 2559
rect 811 2555 812 2559
rect 806 2554 812 2555
rect 884 2552 886 2574
rect 936 2560 938 2581
rect 1010 2579 1016 2580
rect 1010 2575 1011 2579
rect 1015 2575 1016 2579
rect 1010 2574 1016 2575
rect 934 2559 940 2560
rect 934 2555 935 2559
rect 939 2555 940 2559
rect 934 2554 940 2555
rect 1012 2552 1014 2574
rect 1072 2560 1074 2581
rect 1070 2559 1076 2560
rect 1070 2555 1071 2559
rect 1075 2555 1076 2559
rect 1070 2554 1076 2555
rect 1200 2552 1202 2602
rect 1328 2587 1330 2624
rect 1344 2608 1346 2706
rect 1422 2704 1423 2708
rect 1427 2704 1428 2708
rect 1422 2703 1428 2704
rect 1598 2708 1604 2709
rect 1598 2704 1599 2708
rect 1603 2704 1604 2708
rect 2006 2707 2007 2711
rect 2011 2707 2012 2711
rect 2006 2706 2012 2707
rect 1598 2703 1604 2704
rect 1424 2679 1426 2703
rect 1600 2679 1602 2703
rect 2008 2679 2010 2706
rect 2048 2699 2050 2746
rect 2070 2744 2071 2748
rect 2075 2744 2076 2748
rect 2070 2743 2076 2744
rect 2072 2699 2074 2743
rect 2047 2698 2051 2699
rect 2047 2693 2051 2694
rect 2071 2698 2075 2699
rect 2071 2693 2075 2694
rect 2095 2698 2099 2699
rect 2095 2693 2099 2694
rect 1423 2678 1427 2679
rect 1423 2673 1427 2674
rect 1511 2678 1515 2679
rect 1511 2673 1515 2674
rect 1599 2678 1603 2679
rect 1599 2673 1603 2674
rect 1703 2678 1707 2679
rect 1703 2673 1707 2674
rect 2007 2678 2011 2679
rect 2007 2673 2011 2674
rect 1512 2649 1514 2673
rect 1704 2649 1706 2673
rect 1510 2648 1516 2649
rect 1510 2644 1511 2648
rect 1515 2644 1516 2648
rect 1510 2643 1516 2644
rect 1702 2648 1708 2649
rect 1702 2644 1703 2648
rect 1707 2644 1708 2648
rect 2008 2646 2010 2673
rect 2048 2666 2050 2693
rect 2096 2669 2098 2693
rect 2094 2668 2100 2669
rect 2046 2665 2052 2666
rect 2046 2661 2047 2665
rect 2051 2661 2052 2665
rect 2094 2664 2095 2668
rect 2099 2664 2100 2668
rect 2094 2663 2100 2664
rect 2046 2660 2052 2661
rect 2094 2649 2100 2650
rect 2046 2648 2052 2649
rect 1702 2643 1708 2644
rect 2006 2645 2012 2646
rect 2006 2641 2007 2645
rect 2011 2641 2012 2645
rect 2046 2644 2047 2648
rect 2051 2644 2052 2648
rect 2094 2645 2095 2649
rect 2099 2645 2100 2649
rect 2094 2644 2100 2645
rect 2046 2643 2052 2644
rect 2006 2640 2012 2641
rect 1402 2639 1408 2640
rect 1402 2635 1403 2639
rect 1407 2635 1408 2639
rect 1402 2634 1408 2635
rect 1586 2639 1592 2640
rect 1586 2635 1587 2639
rect 1591 2635 1592 2639
rect 1586 2634 1592 2635
rect 1778 2639 1784 2640
rect 1778 2635 1779 2639
rect 1783 2635 1784 2639
rect 1778 2634 1784 2635
rect 1404 2608 1406 2634
rect 1510 2629 1516 2630
rect 1510 2625 1511 2629
rect 1515 2625 1516 2629
rect 1510 2624 1516 2625
rect 1342 2607 1348 2608
rect 1342 2603 1343 2607
rect 1347 2603 1348 2607
rect 1342 2602 1348 2603
rect 1402 2607 1408 2608
rect 1402 2603 1403 2607
rect 1407 2603 1408 2607
rect 1402 2602 1408 2603
rect 1512 2587 1514 2624
rect 1588 2608 1590 2634
rect 1702 2629 1708 2630
rect 1702 2625 1703 2629
rect 1707 2625 1708 2629
rect 1702 2624 1708 2625
rect 1586 2607 1592 2608
rect 1586 2603 1587 2607
rect 1591 2603 1592 2607
rect 1586 2602 1592 2603
rect 1704 2587 1706 2624
rect 1207 2586 1211 2587
rect 1207 2581 1211 2582
rect 1327 2586 1331 2587
rect 1327 2581 1331 2582
rect 1351 2586 1355 2587
rect 1351 2581 1355 2582
rect 1495 2586 1499 2587
rect 1495 2581 1499 2582
rect 1511 2586 1515 2587
rect 1511 2581 1515 2582
rect 1647 2586 1651 2587
rect 1647 2581 1651 2582
rect 1703 2586 1707 2587
rect 1703 2581 1707 2582
rect 1208 2560 1210 2581
rect 1352 2560 1354 2581
rect 1358 2579 1364 2580
rect 1358 2575 1359 2579
rect 1363 2575 1364 2579
rect 1358 2574 1364 2575
rect 1206 2559 1212 2560
rect 1206 2555 1207 2559
rect 1211 2555 1212 2559
rect 1206 2554 1212 2555
rect 1350 2559 1356 2560
rect 1350 2555 1351 2559
rect 1355 2555 1356 2559
rect 1350 2554 1356 2555
rect 782 2551 788 2552
rect 782 2547 783 2551
rect 787 2547 788 2551
rect 782 2546 788 2547
rect 882 2551 888 2552
rect 882 2547 883 2551
rect 887 2547 888 2551
rect 882 2546 888 2547
rect 1010 2551 1016 2552
rect 1010 2547 1011 2551
rect 1015 2547 1016 2551
rect 1198 2551 1204 2552
rect 1010 2546 1016 2547
rect 1146 2547 1152 2548
rect 1146 2543 1147 2547
rect 1151 2543 1152 2547
rect 1198 2547 1199 2551
rect 1203 2547 1204 2551
rect 1198 2546 1204 2547
rect 1146 2542 1152 2543
rect 806 2540 812 2541
rect 806 2536 807 2540
rect 811 2536 812 2540
rect 806 2535 812 2536
rect 934 2540 940 2541
rect 934 2536 935 2540
rect 939 2536 940 2540
rect 934 2535 940 2536
rect 1070 2540 1076 2541
rect 1070 2536 1071 2540
rect 1075 2536 1076 2540
rect 1070 2535 1076 2536
rect 808 2507 810 2535
rect 936 2507 938 2535
rect 1072 2507 1074 2535
rect 719 2506 723 2507
rect 719 2501 723 2502
rect 807 2506 811 2507
rect 807 2501 811 2502
rect 847 2506 851 2507
rect 847 2501 851 2502
rect 935 2506 939 2507
rect 935 2501 939 2502
rect 983 2506 987 2507
rect 983 2501 987 2502
rect 1071 2506 1075 2507
rect 1071 2501 1075 2502
rect 1127 2506 1131 2507
rect 1127 2501 1131 2502
rect 720 2477 722 2501
rect 848 2477 850 2501
rect 984 2477 986 2501
rect 1128 2477 1130 2501
rect 718 2476 724 2477
rect 718 2472 719 2476
rect 723 2472 724 2476
rect 718 2471 724 2472
rect 846 2476 852 2477
rect 846 2472 847 2476
rect 851 2472 852 2476
rect 846 2471 852 2472
rect 982 2476 988 2477
rect 982 2472 983 2476
rect 987 2472 988 2476
rect 982 2471 988 2472
rect 1126 2476 1132 2477
rect 1126 2472 1127 2476
rect 1131 2472 1132 2476
rect 1126 2471 1132 2472
rect 578 2467 584 2468
rect 578 2463 579 2467
rect 583 2463 584 2467
rect 578 2462 584 2463
rect 682 2467 688 2468
rect 682 2463 683 2467
rect 687 2463 688 2467
rect 682 2462 688 2463
rect 702 2467 708 2468
rect 702 2463 703 2467
rect 707 2463 708 2467
rect 702 2462 708 2463
rect 922 2467 928 2468
rect 922 2463 923 2467
rect 927 2463 928 2467
rect 922 2462 928 2463
rect 930 2467 936 2468
rect 930 2463 931 2467
rect 935 2463 936 2467
rect 930 2462 936 2463
rect 1066 2467 1072 2468
rect 1066 2463 1067 2467
rect 1071 2463 1072 2467
rect 1066 2462 1072 2463
rect 502 2457 508 2458
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 502 2453 503 2457
rect 507 2453 508 2457
rect 502 2452 508 2453
rect 110 2451 116 2452
rect 112 2415 114 2451
rect 504 2415 506 2452
rect 580 2444 582 2462
rect 606 2457 612 2458
rect 606 2453 607 2457
rect 611 2453 612 2457
rect 606 2452 612 2453
rect 578 2443 584 2444
rect 578 2439 579 2443
rect 583 2439 584 2443
rect 578 2438 584 2439
rect 608 2415 610 2452
rect 684 2436 686 2462
rect 718 2457 724 2458
rect 718 2453 719 2457
rect 723 2453 724 2457
rect 718 2452 724 2453
rect 846 2457 852 2458
rect 846 2453 847 2457
rect 851 2453 852 2457
rect 846 2452 852 2453
rect 618 2435 624 2436
rect 618 2431 619 2435
rect 623 2431 624 2435
rect 618 2430 624 2431
rect 682 2435 688 2436
rect 682 2431 683 2435
rect 687 2431 688 2435
rect 682 2430 688 2431
rect 111 2414 115 2415
rect 111 2409 115 2410
rect 503 2414 507 2415
rect 503 2409 507 2410
rect 535 2414 539 2415
rect 535 2409 539 2410
rect 607 2414 611 2415
rect 607 2409 611 2410
rect 112 2389 114 2409
rect 110 2388 116 2389
rect 536 2388 538 2409
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 534 2387 540 2388
rect 534 2383 535 2387
rect 539 2383 540 2387
rect 534 2382 540 2383
rect 620 2380 622 2430
rect 720 2415 722 2452
rect 848 2415 850 2452
rect 924 2416 926 2462
rect 932 2436 934 2462
rect 982 2457 988 2458
rect 982 2453 983 2457
rect 987 2453 988 2457
rect 982 2452 988 2453
rect 930 2435 936 2436
rect 930 2431 931 2435
rect 935 2431 936 2435
rect 930 2430 936 2431
rect 922 2415 928 2416
rect 984 2415 986 2452
rect 1068 2436 1070 2462
rect 1126 2457 1132 2458
rect 1126 2453 1127 2457
rect 1131 2453 1132 2457
rect 1126 2452 1132 2453
rect 1066 2435 1072 2436
rect 1066 2431 1067 2435
rect 1071 2431 1072 2435
rect 1066 2430 1072 2431
rect 1128 2415 1130 2452
rect 1148 2436 1150 2542
rect 1206 2540 1212 2541
rect 1206 2536 1207 2540
rect 1211 2536 1212 2540
rect 1206 2535 1212 2536
rect 1350 2540 1356 2541
rect 1350 2536 1351 2540
rect 1355 2536 1356 2540
rect 1350 2535 1356 2536
rect 1208 2507 1210 2535
rect 1352 2507 1354 2535
rect 1207 2506 1211 2507
rect 1207 2501 1211 2502
rect 1279 2506 1283 2507
rect 1279 2501 1283 2502
rect 1351 2506 1355 2507
rect 1351 2501 1355 2502
rect 1280 2477 1282 2501
rect 1360 2499 1362 2574
rect 1496 2560 1498 2581
rect 1578 2579 1584 2580
rect 1578 2575 1579 2579
rect 1583 2575 1584 2579
rect 1578 2574 1584 2575
rect 1494 2559 1500 2560
rect 1494 2555 1495 2559
rect 1499 2555 1500 2559
rect 1494 2554 1500 2555
rect 1580 2552 1582 2574
rect 1648 2560 1650 2581
rect 1780 2580 1782 2634
rect 2006 2628 2012 2629
rect 2006 2624 2007 2628
rect 2011 2624 2012 2628
rect 2006 2623 2012 2624
rect 2008 2587 2010 2623
rect 2048 2615 2050 2643
rect 2096 2615 2098 2644
rect 2164 2628 2166 2754
rect 2198 2748 2204 2749
rect 2198 2744 2199 2748
rect 2203 2744 2204 2748
rect 2198 2743 2204 2744
rect 2342 2748 2348 2749
rect 2342 2744 2343 2748
rect 2347 2744 2348 2748
rect 2342 2743 2348 2744
rect 2200 2699 2202 2743
rect 2344 2699 2346 2743
rect 2199 2698 2203 2699
rect 2199 2693 2203 2694
rect 2263 2698 2267 2699
rect 2263 2693 2267 2694
rect 2343 2698 2347 2699
rect 2343 2693 2347 2694
rect 2264 2669 2266 2693
rect 2262 2668 2268 2669
rect 2262 2664 2263 2668
rect 2267 2664 2268 2668
rect 2262 2663 2268 2664
rect 2412 2660 2414 2782
rect 2420 2760 2422 2782
rect 2480 2768 2482 2789
rect 2554 2787 2560 2788
rect 2554 2783 2555 2787
rect 2559 2783 2560 2787
rect 2554 2782 2560 2783
rect 2478 2767 2484 2768
rect 2478 2763 2479 2767
rect 2483 2763 2484 2767
rect 2478 2762 2484 2763
rect 2556 2760 2558 2782
rect 2608 2768 2610 2789
rect 2606 2767 2612 2768
rect 2606 2763 2607 2767
rect 2611 2763 2612 2767
rect 2606 2762 2612 2763
rect 2684 2760 2686 2794
rect 2727 2789 2731 2790
rect 2839 2789 2843 2790
rect 2887 2794 2891 2795
rect 2887 2789 2891 2790
rect 2943 2794 2947 2795
rect 2962 2794 2968 2795
rect 3047 2794 3051 2795
rect 2943 2789 2947 2790
rect 3047 2789 3051 2790
rect 3095 2794 3099 2795
rect 3095 2789 3099 2790
rect 3143 2794 3147 2795
rect 3143 2789 3147 2790
rect 3239 2794 3243 2795
rect 3239 2789 3243 2790
rect 3287 2794 3291 2795
rect 3287 2789 3291 2790
rect 3343 2794 3347 2795
rect 3343 2789 3347 2790
rect 2728 2768 2730 2789
rect 2822 2787 2828 2788
rect 2822 2783 2823 2787
rect 2827 2783 2828 2787
rect 2822 2782 2828 2783
rect 2726 2767 2732 2768
rect 2726 2763 2727 2767
rect 2731 2763 2732 2767
rect 2726 2762 2732 2763
rect 2824 2760 2826 2782
rect 2840 2768 2842 2789
rect 2922 2779 2928 2780
rect 2922 2775 2923 2779
rect 2927 2775 2928 2779
rect 2922 2774 2928 2775
rect 2838 2767 2844 2768
rect 2838 2763 2839 2767
rect 2843 2763 2844 2767
rect 2838 2762 2844 2763
rect 2924 2760 2926 2774
rect 2944 2768 2946 2789
rect 3048 2768 3050 2789
rect 3130 2787 3136 2788
rect 3130 2783 3131 2787
rect 3135 2783 3136 2787
rect 3130 2782 3136 2783
rect 2942 2767 2948 2768
rect 2942 2763 2943 2767
rect 2947 2763 2948 2767
rect 2942 2762 2948 2763
rect 3046 2767 3052 2768
rect 3046 2763 3047 2767
rect 3051 2763 3052 2767
rect 3046 2762 3052 2763
rect 3132 2760 3134 2782
rect 3144 2768 3146 2789
rect 3240 2768 3242 2789
rect 3344 2768 3346 2789
rect 3356 2788 3358 2826
rect 3372 2800 3374 2826
rect 3478 2821 3484 2822
rect 3478 2817 3479 2821
rect 3483 2817 3484 2821
rect 3478 2816 3484 2817
rect 3670 2821 3676 2822
rect 3670 2817 3671 2821
rect 3675 2817 3676 2821
rect 3670 2816 3676 2817
rect 3370 2799 3376 2800
rect 3370 2795 3371 2799
rect 3375 2795 3376 2799
rect 3480 2795 3482 2816
rect 3522 2799 3528 2800
rect 3522 2795 3523 2799
rect 3527 2795 3528 2799
rect 3672 2795 3674 2816
rect 3756 2800 3758 2826
rect 3838 2821 3844 2822
rect 3838 2817 3839 2821
rect 3843 2817 3844 2821
rect 3838 2816 3844 2817
rect 3754 2799 3760 2800
rect 3754 2795 3755 2799
rect 3759 2795 3760 2799
rect 3840 2795 3842 2816
rect 3908 2800 3910 2831
rect 3942 2820 3948 2821
rect 3942 2816 3943 2820
rect 3947 2816 3948 2820
rect 3942 2815 3948 2816
rect 3906 2799 3912 2800
rect 3906 2795 3907 2799
rect 3911 2795 3912 2799
rect 3944 2795 3946 2815
rect 3370 2794 3376 2795
rect 3447 2794 3451 2795
rect 3447 2789 3451 2790
rect 3479 2794 3483 2795
rect 3522 2794 3528 2795
rect 3551 2794 3555 2795
rect 3479 2789 3483 2790
rect 3354 2787 3360 2788
rect 3354 2783 3355 2787
rect 3359 2783 3360 2787
rect 3354 2782 3360 2783
rect 3418 2787 3424 2788
rect 3418 2783 3419 2787
rect 3423 2783 3424 2787
rect 3418 2782 3424 2783
rect 3142 2767 3148 2768
rect 3142 2763 3143 2767
rect 3147 2763 3148 2767
rect 3142 2762 3148 2763
rect 3238 2767 3244 2768
rect 3238 2763 3239 2767
rect 3243 2763 3244 2767
rect 3238 2762 3244 2763
rect 3342 2767 3348 2768
rect 3342 2763 3343 2767
rect 3347 2763 3348 2767
rect 3342 2762 3348 2763
rect 3420 2760 3422 2782
rect 3448 2768 3450 2789
rect 3446 2767 3452 2768
rect 3446 2763 3447 2767
rect 3451 2763 3452 2767
rect 3446 2762 3452 2763
rect 3524 2760 3526 2794
rect 3551 2789 3555 2790
rect 3647 2794 3651 2795
rect 3647 2789 3651 2790
rect 3671 2794 3675 2795
rect 3671 2789 3675 2790
rect 3743 2794 3747 2795
rect 3754 2794 3760 2795
rect 3839 2794 3843 2795
rect 3906 2794 3912 2795
rect 3943 2794 3947 2795
rect 3743 2789 3747 2790
rect 3839 2789 3843 2790
rect 3943 2789 3947 2790
rect 3530 2779 3536 2780
rect 3530 2775 3531 2779
rect 3535 2775 3536 2779
rect 3530 2774 3536 2775
rect 3532 2760 3534 2774
rect 3552 2768 3554 2789
rect 3648 2768 3650 2789
rect 3744 2768 3746 2789
rect 3818 2787 3824 2788
rect 3818 2783 3819 2787
rect 3823 2783 3824 2787
rect 3818 2782 3824 2783
rect 3550 2767 3556 2768
rect 3550 2763 3551 2767
rect 3555 2763 3556 2767
rect 3550 2762 3556 2763
rect 3646 2767 3652 2768
rect 3646 2763 3647 2767
rect 3651 2763 3652 2767
rect 3646 2762 3652 2763
rect 3742 2767 3748 2768
rect 3742 2763 3743 2767
rect 3747 2763 3748 2767
rect 3742 2762 3748 2763
rect 3820 2760 3822 2782
rect 3826 2779 3832 2780
rect 3826 2775 3827 2779
rect 3831 2775 3832 2779
rect 3826 2774 3832 2775
rect 3828 2760 3830 2774
rect 3840 2768 3842 2789
rect 3944 2769 3946 2789
rect 3942 2768 3948 2769
rect 3838 2767 3844 2768
rect 3838 2763 3839 2767
rect 3843 2763 3844 2767
rect 3942 2764 3943 2768
rect 3947 2764 3948 2768
rect 3942 2763 3948 2764
rect 3838 2762 3844 2763
rect 2418 2759 2424 2760
rect 2418 2755 2419 2759
rect 2423 2755 2424 2759
rect 2418 2754 2424 2755
rect 2554 2759 2560 2760
rect 2554 2755 2555 2759
rect 2559 2755 2560 2759
rect 2554 2754 2560 2755
rect 2682 2759 2688 2760
rect 2682 2755 2683 2759
rect 2687 2755 2688 2759
rect 2682 2754 2688 2755
rect 2822 2759 2828 2760
rect 2822 2755 2823 2759
rect 2827 2755 2828 2759
rect 2922 2759 2928 2760
rect 2822 2754 2828 2755
rect 2914 2755 2920 2756
rect 2914 2751 2915 2755
rect 2919 2751 2920 2755
rect 2922 2755 2923 2759
rect 2927 2755 2928 2759
rect 2922 2754 2928 2755
rect 3130 2759 3136 2760
rect 3130 2755 3131 2759
rect 3135 2755 3136 2759
rect 3130 2754 3136 2755
rect 3418 2759 3424 2760
rect 3418 2755 3419 2759
rect 3423 2755 3424 2759
rect 3418 2754 3424 2755
rect 3522 2759 3528 2760
rect 3522 2755 3523 2759
rect 3527 2755 3528 2759
rect 3522 2754 3528 2755
rect 3530 2759 3536 2760
rect 3530 2755 3531 2759
rect 3535 2755 3536 2759
rect 3530 2754 3536 2755
rect 3818 2759 3824 2760
rect 3818 2755 3819 2759
rect 3823 2755 3824 2759
rect 3818 2754 3824 2755
rect 3826 2759 3832 2760
rect 3826 2755 3827 2759
rect 3831 2755 3832 2759
rect 3826 2754 3832 2755
rect 2914 2750 2920 2751
rect 3942 2751 3948 2752
rect 2478 2748 2484 2749
rect 2478 2744 2479 2748
rect 2483 2744 2484 2748
rect 2478 2743 2484 2744
rect 2606 2748 2612 2749
rect 2606 2744 2607 2748
rect 2611 2744 2612 2748
rect 2606 2743 2612 2744
rect 2726 2748 2732 2749
rect 2726 2744 2727 2748
rect 2731 2744 2732 2748
rect 2726 2743 2732 2744
rect 2838 2748 2844 2749
rect 2838 2744 2839 2748
rect 2843 2744 2844 2748
rect 2838 2743 2844 2744
rect 2480 2699 2482 2743
rect 2608 2699 2610 2743
rect 2728 2699 2730 2743
rect 2840 2699 2842 2743
rect 2439 2698 2443 2699
rect 2439 2693 2443 2694
rect 2479 2698 2483 2699
rect 2479 2693 2483 2694
rect 2607 2698 2611 2699
rect 2607 2693 2611 2694
rect 2615 2698 2619 2699
rect 2615 2693 2619 2694
rect 2727 2698 2731 2699
rect 2727 2693 2731 2694
rect 2783 2698 2787 2699
rect 2783 2693 2787 2694
rect 2839 2698 2843 2699
rect 2839 2693 2843 2694
rect 2440 2669 2442 2693
rect 2616 2669 2618 2693
rect 2784 2669 2786 2693
rect 2438 2668 2444 2669
rect 2438 2664 2439 2668
rect 2443 2664 2444 2668
rect 2438 2663 2444 2664
rect 2614 2668 2620 2669
rect 2614 2664 2615 2668
rect 2619 2664 2620 2668
rect 2614 2663 2620 2664
rect 2782 2668 2788 2669
rect 2782 2664 2783 2668
rect 2787 2664 2788 2668
rect 2782 2663 2788 2664
rect 2170 2659 2176 2660
rect 2170 2655 2171 2659
rect 2175 2655 2176 2659
rect 2170 2654 2176 2655
rect 2330 2659 2336 2660
rect 2330 2655 2331 2659
rect 2335 2655 2336 2659
rect 2330 2654 2336 2655
rect 2410 2659 2416 2660
rect 2410 2655 2411 2659
rect 2415 2655 2416 2659
rect 2410 2654 2416 2655
rect 2522 2659 2528 2660
rect 2522 2655 2523 2659
rect 2527 2655 2528 2659
rect 2522 2654 2528 2655
rect 2172 2628 2174 2654
rect 2262 2649 2268 2650
rect 2262 2645 2263 2649
rect 2267 2645 2268 2649
rect 2262 2644 2268 2645
rect 2162 2627 2168 2628
rect 2162 2623 2163 2627
rect 2167 2623 2168 2627
rect 2162 2622 2168 2623
rect 2170 2627 2176 2628
rect 2170 2623 2171 2627
rect 2175 2623 2176 2627
rect 2170 2622 2176 2623
rect 2264 2615 2266 2644
rect 2047 2614 2051 2615
rect 2047 2609 2051 2610
rect 2095 2614 2099 2615
rect 2095 2609 2099 2610
rect 2215 2614 2219 2615
rect 2215 2609 2219 2610
rect 2263 2614 2267 2615
rect 2263 2609 2267 2610
rect 2048 2589 2050 2609
rect 2046 2588 2052 2589
rect 2216 2588 2218 2609
rect 2332 2608 2334 2654
rect 2438 2649 2444 2650
rect 2438 2645 2439 2649
rect 2443 2645 2444 2649
rect 2438 2644 2444 2645
rect 2440 2615 2442 2644
rect 2524 2628 2526 2654
rect 2614 2649 2620 2650
rect 2614 2645 2615 2649
rect 2619 2645 2620 2649
rect 2614 2644 2620 2645
rect 2782 2649 2788 2650
rect 2782 2645 2783 2649
rect 2787 2645 2788 2649
rect 2782 2644 2788 2645
rect 2522 2627 2528 2628
rect 2522 2623 2523 2627
rect 2527 2623 2528 2627
rect 2522 2622 2528 2623
rect 2616 2615 2618 2644
rect 2746 2627 2752 2628
rect 2746 2623 2747 2627
rect 2751 2623 2752 2627
rect 2746 2622 2752 2623
rect 2367 2614 2371 2615
rect 2367 2609 2371 2610
rect 2439 2614 2443 2615
rect 2439 2609 2443 2610
rect 2519 2614 2523 2615
rect 2519 2609 2523 2610
rect 2615 2614 2619 2615
rect 2615 2609 2619 2610
rect 2671 2614 2675 2615
rect 2671 2609 2675 2610
rect 2330 2607 2336 2608
rect 2330 2603 2331 2607
rect 2335 2603 2336 2607
rect 2330 2602 2336 2603
rect 2368 2588 2370 2609
rect 2418 2607 2424 2608
rect 2418 2603 2419 2607
rect 2423 2603 2424 2607
rect 2418 2602 2424 2603
rect 2494 2607 2500 2608
rect 2494 2603 2495 2607
rect 2499 2603 2500 2607
rect 2494 2602 2500 2603
rect 1799 2586 1803 2587
rect 1799 2581 1803 2582
rect 2007 2586 2011 2587
rect 2046 2584 2047 2588
rect 2051 2584 2052 2588
rect 2046 2583 2052 2584
rect 2214 2587 2220 2588
rect 2214 2583 2215 2587
rect 2219 2583 2220 2587
rect 2214 2582 2220 2583
rect 2366 2587 2372 2588
rect 2366 2583 2367 2587
rect 2371 2583 2372 2587
rect 2366 2582 2372 2583
rect 2007 2581 2011 2582
rect 1730 2579 1736 2580
rect 1730 2575 1731 2579
rect 1735 2575 1736 2579
rect 1730 2574 1736 2575
rect 1778 2579 1784 2580
rect 1778 2575 1779 2579
rect 1783 2575 1784 2579
rect 1778 2574 1784 2575
rect 1646 2559 1652 2560
rect 1646 2555 1647 2559
rect 1651 2555 1652 2559
rect 1646 2554 1652 2555
rect 1732 2552 1734 2574
rect 1800 2560 1802 2581
rect 2008 2561 2010 2581
rect 2358 2575 2364 2576
rect 2046 2571 2052 2572
rect 2046 2567 2047 2571
rect 2051 2567 2052 2571
rect 2358 2571 2359 2575
rect 2363 2571 2364 2575
rect 2358 2570 2364 2571
rect 2046 2566 2052 2567
rect 2214 2568 2220 2569
rect 2006 2560 2012 2561
rect 1798 2559 1804 2560
rect 1798 2555 1799 2559
rect 1803 2555 1804 2559
rect 2006 2556 2007 2560
rect 2011 2556 2012 2560
rect 2006 2555 2012 2556
rect 1798 2554 1804 2555
rect 1578 2551 1584 2552
rect 1570 2547 1576 2548
rect 1570 2543 1571 2547
rect 1575 2543 1576 2547
rect 1578 2547 1579 2551
rect 1583 2547 1584 2551
rect 1578 2546 1584 2547
rect 1730 2551 1736 2552
rect 1730 2547 1731 2551
rect 1735 2547 1736 2551
rect 1730 2546 1736 2547
rect 1570 2542 1576 2543
rect 2006 2543 2012 2544
rect 1494 2540 1500 2541
rect 1494 2536 1495 2540
rect 1499 2536 1500 2540
rect 1494 2535 1500 2536
rect 1496 2507 1498 2535
rect 1431 2506 1435 2507
rect 1431 2501 1435 2502
rect 1495 2506 1499 2507
rect 1495 2501 1499 2502
rect 1356 2497 1362 2499
rect 1278 2476 1284 2477
rect 1278 2472 1279 2476
rect 1283 2472 1284 2476
rect 1278 2471 1284 2472
rect 1356 2468 1358 2497
rect 1432 2477 1434 2501
rect 1430 2476 1436 2477
rect 1430 2472 1431 2476
rect 1435 2472 1436 2476
rect 1430 2471 1436 2472
rect 1354 2467 1360 2468
rect 1354 2463 1355 2467
rect 1359 2463 1360 2467
rect 1354 2462 1360 2463
rect 1362 2467 1368 2468
rect 1362 2463 1363 2467
rect 1367 2463 1368 2467
rect 1362 2462 1368 2463
rect 1278 2457 1284 2458
rect 1278 2453 1279 2457
rect 1283 2453 1284 2457
rect 1278 2452 1284 2453
rect 1146 2435 1152 2436
rect 1146 2431 1147 2435
rect 1151 2431 1152 2435
rect 1146 2430 1152 2431
rect 1280 2415 1282 2452
rect 1364 2436 1366 2462
rect 1430 2457 1436 2458
rect 1430 2453 1431 2457
rect 1435 2453 1436 2457
rect 1430 2452 1436 2453
rect 1362 2435 1368 2436
rect 1362 2431 1363 2435
rect 1367 2431 1368 2435
rect 1362 2430 1368 2431
rect 1432 2415 1434 2452
rect 1572 2436 1574 2542
rect 1646 2540 1652 2541
rect 1646 2536 1647 2540
rect 1651 2536 1652 2540
rect 1646 2535 1652 2536
rect 1798 2540 1804 2541
rect 1798 2536 1799 2540
rect 1803 2536 1804 2540
rect 2006 2539 2007 2543
rect 2011 2539 2012 2543
rect 2006 2538 2012 2539
rect 1798 2535 1804 2536
rect 1648 2507 1650 2535
rect 1800 2507 1802 2535
rect 2008 2507 2010 2538
rect 2048 2535 2050 2566
rect 2214 2564 2215 2568
rect 2219 2564 2220 2568
rect 2214 2563 2220 2564
rect 2216 2535 2218 2563
rect 2047 2534 2051 2535
rect 2047 2529 2051 2530
rect 2095 2534 2099 2535
rect 2095 2529 2099 2530
rect 2215 2534 2219 2535
rect 2215 2529 2219 2530
rect 2343 2534 2347 2535
rect 2343 2529 2347 2530
rect 1583 2506 1587 2507
rect 1583 2501 1587 2502
rect 1647 2506 1651 2507
rect 1647 2501 1651 2502
rect 1743 2506 1747 2507
rect 1743 2501 1747 2502
rect 1799 2506 1803 2507
rect 1799 2501 1803 2502
rect 1903 2506 1907 2507
rect 1903 2501 1907 2502
rect 2007 2506 2011 2507
rect 2048 2502 2050 2529
rect 2096 2505 2098 2529
rect 2216 2505 2218 2529
rect 2344 2505 2346 2529
rect 2094 2504 2100 2505
rect 2007 2501 2011 2502
rect 2046 2501 2052 2502
rect 1584 2477 1586 2501
rect 1744 2477 1746 2501
rect 1904 2477 1906 2501
rect 1582 2476 1588 2477
rect 1582 2472 1583 2476
rect 1587 2472 1588 2476
rect 1582 2471 1588 2472
rect 1742 2476 1748 2477
rect 1742 2472 1743 2476
rect 1747 2472 1748 2476
rect 1742 2471 1748 2472
rect 1902 2476 1908 2477
rect 1902 2472 1903 2476
rect 1907 2472 1908 2476
rect 2008 2474 2010 2501
rect 2046 2497 2047 2501
rect 2051 2497 2052 2501
rect 2094 2500 2095 2504
rect 2099 2500 2100 2504
rect 2094 2499 2100 2500
rect 2214 2504 2220 2505
rect 2214 2500 2215 2504
rect 2219 2500 2220 2504
rect 2214 2499 2220 2500
rect 2342 2504 2348 2505
rect 2342 2500 2343 2504
rect 2347 2500 2348 2504
rect 2342 2499 2348 2500
rect 2046 2496 2052 2497
rect 2170 2495 2176 2496
rect 2170 2491 2171 2495
rect 2175 2491 2176 2495
rect 2170 2490 2176 2491
rect 2290 2495 2296 2496
rect 2290 2491 2291 2495
rect 2295 2491 2296 2495
rect 2290 2490 2296 2491
rect 2094 2485 2100 2486
rect 2046 2484 2052 2485
rect 2046 2480 2047 2484
rect 2051 2480 2052 2484
rect 2094 2481 2095 2485
rect 2099 2481 2100 2485
rect 2094 2480 2100 2481
rect 2046 2479 2052 2480
rect 1902 2471 1908 2472
rect 2006 2473 2012 2474
rect 2006 2469 2007 2473
rect 2011 2469 2012 2473
rect 2006 2468 2012 2469
rect 1658 2467 1664 2468
rect 1658 2463 1659 2467
rect 1663 2463 1664 2467
rect 1658 2462 1664 2463
rect 1818 2467 1824 2468
rect 1818 2463 1819 2467
rect 1823 2463 1824 2467
rect 1818 2462 1824 2463
rect 1970 2467 1976 2468
rect 1970 2463 1971 2467
rect 1975 2463 1976 2467
rect 1970 2462 1976 2463
rect 1582 2457 1588 2458
rect 1582 2453 1583 2457
rect 1587 2453 1588 2457
rect 1582 2452 1588 2453
rect 1570 2435 1576 2436
rect 1570 2431 1571 2435
rect 1575 2431 1576 2435
rect 1570 2430 1576 2431
rect 1584 2415 1586 2452
rect 1660 2436 1662 2462
rect 1742 2457 1748 2458
rect 1742 2453 1743 2457
rect 1747 2453 1748 2457
rect 1742 2452 1748 2453
rect 1658 2435 1664 2436
rect 1658 2431 1659 2435
rect 1663 2431 1664 2435
rect 1658 2430 1664 2431
rect 1744 2415 1746 2452
rect 1820 2436 1822 2462
rect 1902 2457 1908 2458
rect 1902 2453 1903 2457
rect 1907 2453 1908 2457
rect 1902 2452 1908 2453
rect 1818 2435 1824 2436
rect 1818 2431 1819 2435
rect 1823 2431 1824 2435
rect 1818 2430 1824 2431
rect 1904 2415 1906 2452
rect 671 2414 675 2415
rect 671 2409 675 2410
rect 719 2414 723 2415
rect 719 2409 723 2410
rect 815 2414 819 2415
rect 815 2409 819 2410
rect 847 2414 851 2415
rect 922 2411 923 2415
rect 927 2411 928 2415
rect 922 2410 928 2411
rect 959 2414 963 2415
rect 847 2409 851 2410
rect 959 2409 963 2410
rect 983 2414 987 2415
rect 983 2409 987 2410
rect 1103 2414 1107 2415
rect 1103 2409 1107 2410
rect 1127 2414 1131 2415
rect 1127 2409 1131 2410
rect 1247 2414 1251 2415
rect 1247 2409 1251 2410
rect 1279 2414 1283 2415
rect 1279 2409 1283 2410
rect 1391 2414 1395 2415
rect 1391 2409 1395 2410
rect 1431 2414 1435 2415
rect 1431 2409 1435 2410
rect 1527 2414 1531 2415
rect 1527 2409 1531 2410
rect 1583 2414 1587 2415
rect 1583 2409 1587 2410
rect 1655 2414 1659 2415
rect 1655 2409 1659 2410
rect 1743 2414 1747 2415
rect 1743 2409 1747 2410
rect 1791 2414 1795 2415
rect 1791 2409 1795 2410
rect 1903 2414 1907 2415
rect 1903 2409 1907 2410
rect 672 2388 674 2409
rect 730 2407 736 2408
rect 730 2403 731 2407
rect 735 2403 736 2407
rect 730 2402 736 2403
rect 670 2387 676 2388
rect 670 2383 671 2387
rect 675 2383 676 2387
rect 670 2382 676 2383
rect 618 2379 624 2380
rect 618 2375 619 2379
rect 623 2375 624 2379
rect 618 2374 624 2375
rect 110 2371 116 2372
rect 110 2367 111 2371
rect 115 2367 116 2371
rect 110 2366 116 2367
rect 534 2368 540 2369
rect 112 2335 114 2366
rect 534 2364 535 2368
rect 539 2364 540 2368
rect 534 2363 540 2364
rect 670 2368 676 2369
rect 670 2364 671 2368
rect 675 2364 676 2368
rect 670 2363 676 2364
rect 536 2335 538 2363
rect 672 2335 674 2363
rect 111 2334 115 2335
rect 111 2329 115 2330
rect 535 2334 539 2335
rect 535 2329 539 2330
rect 647 2334 651 2335
rect 647 2329 651 2330
rect 671 2334 675 2335
rect 671 2329 675 2330
rect 112 2302 114 2329
rect 536 2305 538 2329
rect 648 2305 650 2329
rect 534 2304 540 2305
rect 110 2301 116 2302
rect 110 2297 111 2301
rect 115 2297 116 2301
rect 534 2300 535 2304
rect 539 2300 540 2304
rect 534 2299 540 2300
rect 646 2304 652 2305
rect 646 2300 647 2304
rect 651 2300 652 2304
rect 646 2299 652 2300
rect 110 2296 116 2297
rect 732 2296 734 2402
rect 816 2388 818 2409
rect 960 2388 962 2409
rect 1034 2407 1040 2408
rect 1034 2403 1035 2407
rect 1039 2403 1040 2407
rect 1034 2402 1040 2403
rect 814 2387 820 2388
rect 814 2383 815 2387
rect 819 2383 820 2387
rect 814 2382 820 2383
rect 958 2387 964 2388
rect 958 2383 959 2387
rect 963 2383 964 2387
rect 958 2382 964 2383
rect 1036 2380 1038 2402
rect 1042 2399 1048 2400
rect 1042 2395 1043 2399
rect 1047 2395 1048 2399
rect 1042 2394 1048 2395
rect 1044 2380 1046 2394
rect 1104 2388 1106 2409
rect 1248 2388 1250 2409
rect 1322 2407 1328 2408
rect 1322 2403 1323 2407
rect 1327 2403 1328 2407
rect 1322 2402 1328 2403
rect 1102 2387 1108 2388
rect 1102 2383 1103 2387
rect 1107 2383 1108 2387
rect 1102 2382 1108 2383
rect 1246 2387 1252 2388
rect 1246 2383 1247 2387
rect 1251 2383 1252 2387
rect 1246 2382 1252 2383
rect 1324 2380 1326 2402
rect 1378 2399 1384 2400
rect 1378 2395 1379 2399
rect 1383 2395 1384 2399
rect 1378 2394 1384 2395
rect 1034 2379 1040 2380
rect 1034 2375 1035 2379
rect 1039 2375 1040 2379
rect 1034 2374 1040 2375
rect 1042 2379 1048 2380
rect 1042 2375 1043 2379
rect 1047 2375 1048 2379
rect 1042 2374 1048 2375
rect 1322 2379 1328 2380
rect 1322 2375 1323 2379
rect 1327 2375 1328 2379
rect 1322 2374 1328 2375
rect 882 2371 888 2372
rect 814 2368 820 2369
rect 814 2364 815 2368
rect 819 2364 820 2368
rect 882 2367 883 2371
rect 887 2367 888 2371
rect 882 2366 888 2367
rect 958 2368 964 2369
rect 814 2363 820 2364
rect 816 2335 818 2363
rect 767 2334 771 2335
rect 767 2329 771 2330
rect 815 2334 819 2335
rect 815 2329 819 2330
rect 768 2305 770 2329
rect 766 2304 772 2305
rect 766 2300 767 2304
rect 771 2300 772 2304
rect 766 2299 772 2300
rect 610 2295 616 2296
rect 610 2291 611 2295
rect 615 2291 616 2295
rect 610 2290 616 2291
rect 730 2295 736 2296
rect 730 2291 731 2295
rect 735 2291 736 2295
rect 730 2290 736 2291
rect 534 2285 540 2286
rect 110 2284 116 2285
rect 110 2280 111 2284
rect 115 2280 116 2284
rect 534 2281 535 2285
rect 539 2281 540 2285
rect 534 2280 540 2281
rect 110 2279 116 2280
rect 112 2255 114 2279
rect 490 2263 496 2264
rect 490 2259 491 2263
rect 495 2259 496 2263
rect 490 2258 496 2259
rect 111 2254 115 2255
rect 111 2249 115 2250
rect 415 2254 419 2255
rect 415 2249 419 2250
rect 112 2229 114 2249
rect 110 2228 116 2229
rect 416 2228 418 2249
rect 110 2224 111 2228
rect 115 2224 116 2228
rect 110 2223 116 2224
rect 414 2227 420 2228
rect 414 2223 415 2227
rect 419 2223 420 2227
rect 414 2222 420 2223
rect 492 2220 494 2258
rect 536 2255 538 2280
rect 612 2264 614 2290
rect 646 2285 652 2286
rect 646 2281 647 2285
rect 651 2281 652 2285
rect 646 2280 652 2281
rect 766 2285 772 2286
rect 766 2281 767 2285
rect 771 2281 772 2285
rect 766 2280 772 2281
rect 610 2263 616 2264
rect 610 2259 611 2263
rect 615 2259 616 2263
rect 610 2258 616 2259
rect 648 2255 650 2280
rect 768 2255 770 2280
rect 884 2264 886 2366
rect 958 2364 959 2368
rect 963 2364 964 2368
rect 958 2363 964 2364
rect 1102 2368 1108 2369
rect 1102 2364 1103 2368
rect 1107 2364 1108 2368
rect 1102 2363 1108 2364
rect 1246 2368 1252 2369
rect 1246 2364 1247 2368
rect 1251 2364 1252 2368
rect 1246 2363 1252 2364
rect 960 2335 962 2363
rect 1104 2335 1106 2363
rect 1248 2335 1250 2363
rect 895 2334 899 2335
rect 895 2329 899 2330
rect 959 2334 963 2335
rect 959 2329 963 2330
rect 1031 2334 1035 2335
rect 1031 2329 1035 2330
rect 1103 2334 1107 2335
rect 1103 2329 1107 2330
rect 1167 2334 1171 2335
rect 1167 2329 1171 2330
rect 1247 2334 1251 2335
rect 1247 2329 1251 2330
rect 1295 2334 1299 2335
rect 1295 2329 1299 2330
rect 896 2305 898 2329
rect 1032 2305 1034 2329
rect 1168 2305 1170 2329
rect 1296 2305 1298 2329
rect 894 2304 900 2305
rect 894 2300 895 2304
rect 899 2300 900 2304
rect 894 2299 900 2300
rect 1030 2304 1036 2305
rect 1030 2300 1031 2304
rect 1035 2300 1036 2304
rect 1030 2299 1036 2300
rect 1166 2304 1172 2305
rect 1166 2300 1167 2304
rect 1171 2300 1172 2304
rect 1166 2299 1172 2300
rect 1294 2304 1300 2305
rect 1294 2300 1295 2304
rect 1299 2300 1300 2304
rect 1294 2299 1300 2300
rect 1380 2296 1382 2394
rect 1392 2388 1394 2409
rect 1466 2407 1472 2408
rect 1466 2403 1467 2407
rect 1471 2403 1472 2407
rect 1466 2402 1472 2403
rect 1390 2387 1396 2388
rect 1390 2383 1391 2387
rect 1395 2383 1396 2387
rect 1390 2382 1396 2383
rect 1468 2380 1470 2402
rect 1528 2388 1530 2409
rect 1656 2388 1658 2409
rect 1730 2407 1736 2408
rect 1730 2403 1731 2407
rect 1735 2403 1736 2407
rect 1730 2402 1736 2403
rect 1526 2387 1532 2388
rect 1526 2383 1527 2387
rect 1531 2383 1532 2387
rect 1526 2382 1532 2383
rect 1654 2387 1660 2388
rect 1654 2383 1655 2387
rect 1659 2383 1660 2387
rect 1654 2382 1660 2383
rect 1732 2380 1734 2402
rect 1792 2388 1794 2409
rect 1874 2399 1880 2400
rect 1874 2395 1875 2399
rect 1879 2395 1880 2399
rect 1874 2394 1880 2395
rect 1790 2387 1796 2388
rect 1790 2383 1791 2387
rect 1795 2383 1796 2387
rect 1790 2382 1796 2383
rect 1876 2380 1878 2394
rect 1904 2388 1906 2409
rect 1972 2408 1974 2462
rect 2006 2456 2012 2457
rect 2006 2452 2007 2456
rect 2011 2452 2012 2456
rect 2006 2451 2012 2452
rect 2008 2415 2010 2451
rect 2048 2447 2050 2479
rect 2096 2447 2098 2480
rect 2172 2464 2174 2490
rect 2214 2485 2220 2486
rect 2214 2481 2215 2485
rect 2219 2481 2220 2485
rect 2214 2480 2220 2481
rect 2146 2463 2152 2464
rect 2146 2459 2147 2463
rect 2151 2459 2152 2463
rect 2146 2458 2152 2459
rect 2170 2463 2176 2464
rect 2170 2459 2171 2463
rect 2175 2459 2176 2463
rect 2170 2458 2176 2459
rect 2047 2446 2051 2447
rect 2047 2441 2051 2442
rect 2071 2446 2075 2447
rect 2071 2441 2075 2442
rect 2095 2446 2099 2447
rect 2095 2441 2099 2442
rect 2048 2421 2050 2441
rect 2046 2420 2052 2421
rect 2072 2420 2074 2441
rect 2046 2416 2047 2420
rect 2051 2416 2052 2420
rect 2046 2415 2052 2416
rect 2070 2419 2076 2420
rect 2070 2415 2071 2419
rect 2075 2415 2076 2419
rect 2007 2414 2011 2415
rect 2070 2414 2076 2415
rect 2148 2412 2150 2458
rect 2216 2447 2218 2480
rect 2292 2464 2294 2490
rect 2342 2485 2348 2486
rect 2342 2481 2343 2485
rect 2347 2481 2348 2485
rect 2342 2480 2348 2481
rect 2290 2463 2296 2464
rect 2290 2459 2291 2463
rect 2295 2459 2296 2463
rect 2290 2458 2296 2459
rect 2344 2447 2346 2480
rect 2360 2476 2362 2570
rect 2366 2568 2372 2569
rect 2366 2564 2367 2568
rect 2371 2564 2372 2568
rect 2366 2563 2372 2564
rect 2368 2535 2370 2563
rect 2367 2534 2371 2535
rect 2367 2529 2371 2530
rect 2420 2496 2422 2602
rect 2496 2580 2498 2602
rect 2520 2588 2522 2609
rect 2594 2607 2600 2608
rect 2594 2603 2595 2607
rect 2599 2603 2600 2607
rect 2594 2602 2600 2603
rect 2518 2587 2524 2588
rect 2518 2583 2519 2587
rect 2523 2583 2524 2587
rect 2518 2582 2524 2583
rect 2596 2580 2598 2602
rect 2672 2588 2674 2609
rect 2670 2587 2676 2588
rect 2670 2583 2671 2587
rect 2675 2583 2676 2587
rect 2670 2582 2676 2583
rect 2748 2580 2750 2622
rect 2784 2615 2786 2644
rect 2916 2628 2918 2750
rect 2942 2748 2948 2749
rect 2942 2744 2943 2748
rect 2947 2744 2948 2748
rect 2942 2743 2948 2744
rect 3046 2748 3052 2749
rect 3046 2744 3047 2748
rect 3051 2744 3052 2748
rect 3046 2743 3052 2744
rect 3142 2748 3148 2749
rect 3142 2744 3143 2748
rect 3147 2744 3148 2748
rect 3142 2743 3148 2744
rect 3238 2748 3244 2749
rect 3238 2744 3239 2748
rect 3243 2744 3244 2748
rect 3238 2743 3244 2744
rect 3342 2748 3348 2749
rect 3342 2744 3343 2748
rect 3347 2744 3348 2748
rect 3342 2743 3348 2744
rect 3446 2748 3452 2749
rect 3446 2744 3447 2748
rect 3451 2744 3452 2748
rect 3446 2743 3452 2744
rect 3550 2748 3556 2749
rect 3550 2744 3551 2748
rect 3555 2744 3556 2748
rect 3550 2743 3556 2744
rect 3646 2748 3652 2749
rect 3646 2744 3647 2748
rect 3651 2744 3652 2748
rect 3646 2743 3652 2744
rect 3742 2748 3748 2749
rect 3742 2744 3743 2748
rect 3747 2744 3748 2748
rect 3742 2743 3748 2744
rect 3838 2748 3844 2749
rect 3838 2744 3839 2748
rect 3843 2744 3844 2748
rect 3942 2747 3943 2751
rect 3947 2747 3948 2751
rect 3942 2746 3948 2747
rect 3838 2743 3844 2744
rect 2944 2699 2946 2743
rect 3048 2699 3050 2743
rect 3144 2699 3146 2743
rect 3240 2699 3242 2743
rect 3344 2699 3346 2743
rect 3448 2699 3450 2743
rect 3552 2699 3554 2743
rect 3648 2699 3650 2743
rect 3744 2699 3746 2743
rect 3840 2699 3842 2743
rect 3944 2699 3946 2746
rect 2943 2698 2947 2699
rect 2943 2693 2947 2694
rect 3047 2698 3051 2699
rect 3047 2693 3051 2694
rect 3095 2698 3099 2699
rect 3095 2693 3099 2694
rect 3143 2698 3147 2699
rect 3143 2693 3147 2694
rect 3239 2698 3243 2699
rect 3239 2693 3243 2694
rect 3343 2698 3347 2699
rect 3343 2693 3347 2694
rect 3383 2698 3387 2699
rect 3383 2693 3387 2694
rect 3447 2698 3451 2699
rect 3447 2693 3451 2694
rect 3535 2698 3539 2699
rect 3535 2693 3539 2694
rect 3551 2698 3555 2699
rect 3551 2693 3555 2694
rect 3647 2698 3651 2699
rect 3647 2693 3651 2694
rect 3743 2698 3747 2699
rect 3743 2693 3747 2694
rect 3839 2698 3843 2699
rect 3839 2693 3843 2694
rect 3943 2698 3947 2699
rect 3943 2693 3947 2694
rect 2944 2669 2946 2693
rect 3096 2669 3098 2693
rect 3240 2669 3242 2693
rect 3384 2669 3386 2693
rect 3536 2669 3538 2693
rect 2942 2668 2948 2669
rect 2942 2664 2943 2668
rect 2947 2664 2948 2668
rect 2942 2663 2948 2664
rect 3094 2668 3100 2669
rect 3094 2664 3095 2668
rect 3099 2664 3100 2668
rect 3094 2663 3100 2664
rect 3238 2668 3244 2669
rect 3238 2664 3239 2668
rect 3243 2664 3244 2668
rect 3238 2663 3244 2664
rect 3382 2668 3388 2669
rect 3382 2664 3383 2668
rect 3387 2664 3388 2668
rect 3382 2663 3388 2664
rect 3534 2668 3540 2669
rect 3534 2664 3535 2668
rect 3539 2664 3540 2668
rect 3944 2666 3946 2693
rect 3534 2663 3540 2664
rect 3942 2665 3948 2666
rect 3942 2661 3943 2665
rect 3947 2661 3948 2665
rect 3942 2660 3948 2661
rect 3018 2659 3024 2660
rect 3018 2655 3019 2659
rect 3023 2655 3024 2659
rect 3018 2654 3024 2655
rect 3170 2659 3176 2660
rect 3170 2655 3171 2659
rect 3175 2655 3176 2659
rect 3170 2654 3176 2655
rect 3314 2659 3320 2660
rect 3314 2655 3315 2659
rect 3319 2655 3320 2659
rect 3314 2654 3320 2655
rect 3458 2659 3464 2660
rect 3458 2655 3459 2659
rect 3463 2655 3464 2659
rect 3458 2654 3464 2655
rect 3466 2659 3472 2660
rect 3466 2655 3467 2659
rect 3471 2655 3472 2659
rect 3466 2654 3472 2655
rect 2942 2649 2948 2650
rect 2942 2645 2943 2649
rect 2947 2645 2948 2649
rect 2942 2644 2948 2645
rect 2914 2627 2920 2628
rect 2914 2623 2915 2627
rect 2919 2623 2920 2627
rect 2914 2622 2920 2623
rect 2944 2615 2946 2644
rect 3020 2628 3022 2654
rect 3094 2649 3100 2650
rect 3094 2645 3095 2649
rect 3099 2645 3100 2649
rect 3094 2644 3100 2645
rect 3018 2627 3024 2628
rect 3018 2623 3019 2627
rect 3023 2623 3024 2627
rect 3018 2622 3024 2623
rect 3096 2615 3098 2644
rect 3172 2628 3174 2654
rect 3238 2649 3244 2650
rect 3238 2645 3239 2649
rect 3243 2645 3244 2649
rect 3238 2644 3244 2645
rect 3170 2627 3176 2628
rect 3170 2623 3171 2627
rect 3175 2623 3176 2627
rect 3170 2622 3176 2623
rect 3240 2615 3242 2644
rect 3316 2628 3318 2654
rect 3382 2649 3388 2650
rect 3382 2645 3383 2649
rect 3387 2645 3388 2649
rect 3382 2644 3388 2645
rect 3314 2627 3320 2628
rect 3314 2623 3315 2627
rect 3319 2623 3320 2627
rect 3314 2622 3320 2623
rect 3384 2615 3386 2644
rect 3460 2628 3462 2654
rect 3458 2627 3464 2628
rect 3458 2623 3459 2627
rect 3463 2623 3464 2627
rect 3458 2622 3464 2623
rect 2783 2614 2787 2615
rect 2783 2609 2787 2610
rect 2815 2614 2819 2615
rect 2815 2609 2819 2610
rect 2943 2614 2947 2615
rect 2943 2609 2947 2610
rect 2951 2614 2955 2615
rect 2951 2609 2955 2610
rect 3087 2614 3091 2615
rect 3087 2609 3091 2610
rect 3095 2614 3099 2615
rect 3095 2609 3099 2610
rect 3223 2614 3227 2615
rect 3223 2609 3227 2610
rect 3239 2614 3243 2615
rect 3239 2609 3243 2610
rect 3367 2614 3371 2615
rect 3367 2609 3371 2610
rect 3383 2614 3387 2615
rect 3383 2609 3387 2610
rect 2816 2588 2818 2609
rect 2952 2588 2954 2609
rect 3034 2607 3040 2608
rect 3034 2603 3035 2607
rect 3039 2603 3040 2607
rect 3034 2602 3040 2603
rect 2814 2587 2820 2588
rect 2814 2583 2815 2587
rect 2819 2583 2820 2587
rect 2814 2582 2820 2583
rect 2950 2587 2956 2588
rect 2950 2583 2951 2587
rect 2955 2583 2956 2587
rect 2950 2582 2956 2583
rect 3036 2580 3038 2602
rect 3088 2588 3090 2609
rect 3170 2607 3176 2608
rect 3170 2603 3171 2607
rect 3175 2603 3176 2607
rect 3170 2602 3176 2603
rect 3086 2587 3092 2588
rect 3086 2583 3087 2587
rect 3091 2583 3092 2587
rect 3086 2582 3092 2583
rect 3172 2580 3174 2602
rect 3224 2588 3226 2609
rect 3306 2607 3312 2608
rect 3306 2603 3307 2607
rect 3311 2603 3312 2607
rect 3306 2602 3312 2603
rect 3222 2587 3228 2588
rect 3222 2583 3223 2587
rect 3227 2583 3228 2587
rect 3222 2582 3228 2583
rect 3308 2580 3310 2602
rect 3368 2588 3370 2609
rect 3468 2608 3470 2654
rect 3534 2649 3540 2650
rect 3534 2645 3535 2649
rect 3539 2645 3540 2649
rect 3534 2644 3540 2645
rect 3942 2648 3948 2649
rect 3942 2644 3943 2648
rect 3947 2644 3948 2648
rect 3536 2615 3538 2644
rect 3942 2643 3948 2644
rect 3944 2615 3946 2643
rect 3535 2614 3539 2615
rect 3535 2609 3539 2610
rect 3943 2614 3947 2615
rect 3943 2609 3947 2610
rect 3466 2607 3472 2608
rect 3466 2603 3467 2607
rect 3471 2603 3472 2607
rect 3466 2602 3472 2603
rect 3944 2589 3946 2609
rect 3942 2588 3948 2589
rect 3366 2587 3372 2588
rect 3366 2583 3367 2587
rect 3371 2583 3372 2587
rect 3942 2584 3943 2588
rect 3947 2584 3948 2588
rect 3942 2583 3948 2584
rect 3366 2582 3372 2583
rect 2494 2579 2500 2580
rect 2494 2575 2495 2579
rect 2499 2575 2500 2579
rect 2494 2574 2500 2575
rect 2594 2579 2600 2580
rect 2594 2575 2595 2579
rect 2599 2575 2600 2579
rect 2594 2574 2600 2575
rect 2746 2579 2752 2580
rect 2746 2575 2747 2579
rect 2751 2575 2752 2579
rect 2746 2574 2752 2575
rect 2786 2579 2792 2580
rect 2786 2575 2787 2579
rect 2791 2575 2792 2579
rect 2786 2574 2792 2575
rect 3034 2579 3040 2580
rect 3034 2575 3035 2579
rect 3039 2575 3040 2579
rect 3034 2574 3040 2575
rect 3170 2579 3176 2580
rect 3170 2575 3171 2579
rect 3175 2575 3176 2579
rect 3170 2574 3176 2575
rect 3306 2579 3312 2580
rect 3306 2575 3307 2579
rect 3311 2575 3312 2579
rect 3306 2574 3312 2575
rect 2518 2568 2524 2569
rect 2518 2564 2519 2568
rect 2523 2564 2524 2568
rect 2518 2563 2524 2564
rect 2670 2568 2676 2569
rect 2670 2564 2671 2568
rect 2675 2564 2676 2568
rect 2670 2563 2676 2564
rect 2520 2535 2522 2563
rect 2672 2535 2674 2563
rect 2471 2534 2475 2535
rect 2471 2529 2475 2530
rect 2519 2534 2523 2535
rect 2519 2529 2523 2530
rect 2599 2534 2603 2535
rect 2599 2529 2603 2530
rect 2671 2534 2675 2535
rect 2671 2529 2675 2530
rect 2719 2534 2723 2535
rect 2719 2529 2723 2530
rect 2472 2505 2474 2529
rect 2600 2505 2602 2529
rect 2720 2505 2722 2529
rect 2470 2504 2476 2505
rect 2470 2500 2471 2504
rect 2475 2500 2476 2504
rect 2470 2499 2476 2500
rect 2598 2504 2604 2505
rect 2598 2500 2599 2504
rect 2603 2500 2604 2504
rect 2598 2499 2604 2500
rect 2718 2504 2724 2505
rect 2718 2500 2719 2504
rect 2723 2500 2724 2504
rect 2718 2499 2724 2500
rect 2418 2495 2424 2496
rect 2418 2491 2419 2495
rect 2423 2491 2424 2495
rect 2418 2490 2424 2491
rect 2546 2495 2552 2496
rect 2546 2491 2547 2495
rect 2551 2491 2552 2495
rect 2546 2490 2552 2491
rect 2666 2495 2672 2496
rect 2666 2491 2667 2495
rect 2671 2491 2672 2495
rect 2666 2490 2672 2491
rect 2470 2485 2476 2486
rect 2470 2481 2471 2485
rect 2475 2481 2476 2485
rect 2470 2480 2476 2481
rect 2358 2475 2364 2476
rect 2358 2471 2359 2475
rect 2363 2471 2364 2475
rect 2358 2470 2364 2471
rect 2472 2447 2474 2480
rect 2548 2464 2550 2490
rect 2598 2485 2604 2486
rect 2598 2481 2599 2485
rect 2603 2481 2604 2485
rect 2598 2480 2604 2481
rect 2546 2463 2552 2464
rect 2546 2459 2547 2463
rect 2551 2459 2552 2463
rect 2546 2458 2552 2459
rect 2600 2447 2602 2480
rect 2191 2446 2195 2447
rect 2191 2441 2195 2442
rect 2215 2446 2219 2447
rect 2215 2441 2219 2442
rect 2319 2446 2323 2447
rect 2319 2441 2323 2442
rect 2343 2446 2347 2447
rect 2343 2441 2347 2442
rect 2439 2446 2443 2447
rect 2439 2441 2443 2442
rect 2471 2446 2475 2447
rect 2471 2441 2475 2442
rect 2559 2446 2563 2447
rect 2559 2441 2563 2442
rect 2599 2446 2603 2447
rect 2599 2441 2603 2442
rect 2192 2420 2194 2441
rect 2242 2439 2248 2440
rect 2242 2435 2243 2439
rect 2247 2435 2248 2439
rect 2242 2434 2248 2435
rect 2266 2439 2272 2440
rect 2266 2435 2267 2439
rect 2271 2435 2272 2439
rect 2266 2434 2272 2435
rect 2190 2419 2196 2420
rect 2190 2415 2191 2419
rect 2195 2415 2196 2419
rect 2190 2414 2196 2415
rect 2007 2409 2011 2410
rect 2146 2411 2152 2412
rect 1970 2407 1976 2408
rect 1970 2403 1971 2407
rect 1975 2403 1976 2407
rect 1970 2402 1976 2403
rect 2008 2389 2010 2409
rect 2146 2407 2147 2411
rect 2151 2407 2152 2411
rect 2146 2406 2152 2407
rect 2046 2403 2052 2404
rect 2046 2399 2047 2403
rect 2051 2399 2052 2403
rect 2046 2398 2052 2399
rect 2070 2400 2076 2401
rect 2006 2388 2012 2389
rect 1902 2387 1908 2388
rect 1902 2383 1903 2387
rect 1907 2383 1908 2387
rect 2006 2384 2007 2388
rect 2011 2384 2012 2388
rect 2006 2383 2012 2384
rect 1902 2382 1908 2383
rect 1466 2379 1472 2380
rect 1466 2375 1467 2379
rect 1471 2375 1472 2379
rect 1466 2374 1472 2375
rect 1730 2379 1736 2380
rect 1730 2375 1731 2379
rect 1735 2375 1736 2379
rect 1874 2379 1880 2380
rect 1730 2374 1736 2375
rect 1866 2375 1872 2376
rect 1866 2371 1867 2375
rect 1871 2371 1872 2375
rect 1874 2375 1875 2379
rect 1879 2375 1880 2379
rect 1874 2374 1880 2375
rect 1866 2370 1872 2371
rect 2006 2371 2012 2372
rect 1390 2368 1396 2369
rect 1390 2364 1391 2368
rect 1395 2364 1396 2368
rect 1390 2363 1396 2364
rect 1526 2368 1532 2369
rect 1526 2364 1527 2368
rect 1531 2364 1532 2368
rect 1526 2363 1532 2364
rect 1654 2368 1660 2369
rect 1654 2364 1655 2368
rect 1659 2364 1660 2368
rect 1654 2363 1660 2364
rect 1790 2368 1796 2369
rect 1790 2364 1791 2368
rect 1795 2364 1796 2368
rect 1790 2363 1796 2364
rect 1392 2335 1394 2363
rect 1528 2335 1530 2363
rect 1656 2335 1658 2363
rect 1792 2335 1794 2363
rect 1391 2334 1395 2335
rect 1391 2329 1395 2330
rect 1423 2334 1427 2335
rect 1423 2329 1427 2330
rect 1527 2334 1531 2335
rect 1527 2329 1531 2330
rect 1551 2334 1555 2335
rect 1551 2329 1555 2330
rect 1655 2334 1659 2335
rect 1655 2329 1659 2330
rect 1671 2334 1675 2335
rect 1671 2329 1675 2330
rect 1791 2334 1795 2335
rect 1791 2329 1795 2330
rect 1799 2334 1803 2335
rect 1799 2329 1803 2330
rect 1424 2305 1426 2329
rect 1552 2305 1554 2329
rect 1672 2305 1674 2329
rect 1800 2305 1802 2329
rect 1422 2304 1428 2305
rect 1422 2300 1423 2304
rect 1427 2300 1428 2304
rect 1422 2299 1428 2300
rect 1550 2304 1556 2305
rect 1550 2300 1551 2304
rect 1555 2300 1556 2304
rect 1550 2299 1556 2300
rect 1670 2304 1676 2305
rect 1670 2300 1671 2304
rect 1675 2300 1676 2304
rect 1670 2299 1676 2300
rect 1798 2304 1804 2305
rect 1798 2300 1799 2304
rect 1803 2300 1804 2304
rect 1798 2299 1804 2300
rect 970 2295 976 2296
rect 970 2291 971 2295
rect 975 2291 976 2295
rect 970 2290 976 2291
rect 1106 2295 1112 2296
rect 1106 2291 1107 2295
rect 1111 2291 1112 2295
rect 1106 2290 1112 2291
rect 1114 2295 1120 2296
rect 1114 2291 1115 2295
rect 1119 2291 1120 2295
rect 1114 2290 1120 2291
rect 1370 2295 1376 2296
rect 1370 2291 1371 2295
rect 1375 2291 1376 2295
rect 1370 2290 1376 2291
rect 1378 2295 1384 2296
rect 1378 2291 1379 2295
rect 1383 2291 1384 2295
rect 1378 2290 1384 2291
rect 1506 2295 1512 2296
rect 1506 2291 1507 2295
rect 1511 2291 1512 2295
rect 1506 2290 1512 2291
rect 1634 2295 1640 2296
rect 1634 2291 1635 2295
rect 1639 2291 1640 2295
rect 1634 2290 1640 2291
rect 894 2285 900 2286
rect 894 2281 895 2285
rect 899 2281 900 2285
rect 894 2280 900 2281
rect 882 2263 888 2264
rect 882 2259 883 2263
rect 887 2259 888 2263
rect 882 2258 888 2259
rect 896 2255 898 2280
rect 972 2264 974 2290
rect 1030 2285 1036 2286
rect 1030 2281 1031 2285
rect 1035 2281 1036 2285
rect 1030 2280 1036 2281
rect 970 2263 976 2264
rect 970 2259 971 2263
rect 975 2259 976 2263
rect 970 2258 976 2259
rect 1032 2255 1034 2280
rect 1108 2264 1110 2290
rect 1106 2263 1112 2264
rect 1106 2259 1107 2263
rect 1111 2259 1112 2263
rect 1106 2258 1112 2259
rect 1116 2256 1118 2290
rect 1166 2285 1172 2286
rect 1166 2281 1167 2285
rect 1171 2281 1172 2285
rect 1166 2280 1172 2281
rect 1294 2285 1300 2286
rect 1294 2281 1295 2285
rect 1299 2281 1300 2285
rect 1294 2280 1300 2281
rect 1114 2255 1120 2256
rect 1168 2255 1170 2280
rect 1296 2255 1298 2280
rect 1372 2264 1374 2290
rect 1422 2285 1428 2286
rect 1422 2281 1423 2285
rect 1427 2281 1428 2285
rect 1422 2280 1428 2281
rect 1370 2263 1376 2264
rect 1370 2259 1371 2263
rect 1375 2259 1376 2263
rect 1370 2258 1376 2259
rect 1424 2255 1426 2280
rect 1508 2272 1510 2290
rect 1550 2285 1556 2286
rect 1550 2281 1551 2285
rect 1555 2281 1556 2285
rect 1550 2280 1556 2281
rect 1506 2271 1512 2272
rect 1506 2267 1507 2271
rect 1511 2267 1512 2271
rect 1506 2266 1512 2267
rect 1552 2255 1554 2280
rect 1636 2264 1638 2290
rect 1670 2285 1676 2286
rect 1670 2281 1671 2285
rect 1675 2281 1676 2285
rect 1670 2280 1676 2281
rect 1798 2285 1804 2286
rect 1798 2281 1799 2285
rect 1803 2281 1804 2285
rect 1798 2280 1804 2281
rect 1634 2263 1640 2264
rect 1634 2259 1635 2263
rect 1639 2259 1640 2263
rect 1634 2258 1640 2259
rect 1642 2263 1648 2264
rect 1642 2259 1643 2263
rect 1647 2259 1648 2263
rect 1642 2258 1648 2259
rect 535 2254 539 2255
rect 535 2249 539 2250
rect 647 2254 651 2255
rect 647 2249 651 2250
rect 671 2254 675 2255
rect 671 2249 675 2250
rect 767 2254 771 2255
rect 767 2249 771 2250
rect 823 2254 827 2255
rect 823 2249 827 2250
rect 895 2254 899 2255
rect 895 2249 899 2250
rect 991 2254 995 2255
rect 991 2249 995 2250
rect 1031 2254 1035 2255
rect 1114 2251 1115 2255
rect 1119 2251 1120 2255
rect 1114 2250 1120 2251
rect 1167 2254 1171 2255
rect 1031 2249 1035 2250
rect 1167 2249 1171 2250
rect 1175 2254 1179 2255
rect 1175 2249 1179 2250
rect 1295 2254 1299 2255
rect 1295 2249 1299 2250
rect 1367 2254 1371 2255
rect 1367 2249 1371 2250
rect 1423 2254 1427 2255
rect 1423 2249 1427 2250
rect 1551 2254 1555 2255
rect 1551 2249 1555 2250
rect 1567 2254 1571 2255
rect 1567 2249 1571 2250
rect 498 2247 504 2248
rect 498 2243 499 2247
rect 503 2243 504 2247
rect 498 2242 504 2243
rect 500 2220 502 2242
rect 536 2228 538 2249
rect 618 2247 624 2248
rect 618 2243 619 2247
rect 623 2243 624 2247
rect 618 2242 624 2243
rect 534 2227 540 2228
rect 534 2223 535 2227
rect 539 2223 540 2227
rect 534 2222 540 2223
rect 620 2220 622 2242
rect 672 2228 674 2249
rect 778 2247 784 2248
rect 778 2243 779 2247
rect 783 2243 784 2247
rect 778 2242 784 2243
rect 670 2227 676 2228
rect 670 2223 671 2227
rect 675 2223 676 2227
rect 670 2222 676 2223
rect 490 2219 496 2220
rect 490 2215 491 2219
rect 495 2215 496 2219
rect 490 2214 496 2215
rect 498 2219 504 2220
rect 498 2215 499 2219
rect 503 2215 504 2219
rect 498 2214 504 2215
rect 618 2219 624 2220
rect 618 2215 619 2219
rect 623 2215 624 2219
rect 618 2214 624 2215
rect 110 2211 116 2212
rect 110 2207 111 2211
rect 115 2207 116 2211
rect 110 2206 116 2207
rect 414 2208 420 2209
rect 112 2171 114 2206
rect 414 2204 415 2208
rect 419 2204 420 2208
rect 414 2203 420 2204
rect 534 2208 540 2209
rect 534 2204 535 2208
rect 539 2204 540 2208
rect 534 2203 540 2204
rect 670 2208 676 2209
rect 670 2204 671 2208
rect 675 2204 676 2208
rect 670 2203 676 2204
rect 416 2171 418 2203
rect 536 2171 538 2203
rect 672 2171 674 2203
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 135 2170 139 2171
rect 135 2165 139 2166
rect 247 2170 251 2171
rect 247 2165 251 2166
rect 391 2170 395 2171
rect 391 2165 395 2166
rect 415 2170 419 2171
rect 415 2165 419 2166
rect 535 2170 539 2171
rect 535 2165 539 2166
rect 551 2170 555 2171
rect 551 2165 555 2166
rect 671 2170 675 2171
rect 671 2165 675 2166
rect 711 2170 715 2171
rect 711 2165 715 2166
rect 112 2138 114 2165
rect 136 2141 138 2165
rect 248 2141 250 2165
rect 392 2141 394 2165
rect 552 2141 554 2165
rect 712 2141 714 2165
rect 134 2140 140 2141
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 246 2140 252 2141
rect 246 2136 247 2140
rect 251 2136 252 2140
rect 246 2135 252 2136
rect 390 2140 396 2141
rect 390 2136 391 2140
rect 395 2136 396 2140
rect 390 2135 396 2136
rect 550 2140 556 2141
rect 550 2136 551 2140
rect 555 2136 556 2140
rect 550 2135 556 2136
rect 710 2140 716 2141
rect 710 2136 711 2140
rect 715 2136 716 2140
rect 710 2135 716 2136
rect 110 2132 116 2133
rect 780 2132 782 2242
rect 824 2228 826 2249
rect 992 2228 994 2249
rect 1066 2247 1072 2248
rect 1066 2243 1067 2247
rect 1071 2243 1072 2247
rect 1066 2242 1072 2243
rect 822 2227 828 2228
rect 822 2223 823 2227
rect 827 2223 828 2227
rect 822 2222 828 2223
rect 990 2227 996 2228
rect 990 2223 991 2227
rect 995 2223 996 2227
rect 990 2222 996 2223
rect 1068 2220 1070 2242
rect 1176 2228 1178 2249
rect 1250 2247 1256 2248
rect 1250 2243 1251 2247
rect 1255 2243 1256 2247
rect 1250 2242 1256 2243
rect 1174 2227 1180 2228
rect 1174 2223 1175 2227
rect 1179 2223 1180 2227
rect 1174 2222 1180 2223
rect 1252 2220 1254 2242
rect 1368 2228 1370 2249
rect 1568 2228 1570 2249
rect 1366 2227 1372 2228
rect 1366 2223 1367 2227
rect 1371 2223 1372 2227
rect 1366 2222 1372 2223
rect 1566 2227 1572 2228
rect 1566 2223 1567 2227
rect 1571 2223 1572 2227
rect 1566 2222 1572 2223
rect 1644 2220 1646 2258
rect 1672 2255 1674 2280
rect 1800 2255 1802 2280
rect 1868 2264 1870 2370
rect 1902 2368 1908 2369
rect 1902 2364 1903 2368
rect 1907 2364 1908 2368
rect 2006 2367 2007 2371
rect 2011 2367 2012 2371
rect 2048 2367 2050 2398
rect 2070 2396 2071 2400
rect 2075 2396 2076 2400
rect 2070 2395 2076 2396
rect 2190 2400 2196 2401
rect 2190 2396 2191 2400
rect 2195 2396 2196 2400
rect 2190 2395 2196 2396
rect 2072 2367 2074 2395
rect 2192 2367 2194 2395
rect 2006 2366 2012 2367
rect 2047 2366 2051 2367
rect 1902 2363 1908 2364
rect 1904 2335 1906 2363
rect 2008 2335 2010 2366
rect 2047 2361 2051 2362
rect 2071 2366 2075 2367
rect 2071 2361 2075 2362
rect 2167 2366 2171 2367
rect 2167 2361 2171 2362
rect 2191 2366 2195 2367
rect 2191 2361 2195 2362
rect 1903 2334 1907 2335
rect 1903 2329 1907 2330
rect 2007 2334 2011 2335
rect 2048 2334 2050 2361
rect 2168 2337 2170 2361
rect 2166 2336 2172 2337
rect 2007 2329 2011 2330
rect 2046 2333 2052 2334
rect 2046 2329 2047 2333
rect 2051 2329 2052 2333
rect 2166 2332 2167 2336
rect 2171 2332 2172 2336
rect 2166 2331 2172 2332
rect 1904 2305 1906 2329
rect 1902 2304 1908 2305
rect 1902 2300 1903 2304
rect 1907 2300 1908 2304
rect 2008 2302 2010 2329
rect 2046 2328 2052 2329
rect 2244 2328 2246 2434
rect 2268 2412 2270 2434
rect 2274 2431 2280 2432
rect 2274 2427 2275 2431
rect 2279 2427 2280 2431
rect 2274 2426 2280 2427
rect 2276 2412 2278 2426
rect 2320 2420 2322 2441
rect 2440 2420 2442 2441
rect 2522 2439 2528 2440
rect 2522 2435 2523 2439
rect 2527 2435 2528 2439
rect 2522 2434 2528 2435
rect 2318 2419 2324 2420
rect 2318 2415 2319 2419
rect 2323 2415 2324 2419
rect 2318 2414 2324 2415
rect 2438 2419 2444 2420
rect 2438 2415 2439 2419
rect 2443 2415 2444 2419
rect 2438 2414 2444 2415
rect 2524 2412 2526 2434
rect 2560 2420 2562 2441
rect 2668 2440 2670 2490
rect 2718 2485 2724 2486
rect 2718 2481 2719 2485
rect 2723 2481 2724 2485
rect 2718 2480 2724 2481
rect 2720 2447 2722 2480
rect 2788 2464 2790 2574
rect 3942 2571 3948 2572
rect 2814 2568 2820 2569
rect 2814 2564 2815 2568
rect 2819 2564 2820 2568
rect 2814 2563 2820 2564
rect 2950 2568 2956 2569
rect 2950 2564 2951 2568
rect 2955 2564 2956 2568
rect 2950 2563 2956 2564
rect 3086 2568 3092 2569
rect 3086 2564 3087 2568
rect 3091 2564 3092 2568
rect 3086 2563 3092 2564
rect 3222 2568 3228 2569
rect 3222 2564 3223 2568
rect 3227 2564 3228 2568
rect 3222 2563 3228 2564
rect 3366 2568 3372 2569
rect 3366 2564 3367 2568
rect 3371 2564 3372 2568
rect 3942 2567 3943 2571
rect 3947 2567 3948 2571
rect 3942 2566 3948 2567
rect 3366 2563 3372 2564
rect 2816 2535 2818 2563
rect 2952 2535 2954 2563
rect 3088 2535 3090 2563
rect 3224 2535 3226 2563
rect 3368 2535 3370 2563
rect 3944 2535 3946 2566
rect 2815 2534 2819 2535
rect 2815 2529 2819 2530
rect 2839 2534 2843 2535
rect 2839 2529 2843 2530
rect 2951 2534 2955 2535
rect 2951 2529 2955 2530
rect 2967 2534 2971 2535
rect 2967 2529 2971 2530
rect 3087 2534 3091 2535
rect 3087 2529 3091 2530
rect 3095 2534 3099 2535
rect 3095 2529 3099 2530
rect 3223 2534 3227 2535
rect 3223 2529 3227 2530
rect 3367 2534 3371 2535
rect 3367 2529 3371 2530
rect 3943 2534 3947 2535
rect 3943 2529 3947 2530
rect 2840 2505 2842 2529
rect 2968 2505 2970 2529
rect 3096 2505 3098 2529
rect 3224 2505 3226 2529
rect 2838 2504 2844 2505
rect 2838 2500 2839 2504
rect 2843 2500 2844 2504
rect 2838 2499 2844 2500
rect 2966 2504 2972 2505
rect 2966 2500 2967 2504
rect 2971 2500 2972 2504
rect 2966 2499 2972 2500
rect 3094 2504 3100 2505
rect 3094 2500 3095 2504
rect 3099 2500 3100 2504
rect 3094 2499 3100 2500
rect 3222 2504 3228 2505
rect 3222 2500 3223 2504
rect 3227 2500 3228 2504
rect 3944 2502 3946 2529
rect 3222 2499 3228 2500
rect 3942 2501 3948 2502
rect 3942 2497 3943 2501
rect 3947 2497 3948 2501
rect 3942 2496 3948 2497
rect 2794 2495 2800 2496
rect 2794 2491 2795 2495
rect 2799 2491 2800 2495
rect 2794 2490 2800 2491
rect 2914 2495 2920 2496
rect 2914 2491 2915 2495
rect 2919 2491 2920 2495
rect 2914 2490 2920 2491
rect 3042 2495 3048 2496
rect 3042 2491 3043 2495
rect 3047 2491 3048 2495
rect 3042 2490 3048 2491
rect 3170 2495 3176 2496
rect 3170 2491 3171 2495
rect 3175 2491 3176 2495
rect 3170 2490 3176 2491
rect 3214 2495 3220 2496
rect 3214 2491 3215 2495
rect 3219 2491 3220 2495
rect 3214 2490 3220 2491
rect 2796 2464 2798 2490
rect 2838 2485 2844 2486
rect 2838 2481 2839 2485
rect 2843 2481 2844 2485
rect 2838 2480 2844 2481
rect 2786 2463 2792 2464
rect 2786 2459 2787 2463
rect 2791 2459 2792 2463
rect 2786 2458 2792 2459
rect 2794 2463 2800 2464
rect 2794 2459 2795 2463
rect 2799 2459 2800 2463
rect 2794 2458 2800 2459
rect 2840 2447 2842 2480
rect 2916 2464 2918 2490
rect 2966 2485 2972 2486
rect 2966 2481 2967 2485
rect 2971 2481 2972 2485
rect 2966 2480 2972 2481
rect 2914 2463 2920 2464
rect 2914 2459 2915 2463
rect 2919 2459 2920 2463
rect 2914 2458 2920 2459
rect 2968 2447 2970 2480
rect 3044 2464 3046 2490
rect 3094 2485 3100 2486
rect 3094 2481 3095 2485
rect 3099 2481 3100 2485
rect 3094 2480 3100 2481
rect 3042 2463 3048 2464
rect 3042 2459 3043 2463
rect 3047 2459 3048 2463
rect 3042 2458 3048 2459
rect 3096 2447 3098 2480
rect 3172 2464 3174 2490
rect 3170 2463 3176 2464
rect 3170 2459 3171 2463
rect 3175 2459 3176 2463
rect 3170 2458 3176 2459
rect 2679 2446 2683 2447
rect 2679 2441 2683 2442
rect 2719 2446 2723 2447
rect 2719 2441 2723 2442
rect 2791 2446 2795 2447
rect 2791 2441 2795 2442
rect 2839 2446 2843 2447
rect 2839 2441 2843 2442
rect 2911 2446 2915 2447
rect 2911 2441 2915 2442
rect 2967 2446 2971 2447
rect 2967 2441 2971 2442
rect 3031 2446 3035 2447
rect 3031 2441 3035 2442
rect 3095 2446 3099 2447
rect 3095 2441 3099 2442
rect 3151 2446 3155 2447
rect 3151 2441 3155 2442
rect 2666 2439 2672 2440
rect 2666 2435 2667 2439
rect 2671 2435 2672 2439
rect 2666 2434 2672 2435
rect 2680 2420 2682 2441
rect 2762 2439 2768 2440
rect 2762 2435 2763 2439
rect 2767 2435 2768 2439
rect 2762 2434 2768 2435
rect 2558 2419 2564 2420
rect 2558 2415 2559 2419
rect 2563 2415 2564 2419
rect 2558 2414 2564 2415
rect 2678 2419 2684 2420
rect 2678 2415 2679 2419
rect 2683 2415 2684 2419
rect 2678 2414 2684 2415
rect 2764 2412 2766 2434
rect 2792 2420 2794 2441
rect 2874 2439 2880 2440
rect 2874 2435 2875 2439
rect 2879 2435 2880 2439
rect 2874 2434 2880 2435
rect 2790 2419 2796 2420
rect 2790 2415 2791 2419
rect 2795 2415 2796 2419
rect 2790 2414 2796 2415
rect 2876 2412 2878 2434
rect 2912 2420 2914 2441
rect 2994 2439 3000 2440
rect 2994 2435 2995 2439
rect 2999 2435 3000 2439
rect 2994 2434 3000 2435
rect 2910 2419 2916 2420
rect 2910 2415 2911 2419
rect 2915 2415 2916 2419
rect 2910 2414 2916 2415
rect 2996 2412 2998 2434
rect 3032 2420 3034 2441
rect 3114 2439 3120 2440
rect 3114 2435 3115 2439
rect 3119 2435 3120 2439
rect 3114 2434 3120 2435
rect 3030 2419 3036 2420
rect 3030 2415 3031 2419
rect 3035 2415 3036 2419
rect 3030 2414 3036 2415
rect 3116 2412 3118 2434
rect 3152 2420 3154 2441
rect 3216 2440 3218 2490
rect 3222 2485 3228 2486
rect 3222 2481 3223 2485
rect 3227 2481 3228 2485
rect 3222 2480 3228 2481
rect 3942 2484 3948 2485
rect 3942 2480 3943 2484
rect 3947 2480 3948 2484
rect 3224 2447 3226 2480
rect 3942 2479 3948 2480
rect 3944 2447 3946 2479
rect 3223 2446 3227 2447
rect 3223 2441 3227 2442
rect 3943 2446 3947 2447
rect 3943 2441 3947 2442
rect 3214 2439 3220 2440
rect 3214 2435 3215 2439
rect 3219 2435 3220 2439
rect 3214 2434 3220 2435
rect 3944 2421 3946 2441
rect 3942 2420 3948 2421
rect 3150 2419 3156 2420
rect 3150 2415 3151 2419
rect 3155 2415 3156 2419
rect 3942 2416 3943 2420
rect 3947 2416 3948 2420
rect 3942 2415 3948 2416
rect 3150 2414 3156 2415
rect 2266 2411 2272 2412
rect 2266 2407 2267 2411
rect 2271 2407 2272 2411
rect 2266 2406 2272 2407
rect 2274 2411 2280 2412
rect 2274 2407 2275 2411
rect 2279 2407 2280 2411
rect 2274 2406 2280 2407
rect 2422 2411 2428 2412
rect 2422 2407 2423 2411
rect 2427 2407 2428 2411
rect 2422 2406 2428 2407
rect 2522 2411 2528 2412
rect 2522 2407 2523 2411
rect 2527 2407 2528 2411
rect 2522 2406 2528 2407
rect 2642 2411 2648 2412
rect 2642 2407 2643 2411
rect 2647 2407 2648 2411
rect 2642 2406 2648 2407
rect 2762 2411 2768 2412
rect 2762 2407 2763 2411
rect 2767 2407 2768 2411
rect 2762 2406 2768 2407
rect 2874 2411 2880 2412
rect 2874 2407 2875 2411
rect 2879 2407 2880 2411
rect 2874 2406 2880 2407
rect 2994 2411 3000 2412
rect 2994 2407 2995 2411
rect 2999 2407 3000 2411
rect 2994 2406 3000 2407
rect 3114 2411 3120 2412
rect 3114 2407 3115 2411
rect 3119 2407 3120 2411
rect 3114 2406 3120 2407
rect 2318 2400 2324 2401
rect 2318 2396 2319 2400
rect 2323 2396 2324 2400
rect 2318 2395 2324 2396
rect 2320 2367 2322 2395
rect 2319 2366 2323 2367
rect 2319 2361 2323 2362
rect 2359 2366 2363 2367
rect 2359 2361 2363 2362
rect 2360 2337 2362 2361
rect 2358 2336 2364 2337
rect 2358 2332 2359 2336
rect 2363 2332 2364 2336
rect 2358 2331 2364 2332
rect 2242 2327 2248 2328
rect 2242 2323 2243 2327
rect 2247 2323 2248 2327
rect 2242 2322 2248 2323
rect 2350 2327 2356 2328
rect 2350 2323 2351 2327
rect 2355 2323 2356 2327
rect 2350 2322 2356 2323
rect 2166 2317 2172 2318
rect 2046 2316 2052 2317
rect 2046 2312 2047 2316
rect 2051 2312 2052 2316
rect 2166 2313 2167 2317
rect 2171 2313 2172 2317
rect 2166 2312 2172 2313
rect 2046 2311 2052 2312
rect 1902 2299 1908 2300
rect 2006 2301 2012 2302
rect 2006 2297 2007 2301
rect 2011 2297 2012 2301
rect 2006 2296 2012 2297
rect 1874 2295 1880 2296
rect 1874 2291 1875 2295
rect 1879 2291 1880 2295
rect 2048 2291 2050 2311
rect 2168 2291 2170 2312
rect 2234 2295 2240 2296
rect 2234 2291 2235 2295
rect 2239 2291 2240 2295
rect 1874 2290 1880 2291
rect 2047 2290 2051 2291
rect 1876 2264 1878 2290
rect 1902 2285 1908 2286
rect 2047 2285 2051 2286
rect 2071 2290 2075 2291
rect 2071 2285 2075 2286
rect 2167 2290 2171 2291
rect 2234 2290 2240 2291
rect 2287 2290 2291 2291
rect 2167 2285 2171 2286
rect 1902 2281 1903 2285
rect 1907 2281 1908 2285
rect 1902 2280 1908 2281
rect 2006 2284 2012 2285
rect 2006 2280 2007 2284
rect 2011 2280 2012 2284
rect 1866 2263 1872 2264
rect 1866 2259 1867 2263
rect 1871 2259 1872 2263
rect 1866 2258 1872 2259
rect 1874 2263 1880 2264
rect 1874 2259 1875 2263
rect 1879 2259 1880 2263
rect 1874 2258 1880 2259
rect 1904 2255 1906 2280
rect 2006 2279 2012 2280
rect 2008 2255 2010 2279
rect 2048 2265 2050 2285
rect 2046 2264 2052 2265
rect 2072 2264 2074 2285
rect 2146 2283 2152 2284
rect 2146 2279 2147 2283
rect 2151 2279 2152 2283
rect 2146 2278 2152 2279
rect 2046 2260 2047 2264
rect 2051 2260 2052 2264
rect 2046 2259 2052 2260
rect 2070 2263 2076 2264
rect 2070 2259 2071 2263
rect 2075 2259 2076 2263
rect 2070 2258 2076 2259
rect 2148 2256 2150 2278
rect 2168 2264 2170 2285
rect 2236 2272 2238 2290
rect 2287 2285 2291 2286
rect 2234 2271 2240 2272
rect 2234 2267 2235 2271
rect 2239 2267 2240 2271
rect 2234 2266 2240 2267
rect 2288 2264 2290 2285
rect 2352 2284 2354 2322
rect 2358 2317 2364 2318
rect 2358 2313 2359 2317
rect 2363 2313 2364 2317
rect 2358 2312 2364 2313
rect 2360 2291 2362 2312
rect 2424 2300 2426 2406
rect 2438 2400 2444 2401
rect 2438 2396 2439 2400
rect 2443 2396 2444 2400
rect 2438 2395 2444 2396
rect 2558 2400 2564 2401
rect 2558 2396 2559 2400
rect 2563 2396 2564 2400
rect 2558 2395 2564 2396
rect 2440 2367 2442 2395
rect 2560 2367 2562 2395
rect 2439 2366 2443 2367
rect 2439 2361 2443 2362
rect 2535 2366 2539 2367
rect 2535 2361 2539 2362
rect 2559 2366 2563 2367
rect 2559 2361 2563 2362
rect 2536 2337 2538 2361
rect 2534 2336 2540 2337
rect 2534 2332 2535 2336
rect 2539 2332 2540 2336
rect 2534 2331 2540 2332
rect 2534 2317 2540 2318
rect 2534 2313 2535 2317
rect 2539 2313 2540 2317
rect 2534 2312 2540 2313
rect 2422 2299 2428 2300
rect 2422 2295 2423 2299
rect 2427 2295 2428 2299
rect 2422 2294 2428 2295
rect 2536 2291 2538 2312
rect 2644 2296 2646 2406
rect 3942 2403 3948 2404
rect 2678 2400 2684 2401
rect 2678 2396 2679 2400
rect 2683 2396 2684 2400
rect 2678 2395 2684 2396
rect 2790 2400 2796 2401
rect 2790 2396 2791 2400
rect 2795 2396 2796 2400
rect 2790 2395 2796 2396
rect 2910 2400 2916 2401
rect 2910 2396 2911 2400
rect 2915 2396 2916 2400
rect 2910 2395 2916 2396
rect 3030 2400 3036 2401
rect 3030 2396 3031 2400
rect 3035 2396 3036 2400
rect 3030 2395 3036 2396
rect 3150 2400 3156 2401
rect 3150 2396 3151 2400
rect 3155 2396 3156 2400
rect 3942 2399 3943 2403
rect 3947 2399 3948 2403
rect 3942 2398 3948 2399
rect 3150 2395 3156 2396
rect 2680 2367 2682 2395
rect 2792 2367 2794 2395
rect 2912 2367 2914 2395
rect 3032 2367 3034 2395
rect 3152 2367 3154 2395
rect 3944 2367 3946 2398
rect 2679 2366 2683 2367
rect 2679 2361 2683 2362
rect 2703 2366 2707 2367
rect 2703 2361 2707 2362
rect 2791 2366 2795 2367
rect 2791 2361 2795 2362
rect 2871 2366 2875 2367
rect 2871 2361 2875 2362
rect 2911 2366 2915 2367
rect 2911 2361 2915 2362
rect 3031 2366 3035 2367
rect 3031 2361 3035 2362
rect 3151 2366 3155 2367
rect 3151 2361 3155 2362
rect 3199 2366 3203 2367
rect 3199 2361 3203 2362
rect 3943 2366 3947 2367
rect 3943 2361 3947 2362
rect 2704 2337 2706 2361
rect 2872 2337 2874 2361
rect 3032 2337 3034 2361
rect 3200 2337 3202 2361
rect 2702 2336 2708 2337
rect 2702 2332 2703 2336
rect 2707 2332 2708 2336
rect 2702 2331 2708 2332
rect 2870 2336 2876 2337
rect 2870 2332 2871 2336
rect 2875 2332 2876 2336
rect 2870 2331 2876 2332
rect 3030 2336 3036 2337
rect 3030 2332 3031 2336
rect 3035 2332 3036 2336
rect 3030 2331 3036 2332
rect 3198 2336 3204 2337
rect 3198 2332 3199 2336
rect 3203 2332 3204 2336
rect 3944 2334 3946 2361
rect 3198 2331 3204 2332
rect 3942 2333 3948 2334
rect 3942 2329 3943 2333
rect 3947 2329 3948 2333
rect 3942 2328 3948 2329
rect 2670 2327 2676 2328
rect 2670 2323 2671 2327
rect 2675 2323 2676 2327
rect 2670 2322 2676 2323
rect 2778 2327 2784 2328
rect 2778 2323 2779 2327
rect 2783 2323 2784 2327
rect 2778 2322 2784 2323
rect 2946 2327 2952 2328
rect 2946 2323 2947 2327
rect 2951 2323 2952 2327
rect 2946 2322 2952 2323
rect 3106 2327 3112 2328
rect 3106 2323 3107 2327
rect 3111 2323 3112 2327
rect 3106 2322 3112 2323
rect 3114 2327 3120 2328
rect 3114 2323 3115 2327
rect 3119 2323 3120 2327
rect 3114 2322 3120 2323
rect 2672 2296 2674 2322
rect 2702 2317 2708 2318
rect 2702 2313 2703 2317
rect 2707 2313 2708 2317
rect 2702 2312 2708 2313
rect 2642 2295 2648 2296
rect 2642 2291 2643 2295
rect 2647 2291 2648 2295
rect 2359 2290 2363 2291
rect 2359 2285 2363 2286
rect 2423 2290 2427 2291
rect 2423 2285 2427 2286
rect 2535 2290 2539 2291
rect 2535 2285 2539 2286
rect 2559 2290 2563 2291
rect 2642 2290 2648 2291
rect 2670 2295 2676 2296
rect 2670 2291 2671 2295
rect 2675 2291 2676 2295
rect 2704 2291 2706 2312
rect 2780 2296 2782 2322
rect 2870 2317 2876 2318
rect 2870 2313 2871 2317
rect 2875 2313 2876 2317
rect 2870 2312 2876 2313
rect 2778 2295 2784 2296
rect 2778 2291 2779 2295
rect 2783 2291 2784 2295
rect 2872 2291 2874 2312
rect 2948 2296 2950 2322
rect 3030 2317 3036 2318
rect 3030 2313 3031 2317
rect 3035 2313 3036 2317
rect 3030 2312 3036 2313
rect 2946 2295 2952 2296
rect 2946 2291 2947 2295
rect 2951 2291 2952 2295
rect 3032 2291 3034 2312
rect 3108 2296 3110 2322
rect 3106 2295 3112 2296
rect 3106 2291 3107 2295
rect 3111 2291 3112 2295
rect 2670 2290 2676 2291
rect 2703 2290 2707 2291
rect 2778 2290 2784 2291
rect 2839 2290 2843 2291
rect 2559 2285 2563 2286
rect 2703 2285 2707 2286
rect 2839 2285 2843 2286
rect 2871 2290 2875 2291
rect 2946 2290 2952 2291
rect 2983 2290 2987 2291
rect 2871 2285 2875 2286
rect 2983 2285 2987 2286
rect 3031 2290 3035 2291
rect 3106 2290 3112 2291
rect 3031 2285 3035 2286
rect 2350 2283 2356 2284
rect 2350 2279 2351 2283
rect 2355 2279 2356 2283
rect 2350 2278 2356 2279
rect 2370 2283 2376 2284
rect 2370 2279 2371 2283
rect 2375 2279 2376 2283
rect 2370 2278 2376 2279
rect 2166 2263 2172 2264
rect 2166 2259 2167 2263
rect 2171 2259 2172 2263
rect 2166 2258 2172 2259
rect 2286 2263 2292 2264
rect 2286 2259 2287 2263
rect 2291 2259 2292 2263
rect 2286 2258 2292 2259
rect 2146 2255 2152 2256
rect 1671 2254 1675 2255
rect 1671 2249 1675 2250
rect 1767 2254 1771 2255
rect 1767 2249 1771 2250
rect 1799 2254 1803 2255
rect 1799 2249 1803 2250
rect 1903 2254 1907 2255
rect 1903 2249 1907 2250
rect 2007 2254 2011 2255
rect 2146 2251 2147 2255
rect 2151 2251 2152 2255
rect 2146 2250 2152 2251
rect 2154 2255 2160 2256
rect 2154 2251 2155 2255
rect 2159 2251 2160 2255
rect 2154 2250 2160 2251
rect 2362 2251 2368 2252
rect 2007 2249 2011 2250
rect 1650 2247 1656 2248
rect 1650 2243 1651 2247
rect 1655 2243 1656 2247
rect 1650 2242 1656 2243
rect 1754 2247 1760 2248
rect 1754 2243 1755 2247
rect 1759 2243 1760 2247
rect 1754 2242 1760 2243
rect 1652 2220 1654 2242
rect 1066 2219 1072 2220
rect 1066 2215 1067 2219
rect 1071 2215 1072 2219
rect 1066 2214 1072 2215
rect 1250 2219 1256 2220
rect 1250 2215 1251 2219
rect 1255 2215 1256 2219
rect 1250 2214 1256 2215
rect 1258 2219 1264 2220
rect 1258 2215 1259 2219
rect 1263 2215 1264 2219
rect 1258 2214 1264 2215
rect 1642 2219 1648 2220
rect 1642 2215 1643 2219
rect 1647 2215 1648 2219
rect 1642 2214 1648 2215
rect 1650 2219 1656 2220
rect 1650 2215 1651 2219
rect 1655 2215 1656 2219
rect 1650 2214 1656 2215
rect 822 2208 828 2209
rect 822 2204 823 2208
rect 827 2204 828 2208
rect 822 2203 828 2204
rect 990 2208 996 2209
rect 990 2204 991 2208
rect 995 2204 996 2208
rect 990 2203 996 2204
rect 1174 2208 1180 2209
rect 1174 2204 1175 2208
rect 1179 2204 1180 2208
rect 1174 2203 1180 2204
rect 824 2171 826 2203
rect 992 2171 994 2203
rect 1176 2171 1178 2203
rect 823 2170 827 2171
rect 823 2165 827 2166
rect 871 2170 875 2171
rect 871 2165 875 2166
rect 991 2170 995 2171
rect 991 2165 995 2166
rect 1031 2170 1035 2171
rect 1031 2165 1035 2166
rect 1175 2170 1179 2171
rect 1175 2165 1179 2166
rect 1191 2170 1195 2171
rect 1191 2165 1195 2166
rect 872 2141 874 2165
rect 1032 2141 1034 2165
rect 1192 2141 1194 2165
rect 870 2140 876 2141
rect 870 2136 871 2140
rect 875 2136 876 2140
rect 870 2135 876 2136
rect 1030 2140 1036 2141
rect 1030 2136 1031 2140
rect 1035 2136 1036 2140
rect 1030 2135 1036 2136
rect 1190 2140 1196 2141
rect 1190 2136 1191 2140
rect 1195 2136 1196 2140
rect 1190 2135 1196 2136
rect 322 2131 328 2132
rect 322 2127 323 2131
rect 327 2127 328 2131
rect 322 2126 328 2127
rect 466 2131 472 2132
rect 466 2127 467 2131
rect 471 2127 472 2131
rect 466 2126 472 2127
rect 626 2131 632 2132
rect 626 2127 627 2131
rect 631 2127 632 2131
rect 626 2126 632 2127
rect 778 2131 784 2132
rect 778 2127 779 2131
rect 783 2127 784 2131
rect 778 2126 784 2127
rect 938 2131 944 2132
rect 938 2127 939 2131
rect 943 2127 944 2131
rect 938 2126 944 2127
rect 954 2131 960 2132
rect 954 2127 955 2131
rect 959 2127 960 2131
rect 954 2126 960 2127
rect 134 2121 140 2122
rect 110 2120 116 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 134 2117 135 2121
rect 139 2117 140 2121
rect 134 2116 140 2117
rect 246 2121 252 2122
rect 246 2117 247 2121
rect 251 2117 252 2121
rect 246 2116 252 2117
rect 110 2115 116 2116
rect 112 2087 114 2115
rect 136 2087 138 2116
rect 210 2099 216 2100
rect 210 2095 211 2099
rect 215 2095 216 2099
rect 210 2094 216 2095
rect 111 2086 115 2087
rect 111 2081 115 2082
rect 135 2086 139 2087
rect 135 2081 139 2082
rect 112 2061 114 2081
rect 110 2060 116 2061
rect 136 2060 138 2081
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 134 2059 140 2060
rect 134 2055 135 2059
rect 139 2055 140 2059
rect 134 2054 140 2055
rect 212 2052 214 2094
rect 248 2087 250 2116
rect 324 2100 326 2126
rect 390 2121 396 2122
rect 390 2117 391 2121
rect 395 2117 396 2121
rect 390 2116 396 2117
rect 322 2099 328 2100
rect 322 2095 323 2099
rect 327 2095 328 2099
rect 322 2094 328 2095
rect 392 2087 394 2116
rect 468 2100 470 2126
rect 550 2121 556 2122
rect 550 2117 551 2121
rect 555 2117 556 2121
rect 550 2116 556 2117
rect 466 2099 472 2100
rect 466 2095 467 2099
rect 471 2095 472 2099
rect 466 2094 472 2095
rect 552 2087 554 2116
rect 628 2100 630 2126
rect 710 2121 716 2122
rect 710 2117 711 2121
rect 715 2117 716 2121
rect 710 2116 716 2117
rect 870 2121 876 2122
rect 870 2117 871 2121
rect 875 2117 876 2121
rect 870 2116 876 2117
rect 626 2099 632 2100
rect 626 2095 627 2099
rect 631 2095 632 2099
rect 626 2094 632 2095
rect 712 2087 714 2116
rect 872 2087 874 2116
rect 247 2086 251 2087
rect 247 2081 251 2082
rect 391 2086 395 2087
rect 391 2081 395 2082
rect 399 2086 403 2087
rect 399 2081 403 2082
rect 551 2086 555 2087
rect 551 2081 555 2082
rect 703 2086 707 2087
rect 703 2081 707 2082
rect 711 2086 715 2087
rect 711 2081 715 2082
rect 847 2086 851 2087
rect 847 2081 851 2082
rect 871 2086 875 2087
rect 871 2081 875 2082
rect 218 2079 224 2080
rect 218 2075 219 2079
rect 223 2075 224 2079
rect 218 2074 224 2075
rect 220 2052 222 2074
rect 248 2060 250 2081
rect 378 2079 384 2080
rect 378 2075 379 2079
rect 383 2075 384 2079
rect 378 2074 384 2075
rect 246 2059 252 2060
rect 246 2055 247 2059
rect 251 2055 252 2059
rect 246 2054 252 2055
rect 380 2052 382 2074
rect 400 2060 402 2081
rect 482 2079 488 2080
rect 482 2075 483 2079
rect 487 2075 488 2079
rect 482 2074 488 2075
rect 398 2059 404 2060
rect 398 2055 399 2059
rect 403 2055 404 2059
rect 398 2054 404 2055
rect 484 2052 486 2074
rect 552 2060 554 2081
rect 634 2079 640 2080
rect 634 2075 635 2079
rect 639 2075 640 2079
rect 634 2074 640 2075
rect 550 2059 556 2060
rect 550 2055 551 2059
rect 555 2055 556 2059
rect 550 2054 556 2055
rect 636 2052 638 2074
rect 704 2060 706 2081
rect 848 2060 850 2081
rect 940 2080 942 2126
rect 956 2100 958 2126
rect 1030 2121 1036 2122
rect 1030 2117 1031 2121
rect 1035 2117 1036 2121
rect 1030 2116 1036 2117
rect 1190 2121 1196 2122
rect 1190 2117 1191 2121
rect 1195 2117 1196 2121
rect 1190 2116 1196 2117
rect 954 2099 960 2100
rect 954 2095 955 2099
rect 959 2095 960 2099
rect 954 2094 960 2095
rect 1032 2087 1034 2116
rect 1192 2087 1194 2116
rect 1260 2100 1262 2214
rect 1366 2208 1372 2209
rect 1366 2204 1367 2208
rect 1371 2204 1372 2208
rect 1366 2203 1372 2204
rect 1566 2208 1572 2209
rect 1566 2204 1567 2208
rect 1571 2204 1572 2208
rect 1566 2203 1572 2204
rect 1368 2171 1370 2203
rect 1568 2171 1570 2203
rect 1351 2170 1355 2171
rect 1351 2165 1355 2166
rect 1367 2170 1371 2171
rect 1367 2165 1371 2166
rect 1511 2170 1515 2171
rect 1511 2165 1515 2166
rect 1567 2170 1571 2171
rect 1567 2165 1571 2166
rect 1679 2170 1683 2171
rect 1679 2165 1683 2166
rect 1352 2141 1354 2165
rect 1512 2141 1514 2165
rect 1680 2141 1682 2165
rect 1350 2140 1356 2141
rect 1350 2136 1351 2140
rect 1355 2136 1356 2140
rect 1350 2135 1356 2136
rect 1510 2140 1516 2141
rect 1510 2136 1511 2140
rect 1515 2136 1516 2140
rect 1510 2135 1516 2136
rect 1678 2140 1684 2141
rect 1678 2136 1679 2140
rect 1683 2136 1684 2140
rect 1678 2135 1684 2136
rect 1756 2132 1758 2242
rect 1768 2228 1770 2249
rect 2008 2229 2010 2249
rect 2046 2247 2052 2248
rect 2046 2243 2047 2247
rect 2051 2243 2052 2247
rect 2046 2242 2052 2243
rect 2070 2244 2076 2245
rect 2006 2228 2012 2229
rect 1766 2227 1772 2228
rect 1766 2223 1767 2227
rect 1771 2223 1772 2227
rect 2006 2224 2007 2228
rect 2011 2224 2012 2228
rect 2006 2223 2012 2224
rect 1766 2222 1772 2223
rect 2048 2215 2050 2242
rect 2070 2240 2071 2244
rect 2075 2240 2076 2244
rect 2070 2239 2076 2240
rect 2072 2215 2074 2239
rect 2047 2214 2051 2215
rect 2006 2211 2012 2212
rect 1766 2208 1772 2209
rect 1766 2204 1767 2208
rect 1771 2204 1772 2208
rect 2006 2207 2007 2211
rect 2011 2207 2012 2211
rect 2047 2209 2051 2210
rect 2071 2214 2075 2215
rect 2071 2209 2075 2210
rect 2006 2206 2012 2207
rect 1766 2203 1772 2204
rect 1768 2171 1770 2203
rect 2008 2171 2010 2206
rect 2048 2182 2050 2209
rect 2072 2185 2074 2209
rect 2070 2184 2076 2185
rect 2046 2181 2052 2182
rect 2046 2177 2047 2181
rect 2051 2177 2052 2181
rect 2070 2180 2071 2184
rect 2075 2180 2076 2184
rect 2070 2179 2076 2180
rect 2046 2176 2052 2177
rect 1767 2170 1771 2171
rect 1767 2165 1771 2166
rect 2007 2170 2011 2171
rect 2007 2165 2011 2166
rect 2070 2165 2076 2166
rect 2008 2138 2010 2165
rect 2046 2164 2052 2165
rect 2046 2160 2047 2164
rect 2051 2160 2052 2164
rect 2070 2161 2071 2165
rect 2075 2161 2076 2165
rect 2070 2160 2076 2161
rect 2046 2159 2052 2160
rect 2006 2137 2012 2138
rect 2006 2133 2007 2137
rect 2011 2133 2012 2137
rect 2006 2132 2012 2133
rect 1426 2131 1432 2132
rect 1426 2127 1427 2131
rect 1431 2127 1432 2131
rect 1426 2126 1432 2127
rect 1586 2131 1592 2132
rect 1586 2127 1587 2131
rect 1591 2127 1592 2131
rect 1586 2126 1592 2127
rect 1754 2131 1760 2132
rect 1754 2127 1755 2131
rect 1759 2127 1760 2131
rect 1754 2126 1760 2127
rect 1350 2121 1356 2122
rect 1350 2117 1351 2121
rect 1355 2117 1356 2121
rect 1350 2116 1356 2117
rect 1258 2099 1264 2100
rect 1258 2095 1259 2099
rect 1263 2095 1264 2099
rect 1258 2094 1264 2095
rect 1352 2087 1354 2116
rect 1428 2100 1430 2126
rect 1510 2121 1516 2122
rect 1510 2117 1511 2121
rect 1515 2117 1516 2121
rect 1510 2116 1516 2117
rect 1426 2099 1432 2100
rect 1426 2095 1427 2099
rect 1431 2095 1432 2099
rect 1426 2094 1432 2095
rect 1512 2087 1514 2116
rect 1588 2100 1590 2126
rect 1678 2121 1684 2122
rect 1678 2117 1679 2121
rect 1683 2117 1684 2121
rect 1678 2116 1684 2117
rect 2006 2120 2012 2121
rect 2006 2116 2007 2120
rect 2011 2116 2012 2120
rect 1586 2099 1592 2100
rect 1586 2095 1587 2099
rect 1591 2095 1592 2099
rect 1586 2094 1592 2095
rect 1680 2087 1682 2116
rect 2006 2115 2012 2116
rect 2048 2115 2050 2159
rect 2072 2115 2074 2160
rect 2156 2144 2158 2250
rect 2362 2247 2363 2251
rect 2367 2247 2368 2251
rect 2362 2246 2368 2247
rect 2166 2244 2172 2245
rect 2166 2240 2167 2244
rect 2171 2240 2172 2244
rect 2166 2239 2172 2240
rect 2286 2244 2292 2245
rect 2286 2240 2287 2244
rect 2291 2240 2292 2244
rect 2286 2239 2292 2240
rect 2168 2215 2170 2239
rect 2288 2215 2290 2239
rect 2167 2214 2171 2215
rect 2167 2209 2171 2210
rect 2287 2214 2291 2215
rect 2287 2209 2291 2210
rect 2295 2214 2299 2215
rect 2295 2209 2299 2210
rect 2296 2185 2298 2209
rect 2294 2184 2300 2185
rect 2294 2180 2295 2184
rect 2299 2180 2300 2184
rect 2294 2179 2300 2180
rect 2294 2165 2300 2166
rect 2294 2161 2295 2165
rect 2299 2161 2300 2165
rect 2294 2160 2300 2161
rect 2154 2143 2160 2144
rect 2154 2139 2155 2143
rect 2159 2139 2160 2143
rect 2154 2138 2160 2139
rect 2296 2115 2298 2160
rect 2364 2144 2366 2246
rect 2372 2192 2374 2278
rect 2424 2264 2426 2285
rect 2498 2283 2504 2284
rect 2498 2279 2499 2283
rect 2503 2279 2504 2283
rect 2498 2278 2504 2279
rect 2422 2263 2428 2264
rect 2422 2259 2423 2263
rect 2427 2259 2428 2263
rect 2422 2258 2428 2259
rect 2500 2256 2502 2278
rect 2560 2264 2562 2285
rect 2634 2283 2640 2284
rect 2634 2279 2635 2283
rect 2639 2279 2640 2283
rect 2634 2278 2640 2279
rect 2558 2263 2564 2264
rect 2558 2259 2559 2263
rect 2563 2259 2564 2263
rect 2558 2258 2564 2259
rect 2636 2256 2638 2278
rect 2704 2264 2706 2285
rect 2840 2264 2842 2285
rect 2914 2283 2920 2284
rect 2914 2279 2915 2283
rect 2919 2279 2920 2283
rect 2914 2278 2920 2279
rect 2702 2263 2708 2264
rect 2702 2259 2703 2263
rect 2707 2259 2708 2263
rect 2702 2258 2708 2259
rect 2838 2263 2844 2264
rect 2838 2259 2839 2263
rect 2843 2259 2844 2263
rect 2838 2258 2844 2259
rect 2916 2256 2918 2278
rect 2984 2264 2986 2285
rect 3058 2283 3064 2284
rect 3058 2279 3059 2283
rect 3063 2279 3064 2283
rect 3058 2278 3064 2279
rect 2982 2263 2988 2264
rect 2982 2259 2983 2263
rect 2987 2259 2988 2263
rect 2982 2258 2988 2259
rect 3060 2256 3062 2278
rect 3116 2276 3118 2322
rect 3198 2317 3204 2318
rect 3198 2313 3199 2317
rect 3203 2313 3204 2317
rect 3198 2312 3204 2313
rect 3942 2316 3948 2317
rect 3942 2312 3943 2316
rect 3947 2312 3948 2316
rect 3200 2291 3202 2312
rect 3942 2311 3948 2312
rect 3944 2291 3946 2311
rect 3127 2290 3131 2291
rect 3127 2285 3131 2286
rect 3199 2290 3203 2291
rect 3199 2285 3203 2286
rect 3271 2290 3275 2291
rect 3271 2285 3275 2286
rect 3943 2290 3947 2291
rect 3943 2285 3947 2286
rect 3114 2275 3120 2276
rect 3114 2271 3115 2275
rect 3119 2271 3120 2275
rect 3114 2270 3120 2271
rect 3128 2264 3130 2285
rect 3250 2283 3256 2284
rect 3250 2279 3251 2283
rect 3255 2279 3256 2283
rect 3250 2278 3256 2279
rect 3126 2263 3132 2264
rect 3126 2259 3127 2263
rect 3131 2259 3132 2263
rect 3126 2258 3132 2259
rect 3252 2256 3254 2278
rect 3272 2264 3274 2285
rect 3944 2265 3946 2285
rect 3942 2264 3948 2265
rect 3270 2263 3276 2264
rect 3270 2259 3271 2263
rect 3275 2259 3276 2263
rect 3942 2260 3943 2264
rect 3947 2260 3948 2264
rect 3942 2259 3948 2260
rect 3270 2258 3276 2259
rect 2498 2255 2504 2256
rect 2498 2251 2499 2255
rect 2503 2251 2504 2255
rect 2498 2250 2504 2251
rect 2634 2255 2640 2256
rect 2634 2251 2635 2255
rect 2639 2251 2640 2255
rect 2634 2250 2640 2251
rect 2914 2255 2920 2256
rect 2914 2251 2915 2255
rect 2919 2251 2920 2255
rect 2914 2250 2920 2251
rect 3058 2255 3064 2256
rect 3058 2251 3059 2255
rect 3063 2251 3064 2255
rect 3058 2250 3064 2251
rect 3250 2255 3256 2256
rect 3250 2251 3251 2255
rect 3255 2251 3256 2255
rect 3250 2250 3256 2251
rect 3258 2255 3264 2256
rect 3258 2251 3259 2255
rect 3263 2251 3264 2255
rect 3258 2250 3264 2251
rect 2422 2244 2428 2245
rect 2422 2240 2423 2244
rect 2427 2240 2428 2244
rect 2422 2239 2428 2240
rect 2558 2244 2564 2245
rect 2558 2240 2559 2244
rect 2563 2240 2564 2244
rect 2558 2239 2564 2240
rect 2702 2244 2708 2245
rect 2702 2240 2703 2244
rect 2707 2240 2708 2244
rect 2702 2239 2708 2240
rect 2838 2244 2844 2245
rect 2838 2240 2839 2244
rect 2843 2240 2844 2244
rect 2838 2239 2844 2240
rect 2982 2244 2988 2245
rect 2982 2240 2983 2244
rect 2987 2240 2988 2244
rect 2982 2239 2988 2240
rect 3126 2244 3132 2245
rect 3126 2240 3127 2244
rect 3131 2240 3132 2244
rect 3126 2239 3132 2240
rect 2424 2215 2426 2239
rect 2560 2215 2562 2239
rect 2704 2215 2706 2239
rect 2840 2215 2842 2239
rect 2984 2215 2986 2239
rect 3128 2215 3130 2239
rect 2423 2214 2427 2215
rect 2423 2209 2427 2210
rect 2503 2214 2507 2215
rect 2503 2209 2507 2210
rect 2559 2214 2563 2215
rect 2559 2209 2563 2210
rect 2687 2214 2691 2215
rect 2687 2209 2691 2210
rect 2703 2214 2707 2215
rect 2703 2209 2707 2210
rect 2839 2214 2843 2215
rect 2839 2209 2843 2210
rect 2863 2214 2867 2215
rect 2863 2209 2867 2210
rect 2983 2214 2987 2215
rect 2983 2209 2987 2210
rect 3023 2214 3027 2215
rect 3023 2209 3027 2210
rect 3127 2214 3131 2215
rect 3127 2209 3131 2210
rect 3175 2214 3179 2215
rect 3175 2209 3179 2210
rect 2370 2191 2376 2192
rect 2370 2187 2371 2191
rect 2375 2187 2376 2191
rect 2370 2186 2376 2187
rect 2504 2185 2506 2209
rect 2688 2185 2690 2209
rect 2864 2185 2866 2209
rect 3024 2185 3026 2209
rect 3176 2185 3178 2209
rect 2502 2184 2508 2185
rect 2502 2180 2503 2184
rect 2507 2180 2508 2184
rect 2502 2179 2508 2180
rect 2686 2184 2692 2185
rect 2686 2180 2687 2184
rect 2691 2180 2692 2184
rect 2686 2179 2692 2180
rect 2862 2184 2868 2185
rect 2862 2180 2863 2184
rect 2867 2180 2868 2184
rect 2862 2179 2868 2180
rect 3022 2184 3028 2185
rect 3022 2180 3023 2184
rect 3027 2180 3028 2184
rect 3022 2179 3028 2180
rect 3174 2184 3180 2185
rect 3174 2180 3175 2184
rect 3179 2180 3180 2184
rect 3174 2179 3180 2180
rect 2370 2175 2376 2176
rect 2370 2171 2371 2175
rect 2375 2171 2376 2175
rect 2370 2170 2376 2171
rect 2578 2175 2584 2176
rect 2578 2171 2579 2175
rect 2583 2171 2584 2175
rect 2578 2170 2584 2171
rect 2754 2175 2760 2176
rect 2754 2171 2755 2175
rect 2759 2171 2760 2175
rect 2754 2170 2760 2171
rect 2938 2175 2944 2176
rect 2938 2171 2939 2175
rect 2943 2171 2944 2175
rect 2938 2170 2944 2171
rect 3098 2175 3104 2176
rect 3098 2171 3099 2175
rect 3103 2171 3104 2175
rect 3098 2170 3104 2171
rect 3250 2175 3256 2176
rect 3250 2171 3251 2175
rect 3255 2171 3256 2175
rect 3250 2170 3256 2171
rect 2372 2144 2374 2170
rect 2502 2165 2508 2166
rect 2502 2161 2503 2165
rect 2507 2161 2508 2165
rect 2502 2160 2508 2161
rect 2362 2143 2368 2144
rect 2362 2139 2363 2143
rect 2367 2139 2368 2143
rect 2362 2138 2368 2139
rect 2370 2143 2376 2144
rect 2370 2139 2371 2143
rect 2375 2139 2376 2143
rect 2370 2138 2376 2139
rect 2504 2115 2506 2160
rect 2580 2144 2582 2170
rect 2686 2165 2692 2166
rect 2686 2161 2687 2165
rect 2691 2161 2692 2165
rect 2686 2160 2692 2161
rect 2578 2143 2584 2144
rect 2578 2139 2579 2143
rect 2583 2139 2584 2143
rect 2578 2138 2584 2139
rect 2688 2115 2690 2160
rect 2008 2087 2010 2115
rect 2047 2114 2051 2115
rect 2047 2109 2051 2110
rect 2071 2114 2075 2115
rect 2071 2109 2075 2110
rect 2295 2114 2299 2115
rect 2295 2109 2299 2110
rect 2399 2114 2403 2115
rect 2399 2109 2403 2110
rect 2495 2114 2499 2115
rect 2495 2109 2499 2110
rect 2503 2114 2507 2115
rect 2503 2109 2507 2110
rect 2591 2114 2595 2115
rect 2591 2109 2595 2110
rect 2687 2114 2691 2115
rect 2687 2109 2691 2110
rect 2048 2089 2050 2109
rect 2046 2088 2052 2089
rect 2400 2088 2402 2109
rect 2474 2107 2480 2108
rect 2474 2103 2475 2107
rect 2479 2103 2480 2107
rect 2474 2102 2480 2103
rect 991 2086 995 2087
rect 991 2081 995 2082
rect 1031 2086 1035 2087
rect 1031 2081 1035 2082
rect 1127 2086 1131 2087
rect 1127 2081 1131 2082
rect 1191 2086 1195 2087
rect 1191 2081 1195 2082
rect 1255 2086 1259 2087
rect 1255 2081 1259 2082
rect 1351 2086 1355 2087
rect 1351 2081 1355 2082
rect 1383 2086 1387 2087
rect 1383 2081 1387 2082
rect 1511 2086 1515 2087
rect 1511 2081 1515 2082
rect 1519 2086 1523 2087
rect 1519 2081 1523 2082
rect 1679 2086 1683 2087
rect 1679 2081 1683 2082
rect 2007 2086 2011 2087
rect 2046 2084 2047 2088
rect 2051 2084 2052 2088
rect 2046 2083 2052 2084
rect 2398 2087 2404 2088
rect 2398 2083 2399 2087
rect 2403 2083 2404 2087
rect 2398 2082 2404 2083
rect 2007 2081 2011 2082
rect 878 2079 884 2080
rect 878 2075 879 2079
rect 883 2075 884 2079
rect 878 2074 884 2075
rect 938 2079 944 2080
rect 938 2075 939 2079
rect 943 2075 944 2079
rect 938 2074 944 2075
rect 970 2079 976 2080
rect 970 2075 971 2079
rect 975 2075 976 2079
rect 970 2074 976 2075
rect 702 2059 708 2060
rect 702 2055 703 2059
rect 707 2055 708 2059
rect 702 2054 708 2055
rect 846 2059 852 2060
rect 846 2055 847 2059
rect 851 2055 852 2059
rect 846 2054 852 2055
rect 210 2051 216 2052
rect 210 2047 211 2051
rect 215 2047 216 2051
rect 210 2046 216 2047
rect 218 2051 224 2052
rect 218 2047 219 2051
rect 223 2047 224 2051
rect 218 2046 224 2047
rect 378 2051 384 2052
rect 378 2047 379 2051
rect 383 2047 384 2051
rect 378 2046 384 2047
rect 482 2051 488 2052
rect 482 2047 483 2051
rect 487 2047 488 2051
rect 482 2046 488 2047
rect 634 2051 640 2052
rect 634 2047 635 2051
rect 639 2047 640 2051
rect 634 2046 640 2047
rect 110 2043 116 2044
rect 110 2039 111 2043
rect 115 2039 116 2043
rect 110 2038 116 2039
rect 134 2040 140 2041
rect 112 1995 114 2038
rect 134 2036 135 2040
rect 139 2036 140 2040
rect 134 2035 140 2036
rect 246 2040 252 2041
rect 246 2036 247 2040
rect 251 2036 252 2040
rect 246 2035 252 2036
rect 398 2040 404 2041
rect 398 2036 399 2040
rect 403 2036 404 2040
rect 398 2035 404 2036
rect 550 2040 556 2041
rect 550 2036 551 2040
rect 555 2036 556 2040
rect 550 2035 556 2036
rect 702 2040 708 2041
rect 702 2036 703 2040
rect 707 2036 708 2040
rect 702 2035 708 2036
rect 846 2040 852 2041
rect 846 2036 847 2040
rect 851 2036 852 2040
rect 846 2035 852 2036
rect 136 1995 138 2035
rect 248 1995 250 2035
rect 400 1995 402 2035
rect 552 1995 554 2035
rect 704 1995 706 2035
rect 848 1995 850 2035
rect 111 1994 115 1995
rect 111 1989 115 1990
rect 135 1994 139 1995
rect 135 1989 139 1990
rect 231 1994 235 1995
rect 231 1989 235 1990
rect 247 1994 251 1995
rect 247 1989 251 1990
rect 391 1994 395 1995
rect 391 1989 395 1990
rect 399 1994 403 1995
rect 399 1989 403 1990
rect 551 1994 555 1995
rect 551 1989 555 1990
rect 567 1994 571 1995
rect 567 1989 571 1990
rect 703 1994 707 1995
rect 703 1989 707 1990
rect 751 1994 755 1995
rect 751 1989 755 1990
rect 847 1994 851 1995
rect 847 1989 851 1990
rect 112 1962 114 1989
rect 232 1965 234 1989
rect 392 1965 394 1989
rect 568 1965 570 1989
rect 752 1965 754 1989
rect 230 1964 236 1965
rect 110 1961 116 1962
rect 110 1957 111 1961
rect 115 1957 116 1961
rect 230 1960 231 1964
rect 235 1960 236 1964
rect 230 1959 236 1960
rect 390 1964 396 1965
rect 390 1960 391 1964
rect 395 1960 396 1964
rect 390 1959 396 1960
rect 566 1964 572 1965
rect 566 1960 567 1964
rect 571 1960 572 1964
rect 566 1959 572 1960
rect 750 1964 756 1965
rect 750 1960 751 1964
rect 755 1960 756 1964
rect 750 1959 756 1960
rect 110 1956 116 1957
rect 880 1956 882 2074
rect 972 2052 974 2074
rect 992 2060 994 2081
rect 1066 2079 1072 2080
rect 1066 2075 1067 2079
rect 1071 2075 1072 2079
rect 1066 2074 1072 2075
rect 990 2059 996 2060
rect 990 2055 991 2059
rect 995 2055 996 2059
rect 990 2054 996 2055
rect 1068 2052 1070 2074
rect 1128 2060 1130 2081
rect 1202 2079 1208 2080
rect 1202 2075 1203 2079
rect 1207 2075 1208 2079
rect 1202 2074 1208 2075
rect 1126 2059 1132 2060
rect 1126 2055 1127 2059
rect 1131 2055 1132 2059
rect 1126 2054 1132 2055
rect 1204 2052 1206 2074
rect 1256 2060 1258 2081
rect 1330 2079 1336 2080
rect 1330 2075 1331 2079
rect 1335 2075 1336 2079
rect 1330 2074 1336 2075
rect 1254 2059 1260 2060
rect 1254 2055 1255 2059
rect 1259 2055 1260 2059
rect 1254 2054 1260 2055
rect 1332 2052 1334 2074
rect 1384 2060 1386 2081
rect 1458 2079 1464 2080
rect 1458 2075 1459 2079
rect 1463 2075 1464 2079
rect 1458 2074 1464 2075
rect 1382 2059 1388 2060
rect 1382 2055 1383 2059
rect 1387 2055 1388 2059
rect 1382 2054 1388 2055
rect 1460 2052 1462 2074
rect 1520 2060 1522 2081
rect 2008 2061 2010 2081
rect 2476 2080 2478 2102
rect 2496 2088 2498 2109
rect 2570 2107 2576 2108
rect 2570 2103 2571 2107
rect 2575 2103 2576 2107
rect 2570 2102 2576 2103
rect 2494 2087 2500 2088
rect 2494 2083 2495 2087
rect 2499 2083 2500 2087
rect 2494 2082 2500 2083
rect 2572 2080 2574 2102
rect 2592 2088 2594 2109
rect 2666 2099 2672 2100
rect 2666 2095 2667 2099
rect 2671 2095 2672 2099
rect 2666 2094 2672 2095
rect 2590 2087 2596 2088
rect 2590 2083 2591 2087
rect 2595 2083 2596 2087
rect 2590 2082 2596 2083
rect 2668 2080 2670 2094
rect 2688 2088 2690 2109
rect 2756 2108 2758 2170
rect 2862 2165 2868 2166
rect 2862 2161 2863 2165
rect 2867 2161 2868 2165
rect 2862 2160 2868 2161
rect 2864 2115 2866 2160
rect 2940 2144 2942 2170
rect 3022 2165 3028 2166
rect 3022 2161 3023 2165
rect 3027 2161 3028 2165
rect 3022 2160 3028 2161
rect 2938 2143 2944 2144
rect 2938 2139 2939 2143
rect 2943 2139 2944 2143
rect 2938 2138 2944 2139
rect 2947 2124 2951 2125
rect 2947 2119 2951 2120
rect 2783 2114 2787 2115
rect 2783 2109 2787 2110
rect 2863 2114 2867 2115
rect 2863 2109 2867 2110
rect 2879 2114 2883 2115
rect 2879 2109 2883 2110
rect 2754 2107 2760 2108
rect 2754 2103 2755 2107
rect 2759 2103 2760 2107
rect 2754 2102 2760 2103
rect 2784 2088 2786 2109
rect 2880 2088 2882 2109
rect 2948 2108 2950 2119
rect 3024 2115 3026 2160
rect 3100 2144 3102 2170
rect 3174 2165 3180 2166
rect 3174 2161 3175 2165
rect 3179 2161 3180 2165
rect 3174 2160 3180 2161
rect 3098 2143 3104 2144
rect 3098 2139 3099 2143
rect 3103 2139 3104 2143
rect 3098 2138 3104 2139
rect 3176 2115 3178 2160
rect 3252 2144 3254 2170
rect 3260 2152 3262 2250
rect 3942 2247 3948 2248
rect 3270 2244 3276 2245
rect 3270 2240 3271 2244
rect 3275 2240 3276 2244
rect 3942 2243 3943 2247
rect 3947 2243 3948 2247
rect 3942 2242 3948 2243
rect 3270 2239 3276 2240
rect 3272 2215 3274 2239
rect 3944 2215 3946 2242
rect 3271 2214 3275 2215
rect 3271 2209 3275 2210
rect 3319 2214 3323 2215
rect 3319 2209 3323 2210
rect 3471 2214 3475 2215
rect 3471 2209 3475 2210
rect 3943 2214 3947 2215
rect 3943 2209 3947 2210
rect 3320 2185 3322 2209
rect 3472 2185 3474 2209
rect 3318 2184 3324 2185
rect 3318 2180 3319 2184
rect 3323 2180 3324 2184
rect 3318 2179 3324 2180
rect 3470 2184 3476 2185
rect 3470 2180 3471 2184
rect 3475 2180 3476 2184
rect 3944 2182 3946 2209
rect 3470 2179 3476 2180
rect 3942 2181 3948 2182
rect 3942 2177 3943 2181
rect 3947 2177 3948 2181
rect 3942 2176 3948 2177
rect 3394 2175 3400 2176
rect 3394 2171 3395 2175
rect 3399 2171 3400 2175
rect 3394 2170 3400 2171
rect 3438 2175 3444 2176
rect 3438 2171 3439 2175
rect 3443 2171 3444 2175
rect 3438 2170 3444 2171
rect 3318 2165 3324 2166
rect 3318 2161 3319 2165
rect 3323 2161 3324 2165
rect 3318 2160 3324 2161
rect 3258 2151 3264 2152
rect 3258 2147 3259 2151
rect 3263 2147 3264 2151
rect 3258 2146 3264 2147
rect 3250 2143 3256 2144
rect 3250 2139 3251 2143
rect 3255 2139 3256 2143
rect 3250 2138 3256 2139
rect 3320 2115 3322 2160
rect 3396 2144 3398 2170
rect 3394 2143 3400 2144
rect 3394 2139 3395 2143
rect 3399 2139 3400 2143
rect 3394 2138 3400 2139
rect 3440 2125 3442 2170
rect 3470 2165 3476 2166
rect 3470 2161 3471 2165
rect 3475 2161 3476 2165
rect 3470 2160 3476 2161
rect 3942 2164 3948 2165
rect 3942 2160 3943 2164
rect 3947 2160 3948 2164
rect 3439 2124 3443 2125
rect 3439 2119 3443 2120
rect 3472 2115 3474 2160
rect 3942 2159 3948 2160
rect 3944 2115 3946 2159
rect 2975 2114 2979 2115
rect 2975 2109 2979 2110
rect 3023 2114 3027 2115
rect 3023 2109 3027 2110
rect 3071 2114 3075 2115
rect 3071 2109 3075 2110
rect 3167 2114 3171 2115
rect 3167 2109 3171 2110
rect 3175 2114 3179 2115
rect 3175 2109 3179 2110
rect 3263 2114 3267 2115
rect 3263 2109 3267 2110
rect 3319 2114 3323 2115
rect 3319 2109 3323 2110
rect 3359 2114 3363 2115
rect 3359 2109 3363 2110
rect 3455 2114 3459 2115
rect 3455 2109 3459 2110
rect 3471 2114 3475 2115
rect 3471 2109 3475 2110
rect 3551 2114 3555 2115
rect 3551 2109 3555 2110
rect 3647 2114 3651 2115
rect 3647 2109 3651 2110
rect 3743 2114 3747 2115
rect 3743 2109 3747 2110
rect 3839 2114 3843 2115
rect 3839 2109 3843 2110
rect 3943 2114 3947 2115
rect 3943 2109 3947 2110
rect 2946 2107 2952 2108
rect 2946 2103 2947 2107
rect 2951 2103 2952 2107
rect 2946 2102 2952 2103
rect 2954 2107 2960 2108
rect 2954 2103 2955 2107
rect 2959 2103 2960 2107
rect 2954 2102 2960 2103
rect 2686 2087 2692 2088
rect 2686 2083 2687 2087
rect 2691 2083 2692 2087
rect 2686 2082 2692 2083
rect 2782 2087 2788 2088
rect 2782 2083 2783 2087
rect 2787 2083 2788 2087
rect 2782 2082 2788 2083
rect 2878 2087 2884 2088
rect 2878 2083 2879 2087
rect 2883 2083 2884 2087
rect 2878 2082 2884 2083
rect 2956 2080 2958 2102
rect 2976 2088 2978 2109
rect 3050 2107 3056 2108
rect 3050 2103 3051 2107
rect 3055 2103 3056 2107
rect 3050 2102 3056 2103
rect 2974 2087 2980 2088
rect 2974 2083 2975 2087
rect 2979 2083 2980 2087
rect 2974 2082 2980 2083
rect 3052 2080 3054 2102
rect 3072 2088 3074 2109
rect 3146 2107 3152 2108
rect 3146 2103 3147 2107
rect 3151 2103 3152 2107
rect 3146 2102 3152 2103
rect 3070 2087 3076 2088
rect 3070 2083 3071 2087
rect 3075 2083 3076 2087
rect 3070 2082 3076 2083
rect 3148 2080 3150 2102
rect 3168 2088 3170 2109
rect 3242 2107 3248 2108
rect 3242 2103 3243 2107
rect 3247 2103 3248 2107
rect 3242 2102 3248 2103
rect 3166 2087 3172 2088
rect 3166 2083 3167 2087
rect 3171 2083 3172 2087
rect 3166 2082 3172 2083
rect 3244 2080 3246 2102
rect 3264 2088 3266 2109
rect 3338 2107 3344 2108
rect 3338 2103 3339 2107
rect 3343 2103 3344 2107
rect 3338 2102 3344 2103
rect 3262 2087 3268 2088
rect 3262 2083 3263 2087
rect 3267 2083 3268 2087
rect 3262 2082 3268 2083
rect 3340 2080 3342 2102
rect 3360 2088 3362 2109
rect 3434 2107 3440 2108
rect 3434 2103 3435 2107
rect 3439 2103 3440 2107
rect 3434 2102 3440 2103
rect 3358 2087 3364 2088
rect 3358 2083 3359 2087
rect 3363 2083 3364 2087
rect 3358 2082 3364 2083
rect 3436 2080 3438 2102
rect 3456 2088 3458 2109
rect 3530 2107 3536 2108
rect 3530 2103 3531 2107
rect 3535 2103 3536 2107
rect 3530 2102 3536 2103
rect 3454 2087 3460 2088
rect 3454 2083 3455 2087
rect 3459 2083 3460 2087
rect 3454 2082 3460 2083
rect 3532 2080 3534 2102
rect 3552 2088 3554 2109
rect 3626 2107 3632 2108
rect 3626 2103 3627 2107
rect 3631 2103 3632 2107
rect 3626 2102 3632 2103
rect 3550 2087 3556 2088
rect 3550 2083 3551 2087
rect 3555 2083 3556 2087
rect 3550 2082 3556 2083
rect 3628 2080 3630 2102
rect 3648 2088 3650 2109
rect 3722 2107 3728 2108
rect 3722 2103 3723 2107
rect 3727 2103 3728 2107
rect 3722 2102 3728 2103
rect 3646 2087 3652 2088
rect 3646 2083 3647 2087
rect 3651 2083 3652 2087
rect 3646 2082 3652 2083
rect 3724 2080 3726 2102
rect 3744 2088 3746 2109
rect 3818 2107 3824 2108
rect 3818 2103 3819 2107
rect 3823 2103 3824 2107
rect 3818 2102 3824 2103
rect 3742 2087 3748 2088
rect 3742 2083 3743 2087
rect 3747 2083 3748 2087
rect 3742 2082 3748 2083
rect 3820 2080 3822 2102
rect 3840 2088 3842 2109
rect 3944 2089 3946 2109
rect 3942 2088 3948 2089
rect 3838 2087 3844 2088
rect 3838 2083 3839 2087
rect 3843 2083 3844 2087
rect 3942 2084 3943 2088
rect 3947 2084 3948 2088
rect 3942 2083 3948 2084
rect 3838 2082 3844 2083
rect 2474 2079 2480 2080
rect 2474 2075 2475 2079
rect 2479 2075 2480 2079
rect 2474 2074 2480 2075
rect 2570 2079 2576 2080
rect 2570 2075 2571 2079
rect 2575 2075 2576 2079
rect 2570 2074 2576 2075
rect 2666 2079 2672 2080
rect 2666 2075 2667 2079
rect 2671 2075 2672 2079
rect 2666 2074 2672 2075
rect 2954 2079 2960 2080
rect 2954 2075 2955 2079
rect 2959 2075 2960 2079
rect 2954 2074 2960 2075
rect 3050 2079 3056 2080
rect 3050 2075 3051 2079
rect 3055 2075 3056 2079
rect 3050 2074 3056 2075
rect 3146 2079 3152 2080
rect 3146 2075 3147 2079
rect 3151 2075 3152 2079
rect 3146 2074 3152 2075
rect 3242 2079 3248 2080
rect 3242 2075 3243 2079
rect 3247 2075 3248 2079
rect 3242 2074 3248 2075
rect 3338 2079 3344 2080
rect 3338 2075 3339 2079
rect 3343 2075 3344 2079
rect 3338 2074 3344 2075
rect 3434 2079 3440 2080
rect 3434 2075 3435 2079
rect 3439 2075 3440 2079
rect 3434 2074 3440 2075
rect 3530 2079 3536 2080
rect 3530 2075 3531 2079
rect 3535 2075 3536 2079
rect 3530 2074 3536 2075
rect 3626 2079 3632 2080
rect 3626 2075 3627 2079
rect 3631 2075 3632 2079
rect 3626 2074 3632 2075
rect 3722 2079 3728 2080
rect 3722 2075 3723 2079
rect 3727 2075 3728 2079
rect 3722 2074 3728 2075
rect 3818 2079 3824 2080
rect 3818 2075 3819 2079
rect 3823 2075 3824 2079
rect 3818 2074 3824 2075
rect 3914 2075 3920 2076
rect 2046 2071 2052 2072
rect 2046 2067 2047 2071
rect 2051 2067 2052 2071
rect 3914 2071 3915 2075
rect 3919 2071 3920 2075
rect 3914 2070 3920 2071
rect 3942 2071 3948 2072
rect 2046 2066 2052 2067
rect 2398 2068 2404 2069
rect 2006 2060 2012 2061
rect 1518 2059 1524 2060
rect 1518 2055 1519 2059
rect 1523 2055 1524 2059
rect 2006 2056 2007 2060
rect 2011 2056 2012 2060
rect 2006 2055 2012 2056
rect 1518 2054 1524 2055
rect 970 2051 976 2052
rect 970 2047 971 2051
rect 975 2047 976 2051
rect 970 2046 976 2047
rect 1066 2051 1072 2052
rect 1066 2047 1067 2051
rect 1071 2047 1072 2051
rect 1066 2046 1072 2047
rect 1202 2051 1208 2052
rect 1202 2047 1203 2051
rect 1207 2047 1208 2051
rect 1202 2046 1208 2047
rect 1330 2051 1336 2052
rect 1330 2047 1331 2051
rect 1335 2047 1336 2051
rect 1330 2046 1336 2047
rect 1458 2051 1464 2052
rect 1458 2047 1459 2051
rect 1463 2047 1464 2051
rect 1458 2046 1464 2047
rect 2006 2043 2012 2044
rect 990 2040 996 2041
rect 990 2036 991 2040
rect 995 2036 996 2040
rect 990 2035 996 2036
rect 1126 2040 1132 2041
rect 1126 2036 1127 2040
rect 1131 2036 1132 2040
rect 1126 2035 1132 2036
rect 1254 2040 1260 2041
rect 1254 2036 1255 2040
rect 1259 2036 1260 2040
rect 1254 2035 1260 2036
rect 1382 2040 1388 2041
rect 1382 2036 1383 2040
rect 1387 2036 1388 2040
rect 1382 2035 1388 2036
rect 1518 2040 1524 2041
rect 1518 2036 1519 2040
rect 1523 2036 1524 2040
rect 2006 2039 2007 2043
rect 2011 2039 2012 2043
rect 2048 2039 2050 2066
rect 2398 2064 2399 2068
rect 2403 2064 2404 2068
rect 2398 2063 2404 2064
rect 2494 2068 2500 2069
rect 2494 2064 2495 2068
rect 2499 2064 2500 2068
rect 2494 2063 2500 2064
rect 2590 2068 2596 2069
rect 2590 2064 2591 2068
rect 2595 2064 2596 2068
rect 2590 2063 2596 2064
rect 2686 2068 2692 2069
rect 2686 2064 2687 2068
rect 2691 2064 2692 2068
rect 2686 2063 2692 2064
rect 2782 2068 2788 2069
rect 2782 2064 2783 2068
rect 2787 2064 2788 2068
rect 2782 2063 2788 2064
rect 2878 2068 2884 2069
rect 2878 2064 2879 2068
rect 2883 2064 2884 2068
rect 2878 2063 2884 2064
rect 2974 2068 2980 2069
rect 2974 2064 2975 2068
rect 2979 2064 2980 2068
rect 2974 2063 2980 2064
rect 3070 2068 3076 2069
rect 3070 2064 3071 2068
rect 3075 2064 3076 2068
rect 3070 2063 3076 2064
rect 3166 2068 3172 2069
rect 3166 2064 3167 2068
rect 3171 2064 3172 2068
rect 3166 2063 3172 2064
rect 3262 2068 3268 2069
rect 3262 2064 3263 2068
rect 3267 2064 3268 2068
rect 3262 2063 3268 2064
rect 3358 2068 3364 2069
rect 3358 2064 3359 2068
rect 3363 2064 3364 2068
rect 3358 2063 3364 2064
rect 3454 2068 3460 2069
rect 3454 2064 3455 2068
rect 3459 2064 3460 2068
rect 3454 2063 3460 2064
rect 3550 2068 3556 2069
rect 3550 2064 3551 2068
rect 3555 2064 3556 2068
rect 3550 2063 3556 2064
rect 3646 2068 3652 2069
rect 3646 2064 3647 2068
rect 3651 2064 3652 2068
rect 3646 2063 3652 2064
rect 3742 2068 3748 2069
rect 3742 2064 3743 2068
rect 3747 2064 3748 2068
rect 3742 2063 3748 2064
rect 3838 2068 3844 2069
rect 3838 2064 3839 2068
rect 3843 2064 3844 2068
rect 3838 2063 3844 2064
rect 2400 2039 2402 2063
rect 2496 2039 2498 2063
rect 2592 2039 2594 2063
rect 2688 2039 2690 2063
rect 2784 2039 2786 2063
rect 2880 2039 2882 2063
rect 2976 2039 2978 2063
rect 3072 2039 3074 2063
rect 3168 2039 3170 2063
rect 3264 2039 3266 2063
rect 3360 2039 3362 2063
rect 3456 2039 3458 2063
rect 3552 2039 3554 2063
rect 3648 2039 3650 2063
rect 3744 2039 3746 2063
rect 3840 2039 3842 2063
rect 2006 2038 2012 2039
rect 2047 2038 2051 2039
rect 1518 2035 1524 2036
rect 992 1995 994 2035
rect 1128 1995 1130 2035
rect 1256 1995 1258 2035
rect 1384 1995 1386 2035
rect 1520 1995 1522 2035
rect 2008 1995 2010 2038
rect 2047 2033 2051 2034
rect 2191 2038 2195 2039
rect 2191 2033 2195 2034
rect 2399 2038 2403 2039
rect 2399 2033 2403 2034
rect 2495 2038 2499 2039
rect 2495 2033 2499 2034
rect 2591 2038 2595 2039
rect 2591 2033 2595 2034
rect 2647 2038 2651 2039
rect 2647 2033 2651 2034
rect 2687 2038 2691 2039
rect 2687 2033 2691 2034
rect 2783 2038 2787 2039
rect 2783 2033 2787 2034
rect 2879 2038 2883 2039
rect 2879 2033 2883 2034
rect 2919 2038 2923 2039
rect 2919 2033 2923 2034
rect 2975 2038 2979 2039
rect 2975 2033 2979 2034
rect 3071 2038 3075 2039
rect 3071 2033 3075 2034
rect 3167 2038 3171 2039
rect 3167 2033 3171 2034
rect 3215 2038 3219 2039
rect 3215 2033 3219 2034
rect 3263 2038 3267 2039
rect 3263 2033 3267 2034
rect 3359 2038 3363 2039
rect 3359 2033 3363 2034
rect 3455 2038 3459 2039
rect 3455 2033 3459 2034
rect 3527 2038 3531 2039
rect 3527 2033 3531 2034
rect 3551 2038 3555 2039
rect 3551 2033 3555 2034
rect 3647 2038 3651 2039
rect 3647 2033 3651 2034
rect 3743 2038 3747 2039
rect 3743 2033 3747 2034
rect 3839 2038 3843 2039
rect 3839 2033 3843 2034
rect 2048 2006 2050 2033
rect 2192 2009 2194 2033
rect 2400 2009 2402 2033
rect 2648 2009 2650 2033
rect 2920 2009 2922 2033
rect 3216 2009 3218 2033
rect 3528 2009 3530 2033
rect 3840 2009 3842 2033
rect 2190 2008 2196 2009
rect 2046 2005 2052 2006
rect 2046 2001 2047 2005
rect 2051 2001 2052 2005
rect 2190 2004 2191 2008
rect 2195 2004 2196 2008
rect 2190 2003 2196 2004
rect 2398 2008 2404 2009
rect 2398 2004 2399 2008
rect 2403 2004 2404 2008
rect 2398 2003 2404 2004
rect 2646 2008 2652 2009
rect 2646 2004 2647 2008
rect 2651 2004 2652 2008
rect 2646 2003 2652 2004
rect 2918 2008 2924 2009
rect 2918 2004 2919 2008
rect 2923 2004 2924 2008
rect 2918 2003 2924 2004
rect 3214 2008 3220 2009
rect 3214 2004 3215 2008
rect 3219 2004 3220 2008
rect 3214 2003 3220 2004
rect 3526 2008 3532 2009
rect 3526 2004 3527 2008
rect 3531 2004 3532 2008
rect 3526 2003 3532 2004
rect 3838 2008 3844 2009
rect 3838 2004 3839 2008
rect 3843 2004 3844 2008
rect 3838 2003 3844 2004
rect 2046 2000 2052 2001
rect 2314 1999 2320 2000
rect 2314 1995 2315 1999
rect 2319 1995 2320 1999
rect 943 1994 947 1995
rect 943 1989 947 1990
rect 991 1994 995 1995
rect 991 1989 995 1990
rect 1127 1994 1131 1995
rect 1127 1989 1131 1990
rect 1135 1994 1139 1995
rect 1135 1989 1139 1990
rect 1255 1994 1259 1995
rect 1255 1989 1259 1990
rect 1335 1994 1339 1995
rect 1335 1989 1339 1990
rect 1383 1994 1387 1995
rect 1383 1989 1387 1990
rect 1519 1994 1523 1995
rect 1519 1989 1523 1990
rect 1543 1994 1547 1995
rect 1543 1989 1547 1990
rect 2007 1994 2011 1995
rect 2314 1994 2320 1995
rect 2474 1999 2480 2000
rect 2474 1995 2475 1999
rect 2479 1995 2480 1999
rect 2474 1994 2480 1995
rect 2522 1999 2528 2000
rect 2522 1995 2523 1999
rect 2527 1995 2528 1999
rect 2522 1994 2528 1995
rect 2994 1999 3000 2000
rect 2994 1995 2995 1999
rect 2999 1995 3000 1999
rect 2994 1994 3000 1995
rect 3002 1999 3008 2000
rect 3002 1995 3003 1999
rect 3007 1995 3008 1999
rect 3002 1994 3008 1995
rect 3610 1999 3616 2000
rect 3610 1995 3611 1999
rect 3615 1995 3616 1999
rect 3610 1994 3616 1995
rect 2007 1989 2011 1990
rect 2190 1989 2196 1990
rect 944 1965 946 1989
rect 1136 1965 1138 1989
rect 1336 1965 1338 1989
rect 1544 1965 1546 1989
rect 942 1964 948 1965
rect 942 1960 943 1964
rect 947 1960 948 1964
rect 942 1959 948 1960
rect 1134 1964 1140 1965
rect 1134 1960 1135 1964
rect 1139 1960 1140 1964
rect 1134 1959 1140 1960
rect 1334 1964 1340 1965
rect 1334 1960 1335 1964
rect 1339 1960 1340 1964
rect 1334 1959 1340 1960
rect 1542 1964 1548 1965
rect 1542 1960 1543 1964
rect 1547 1960 1548 1964
rect 2008 1962 2010 1989
rect 2046 1988 2052 1989
rect 2046 1984 2047 1988
rect 2051 1984 2052 1988
rect 2190 1985 2191 1989
rect 2195 1985 2196 1989
rect 2190 1984 2196 1985
rect 2046 1983 2052 1984
rect 1542 1959 1548 1960
rect 2006 1961 2012 1962
rect 2006 1957 2007 1961
rect 2011 1957 2012 1961
rect 2006 1956 2012 1957
rect 314 1955 320 1956
rect 314 1951 315 1955
rect 319 1951 320 1955
rect 314 1950 320 1951
rect 466 1955 472 1956
rect 466 1951 467 1955
rect 471 1951 472 1955
rect 466 1950 472 1951
rect 642 1955 648 1956
rect 642 1951 643 1955
rect 647 1951 648 1955
rect 642 1950 648 1951
rect 826 1955 832 1956
rect 826 1951 827 1955
rect 831 1951 832 1955
rect 826 1950 832 1951
rect 878 1955 884 1956
rect 878 1951 879 1955
rect 883 1951 884 1955
rect 878 1950 884 1951
rect 1210 1955 1216 1956
rect 1210 1951 1211 1955
rect 1215 1951 1216 1955
rect 1210 1950 1216 1951
rect 1402 1955 1408 1956
rect 1402 1951 1403 1955
rect 1407 1951 1408 1955
rect 1402 1950 1408 1951
rect 1458 1955 1464 1956
rect 1458 1951 1459 1955
rect 1463 1951 1464 1955
rect 2048 1951 2050 1983
rect 2192 1951 2194 1984
rect 2316 1968 2318 1994
rect 2398 1989 2404 1990
rect 2398 1985 2399 1989
rect 2403 1985 2404 1989
rect 2398 1984 2404 1985
rect 2314 1967 2320 1968
rect 2314 1963 2315 1967
rect 2319 1963 2320 1967
rect 2314 1962 2320 1963
rect 2400 1951 2402 1984
rect 1458 1950 1464 1951
rect 2047 1950 2051 1951
rect 230 1945 236 1946
rect 110 1944 116 1945
rect 110 1940 111 1944
rect 115 1940 116 1944
rect 230 1941 231 1945
rect 235 1941 236 1945
rect 230 1940 236 1941
rect 110 1939 116 1940
rect 112 1919 114 1939
rect 232 1919 234 1940
rect 316 1924 318 1950
rect 390 1945 396 1946
rect 390 1941 391 1945
rect 395 1941 396 1945
rect 390 1940 396 1941
rect 306 1923 312 1924
rect 306 1919 307 1923
rect 311 1919 312 1923
rect 111 1918 115 1919
rect 111 1913 115 1914
rect 231 1918 235 1919
rect 306 1918 312 1919
rect 314 1923 320 1924
rect 314 1919 315 1923
rect 319 1919 320 1923
rect 392 1919 394 1940
rect 468 1924 470 1950
rect 566 1945 572 1946
rect 566 1941 567 1945
rect 571 1941 572 1945
rect 566 1940 572 1941
rect 466 1923 472 1924
rect 466 1919 467 1923
rect 471 1919 472 1923
rect 568 1919 570 1940
rect 644 1924 646 1950
rect 750 1945 756 1946
rect 750 1941 751 1945
rect 755 1941 756 1945
rect 750 1940 756 1941
rect 642 1923 648 1924
rect 642 1919 643 1923
rect 647 1919 648 1923
rect 752 1919 754 1940
rect 828 1924 830 1950
rect 942 1945 948 1946
rect 942 1941 943 1945
rect 947 1941 948 1945
rect 942 1940 948 1941
rect 1134 1945 1140 1946
rect 1134 1941 1135 1945
rect 1139 1941 1140 1945
rect 1134 1940 1140 1941
rect 826 1923 832 1924
rect 826 1919 827 1923
rect 831 1919 832 1923
rect 944 1919 946 1940
rect 1136 1919 1138 1940
rect 1203 1932 1207 1933
rect 1203 1927 1207 1928
rect 1204 1924 1206 1927
rect 1212 1924 1214 1950
rect 1334 1945 1340 1946
rect 1334 1941 1335 1945
rect 1339 1941 1340 1945
rect 1334 1940 1340 1941
rect 1202 1923 1208 1924
rect 1202 1919 1203 1923
rect 1207 1919 1208 1923
rect 314 1918 320 1919
rect 391 1918 395 1919
rect 466 1918 472 1919
rect 511 1918 515 1919
rect 231 1913 235 1914
rect 112 1893 114 1913
rect 110 1892 116 1893
rect 110 1888 111 1892
rect 115 1888 116 1892
rect 110 1887 116 1888
rect 308 1884 310 1918
rect 391 1913 395 1914
rect 511 1913 515 1914
rect 567 1918 571 1919
rect 567 1913 571 1914
rect 623 1918 627 1919
rect 642 1918 648 1919
rect 743 1918 747 1919
rect 623 1913 627 1914
rect 743 1913 747 1914
rect 751 1918 755 1919
rect 826 1918 832 1919
rect 863 1918 867 1919
rect 751 1913 755 1914
rect 863 1913 867 1914
rect 943 1918 947 1919
rect 943 1913 947 1914
rect 983 1918 987 1919
rect 983 1913 987 1914
rect 1103 1918 1107 1919
rect 1103 1913 1107 1914
rect 1135 1918 1139 1919
rect 1202 1918 1208 1919
rect 1210 1923 1216 1924
rect 1210 1919 1211 1923
rect 1215 1919 1216 1923
rect 1336 1919 1338 1940
rect 1210 1918 1216 1919
rect 1223 1918 1227 1919
rect 1135 1913 1139 1914
rect 1223 1913 1227 1914
rect 1335 1918 1339 1919
rect 1335 1913 1339 1914
rect 512 1892 514 1913
rect 594 1911 600 1912
rect 594 1907 595 1911
rect 599 1907 600 1911
rect 594 1906 600 1907
rect 510 1891 516 1892
rect 510 1887 511 1891
rect 515 1887 516 1891
rect 510 1886 516 1887
rect 596 1884 598 1906
rect 624 1892 626 1913
rect 744 1892 746 1913
rect 864 1892 866 1913
rect 984 1892 986 1913
rect 1104 1892 1106 1913
rect 1110 1911 1116 1912
rect 1110 1907 1111 1911
rect 1115 1907 1116 1911
rect 1110 1906 1116 1907
rect 1190 1911 1196 1912
rect 1190 1907 1191 1911
rect 1195 1907 1196 1911
rect 1190 1906 1196 1907
rect 622 1891 628 1892
rect 622 1887 623 1891
rect 627 1887 628 1891
rect 622 1886 628 1887
rect 742 1891 748 1892
rect 742 1887 743 1891
rect 747 1887 748 1891
rect 742 1886 748 1887
rect 862 1891 868 1892
rect 862 1887 863 1891
rect 867 1887 868 1891
rect 862 1886 868 1887
rect 982 1891 988 1892
rect 982 1887 983 1891
rect 987 1887 988 1891
rect 982 1886 988 1887
rect 1102 1891 1108 1892
rect 1102 1887 1103 1891
rect 1107 1887 1108 1891
rect 1102 1886 1108 1887
rect 306 1883 312 1884
rect 306 1879 307 1883
rect 311 1879 312 1883
rect 306 1878 312 1879
rect 594 1883 600 1884
rect 594 1879 595 1883
rect 599 1879 600 1883
rect 594 1878 600 1879
rect 110 1875 116 1876
rect 110 1871 111 1875
rect 115 1871 116 1875
rect 110 1870 116 1871
rect 510 1872 516 1873
rect 112 1835 114 1870
rect 510 1868 511 1872
rect 515 1868 516 1872
rect 510 1867 516 1868
rect 622 1872 628 1873
rect 622 1868 623 1872
rect 627 1868 628 1872
rect 622 1867 628 1868
rect 742 1872 748 1873
rect 742 1868 743 1872
rect 747 1868 748 1872
rect 742 1867 748 1868
rect 862 1872 868 1873
rect 862 1868 863 1872
rect 867 1868 868 1872
rect 862 1867 868 1868
rect 982 1872 988 1873
rect 982 1868 983 1872
rect 987 1868 988 1872
rect 982 1867 988 1868
rect 1102 1872 1108 1873
rect 1102 1868 1103 1872
rect 1107 1868 1108 1872
rect 1102 1867 1108 1868
rect 512 1835 514 1867
rect 624 1835 626 1867
rect 744 1835 746 1867
rect 864 1835 866 1867
rect 984 1835 986 1867
rect 1104 1835 1106 1867
rect 111 1834 115 1835
rect 111 1829 115 1830
rect 511 1834 515 1835
rect 511 1829 515 1830
rect 615 1834 619 1835
rect 615 1829 619 1830
rect 623 1834 627 1835
rect 623 1829 627 1830
rect 711 1834 715 1835
rect 711 1829 715 1830
rect 743 1834 747 1835
rect 743 1829 747 1830
rect 815 1834 819 1835
rect 815 1829 819 1830
rect 863 1834 867 1835
rect 863 1829 867 1830
rect 927 1834 931 1835
rect 927 1829 931 1830
rect 983 1834 987 1835
rect 983 1829 987 1830
rect 1039 1834 1043 1835
rect 1039 1829 1043 1830
rect 1103 1834 1107 1835
rect 1103 1829 1107 1830
rect 112 1802 114 1829
rect 616 1805 618 1829
rect 712 1805 714 1829
rect 816 1805 818 1829
rect 928 1805 930 1829
rect 1040 1805 1042 1829
rect 614 1804 620 1805
rect 110 1801 116 1802
rect 110 1797 111 1801
rect 115 1797 116 1801
rect 614 1800 615 1804
rect 619 1800 620 1804
rect 614 1799 620 1800
rect 710 1804 716 1805
rect 710 1800 711 1804
rect 715 1800 716 1804
rect 710 1799 716 1800
rect 814 1804 820 1805
rect 814 1800 815 1804
rect 819 1800 820 1804
rect 814 1799 820 1800
rect 926 1804 932 1805
rect 926 1800 927 1804
rect 931 1800 932 1804
rect 926 1799 932 1800
rect 1038 1804 1044 1805
rect 1038 1800 1039 1804
rect 1043 1800 1044 1804
rect 1038 1799 1044 1800
rect 110 1796 116 1797
rect 1112 1796 1114 1906
rect 1192 1884 1194 1906
rect 1224 1892 1226 1913
rect 1306 1911 1312 1912
rect 1306 1907 1307 1911
rect 1311 1907 1312 1911
rect 1306 1906 1312 1907
rect 1222 1891 1228 1892
rect 1222 1887 1223 1891
rect 1227 1887 1228 1891
rect 1222 1886 1228 1887
rect 1308 1884 1310 1906
rect 1336 1892 1338 1913
rect 1404 1912 1406 1950
rect 1460 1933 1462 1950
rect 1542 1945 1548 1946
rect 2047 1945 2051 1946
rect 2071 1950 2075 1951
rect 2071 1945 2075 1946
rect 2191 1950 2195 1951
rect 2191 1945 2195 1946
rect 2239 1950 2243 1951
rect 2239 1945 2243 1946
rect 2399 1950 2403 1951
rect 2399 1945 2403 1946
rect 2447 1950 2451 1951
rect 2447 1945 2451 1946
rect 1542 1941 1543 1945
rect 1547 1941 1548 1945
rect 1542 1940 1548 1941
rect 2006 1944 2012 1945
rect 2006 1940 2007 1944
rect 2011 1940 2012 1944
rect 1459 1932 1463 1933
rect 1459 1927 1463 1928
rect 1530 1923 1536 1924
rect 1530 1919 1531 1923
rect 1535 1919 1536 1923
rect 1544 1919 1546 1940
rect 2006 1939 2012 1940
rect 2008 1919 2010 1939
rect 2048 1925 2050 1945
rect 2046 1924 2052 1925
rect 2072 1924 2074 1945
rect 2146 1943 2152 1944
rect 2146 1939 2147 1943
rect 2151 1939 2152 1943
rect 2146 1938 2152 1939
rect 2046 1920 2047 1924
rect 2051 1920 2052 1924
rect 2046 1919 2052 1920
rect 2070 1923 2076 1924
rect 2070 1919 2071 1923
rect 2075 1919 2076 1923
rect 1455 1918 1459 1919
rect 1530 1918 1536 1919
rect 1543 1918 1547 1919
rect 1455 1913 1459 1914
rect 1402 1911 1408 1912
rect 1402 1907 1403 1911
rect 1407 1907 1408 1911
rect 1402 1906 1408 1907
rect 1456 1892 1458 1913
rect 1334 1891 1340 1892
rect 1334 1887 1335 1891
rect 1339 1887 1340 1891
rect 1334 1886 1340 1887
rect 1454 1891 1460 1892
rect 1454 1887 1455 1891
rect 1459 1887 1460 1891
rect 1454 1886 1460 1887
rect 1532 1884 1534 1918
rect 1543 1913 1547 1914
rect 1575 1918 1579 1919
rect 1575 1913 1579 1914
rect 1695 1918 1699 1919
rect 1695 1913 1699 1914
rect 2007 1918 2011 1919
rect 2070 1918 2076 1919
rect 2148 1916 2150 1938
rect 2240 1924 2242 1945
rect 2448 1924 2450 1945
rect 2476 1944 2478 1994
rect 2524 1976 2526 1994
rect 2646 1989 2652 1990
rect 2646 1985 2647 1989
rect 2651 1985 2652 1989
rect 2646 1984 2652 1985
rect 2918 1989 2924 1990
rect 2918 1985 2919 1989
rect 2923 1985 2924 1989
rect 2918 1984 2924 1985
rect 2522 1975 2528 1976
rect 2522 1971 2523 1975
rect 2527 1971 2528 1975
rect 2522 1970 2528 1971
rect 2648 1951 2650 1984
rect 2920 1951 2922 1984
rect 2996 1968 2998 1994
rect 3004 1976 3006 1994
rect 3214 1989 3220 1990
rect 3214 1985 3215 1989
rect 3219 1985 3220 1989
rect 3214 1984 3220 1985
rect 3526 1989 3532 1990
rect 3526 1985 3527 1989
rect 3531 1985 3532 1989
rect 3526 1984 3532 1985
rect 3002 1975 3008 1976
rect 3002 1971 3003 1975
rect 3007 1971 3008 1975
rect 3002 1970 3008 1971
rect 2994 1967 3000 1968
rect 2994 1963 2995 1967
rect 2999 1963 3000 1967
rect 2994 1962 3000 1963
rect 3216 1951 3218 1984
rect 3528 1951 3530 1984
rect 3612 1968 3614 1994
rect 3838 1989 3844 1990
rect 3838 1985 3839 1989
rect 3843 1985 3844 1989
rect 3838 1984 3844 1985
rect 3610 1967 3616 1968
rect 3610 1963 3611 1967
rect 3615 1963 3616 1967
rect 3610 1962 3616 1963
rect 3840 1951 3842 1984
rect 3916 1968 3918 2070
rect 3942 2067 3943 2071
rect 3947 2067 3948 2071
rect 3942 2066 3948 2067
rect 3944 2039 3946 2066
rect 3943 2038 3947 2039
rect 3943 2033 3947 2034
rect 3944 2006 3946 2033
rect 3942 2005 3948 2006
rect 3942 2001 3943 2005
rect 3947 2001 3948 2005
rect 3942 2000 3948 2001
rect 3942 1988 3948 1989
rect 3942 1984 3943 1988
rect 3947 1984 3948 1988
rect 3942 1983 3948 1984
rect 3914 1967 3920 1968
rect 3914 1963 3915 1967
rect 3919 1963 3920 1967
rect 3914 1962 3920 1963
rect 3944 1951 3946 1983
rect 2647 1950 2651 1951
rect 2647 1945 2651 1946
rect 2671 1950 2675 1951
rect 2671 1945 2675 1946
rect 2895 1950 2899 1951
rect 2895 1945 2899 1946
rect 2919 1950 2923 1951
rect 2919 1945 2923 1946
rect 3127 1950 3131 1951
rect 3127 1945 3131 1946
rect 3215 1950 3219 1951
rect 3215 1945 3219 1946
rect 3359 1950 3363 1951
rect 3359 1945 3363 1946
rect 3527 1950 3531 1951
rect 3527 1945 3531 1946
rect 3591 1950 3595 1951
rect 3591 1945 3595 1946
rect 3831 1950 3835 1951
rect 3831 1945 3835 1946
rect 3839 1950 3843 1951
rect 3839 1945 3843 1946
rect 3943 1950 3947 1951
rect 3943 1945 3947 1946
rect 2474 1943 2480 1944
rect 2474 1939 2475 1943
rect 2479 1939 2480 1943
rect 2474 1938 2480 1939
rect 2522 1943 2528 1944
rect 2522 1939 2523 1943
rect 2527 1939 2528 1943
rect 2522 1938 2528 1939
rect 2238 1923 2244 1924
rect 2238 1919 2239 1923
rect 2243 1919 2244 1923
rect 2238 1918 2244 1919
rect 2446 1923 2452 1924
rect 2446 1919 2447 1923
rect 2451 1919 2452 1923
rect 2446 1918 2452 1919
rect 2524 1916 2526 1938
rect 2672 1924 2674 1945
rect 2746 1943 2752 1944
rect 2746 1939 2747 1943
rect 2751 1939 2752 1943
rect 2746 1938 2752 1939
rect 2670 1923 2676 1924
rect 2670 1919 2671 1923
rect 2675 1919 2676 1923
rect 2670 1918 2676 1919
rect 2748 1916 2750 1938
rect 2778 1935 2784 1936
rect 2778 1931 2779 1935
rect 2783 1931 2784 1935
rect 2778 1930 2784 1931
rect 2780 1916 2782 1930
rect 2896 1924 2898 1945
rect 3128 1924 3130 1945
rect 3360 1924 3362 1945
rect 3442 1943 3448 1944
rect 3442 1939 3443 1943
rect 3447 1939 3448 1943
rect 3442 1938 3448 1939
rect 2894 1923 2900 1924
rect 2894 1919 2895 1923
rect 2899 1919 2900 1923
rect 2894 1918 2900 1919
rect 3126 1923 3132 1924
rect 3126 1919 3127 1923
rect 3131 1919 3132 1923
rect 3126 1918 3132 1919
rect 3358 1923 3364 1924
rect 3358 1919 3359 1923
rect 3363 1919 3364 1923
rect 3358 1918 3364 1919
rect 3444 1916 3446 1938
rect 3592 1924 3594 1945
rect 3654 1943 3660 1944
rect 3654 1939 3655 1943
rect 3659 1939 3660 1943
rect 3654 1938 3660 1939
rect 3590 1923 3596 1924
rect 3590 1919 3591 1923
rect 3595 1919 3596 1923
rect 3590 1918 3596 1919
rect 2007 1913 2011 1914
rect 2146 1915 2152 1916
rect 1576 1892 1578 1913
rect 1696 1892 1698 1913
rect 1714 1911 1720 1912
rect 1714 1907 1715 1911
rect 1719 1907 1720 1911
rect 1714 1906 1720 1907
rect 1574 1891 1580 1892
rect 1574 1887 1575 1891
rect 1579 1887 1580 1891
rect 1574 1886 1580 1887
rect 1694 1891 1700 1892
rect 1694 1887 1695 1891
rect 1699 1887 1700 1891
rect 1694 1886 1700 1887
rect 1190 1883 1196 1884
rect 1178 1879 1184 1880
rect 1178 1875 1179 1879
rect 1183 1875 1184 1879
rect 1190 1879 1191 1883
rect 1195 1879 1196 1883
rect 1190 1878 1196 1879
rect 1306 1883 1312 1884
rect 1306 1879 1307 1883
rect 1311 1879 1312 1883
rect 1306 1878 1312 1879
rect 1530 1883 1536 1884
rect 1530 1879 1531 1883
rect 1535 1879 1536 1883
rect 1530 1878 1536 1879
rect 1178 1874 1184 1875
rect 1159 1834 1163 1835
rect 1159 1829 1163 1830
rect 1160 1805 1162 1829
rect 1158 1804 1164 1805
rect 1158 1800 1159 1804
rect 1163 1800 1164 1804
rect 1158 1799 1164 1800
rect 690 1795 696 1796
rect 690 1791 691 1795
rect 695 1791 696 1795
rect 690 1790 696 1791
rect 786 1795 792 1796
rect 786 1791 787 1795
rect 791 1791 792 1795
rect 786 1790 792 1791
rect 890 1795 896 1796
rect 890 1791 891 1795
rect 895 1791 896 1795
rect 890 1790 896 1791
rect 1002 1795 1008 1796
rect 1002 1791 1003 1795
rect 1007 1791 1008 1795
rect 1002 1790 1008 1791
rect 1110 1795 1116 1796
rect 1110 1791 1111 1795
rect 1115 1791 1116 1795
rect 1110 1790 1116 1791
rect 614 1785 620 1786
rect 110 1784 116 1785
rect 110 1780 111 1784
rect 115 1780 116 1784
rect 614 1781 615 1785
rect 619 1781 620 1785
rect 614 1780 620 1781
rect 110 1779 116 1780
rect 112 1759 114 1779
rect 616 1759 618 1780
rect 692 1764 694 1790
rect 710 1785 716 1786
rect 710 1781 711 1785
rect 715 1781 716 1785
rect 710 1780 716 1781
rect 682 1763 688 1764
rect 682 1759 683 1763
rect 687 1759 688 1763
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 367 1758 371 1759
rect 367 1753 371 1754
rect 495 1758 499 1759
rect 495 1753 499 1754
rect 615 1758 619 1759
rect 615 1753 619 1754
rect 639 1758 643 1759
rect 682 1758 688 1759
rect 690 1763 696 1764
rect 690 1759 691 1763
rect 695 1759 696 1763
rect 712 1759 714 1780
rect 788 1764 790 1790
rect 814 1785 820 1786
rect 814 1781 815 1785
rect 819 1781 820 1785
rect 814 1780 820 1781
rect 786 1763 792 1764
rect 786 1759 787 1763
rect 791 1759 792 1763
rect 816 1759 818 1780
rect 892 1764 894 1790
rect 926 1785 932 1786
rect 926 1781 927 1785
rect 931 1781 932 1785
rect 926 1780 932 1781
rect 890 1763 896 1764
rect 890 1759 891 1763
rect 895 1759 896 1763
rect 928 1759 930 1780
rect 1004 1764 1006 1790
rect 1038 1785 1044 1786
rect 1038 1781 1039 1785
rect 1043 1781 1044 1785
rect 1038 1780 1044 1781
rect 1158 1785 1164 1786
rect 1158 1781 1159 1785
rect 1163 1781 1164 1785
rect 1158 1780 1164 1781
rect 1002 1763 1008 1764
rect 1002 1759 1003 1763
rect 1007 1759 1008 1763
rect 1040 1759 1042 1780
rect 1160 1759 1162 1780
rect 1180 1764 1182 1874
rect 1222 1872 1228 1873
rect 1222 1868 1223 1872
rect 1227 1868 1228 1872
rect 1222 1867 1228 1868
rect 1334 1872 1340 1873
rect 1334 1868 1335 1872
rect 1339 1868 1340 1872
rect 1334 1867 1340 1868
rect 1454 1872 1460 1873
rect 1454 1868 1455 1872
rect 1459 1868 1460 1872
rect 1454 1867 1460 1868
rect 1574 1872 1580 1873
rect 1574 1868 1575 1872
rect 1579 1868 1580 1872
rect 1574 1867 1580 1868
rect 1694 1872 1700 1873
rect 1694 1868 1695 1872
rect 1699 1868 1700 1872
rect 1694 1867 1700 1868
rect 1224 1835 1226 1867
rect 1336 1835 1338 1867
rect 1456 1835 1458 1867
rect 1576 1835 1578 1867
rect 1696 1835 1698 1867
rect 1223 1834 1227 1835
rect 1223 1829 1227 1830
rect 1279 1834 1283 1835
rect 1279 1829 1283 1830
rect 1335 1834 1339 1835
rect 1335 1829 1339 1830
rect 1399 1834 1403 1835
rect 1399 1829 1403 1830
rect 1455 1834 1459 1835
rect 1455 1829 1459 1830
rect 1519 1834 1523 1835
rect 1519 1829 1523 1830
rect 1575 1834 1579 1835
rect 1575 1829 1579 1830
rect 1639 1834 1643 1835
rect 1639 1829 1643 1830
rect 1695 1834 1699 1835
rect 1695 1829 1699 1830
rect 1280 1805 1282 1829
rect 1400 1805 1402 1829
rect 1520 1805 1522 1829
rect 1640 1805 1642 1829
rect 1278 1804 1284 1805
rect 1278 1800 1279 1804
rect 1283 1800 1284 1804
rect 1278 1799 1284 1800
rect 1398 1804 1404 1805
rect 1398 1800 1399 1804
rect 1403 1800 1404 1804
rect 1398 1799 1404 1800
rect 1518 1804 1524 1805
rect 1518 1800 1519 1804
rect 1523 1800 1524 1804
rect 1518 1799 1524 1800
rect 1638 1804 1644 1805
rect 1638 1800 1639 1804
rect 1643 1800 1644 1804
rect 1638 1799 1644 1800
rect 1716 1796 1718 1906
rect 2008 1893 2010 1913
rect 2146 1911 2147 1915
rect 2151 1911 2152 1915
rect 2522 1915 2528 1916
rect 2146 1910 2152 1911
rect 2314 1911 2320 1912
rect 2046 1907 2052 1908
rect 2046 1903 2047 1907
rect 2051 1903 2052 1907
rect 2314 1907 2315 1911
rect 2319 1907 2320 1911
rect 2522 1911 2523 1915
rect 2527 1911 2528 1915
rect 2522 1910 2528 1911
rect 2746 1915 2752 1916
rect 2746 1911 2747 1915
rect 2751 1911 2752 1915
rect 2746 1910 2752 1911
rect 2778 1915 2784 1916
rect 2778 1911 2779 1915
rect 2783 1911 2784 1915
rect 2778 1910 2784 1911
rect 3442 1915 3448 1916
rect 3442 1911 3443 1915
rect 3447 1911 3448 1915
rect 3442 1910 3448 1911
rect 2314 1906 2320 1907
rect 2046 1902 2052 1903
rect 2070 1904 2076 1905
rect 2006 1892 2012 1893
rect 2006 1888 2007 1892
rect 2011 1888 2012 1892
rect 2006 1887 2012 1888
rect 2006 1875 2012 1876
rect 2048 1875 2050 1902
rect 2070 1900 2071 1904
rect 2075 1900 2076 1904
rect 2070 1899 2076 1900
rect 2238 1904 2244 1905
rect 2238 1900 2239 1904
rect 2243 1900 2244 1904
rect 2238 1899 2244 1900
rect 2072 1875 2074 1899
rect 2240 1875 2242 1899
rect 2006 1871 2007 1875
rect 2011 1871 2012 1875
rect 2006 1870 2012 1871
rect 2047 1874 2051 1875
rect 2008 1835 2010 1870
rect 2047 1869 2051 1870
rect 2071 1874 2075 1875
rect 2071 1869 2075 1870
rect 2199 1874 2203 1875
rect 2199 1869 2203 1870
rect 2239 1874 2243 1875
rect 2239 1869 2243 1870
rect 2048 1842 2050 1869
rect 2072 1845 2074 1869
rect 2200 1845 2202 1869
rect 2070 1844 2076 1845
rect 2046 1841 2052 1842
rect 2046 1837 2047 1841
rect 2051 1837 2052 1841
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2070 1839 2076 1840
rect 2198 1844 2204 1845
rect 2198 1840 2199 1844
rect 2203 1840 2204 1844
rect 2198 1839 2204 1840
rect 2046 1836 2052 1837
rect 2138 1835 2144 1836
rect 2007 1834 2011 1835
rect 2138 1831 2139 1835
rect 2143 1831 2144 1835
rect 2138 1830 2144 1831
rect 2154 1835 2160 1836
rect 2154 1831 2155 1835
rect 2159 1831 2160 1835
rect 2154 1830 2160 1831
rect 2007 1829 2011 1830
rect 2008 1802 2010 1829
rect 2070 1825 2076 1826
rect 2046 1824 2052 1825
rect 2046 1820 2047 1824
rect 2051 1820 2052 1824
rect 2070 1821 2071 1825
rect 2075 1821 2076 1825
rect 2070 1820 2076 1821
rect 2046 1819 2052 1820
rect 2006 1801 2012 1802
rect 2006 1797 2007 1801
rect 2011 1797 2012 1801
rect 2006 1796 2012 1797
rect 1234 1795 1240 1796
rect 1234 1791 1235 1795
rect 1239 1791 1240 1795
rect 1234 1790 1240 1791
rect 1354 1795 1360 1796
rect 1354 1791 1355 1795
rect 1359 1791 1360 1795
rect 1354 1790 1360 1791
rect 1390 1795 1396 1796
rect 1390 1791 1391 1795
rect 1395 1791 1396 1795
rect 1390 1790 1396 1791
rect 1594 1795 1600 1796
rect 1594 1791 1595 1795
rect 1599 1791 1600 1795
rect 1594 1790 1600 1791
rect 1714 1795 1720 1796
rect 2048 1795 2050 1819
rect 2072 1795 2074 1820
rect 1714 1791 1715 1795
rect 1719 1791 1720 1795
rect 1714 1790 1720 1791
rect 2047 1794 2051 1795
rect 1236 1764 1238 1790
rect 1278 1785 1284 1786
rect 1278 1781 1279 1785
rect 1283 1781 1284 1785
rect 1278 1780 1284 1781
rect 1178 1763 1184 1764
rect 1178 1759 1179 1763
rect 1183 1759 1184 1763
rect 690 1758 696 1759
rect 711 1758 715 1759
rect 786 1758 792 1759
rect 799 1758 803 1759
rect 639 1753 643 1754
rect 112 1733 114 1753
rect 110 1732 116 1733
rect 368 1732 370 1753
rect 434 1751 440 1752
rect 434 1747 435 1751
rect 439 1747 440 1751
rect 434 1746 440 1747
rect 442 1751 448 1752
rect 442 1747 443 1751
rect 447 1747 448 1751
rect 442 1746 448 1747
rect 110 1728 111 1732
rect 115 1728 116 1732
rect 110 1727 116 1728
rect 366 1731 372 1732
rect 366 1727 367 1731
rect 371 1727 372 1731
rect 366 1726 372 1727
rect 110 1715 116 1716
rect 110 1711 111 1715
rect 115 1711 116 1715
rect 110 1710 116 1711
rect 366 1712 372 1713
rect 112 1679 114 1710
rect 366 1708 367 1712
rect 371 1708 372 1712
rect 366 1707 372 1708
rect 368 1679 370 1707
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 135 1678 139 1679
rect 135 1673 139 1674
rect 247 1678 251 1679
rect 247 1673 251 1674
rect 367 1678 371 1679
rect 367 1673 371 1674
rect 399 1678 403 1679
rect 399 1673 403 1674
rect 112 1646 114 1673
rect 136 1649 138 1673
rect 248 1649 250 1673
rect 400 1649 402 1673
rect 436 1656 438 1746
rect 444 1724 446 1746
rect 496 1732 498 1753
rect 570 1751 576 1752
rect 570 1747 571 1751
rect 575 1747 576 1751
rect 570 1746 576 1747
rect 494 1731 500 1732
rect 494 1727 495 1731
rect 499 1727 500 1731
rect 494 1726 500 1727
rect 572 1724 574 1746
rect 640 1732 642 1753
rect 684 1741 686 1758
rect 711 1753 715 1754
rect 799 1753 803 1754
rect 815 1758 819 1759
rect 890 1758 896 1759
rect 927 1758 931 1759
rect 815 1753 819 1754
rect 927 1753 931 1754
rect 967 1758 971 1759
rect 1002 1758 1008 1759
rect 1039 1758 1043 1759
rect 967 1753 971 1754
rect 1039 1753 1043 1754
rect 1143 1758 1147 1759
rect 1143 1753 1147 1754
rect 1159 1758 1163 1759
rect 1178 1758 1184 1759
rect 1234 1763 1240 1764
rect 1234 1759 1235 1763
rect 1239 1759 1240 1763
rect 1280 1759 1282 1780
rect 1356 1764 1358 1790
rect 1354 1763 1360 1764
rect 1354 1759 1355 1763
rect 1359 1759 1360 1763
rect 1234 1758 1240 1759
rect 1279 1758 1283 1759
rect 1159 1753 1163 1754
rect 1279 1753 1283 1754
rect 1327 1758 1331 1759
rect 1354 1758 1360 1759
rect 1327 1753 1331 1754
rect 770 1751 776 1752
rect 770 1747 771 1751
rect 775 1747 776 1751
rect 770 1746 776 1747
rect 683 1740 687 1741
rect 683 1735 687 1736
rect 638 1731 644 1732
rect 638 1727 639 1731
rect 643 1727 644 1731
rect 638 1726 644 1727
rect 772 1724 774 1746
rect 800 1732 802 1753
rect 874 1751 880 1752
rect 874 1747 875 1751
rect 879 1747 880 1751
rect 874 1746 880 1747
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 876 1724 878 1746
rect 919 1740 923 1741
rect 919 1735 923 1736
rect 920 1724 922 1735
rect 968 1732 970 1753
rect 1144 1732 1146 1753
rect 1328 1732 1330 1753
rect 1392 1752 1394 1790
rect 1398 1785 1404 1786
rect 1398 1781 1399 1785
rect 1403 1781 1404 1785
rect 1398 1780 1404 1781
rect 1518 1785 1524 1786
rect 1518 1781 1519 1785
rect 1523 1781 1524 1785
rect 1518 1780 1524 1781
rect 1400 1759 1402 1780
rect 1520 1759 1522 1780
rect 1596 1764 1598 1790
rect 2047 1789 2051 1790
rect 2071 1794 2075 1795
rect 2071 1789 2075 1790
rect 1638 1785 1644 1786
rect 1638 1781 1639 1785
rect 1643 1781 1644 1785
rect 1638 1780 1644 1781
rect 2006 1784 2012 1785
rect 2006 1780 2007 1784
rect 2011 1780 2012 1784
rect 1586 1763 1592 1764
rect 1586 1759 1587 1763
rect 1591 1759 1592 1763
rect 1399 1758 1403 1759
rect 1399 1753 1403 1754
rect 1511 1758 1515 1759
rect 1511 1753 1515 1754
rect 1519 1758 1523 1759
rect 1586 1758 1592 1759
rect 1594 1763 1600 1764
rect 1594 1759 1595 1763
rect 1599 1759 1600 1763
rect 1640 1759 1642 1780
rect 2006 1779 2012 1780
rect 2008 1759 2010 1779
rect 2048 1769 2050 1789
rect 2046 1768 2052 1769
rect 2072 1768 2074 1789
rect 2140 1788 2142 1830
rect 2156 1804 2158 1830
rect 2198 1825 2204 1826
rect 2198 1821 2199 1825
rect 2203 1821 2204 1825
rect 2198 1820 2204 1821
rect 2154 1803 2160 1804
rect 2154 1799 2155 1803
rect 2159 1799 2160 1803
rect 2154 1798 2160 1799
rect 2200 1795 2202 1820
rect 2316 1804 2318 1906
rect 2446 1904 2452 1905
rect 2446 1900 2447 1904
rect 2451 1900 2452 1904
rect 2446 1899 2452 1900
rect 2670 1904 2676 1905
rect 2670 1900 2671 1904
rect 2675 1900 2676 1904
rect 2670 1899 2676 1900
rect 2894 1904 2900 1905
rect 2894 1900 2895 1904
rect 2899 1900 2900 1904
rect 2894 1899 2900 1900
rect 3126 1904 3132 1905
rect 3126 1900 3127 1904
rect 3131 1900 3132 1904
rect 3126 1899 3132 1900
rect 3358 1904 3364 1905
rect 3358 1900 3359 1904
rect 3363 1900 3364 1904
rect 3358 1899 3364 1900
rect 3590 1904 3596 1905
rect 3590 1900 3591 1904
rect 3595 1900 3596 1904
rect 3590 1899 3596 1900
rect 2448 1875 2450 1899
rect 2672 1875 2674 1899
rect 2896 1875 2898 1899
rect 3128 1875 3130 1899
rect 3360 1875 3362 1899
rect 3592 1875 3594 1899
rect 2367 1874 2371 1875
rect 2367 1869 2371 1870
rect 2447 1874 2451 1875
rect 2447 1869 2451 1870
rect 2543 1874 2547 1875
rect 2543 1869 2547 1870
rect 2671 1874 2675 1875
rect 2671 1869 2675 1870
rect 2719 1874 2723 1875
rect 2719 1869 2723 1870
rect 2887 1874 2891 1875
rect 2887 1869 2891 1870
rect 2895 1874 2899 1875
rect 2895 1869 2899 1870
rect 3039 1874 3043 1875
rect 3039 1869 3043 1870
rect 3127 1874 3131 1875
rect 3127 1869 3131 1870
rect 3183 1874 3187 1875
rect 3183 1869 3187 1870
rect 3319 1874 3323 1875
rect 3319 1869 3323 1870
rect 3359 1874 3363 1875
rect 3359 1869 3363 1870
rect 3455 1874 3459 1875
rect 3455 1869 3459 1870
rect 3583 1874 3587 1875
rect 3583 1869 3587 1870
rect 3591 1874 3595 1875
rect 3591 1869 3595 1870
rect 2368 1845 2370 1869
rect 2544 1845 2546 1869
rect 2720 1845 2722 1869
rect 2888 1845 2890 1869
rect 3040 1845 3042 1869
rect 3184 1845 3186 1869
rect 3320 1845 3322 1869
rect 3456 1845 3458 1869
rect 3584 1845 3586 1869
rect 2366 1844 2372 1845
rect 2366 1840 2367 1844
rect 2371 1840 2372 1844
rect 2366 1839 2372 1840
rect 2542 1844 2548 1845
rect 2542 1840 2543 1844
rect 2547 1840 2548 1844
rect 2542 1839 2548 1840
rect 2718 1844 2724 1845
rect 2718 1840 2719 1844
rect 2723 1840 2724 1844
rect 2718 1839 2724 1840
rect 2886 1844 2892 1845
rect 2886 1840 2887 1844
rect 2891 1840 2892 1844
rect 2886 1839 2892 1840
rect 3038 1844 3044 1845
rect 3038 1840 3039 1844
rect 3043 1840 3044 1844
rect 3038 1839 3044 1840
rect 3182 1844 3188 1845
rect 3182 1840 3183 1844
rect 3187 1840 3188 1844
rect 3182 1839 3188 1840
rect 3318 1844 3324 1845
rect 3318 1840 3319 1844
rect 3323 1840 3324 1844
rect 3318 1839 3324 1840
rect 3454 1844 3460 1845
rect 3454 1840 3455 1844
rect 3459 1840 3460 1844
rect 3454 1839 3460 1840
rect 3582 1844 3588 1845
rect 3582 1840 3583 1844
rect 3587 1840 3588 1844
rect 3582 1839 3588 1840
rect 3656 1836 3658 1938
rect 3832 1924 3834 1945
rect 3944 1925 3946 1945
rect 3942 1924 3948 1925
rect 3830 1923 3836 1924
rect 3830 1919 3831 1923
rect 3835 1919 3836 1923
rect 3942 1920 3943 1924
rect 3947 1920 3948 1924
rect 3942 1919 3948 1920
rect 3830 1918 3836 1919
rect 3914 1911 3920 1912
rect 3914 1907 3915 1911
rect 3919 1907 3920 1911
rect 3914 1906 3920 1907
rect 3942 1907 3948 1908
rect 3830 1904 3836 1905
rect 3830 1900 3831 1904
rect 3835 1900 3836 1904
rect 3830 1899 3836 1900
rect 3832 1875 3834 1899
rect 3711 1874 3715 1875
rect 3711 1869 3715 1870
rect 3831 1874 3835 1875
rect 3831 1869 3835 1870
rect 3839 1874 3843 1875
rect 3839 1869 3843 1870
rect 3712 1845 3714 1869
rect 3840 1845 3842 1869
rect 3710 1844 3716 1845
rect 3710 1840 3711 1844
rect 3715 1840 3716 1844
rect 3710 1839 3716 1840
rect 3838 1844 3844 1845
rect 3838 1840 3839 1844
rect 3843 1840 3844 1844
rect 3838 1839 3844 1840
rect 2442 1835 2448 1836
rect 2442 1831 2443 1835
rect 2447 1831 2448 1835
rect 2442 1830 2448 1831
rect 2618 1835 2624 1836
rect 2618 1831 2619 1835
rect 2623 1831 2624 1835
rect 2618 1830 2624 1831
rect 2658 1835 2664 1836
rect 2658 1831 2659 1835
rect 2663 1831 2664 1835
rect 2658 1830 2664 1831
rect 2962 1835 2968 1836
rect 2962 1831 2963 1835
rect 2967 1831 2968 1835
rect 2962 1830 2968 1831
rect 3114 1835 3120 1836
rect 3114 1831 3115 1835
rect 3119 1831 3120 1835
rect 3114 1830 3120 1831
rect 3258 1835 3264 1836
rect 3258 1831 3259 1835
rect 3263 1831 3264 1835
rect 3258 1830 3264 1831
rect 3394 1835 3400 1836
rect 3394 1831 3395 1835
rect 3399 1831 3400 1835
rect 3394 1830 3400 1831
rect 3522 1835 3528 1836
rect 3522 1831 3523 1835
rect 3527 1831 3528 1835
rect 3522 1830 3528 1831
rect 3654 1835 3660 1836
rect 3654 1831 3655 1835
rect 3659 1831 3660 1835
rect 3654 1830 3660 1831
rect 3666 1835 3672 1836
rect 3666 1831 3667 1835
rect 3671 1831 3672 1835
rect 3666 1830 3672 1831
rect 3906 1835 3912 1836
rect 3906 1831 3907 1835
rect 3911 1831 3912 1835
rect 3906 1830 3912 1831
rect 2366 1825 2372 1826
rect 2366 1821 2367 1825
rect 2371 1821 2372 1825
rect 2366 1820 2372 1821
rect 2314 1803 2320 1804
rect 2314 1799 2315 1803
rect 2319 1799 2320 1803
rect 2314 1798 2320 1799
rect 2368 1795 2370 1820
rect 2444 1804 2446 1830
rect 2542 1825 2548 1826
rect 2542 1821 2543 1825
rect 2547 1821 2548 1825
rect 2542 1820 2548 1821
rect 2442 1803 2448 1804
rect 2442 1799 2443 1803
rect 2447 1799 2448 1803
rect 2442 1798 2448 1799
rect 2544 1795 2546 1820
rect 2620 1804 2622 1830
rect 2660 1812 2662 1830
rect 2718 1825 2724 1826
rect 2718 1821 2719 1825
rect 2723 1821 2724 1825
rect 2718 1820 2724 1821
rect 2886 1825 2892 1826
rect 2886 1821 2887 1825
rect 2891 1821 2892 1825
rect 2886 1820 2892 1821
rect 2658 1811 2664 1812
rect 2658 1807 2659 1811
rect 2663 1807 2664 1811
rect 2658 1806 2664 1807
rect 2618 1803 2624 1804
rect 2618 1799 2619 1803
rect 2623 1799 2624 1803
rect 2618 1798 2624 1799
rect 2720 1795 2722 1820
rect 2888 1795 2890 1820
rect 2964 1804 2966 1830
rect 3038 1825 3044 1826
rect 3038 1821 3039 1825
rect 3043 1821 3044 1825
rect 3038 1820 3044 1821
rect 2962 1803 2968 1804
rect 2962 1799 2963 1803
rect 2967 1799 2968 1803
rect 2962 1798 2968 1799
rect 3040 1795 3042 1820
rect 3116 1804 3118 1830
rect 3182 1825 3188 1826
rect 3182 1821 3183 1825
rect 3187 1821 3188 1825
rect 3182 1820 3188 1821
rect 3114 1803 3120 1804
rect 3114 1799 3115 1803
rect 3119 1799 3120 1803
rect 3114 1798 3120 1799
rect 3184 1795 3186 1820
rect 3260 1804 3262 1830
rect 3318 1825 3324 1826
rect 3318 1821 3319 1825
rect 3323 1821 3324 1825
rect 3318 1820 3324 1821
rect 3258 1803 3264 1804
rect 3258 1799 3259 1803
rect 3263 1799 3264 1803
rect 3258 1798 3264 1799
rect 3320 1795 3322 1820
rect 3396 1804 3398 1830
rect 3454 1825 3460 1826
rect 3454 1821 3455 1825
rect 3459 1821 3460 1825
rect 3454 1820 3460 1821
rect 3394 1803 3400 1804
rect 3394 1799 3395 1803
rect 3399 1799 3400 1803
rect 3394 1798 3400 1799
rect 3456 1795 3458 1820
rect 2183 1794 2187 1795
rect 2183 1789 2187 1790
rect 2199 1794 2203 1795
rect 2199 1789 2203 1790
rect 2327 1794 2331 1795
rect 2327 1789 2331 1790
rect 2367 1794 2371 1795
rect 2367 1789 2371 1790
rect 2487 1794 2491 1795
rect 2487 1789 2491 1790
rect 2543 1794 2547 1795
rect 2543 1789 2547 1790
rect 2655 1794 2659 1795
rect 2655 1789 2659 1790
rect 2719 1794 2723 1795
rect 2719 1789 2723 1790
rect 2831 1794 2835 1795
rect 2831 1789 2835 1790
rect 2887 1794 2891 1795
rect 2887 1789 2891 1790
rect 3023 1794 3027 1795
rect 3023 1789 3027 1790
rect 3039 1794 3043 1795
rect 3039 1789 3043 1790
rect 3183 1794 3187 1795
rect 3183 1789 3187 1790
rect 3223 1794 3227 1795
rect 3223 1789 3227 1790
rect 3319 1794 3323 1795
rect 3319 1789 3323 1790
rect 3431 1794 3435 1795
rect 3431 1789 3435 1790
rect 3455 1794 3459 1795
rect 3455 1789 3459 1790
rect 2138 1787 2144 1788
rect 2138 1783 2139 1787
rect 2143 1783 2144 1787
rect 2138 1782 2144 1783
rect 2146 1787 2152 1788
rect 2146 1783 2147 1787
rect 2151 1783 2152 1787
rect 2146 1782 2152 1783
rect 2046 1764 2047 1768
rect 2051 1764 2052 1768
rect 2046 1763 2052 1764
rect 2070 1767 2076 1768
rect 2070 1763 2071 1767
rect 2075 1763 2076 1767
rect 2070 1762 2076 1763
rect 2148 1760 2150 1782
rect 2184 1768 2186 1789
rect 2258 1787 2264 1788
rect 2258 1783 2259 1787
rect 2263 1783 2264 1787
rect 2258 1782 2264 1783
rect 2182 1767 2188 1768
rect 2182 1763 2183 1767
rect 2187 1763 2188 1767
rect 2182 1762 2188 1763
rect 2260 1760 2262 1782
rect 2328 1768 2330 1789
rect 2402 1787 2408 1788
rect 2402 1783 2403 1787
rect 2407 1783 2408 1787
rect 2402 1782 2408 1783
rect 2326 1767 2332 1768
rect 2326 1763 2327 1767
rect 2331 1763 2332 1767
rect 2326 1762 2332 1763
rect 2404 1760 2406 1782
rect 2488 1768 2490 1789
rect 2562 1787 2568 1788
rect 2562 1783 2563 1787
rect 2567 1783 2568 1787
rect 2562 1782 2568 1783
rect 2486 1767 2492 1768
rect 2486 1763 2487 1767
rect 2491 1763 2492 1767
rect 2486 1762 2492 1763
rect 2564 1760 2566 1782
rect 2656 1768 2658 1789
rect 2832 1768 2834 1789
rect 3024 1768 3026 1789
rect 3106 1787 3112 1788
rect 3106 1783 3107 1787
rect 3111 1783 3112 1787
rect 3106 1782 3112 1783
rect 2654 1767 2660 1768
rect 2654 1763 2655 1767
rect 2659 1763 2660 1767
rect 2654 1762 2660 1763
rect 2830 1767 2836 1768
rect 2830 1763 2831 1767
rect 2835 1763 2836 1767
rect 2830 1762 2836 1763
rect 3022 1767 3028 1768
rect 3022 1763 3023 1767
rect 3027 1763 3028 1767
rect 3022 1762 3028 1763
rect 3108 1760 3110 1782
rect 3224 1768 3226 1789
rect 3306 1787 3312 1788
rect 3306 1783 3307 1787
rect 3311 1783 3312 1787
rect 3306 1782 3312 1783
rect 3222 1767 3228 1768
rect 3222 1763 3223 1767
rect 3227 1763 3228 1767
rect 3222 1762 3228 1763
rect 3308 1760 3310 1782
rect 3432 1768 3434 1789
rect 3524 1788 3526 1830
rect 3582 1825 3588 1826
rect 3582 1821 3583 1825
rect 3587 1821 3588 1825
rect 3582 1820 3588 1821
rect 3584 1795 3586 1820
rect 3668 1804 3670 1830
rect 3710 1825 3716 1826
rect 3710 1821 3711 1825
rect 3715 1821 3716 1825
rect 3710 1820 3716 1821
rect 3838 1825 3844 1826
rect 3838 1821 3839 1825
rect 3843 1821 3844 1825
rect 3838 1820 3844 1821
rect 3666 1803 3672 1804
rect 3666 1799 3667 1803
rect 3671 1799 3672 1803
rect 3666 1798 3672 1799
rect 3712 1795 3714 1820
rect 3722 1803 3728 1804
rect 3722 1799 3723 1803
rect 3727 1799 3728 1803
rect 3722 1798 3728 1799
rect 3583 1794 3587 1795
rect 3583 1789 3587 1790
rect 3647 1794 3651 1795
rect 3647 1789 3651 1790
rect 3711 1794 3715 1795
rect 3711 1789 3715 1790
rect 3522 1787 3528 1788
rect 3522 1783 3523 1787
rect 3527 1783 3528 1787
rect 3522 1782 3528 1783
rect 3648 1768 3650 1789
rect 3430 1767 3436 1768
rect 3430 1763 3431 1767
rect 3435 1763 3436 1767
rect 3430 1762 3436 1763
rect 3646 1767 3652 1768
rect 3646 1763 3647 1767
rect 3651 1763 3652 1767
rect 3646 1762 3652 1763
rect 3724 1760 3726 1798
rect 3840 1795 3842 1820
rect 3839 1794 3843 1795
rect 3839 1789 3843 1790
rect 3738 1787 3744 1788
rect 3738 1783 3739 1787
rect 3743 1783 3744 1787
rect 3738 1782 3744 1783
rect 2146 1759 2152 1760
rect 1594 1758 1600 1759
rect 1639 1758 1643 1759
rect 1519 1753 1523 1754
rect 1390 1751 1396 1752
rect 1390 1747 1391 1751
rect 1395 1747 1396 1751
rect 1390 1746 1396 1747
rect 1512 1732 1514 1753
rect 966 1731 972 1732
rect 966 1727 967 1731
rect 971 1727 972 1731
rect 966 1726 972 1727
rect 1142 1731 1148 1732
rect 1142 1727 1143 1731
rect 1147 1727 1148 1731
rect 1142 1726 1148 1727
rect 1326 1731 1332 1732
rect 1326 1727 1327 1731
rect 1331 1727 1332 1731
rect 1326 1726 1332 1727
rect 1510 1731 1516 1732
rect 1510 1727 1511 1731
rect 1515 1727 1516 1731
rect 1510 1726 1516 1727
rect 1588 1724 1590 1758
rect 1639 1753 1643 1754
rect 1703 1758 1707 1759
rect 1703 1753 1707 1754
rect 2007 1758 2011 1759
rect 2146 1755 2147 1759
rect 2151 1755 2152 1759
rect 2146 1754 2152 1755
rect 2258 1759 2264 1760
rect 2258 1755 2259 1759
rect 2263 1755 2264 1759
rect 2258 1754 2264 1755
rect 2402 1759 2408 1760
rect 2402 1755 2403 1759
rect 2407 1755 2408 1759
rect 2402 1754 2408 1755
rect 2562 1759 2568 1760
rect 2562 1755 2563 1759
rect 2567 1755 2568 1759
rect 2562 1754 2568 1755
rect 2598 1759 2604 1760
rect 2598 1755 2599 1759
rect 2603 1755 2604 1759
rect 3106 1759 3112 1760
rect 2598 1754 2604 1755
rect 2906 1755 2912 1756
rect 2007 1753 2011 1754
rect 1662 1751 1668 1752
rect 1662 1747 1663 1751
rect 1667 1747 1668 1751
rect 1662 1746 1668 1747
rect 1664 1724 1666 1746
rect 1704 1732 1706 1753
rect 1758 1751 1764 1752
rect 1758 1747 1759 1751
rect 1763 1747 1764 1751
rect 1758 1746 1764 1747
rect 1702 1731 1708 1732
rect 1702 1727 1703 1731
rect 1707 1727 1708 1731
rect 1702 1726 1708 1727
rect 442 1723 448 1724
rect 442 1719 443 1723
rect 447 1719 448 1723
rect 442 1718 448 1719
rect 570 1723 576 1724
rect 570 1719 571 1723
rect 575 1719 576 1723
rect 570 1718 576 1719
rect 770 1723 776 1724
rect 770 1719 771 1723
rect 775 1719 776 1723
rect 770 1718 776 1719
rect 874 1723 880 1724
rect 874 1719 875 1723
rect 879 1719 880 1723
rect 874 1718 880 1719
rect 918 1723 924 1724
rect 918 1719 919 1723
rect 923 1719 924 1723
rect 918 1718 924 1719
rect 1054 1723 1060 1724
rect 1054 1719 1055 1723
rect 1059 1719 1060 1723
rect 1054 1718 1060 1719
rect 1586 1723 1592 1724
rect 1586 1719 1587 1723
rect 1591 1719 1592 1723
rect 1586 1718 1592 1719
rect 1662 1723 1668 1724
rect 1662 1719 1663 1723
rect 1667 1719 1668 1723
rect 1662 1718 1668 1719
rect 494 1712 500 1713
rect 494 1708 495 1712
rect 499 1708 500 1712
rect 494 1707 500 1708
rect 638 1712 644 1713
rect 638 1708 639 1712
rect 643 1708 644 1712
rect 638 1707 644 1708
rect 798 1712 804 1713
rect 798 1708 799 1712
rect 803 1708 804 1712
rect 798 1707 804 1708
rect 966 1712 972 1713
rect 966 1708 967 1712
rect 971 1708 972 1712
rect 966 1707 972 1708
rect 496 1679 498 1707
rect 640 1679 642 1707
rect 800 1679 802 1707
rect 968 1679 970 1707
rect 495 1678 499 1679
rect 495 1673 499 1674
rect 567 1678 571 1679
rect 567 1673 571 1674
rect 639 1678 643 1679
rect 639 1673 643 1674
rect 743 1678 747 1679
rect 743 1673 747 1674
rect 799 1678 803 1679
rect 799 1673 803 1674
rect 935 1678 939 1679
rect 935 1673 939 1674
rect 967 1678 971 1679
rect 967 1673 971 1674
rect 434 1655 440 1656
rect 434 1651 435 1655
rect 439 1651 440 1655
rect 434 1650 440 1651
rect 568 1649 570 1673
rect 744 1649 746 1673
rect 936 1649 938 1673
rect 134 1648 140 1649
rect 110 1645 116 1646
rect 110 1641 111 1645
rect 115 1641 116 1645
rect 134 1644 135 1648
rect 139 1644 140 1648
rect 134 1643 140 1644
rect 246 1648 252 1649
rect 246 1644 247 1648
rect 251 1644 252 1648
rect 246 1643 252 1644
rect 398 1648 404 1649
rect 398 1644 399 1648
rect 403 1644 404 1648
rect 398 1643 404 1644
rect 566 1648 572 1649
rect 566 1644 567 1648
rect 571 1644 572 1648
rect 566 1643 572 1644
rect 742 1648 748 1649
rect 742 1644 743 1648
rect 747 1644 748 1648
rect 742 1643 748 1644
rect 934 1648 940 1649
rect 934 1644 935 1648
rect 939 1644 940 1648
rect 934 1643 940 1644
rect 110 1640 116 1641
rect 322 1639 328 1640
rect 322 1635 323 1639
rect 327 1635 328 1639
rect 322 1634 328 1635
rect 474 1639 480 1640
rect 474 1635 475 1639
rect 479 1635 480 1639
rect 474 1634 480 1635
rect 642 1639 648 1640
rect 642 1635 643 1639
rect 647 1635 648 1639
rect 642 1634 648 1635
rect 1010 1639 1016 1640
rect 1010 1635 1011 1639
rect 1015 1635 1016 1639
rect 1010 1634 1016 1635
rect 134 1629 140 1630
rect 110 1628 116 1629
rect 110 1624 111 1628
rect 115 1624 116 1628
rect 134 1625 135 1629
rect 139 1625 140 1629
rect 134 1624 140 1625
rect 246 1629 252 1630
rect 246 1625 247 1629
rect 251 1625 252 1629
rect 246 1624 252 1625
rect 110 1623 116 1624
rect 112 1599 114 1623
rect 136 1599 138 1624
rect 210 1607 216 1608
rect 210 1603 211 1607
rect 215 1603 216 1607
rect 210 1602 216 1603
rect 111 1598 115 1599
rect 111 1593 115 1594
rect 135 1598 139 1599
rect 135 1593 139 1594
rect 112 1573 114 1593
rect 110 1572 116 1573
rect 136 1572 138 1593
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 110 1567 116 1568
rect 134 1571 140 1572
rect 134 1567 135 1571
rect 139 1567 140 1571
rect 134 1566 140 1567
rect 212 1564 214 1602
rect 248 1599 250 1624
rect 324 1608 326 1634
rect 398 1629 404 1630
rect 398 1625 399 1629
rect 403 1625 404 1629
rect 398 1624 404 1625
rect 322 1607 328 1608
rect 322 1603 323 1607
rect 327 1603 328 1607
rect 322 1602 328 1603
rect 400 1599 402 1624
rect 476 1608 478 1634
rect 566 1629 572 1630
rect 566 1625 567 1629
rect 571 1625 572 1629
rect 566 1624 572 1625
rect 474 1607 480 1608
rect 474 1603 475 1607
rect 479 1603 480 1607
rect 474 1602 480 1603
rect 568 1599 570 1624
rect 644 1608 646 1634
rect 742 1629 748 1630
rect 742 1625 743 1629
rect 747 1625 748 1629
rect 742 1624 748 1625
rect 934 1629 940 1630
rect 934 1625 935 1629
rect 939 1625 940 1629
rect 934 1624 940 1625
rect 642 1607 648 1608
rect 642 1603 643 1607
rect 647 1603 648 1607
rect 642 1602 648 1603
rect 744 1599 746 1624
rect 936 1599 938 1624
rect 1012 1608 1014 1634
rect 1056 1616 1058 1718
rect 1142 1712 1148 1713
rect 1142 1708 1143 1712
rect 1147 1708 1148 1712
rect 1142 1707 1148 1708
rect 1326 1712 1332 1713
rect 1326 1708 1327 1712
rect 1331 1708 1332 1712
rect 1326 1707 1332 1708
rect 1510 1712 1516 1713
rect 1510 1708 1511 1712
rect 1515 1708 1516 1712
rect 1510 1707 1516 1708
rect 1702 1712 1708 1713
rect 1702 1708 1703 1712
rect 1707 1708 1708 1712
rect 1702 1707 1708 1708
rect 1144 1679 1146 1707
rect 1328 1679 1330 1707
rect 1512 1679 1514 1707
rect 1704 1679 1706 1707
rect 1135 1678 1139 1679
rect 1135 1673 1139 1674
rect 1143 1678 1147 1679
rect 1143 1673 1147 1674
rect 1327 1678 1331 1679
rect 1327 1673 1331 1674
rect 1343 1678 1347 1679
rect 1343 1673 1347 1674
rect 1511 1678 1515 1679
rect 1511 1673 1515 1674
rect 1551 1678 1555 1679
rect 1551 1673 1555 1674
rect 1703 1678 1707 1679
rect 1703 1673 1707 1674
rect 1136 1649 1138 1673
rect 1344 1649 1346 1673
rect 1552 1649 1554 1673
rect 1134 1648 1140 1649
rect 1134 1644 1135 1648
rect 1139 1644 1140 1648
rect 1134 1643 1140 1644
rect 1342 1648 1348 1649
rect 1342 1644 1343 1648
rect 1347 1644 1348 1648
rect 1342 1643 1348 1644
rect 1550 1648 1556 1649
rect 1550 1644 1551 1648
rect 1555 1644 1556 1648
rect 1550 1643 1556 1644
rect 1760 1640 1762 1746
rect 2008 1733 2010 1753
rect 2046 1751 2052 1752
rect 2046 1747 2047 1751
rect 2051 1747 2052 1751
rect 2046 1746 2052 1747
rect 2070 1748 2076 1749
rect 2006 1732 2012 1733
rect 2006 1728 2007 1732
rect 2011 1728 2012 1732
rect 2006 1727 2012 1728
rect 2006 1715 2012 1716
rect 2006 1711 2007 1715
rect 2011 1711 2012 1715
rect 2048 1711 2050 1746
rect 2070 1744 2071 1748
rect 2075 1744 2076 1748
rect 2070 1743 2076 1744
rect 2182 1748 2188 1749
rect 2182 1744 2183 1748
rect 2187 1744 2188 1748
rect 2182 1743 2188 1744
rect 2326 1748 2332 1749
rect 2326 1744 2327 1748
rect 2331 1744 2332 1748
rect 2326 1743 2332 1744
rect 2486 1748 2492 1749
rect 2486 1744 2487 1748
rect 2491 1744 2492 1748
rect 2486 1743 2492 1744
rect 2072 1711 2074 1743
rect 2184 1711 2186 1743
rect 2328 1711 2330 1743
rect 2488 1711 2490 1743
rect 2006 1710 2012 1711
rect 2047 1710 2051 1711
rect 2008 1679 2010 1710
rect 2047 1705 2051 1706
rect 2071 1710 2075 1711
rect 2071 1705 2075 1706
rect 2183 1710 2187 1711
rect 2183 1705 2187 1706
rect 2223 1710 2227 1711
rect 2223 1705 2227 1706
rect 2327 1710 2331 1711
rect 2327 1705 2331 1706
rect 2439 1710 2443 1711
rect 2439 1705 2443 1706
rect 2487 1710 2491 1711
rect 2487 1705 2491 1706
rect 2559 1710 2563 1711
rect 2559 1705 2563 1706
rect 1767 1678 1771 1679
rect 1767 1673 1771 1674
rect 2007 1678 2011 1679
rect 2048 1678 2050 1705
rect 2224 1681 2226 1705
rect 2328 1681 2330 1705
rect 2440 1681 2442 1705
rect 2560 1681 2562 1705
rect 2222 1680 2228 1681
rect 2007 1673 2011 1674
rect 2046 1677 2052 1678
rect 2046 1673 2047 1677
rect 2051 1673 2052 1677
rect 2222 1676 2223 1680
rect 2227 1676 2228 1680
rect 2222 1675 2228 1676
rect 2326 1680 2332 1681
rect 2326 1676 2327 1680
rect 2331 1676 2332 1680
rect 2326 1675 2332 1676
rect 2438 1680 2444 1681
rect 2438 1676 2439 1680
rect 2443 1676 2444 1680
rect 2438 1675 2444 1676
rect 2558 1680 2564 1681
rect 2558 1676 2559 1680
rect 2563 1676 2564 1680
rect 2558 1675 2564 1676
rect 1768 1649 1770 1673
rect 1766 1648 1772 1649
rect 1766 1644 1767 1648
rect 1771 1644 1772 1648
rect 2008 1646 2010 1673
rect 2046 1672 2052 1673
rect 2298 1671 2304 1672
rect 2298 1667 2299 1671
rect 2303 1667 2304 1671
rect 2298 1666 2304 1667
rect 2402 1671 2408 1672
rect 2402 1667 2403 1671
rect 2407 1667 2408 1671
rect 2402 1666 2408 1667
rect 2514 1671 2520 1672
rect 2514 1667 2515 1671
rect 2519 1667 2520 1671
rect 2514 1666 2520 1667
rect 2222 1661 2228 1662
rect 2046 1660 2052 1661
rect 2046 1656 2047 1660
rect 2051 1656 2052 1660
rect 2222 1657 2223 1661
rect 2227 1657 2228 1661
rect 2222 1656 2228 1657
rect 2046 1655 2052 1656
rect 1766 1643 1772 1644
rect 2006 1645 2012 1646
rect 2006 1641 2007 1645
rect 2011 1641 2012 1645
rect 2006 1640 2012 1641
rect 1210 1639 1216 1640
rect 1210 1635 1211 1639
rect 1215 1635 1216 1639
rect 1210 1634 1216 1635
rect 1410 1639 1416 1640
rect 1410 1635 1411 1639
rect 1415 1635 1416 1639
rect 1410 1634 1416 1635
rect 1666 1639 1672 1640
rect 1666 1635 1667 1639
rect 1671 1635 1672 1639
rect 1666 1634 1672 1635
rect 1758 1639 1764 1640
rect 1758 1635 1759 1639
rect 1763 1635 1764 1639
rect 1758 1634 1764 1635
rect 1134 1629 1140 1630
rect 1134 1625 1135 1629
rect 1139 1625 1140 1629
rect 1134 1624 1140 1625
rect 1054 1615 1060 1616
rect 1054 1611 1055 1615
rect 1059 1611 1060 1615
rect 1054 1610 1060 1611
rect 1010 1607 1016 1608
rect 1010 1603 1011 1607
rect 1015 1603 1016 1607
rect 1010 1602 1016 1603
rect 1136 1599 1138 1624
rect 1212 1608 1214 1634
rect 1342 1629 1348 1630
rect 1342 1625 1343 1629
rect 1347 1625 1348 1629
rect 1342 1624 1348 1625
rect 1210 1607 1216 1608
rect 1210 1603 1211 1607
rect 1215 1603 1216 1607
rect 1210 1602 1216 1603
rect 1344 1599 1346 1624
rect 247 1598 251 1599
rect 247 1593 251 1594
rect 255 1598 259 1599
rect 255 1593 259 1594
rect 399 1598 403 1599
rect 399 1593 403 1594
rect 423 1598 427 1599
rect 423 1593 427 1594
rect 567 1598 571 1599
rect 567 1593 571 1594
rect 615 1598 619 1599
rect 615 1593 619 1594
rect 743 1598 747 1599
rect 743 1593 747 1594
rect 831 1598 835 1599
rect 831 1593 835 1594
rect 935 1598 939 1599
rect 935 1593 939 1594
rect 1063 1598 1067 1599
rect 1063 1593 1067 1594
rect 1135 1598 1139 1599
rect 1135 1593 1139 1594
rect 1311 1598 1315 1599
rect 1311 1593 1315 1594
rect 1343 1598 1347 1599
rect 1343 1593 1347 1594
rect 218 1591 224 1592
rect 218 1587 219 1591
rect 223 1587 224 1591
rect 218 1586 224 1587
rect 220 1564 222 1586
rect 256 1572 258 1593
rect 338 1591 344 1592
rect 338 1587 339 1591
rect 343 1587 344 1591
rect 338 1586 344 1587
rect 254 1571 260 1572
rect 254 1567 255 1571
rect 259 1567 260 1571
rect 254 1566 260 1567
rect 340 1564 342 1586
rect 424 1572 426 1593
rect 574 1591 580 1592
rect 574 1587 575 1591
rect 579 1587 580 1591
rect 574 1586 580 1587
rect 422 1571 428 1572
rect 422 1567 423 1571
rect 427 1567 428 1571
rect 422 1566 428 1567
rect 576 1564 578 1586
rect 616 1572 618 1593
rect 832 1572 834 1593
rect 850 1591 856 1592
rect 850 1587 851 1591
rect 855 1587 856 1591
rect 850 1586 856 1587
rect 614 1571 620 1572
rect 614 1567 615 1571
rect 619 1567 620 1571
rect 614 1566 620 1567
rect 830 1571 836 1572
rect 830 1567 831 1571
rect 835 1567 836 1571
rect 830 1566 836 1567
rect 210 1563 216 1564
rect 210 1559 211 1563
rect 215 1559 216 1563
rect 210 1558 216 1559
rect 218 1563 224 1564
rect 218 1559 219 1563
rect 223 1559 224 1563
rect 218 1558 224 1559
rect 338 1563 344 1564
rect 338 1559 339 1563
rect 343 1559 344 1563
rect 338 1558 344 1559
rect 574 1563 580 1564
rect 574 1559 575 1563
rect 579 1559 580 1563
rect 574 1558 580 1559
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 110 1550 116 1551
rect 134 1552 140 1553
rect 112 1519 114 1550
rect 134 1548 135 1552
rect 139 1548 140 1552
rect 134 1547 140 1548
rect 254 1552 260 1553
rect 254 1548 255 1552
rect 259 1548 260 1552
rect 254 1547 260 1548
rect 422 1552 428 1553
rect 422 1548 423 1552
rect 427 1548 428 1552
rect 422 1547 428 1548
rect 614 1552 620 1553
rect 614 1548 615 1552
rect 619 1548 620 1552
rect 614 1547 620 1548
rect 830 1552 836 1553
rect 830 1548 831 1552
rect 835 1548 836 1552
rect 830 1547 836 1548
rect 136 1519 138 1547
rect 256 1519 258 1547
rect 424 1519 426 1547
rect 616 1519 618 1547
rect 832 1519 834 1547
rect 111 1518 115 1519
rect 111 1513 115 1514
rect 135 1518 139 1519
rect 135 1513 139 1514
rect 239 1518 243 1519
rect 239 1513 243 1514
rect 255 1518 259 1519
rect 255 1513 259 1514
rect 407 1518 411 1519
rect 407 1513 411 1514
rect 423 1518 427 1519
rect 423 1513 427 1514
rect 583 1518 587 1519
rect 583 1513 587 1514
rect 615 1518 619 1519
rect 615 1513 619 1514
rect 775 1518 779 1519
rect 775 1513 779 1514
rect 831 1518 835 1519
rect 831 1513 835 1514
rect 112 1486 114 1513
rect 240 1489 242 1513
rect 408 1489 410 1513
rect 584 1489 586 1513
rect 776 1489 778 1513
rect 238 1488 244 1489
rect 110 1485 116 1486
rect 110 1481 111 1485
rect 115 1481 116 1485
rect 238 1484 239 1488
rect 243 1484 244 1488
rect 238 1483 244 1484
rect 406 1488 412 1489
rect 406 1484 407 1488
rect 411 1484 412 1488
rect 406 1483 412 1484
rect 582 1488 588 1489
rect 582 1484 583 1488
rect 587 1484 588 1488
rect 582 1483 588 1484
rect 774 1488 780 1489
rect 774 1484 775 1488
rect 779 1484 780 1488
rect 774 1483 780 1484
rect 110 1480 116 1481
rect 852 1480 854 1586
rect 1064 1572 1066 1593
rect 1146 1591 1152 1592
rect 1146 1587 1147 1591
rect 1151 1587 1152 1591
rect 1146 1586 1152 1587
rect 1062 1571 1068 1572
rect 1062 1567 1063 1571
rect 1067 1567 1068 1571
rect 1062 1566 1068 1567
rect 1148 1564 1150 1586
rect 1312 1572 1314 1593
rect 1412 1592 1414 1634
rect 1550 1629 1556 1630
rect 1550 1625 1551 1629
rect 1555 1625 1556 1629
rect 1550 1624 1556 1625
rect 1552 1599 1554 1624
rect 1668 1608 1670 1634
rect 2048 1631 2050 1655
rect 2224 1631 2226 1656
rect 2300 1640 2302 1666
rect 2326 1661 2332 1662
rect 2326 1657 2327 1661
rect 2331 1657 2332 1661
rect 2326 1656 2332 1657
rect 2298 1639 2304 1640
rect 2298 1635 2299 1639
rect 2303 1635 2304 1639
rect 2298 1634 2304 1635
rect 2328 1631 2330 1656
rect 2404 1640 2406 1666
rect 2438 1661 2444 1662
rect 2438 1657 2439 1661
rect 2443 1657 2444 1661
rect 2438 1656 2444 1657
rect 2402 1639 2408 1640
rect 2402 1635 2403 1639
rect 2407 1635 2408 1639
rect 2402 1634 2408 1635
rect 2440 1631 2442 1656
rect 2516 1640 2518 1666
rect 2558 1661 2564 1662
rect 2558 1657 2559 1661
rect 2563 1657 2564 1661
rect 2558 1656 2564 1657
rect 2514 1639 2520 1640
rect 2514 1635 2515 1639
rect 2519 1635 2520 1639
rect 2514 1634 2520 1635
rect 2560 1631 2562 1656
rect 2600 1648 2602 1754
rect 2906 1751 2907 1755
rect 2911 1751 2912 1755
rect 3106 1755 3107 1759
rect 3111 1755 3112 1759
rect 3106 1754 3112 1755
rect 3306 1759 3312 1760
rect 3306 1755 3307 1759
rect 3311 1755 3312 1759
rect 3306 1754 3312 1755
rect 3722 1759 3728 1760
rect 3722 1755 3723 1759
rect 3727 1755 3728 1759
rect 3722 1754 3728 1755
rect 2906 1750 2912 1751
rect 2654 1748 2660 1749
rect 2654 1744 2655 1748
rect 2659 1744 2660 1748
rect 2654 1743 2660 1744
rect 2830 1748 2836 1749
rect 2830 1744 2831 1748
rect 2835 1744 2836 1748
rect 2830 1743 2836 1744
rect 2656 1711 2658 1743
rect 2832 1711 2834 1743
rect 2655 1710 2659 1711
rect 2655 1705 2659 1706
rect 2687 1710 2691 1711
rect 2687 1705 2691 1706
rect 2823 1710 2827 1711
rect 2823 1705 2827 1706
rect 2831 1710 2835 1711
rect 2831 1705 2835 1706
rect 2688 1681 2690 1705
rect 2824 1681 2826 1705
rect 2686 1680 2692 1681
rect 2686 1676 2687 1680
rect 2691 1676 2692 1680
rect 2686 1675 2692 1676
rect 2822 1680 2828 1681
rect 2822 1676 2823 1680
rect 2827 1676 2828 1680
rect 2822 1675 2828 1676
rect 2634 1671 2640 1672
rect 2634 1667 2635 1671
rect 2639 1667 2640 1671
rect 2634 1666 2640 1667
rect 2658 1671 2664 1672
rect 2658 1667 2659 1671
rect 2663 1667 2664 1671
rect 2658 1666 2664 1667
rect 2598 1647 2604 1648
rect 2598 1643 2599 1647
rect 2603 1643 2604 1647
rect 2598 1642 2604 1643
rect 2636 1640 2638 1666
rect 2634 1639 2640 1640
rect 2634 1635 2635 1639
rect 2639 1635 2640 1639
rect 2634 1634 2640 1635
rect 2660 1632 2662 1666
rect 2686 1661 2692 1662
rect 2686 1657 2687 1661
rect 2691 1657 2692 1661
rect 2686 1656 2692 1657
rect 2822 1661 2828 1662
rect 2822 1657 2823 1661
rect 2827 1657 2828 1661
rect 2822 1656 2828 1657
rect 2658 1631 2664 1632
rect 2688 1631 2690 1656
rect 2824 1631 2826 1656
rect 2908 1640 2910 1750
rect 3022 1748 3028 1749
rect 3022 1744 3023 1748
rect 3027 1744 3028 1748
rect 3022 1743 3028 1744
rect 3222 1748 3228 1749
rect 3222 1744 3223 1748
rect 3227 1744 3228 1748
rect 3222 1743 3228 1744
rect 3430 1748 3436 1749
rect 3430 1744 3431 1748
rect 3435 1744 3436 1748
rect 3430 1743 3436 1744
rect 3646 1748 3652 1749
rect 3646 1744 3647 1748
rect 3651 1744 3652 1748
rect 3646 1743 3652 1744
rect 3024 1711 3026 1743
rect 3224 1711 3226 1743
rect 3432 1711 3434 1743
rect 3648 1711 3650 1743
rect 2967 1710 2971 1711
rect 2967 1705 2971 1706
rect 3023 1710 3027 1711
rect 3023 1705 3027 1706
rect 3127 1710 3131 1711
rect 3127 1705 3131 1706
rect 3223 1710 3227 1711
rect 3223 1705 3227 1706
rect 3303 1710 3307 1711
rect 3303 1705 3307 1706
rect 3431 1710 3435 1711
rect 3431 1705 3435 1706
rect 3487 1710 3491 1711
rect 3487 1705 3491 1706
rect 3647 1710 3651 1711
rect 3647 1705 3651 1706
rect 3671 1710 3675 1711
rect 3671 1705 3675 1706
rect 2968 1681 2970 1705
rect 3128 1681 3130 1705
rect 3304 1681 3306 1705
rect 3488 1681 3490 1705
rect 3672 1681 3674 1705
rect 2966 1680 2972 1681
rect 2966 1676 2967 1680
rect 2971 1676 2972 1680
rect 2966 1675 2972 1676
rect 3126 1680 3132 1681
rect 3126 1676 3127 1680
rect 3131 1676 3132 1680
rect 3126 1675 3132 1676
rect 3302 1680 3308 1681
rect 3302 1676 3303 1680
rect 3307 1676 3308 1680
rect 3302 1675 3308 1676
rect 3486 1680 3492 1681
rect 3486 1676 3487 1680
rect 3491 1676 3492 1680
rect 3486 1675 3492 1676
rect 3670 1680 3676 1681
rect 3670 1676 3671 1680
rect 3675 1676 3676 1680
rect 3670 1675 3676 1676
rect 3740 1672 3742 1782
rect 3840 1768 3842 1789
rect 3908 1788 3910 1830
rect 3916 1804 3918 1906
rect 3942 1903 3943 1907
rect 3947 1903 3948 1907
rect 3942 1902 3948 1903
rect 3944 1875 3946 1902
rect 3943 1874 3947 1875
rect 3943 1869 3947 1870
rect 3944 1842 3946 1869
rect 3942 1841 3948 1842
rect 3942 1837 3943 1841
rect 3947 1837 3948 1841
rect 3942 1836 3948 1837
rect 3942 1824 3948 1825
rect 3942 1820 3943 1824
rect 3947 1820 3948 1824
rect 3942 1819 3948 1820
rect 3914 1803 3920 1804
rect 3914 1799 3915 1803
rect 3919 1799 3920 1803
rect 3914 1798 3920 1799
rect 3944 1795 3946 1819
rect 3943 1794 3947 1795
rect 3943 1789 3947 1790
rect 3906 1787 3912 1788
rect 3906 1783 3907 1787
rect 3911 1783 3912 1787
rect 3906 1782 3912 1783
rect 3944 1769 3946 1789
rect 3942 1768 3948 1769
rect 3838 1767 3844 1768
rect 3838 1763 3839 1767
rect 3843 1763 3844 1767
rect 3942 1764 3943 1768
rect 3947 1764 3948 1768
rect 3942 1763 3948 1764
rect 3838 1762 3844 1763
rect 3906 1751 3912 1752
rect 3838 1748 3844 1749
rect 3838 1744 3839 1748
rect 3843 1744 3844 1748
rect 3906 1747 3907 1751
rect 3911 1747 3912 1751
rect 3906 1746 3912 1747
rect 3942 1751 3948 1752
rect 3942 1747 3943 1751
rect 3947 1747 3948 1751
rect 3942 1746 3948 1747
rect 3838 1743 3844 1744
rect 3840 1711 3842 1743
rect 3839 1710 3843 1711
rect 3839 1705 3843 1706
rect 3840 1681 3842 1705
rect 3838 1680 3844 1681
rect 3838 1676 3839 1680
rect 3843 1676 3844 1680
rect 3838 1675 3844 1676
rect 2946 1671 2952 1672
rect 2946 1667 2947 1671
rect 2951 1667 2952 1671
rect 2946 1666 2952 1667
rect 3042 1671 3048 1672
rect 3042 1667 3043 1671
rect 3047 1667 3048 1671
rect 3042 1666 3048 1667
rect 3202 1671 3208 1672
rect 3202 1667 3203 1671
rect 3207 1667 3208 1671
rect 3202 1666 3208 1667
rect 3378 1671 3384 1672
rect 3378 1667 3379 1671
rect 3383 1667 3384 1671
rect 3378 1666 3384 1667
rect 3438 1671 3444 1672
rect 3438 1667 3439 1671
rect 3443 1667 3444 1671
rect 3438 1666 3444 1667
rect 3738 1671 3744 1672
rect 3738 1667 3739 1671
rect 3743 1667 3744 1671
rect 3738 1666 3744 1667
rect 2948 1640 2950 1666
rect 2966 1661 2972 1662
rect 2966 1657 2967 1661
rect 2971 1657 2972 1661
rect 2966 1656 2972 1657
rect 2906 1639 2912 1640
rect 2906 1635 2907 1639
rect 2911 1635 2912 1639
rect 2906 1634 2912 1635
rect 2946 1639 2952 1640
rect 2946 1635 2947 1639
rect 2951 1635 2952 1639
rect 2946 1634 2952 1635
rect 2968 1631 2970 1656
rect 3044 1640 3046 1666
rect 3126 1661 3132 1662
rect 3126 1657 3127 1661
rect 3131 1657 3132 1661
rect 3126 1656 3132 1657
rect 3042 1639 3048 1640
rect 3042 1635 3043 1639
rect 3047 1635 3048 1639
rect 3042 1634 3048 1635
rect 3128 1631 3130 1656
rect 3204 1640 3206 1666
rect 3302 1661 3308 1662
rect 3302 1657 3303 1661
rect 3307 1657 3308 1661
rect 3302 1656 3308 1657
rect 3202 1639 3208 1640
rect 3202 1635 3203 1639
rect 3207 1635 3208 1639
rect 3202 1634 3208 1635
rect 3304 1631 3306 1656
rect 3380 1640 3382 1666
rect 3378 1639 3384 1640
rect 3378 1635 3379 1639
rect 3383 1635 3384 1639
rect 3378 1634 3384 1635
rect 3440 1632 3442 1666
rect 3486 1661 3492 1662
rect 3486 1657 3487 1661
rect 3491 1657 3492 1661
rect 3486 1656 3492 1657
rect 3670 1661 3676 1662
rect 3670 1657 3671 1661
rect 3675 1657 3676 1661
rect 3670 1656 3676 1657
rect 3838 1661 3844 1662
rect 3838 1657 3839 1661
rect 3843 1657 3844 1661
rect 3838 1656 3844 1657
rect 3438 1631 3444 1632
rect 3488 1631 3490 1656
rect 3672 1631 3674 1656
rect 3794 1639 3800 1640
rect 3794 1635 3795 1639
rect 3799 1635 3800 1639
rect 3794 1634 3800 1635
rect 2047 1630 2051 1631
rect 1766 1629 1772 1630
rect 1766 1625 1767 1629
rect 1771 1625 1772 1629
rect 1766 1624 1772 1625
rect 2006 1628 2012 1629
rect 2006 1624 2007 1628
rect 2011 1624 2012 1628
rect 2047 1625 2051 1626
rect 2223 1630 2227 1631
rect 2223 1625 2227 1626
rect 2327 1630 2331 1631
rect 2327 1625 2331 1626
rect 2391 1630 2395 1631
rect 2391 1625 2395 1626
rect 2439 1630 2443 1631
rect 2439 1625 2443 1626
rect 2503 1630 2507 1631
rect 2503 1625 2507 1626
rect 2559 1630 2563 1631
rect 2559 1625 2563 1626
rect 2615 1630 2619 1631
rect 2658 1627 2659 1631
rect 2663 1627 2664 1631
rect 2658 1626 2664 1627
rect 2687 1630 2691 1631
rect 2615 1625 2619 1626
rect 2687 1625 2691 1626
rect 2735 1630 2739 1631
rect 2735 1625 2739 1626
rect 2823 1630 2827 1631
rect 2823 1625 2827 1626
rect 2855 1630 2859 1631
rect 2855 1625 2859 1626
rect 2967 1630 2971 1631
rect 2967 1625 2971 1626
rect 2975 1630 2979 1631
rect 2975 1625 2979 1626
rect 3095 1630 3099 1631
rect 3095 1625 3099 1626
rect 3127 1630 3131 1631
rect 3127 1625 3131 1626
rect 3215 1630 3219 1631
rect 3215 1625 3219 1626
rect 3303 1630 3307 1631
rect 3303 1625 3307 1626
rect 3335 1630 3339 1631
rect 3438 1627 3439 1631
rect 3443 1627 3444 1631
rect 3438 1626 3444 1627
rect 3455 1630 3459 1631
rect 3335 1625 3339 1626
rect 3455 1625 3459 1626
rect 3487 1630 3491 1631
rect 3487 1625 3491 1626
rect 3671 1630 3675 1631
rect 3671 1625 3675 1626
rect 1642 1607 1648 1608
rect 1642 1603 1643 1607
rect 1647 1603 1648 1607
rect 1642 1602 1648 1603
rect 1666 1607 1672 1608
rect 1666 1603 1667 1607
rect 1671 1603 1672 1607
rect 1666 1602 1672 1603
rect 1551 1598 1555 1599
rect 1551 1593 1555 1594
rect 1567 1598 1571 1599
rect 1567 1593 1571 1594
rect 1410 1591 1416 1592
rect 1410 1587 1411 1591
rect 1415 1587 1416 1591
rect 1410 1586 1416 1587
rect 1568 1572 1570 1593
rect 1310 1571 1316 1572
rect 1310 1567 1311 1571
rect 1315 1567 1316 1571
rect 1310 1566 1316 1567
rect 1566 1571 1572 1572
rect 1566 1567 1567 1571
rect 1571 1567 1572 1571
rect 1566 1566 1572 1567
rect 1644 1564 1646 1602
rect 1768 1599 1770 1624
rect 2006 1623 2012 1624
rect 2008 1599 2010 1623
rect 2048 1605 2050 1625
rect 2046 1604 2052 1605
rect 2392 1604 2394 1625
rect 2466 1623 2472 1624
rect 2466 1619 2467 1623
rect 2471 1619 2472 1623
rect 2466 1618 2472 1619
rect 2046 1600 2047 1604
rect 2051 1600 2052 1604
rect 2046 1599 2052 1600
rect 2390 1603 2396 1604
rect 2390 1599 2391 1603
rect 2395 1599 2396 1603
rect 1767 1598 1771 1599
rect 1767 1593 1771 1594
rect 1831 1598 1835 1599
rect 1831 1593 1835 1594
rect 2007 1598 2011 1599
rect 2390 1598 2396 1599
rect 2468 1596 2470 1618
rect 2504 1604 2506 1625
rect 2578 1623 2584 1624
rect 2578 1619 2579 1623
rect 2583 1619 2584 1623
rect 2578 1618 2584 1619
rect 2502 1603 2508 1604
rect 2502 1599 2503 1603
rect 2507 1599 2508 1603
rect 2502 1598 2508 1599
rect 2580 1596 2582 1618
rect 2616 1604 2618 1625
rect 2726 1623 2732 1624
rect 2726 1619 2727 1623
rect 2731 1619 2732 1623
rect 2726 1618 2732 1619
rect 2614 1603 2620 1604
rect 2614 1599 2615 1603
rect 2619 1599 2620 1603
rect 2614 1598 2620 1599
rect 2728 1596 2730 1618
rect 2736 1604 2738 1625
rect 2810 1623 2816 1624
rect 2810 1619 2811 1623
rect 2815 1619 2816 1623
rect 2810 1618 2816 1619
rect 2734 1603 2740 1604
rect 2734 1599 2735 1603
rect 2739 1599 2740 1603
rect 2734 1598 2740 1599
rect 2812 1596 2814 1618
rect 2856 1604 2858 1625
rect 2976 1604 2978 1625
rect 3050 1623 3056 1624
rect 3050 1619 3051 1623
rect 3055 1619 3056 1623
rect 3050 1618 3056 1619
rect 2854 1603 2860 1604
rect 2854 1599 2855 1603
rect 2859 1599 2860 1603
rect 2854 1598 2860 1599
rect 2974 1603 2980 1604
rect 2974 1599 2975 1603
rect 2979 1599 2980 1603
rect 2974 1598 2980 1599
rect 3052 1596 3054 1618
rect 3096 1604 3098 1625
rect 3170 1623 3176 1624
rect 3170 1619 3171 1623
rect 3175 1619 3176 1623
rect 3170 1618 3176 1619
rect 3094 1603 3100 1604
rect 3094 1599 3095 1603
rect 3099 1599 3100 1603
rect 3094 1598 3100 1599
rect 3172 1596 3174 1618
rect 3216 1604 3218 1625
rect 3290 1623 3296 1624
rect 3290 1619 3291 1623
rect 3295 1619 3296 1623
rect 3290 1618 3296 1619
rect 3214 1603 3220 1604
rect 3214 1599 3215 1603
rect 3219 1599 3220 1603
rect 3214 1598 3220 1599
rect 3292 1596 3294 1618
rect 3336 1604 3338 1625
rect 3410 1623 3416 1624
rect 3410 1619 3411 1623
rect 3415 1619 3416 1623
rect 3410 1618 3416 1619
rect 3334 1603 3340 1604
rect 3334 1599 3335 1603
rect 3339 1599 3340 1603
rect 3334 1598 3340 1599
rect 3412 1596 3414 1618
rect 3456 1604 3458 1625
rect 3454 1603 3460 1604
rect 3454 1599 3455 1603
rect 3459 1599 3460 1603
rect 3454 1598 3460 1599
rect 2007 1593 2011 1594
rect 2466 1595 2472 1596
rect 1650 1591 1656 1592
rect 1650 1587 1651 1591
rect 1655 1587 1656 1591
rect 1650 1586 1656 1587
rect 1810 1591 1816 1592
rect 1810 1587 1811 1591
rect 1815 1587 1816 1591
rect 1810 1586 1816 1587
rect 1652 1564 1654 1586
rect 1034 1563 1040 1564
rect 1034 1559 1035 1563
rect 1039 1559 1040 1563
rect 1034 1558 1040 1559
rect 1146 1563 1152 1564
rect 1146 1559 1147 1563
rect 1151 1559 1152 1563
rect 1146 1558 1152 1559
rect 1642 1563 1648 1564
rect 1642 1559 1643 1563
rect 1647 1559 1648 1563
rect 1642 1558 1648 1559
rect 1650 1563 1656 1564
rect 1650 1559 1651 1563
rect 1655 1559 1656 1563
rect 1650 1558 1656 1559
rect 967 1518 971 1519
rect 967 1513 971 1514
rect 968 1489 970 1513
rect 966 1488 972 1489
rect 966 1484 967 1488
rect 971 1484 972 1488
rect 966 1483 972 1484
rect 482 1479 488 1480
rect 482 1475 483 1479
rect 487 1475 488 1479
rect 482 1474 488 1475
rect 658 1479 664 1480
rect 658 1475 659 1479
rect 663 1475 664 1479
rect 658 1474 664 1475
rect 850 1479 856 1480
rect 850 1475 851 1479
rect 855 1475 856 1479
rect 850 1474 856 1475
rect 238 1469 244 1470
rect 110 1468 116 1469
rect 110 1464 111 1468
rect 115 1464 116 1468
rect 238 1465 239 1469
rect 243 1465 244 1469
rect 238 1464 244 1465
rect 406 1469 412 1470
rect 406 1465 407 1469
rect 411 1465 412 1469
rect 406 1464 412 1465
rect 110 1463 116 1464
rect 112 1435 114 1463
rect 240 1435 242 1464
rect 408 1435 410 1464
rect 484 1448 486 1474
rect 582 1469 588 1470
rect 582 1465 583 1469
rect 587 1465 588 1469
rect 582 1464 588 1465
rect 482 1447 488 1448
rect 482 1443 483 1447
rect 487 1443 488 1447
rect 482 1442 488 1443
rect 584 1435 586 1464
rect 660 1448 662 1474
rect 774 1469 780 1470
rect 774 1465 775 1469
rect 779 1465 780 1469
rect 774 1464 780 1465
rect 966 1469 972 1470
rect 966 1465 967 1469
rect 971 1465 972 1469
rect 966 1464 972 1465
rect 658 1447 664 1448
rect 658 1443 659 1447
rect 663 1443 664 1447
rect 658 1442 664 1443
rect 776 1435 778 1464
rect 968 1435 970 1464
rect 1036 1448 1038 1558
rect 1062 1552 1068 1553
rect 1062 1548 1063 1552
rect 1067 1548 1068 1552
rect 1062 1547 1068 1548
rect 1310 1552 1316 1553
rect 1310 1548 1311 1552
rect 1315 1548 1316 1552
rect 1310 1547 1316 1548
rect 1566 1552 1572 1553
rect 1566 1548 1567 1552
rect 1571 1548 1572 1552
rect 1566 1547 1572 1548
rect 1064 1519 1066 1547
rect 1312 1519 1314 1547
rect 1568 1519 1570 1547
rect 1063 1518 1067 1519
rect 1063 1513 1067 1514
rect 1159 1518 1163 1519
rect 1159 1513 1163 1514
rect 1311 1518 1315 1519
rect 1311 1513 1315 1514
rect 1351 1518 1355 1519
rect 1351 1513 1355 1514
rect 1543 1518 1547 1519
rect 1543 1513 1547 1514
rect 1567 1518 1571 1519
rect 1567 1513 1571 1514
rect 1735 1518 1739 1519
rect 1735 1513 1739 1514
rect 1160 1489 1162 1513
rect 1352 1489 1354 1513
rect 1544 1489 1546 1513
rect 1736 1489 1738 1513
rect 1158 1488 1164 1489
rect 1158 1484 1159 1488
rect 1163 1484 1164 1488
rect 1158 1483 1164 1484
rect 1350 1488 1356 1489
rect 1350 1484 1351 1488
rect 1355 1484 1356 1488
rect 1350 1483 1356 1484
rect 1542 1488 1548 1489
rect 1542 1484 1543 1488
rect 1547 1484 1548 1488
rect 1542 1483 1548 1484
rect 1734 1488 1740 1489
rect 1734 1484 1735 1488
rect 1739 1484 1740 1488
rect 1734 1483 1740 1484
rect 1812 1480 1814 1586
rect 1832 1572 1834 1593
rect 2008 1573 2010 1593
rect 2466 1591 2467 1595
rect 2471 1591 2472 1595
rect 2466 1590 2472 1591
rect 2578 1595 2584 1596
rect 2578 1591 2579 1595
rect 2583 1591 2584 1595
rect 2578 1590 2584 1591
rect 2726 1595 2732 1596
rect 2726 1591 2727 1595
rect 2731 1591 2732 1595
rect 2726 1590 2732 1591
rect 2810 1595 2816 1596
rect 2810 1591 2811 1595
rect 2815 1591 2816 1595
rect 2810 1590 2816 1591
rect 2818 1595 2824 1596
rect 2818 1591 2819 1595
rect 2823 1591 2824 1595
rect 2818 1590 2824 1591
rect 3050 1595 3056 1596
rect 3050 1591 3051 1595
rect 3055 1591 3056 1595
rect 3050 1590 3056 1591
rect 3170 1595 3176 1596
rect 3170 1591 3171 1595
rect 3175 1591 3176 1595
rect 3170 1590 3176 1591
rect 3290 1595 3296 1596
rect 3290 1591 3291 1595
rect 3295 1591 3296 1595
rect 3290 1590 3296 1591
rect 3410 1595 3416 1596
rect 3410 1591 3411 1595
rect 3415 1591 3416 1595
rect 3410 1590 3416 1591
rect 3418 1595 3424 1596
rect 3418 1591 3419 1595
rect 3423 1591 3424 1595
rect 3418 1590 3424 1591
rect 2046 1587 2052 1588
rect 2046 1583 2047 1587
rect 2051 1583 2052 1587
rect 2046 1582 2052 1583
rect 2390 1584 2396 1585
rect 2006 1572 2012 1573
rect 1830 1571 1836 1572
rect 1830 1567 1831 1571
rect 1835 1567 1836 1571
rect 2006 1568 2007 1572
rect 2011 1568 2012 1572
rect 2006 1567 2012 1568
rect 1830 1566 1836 1567
rect 2006 1555 2012 1556
rect 2048 1555 2050 1582
rect 2390 1580 2391 1584
rect 2395 1580 2396 1584
rect 2390 1579 2396 1580
rect 2502 1584 2508 1585
rect 2502 1580 2503 1584
rect 2507 1580 2508 1584
rect 2502 1579 2508 1580
rect 2614 1584 2620 1585
rect 2614 1580 2615 1584
rect 2619 1580 2620 1584
rect 2614 1579 2620 1580
rect 2734 1584 2740 1585
rect 2734 1580 2735 1584
rect 2739 1580 2740 1584
rect 2734 1579 2740 1580
rect 2392 1555 2394 1579
rect 2504 1555 2506 1579
rect 2616 1555 2618 1579
rect 2736 1555 2738 1579
rect 1830 1552 1836 1553
rect 1830 1548 1831 1552
rect 1835 1548 1836 1552
rect 2006 1551 2007 1555
rect 2011 1551 2012 1555
rect 2006 1550 2012 1551
rect 2047 1554 2051 1555
rect 1830 1547 1836 1548
rect 1832 1519 1834 1547
rect 2008 1519 2010 1550
rect 2047 1549 2051 1550
rect 2391 1554 2395 1555
rect 2391 1549 2395 1550
rect 2503 1554 2507 1555
rect 2503 1549 2507 1550
rect 2543 1554 2547 1555
rect 2543 1549 2547 1550
rect 2615 1554 2619 1555
rect 2615 1549 2619 1550
rect 2671 1554 2675 1555
rect 2671 1549 2675 1550
rect 2735 1554 2739 1555
rect 2735 1549 2739 1550
rect 2799 1554 2803 1555
rect 2799 1549 2803 1550
rect 2048 1522 2050 1549
rect 2544 1525 2546 1549
rect 2672 1525 2674 1549
rect 2800 1525 2802 1549
rect 2542 1524 2548 1525
rect 2046 1521 2052 1522
rect 1831 1518 1835 1519
rect 1831 1513 1835 1514
rect 1903 1518 1907 1519
rect 1903 1513 1907 1514
rect 2007 1518 2011 1519
rect 2046 1517 2047 1521
rect 2051 1517 2052 1521
rect 2542 1520 2543 1524
rect 2547 1520 2548 1524
rect 2542 1519 2548 1520
rect 2670 1524 2676 1525
rect 2670 1520 2671 1524
rect 2675 1520 2676 1524
rect 2670 1519 2676 1520
rect 2798 1524 2804 1525
rect 2798 1520 2799 1524
rect 2803 1520 2804 1524
rect 2798 1519 2804 1520
rect 2046 1516 2052 1517
rect 2007 1513 2011 1514
rect 2618 1515 2624 1516
rect 1904 1489 1906 1513
rect 1902 1488 1908 1489
rect 1902 1484 1903 1488
rect 1907 1484 1908 1488
rect 2008 1486 2010 1513
rect 2618 1511 2619 1515
rect 2623 1511 2624 1515
rect 2618 1510 2624 1511
rect 2746 1515 2752 1516
rect 2746 1511 2747 1515
rect 2751 1511 2752 1515
rect 2746 1510 2752 1511
rect 2542 1505 2548 1506
rect 2046 1504 2052 1505
rect 2046 1500 2047 1504
rect 2051 1500 2052 1504
rect 2542 1501 2543 1505
rect 2547 1501 2548 1505
rect 2542 1500 2548 1501
rect 2046 1499 2052 1500
rect 1902 1483 1908 1484
rect 2006 1485 2012 1486
rect 2006 1481 2007 1485
rect 2011 1481 2012 1485
rect 2006 1480 2012 1481
rect 1042 1479 1048 1480
rect 1042 1475 1043 1479
rect 1047 1475 1048 1479
rect 1042 1474 1048 1475
rect 1234 1479 1240 1480
rect 1234 1475 1235 1479
rect 1239 1475 1240 1479
rect 1234 1474 1240 1475
rect 1442 1479 1448 1480
rect 1442 1475 1443 1479
rect 1447 1475 1448 1479
rect 1442 1474 1448 1475
rect 1618 1479 1624 1480
rect 1618 1475 1619 1479
rect 1623 1475 1624 1479
rect 1618 1474 1624 1475
rect 1810 1479 1816 1480
rect 1810 1475 1811 1479
rect 1815 1475 1816 1479
rect 1810 1474 1816 1475
rect 1818 1479 1824 1480
rect 1818 1475 1819 1479
rect 1823 1475 1824 1479
rect 1818 1474 1824 1475
rect 1044 1448 1046 1474
rect 1158 1469 1164 1470
rect 1158 1465 1159 1469
rect 1163 1465 1164 1469
rect 1158 1464 1164 1465
rect 1034 1447 1040 1448
rect 1034 1443 1035 1447
rect 1039 1443 1040 1447
rect 1034 1442 1040 1443
rect 1042 1447 1048 1448
rect 1042 1443 1043 1447
rect 1047 1443 1048 1447
rect 1042 1442 1048 1443
rect 1160 1435 1162 1464
rect 1236 1448 1238 1474
rect 1350 1469 1356 1470
rect 1350 1465 1351 1469
rect 1355 1465 1356 1469
rect 1350 1464 1356 1465
rect 1234 1447 1240 1448
rect 1234 1443 1235 1447
rect 1239 1443 1240 1447
rect 1234 1442 1240 1443
rect 1352 1435 1354 1464
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 239 1434 243 1435
rect 239 1429 243 1430
rect 407 1434 411 1435
rect 407 1429 411 1430
rect 463 1434 467 1435
rect 463 1429 467 1430
rect 583 1434 587 1435
rect 583 1429 587 1430
rect 711 1434 715 1435
rect 711 1429 715 1430
rect 775 1434 779 1435
rect 775 1429 779 1430
rect 855 1434 859 1435
rect 855 1429 859 1430
rect 967 1434 971 1435
rect 967 1429 971 1430
rect 1007 1434 1011 1435
rect 1007 1429 1011 1430
rect 1159 1434 1163 1435
rect 1159 1429 1163 1430
rect 1167 1434 1171 1435
rect 1167 1429 1171 1430
rect 1335 1434 1339 1435
rect 1335 1429 1339 1430
rect 1351 1434 1355 1435
rect 1351 1429 1355 1430
rect 112 1409 114 1429
rect 110 1408 116 1409
rect 464 1408 466 1429
rect 584 1408 586 1429
rect 670 1427 676 1428
rect 670 1423 671 1427
rect 675 1423 676 1427
rect 670 1422 676 1423
rect 110 1404 111 1408
rect 115 1404 116 1408
rect 110 1403 116 1404
rect 462 1407 468 1408
rect 462 1403 463 1407
rect 467 1403 468 1407
rect 462 1402 468 1403
rect 582 1407 588 1408
rect 582 1403 583 1407
rect 587 1403 588 1407
rect 582 1402 588 1403
rect 672 1400 674 1422
rect 712 1408 714 1429
rect 856 1408 858 1429
rect 938 1427 944 1428
rect 938 1423 939 1427
rect 943 1423 944 1427
rect 938 1422 944 1423
rect 710 1407 716 1408
rect 710 1403 711 1407
rect 715 1403 716 1407
rect 710 1402 716 1403
rect 854 1407 860 1408
rect 854 1403 855 1407
rect 859 1403 860 1407
rect 854 1402 860 1403
rect 940 1400 942 1422
rect 1008 1408 1010 1429
rect 1114 1427 1120 1428
rect 1114 1423 1115 1427
rect 1119 1423 1120 1427
rect 1114 1422 1120 1423
rect 1006 1407 1012 1408
rect 1006 1403 1007 1407
rect 1011 1403 1012 1407
rect 1006 1402 1012 1403
rect 670 1399 676 1400
rect 670 1395 671 1399
rect 675 1395 676 1399
rect 670 1394 676 1395
rect 938 1399 944 1400
rect 938 1395 939 1399
rect 943 1395 944 1399
rect 938 1394 944 1395
rect 110 1391 116 1392
rect 110 1387 111 1391
rect 115 1387 116 1391
rect 110 1386 116 1387
rect 462 1388 468 1389
rect 112 1359 114 1386
rect 462 1384 463 1388
rect 467 1384 468 1388
rect 462 1383 468 1384
rect 582 1388 588 1389
rect 582 1384 583 1388
rect 587 1384 588 1388
rect 582 1383 588 1384
rect 710 1388 716 1389
rect 710 1384 711 1388
rect 715 1384 716 1388
rect 710 1383 716 1384
rect 854 1388 860 1389
rect 854 1384 855 1388
rect 859 1384 860 1388
rect 854 1383 860 1384
rect 1006 1388 1012 1389
rect 1006 1384 1007 1388
rect 1011 1384 1012 1388
rect 1006 1383 1012 1384
rect 464 1359 466 1383
rect 584 1359 586 1383
rect 712 1359 714 1383
rect 856 1359 858 1383
rect 1008 1359 1010 1383
rect 111 1358 115 1359
rect 111 1353 115 1354
rect 463 1358 467 1359
rect 463 1353 467 1354
rect 583 1358 587 1359
rect 583 1353 587 1354
rect 655 1358 659 1359
rect 655 1353 659 1354
rect 711 1358 715 1359
rect 711 1353 715 1354
rect 767 1358 771 1359
rect 767 1353 771 1354
rect 855 1358 859 1359
rect 855 1353 859 1354
rect 887 1358 891 1359
rect 887 1353 891 1354
rect 1007 1358 1011 1359
rect 1007 1353 1011 1354
rect 1015 1358 1019 1359
rect 1015 1353 1019 1354
rect 112 1326 114 1353
rect 656 1329 658 1353
rect 768 1329 770 1353
rect 888 1329 890 1353
rect 1016 1329 1018 1353
rect 654 1328 660 1329
rect 110 1325 116 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 654 1324 655 1328
rect 659 1324 660 1328
rect 654 1323 660 1324
rect 766 1328 772 1329
rect 766 1324 767 1328
rect 771 1324 772 1328
rect 766 1323 772 1324
rect 886 1328 892 1329
rect 886 1324 887 1328
rect 891 1324 892 1328
rect 886 1323 892 1324
rect 1014 1328 1020 1329
rect 1014 1324 1015 1328
rect 1019 1324 1020 1328
rect 1014 1323 1020 1324
rect 110 1320 116 1321
rect 1116 1320 1118 1422
rect 1168 1408 1170 1429
rect 1250 1427 1256 1428
rect 1250 1423 1251 1427
rect 1255 1423 1256 1427
rect 1250 1422 1256 1423
rect 1166 1407 1172 1408
rect 1166 1403 1167 1407
rect 1171 1403 1172 1407
rect 1166 1402 1172 1403
rect 1252 1400 1254 1422
rect 1336 1408 1338 1429
rect 1444 1428 1446 1474
rect 1542 1469 1548 1470
rect 1542 1465 1543 1469
rect 1547 1465 1548 1469
rect 1542 1464 1548 1465
rect 1544 1435 1546 1464
rect 1620 1448 1622 1474
rect 1734 1469 1740 1470
rect 1734 1465 1735 1469
rect 1739 1465 1740 1469
rect 1734 1464 1740 1465
rect 1618 1447 1624 1448
rect 1618 1443 1619 1447
rect 1623 1443 1624 1447
rect 1618 1442 1624 1443
rect 1736 1435 1738 1464
rect 1820 1456 1822 1474
rect 1902 1469 1908 1470
rect 1902 1465 1903 1469
rect 1907 1465 1908 1469
rect 1902 1464 1908 1465
rect 2006 1468 2012 1469
rect 2006 1464 2007 1468
rect 2011 1464 2012 1468
rect 2048 1467 2050 1499
rect 2544 1467 2546 1500
rect 2620 1484 2622 1510
rect 2670 1505 2676 1506
rect 2670 1501 2671 1505
rect 2675 1501 2676 1505
rect 2670 1500 2676 1501
rect 2618 1483 2624 1484
rect 2618 1479 2619 1483
rect 2623 1479 2624 1483
rect 2618 1478 2624 1479
rect 2672 1467 2674 1500
rect 2748 1484 2750 1510
rect 2798 1505 2804 1506
rect 2798 1501 2799 1505
rect 2803 1501 2804 1505
rect 2798 1500 2804 1501
rect 2746 1483 2752 1484
rect 2746 1479 2747 1483
rect 2751 1479 2752 1483
rect 2746 1478 2752 1479
rect 2800 1467 2802 1500
rect 2820 1492 2822 1590
rect 2854 1584 2860 1585
rect 2854 1580 2855 1584
rect 2859 1580 2860 1584
rect 2854 1579 2860 1580
rect 2974 1584 2980 1585
rect 2974 1580 2975 1584
rect 2979 1580 2980 1584
rect 2974 1579 2980 1580
rect 3094 1584 3100 1585
rect 3094 1580 3095 1584
rect 3099 1580 3100 1584
rect 3094 1579 3100 1580
rect 3214 1584 3220 1585
rect 3214 1580 3215 1584
rect 3219 1580 3220 1584
rect 3214 1579 3220 1580
rect 3334 1584 3340 1585
rect 3334 1580 3335 1584
rect 3339 1580 3340 1584
rect 3334 1579 3340 1580
rect 2856 1555 2858 1579
rect 2976 1555 2978 1579
rect 3096 1555 3098 1579
rect 3216 1555 3218 1579
rect 3336 1555 3338 1579
rect 2855 1554 2859 1555
rect 2855 1549 2859 1550
rect 2935 1554 2939 1555
rect 2935 1549 2939 1550
rect 2975 1554 2979 1555
rect 2975 1549 2979 1550
rect 3071 1554 3075 1555
rect 3071 1549 3075 1550
rect 3095 1554 3099 1555
rect 3095 1549 3099 1550
rect 3207 1554 3211 1555
rect 3207 1549 3211 1550
rect 3215 1554 3219 1555
rect 3215 1549 3219 1550
rect 3335 1554 3339 1555
rect 3335 1549 3339 1550
rect 2936 1525 2938 1549
rect 3072 1525 3074 1549
rect 3208 1525 3210 1549
rect 3336 1525 3338 1549
rect 2934 1524 2940 1525
rect 2934 1520 2935 1524
rect 2939 1520 2940 1524
rect 2934 1519 2940 1520
rect 3070 1524 3076 1525
rect 3070 1520 3071 1524
rect 3075 1520 3076 1524
rect 3070 1519 3076 1520
rect 3206 1524 3212 1525
rect 3206 1520 3207 1524
rect 3211 1520 3212 1524
rect 3206 1519 3212 1520
rect 3334 1524 3340 1525
rect 3334 1520 3335 1524
rect 3339 1520 3340 1524
rect 3334 1519 3340 1520
rect 2874 1515 2880 1516
rect 2874 1511 2875 1515
rect 2879 1511 2880 1515
rect 2874 1510 2880 1511
rect 3010 1515 3016 1516
rect 3010 1511 3011 1515
rect 3015 1511 3016 1515
rect 3010 1510 3016 1511
rect 3146 1515 3152 1516
rect 3146 1511 3147 1515
rect 3151 1511 3152 1515
rect 3146 1510 3152 1511
rect 3282 1515 3288 1516
rect 3282 1511 3283 1515
rect 3287 1511 3288 1515
rect 3282 1510 3288 1511
rect 3410 1515 3416 1516
rect 3410 1511 3411 1515
rect 3415 1511 3416 1515
rect 3410 1510 3416 1511
rect 2818 1491 2824 1492
rect 2818 1487 2819 1491
rect 2823 1487 2824 1491
rect 2818 1486 2824 1487
rect 2876 1484 2878 1510
rect 2934 1505 2940 1506
rect 2934 1501 2935 1505
rect 2939 1501 2940 1505
rect 2934 1500 2940 1501
rect 2874 1483 2880 1484
rect 2874 1479 2875 1483
rect 2879 1479 2880 1483
rect 2874 1478 2880 1479
rect 2936 1467 2938 1500
rect 3012 1484 3014 1510
rect 3070 1505 3076 1506
rect 3070 1501 3071 1505
rect 3075 1501 3076 1505
rect 3070 1500 3076 1501
rect 3010 1483 3016 1484
rect 3010 1479 3011 1483
rect 3015 1479 3016 1483
rect 3010 1478 3016 1479
rect 3072 1467 3074 1500
rect 1818 1455 1824 1456
rect 1818 1451 1819 1455
rect 1823 1451 1824 1455
rect 1818 1450 1824 1451
rect 1904 1435 1906 1464
rect 2006 1463 2012 1464
rect 2047 1466 2051 1467
rect 1946 1447 1952 1448
rect 1946 1443 1947 1447
rect 1951 1443 1952 1447
rect 1946 1442 1952 1443
rect 1511 1434 1515 1435
rect 1511 1429 1515 1430
rect 1543 1434 1547 1435
rect 1543 1429 1547 1430
rect 1687 1434 1691 1435
rect 1687 1429 1691 1430
rect 1735 1434 1739 1435
rect 1735 1429 1739 1430
rect 1871 1434 1875 1435
rect 1871 1429 1875 1430
rect 1903 1434 1907 1435
rect 1903 1429 1907 1430
rect 1442 1427 1448 1428
rect 1442 1423 1443 1427
rect 1447 1423 1448 1427
rect 1442 1422 1448 1423
rect 1512 1408 1514 1429
rect 1688 1408 1690 1429
rect 1822 1427 1828 1428
rect 1822 1423 1823 1427
rect 1827 1423 1828 1427
rect 1822 1422 1828 1423
rect 1830 1427 1836 1428
rect 1830 1423 1831 1427
rect 1835 1423 1836 1427
rect 1830 1422 1836 1423
rect 1334 1407 1340 1408
rect 1334 1403 1335 1407
rect 1339 1403 1340 1407
rect 1334 1402 1340 1403
rect 1510 1407 1516 1408
rect 1510 1403 1511 1407
rect 1515 1403 1516 1407
rect 1510 1402 1516 1403
rect 1686 1407 1692 1408
rect 1686 1403 1687 1407
rect 1691 1403 1692 1407
rect 1686 1402 1692 1403
rect 1250 1399 1256 1400
rect 1242 1395 1248 1396
rect 1242 1391 1243 1395
rect 1247 1391 1248 1395
rect 1250 1395 1251 1399
rect 1255 1395 1256 1399
rect 1250 1394 1256 1395
rect 1242 1390 1248 1391
rect 1166 1388 1172 1389
rect 1166 1384 1167 1388
rect 1171 1384 1172 1388
rect 1166 1383 1172 1384
rect 1168 1359 1170 1383
rect 1143 1358 1147 1359
rect 1143 1353 1147 1354
rect 1167 1358 1171 1359
rect 1167 1353 1171 1354
rect 1144 1329 1146 1353
rect 1142 1328 1148 1329
rect 1142 1324 1143 1328
rect 1147 1324 1148 1328
rect 1142 1323 1148 1324
rect 730 1319 736 1320
rect 730 1315 731 1319
rect 735 1315 736 1319
rect 730 1314 736 1315
rect 842 1319 848 1320
rect 842 1315 843 1319
rect 847 1315 848 1319
rect 842 1314 848 1315
rect 962 1319 968 1320
rect 962 1315 963 1319
rect 967 1315 968 1319
rect 962 1314 968 1315
rect 1090 1319 1096 1320
rect 1090 1315 1091 1319
rect 1095 1315 1096 1319
rect 1090 1314 1096 1315
rect 1114 1319 1120 1320
rect 1114 1315 1115 1319
rect 1119 1315 1120 1319
rect 1114 1314 1120 1315
rect 654 1309 660 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 654 1305 655 1309
rect 659 1305 660 1309
rect 654 1304 660 1305
rect 110 1303 116 1304
rect 112 1279 114 1303
rect 656 1279 658 1304
rect 732 1288 734 1314
rect 766 1309 772 1310
rect 766 1305 767 1309
rect 771 1305 772 1309
rect 766 1304 772 1305
rect 730 1287 736 1288
rect 730 1283 731 1287
rect 735 1283 736 1287
rect 730 1282 736 1283
rect 768 1279 770 1304
rect 844 1288 846 1314
rect 886 1309 892 1310
rect 886 1305 887 1309
rect 891 1305 892 1309
rect 886 1304 892 1305
rect 842 1287 848 1288
rect 842 1283 843 1287
rect 847 1283 848 1287
rect 842 1282 848 1283
rect 888 1279 890 1304
rect 964 1288 966 1314
rect 1014 1309 1020 1310
rect 1014 1305 1015 1309
rect 1019 1305 1020 1309
rect 1014 1304 1020 1305
rect 962 1287 968 1288
rect 962 1283 963 1287
rect 967 1283 968 1287
rect 962 1282 968 1283
rect 1016 1279 1018 1304
rect 1092 1288 1094 1314
rect 1142 1309 1148 1310
rect 1142 1305 1143 1309
rect 1147 1305 1148 1309
rect 1142 1304 1148 1305
rect 1090 1287 1096 1288
rect 1090 1283 1091 1287
rect 1095 1283 1096 1287
rect 1090 1282 1096 1283
rect 1144 1279 1146 1304
rect 1244 1288 1246 1390
rect 1334 1388 1340 1389
rect 1334 1384 1335 1388
rect 1339 1384 1340 1388
rect 1334 1383 1340 1384
rect 1510 1388 1516 1389
rect 1510 1384 1511 1388
rect 1515 1384 1516 1388
rect 1510 1383 1516 1384
rect 1686 1388 1692 1389
rect 1686 1384 1687 1388
rect 1691 1384 1692 1388
rect 1686 1383 1692 1384
rect 1336 1359 1338 1383
rect 1512 1359 1514 1383
rect 1688 1359 1690 1383
rect 1279 1358 1283 1359
rect 1279 1353 1283 1354
rect 1335 1358 1339 1359
rect 1335 1353 1339 1354
rect 1415 1358 1419 1359
rect 1415 1353 1419 1354
rect 1511 1358 1515 1359
rect 1511 1353 1515 1354
rect 1559 1358 1563 1359
rect 1559 1353 1563 1354
rect 1687 1358 1691 1359
rect 1687 1353 1691 1354
rect 1703 1358 1707 1359
rect 1703 1353 1707 1354
rect 1280 1329 1282 1353
rect 1416 1329 1418 1353
rect 1560 1329 1562 1353
rect 1704 1329 1706 1353
rect 1278 1328 1284 1329
rect 1278 1324 1279 1328
rect 1283 1324 1284 1328
rect 1278 1323 1284 1324
rect 1414 1328 1420 1329
rect 1414 1324 1415 1328
rect 1419 1324 1420 1328
rect 1414 1323 1420 1324
rect 1558 1328 1564 1329
rect 1558 1324 1559 1328
rect 1563 1324 1564 1328
rect 1558 1323 1564 1324
rect 1702 1328 1708 1329
rect 1702 1324 1703 1328
rect 1707 1324 1708 1328
rect 1702 1323 1708 1324
rect 1824 1320 1826 1422
rect 1832 1400 1834 1422
rect 1872 1408 1874 1429
rect 1870 1407 1876 1408
rect 1870 1403 1871 1407
rect 1875 1403 1876 1407
rect 1870 1402 1876 1403
rect 1948 1400 1950 1442
rect 2008 1435 2010 1463
rect 2047 1461 2051 1462
rect 2519 1466 2523 1467
rect 2519 1461 2523 1462
rect 2543 1466 2547 1467
rect 2543 1461 2547 1462
rect 2631 1466 2635 1467
rect 2631 1461 2635 1462
rect 2671 1466 2675 1467
rect 2671 1461 2675 1462
rect 2759 1466 2763 1467
rect 2759 1461 2763 1462
rect 2799 1466 2803 1467
rect 2799 1461 2803 1462
rect 2895 1466 2899 1467
rect 2895 1461 2899 1462
rect 2935 1466 2939 1467
rect 2935 1461 2939 1462
rect 3031 1466 3035 1467
rect 3031 1461 3035 1462
rect 3071 1466 3075 1467
rect 3071 1461 3075 1462
rect 2048 1441 2050 1461
rect 2046 1440 2052 1441
rect 2520 1440 2522 1461
rect 2594 1459 2600 1460
rect 2594 1455 2595 1459
rect 2599 1455 2600 1459
rect 2594 1454 2600 1455
rect 2046 1436 2047 1440
rect 2051 1436 2052 1440
rect 2046 1435 2052 1436
rect 2518 1439 2524 1440
rect 2518 1435 2519 1439
rect 2523 1435 2524 1439
rect 2007 1434 2011 1435
rect 2518 1434 2524 1435
rect 2596 1432 2598 1454
rect 2632 1440 2634 1461
rect 2714 1451 2720 1452
rect 2714 1447 2715 1451
rect 2719 1447 2720 1451
rect 2714 1446 2720 1447
rect 2630 1439 2636 1440
rect 2630 1435 2631 1439
rect 2635 1435 2636 1439
rect 2630 1434 2636 1435
rect 2716 1432 2718 1446
rect 2760 1440 2762 1461
rect 2886 1459 2892 1460
rect 2886 1455 2887 1459
rect 2891 1455 2892 1459
rect 2886 1454 2892 1455
rect 2758 1439 2764 1440
rect 2758 1435 2759 1439
rect 2763 1435 2764 1439
rect 2758 1434 2764 1435
rect 2888 1432 2890 1454
rect 2896 1440 2898 1461
rect 2978 1459 2984 1460
rect 2978 1455 2979 1459
rect 2983 1455 2984 1459
rect 2978 1454 2984 1455
rect 2894 1439 2900 1440
rect 2894 1435 2895 1439
rect 2899 1435 2900 1439
rect 2894 1434 2900 1435
rect 2980 1432 2982 1454
rect 3032 1440 3034 1461
rect 3148 1460 3150 1510
rect 3206 1505 3212 1506
rect 3206 1501 3207 1505
rect 3211 1501 3212 1505
rect 3206 1500 3212 1501
rect 3208 1467 3210 1500
rect 3284 1484 3286 1510
rect 3334 1505 3340 1506
rect 3334 1501 3335 1505
rect 3339 1501 3340 1505
rect 3334 1500 3340 1501
rect 3282 1483 3288 1484
rect 3282 1479 3283 1483
rect 3287 1479 3288 1483
rect 3282 1478 3288 1479
rect 3336 1467 3338 1500
rect 3412 1484 3414 1510
rect 3420 1492 3422 1590
rect 3454 1584 3460 1585
rect 3454 1580 3455 1584
rect 3459 1580 3460 1584
rect 3454 1579 3460 1580
rect 3456 1555 3458 1579
rect 3455 1554 3459 1555
rect 3455 1549 3459 1550
rect 3463 1554 3467 1555
rect 3463 1549 3467 1550
rect 3591 1554 3595 1555
rect 3591 1549 3595 1550
rect 3727 1554 3731 1555
rect 3727 1549 3731 1550
rect 3464 1525 3466 1549
rect 3592 1525 3594 1549
rect 3728 1525 3730 1549
rect 3462 1524 3468 1525
rect 3462 1520 3463 1524
rect 3467 1520 3468 1524
rect 3462 1519 3468 1520
rect 3590 1524 3596 1525
rect 3590 1520 3591 1524
rect 3595 1520 3596 1524
rect 3590 1519 3596 1520
rect 3726 1524 3732 1525
rect 3726 1520 3727 1524
rect 3731 1520 3732 1524
rect 3726 1519 3732 1520
rect 3796 1516 3798 1634
rect 3840 1631 3842 1656
rect 3908 1640 3910 1746
rect 3944 1711 3946 1746
rect 3943 1710 3947 1711
rect 3943 1705 3947 1706
rect 3944 1678 3946 1705
rect 3942 1677 3948 1678
rect 3942 1673 3943 1677
rect 3947 1673 3948 1677
rect 3942 1672 3948 1673
rect 3914 1671 3920 1672
rect 3914 1667 3915 1671
rect 3919 1667 3920 1671
rect 3914 1666 3920 1667
rect 3906 1639 3912 1640
rect 3906 1635 3907 1639
rect 3911 1635 3912 1639
rect 3906 1634 3912 1635
rect 3839 1630 3843 1631
rect 3839 1625 3843 1626
rect 3839 1554 3843 1555
rect 3839 1549 3843 1550
rect 3840 1525 3842 1549
rect 3838 1524 3844 1525
rect 3838 1520 3839 1524
rect 3843 1520 3844 1524
rect 3838 1519 3844 1520
rect 3538 1515 3544 1516
rect 3538 1511 3539 1515
rect 3543 1511 3544 1515
rect 3538 1510 3544 1511
rect 3794 1515 3800 1516
rect 3794 1511 3795 1515
rect 3799 1511 3800 1515
rect 3794 1510 3800 1511
rect 3906 1515 3912 1516
rect 3906 1511 3907 1515
rect 3911 1511 3912 1515
rect 3906 1510 3912 1511
rect 3462 1505 3468 1506
rect 3462 1501 3463 1505
rect 3467 1501 3468 1505
rect 3462 1500 3468 1501
rect 3418 1491 3424 1492
rect 3418 1487 3419 1491
rect 3423 1487 3424 1491
rect 3418 1486 3424 1487
rect 3410 1483 3416 1484
rect 3410 1479 3411 1483
rect 3415 1479 3416 1483
rect 3410 1478 3416 1479
rect 3464 1467 3466 1500
rect 3540 1484 3542 1510
rect 3590 1505 3596 1506
rect 3590 1501 3591 1505
rect 3595 1501 3596 1505
rect 3590 1500 3596 1501
rect 3726 1505 3732 1506
rect 3726 1501 3727 1505
rect 3731 1501 3732 1505
rect 3726 1500 3732 1501
rect 3838 1505 3844 1506
rect 3838 1501 3839 1505
rect 3843 1501 3844 1505
rect 3838 1500 3844 1501
rect 3538 1483 3544 1484
rect 3538 1479 3539 1483
rect 3543 1479 3544 1483
rect 3538 1478 3544 1479
rect 3592 1467 3594 1500
rect 3728 1467 3730 1500
rect 3790 1483 3796 1484
rect 3790 1479 3791 1483
rect 3795 1479 3796 1483
rect 3790 1478 3796 1479
rect 3792 1475 3794 1478
rect 3792 1473 3802 1475
rect 3175 1466 3179 1467
rect 3175 1461 3179 1462
rect 3207 1466 3211 1467
rect 3207 1461 3211 1462
rect 3311 1466 3315 1467
rect 3311 1461 3315 1462
rect 3335 1466 3339 1467
rect 3335 1461 3339 1462
rect 3447 1466 3451 1467
rect 3447 1461 3451 1462
rect 3463 1466 3467 1467
rect 3463 1461 3467 1462
rect 3583 1466 3587 1467
rect 3583 1461 3587 1462
rect 3591 1466 3595 1467
rect 3591 1461 3595 1462
rect 3719 1466 3723 1467
rect 3719 1461 3723 1462
rect 3727 1466 3731 1467
rect 3727 1461 3731 1462
rect 3146 1459 3152 1460
rect 3146 1455 3147 1459
rect 3151 1455 3152 1459
rect 3146 1454 3152 1455
rect 3176 1440 3178 1461
rect 3312 1440 3314 1461
rect 3386 1459 3392 1460
rect 3386 1455 3387 1459
rect 3391 1455 3392 1459
rect 3386 1454 3392 1455
rect 3030 1439 3036 1440
rect 3030 1435 3031 1439
rect 3035 1435 3036 1439
rect 3030 1434 3036 1435
rect 3174 1439 3180 1440
rect 3174 1435 3175 1439
rect 3179 1435 3180 1439
rect 3174 1434 3180 1435
rect 3310 1439 3316 1440
rect 3310 1435 3311 1439
rect 3315 1435 3316 1439
rect 3310 1434 3316 1435
rect 3388 1432 3390 1454
rect 3448 1440 3450 1461
rect 3530 1451 3536 1452
rect 3530 1447 3531 1451
rect 3535 1447 3536 1451
rect 3530 1446 3536 1447
rect 3446 1439 3452 1440
rect 3446 1435 3447 1439
rect 3451 1435 3452 1439
rect 3446 1434 3452 1435
rect 3532 1432 3534 1446
rect 3584 1440 3586 1461
rect 3666 1459 3672 1460
rect 3666 1455 3667 1459
rect 3671 1455 3672 1459
rect 3666 1454 3672 1455
rect 3582 1439 3588 1440
rect 3582 1435 3583 1439
rect 3587 1435 3588 1439
rect 3582 1434 3588 1435
rect 3668 1432 3670 1454
rect 3720 1440 3722 1461
rect 3718 1439 3724 1440
rect 3718 1435 3719 1439
rect 3723 1435 3724 1439
rect 3718 1434 3724 1435
rect 2007 1429 2011 1430
rect 2594 1431 2600 1432
rect 2008 1409 2010 1429
rect 2594 1427 2595 1431
rect 2599 1427 2600 1431
rect 2714 1431 2720 1432
rect 2594 1426 2600 1427
rect 2706 1427 2712 1428
rect 2046 1423 2052 1424
rect 2046 1419 2047 1423
rect 2051 1419 2052 1423
rect 2706 1423 2707 1427
rect 2711 1423 2712 1427
rect 2714 1427 2715 1431
rect 2719 1427 2720 1431
rect 2714 1426 2720 1427
rect 2886 1431 2892 1432
rect 2886 1427 2887 1431
rect 2891 1427 2892 1431
rect 2886 1426 2892 1427
rect 2978 1431 2984 1432
rect 2978 1427 2979 1431
rect 2983 1427 2984 1431
rect 2978 1426 2984 1427
rect 3386 1431 3392 1432
rect 3386 1427 3387 1431
rect 3391 1427 3392 1431
rect 3386 1426 3392 1427
rect 3530 1431 3536 1432
rect 3530 1427 3531 1431
rect 3535 1427 3536 1431
rect 3530 1426 3536 1427
rect 3666 1431 3672 1432
rect 3666 1427 3667 1431
rect 3671 1427 3672 1431
rect 3666 1426 3672 1427
rect 2706 1422 2712 1423
rect 3574 1423 3580 1424
rect 2046 1418 2052 1419
rect 2518 1420 2524 1421
rect 2006 1408 2012 1409
rect 2006 1404 2007 1408
rect 2011 1404 2012 1408
rect 2006 1403 2012 1404
rect 1830 1399 1836 1400
rect 1830 1395 1831 1399
rect 1835 1395 1836 1399
rect 1830 1394 1836 1395
rect 1946 1399 1952 1400
rect 1946 1395 1947 1399
rect 1951 1395 1952 1399
rect 1946 1394 1952 1395
rect 2006 1391 2012 1392
rect 2048 1391 2050 1418
rect 2518 1416 2519 1420
rect 2523 1416 2524 1420
rect 2518 1415 2524 1416
rect 2630 1420 2636 1421
rect 2630 1416 2631 1420
rect 2635 1416 2636 1420
rect 2630 1415 2636 1416
rect 2520 1391 2522 1415
rect 2632 1391 2634 1415
rect 1870 1388 1876 1389
rect 1870 1384 1871 1388
rect 1875 1384 1876 1388
rect 2006 1387 2007 1391
rect 2011 1387 2012 1391
rect 2006 1386 2012 1387
rect 2047 1390 2051 1391
rect 1870 1383 1876 1384
rect 1872 1359 1874 1383
rect 2008 1359 2010 1386
rect 2047 1385 2051 1386
rect 2399 1390 2403 1391
rect 2399 1385 2403 1386
rect 2519 1390 2523 1391
rect 2519 1385 2523 1386
rect 2535 1390 2539 1391
rect 2535 1385 2539 1386
rect 2631 1390 2635 1391
rect 2631 1385 2635 1386
rect 2679 1390 2683 1391
rect 2679 1385 2683 1386
rect 1847 1358 1851 1359
rect 1847 1353 1851 1354
rect 1871 1358 1875 1359
rect 1871 1353 1875 1354
rect 2007 1358 2011 1359
rect 2048 1358 2050 1385
rect 2400 1361 2402 1385
rect 2536 1361 2538 1385
rect 2680 1361 2682 1385
rect 2398 1360 2404 1361
rect 2007 1353 2011 1354
rect 2046 1357 2052 1358
rect 2046 1353 2047 1357
rect 2051 1353 2052 1357
rect 2398 1356 2399 1360
rect 2403 1356 2404 1360
rect 2398 1355 2404 1356
rect 2534 1360 2540 1361
rect 2534 1356 2535 1360
rect 2539 1356 2540 1360
rect 2534 1355 2540 1356
rect 2678 1360 2684 1361
rect 2678 1356 2679 1360
rect 2683 1356 2684 1360
rect 2678 1355 2684 1356
rect 1848 1329 1850 1353
rect 1846 1328 1852 1329
rect 1846 1324 1847 1328
rect 1851 1324 1852 1328
rect 2008 1326 2010 1353
rect 2046 1352 2052 1353
rect 2474 1351 2480 1352
rect 2474 1347 2475 1351
rect 2479 1347 2480 1351
rect 2474 1346 2480 1347
rect 2482 1351 2488 1352
rect 2482 1347 2483 1351
rect 2487 1347 2488 1351
rect 2482 1346 2488 1347
rect 2398 1341 2404 1342
rect 2046 1340 2052 1341
rect 2046 1336 2047 1340
rect 2051 1336 2052 1340
rect 2398 1337 2399 1341
rect 2403 1337 2404 1341
rect 2398 1336 2404 1337
rect 2046 1335 2052 1336
rect 1846 1323 1852 1324
rect 2006 1325 2012 1326
rect 2006 1321 2007 1325
rect 2011 1321 2012 1325
rect 2006 1320 2012 1321
rect 1354 1319 1360 1320
rect 1354 1315 1355 1319
rect 1359 1315 1360 1319
rect 1354 1314 1360 1315
rect 1482 1319 1488 1320
rect 1482 1315 1483 1319
rect 1487 1315 1488 1319
rect 1482 1314 1488 1315
rect 1634 1319 1640 1320
rect 1634 1315 1635 1319
rect 1639 1315 1640 1319
rect 1634 1314 1640 1315
rect 1778 1319 1784 1320
rect 1778 1315 1779 1319
rect 1783 1315 1784 1319
rect 1778 1314 1784 1315
rect 1822 1319 1828 1320
rect 1822 1315 1823 1319
rect 1827 1315 1828 1319
rect 1822 1314 1828 1315
rect 1278 1309 1284 1310
rect 1278 1305 1279 1309
rect 1283 1305 1284 1309
rect 1278 1304 1284 1305
rect 1242 1287 1248 1288
rect 1242 1283 1243 1287
rect 1247 1283 1248 1287
rect 1242 1282 1248 1283
rect 1280 1279 1282 1304
rect 1356 1288 1358 1314
rect 1414 1309 1420 1310
rect 1414 1305 1415 1309
rect 1419 1305 1420 1309
rect 1414 1304 1420 1305
rect 1354 1287 1360 1288
rect 1354 1283 1355 1287
rect 1359 1283 1360 1287
rect 1354 1282 1360 1283
rect 1416 1279 1418 1304
rect 111 1278 115 1279
rect 111 1273 115 1274
rect 439 1278 443 1279
rect 439 1273 443 1274
rect 551 1278 555 1279
rect 551 1273 555 1274
rect 655 1278 659 1279
rect 655 1273 659 1274
rect 671 1278 675 1279
rect 671 1273 675 1274
rect 767 1278 771 1279
rect 767 1273 771 1274
rect 799 1278 803 1279
rect 799 1273 803 1274
rect 887 1278 891 1279
rect 887 1273 891 1274
rect 935 1278 939 1279
rect 935 1273 939 1274
rect 1015 1278 1019 1279
rect 1015 1273 1019 1274
rect 1079 1278 1083 1279
rect 1079 1273 1083 1274
rect 1143 1278 1147 1279
rect 1143 1273 1147 1274
rect 1231 1278 1235 1279
rect 1231 1273 1235 1274
rect 1279 1278 1283 1279
rect 1279 1273 1283 1274
rect 1391 1278 1395 1279
rect 1391 1273 1395 1274
rect 1415 1278 1419 1279
rect 1415 1273 1419 1274
rect 112 1253 114 1273
rect 110 1252 116 1253
rect 440 1252 442 1273
rect 514 1271 520 1272
rect 514 1267 515 1271
rect 519 1267 520 1271
rect 514 1266 520 1267
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 438 1251 444 1252
rect 438 1247 439 1251
rect 443 1247 444 1251
rect 438 1246 444 1247
rect 516 1244 518 1266
rect 552 1252 554 1273
rect 626 1271 632 1272
rect 626 1267 627 1271
rect 631 1267 632 1271
rect 626 1266 632 1267
rect 550 1251 556 1252
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 550 1246 556 1247
rect 628 1244 630 1266
rect 672 1252 674 1273
rect 746 1271 752 1272
rect 746 1267 747 1271
rect 751 1267 752 1271
rect 746 1266 752 1267
rect 738 1263 744 1264
rect 738 1259 739 1263
rect 743 1259 744 1263
rect 738 1258 744 1259
rect 670 1251 676 1252
rect 670 1247 671 1251
rect 675 1247 676 1251
rect 670 1246 676 1247
rect 514 1243 520 1244
rect 514 1239 515 1243
rect 519 1239 520 1243
rect 514 1238 520 1239
rect 626 1243 632 1244
rect 626 1239 627 1243
rect 631 1239 632 1243
rect 626 1238 632 1239
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 438 1232 444 1233
rect 112 1203 114 1230
rect 438 1228 439 1232
rect 443 1228 444 1232
rect 438 1227 444 1228
rect 550 1232 556 1233
rect 550 1228 551 1232
rect 555 1228 556 1232
rect 550 1227 556 1228
rect 670 1232 676 1233
rect 670 1228 671 1232
rect 675 1228 676 1232
rect 670 1227 676 1228
rect 440 1203 442 1227
rect 552 1203 554 1227
rect 672 1203 674 1227
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 167 1202 171 1203
rect 167 1197 171 1198
rect 303 1202 307 1203
rect 303 1197 307 1198
rect 439 1202 443 1203
rect 439 1197 443 1198
rect 463 1202 467 1203
rect 463 1197 467 1198
rect 551 1202 555 1203
rect 551 1197 555 1198
rect 631 1202 635 1203
rect 631 1197 635 1198
rect 671 1202 675 1203
rect 671 1197 675 1198
rect 112 1170 114 1197
rect 168 1173 170 1197
rect 304 1173 306 1197
rect 464 1173 466 1197
rect 632 1173 634 1197
rect 166 1172 172 1173
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 166 1168 167 1172
rect 171 1168 172 1172
rect 166 1167 172 1168
rect 302 1172 308 1173
rect 302 1168 303 1172
rect 307 1168 308 1172
rect 302 1167 308 1168
rect 462 1172 468 1173
rect 462 1168 463 1172
rect 467 1168 468 1172
rect 462 1167 468 1168
rect 630 1172 636 1173
rect 630 1168 631 1172
rect 635 1168 636 1172
rect 630 1167 636 1168
rect 110 1164 116 1165
rect 740 1164 742 1258
rect 748 1244 750 1266
rect 800 1252 802 1273
rect 874 1271 880 1272
rect 874 1267 875 1271
rect 879 1267 880 1271
rect 874 1266 880 1267
rect 798 1251 804 1252
rect 798 1247 799 1251
rect 803 1247 804 1251
rect 798 1246 804 1247
rect 876 1244 878 1266
rect 936 1252 938 1273
rect 1080 1252 1082 1273
rect 1214 1271 1220 1272
rect 1214 1267 1215 1271
rect 1219 1267 1220 1271
rect 1214 1266 1220 1267
rect 934 1251 940 1252
rect 934 1247 935 1251
rect 939 1247 940 1251
rect 934 1246 940 1247
rect 1078 1251 1084 1252
rect 1078 1247 1079 1251
rect 1083 1247 1084 1251
rect 1078 1246 1084 1247
rect 1216 1244 1218 1266
rect 1232 1252 1234 1273
rect 1314 1271 1320 1272
rect 1314 1267 1315 1271
rect 1319 1267 1320 1271
rect 1314 1266 1320 1267
rect 1230 1251 1236 1252
rect 1230 1247 1231 1251
rect 1235 1247 1236 1251
rect 1230 1246 1236 1247
rect 1316 1244 1318 1266
rect 1392 1252 1394 1273
rect 1484 1272 1486 1314
rect 1558 1309 1564 1310
rect 1558 1305 1559 1309
rect 1563 1305 1564 1309
rect 1558 1304 1564 1305
rect 1560 1279 1562 1304
rect 1636 1288 1638 1314
rect 1702 1309 1708 1310
rect 1702 1305 1703 1309
rect 1707 1305 1708 1309
rect 1702 1304 1708 1305
rect 1626 1287 1632 1288
rect 1626 1283 1627 1287
rect 1631 1283 1632 1287
rect 1626 1282 1632 1283
rect 1634 1287 1640 1288
rect 1634 1283 1635 1287
rect 1639 1283 1640 1287
rect 1634 1282 1640 1283
rect 1551 1278 1555 1279
rect 1551 1273 1555 1274
rect 1559 1278 1563 1279
rect 1559 1273 1563 1274
rect 1482 1271 1488 1272
rect 1482 1267 1483 1271
rect 1487 1267 1488 1271
rect 1482 1266 1488 1267
rect 1552 1252 1554 1273
rect 1390 1251 1396 1252
rect 1390 1247 1391 1251
rect 1395 1247 1396 1251
rect 1390 1246 1396 1247
rect 1550 1251 1556 1252
rect 1550 1247 1551 1251
rect 1555 1247 1556 1251
rect 1550 1246 1556 1247
rect 1628 1244 1630 1282
rect 1704 1279 1706 1304
rect 1780 1288 1782 1314
rect 2048 1311 2050 1335
rect 2400 1311 2402 1336
rect 2047 1310 2051 1311
rect 1846 1309 1852 1310
rect 1846 1305 1847 1309
rect 1851 1305 1852 1309
rect 1846 1304 1852 1305
rect 2006 1308 2012 1309
rect 2006 1304 2007 1308
rect 2011 1304 2012 1308
rect 2047 1305 2051 1306
rect 2247 1310 2251 1311
rect 2247 1305 2251 1306
rect 2375 1310 2379 1311
rect 2375 1305 2379 1306
rect 2399 1310 2403 1311
rect 2399 1305 2403 1306
rect 1778 1287 1784 1288
rect 1778 1283 1779 1287
rect 1783 1283 1784 1287
rect 1778 1282 1784 1283
rect 1848 1279 1850 1304
rect 2006 1303 2012 1304
rect 2008 1279 2010 1303
rect 2048 1285 2050 1305
rect 2046 1284 2052 1285
rect 2248 1284 2250 1305
rect 2366 1303 2372 1304
rect 2366 1299 2367 1303
rect 2371 1299 2372 1303
rect 2366 1298 2372 1299
rect 2046 1280 2047 1284
rect 2051 1280 2052 1284
rect 2046 1279 2052 1280
rect 2246 1283 2252 1284
rect 2246 1279 2247 1283
rect 2251 1279 2252 1283
rect 1703 1278 1707 1279
rect 1703 1273 1707 1274
rect 1719 1278 1723 1279
rect 1719 1273 1723 1274
rect 1847 1278 1851 1279
rect 1847 1273 1851 1274
rect 2007 1278 2011 1279
rect 2246 1278 2252 1279
rect 2368 1276 2370 1298
rect 2376 1284 2378 1305
rect 2476 1304 2478 1346
rect 2484 1320 2486 1346
rect 2534 1341 2540 1342
rect 2534 1337 2535 1341
rect 2539 1337 2540 1341
rect 2534 1336 2540 1337
rect 2678 1341 2684 1342
rect 2678 1337 2679 1341
rect 2683 1337 2684 1341
rect 2678 1336 2684 1337
rect 2482 1319 2488 1320
rect 2482 1315 2483 1319
rect 2487 1315 2488 1319
rect 2482 1314 2488 1315
rect 2536 1311 2538 1336
rect 2680 1311 2682 1336
rect 2708 1320 2710 1422
rect 2758 1420 2764 1421
rect 2758 1416 2759 1420
rect 2763 1416 2764 1420
rect 2758 1415 2764 1416
rect 2894 1420 2900 1421
rect 2894 1416 2895 1420
rect 2899 1416 2900 1420
rect 2894 1415 2900 1416
rect 3030 1420 3036 1421
rect 3030 1416 3031 1420
rect 3035 1416 3036 1420
rect 3030 1415 3036 1416
rect 3174 1420 3180 1421
rect 3174 1416 3175 1420
rect 3179 1416 3180 1420
rect 3174 1415 3180 1416
rect 3310 1420 3316 1421
rect 3310 1416 3311 1420
rect 3315 1416 3316 1420
rect 3310 1415 3316 1416
rect 3446 1420 3452 1421
rect 3446 1416 3447 1420
rect 3451 1416 3452 1420
rect 3574 1419 3575 1423
rect 3579 1419 3580 1423
rect 3574 1418 3580 1419
rect 3582 1420 3588 1421
rect 3446 1415 3452 1416
rect 2760 1391 2762 1415
rect 2896 1391 2898 1415
rect 3032 1391 3034 1415
rect 3176 1391 3178 1415
rect 3312 1391 3314 1415
rect 3448 1391 3450 1415
rect 2759 1390 2763 1391
rect 2759 1385 2763 1386
rect 2823 1390 2827 1391
rect 2823 1385 2827 1386
rect 2895 1390 2899 1391
rect 2895 1385 2899 1386
rect 2967 1390 2971 1391
rect 2967 1385 2971 1386
rect 3031 1390 3035 1391
rect 3031 1385 3035 1386
rect 3111 1390 3115 1391
rect 3111 1385 3115 1386
rect 3175 1390 3179 1391
rect 3175 1385 3179 1386
rect 3255 1390 3259 1391
rect 3255 1385 3259 1386
rect 3311 1390 3315 1391
rect 3311 1385 3315 1386
rect 3407 1390 3411 1391
rect 3407 1385 3411 1386
rect 3447 1390 3451 1391
rect 3447 1385 3451 1386
rect 3559 1390 3563 1391
rect 3559 1385 3563 1386
rect 2824 1361 2826 1385
rect 2968 1361 2970 1385
rect 3112 1361 3114 1385
rect 3256 1361 3258 1385
rect 3408 1361 3410 1385
rect 3560 1361 3562 1385
rect 3576 1379 3578 1418
rect 3582 1416 3583 1420
rect 3587 1416 3588 1420
rect 3582 1415 3588 1416
rect 3718 1420 3724 1421
rect 3718 1416 3719 1420
rect 3723 1416 3724 1420
rect 3718 1415 3724 1416
rect 3584 1391 3586 1415
rect 3720 1391 3722 1415
rect 3583 1390 3587 1391
rect 3583 1385 3587 1386
rect 3711 1390 3715 1391
rect 3711 1385 3715 1386
rect 3719 1390 3723 1391
rect 3719 1385 3723 1386
rect 3576 1377 3586 1379
rect 2822 1360 2828 1361
rect 2822 1356 2823 1360
rect 2827 1356 2828 1360
rect 2822 1355 2828 1356
rect 2966 1360 2972 1361
rect 2966 1356 2967 1360
rect 2971 1356 2972 1360
rect 2966 1355 2972 1356
rect 3110 1360 3116 1361
rect 3110 1356 3111 1360
rect 3115 1356 3116 1360
rect 3110 1355 3116 1356
rect 3254 1360 3260 1361
rect 3254 1356 3255 1360
rect 3259 1356 3260 1360
rect 3254 1355 3260 1356
rect 3406 1360 3412 1361
rect 3406 1356 3407 1360
rect 3411 1356 3412 1360
rect 3406 1355 3412 1356
rect 3558 1360 3564 1361
rect 3558 1356 3559 1360
rect 3563 1356 3564 1360
rect 3558 1355 3564 1356
rect 2754 1351 2760 1352
rect 2754 1347 2755 1351
rect 2759 1347 2760 1351
rect 2754 1346 2760 1347
rect 2898 1351 2904 1352
rect 2898 1347 2899 1351
rect 2903 1347 2904 1351
rect 2898 1346 2904 1347
rect 2922 1351 2928 1352
rect 2922 1347 2923 1351
rect 2927 1347 2928 1351
rect 2922 1346 2928 1347
rect 3050 1351 3056 1352
rect 3050 1347 3051 1351
rect 3055 1347 3056 1351
rect 3050 1346 3056 1347
rect 3194 1351 3200 1352
rect 3194 1347 3195 1351
rect 3199 1347 3200 1351
rect 3194 1346 3200 1347
rect 3338 1351 3344 1352
rect 3338 1347 3339 1351
rect 3343 1347 3344 1351
rect 3338 1346 3344 1347
rect 2756 1320 2758 1346
rect 2822 1341 2828 1342
rect 2822 1337 2823 1341
rect 2827 1337 2828 1341
rect 2822 1336 2828 1337
rect 2706 1319 2712 1320
rect 2706 1315 2707 1319
rect 2711 1315 2712 1319
rect 2706 1314 2712 1315
rect 2754 1319 2760 1320
rect 2754 1315 2755 1319
rect 2759 1315 2760 1319
rect 2754 1314 2760 1315
rect 2824 1311 2826 1336
rect 2900 1320 2902 1346
rect 2924 1328 2926 1346
rect 2966 1341 2972 1342
rect 2966 1337 2967 1341
rect 2971 1337 2972 1341
rect 2966 1336 2972 1337
rect 2922 1327 2928 1328
rect 2922 1323 2923 1327
rect 2927 1323 2928 1327
rect 2922 1322 2928 1323
rect 2898 1319 2904 1320
rect 2898 1315 2899 1319
rect 2903 1315 2904 1319
rect 2898 1314 2904 1315
rect 2968 1311 2970 1336
rect 2511 1310 2515 1311
rect 2511 1305 2515 1306
rect 2535 1310 2539 1311
rect 2535 1305 2539 1306
rect 2647 1310 2651 1311
rect 2647 1305 2651 1306
rect 2679 1310 2683 1311
rect 2679 1305 2683 1306
rect 2791 1310 2795 1311
rect 2791 1305 2795 1306
rect 2823 1310 2827 1311
rect 2823 1305 2827 1306
rect 2943 1310 2947 1311
rect 2943 1305 2947 1306
rect 2967 1310 2971 1311
rect 2967 1305 2971 1306
rect 2474 1303 2480 1304
rect 2474 1299 2475 1303
rect 2479 1299 2480 1303
rect 2474 1298 2480 1299
rect 2512 1284 2514 1305
rect 2586 1303 2592 1304
rect 2586 1299 2587 1303
rect 2591 1299 2592 1303
rect 2586 1298 2592 1299
rect 2374 1283 2380 1284
rect 2374 1279 2375 1283
rect 2379 1279 2380 1283
rect 2374 1278 2380 1279
rect 2510 1283 2516 1284
rect 2510 1279 2511 1283
rect 2515 1279 2516 1283
rect 2510 1278 2516 1279
rect 2588 1276 2590 1298
rect 2648 1284 2650 1305
rect 2722 1303 2728 1304
rect 2722 1299 2723 1303
rect 2727 1299 2728 1303
rect 2722 1298 2728 1299
rect 2646 1283 2652 1284
rect 2646 1279 2647 1283
rect 2651 1279 2652 1283
rect 2646 1278 2652 1279
rect 2724 1276 2726 1298
rect 2730 1295 2736 1296
rect 2730 1291 2731 1295
rect 2735 1291 2736 1295
rect 2730 1290 2736 1291
rect 2732 1276 2734 1290
rect 2792 1284 2794 1305
rect 2944 1284 2946 1305
rect 3052 1304 3054 1346
rect 3110 1341 3116 1342
rect 3110 1337 3111 1341
rect 3115 1337 3116 1341
rect 3110 1336 3116 1337
rect 3112 1311 3114 1336
rect 3196 1320 3198 1346
rect 3254 1341 3260 1342
rect 3254 1337 3255 1341
rect 3259 1337 3260 1341
rect 3254 1336 3260 1337
rect 3194 1319 3200 1320
rect 3194 1315 3195 1319
rect 3199 1315 3200 1319
rect 3194 1314 3200 1315
rect 3256 1311 3258 1336
rect 3340 1320 3342 1346
rect 3406 1341 3412 1342
rect 3406 1337 3407 1341
rect 3411 1337 3412 1341
rect 3406 1336 3412 1337
rect 3558 1341 3564 1342
rect 3558 1337 3559 1341
rect 3563 1337 3564 1341
rect 3558 1336 3564 1337
rect 3338 1319 3344 1320
rect 3338 1315 3339 1319
rect 3343 1315 3344 1319
rect 3338 1314 3344 1315
rect 3408 1311 3410 1336
rect 3560 1311 3562 1336
rect 3584 1320 3586 1377
rect 3712 1361 3714 1385
rect 3710 1360 3716 1361
rect 3710 1356 3711 1360
rect 3715 1356 3716 1360
rect 3710 1355 3716 1356
rect 3800 1352 3802 1473
rect 3840 1467 3842 1500
rect 3839 1466 3843 1467
rect 3839 1461 3843 1462
rect 3840 1440 3842 1461
rect 3908 1460 3910 1510
rect 3916 1484 3918 1666
rect 3942 1660 3948 1661
rect 3942 1656 3943 1660
rect 3947 1656 3948 1660
rect 3942 1655 3948 1656
rect 3944 1631 3946 1655
rect 3943 1630 3947 1631
rect 3943 1625 3947 1626
rect 3944 1605 3946 1625
rect 3942 1604 3948 1605
rect 3942 1600 3943 1604
rect 3947 1600 3948 1604
rect 3942 1599 3948 1600
rect 3942 1587 3948 1588
rect 3942 1583 3943 1587
rect 3947 1583 3948 1587
rect 3942 1582 3948 1583
rect 3944 1555 3946 1582
rect 3943 1554 3947 1555
rect 3943 1549 3947 1550
rect 3944 1522 3946 1549
rect 3942 1521 3948 1522
rect 3942 1517 3943 1521
rect 3947 1517 3948 1521
rect 3942 1516 3948 1517
rect 3942 1504 3948 1505
rect 3942 1500 3943 1504
rect 3947 1500 3948 1504
rect 3942 1499 3948 1500
rect 3914 1483 3920 1484
rect 3914 1479 3915 1483
rect 3919 1479 3920 1483
rect 3914 1478 3920 1479
rect 3944 1467 3946 1499
rect 3943 1466 3947 1467
rect 3943 1461 3947 1462
rect 3906 1459 3912 1460
rect 3906 1455 3907 1459
rect 3911 1455 3912 1459
rect 3906 1454 3912 1455
rect 3944 1441 3946 1461
rect 3942 1440 3948 1441
rect 3838 1439 3844 1440
rect 3838 1435 3839 1439
rect 3843 1435 3844 1439
rect 3942 1436 3943 1440
rect 3947 1436 3948 1440
rect 3942 1435 3948 1436
rect 3838 1434 3844 1435
rect 3906 1423 3912 1424
rect 3838 1420 3844 1421
rect 3838 1416 3839 1420
rect 3843 1416 3844 1420
rect 3906 1419 3907 1423
rect 3911 1419 3912 1423
rect 3906 1418 3912 1419
rect 3942 1423 3948 1424
rect 3942 1419 3943 1423
rect 3947 1419 3948 1423
rect 3942 1418 3948 1419
rect 3838 1415 3844 1416
rect 3840 1391 3842 1415
rect 3839 1390 3843 1391
rect 3839 1385 3843 1386
rect 3840 1361 3842 1385
rect 3838 1360 3844 1361
rect 3838 1356 3839 1360
rect 3843 1356 3844 1360
rect 3838 1355 3844 1356
rect 3634 1351 3640 1352
rect 3634 1347 3635 1351
rect 3639 1347 3640 1351
rect 3634 1346 3640 1347
rect 3798 1351 3804 1352
rect 3798 1347 3799 1351
rect 3803 1347 3804 1351
rect 3798 1346 3804 1347
rect 3636 1320 3638 1346
rect 3710 1341 3716 1342
rect 3710 1337 3711 1341
rect 3715 1337 3716 1341
rect 3710 1336 3716 1337
rect 3838 1341 3844 1342
rect 3838 1337 3839 1341
rect 3843 1337 3844 1341
rect 3838 1336 3844 1337
rect 3582 1319 3588 1320
rect 3582 1315 3583 1319
rect 3587 1315 3588 1319
rect 3582 1314 3588 1315
rect 3634 1319 3640 1320
rect 3634 1315 3635 1319
rect 3639 1315 3640 1319
rect 3634 1314 3640 1315
rect 3712 1311 3714 1336
rect 3840 1311 3842 1336
rect 3111 1310 3115 1311
rect 3111 1305 3115 1306
rect 3255 1310 3259 1311
rect 3255 1305 3259 1306
rect 3287 1310 3291 1311
rect 3287 1305 3291 1306
rect 3407 1310 3411 1311
rect 3407 1305 3411 1306
rect 3471 1310 3475 1311
rect 3471 1305 3475 1306
rect 3559 1310 3563 1311
rect 3559 1305 3563 1306
rect 3663 1310 3667 1311
rect 3663 1305 3667 1306
rect 3711 1310 3715 1311
rect 3711 1305 3715 1306
rect 3839 1310 3843 1311
rect 3839 1305 3843 1306
rect 3050 1303 3056 1304
rect 3050 1299 3051 1303
rect 3055 1299 3056 1303
rect 3050 1298 3056 1299
rect 3078 1303 3084 1304
rect 3078 1299 3079 1303
rect 3083 1299 3084 1303
rect 3078 1298 3084 1299
rect 2790 1283 2796 1284
rect 2790 1279 2791 1283
rect 2795 1279 2796 1283
rect 2790 1278 2796 1279
rect 2942 1283 2948 1284
rect 2942 1279 2943 1283
rect 2947 1279 2948 1283
rect 2942 1278 2948 1279
rect 3080 1276 3082 1298
rect 3112 1284 3114 1305
rect 3186 1303 3192 1304
rect 3186 1299 3187 1303
rect 3191 1299 3192 1303
rect 3186 1298 3192 1299
rect 3110 1283 3116 1284
rect 3110 1279 3111 1283
rect 3115 1279 3116 1283
rect 3110 1278 3116 1279
rect 3188 1276 3190 1298
rect 3288 1284 3290 1305
rect 3362 1303 3368 1304
rect 3362 1299 3363 1303
rect 3367 1299 3368 1303
rect 3362 1298 3368 1299
rect 3286 1283 3292 1284
rect 3286 1279 3287 1283
rect 3291 1279 3292 1283
rect 3286 1278 3292 1279
rect 3364 1276 3366 1298
rect 3472 1284 3474 1305
rect 3546 1303 3552 1304
rect 3546 1299 3547 1303
rect 3551 1299 3552 1303
rect 3546 1298 3552 1299
rect 3470 1283 3476 1284
rect 3470 1279 3471 1283
rect 3475 1279 3476 1283
rect 3470 1278 3476 1279
rect 3548 1276 3550 1298
rect 3664 1284 3666 1305
rect 3840 1284 3842 1305
rect 3908 1304 3910 1418
rect 3944 1391 3946 1418
rect 3943 1390 3947 1391
rect 3943 1385 3947 1386
rect 3944 1358 3946 1385
rect 3942 1357 3948 1358
rect 3942 1353 3943 1357
rect 3947 1353 3948 1357
rect 3942 1352 3948 1353
rect 3942 1340 3948 1341
rect 3942 1336 3943 1340
rect 3947 1336 3948 1340
rect 3942 1335 3948 1336
rect 3914 1319 3920 1320
rect 3914 1315 3915 1319
rect 3919 1315 3920 1319
rect 3914 1314 3920 1315
rect 3906 1303 3912 1304
rect 3906 1299 3907 1303
rect 3911 1299 3912 1303
rect 3906 1298 3912 1299
rect 3662 1283 3668 1284
rect 3662 1279 3663 1283
rect 3667 1279 3668 1283
rect 3662 1278 3668 1279
rect 3838 1283 3844 1284
rect 3838 1279 3839 1283
rect 3843 1279 3844 1283
rect 3838 1278 3844 1279
rect 3916 1276 3918 1314
rect 3944 1311 3946 1335
rect 3943 1310 3947 1311
rect 3943 1305 3947 1306
rect 3944 1285 3946 1305
rect 3942 1284 3948 1285
rect 3942 1280 3943 1284
rect 3947 1280 3948 1284
rect 3942 1279 3948 1280
rect 2007 1273 2011 1274
rect 2366 1275 2372 1276
rect 1720 1252 1722 1273
rect 1770 1271 1776 1272
rect 1770 1267 1771 1271
rect 1775 1267 1776 1271
rect 1770 1266 1776 1267
rect 1718 1251 1724 1252
rect 1718 1247 1719 1251
rect 1723 1247 1724 1251
rect 1718 1246 1724 1247
rect 746 1243 752 1244
rect 746 1239 747 1243
rect 751 1239 752 1243
rect 746 1238 752 1239
rect 874 1243 880 1244
rect 874 1239 875 1243
rect 879 1239 880 1243
rect 874 1238 880 1239
rect 1070 1243 1076 1244
rect 1070 1239 1071 1243
rect 1075 1239 1076 1243
rect 1070 1238 1076 1239
rect 1214 1243 1220 1244
rect 1214 1239 1215 1243
rect 1219 1239 1220 1243
rect 1214 1238 1220 1239
rect 1314 1243 1320 1244
rect 1314 1239 1315 1243
rect 1319 1239 1320 1243
rect 1314 1238 1320 1239
rect 1626 1243 1632 1244
rect 1626 1239 1627 1243
rect 1631 1239 1632 1243
rect 1626 1238 1632 1239
rect 798 1232 804 1233
rect 798 1228 799 1232
rect 803 1228 804 1232
rect 798 1227 804 1228
rect 934 1232 940 1233
rect 934 1228 935 1232
rect 939 1228 940 1232
rect 934 1227 940 1228
rect 800 1203 802 1227
rect 936 1203 938 1227
rect 799 1202 803 1203
rect 799 1197 803 1198
rect 807 1202 811 1203
rect 807 1197 811 1198
rect 935 1202 939 1203
rect 935 1197 939 1198
rect 983 1202 987 1203
rect 983 1197 987 1198
rect 808 1173 810 1197
rect 984 1173 986 1197
rect 806 1172 812 1173
rect 806 1168 807 1172
rect 811 1168 812 1172
rect 806 1167 812 1168
rect 982 1172 988 1173
rect 982 1168 983 1172
rect 987 1168 988 1172
rect 982 1167 988 1168
rect 242 1163 248 1164
rect 242 1159 243 1163
rect 247 1159 248 1163
rect 242 1158 248 1159
rect 378 1163 384 1164
rect 378 1159 379 1163
rect 383 1159 384 1163
rect 378 1158 384 1159
rect 538 1163 544 1164
rect 538 1159 539 1163
rect 543 1159 544 1163
rect 538 1158 544 1159
rect 706 1163 712 1164
rect 706 1159 707 1163
rect 711 1159 712 1163
rect 706 1158 712 1159
rect 738 1163 744 1164
rect 738 1159 739 1163
rect 743 1159 744 1163
rect 738 1158 744 1159
rect 166 1153 172 1154
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 166 1149 167 1153
rect 171 1149 172 1153
rect 166 1148 172 1149
rect 110 1147 116 1148
rect 112 1123 114 1147
rect 168 1123 170 1148
rect 244 1132 246 1158
rect 302 1153 308 1154
rect 302 1149 303 1153
rect 307 1149 308 1153
rect 302 1148 308 1149
rect 242 1131 248 1132
rect 242 1127 243 1131
rect 247 1127 248 1131
rect 242 1126 248 1127
rect 304 1123 306 1148
rect 380 1132 382 1158
rect 462 1153 468 1154
rect 462 1149 463 1153
rect 467 1149 468 1153
rect 462 1148 468 1149
rect 378 1131 384 1132
rect 378 1127 379 1131
rect 383 1127 384 1131
rect 378 1126 384 1127
rect 464 1123 466 1148
rect 540 1132 542 1158
rect 630 1153 636 1154
rect 630 1149 631 1153
rect 635 1149 636 1153
rect 630 1148 636 1149
rect 538 1131 544 1132
rect 538 1127 539 1131
rect 543 1127 544 1131
rect 538 1126 544 1127
rect 618 1123 624 1124
rect 632 1123 634 1148
rect 708 1132 710 1158
rect 806 1153 812 1154
rect 806 1149 807 1153
rect 811 1149 812 1153
rect 806 1148 812 1149
rect 982 1153 988 1154
rect 982 1149 983 1153
rect 987 1149 988 1153
rect 982 1148 988 1149
rect 706 1131 712 1132
rect 706 1127 707 1131
rect 711 1127 712 1131
rect 706 1126 712 1127
rect 808 1123 810 1148
rect 984 1123 986 1148
rect 1072 1132 1074 1238
rect 1078 1232 1084 1233
rect 1078 1228 1079 1232
rect 1083 1228 1084 1232
rect 1078 1227 1084 1228
rect 1230 1232 1236 1233
rect 1230 1228 1231 1232
rect 1235 1228 1236 1232
rect 1230 1227 1236 1228
rect 1390 1232 1396 1233
rect 1390 1228 1391 1232
rect 1395 1228 1396 1232
rect 1390 1227 1396 1228
rect 1550 1232 1556 1233
rect 1550 1228 1551 1232
rect 1555 1228 1556 1232
rect 1550 1227 1556 1228
rect 1718 1232 1724 1233
rect 1718 1228 1719 1232
rect 1723 1228 1724 1232
rect 1718 1227 1724 1228
rect 1080 1203 1082 1227
rect 1232 1203 1234 1227
rect 1392 1203 1394 1227
rect 1552 1203 1554 1227
rect 1720 1203 1722 1227
rect 1079 1202 1083 1203
rect 1079 1197 1083 1198
rect 1159 1202 1163 1203
rect 1159 1197 1163 1198
rect 1231 1202 1235 1203
rect 1231 1197 1235 1198
rect 1335 1202 1339 1203
rect 1335 1197 1339 1198
rect 1391 1202 1395 1203
rect 1391 1197 1395 1198
rect 1511 1202 1515 1203
rect 1511 1197 1515 1198
rect 1551 1202 1555 1203
rect 1551 1197 1555 1198
rect 1695 1202 1699 1203
rect 1695 1197 1699 1198
rect 1719 1202 1723 1203
rect 1719 1197 1723 1198
rect 1160 1173 1162 1197
rect 1336 1173 1338 1197
rect 1512 1173 1514 1197
rect 1696 1173 1698 1197
rect 1158 1172 1164 1173
rect 1158 1168 1159 1172
rect 1163 1168 1164 1172
rect 1158 1167 1164 1168
rect 1334 1172 1340 1173
rect 1334 1168 1335 1172
rect 1339 1168 1340 1172
rect 1334 1167 1340 1168
rect 1510 1172 1516 1173
rect 1510 1168 1511 1172
rect 1515 1168 1516 1172
rect 1510 1167 1516 1168
rect 1694 1172 1700 1173
rect 1694 1168 1695 1172
rect 1699 1168 1700 1172
rect 1694 1167 1700 1168
rect 1772 1164 1774 1266
rect 2008 1253 2010 1273
rect 2322 1271 2328 1272
rect 2046 1267 2052 1268
rect 2046 1263 2047 1267
rect 2051 1263 2052 1267
rect 2322 1267 2323 1271
rect 2327 1267 2328 1271
rect 2366 1271 2367 1275
rect 2371 1271 2372 1275
rect 2366 1270 2372 1271
rect 2586 1275 2592 1276
rect 2586 1271 2587 1275
rect 2591 1271 2592 1275
rect 2586 1270 2592 1271
rect 2722 1275 2728 1276
rect 2722 1271 2723 1275
rect 2727 1271 2728 1275
rect 2722 1270 2728 1271
rect 2730 1275 2736 1276
rect 2730 1271 2731 1275
rect 2735 1271 2736 1275
rect 2730 1270 2736 1271
rect 3078 1275 3084 1276
rect 3078 1271 3079 1275
rect 3083 1271 3084 1275
rect 3078 1270 3084 1271
rect 3186 1275 3192 1276
rect 3186 1271 3187 1275
rect 3191 1271 3192 1275
rect 3186 1270 3192 1271
rect 3362 1275 3368 1276
rect 3362 1271 3363 1275
rect 3367 1271 3368 1275
rect 3362 1270 3368 1271
rect 3546 1275 3552 1276
rect 3546 1271 3547 1275
rect 3551 1271 3552 1275
rect 3546 1270 3552 1271
rect 3610 1275 3616 1276
rect 3610 1271 3611 1275
rect 3615 1271 3616 1275
rect 3610 1270 3616 1271
rect 3914 1275 3920 1276
rect 3914 1271 3915 1275
rect 3919 1271 3920 1275
rect 3914 1270 3920 1271
rect 2322 1266 2328 1267
rect 2046 1262 2052 1263
rect 2246 1264 2252 1265
rect 2006 1252 2012 1253
rect 2006 1248 2007 1252
rect 2011 1248 2012 1252
rect 2006 1247 2012 1248
rect 2006 1235 2012 1236
rect 2006 1231 2007 1235
rect 2011 1231 2012 1235
rect 2048 1231 2050 1262
rect 2246 1260 2247 1264
rect 2251 1260 2252 1264
rect 2246 1259 2252 1260
rect 2248 1231 2250 1259
rect 2006 1230 2012 1231
rect 2047 1230 2051 1231
rect 2008 1203 2010 1230
rect 2047 1225 2051 1226
rect 2071 1230 2075 1231
rect 2071 1225 2075 1226
rect 2183 1230 2187 1231
rect 2183 1225 2187 1226
rect 2247 1230 2251 1231
rect 2247 1225 2251 1226
rect 2303 1230 2307 1231
rect 2303 1225 2307 1226
rect 2007 1202 2011 1203
rect 2048 1198 2050 1225
rect 2072 1201 2074 1225
rect 2184 1201 2186 1225
rect 2304 1201 2306 1225
rect 2070 1200 2076 1201
rect 2007 1197 2011 1198
rect 2046 1197 2052 1198
rect 2008 1170 2010 1197
rect 2046 1193 2047 1197
rect 2051 1193 2052 1197
rect 2070 1196 2071 1200
rect 2075 1196 2076 1200
rect 2070 1195 2076 1196
rect 2182 1200 2188 1201
rect 2182 1196 2183 1200
rect 2187 1196 2188 1200
rect 2182 1195 2188 1196
rect 2302 1200 2308 1201
rect 2302 1196 2303 1200
rect 2307 1196 2308 1200
rect 2302 1195 2308 1196
rect 2046 1192 2052 1193
rect 2146 1191 2152 1192
rect 2146 1187 2147 1191
rect 2151 1187 2152 1191
rect 2146 1186 2152 1187
rect 2258 1191 2264 1192
rect 2258 1187 2259 1191
rect 2263 1187 2264 1191
rect 2258 1186 2264 1187
rect 2070 1181 2076 1182
rect 2046 1180 2052 1181
rect 2046 1176 2047 1180
rect 2051 1176 2052 1180
rect 2070 1177 2071 1181
rect 2075 1177 2076 1181
rect 2070 1176 2076 1177
rect 2046 1175 2052 1176
rect 2006 1169 2012 1170
rect 2006 1165 2007 1169
rect 2011 1165 2012 1169
rect 2006 1164 2012 1165
rect 1122 1163 1128 1164
rect 1122 1159 1123 1163
rect 1127 1159 1128 1163
rect 1122 1158 1128 1159
rect 1234 1163 1240 1164
rect 1234 1159 1235 1163
rect 1239 1159 1240 1163
rect 1234 1158 1240 1159
rect 1410 1163 1416 1164
rect 1410 1159 1411 1163
rect 1415 1159 1416 1163
rect 1410 1158 1416 1159
rect 1586 1163 1592 1164
rect 1586 1159 1587 1163
rect 1591 1159 1592 1163
rect 1586 1158 1592 1159
rect 1770 1163 1776 1164
rect 1770 1159 1771 1163
rect 1775 1159 1776 1163
rect 1770 1158 1776 1159
rect 1124 1132 1126 1158
rect 1158 1153 1164 1154
rect 1158 1149 1159 1153
rect 1163 1149 1164 1153
rect 1158 1148 1164 1149
rect 1070 1131 1076 1132
rect 1070 1127 1071 1131
rect 1075 1127 1076 1131
rect 1070 1126 1076 1127
rect 1122 1131 1128 1132
rect 1122 1127 1123 1131
rect 1127 1127 1128 1131
rect 1122 1126 1128 1127
rect 1160 1123 1162 1148
rect 111 1122 115 1123
rect 111 1117 115 1118
rect 135 1122 139 1123
rect 135 1117 139 1118
rect 167 1122 171 1123
rect 167 1117 171 1118
rect 239 1122 243 1123
rect 239 1117 243 1118
rect 303 1122 307 1123
rect 303 1117 307 1118
rect 375 1122 379 1123
rect 375 1117 379 1118
rect 463 1122 467 1123
rect 463 1117 467 1118
rect 527 1122 531 1123
rect 618 1119 619 1123
rect 623 1119 624 1123
rect 618 1118 624 1119
rect 631 1122 635 1123
rect 527 1117 531 1118
rect 112 1097 114 1117
rect 110 1096 116 1097
rect 136 1096 138 1117
rect 202 1115 208 1116
rect 202 1111 203 1115
rect 207 1111 208 1115
rect 202 1110 208 1111
rect 210 1115 216 1116
rect 210 1111 211 1115
rect 215 1111 216 1115
rect 210 1110 216 1111
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 134 1095 140 1096
rect 134 1091 135 1095
rect 139 1091 140 1095
rect 134 1090 140 1091
rect 110 1079 116 1080
rect 110 1075 111 1079
rect 115 1075 116 1079
rect 110 1074 116 1075
rect 134 1076 140 1077
rect 112 1047 114 1074
rect 134 1072 135 1076
rect 139 1072 140 1076
rect 134 1071 140 1072
rect 136 1047 138 1071
rect 111 1046 115 1047
rect 111 1041 115 1042
rect 135 1046 139 1047
rect 135 1041 139 1042
rect 112 1014 114 1041
rect 136 1017 138 1041
rect 204 1024 206 1110
rect 212 1088 214 1110
rect 240 1096 242 1117
rect 314 1115 320 1116
rect 314 1111 315 1115
rect 319 1111 320 1115
rect 314 1110 320 1111
rect 238 1095 244 1096
rect 238 1091 239 1095
rect 243 1091 244 1095
rect 238 1090 244 1091
rect 316 1088 318 1110
rect 376 1096 378 1117
rect 450 1115 456 1116
rect 450 1111 451 1115
rect 455 1111 456 1115
rect 450 1110 456 1111
rect 374 1095 380 1096
rect 374 1091 375 1095
rect 379 1091 380 1095
rect 374 1090 380 1091
rect 452 1088 454 1110
rect 528 1096 530 1117
rect 602 1115 608 1116
rect 602 1111 603 1115
rect 607 1111 608 1115
rect 602 1110 608 1111
rect 526 1095 532 1096
rect 526 1091 527 1095
rect 531 1091 532 1095
rect 526 1090 532 1091
rect 604 1088 606 1110
rect 620 1088 622 1118
rect 631 1117 635 1118
rect 695 1122 699 1123
rect 695 1117 699 1118
rect 807 1122 811 1123
rect 807 1117 811 1118
rect 863 1122 867 1123
rect 863 1117 867 1118
rect 983 1122 987 1123
rect 983 1117 987 1118
rect 1039 1122 1043 1123
rect 1039 1117 1043 1118
rect 1159 1122 1163 1123
rect 1159 1117 1163 1118
rect 1215 1122 1219 1123
rect 1215 1117 1219 1118
rect 696 1096 698 1117
rect 864 1096 866 1117
rect 946 1115 952 1116
rect 946 1111 947 1115
rect 951 1111 952 1115
rect 946 1110 952 1111
rect 694 1095 700 1096
rect 694 1091 695 1095
rect 699 1091 700 1095
rect 694 1090 700 1091
rect 862 1095 868 1096
rect 862 1091 863 1095
rect 867 1091 868 1095
rect 862 1090 868 1091
rect 948 1088 950 1110
rect 1040 1096 1042 1117
rect 1216 1096 1218 1117
rect 1236 1116 1238 1158
rect 1334 1153 1340 1154
rect 1334 1149 1335 1153
rect 1339 1149 1340 1153
rect 1334 1148 1340 1149
rect 1336 1123 1338 1148
rect 1412 1132 1414 1158
rect 1510 1153 1516 1154
rect 1510 1149 1511 1153
rect 1515 1149 1516 1153
rect 1510 1148 1516 1149
rect 1410 1131 1416 1132
rect 1410 1127 1411 1131
rect 1415 1127 1416 1131
rect 1410 1126 1416 1127
rect 1512 1123 1514 1148
rect 1588 1132 1590 1158
rect 1694 1153 1700 1154
rect 1694 1149 1695 1153
rect 1699 1149 1700 1153
rect 1694 1148 1700 1149
rect 2006 1152 2012 1153
rect 2006 1148 2007 1152
rect 2011 1148 2012 1152
rect 2048 1151 2050 1175
rect 2072 1151 2074 1176
rect 2148 1160 2150 1186
rect 2182 1181 2188 1182
rect 2182 1177 2183 1181
rect 2187 1177 2188 1181
rect 2182 1176 2188 1177
rect 2146 1159 2152 1160
rect 2146 1155 2147 1159
rect 2151 1155 2152 1159
rect 2146 1154 2152 1155
rect 2184 1151 2186 1176
rect 1586 1131 1592 1132
rect 1586 1127 1587 1131
rect 1591 1127 1592 1131
rect 1586 1126 1592 1127
rect 1696 1123 1698 1148
rect 2006 1147 2012 1148
rect 2047 1150 2051 1151
rect 2008 1123 2010 1147
rect 2047 1145 2051 1146
rect 2071 1150 2075 1151
rect 2071 1145 2075 1146
rect 2183 1150 2187 1151
rect 2183 1145 2187 1146
rect 2199 1150 2203 1151
rect 2199 1145 2203 1146
rect 2048 1125 2050 1145
rect 2046 1124 2052 1125
rect 2072 1124 2074 1145
rect 2200 1124 2202 1145
rect 2260 1144 2262 1186
rect 2302 1181 2308 1182
rect 2302 1177 2303 1181
rect 2307 1177 2308 1181
rect 2302 1176 2308 1177
rect 2304 1151 2306 1176
rect 2324 1160 2326 1266
rect 2374 1264 2380 1265
rect 2374 1260 2375 1264
rect 2379 1260 2380 1264
rect 2374 1259 2380 1260
rect 2510 1264 2516 1265
rect 2510 1260 2511 1264
rect 2515 1260 2516 1264
rect 2510 1259 2516 1260
rect 2646 1264 2652 1265
rect 2646 1260 2647 1264
rect 2651 1260 2652 1264
rect 2646 1259 2652 1260
rect 2790 1264 2796 1265
rect 2790 1260 2791 1264
rect 2795 1260 2796 1264
rect 2790 1259 2796 1260
rect 2942 1264 2948 1265
rect 2942 1260 2943 1264
rect 2947 1260 2948 1264
rect 2942 1259 2948 1260
rect 3110 1264 3116 1265
rect 3110 1260 3111 1264
rect 3115 1260 3116 1264
rect 3110 1259 3116 1260
rect 3286 1264 3292 1265
rect 3286 1260 3287 1264
rect 3291 1260 3292 1264
rect 3286 1259 3292 1260
rect 3470 1264 3476 1265
rect 3470 1260 3471 1264
rect 3475 1260 3476 1264
rect 3470 1259 3476 1260
rect 2376 1231 2378 1259
rect 2512 1231 2514 1259
rect 2648 1231 2650 1259
rect 2792 1231 2794 1259
rect 2944 1231 2946 1259
rect 3112 1231 3114 1259
rect 3288 1231 3290 1259
rect 3472 1231 3474 1259
rect 2375 1230 2379 1231
rect 2375 1225 2379 1226
rect 2431 1230 2435 1231
rect 2431 1225 2435 1226
rect 2511 1230 2515 1231
rect 2511 1225 2515 1226
rect 2559 1230 2563 1231
rect 2559 1225 2563 1226
rect 2647 1230 2651 1231
rect 2647 1225 2651 1226
rect 2711 1230 2715 1231
rect 2711 1225 2715 1226
rect 2791 1230 2795 1231
rect 2791 1225 2795 1226
rect 2887 1230 2891 1231
rect 2887 1225 2891 1226
rect 2943 1230 2947 1231
rect 2943 1225 2947 1226
rect 3087 1230 3091 1231
rect 3087 1225 3091 1226
rect 3111 1230 3115 1231
rect 3111 1225 3115 1226
rect 3287 1230 3291 1231
rect 3287 1225 3291 1226
rect 3311 1230 3315 1231
rect 3311 1225 3315 1226
rect 3471 1230 3475 1231
rect 3471 1225 3475 1226
rect 3543 1230 3547 1231
rect 3543 1225 3547 1226
rect 2432 1201 2434 1225
rect 2560 1201 2562 1225
rect 2712 1201 2714 1225
rect 2888 1201 2890 1225
rect 3088 1201 3090 1225
rect 3312 1201 3314 1225
rect 3544 1201 3546 1225
rect 2430 1200 2436 1201
rect 2430 1196 2431 1200
rect 2435 1196 2436 1200
rect 2430 1195 2436 1196
rect 2558 1200 2564 1201
rect 2558 1196 2559 1200
rect 2563 1196 2564 1200
rect 2558 1195 2564 1196
rect 2710 1200 2716 1201
rect 2710 1196 2711 1200
rect 2715 1196 2716 1200
rect 2710 1195 2716 1196
rect 2886 1200 2892 1201
rect 2886 1196 2887 1200
rect 2891 1196 2892 1200
rect 2886 1195 2892 1196
rect 3086 1200 3092 1201
rect 3086 1196 3087 1200
rect 3091 1196 3092 1200
rect 3086 1195 3092 1196
rect 3310 1200 3316 1201
rect 3310 1196 3311 1200
rect 3315 1196 3316 1200
rect 3310 1195 3316 1196
rect 3542 1200 3548 1201
rect 3542 1196 3543 1200
rect 3547 1196 3548 1200
rect 3542 1195 3548 1196
rect 2378 1191 2384 1192
rect 2378 1187 2379 1191
rect 2383 1187 2384 1191
rect 2378 1186 2384 1187
rect 2506 1191 2512 1192
rect 2506 1187 2507 1191
rect 2511 1187 2512 1191
rect 2506 1186 2512 1187
rect 2514 1191 2520 1192
rect 2514 1187 2515 1191
rect 2519 1187 2520 1191
rect 2514 1186 2520 1187
rect 2778 1191 2784 1192
rect 2778 1187 2779 1191
rect 2783 1187 2784 1191
rect 2778 1186 2784 1187
rect 2794 1191 2800 1192
rect 2794 1187 2795 1191
rect 2799 1187 2800 1191
rect 2794 1186 2800 1187
rect 2970 1191 2976 1192
rect 2970 1187 2971 1191
rect 2975 1187 2976 1191
rect 2970 1186 2976 1187
rect 3170 1191 3176 1192
rect 3170 1187 3171 1191
rect 3175 1187 3176 1191
rect 3170 1186 3176 1187
rect 3394 1191 3400 1192
rect 3394 1187 3395 1191
rect 3399 1187 3400 1191
rect 3394 1186 3400 1187
rect 2380 1160 2382 1186
rect 2430 1181 2436 1182
rect 2430 1177 2431 1181
rect 2435 1177 2436 1181
rect 2430 1176 2436 1177
rect 2322 1159 2328 1160
rect 2322 1155 2323 1159
rect 2327 1155 2328 1159
rect 2322 1154 2328 1155
rect 2378 1159 2384 1160
rect 2378 1155 2379 1159
rect 2383 1155 2384 1159
rect 2378 1154 2384 1155
rect 2432 1151 2434 1176
rect 2508 1160 2510 1186
rect 2516 1168 2518 1186
rect 2558 1181 2564 1182
rect 2558 1177 2559 1181
rect 2563 1177 2564 1181
rect 2558 1176 2564 1177
rect 2710 1181 2716 1182
rect 2710 1177 2711 1181
rect 2715 1177 2716 1181
rect 2710 1176 2716 1177
rect 2514 1167 2520 1168
rect 2514 1163 2515 1167
rect 2519 1163 2520 1167
rect 2514 1162 2520 1163
rect 2506 1159 2512 1160
rect 2506 1155 2507 1159
rect 2511 1155 2512 1159
rect 2506 1154 2512 1155
rect 2560 1151 2562 1176
rect 2712 1151 2714 1176
rect 2303 1150 2307 1151
rect 2303 1145 2307 1146
rect 2351 1150 2355 1151
rect 2351 1145 2355 1146
rect 2431 1150 2435 1151
rect 2431 1145 2435 1146
rect 2511 1150 2515 1151
rect 2511 1145 2515 1146
rect 2559 1150 2563 1151
rect 2559 1145 2563 1146
rect 2679 1150 2683 1151
rect 2679 1145 2683 1146
rect 2711 1150 2715 1151
rect 2711 1145 2715 1146
rect 2258 1143 2264 1144
rect 2258 1139 2259 1143
rect 2263 1139 2264 1143
rect 2258 1138 2264 1139
rect 2274 1143 2280 1144
rect 2274 1139 2275 1143
rect 2279 1139 2280 1143
rect 2274 1138 2280 1139
rect 1335 1122 1339 1123
rect 1335 1117 1339 1118
rect 1391 1122 1395 1123
rect 1391 1117 1395 1118
rect 1511 1122 1515 1123
rect 1511 1117 1515 1118
rect 1567 1122 1571 1123
rect 1567 1117 1571 1118
rect 1695 1122 1699 1123
rect 1695 1117 1699 1118
rect 1743 1122 1747 1123
rect 1743 1117 1747 1118
rect 1903 1122 1907 1123
rect 1903 1117 1907 1118
rect 2007 1122 2011 1123
rect 2046 1120 2047 1124
rect 2051 1120 2052 1124
rect 2046 1119 2052 1120
rect 2070 1123 2076 1124
rect 2070 1119 2071 1123
rect 2075 1119 2076 1123
rect 2070 1118 2076 1119
rect 2198 1123 2204 1124
rect 2198 1119 2199 1123
rect 2203 1119 2204 1123
rect 2198 1118 2204 1119
rect 2007 1117 2011 1118
rect 1234 1115 1240 1116
rect 1234 1111 1235 1115
rect 1239 1111 1240 1115
rect 1234 1110 1240 1111
rect 1392 1096 1394 1117
rect 1454 1115 1460 1116
rect 1454 1111 1455 1115
rect 1459 1111 1460 1115
rect 1454 1110 1460 1111
rect 1466 1115 1472 1116
rect 1466 1111 1467 1115
rect 1471 1111 1472 1115
rect 1466 1110 1472 1111
rect 1038 1095 1044 1096
rect 1038 1091 1039 1095
rect 1043 1091 1044 1095
rect 1038 1090 1044 1091
rect 1214 1095 1220 1096
rect 1214 1091 1215 1095
rect 1219 1091 1220 1095
rect 1214 1090 1220 1091
rect 1390 1095 1396 1096
rect 1390 1091 1391 1095
rect 1395 1091 1396 1095
rect 1390 1090 1396 1091
rect 210 1087 216 1088
rect 210 1083 211 1087
rect 215 1083 216 1087
rect 210 1082 216 1083
rect 314 1087 320 1088
rect 314 1083 315 1087
rect 319 1083 320 1087
rect 314 1082 320 1083
rect 450 1087 456 1088
rect 450 1083 451 1087
rect 455 1083 456 1087
rect 450 1082 456 1083
rect 602 1087 608 1088
rect 602 1083 603 1087
rect 607 1083 608 1087
rect 602 1082 608 1083
rect 618 1087 624 1088
rect 618 1083 619 1087
rect 623 1083 624 1087
rect 946 1087 952 1088
rect 618 1082 624 1083
rect 938 1083 944 1084
rect 938 1079 939 1083
rect 943 1079 944 1083
rect 946 1083 947 1087
rect 951 1083 952 1087
rect 946 1082 952 1083
rect 938 1078 944 1079
rect 238 1076 244 1077
rect 238 1072 239 1076
rect 243 1072 244 1076
rect 238 1071 244 1072
rect 374 1076 380 1077
rect 374 1072 375 1076
rect 379 1072 380 1076
rect 374 1071 380 1072
rect 526 1076 532 1077
rect 526 1072 527 1076
rect 531 1072 532 1076
rect 526 1071 532 1072
rect 694 1076 700 1077
rect 694 1072 695 1076
rect 699 1072 700 1076
rect 694 1071 700 1072
rect 862 1076 868 1077
rect 862 1072 863 1076
rect 867 1072 868 1076
rect 862 1071 868 1072
rect 240 1047 242 1071
rect 376 1047 378 1071
rect 528 1047 530 1071
rect 696 1047 698 1071
rect 864 1047 866 1071
rect 239 1046 243 1047
rect 239 1041 243 1042
rect 287 1046 291 1047
rect 287 1041 291 1042
rect 375 1046 379 1047
rect 375 1041 379 1042
rect 471 1046 475 1047
rect 471 1041 475 1042
rect 527 1046 531 1047
rect 527 1041 531 1042
rect 655 1046 659 1047
rect 655 1041 659 1042
rect 695 1046 699 1047
rect 695 1041 699 1042
rect 839 1046 843 1047
rect 839 1041 843 1042
rect 863 1046 867 1047
rect 863 1041 867 1042
rect 202 1023 208 1024
rect 202 1019 203 1023
rect 207 1019 208 1023
rect 202 1018 208 1019
rect 288 1017 290 1041
rect 472 1017 474 1041
rect 656 1017 658 1041
rect 840 1017 842 1041
rect 134 1016 140 1017
rect 110 1013 116 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 134 1012 135 1016
rect 139 1012 140 1016
rect 134 1011 140 1012
rect 286 1016 292 1017
rect 286 1012 287 1016
rect 291 1012 292 1016
rect 286 1011 292 1012
rect 470 1016 476 1017
rect 470 1012 471 1016
rect 475 1012 476 1016
rect 470 1011 476 1012
rect 654 1016 660 1017
rect 654 1012 655 1016
rect 659 1012 660 1016
rect 654 1011 660 1012
rect 838 1016 844 1017
rect 838 1012 839 1016
rect 843 1012 844 1016
rect 838 1011 844 1012
rect 110 1008 116 1009
rect 222 1007 228 1008
rect 222 1003 223 1007
rect 227 1003 228 1007
rect 222 1002 228 1003
rect 362 1007 368 1008
rect 362 1003 363 1007
rect 367 1003 368 1007
rect 362 1002 368 1003
rect 546 1007 552 1008
rect 546 1003 547 1007
rect 551 1003 552 1007
rect 546 1002 552 1003
rect 134 997 140 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 134 993 135 997
rect 139 993 140 997
rect 134 992 140 993
rect 110 991 116 992
rect 112 967 114 991
rect 136 967 138 992
rect 224 976 226 1002
rect 286 997 292 998
rect 286 993 287 997
rect 291 993 292 997
rect 286 992 292 993
rect 210 975 216 976
rect 210 971 211 975
rect 215 971 216 975
rect 210 970 216 971
rect 222 975 228 976
rect 222 971 223 975
rect 227 971 228 975
rect 222 970 228 971
rect 111 966 115 967
rect 111 961 115 962
rect 135 966 139 967
rect 135 961 139 962
rect 112 941 114 961
rect 110 940 116 941
rect 136 940 138 961
rect 110 936 111 940
rect 115 936 116 940
rect 110 935 116 936
rect 134 939 140 940
rect 134 935 135 939
rect 139 935 140 939
rect 134 934 140 935
rect 212 932 214 970
rect 288 967 290 992
rect 364 976 366 1002
rect 470 997 476 998
rect 470 993 471 997
rect 475 993 476 997
rect 470 992 476 993
rect 362 975 368 976
rect 362 971 363 975
rect 367 971 368 975
rect 362 970 368 971
rect 472 967 474 992
rect 548 976 550 1002
rect 654 997 660 998
rect 654 993 655 997
rect 659 993 660 997
rect 654 992 660 993
rect 838 997 844 998
rect 838 993 839 997
rect 843 993 844 997
rect 838 992 844 993
rect 546 975 552 976
rect 546 971 547 975
rect 551 971 552 975
rect 546 970 552 971
rect 656 967 658 992
rect 840 967 842 992
rect 940 976 942 1078
rect 1038 1076 1044 1077
rect 1038 1072 1039 1076
rect 1043 1072 1044 1076
rect 1038 1071 1044 1072
rect 1214 1076 1220 1077
rect 1214 1072 1215 1076
rect 1219 1072 1220 1076
rect 1214 1071 1220 1072
rect 1390 1076 1396 1077
rect 1390 1072 1391 1076
rect 1395 1072 1396 1076
rect 1390 1071 1396 1072
rect 1040 1047 1042 1071
rect 1216 1047 1218 1071
rect 1392 1047 1394 1071
rect 1015 1046 1019 1047
rect 1015 1041 1019 1042
rect 1039 1046 1043 1047
rect 1039 1041 1043 1042
rect 1199 1046 1203 1047
rect 1199 1041 1203 1042
rect 1215 1046 1219 1047
rect 1215 1041 1219 1042
rect 1383 1046 1387 1047
rect 1383 1041 1387 1042
rect 1391 1046 1395 1047
rect 1391 1041 1395 1042
rect 1016 1017 1018 1041
rect 1200 1017 1202 1041
rect 1384 1017 1386 1041
rect 1014 1016 1020 1017
rect 1014 1012 1015 1016
rect 1019 1012 1020 1016
rect 1014 1011 1020 1012
rect 1198 1016 1204 1017
rect 1198 1012 1199 1016
rect 1203 1012 1204 1016
rect 1198 1011 1204 1012
rect 1382 1016 1388 1017
rect 1382 1012 1383 1016
rect 1387 1012 1388 1016
rect 1382 1011 1388 1012
rect 1456 1008 1458 1110
rect 1468 1088 1470 1110
rect 1568 1096 1570 1117
rect 1744 1096 1746 1117
rect 1818 1107 1824 1108
rect 1818 1103 1819 1107
rect 1823 1103 1824 1107
rect 1818 1102 1824 1103
rect 1566 1095 1572 1096
rect 1566 1091 1567 1095
rect 1571 1091 1572 1095
rect 1566 1090 1572 1091
rect 1742 1095 1748 1096
rect 1742 1091 1743 1095
rect 1747 1091 1748 1095
rect 1742 1090 1748 1091
rect 1820 1088 1822 1102
rect 1904 1096 1906 1117
rect 2008 1097 2010 1117
rect 2276 1116 2278 1138
rect 2352 1124 2354 1145
rect 2482 1143 2488 1144
rect 2482 1139 2483 1143
rect 2487 1139 2488 1143
rect 2482 1138 2488 1139
rect 2350 1123 2356 1124
rect 2350 1119 2351 1123
rect 2355 1119 2356 1123
rect 2350 1118 2356 1119
rect 2484 1116 2486 1138
rect 2490 1135 2496 1136
rect 2490 1131 2491 1135
rect 2495 1131 2496 1135
rect 2490 1130 2496 1131
rect 2492 1116 2494 1130
rect 2512 1124 2514 1145
rect 2680 1124 2682 1145
rect 2780 1144 2782 1186
rect 2796 1160 2798 1186
rect 2886 1181 2892 1182
rect 2886 1177 2887 1181
rect 2891 1177 2892 1181
rect 2886 1176 2892 1177
rect 2794 1159 2800 1160
rect 2794 1155 2795 1159
rect 2799 1155 2800 1159
rect 2794 1154 2800 1155
rect 2888 1151 2890 1176
rect 2972 1160 2974 1186
rect 3086 1181 3092 1182
rect 3086 1177 3087 1181
rect 3091 1177 3092 1181
rect 3086 1176 3092 1177
rect 2970 1159 2976 1160
rect 2970 1155 2971 1159
rect 2975 1155 2976 1159
rect 2970 1154 2976 1155
rect 3088 1151 3090 1176
rect 3172 1160 3174 1186
rect 3310 1181 3316 1182
rect 3310 1177 3311 1181
rect 3315 1177 3316 1181
rect 3310 1176 3316 1177
rect 3170 1159 3176 1160
rect 3170 1155 3171 1159
rect 3175 1155 3176 1159
rect 3170 1154 3176 1155
rect 3312 1151 3314 1176
rect 3396 1160 3398 1186
rect 3542 1181 3548 1182
rect 3542 1177 3543 1181
rect 3547 1177 3548 1181
rect 3542 1176 3548 1177
rect 3394 1159 3400 1160
rect 3394 1155 3395 1159
rect 3399 1155 3400 1159
rect 3394 1154 3400 1155
rect 3544 1151 3546 1176
rect 3612 1160 3614 1270
rect 3942 1267 3948 1268
rect 3662 1264 3668 1265
rect 3662 1260 3663 1264
rect 3667 1260 3668 1264
rect 3662 1259 3668 1260
rect 3838 1264 3844 1265
rect 3838 1260 3839 1264
rect 3843 1260 3844 1264
rect 3942 1263 3943 1267
rect 3947 1263 3948 1267
rect 3942 1262 3948 1263
rect 3838 1259 3844 1260
rect 3664 1231 3666 1259
rect 3840 1231 3842 1259
rect 3944 1231 3946 1262
rect 3663 1230 3667 1231
rect 3663 1225 3667 1226
rect 3783 1230 3787 1231
rect 3783 1225 3787 1226
rect 3839 1230 3843 1231
rect 3839 1225 3843 1226
rect 3943 1230 3947 1231
rect 3943 1225 3947 1226
rect 3784 1201 3786 1225
rect 3782 1200 3788 1201
rect 3782 1196 3783 1200
rect 3787 1196 3788 1200
rect 3944 1198 3946 1225
rect 3782 1195 3788 1196
rect 3942 1197 3948 1198
rect 3942 1193 3943 1197
rect 3947 1193 3948 1197
rect 3942 1192 3948 1193
rect 3858 1191 3864 1192
rect 3858 1187 3859 1191
rect 3863 1187 3864 1191
rect 3858 1186 3864 1187
rect 3782 1181 3788 1182
rect 3782 1177 3783 1181
rect 3787 1177 3788 1181
rect 3782 1176 3788 1177
rect 3610 1159 3616 1160
rect 3610 1155 3611 1159
rect 3615 1155 3616 1159
rect 3610 1154 3616 1155
rect 3754 1159 3760 1160
rect 3754 1155 3755 1159
rect 3759 1155 3760 1159
rect 3754 1154 3760 1155
rect 2871 1150 2875 1151
rect 2871 1145 2875 1146
rect 2887 1150 2891 1151
rect 2887 1145 2891 1146
rect 3087 1150 3091 1151
rect 3087 1145 3091 1146
rect 3311 1150 3315 1151
rect 3311 1145 3315 1146
rect 3319 1150 3323 1151
rect 3319 1145 3323 1146
rect 3543 1150 3547 1151
rect 3543 1145 3547 1146
rect 3559 1150 3563 1151
rect 3559 1145 3563 1146
rect 2778 1143 2784 1144
rect 2778 1139 2779 1143
rect 2783 1139 2784 1143
rect 2778 1138 2784 1139
rect 2786 1143 2792 1144
rect 2786 1139 2787 1143
rect 2791 1139 2792 1143
rect 2786 1138 2792 1139
rect 2510 1123 2516 1124
rect 2510 1119 2511 1123
rect 2515 1119 2516 1123
rect 2510 1118 2516 1119
rect 2678 1123 2684 1124
rect 2678 1119 2679 1123
rect 2683 1119 2684 1123
rect 2678 1118 2684 1119
rect 2788 1116 2790 1138
rect 2872 1124 2874 1145
rect 2946 1143 2952 1144
rect 2946 1139 2947 1143
rect 2951 1139 2952 1143
rect 2946 1138 2952 1139
rect 2870 1123 2876 1124
rect 2870 1119 2871 1123
rect 2875 1119 2876 1123
rect 2870 1118 2876 1119
rect 2948 1116 2950 1138
rect 3088 1124 3090 1145
rect 3162 1143 3168 1144
rect 3162 1139 3163 1143
rect 3167 1139 3168 1143
rect 3162 1138 3168 1139
rect 3086 1123 3092 1124
rect 3086 1119 3087 1123
rect 3091 1119 3092 1123
rect 3086 1118 3092 1119
rect 3164 1116 3166 1138
rect 3320 1124 3322 1145
rect 3394 1143 3400 1144
rect 3394 1139 3395 1143
rect 3399 1139 3400 1143
rect 3394 1138 3400 1139
rect 3318 1123 3324 1124
rect 3318 1119 3319 1123
rect 3323 1119 3324 1123
rect 3318 1118 3324 1119
rect 3396 1116 3398 1138
rect 3560 1124 3562 1145
rect 3558 1123 3564 1124
rect 3558 1119 3559 1123
rect 3563 1119 3564 1123
rect 3558 1118 3564 1119
rect 2274 1115 2280 1116
rect 2274 1111 2275 1115
rect 2279 1111 2280 1115
rect 2274 1110 2280 1111
rect 2482 1115 2488 1116
rect 2482 1111 2483 1115
rect 2487 1111 2488 1115
rect 2482 1110 2488 1111
rect 2490 1115 2496 1116
rect 2490 1111 2491 1115
rect 2495 1111 2496 1115
rect 2490 1110 2496 1111
rect 2786 1115 2792 1116
rect 2786 1111 2787 1115
rect 2791 1111 2792 1115
rect 2786 1110 2792 1111
rect 2946 1115 2952 1116
rect 2946 1111 2947 1115
rect 2951 1111 2952 1115
rect 2946 1110 2952 1111
rect 3162 1115 3168 1116
rect 3162 1111 3163 1115
rect 3167 1111 3168 1115
rect 3162 1110 3168 1111
rect 3394 1115 3400 1116
rect 3394 1111 3395 1115
rect 3399 1111 3400 1115
rect 3394 1110 3400 1111
rect 3402 1115 3408 1116
rect 3402 1111 3403 1115
rect 3407 1111 3408 1115
rect 3402 1110 3408 1111
rect 2046 1107 2052 1108
rect 2046 1103 2047 1107
rect 2051 1103 2052 1107
rect 2046 1102 2052 1103
rect 2070 1104 2076 1105
rect 2006 1096 2012 1097
rect 1902 1095 1908 1096
rect 1902 1091 1903 1095
rect 1907 1091 1908 1095
rect 2006 1092 2007 1096
rect 2011 1092 2012 1096
rect 2006 1091 2012 1092
rect 1902 1090 1908 1091
rect 1466 1087 1472 1088
rect 1466 1083 1467 1087
rect 1471 1083 1472 1087
rect 1466 1082 1472 1083
rect 1818 1087 1824 1088
rect 1818 1083 1819 1087
rect 1823 1083 1824 1087
rect 1818 1082 1824 1083
rect 2006 1079 2012 1080
rect 1566 1076 1572 1077
rect 1566 1072 1567 1076
rect 1571 1072 1572 1076
rect 1566 1071 1572 1072
rect 1742 1076 1748 1077
rect 1742 1072 1743 1076
rect 1747 1072 1748 1076
rect 1742 1071 1748 1072
rect 1902 1076 1908 1077
rect 1902 1072 1903 1076
rect 1907 1072 1908 1076
rect 2006 1075 2007 1079
rect 2011 1075 2012 1079
rect 2006 1074 2012 1075
rect 1902 1071 1908 1072
rect 1568 1047 1570 1071
rect 1744 1047 1746 1071
rect 1904 1047 1906 1071
rect 2008 1047 2010 1074
rect 2048 1063 2050 1102
rect 2070 1100 2071 1104
rect 2075 1100 2076 1104
rect 2070 1099 2076 1100
rect 2198 1104 2204 1105
rect 2198 1100 2199 1104
rect 2203 1100 2204 1104
rect 2198 1099 2204 1100
rect 2350 1104 2356 1105
rect 2350 1100 2351 1104
rect 2355 1100 2356 1104
rect 2350 1099 2356 1100
rect 2510 1104 2516 1105
rect 2510 1100 2511 1104
rect 2515 1100 2516 1104
rect 2510 1099 2516 1100
rect 2678 1104 2684 1105
rect 2678 1100 2679 1104
rect 2683 1100 2684 1104
rect 2678 1099 2684 1100
rect 2870 1104 2876 1105
rect 2870 1100 2871 1104
rect 2875 1100 2876 1104
rect 2870 1099 2876 1100
rect 3086 1104 3092 1105
rect 3086 1100 3087 1104
rect 3091 1100 3092 1104
rect 3086 1099 3092 1100
rect 3318 1104 3324 1105
rect 3318 1100 3319 1104
rect 3323 1100 3324 1104
rect 3318 1099 3324 1100
rect 2072 1063 2074 1099
rect 2134 1087 2140 1088
rect 2134 1083 2135 1087
rect 2139 1083 2140 1087
rect 2134 1082 2140 1083
rect 2047 1062 2051 1063
rect 2047 1057 2051 1058
rect 2071 1062 2075 1063
rect 2071 1057 2075 1058
rect 1567 1046 1571 1047
rect 1567 1041 1571 1042
rect 1743 1046 1747 1047
rect 1743 1041 1747 1042
rect 1903 1046 1907 1047
rect 1903 1041 1907 1042
rect 2007 1046 2011 1047
rect 2007 1041 2011 1042
rect 1568 1017 1570 1041
rect 1566 1016 1572 1017
rect 1566 1012 1567 1016
rect 1571 1012 1572 1016
rect 2008 1014 2010 1041
rect 2048 1030 2050 1057
rect 2072 1033 2074 1057
rect 2070 1032 2076 1033
rect 2046 1029 2052 1030
rect 2046 1025 2047 1029
rect 2051 1025 2052 1029
rect 2070 1028 2071 1032
rect 2075 1028 2076 1032
rect 2070 1027 2076 1028
rect 2046 1024 2052 1025
rect 1566 1011 1572 1012
rect 2006 1013 2012 1014
rect 2070 1013 2076 1014
rect 2006 1009 2007 1013
rect 2011 1009 2012 1013
rect 2006 1008 2012 1009
rect 2046 1012 2052 1013
rect 2046 1008 2047 1012
rect 2051 1008 2052 1012
rect 2070 1009 2071 1013
rect 2075 1009 2076 1013
rect 2070 1008 2076 1009
rect 978 1007 984 1008
rect 978 1003 979 1007
rect 983 1003 984 1007
rect 978 1002 984 1003
rect 1006 1007 1012 1008
rect 1006 1003 1007 1007
rect 1011 1003 1012 1007
rect 1006 1002 1012 1003
rect 1274 1007 1280 1008
rect 1274 1003 1275 1007
rect 1279 1003 1280 1007
rect 1274 1002 1280 1003
rect 1454 1007 1460 1008
rect 1454 1003 1455 1007
rect 1459 1003 1460 1007
rect 1454 1002 1460 1003
rect 1466 1007 1472 1008
rect 2046 1007 2052 1008
rect 1466 1003 1467 1007
rect 1471 1003 1472 1007
rect 1466 1002 1472 1003
rect 980 976 982 1002
rect 938 975 944 976
rect 938 971 939 975
rect 943 971 944 975
rect 938 970 944 971
rect 978 975 984 976
rect 978 971 979 975
rect 983 971 984 975
rect 978 970 984 971
rect 287 966 291 967
rect 287 961 291 962
rect 295 966 299 967
rect 295 961 299 962
rect 471 966 475 967
rect 471 961 475 962
rect 639 966 643 967
rect 639 961 643 962
rect 655 966 659 967
rect 655 961 659 962
rect 799 966 803 967
rect 799 961 803 962
rect 839 966 843 967
rect 839 961 843 962
rect 951 966 955 967
rect 951 961 955 962
rect 270 959 276 960
rect 270 955 271 959
rect 275 955 276 959
rect 270 954 276 955
rect 272 932 274 954
rect 296 940 298 961
rect 430 959 436 960
rect 430 955 431 959
rect 435 955 436 959
rect 430 954 436 955
rect 294 939 300 940
rect 294 935 295 939
rect 299 935 300 939
rect 294 934 300 935
rect 210 931 216 932
rect 210 927 211 931
rect 215 927 216 931
rect 210 926 216 927
rect 270 931 276 932
rect 270 927 271 931
rect 275 927 276 931
rect 270 926 276 927
rect 110 923 116 924
rect 110 919 111 923
rect 115 919 116 923
rect 110 918 116 919
rect 134 920 140 921
rect 112 891 114 918
rect 134 916 135 920
rect 139 916 140 920
rect 134 915 140 916
rect 294 920 300 921
rect 294 916 295 920
rect 299 916 300 920
rect 294 915 300 916
rect 136 891 138 915
rect 296 891 298 915
rect 111 890 115 891
rect 111 885 115 886
rect 135 890 139 891
rect 135 885 139 886
rect 159 890 163 891
rect 159 885 163 886
rect 295 890 299 891
rect 295 885 299 886
rect 319 890 323 891
rect 319 885 323 886
rect 112 858 114 885
rect 160 861 162 885
rect 320 861 322 885
rect 158 860 164 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 158 856 159 860
rect 163 856 164 860
rect 158 855 164 856
rect 318 860 324 861
rect 318 856 319 860
rect 323 856 324 860
rect 318 855 324 856
rect 110 852 116 853
rect 432 852 434 954
rect 472 940 474 961
rect 640 940 642 961
rect 800 940 802 961
rect 882 959 888 960
rect 882 955 883 959
rect 887 955 888 959
rect 882 954 888 955
rect 470 939 476 940
rect 470 935 471 939
rect 475 935 476 939
rect 470 934 476 935
rect 638 939 644 940
rect 638 935 639 939
rect 643 935 644 939
rect 638 934 644 935
rect 798 939 804 940
rect 798 935 799 939
rect 803 935 804 939
rect 798 934 804 935
rect 884 932 886 954
rect 952 940 954 961
rect 1008 960 1010 1002
rect 1014 997 1020 998
rect 1014 993 1015 997
rect 1019 993 1020 997
rect 1014 992 1020 993
rect 1198 997 1204 998
rect 1198 993 1199 997
rect 1203 993 1204 997
rect 1198 992 1204 993
rect 1016 967 1018 992
rect 1200 967 1202 992
rect 1276 976 1278 1002
rect 1382 997 1388 998
rect 1382 993 1383 997
rect 1387 993 1388 997
rect 1382 992 1388 993
rect 1274 975 1280 976
rect 1274 971 1275 975
rect 1279 971 1280 975
rect 1274 970 1280 971
rect 1384 967 1386 992
rect 1468 984 1470 1002
rect 1566 997 1572 998
rect 1566 993 1567 997
rect 1571 993 1572 997
rect 1566 992 1572 993
rect 2006 996 2012 997
rect 2006 992 2007 996
rect 2011 992 2012 996
rect 1466 983 1472 984
rect 1466 979 1467 983
rect 1471 979 1472 983
rect 1466 978 1472 979
rect 1568 967 1570 992
rect 2006 991 2012 992
rect 1582 975 1588 976
rect 1582 971 1583 975
rect 1587 971 1588 975
rect 1582 970 1588 971
rect 1015 966 1019 967
rect 1015 961 1019 962
rect 1087 966 1091 967
rect 1087 961 1091 962
rect 1199 966 1203 967
rect 1199 961 1203 962
rect 1223 966 1227 967
rect 1223 961 1227 962
rect 1359 966 1363 967
rect 1359 961 1363 962
rect 1383 966 1387 967
rect 1383 961 1387 962
rect 1495 966 1499 967
rect 1495 961 1499 962
rect 1567 966 1571 967
rect 1567 961 1571 962
rect 1006 959 1012 960
rect 1006 955 1007 959
rect 1011 955 1012 959
rect 1006 954 1012 955
rect 1088 940 1090 961
rect 1162 959 1168 960
rect 1162 955 1163 959
rect 1167 955 1168 959
rect 1162 954 1168 955
rect 950 939 956 940
rect 950 935 951 939
rect 955 935 956 939
rect 950 934 956 935
rect 1086 939 1092 940
rect 1086 935 1087 939
rect 1091 935 1092 939
rect 1086 934 1092 935
rect 1164 932 1166 954
rect 1224 940 1226 961
rect 1298 959 1304 960
rect 1298 955 1299 959
rect 1303 955 1304 959
rect 1298 954 1304 955
rect 1222 939 1228 940
rect 1222 935 1223 939
rect 1227 935 1228 939
rect 1222 934 1228 935
rect 1300 932 1302 954
rect 1314 951 1320 952
rect 1314 947 1315 951
rect 1319 947 1320 951
rect 1314 946 1320 947
rect 882 931 888 932
rect 714 927 720 928
rect 714 923 715 927
rect 719 923 720 927
rect 882 927 883 931
rect 887 927 888 931
rect 882 926 888 927
rect 1162 931 1168 932
rect 1162 927 1163 931
rect 1167 927 1168 931
rect 1162 926 1168 927
rect 1298 931 1304 932
rect 1298 927 1299 931
rect 1303 927 1304 931
rect 1298 926 1304 927
rect 714 922 720 923
rect 470 920 476 921
rect 470 916 471 920
rect 475 916 476 920
rect 470 915 476 916
rect 638 920 644 921
rect 638 916 639 920
rect 643 916 644 920
rect 638 915 644 916
rect 472 891 474 915
rect 640 891 642 915
rect 471 890 475 891
rect 471 885 475 886
rect 615 890 619 891
rect 615 885 619 886
rect 639 890 643 891
rect 639 885 643 886
rect 472 861 474 885
rect 616 861 618 885
rect 470 860 476 861
rect 470 856 471 860
rect 475 856 476 860
rect 470 855 476 856
rect 614 860 620 861
rect 614 856 615 860
rect 619 856 620 860
rect 614 855 620 856
rect 234 851 240 852
rect 234 847 235 851
rect 239 847 240 851
rect 234 846 240 847
rect 430 851 436 852
rect 430 847 431 851
rect 435 847 436 851
rect 430 846 436 847
rect 546 851 552 852
rect 546 847 547 851
rect 551 847 552 851
rect 546 846 552 847
rect 554 851 560 852
rect 554 847 555 851
rect 559 847 560 851
rect 554 846 560 847
rect 698 851 704 852
rect 698 847 699 851
rect 703 847 704 851
rect 698 846 704 847
rect 158 841 164 842
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 158 837 159 841
rect 163 837 164 841
rect 158 836 164 837
rect 110 835 116 836
rect 112 815 114 835
rect 160 815 162 836
rect 236 820 238 846
rect 318 841 324 842
rect 318 837 319 841
rect 323 837 324 841
rect 318 836 324 837
rect 470 841 476 842
rect 470 837 471 841
rect 475 837 476 841
rect 470 836 476 837
rect 214 819 220 820
rect 214 815 215 819
rect 219 815 220 819
rect 234 819 240 820
rect 234 815 235 819
rect 239 815 240 819
rect 320 815 322 836
rect 472 815 474 836
rect 111 814 115 815
rect 111 809 115 810
rect 159 814 163 815
rect 214 814 220 815
rect 223 814 227 815
rect 234 814 240 815
rect 319 814 323 815
rect 159 809 163 810
rect 112 789 114 809
rect 110 788 116 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 216 780 218 814
rect 223 809 227 810
rect 319 809 323 810
rect 383 814 387 815
rect 383 809 387 810
rect 471 814 475 815
rect 471 809 475 810
rect 535 814 539 815
rect 535 809 539 810
rect 224 788 226 809
rect 306 807 312 808
rect 306 803 307 807
rect 311 803 312 807
rect 306 802 312 803
rect 222 787 228 788
rect 222 783 223 787
rect 227 783 228 787
rect 222 782 228 783
rect 308 780 310 802
rect 384 788 386 809
rect 402 807 408 808
rect 402 803 403 807
rect 407 803 408 807
rect 402 802 408 803
rect 382 787 388 788
rect 382 783 383 787
rect 387 783 388 787
rect 382 782 388 783
rect 214 779 220 780
rect 214 775 215 779
rect 219 775 220 779
rect 214 774 220 775
rect 306 779 312 780
rect 306 775 307 779
rect 311 775 312 779
rect 306 774 312 775
rect 110 771 116 772
rect 110 767 111 771
rect 115 767 116 771
rect 110 766 116 767
rect 222 768 228 769
rect 112 735 114 766
rect 222 764 223 768
rect 227 764 228 768
rect 222 763 228 764
rect 382 768 388 769
rect 382 764 383 768
rect 387 764 388 768
rect 382 763 388 764
rect 224 735 226 763
rect 384 735 386 763
rect 111 734 115 735
rect 111 729 115 730
rect 223 734 227 735
rect 223 729 227 730
rect 311 734 315 735
rect 311 729 315 730
rect 383 734 387 735
rect 383 729 387 730
rect 112 702 114 729
rect 312 705 314 729
rect 310 704 316 705
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 310 700 311 704
rect 315 700 316 704
rect 310 699 316 700
rect 110 696 116 697
rect 404 696 406 802
rect 536 788 538 809
rect 548 808 550 846
rect 556 820 558 846
rect 614 841 620 842
rect 614 837 615 841
rect 619 837 620 841
rect 614 836 620 837
rect 554 819 560 820
rect 554 815 555 819
rect 559 815 560 819
rect 616 815 618 836
rect 700 820 702 846
rect 716 820 718 922
rect 798 920 804 921
rect 798 916 799 920
rect 803 916 804 920
rect 798 915 804 916
rect 950 920 956 921
rect 950 916 951 920
rect 955 916 956 920
rect 950 915 956 916
rect 1086 920 1092 921
rect 1086 916 1087 920
rect 1091 916 1092 920
rect 1086 915 1092 916
rect 1222 920 1228 921
rect 1222 916 1223 920
rect 1227 916 1228 920
rect 1222 915 1228 916
rect 800 891 802 915
rect 952 891 954 915
rect 1088 891 1090 915
rect 1224 891 1226 915
rect 751 890 755 891
rect 751 885 755 886
rect 799 890 803 891
rect 799 885 803 886
rect 879 890 883 891
rect 879 885 883 886
rect 951 890 955 891
rect 951 885 955 886
rect 999 890 1003 891
rect 999 885 1003 886
rect 1087 890 1091 891
rect 1087 885 1091 886
rect 1111 890 1115 891
rect 1111 885 1115 886
rect 1223 890 1227 891
rect 1223 885 1227 886
rect 1231 890 1235 891
rect 1231 885 1235 886
rect 752 861 754 885
rect 880 861 882 885
rect 1000 861 1002 885
rect 1112 861 1114 885
rect 1232 861 1234 885
rect 750 860 756 861
rect 750 856 751 860
rect 755 856 756 860
rect 750 855 756 856
rect 878 860 884 861
rect 878 856 879 860
rect 883 856 884 860
rect 878 855 884 856
rect 998 860 1004 861
rect 998 856 999 860
rect 1003 856 1004 860
rect 998 855 1004 856
rect 1110 860 1116 861
rect 1110 856 1111 860
rect 1115 856 1116 860
rect 1110 855 1116 856
rect 1230 860 1236 861
rect 1230 856 1231 860
rect 1235 856 1236 860
rect 1230 855 1236 856
rect 1316 852 1318 946
rect 1360 940 1362 961
rect 1434 959 1440 960
rect 1434 955 1435 959
rect 1439 955 1440 959
rect 1434 954 1440 955
rect 1358 939 1364 940
rect 1358 935 1359 939
rect 1363 935 1364 939
rect 1358 934 1364 935
rect 1436 932 1438 954
rect 1496 940 1498 961
rect 1494 939 1500 940
rect 1494 935 1495 939
rect 1499 935 1500 939
rect 1494 934 1500 935
rect 1584 932 1586 970
rect 2008 967 2010 991
rect 2048 983 2050 1007
rect 2072 983 2074 1008
rect 2136 992 2138 1082
rect 2200 1063 2202 1099
rect 2352 1063 2354 1099
rect 2512 1063 2514 1099
rect 2680 1063 2682 1099
rect 2872 1063 2874 1099
rect 3088 1063 3090 1099
rect 3320 1063 3322 1099
rect 2199 1062 2203 1063
rect 2199 1057 2203 1058
rect 2263 1062 2267 1063
rect 2263 1057 2267 1058
rect 2351 1062 2355 1063
rect 2351 1057 2355 1058
rect 2487 1062 2491 1063
rect 2487 1057 2491 1058
rect 2511 1062 2515 1063
rect 2511 1057 2515 1058
rect 2679 1062 2683 1063
rect 2679 1057 2683 1058
rect 2703 1062 2707 1063
rect 2703 1057 2707 1058
rect 2871 1062 2875 1063
rect 2871 1057 2875 1058
rect 2919 1062 2923 1063
rect 2919 1057 2923 1058
rect 3087 1062 3091 1063
rect 3087 1057 3091 1058
rect 3119 1062 3123 1063
rect 3119 1057 3123 1058
rect 3311 1062 3315 1063
rect 3311 1057 3315 1058
rect 3319 1062 3323 1063
rect 3319 1057 3323 1058
rect 2264 1033 2266 1057
rect 2488 1033 2490 1057
rect 2704 1033 2706 1057
rect 2920 1033 2922 1057
rect 3120 1033 3122 1057
rect 3312 1033 3314 1057
rect 2262 1032 2268 1033
rect 2262 1028 2263 1032
rect 2267 1028 2268 1032
rect 2262 1027 2268 1028
rect 2486 1032 2492 1033
rect 2486 1028 2487 1032
rect 2491 1028 2492 1032
rect 2486 1027 2492 1028
rect 2702 1032 2708 1033
rect 2702 1028 2703 1032
rect 2707 1028 2708 1032
rect 2702 1027 2708 1028
rect 2918 1032 2924 1033
rect 2918 1028 2919 1032
rect 2923 1028 2924 1032
rect 2918 1027 2924 1028
rect 3118 1032 3124 1033
rect 3118 1028 3119 1032
rect 3123 1028 3124 1032
rect 3118 1027 3124 1028
rect 3310 1032 3316 1033
rect 3310 1028 3311 1032
rect 3315 1028 3316 1032
rect 3310 1027 3316 1028
rect 2146 1023 2152 1024
rect 2146 1019 2147 1023
rect 2151 1019 2152 1023
rect 2146 1018 2152 1019
rect 2338 1023 2344 1024
rect 2338 1019 2339 1023
rect 2343 1019 2344 1023
rect 2338 1018 2344 1019
rect 2562 1023 2568 1024
rect 2562 1019 2563 1023
rect 2567 1019 2568 1023
rect 2562 1018 2568 1019
rect 2570 1023 2576 1024
rect 2570 1019 2571 1023
rect 2575 1019 2576 1023
rect 2570 1018 2576 1019
rect 3002 1023 3008 1024
rect 3002 1019 3003 1023
rect 3007 1019 3008 1023
rect 3002 1018 3008 1019
rect 3202 1023 3208 1024
rect 3202 1019 3203 1023
rect 3207 1019 3208 1023
rect 3202 1018 3208 1019
rect 2148 992 2150 1018
rect 2262 1013 2268 1014
rect 2262 1009 2263 1013
rect 2267 1009 2268 1013
rect 2262 1008 2268 1009
rect 2134 991 2140 992
rect 2134 987 2135 991
rect 2139 987 2140 991
rect 2134 986 2140 987
rect 2146 991 2152 992
rect 2146 987 2147 991
rect 2151 987 2152 991
rect 2146 986 2152 987
rect 2264 983 2266 1008
rect 2340 992 2342 1018
rect 2486 1013 2492 1014
rect 2486 1009 2487 1013
rect 2491 1009 2492 1013
rect 2486 1008 2492 1009
rect 2338 991 2344 992
rect 2338 987 2339 991
rect 2343 987 2344 991
rect 2338 986 2344 987
rect 2488 983 2490 1008
rect 2564 992 2566 1018
rect 2562 991 2568 992
rect 2562 987 2563 991
rect 2567 987 2568 991
rect 2562 986 2568 987
rect 2572 984 2574 1018
rect 2702 1013 2708 1014
rect 2702 1009 2703 1013
rect 2707 1009 2708 1013
rect 2702 1008 2708 1009
rect 2918 1013 2924 1014
rect 2918 1009 2919 1013
rect 2923 1009 2924 1013
rect 2918 1008 2924 1009
rect 2570 983 2576 984
rect 2704 983 2706 1008
rect 2920 983 2922 1008
rect 3004 992 3006 1018
rect 3038 1015 3044 1016
rect 3038 1011 3039 1015
rect 3043 1011 3044 1015
rect 3038 1010 3044 1011
rect 3118 1013 3124 1014
rect 3002 991 3008 992
rect 3002 987 3003 991
rect 3007 987 3008 991
rect 3002 986 3008 987
rect 2047 982 2051 983
rect 2047 977 2051 978
rect 2071 982 2075 983
rect 2071 977 2075 978
rect 2263 982 2267 983
rect 2263 977 2267 978
rect 2303 982 2307 983
rect 2303 977 2307 978
rect 2455 982 2459 983
rect 2455 977 2459 978
rect 2487 982 2491 983
rect 2570 979 2571 983
rect 2575 979 2576 983
rect 2570 978 2576 979
rect 2615 982 2619 983
rect 2487 977 2491 978
rect 2615 977 2619 978
rect 2703 982 2707 983
rect 2703 977 2707 978
rect 2783 982 2787 983
rect 2783 977 2787 978
rect 2919 982 2923 983
rect 2919 977 2923 978
rect 2951 982 2955 983
rect 2951 977 2955 978
rect 2007 966 2011 967
rect 2007 961 2011 962
rect 2008 941 2010 961
rect 2048 957 2050 977
rect 2046 956 2052 957
rect 2304 956 2306 977
rect 2378 975 2384 976
rect 2378 971 2379 975
rect 2383 971 2384 975
rect 2378 970 2384 971
rect 2046 952 2047 956
rect 2051 952 2052 956
rect 2046 951 2052 952
rect 2302 955 2308 956
rect 2302 951 2303 955
rect 2307 951 2308 955
rect 2302 950 2308 951
rect 2380 948 2382 970
rect 2456 956 2458 977
rect 2530 975 2536 976
rect 2530 971 2531 975
rect 2535 971 2536 975
rect 2530 970 2536 971
rect 2454 955 2460 956
rect 2454 951 2455 955
rect 2459 951 2460 955
rect 2454 950 2460 951
rect 2532 948 2534 970
rect 2616 956 2618 977
rect 2690 975 2696 976
rect 2690 971 2691 975
rect 2695 971 2696 975
rect 2690 970 2696 971
rect 2614 955 2620 956
rect 2614 951 2615 955
rect 2619 951 2620 955
rect 2614 950 2620 951
rect 2692 948 2694 970
rect 2784 956 2786 977
rect 2858 975 2864 976
rect 2858 971 2859 975
rect 2863 971 2864 975
rect 2858 970 2864 971
rect 2782 955 2788 956
rect 2782 951 2783 955
rect 2787 951 2788 955
rect 2782 950 2788 951
rect 2860 948 2862 970
rect 2952 956 2954 977
rect 3040 976 3042 1010
rect 3118 1009 3119 1013
rect 3123 1009 3124 1013
rect 3118 1008 3124 1009
rect 3120 983 3122 1008
rect 3204 992 3206 1018
rect 3310 1013 3316 1014
rect 3310 1009 3311 1013
rect 3315 1009 3316 1013
rect 3310 1008 3316 1009
rect 3202 991 3208 992
rect 3202 987 3203 991
rect 3207 987 3208 991
rect 3202 986 3208 987
rect 3312 983 3314 1008
rect 3404 992 3406 1110
rect 3558 1104 3564 1105
rect 3558 1100 3559 1104
rect 3563 1100 3564 1104
rect 3558 1099 3564 1100
rect 3560 1063 3562 1099
rect 3495 1062 3499 1063
rect 3495 1057 3499 1058
rect 3559 1062 3563 1063
rect 3559 1057 3563 1058
rect 3679 1062 3683 1063
rect 3679 1057 3683 1058
rect 3496 1033 3498 1057
rect 3680 1033 3682 1057
rect 3494 1032 3500 1033
rect 3494 1028 3495 1032
rect 3499 1028 3500 1032
rect 3494 1027 3500 1028
rect 3678 1032 3684 1033
rect 3678 1028 3679 1032
rect 3683 1028 3684 1032
rect 3678 1027 3684 1028
rect 3756 1024 3758 1154
rect 3784 1151 3786 1176
rect 3783 1150 3787 1151
rect 3783 1145 3787 1146
rect 3807 1150 3811 1151
rect 3807 1145 3811 1146
rect 3808 1124 3810 1145
rect 3860 1144 3862 1186
rect 3942 1180 3948 1181
rect 3942 1176 3943 1180
rect 3947 1176 3948 1180
rect 3942 1175 3948 1176
rect 3944 1151 3946 1175
rect 3943 1150 3947 1151
rect 3943 1145 3947 1146
rect 3858 1143 3864 1144
rect 3858 1139 3859 1143
rect 3863 1139 3864 1143
rect 3858 1138 3864 1139
rect 3944 1125 3946 1145
rect 3942 1124 3948 1125
rect 3806 1123 3812 1124
rect 3806 1119 3807 1123
rect 3811 1119 3812 1123
rect 3942 1120 3943 1124
rect 3947 1120 3948 1124
rect 3942 1119 3948 1120
rect 3806 1118 3812 1119
rect 3882 1111 3888 1112
rect 3882 1107 3883 1111
rect 3887 1107 3888 1111
rect 3882 1106 3888 1107
rect 3942 1107 3948 1108
rect 3806 1104 3812 1105
rect 3806 1100 3807 1104
rect 3811 1100 3812 1104
rect 3806 1099 3812 1100
rect 3808 1063 3810 1099
rect 3807 1062 3811 1063
rect 3807 1057 3811 1058
rect 3839 1062 3843 1063
rect 3839 1057 3843 1058
rect 3840 1033 3842 1057
rect 3838 1032 3844 1033
rect 3838 1028 3839 1032
rect 3843 1028 3844 1032
rect 3838 1027 3844 1028
rect 3570 1023 3576 1024
rect 3570 1019 3571 1023
rect 3575 1019 3576 1023
rect 3570 1018 3576 1019
rect 3754 1023 3760 1024
rect 3754 1019 3755 1023
rect 3759 1019 3760 1023
rect 3754 1018 3760 1019
rect 3494 1013 3500 1014
rect 3494 1009 3495 1013
rect 3499 1009 3500 1013
rect 3494 1008 3500 1009
rect 3402 991 3408 992
rect 3402 987 3403 991
rect 3407 987 3408 991
rect 3402 986 3408 987
rect 3496 983 3498 1008
rect 3572 992 3574 1018
rect 3678 1013 3684 1014
rect 3678 1009 3679 1013
rect 3683 1009 3684 1013
rect 3678 1008 3684 1009
rect 3838 1013 3844 1014
rect 3838 1009 3839 1013
rect 3843 1009 3844 1013
rect 3838 1008 3844 1009
rect 3550 991 3556 992
rect 3550 987 3551 991
rect 3555 987 3556 991
rect 3550 986 3556 987
rect 3570 991 3576 992
rect 3570 987 3571 991
rect 3575 987 3576 991
rect 3570 986 3576 987
rect 3111 982 3115 983
rect 3111 977 3115 978
rect 3119 982 3123 983
rect 3119 977 3123 978
rect 3263 982 3267 983
rect 3263 977 3267 978
rect 3311 982 3315 983
rect 3311 977 3315 978
rect 3415 982 3419 983
rect 3415 977 3419 978
rect 3495 982 3499 983
rect 3495 977 3499 978
rect 3038 975 3044 976
rect 3038 971 3039 975
rect 3043 971 3044 975
rect 3038 970 3044 971
rect 3112 956 3114 977
rect 3186 975 3192 976
rect 3186 971 3187 975
rect 3191 971 3192 975
rect 3186 970 3192 971
rect 2950 955 2956 956
rect 2950 951 2951 955
rect 2955 951 2956 955
rect 2950 950 2956 951
rect 3110 955 3116 956
rect 3110 951 3111 955
rect 3115 951 3116 955
rect 3110 950 3116 951
rect 3188 948 3190 970
rect 3264 956 3266 977
rect 3338 975 3344 976
rect 3338 971 3339 975
rect 3343 971 3344 975
rect 3338 970 3344 971
rect 3262 955 3268 956
rect 3262 951 3263 955
rect 3267 951 3268 955
rect 3262 950 3268 951
rect 3340 948 3342 970
rect 3416 956 3418 977
rect 3538 975 3544 976
rect 3538 971 3539 975
rect 3543 971 3544 975
rect 3538 970 3544 971
rect 3414 955 3420 956
rect 3414 951 3415 955
rect 3419 951 3420 955
rect 3414 950 3420 951
rect 3540 948 3542 970
rect 3552 948 3554 986
rect 3680 983 3682 1008
rect 3840 983 3842 1008
rect 3884 992 3886 1106
rect 3942 1103 3943 1107
rect 3947 1103 3948 1107
rect 3942 1102 3948 1103
rect 3944 1063 3946 1102
rect 3943 1062 3947 1063
rect 3943 1057 3947 1058
rect 3944 1030 3946 1057
rect 3942 1029 3948 1030
rect 3942 1025 3943 1029
rect 3947 1025 3948 1029
rect 3942 1024 3948 1025
rect 3906 1023 3912 1024
rect 3906 1019 3907 1023
rect 3911 1019 3912 1023
rect 3906 1018 3912 1019
rect 3882 991 3888 992
rect 3882 987 3883 991
rect 3887 987 3888 991
rect 3882 986 3888 987
rect 3559 982 3563 983
rect 3559 977 3563 978
rect 3679 982 3683 983
rect 3679 977 3683 978
rect 3711 982 3715 983
rect 3711 977 3715 978
rect 3839 982 3843 983
rect 3839 977 3843 978
rect 3560 956 3562 977
rect 3712 956 3714 977
rect 3794 975 3800 976
rect 3794 971 3795 975
rect 3799 971 3800 975
rect 3794 970 3800 971
rect 3558 955 3564 956
rect 3558 951 3559 955
rect 3563 951 3564 955
rect 3558 950 3564 951
rect 3710 955 3716 956
rect 3710 951 3711 955
rect 3715 951 3716 955
rect 3710 950 3716 951
rect 2378 947 2384 948
rect 2378 943 2379 947
rect 2383 943 2384 947
rect 2378 942 2384 943
rect 2530 947 2536 948
rect 2530 943 2531 947
rect 2535 943 2536 947
rect 2530 942 2536 943
rect 2690 947 2696 948
rect 2690 943 2691 947
rect 2695 943 2696 947
rect 2690 942 2696 943
rect 2858 947 2864 948
rect 2858 943 2859 947
rect 2863 943 2864 947
rect 2858 942 2864 943
rect 2906 947 2912 948
rect 2906 943 2907 947
rect 2911 943 2912 947
rect 2906 942 2912 943
rect 3186 947 3192 948
rect 3186 943 3187 947
rect 3191 943 3192 947
rect 3186 942 3192 943
rect 3338 947 3344 948
rect 3338 943 3339 947
rect 3343 943 3344 947
rect 3338 942 3344 943
rect 3538 947 3544 948
rect 3538 943 3539 947
rect 3543 943 3544 947
rect 3538 942 3544 943
rect 3550 947 3556 948
rect 3550 943 3551 947
rect 3555 943 3556 947
rect 3550 942 3556 943
rect 3642 947 3648 948
rect 3642 943 3643 947
rect 3647 943 3648 947
rect 3642 942 3648 943
rect 2006 940 2012 941
rect 2006 936 2007 940
rect 2011 936 2012 940
rect 2006 935 2012 936
rect 2046 939 2052 940
rect 2046 935 2047 939
rect 2051 935 2052 939
rect 2046 934 2052 935
rect 2302 936 2308 937
rect 1434 931 1440 932
rect 1434 927 1435 931
rect 1439 927 1440 931
rect 1434 926 1440 927
rect 1582 931 1588 932
rect 1582 927 1583 931
rect 1587 927 1588 931
rect 1582 926 1588 927
rect 2006 923 2012 924
rect 1358 920 1364 921
rect 1358 916 1359 920
rect 1363 916 1364 920
rect 1358 915 1364 916
rect 1494 920 1500 921
rect 1494 916 1495 920
rect 1499 916 1500 920
rect 2006 919 2007 923
rect 2011 919 2012 923
rect 2006 918 2012 919
rect 1494 915 1500 916
rect 1360 891 1362 915
rect 1496 891 1498 915
rect 2008 891 2010 918
rect 2048 903 2050 934
rect 2302 932 2303 936
rect 2307 932 2308 936
rect 2302 931 2308 932
rect 2454 936 2460 937
rect 2454 932 2455 936
rect 2459 932 2460 936
rect 2454 931 2460 932
rect 2614 936 2620 937
rect 2614 932 2615 936
rect 2619 932 2620 936
rect 2614 931 2620 932
rect 2782 936 2788 937
rect 2782 932 2783 936
rect 2787 932 2788 936
rect 2782 931 2788 932
rect 2304 903 2306 931
rect 2456 903 2458 931
rect 2616 903 2618 931
rect 2784 903 2786 931
rect 2047 902 2051 903
rect 2047 897 2051 898
rect 2303 902 2307 903
rect 2303 897 2307 898
rect 2455 902 2459 903
rect 2455 897 2459 898
rect 2559 902 2563 903
rect 2559 897 2563 898
rect 2615 902 2619 903
rect 2615 897 2619 898
rect 2679 902 2683 903
rect 2679 897 2683 898
rect 2783 902 2787 903
rect 2783 897 2787 898
rect 2807 902 2811 903
rect 2807 897 2811 898
rect 1351 890 1355 891
rect 1351 885 1355 886
rect 1359 890 1363 891
rect 1359 885 1363 886
rect 1495 890 1499 891
rect 1495 885 1499 886
rect 2007 890 2011 891
rect 2007 885 2011 886
rect 1352 861 1354 885
rect 1350 860 1356 861
rect 1350 856 1351 860
rect 1355 856 1356 860
rect 2008 858 2010 885
rect 2048 870 2050 897
rect 2560 873 2562 897
rect 2680 873 2682 897
rect 2808 873 2810 897
rect 2558 872 2564 873
rect 2046 869 2052 870
rect 2046 865 2047 869
rect 2051 865 2052 869
rect 2558 868 2559 872
rect 2563 868 2564 872
rect 2558 867 2564 868
rect 2678 872 2684 873
rect 2678 868 2679 872
rect 2683 868 2684 872
rect 2678 867 2684 868
rect 2806 872 2812 873
rect 2806 868 2807 872
rect 2811 868 2812 872
rect 2806 867 2812 868
rect 2046 864 2052 865
rect 2634 863 2640 864
rect 2634 859 2635 863
rect 2639 859 2640 863
rect 2634 858 2640 859
rect 2754 863 2760 864
rect 2754 859 2755 863
rect 2759 859 2760 863
rect 2754 858 2760 859
rect 2882 863 2888 864
rect 2882 859 2883 863
rect 2887 859 2888 863
rect 2882 858 2888 859
rect 1350 855 1356 856
rect 2006 857 2012 858
rect 2006 853 2007 857
rect 2011 853 2012 857
rect 2558 853 2564 854
rect 2006 852 2012 853
rect 2046 852 2052 853
rect 990 851 996 852
rect 990 847 991 851
rect 995 847 996 851
rect 990 846 996 847
rect 1098 851 1104 852
rect 1098 847 1099 851
rect 1103 847 1104 851
rect 1098 846 1104 847
rect 1186 851 1192 852
rect 1186 847 1187 851
rect 1191 847 1192 851
rect 1186 846 1192 847
rect 1306 851 1312 852
rect 1306 847 1307 851
rect 1311 847 1312 851
rect 1306 846 1312 847
rect 1314 851 1320 852
rect 1314 847 1315 851
rect 1319 847 1320 851
rect 2046 848 2047 852
rect 2051 848 2052 852
rect 2558 849 2559 853
rect 2563 849 2564 853
rect 2558 848 2564 849
rect 2046 847 2052 848
rect 1314 846 1320 847
rect 750 841 756 842
rect 750 837 751 841
rect 755 837 756 841
rect 750 836 756 837
rect 878 841 884 842
rect 878 837 879 841
rect 883 837 884 841
rect 878 836 884 837
rect 698 819 704 820
rect 698 815 699 819
rect 703 815 704 819
rect 554 814 560 815
rect 615 814 619 815
rect 615 809 619 810
rect 679 814 683 815
rect 698 814 704 815
rect 714 819 720 820
rect 714 815 715 819
rect 719 815 720 819
rect 752 815 754 836
rect 880 815 882 836
rect 992 820 994 846
rect 998 841 1004 842
rect 998 837 999 841
rect 1003 837 1004 841
rect 998 836 1004 837
rect 942 819 948 820
rect 942 815 943 819
rect 947 815 948 819
rect 990 819 996 820
rect 990 815 991 819
rect 995 815 996 819
rect 1000 815 1002 836
rect 1100 820 1102 846
rect 1110 841 1116 842
rect 1110 837 1111 841
rect 1115 837 1116 841
rect 1110 836 1116 837
rect 1098 819 1104 820
rect 1098 815 1099 819
rect 1103 815 1104 819
rect 1112 815 1114 836
rect 1188 820 1190 846
rect 1230 841 1236 842
rect 1230 837 1231 841
rect 1235 837 1236 841
rect 1230 836 1236 837
rect 1186 819 1192 820
rect 1186 815 1187 819
rect 1191 815 1192 819
rect 1232 815 1234 836
rect 1308 820 1310 846
rect 1350 841 1356 842
rect 1350 837 1351 841
rect 1355 837 1356 841
rect 1350 836 1356 837
rect 2006 840 2012 841
rect 2006 836 2007 840
rect 2011 836 2012 840
rect 1306 819 1312 820
rect 1306 815 1307 819
rect 1311 815 1312 819
rect 1352 815 1354 836
rect 2006 835 2012 836
rect 2008 815 2010 835
rect 2048 823 2050 847
rect 2560 823 2562 848
rect 2636 832 2638 858
rect 2678 853 2684 854
rect 2678 849 2679 853
rect 2683 849 2684 853
rect 2678 848 2684 849
rect 2634 831 2640 832
rect 2634 827 2635 831
rect 2639 827 2640 831
rect 2634 826 2640 827
rect 2680 823 2682 848
rect 2756 832 2758 858
rect 2806 853 2812 854
rect 2806 849 2807 853
rect 2811 849 2812 853
rect 2806 848 2812 849
rect 2754 831 2760 832
rect 2754 827 2755 831
rect 2759 827 2760 831
rect 2754 826 2760 827
rect 2808 823 2810 848
rect 2884 832 2886 858
rect 2908 840 2910 942
rect 2950 936 2956 937
rect 2950 932 2951 936
rect 2955 932 2956 936
rect 2950 931 2956 932
rect 3110 936 3116 937
rect 3110 932 3111 936
rect 3115 932 3116 936
rect 3110 931 3116 932
rect 3262 936 3268 937
rect 3262 932 3263 936
rect 3267 932 3268 936
rect 3262 931 3268 932
rect 3414 936 3420 937
rect 3414 932 3415 936
rect 3419 932 3420 936
rect 3414 931 3420 932
rect 3558 936 3564 937
rect 3558 932 3559 936
rect 3563 932 3564 936
rect 3558 931 3564 932
rect 2952 903 2954 931
rect 3112 903 3114 931
rect 3264 903 3266 931
rect 3416 903 3418 931
rect 3560 903 3562 931
rect 2943 902 2947 903
rect 2943 897 2947 898
rect 2951 902 2955 903
rect 2951 897 2955 898
rect 3079 902 3083 903
rect 3079 897 3083 898
rect 3111 902 3115 903
rect 3111 897 3115 898
rect 3207 902 3211 903
rect 3207 897 3211 898
rect 3263 902 3267 903
rect 3263 897 3267 898
rect 3335 902 3339 903
rect 3335 897 3339 898
rect 3415 902 3419 903
rect 3415 897 3419 898
rect 3463 902 3467 903
rect 3463 897 3467 898
rect 3559 902 3563 903
rect 3559 897 3563 898
rect 3591 902 3595 903
rect 3591 897 3595 898
rect 2944 873 2946 897
rect 3080 873 3082 897
rect 3208 873 3210 897
rect 3336 873 3338 897
rect 3464 873 3466 897
rect 3592 873 3594 897
rect 2942 872 2948 873
rect 2942 868 2943 872
rect 2947 868 2948 872
rect 2942 867 2948 868
rect 3078 872 3084 873
rect 3078 868 3079 872
rect 3083 868 3084 872
rect 3078 867 3084 868
rect 3206 872 3212 873
rect 3206 868 3207 872
rect 3211 868 3212 872
rect 3206 867 3212 868
rect 3334 872 3340 873
rect 3334 868 3335 872
rect 3339 868 3340 872
rect 3334 867 3340 868
rect 3462 872 3468 873
rect 3462 868 3463 872
rect 3467 868 3468 872
rect 3462 867 3468 868
rect 3590 872 3596 873
rect 3590 868 3591 872
rect 3595 868 3596 872
rect 3590 867 3596 868
rect 3018 863 3024 864
rect 3018 859 3019 863
rect 3023 859 3024 863
rect 3018 858 3024 859
rect 3026 863 3032 864
rect 3026 859 3027 863
rect 3031 859 3032 863
rect 3026 858 3032 859
rect 3162 863 3168 864
rect 3162 859 3163 863
rect 3167 859 3168 863
rect 3162 858 3168 859
rect 3290 863 3296 864
rect 3290 859 3291 863
rect 3295 859 3296 863
rect 3290 858 3296 859
rect 3418 863 3424 864
rect 3418 859 3419 863
rect 3423 859 3424 863
rect 3418 858 3424 859
rect 2942 853 2948 854
rect 2942 849 2943 853
rect 2947 849 2948 853
rect 2942 848 2948 849
rect 2906 839 2912 840
rect 2906 835 2907 839
rect 2911 835 2912 839
rect 2906 834 2912 835
rect 2882 831 2888 832
rect 2882 827 2883 831
rect 2887 827 2888 831
rect 2882 826 2888 827
rect 2944 823 2946 848
rect 3020 832 3022 858
rect 3018 831 3024 832
rect 3018 827 3019 831
rect 3023 827 3024 831
rect 3018 826 3024 827
rect 2047 822 2051 823
rect 2047 817 2051 818
rect 2335 822 2339 823
rect 2335 817 2339 818
rect 2471 822 2475 823
rect 2471 817 2475 818
rect 2559 822 2563 823
rect 2559 817 2563 818
rect 2615 822 2619 823
rect 2615 817 2619 818
rect 2679 822 2683 823
rect 2679 817 2683 818
rect 2767 822 2771 823
rect 2767 817 2771 818
rect 2807 822 2811 823
rect 2807 817 2811 818
rect 2919 822 2923 823
rect 2919 817 2923 818
rect 2943 822 2947 823
rect 2943 817 2947 818
rect 714 814 720 815
rect 751 814 755 815
rect 679 809 683 810
rect 751 809 755 810
rect 815 814 819 815
rect 815 809 819 810
rect 879 814 883 815
rect 942 814 948 815
rect 951 814 955 815
rect 990 814 996 815
rect 999 814 1003 815
rect 879 809 883 810
rect 546 807 552 808
rect 546 803 547 807
rect 551 803 552 807
rect 546 802 552 803
rect 634 807 640 808
rect 634 803 635 807
rect 639 803 640 807
rect 634 802 640 803
rect 534 787 540 788
rect 534 783 535 787
rect 539 783 540 787
rect 534 782 540 783
rect 636 780 638 802
rect 680 788 682 809
rect 798 807 804 808
rect 798 803 799 807
rect 803 803 804 807
rect 798 802 804 803
rect 678 787 684 788
rect 678 783 679 787
rect 683 783 684 787
rect 678 782 684 783
rect 800 780 802 802
rect 816 788 818 809
rect 814 787 820 788
rect 814 783 815 787
rect 819 783 820 787
rect 814 782 820 783
rect 944 780 946 814
rect 951 809 955 810
rect 999 809 1003 810
rect 1079 814 1083 815
rect 1098 814 1104 815
rect 1111 814 1115 815
rect 1186 814 1192 815
rect 1199 814 1203 815
rect 1079 809 1083 810
rect 1111 809 1115 810
rect 1199 809 1203 810
rect 1231 814 1235 815
rect 1306 814 1312 815
rect 1327 814 1331 815
rect 1231 809 1235 810
rect 1327 809 1331 810
rect 1351 814 1355 815
rect 1351 809 1355 810
rect 1455 814 1459 815
rect 1455 809 1459 810
rect 2007 814 2011 815
rect 2007 809 2011 810
rect 952 788 954 809
rect 1066 807 1072 808
rect 1066 803 1067 807
rect 1071 803 1072 807
rect 1066 802 1072 803
rect 950 787 956 788
rect 950 783 951 787
rect 955 783 956 787
rect 950 782 956 783
rect 1068 780 1070 802
rect 1080 788 1082 809
rect 1178 807 1184 808
rect 1178 803 1179 807
rect 1183 803 1184 807
rect 1178 802 1184 803
rect 1078 787 1084 788
rect 1078 783 1079 787
rect 1083 783 1084 787
rect 1078 782 1084 783
rect 1180 780 1182 802
rect 1200 788 1202 809
rect 1328 788 1330 809
rect 1370 807 1376 808
rect 1370 803 1371 807
rect 1375 803 1376 807
rect 1370 802 1376 803
rect 1402 807 1408 808
rect 1402 803 1403 807
rect 1407 803 1408 807
rect 1402 802 1408 803
rect 1198 787 1204 788
rect 1198 783 1199 787
rect 1203 783 1204 787
rect 1198 782 1204 783
rect 1326 787 1332 788
rect 1326 783 1327 787
rect 1331 783 1332 787
rect 1326 782 1332 783
rect 634 779 640 780
rect 634 775 635 779
rect 639 775 640 779
rect 634 774 640 775
rect 798 779 804 780
rect 798 775 799 779
rect 803 775 804 779
rect 942 779 948 780
rect 798 774 804 775
rect 890 775 896 776
rect 890 771 891 775
rect 895 771 896 775
rect 942 775 943 779
rect 947 775 948 779
rect 942 774 948 775
rect 1066 779 1072 780
rect 1066 775 1067 779
rect 1071 775 1072 779
rect 1066 774 1072 775
rect 1178 779 1184 780
rect 1178 775 1179 779
rect 1183 775 1184 779
rect 1178 774 1184 775
rect 890 770 896 771
rect 534 768 540 769
rect 534 764 535 768
rect 539 764 540 768
rect 534 763 540 764
rect 678 768 684 769
rect 678 764 679 768
rect 683 764 684 768
rect 678 763 684 764
rect 814 768 820 769
rect 814 764 815 768
rect 819 764 820 768
rect 814 763 820 764
rect 536 735 538 763
rect 680 735 682 763
rect 816 735 818 763
rect 471 734 475 735
rect 471 729 475 730
rect 535 734 539 735
rect 535 729 539 730
rect 639 734 643 735
rect 639 729 643 730
rect 679 734 683 735
rect 679 729 683 730
rect 807 734 811 735
rect 807 729 811 730
rect 815 734 819 735
rect 815 729 819 730
rect 472 705 474 729
rect 640 705 642 729
rect 808 705 810 729
rect 470 704 476 705
rect 470 700 471 704
rect 475 700 476 704
rect 470 699 476 700
rect 638 704 644 705
rect 638 700 639 704
rect 643 700 644 704
rect 638 699 644 700
rect 806 704 812 705
rect 806 700 807 704
rect 811 700 812 704
rect 806 699 812 700
rect 402 695 408 696
rect 402 691 403 695
rect 407 691 408 695
rect 402 690 408 691
rect 546 695 552 696
rect 546 691 547 695
rect 551 691 552 695
rect 546 690 552 691
rect 554 695 560 696
rect 554 691 555 695
rect 559 691 560 695
rect 554 690 560 691
rect 310 685 316 686
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 310 681 311 685
rect 315 681 316 685
rect 310 680 316 681
rect 470 685 476 686
rect 470 681 471 685
rect 475 681 476 685
rect 470 680 476 681
rect 110 679 116 680
rect 112 659 114 679
rect 312 659 314 680
rect 472 659 474 680
rect 548 664 550 690
rect 556 672 558 690
rect 638 685 644 686
rect 638 681 639 685
rect 643 681 644 685
rect 638 680 644 681
rect 806 685 812 686
rect 806 681 807 685
rect 811 681 812 685
rect 806 680 812 681
rect 554 671 560 672
rect 554 667 555 671
rect 559 667 560 671
rect 554 666 560 667
rect 522 663 528 664
rect 522 659 523 663
rect 527 659 528 663
rect 111 658 115 659
rect 111 653 115 654
rect 295 658 299 659
rect 295 653 299 654
rect 311 658 315 659
rect 311 653 315 654
rect 447 658 451 659
rect 447 653 451 654
rect 471 658 475 659
rect 522 658 528 659
rect 546 663 552 664
rect 546 659 547 663
rect 551 659 552 663
rect 640 659 642 680
rect 808 659 810 680
rect 892 664 894 770
rect 950 768 956 769
rect 950 764 951 768
rect 955 764 956 768
rect 950 763 956 764
rect 1078 768 1084 769
rect 1078 764 1079 768
rect 1083 764 1084 768
rect 1078 763 1084 764
rect 1198 768 1204 769
rect 1198 764 1199 768
rect 1203 764 1204 768
rect 1198 763 1204 764
rect 1326 768 1332 769
rect 1326 764 1327 768
rect 1331 764 1332 768
rect 1326 763 1332 764
rect 952 735 954 763
rect 1080 735 1082 763
rect 1200 735 1202 763
rect 1328 735 1330 763
rect 951 734 955 735
rect 951 729 955 730
rect 975 734 979 735
rect 975 729 979 730
rect 1079 734 1083 735
rect 1079 729 1083 730
rect 1135 734 1139 735
rect 1135 729 1139 730
rect 1199 734 1203 735
rect 1199 729 1203 730
rect 1295 734 1299 735
rect 1295 729 1299 730
rect 1327 734 1331 735
rect 1327 729 1331 730
rect 976 705 978 729
rect 1136 705 1138 729
rect 1296 705 1298 729
rect 974 704 980 705
rect 974 700 975 704
rect 979 700 980 704
rect 974 699 980 700
rect 1134 704 1140 705
rect 1134 700 1135 704
rect 1139 700 1140 704
rect 1134 699 1140 700
rect 1294 704 1300 705
rect 1294 700 1295 704
rect 1299 700 1300 704
rect 1294 699 1300 700
rect 1372 696 1374 802
rect 1404 780 1406 802
rect 1410 799 1416 800
rect 1410 795 1411 799
rect 1415 795 1416 799
rect 1410 794 1416 795
rect 1412 780 1414 794
rect 1456 788 1458 809
rect 2008 789 2010 809
rect 2048 797 2050 817
rect 2046 796 2052 797
rect 2336 796 2338 817
rect 2410 815 2416 816
rect 2410 811 2411 815
rect 2415 811 2416 815
rect 2410 810 2416 811
rect 2046 792 2047 796
rect 2051 792 2052 796
rect 2046 791 2052 792
rect 2334 795 2340 796
rect 2334 791 2335 795
rect 2339 791 2340 795
rect 2334 790 2340 791
rect 2006 788 2012 789
rect 2412 788 2414 810
rect 2472 796 2474 817
rect 2546 815 2552 816
rect 2546 811 2547 815
rect 2551 811 2552 815
rect 2546 810 2552 811
rect 2470 795 2476 796
rect 2470 791 2471 795
rect 2475 791 2476 795
rect 2470 790 2476 791
rect 2548 788 2550 810
rect 2616 796 2618 817
rect 2718 807 2724 808
rect 2718 803 2719 807
rect 2723 803 2724 807
rect 2718 802 2724 803
rect 2614 795 2620 796
rect 2614 791 2615 795
rect 2619 791 2620 795
rect 2614 790 2620 791
rect 2720 788 2722 802
rect 2768 796 2770 817
rect 2854 815 2860 816
rect 2854 811 2855 815
rect 2859 811 2860 815
rect 2854 810 2860 811
rect 2766 795 2772 796
rect 2766 791 2767 795
rect 2771 791 2772 795
rect 2766 790 2772 791
rect 2856 788 2858 810
rect 2920 796 2922 817
rect 3028 816 3030 858
rect 3078 853 3084 854
rect 3078 849 3079 853
rect 3083 849 3084 853
rect 3078 848 3084 849
rect 3080 823 3082 848
rect 3079 822 3083 823
rect 3079 817 3083 818
rect 3026 815 3032 816
rect 3026 811 3027 815
rect 3031 811 3032 815
rect 3026 810 3032 811
rect 3080 796 3082 817
rect 3164 816 3166 858
rect 3206 853 3212 854
rect 3206 849 3207 853
rect 3211 849 3212 853
rect 3206 848 3212 849
rect 3208 823 3210 848
rect 3292 832 3294 858
rect 3334 853 3340 854
rect 3334 849 3335 853
rect 3339 849 3340 853
rect 3334 848 3340 849
rect 3290 831 3296 832
rect 3290 827 3291 831
rect 3295 827 3296 831
rect 3290 826 3296 827
rect 3336 823 3338 848
rect 3420 832 3422 858
rect 3462 853 3468 854
rect 3462 849 3463 853
rect 3467 849 3468 853
rect 3462 848 3468 849
rect 3590 853 3596 854
rect 3590 849 3591 853
rect 3595 849 3596 853
rect 3590 848 3596 849
rect 3418 831 3424 832
rect 3418 827 3419 831
rect 3423 827 3424 831
rect 3418 826 3424 827
rect 3464 823 3466 848
rect 3592 823 3594 848
rect 3644 840 3646 942
rect 3710 936 3716 937
rect 3710 932 3711 936
rect 3715 932 3716 936
rect 3710 931 3716 932
rect 3712 903 3714 931
rect 3711 902 3715 903
rect 3711 897 3715 898
rect 3727 902 3731 903
rect 3727 897 3731 898
rect 3728 873 3730 897
rect 3726 872 3732 873
rect 3726 868 3727 872
rect 3731 868 3732 872
rect 3726 867 3732 868
rect 3796 864 3798 970
rect 3840 956 3842 977
rect 3908 976 3910 1018
rect 3942 1012 3948 1013
rect 3942 1008 3943 1012
rect 3947 1008 3948 1012
rect 3942 1007 3948 1008
rect 3944 983 3946 1007
rect 3943 982 3947 983
rect 3943 977 3947 978
rect 3906 975 3912 976
rect 3906 971 3907 975
rect 3911 971 3912 975
rect 3906 970 3912 971
rect 3944 957 3946 977
rect 3942 956 3948 957
rect 3838 955 3844 956
rect 3838 951 3839 955
rect 3843 951 3844 955
rect 3942 952 3943 956
rect 3947 952 3948 956
rect 3942 951 3948 952
rect 3838 950 3844 951
rect 3914 943 3920 944
rect 3914 939 3915 943
rect 3919 939 3920 943
rect 3914 938 3920 939
rect 3942 939 3948 940
rect 3838 936 3844 937
rect 3838 932 3839 936
rect 3843 932 3844 936
rect 3838 931 3844 932
rect 3840 903 3842 931
rect 3839 902 3843 903
rect 3839 897 3843 898
rect 3840 873 3842 897
rect 3838 872 3844 873
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 3838 867 3844 868
rect 3666 863 3672 864
rect 3666 859 3667 863
rect 3671 859 3672 863
rect 3666 858 3672 859
rect 3794 863 3800 864
rect 3794 859 3795 863
rect 3799 859 3800 863
rect 3794 858 3800 859
rect 3906 863 3912 864
rect 3906 859 3907 863
rect 3911 859 3912 863
rect 3906 858 3912 859
rect 3642 839 3648 840
rect 3642 835 3643 839
rect 3647 835 3648 839
rect 3642 834 3648 835
rect 3668 832 3670 858
rect 3726 853 3732 854
rect 3726 849 3727 853
rect 3731 849 3732 853
rect 3726 848 3732 849
rect 3838 853 3844 854
rect 3838 849 3839 853
rect 3843 849 3844 853
rect 3838 848 3844 849
rect 3618 831 3624 832
rect 3618 827 3619 831
rect 3623 827 3624 831
rect 3618 826 3624 827
rect 3666 831 3672 832
rect 3666 827 3667 831
rect 3671 827 3672 831
rect 3666 826 3672 827
rect 3207 822 3211 823
rect 3207 817 3211 818
rect 3239 822 3243 823
rect 3239 817 3243 818
rect 3335 822 3339 823
rect 3335 817 3339 818
rect 3391 822 3395 823
rect 3391 817 3395 818
rect 3463 822 3467 823
rect 3463 817 3467 818
rect 3543 822 3547 823
rect 3543 817 3547 818
rect 3591 822 3595 823
rect 3591 817 3595 818
rect 3162 815 3168 816
rect 3162 811 3163 815
rect 3167 811 3168 815
rect 3162 810 3168 811
rect 3240 796 3242 817
rect 3314 815 3320 816
rect 3314 811 3315 815
rect 3319 811 3320 815
rect 3314 810 3320 811
rect 2918 795 2924 796
rect 2918 791 2919 795
rect 2923 791 2924 795
rect 2918 790 2924 791
rect 3078 795 3084 796
rect 3078 791 3079 795
rect 3083 791 3084 795
rect 3078 790 3084 791
rect 3238 795 3244 796
rect 3238 791 3239 795
rect 3243 791 3244 795
rect 3238 790 3244 791
rect 3316 788 3318 810
rect 3392 796 3394 817
rect 3544 796 3546 817
rect 3390 795 3396 796
rect 3390 791 3391 795
rect 3395 791 3396 795
rect 3390 790 3396 791
rect 3542 795 3548 796
rect 3542 791 3543 795
rect 3547 791 3548 795
rect 3542 790 3548 791
rect 3620 788 3622 826
rect 3728 823 3730 848
rect 3840 823 3842 848
rect 3703 822 3707 823
rect 3703 817 3707 818
rect 3727 822 3731 823
rect 3727 817 3731 818
rect 3839 822 3843 823
rect 3839 817 3843 818
rect 3642 815 3648 816
rect 3642 811 3643 815
rect 3647 811 3648 815
rect 3642 810 3648 811
rect 3644 788 3646 810
rect 3704 796 3706 817
rect 3770 815 3776 816
rect 3770 811 3771 815
rect 3775 811 3776 815
rect 3770 810 3776 811
rect 3702 795 3708 796
rect 3702 791 3703 795
rect 3707 791 3708 795
rect 3702 790 3708 791
rect 1454 787 1460 788
rect 1454 783 1455 787
rect 1459 783 1460 787
rect 2006 784 2007 788
rect 2011 784 2012 788
rect 2006 783 2012 784
rect 2410 787 2416 788
rect 2410 783 2411 787
rect 2415 783 2416 787
rect 1454 782 1460 783
rect 2410 782 2416 783
rect 2546 787 2552 788
rect 2546 783 2547 787
rect 2551 783 2552 787
rect 2718 787 2724 788
rect 2546 782 2552 783
rect 2690 783 2696 784
rect 1402 779 1408 780
rect 1402 775 1403 779
rect 1407 775 1408 779
rect 1402 774 1408 775
rect 1410 779 1416 780
rect 1410 775 1411 779
rect 1415 775 1416 779
rect 1410 774 1416 775
rect 2046 779 2052 780
rect 2046 775 2047 779
rect 2051 775 2052 779
rect 2690 779 2691 783
rect 2695 779 2696 783
rect 2718 783 2719 787
rect 2723 783 2724 787
rect 2718 782 2724 783
rect 2854 787 2860 788
rect 2854 783 2855 787
rect 2859 783 2860 787
rect 2854 782 2860 783
rect 3314 787 3320 788
rect 3314 783 3315 787
rect 3319 783 3320 787
rect 3618 787 3624 788
rect 3314 782 3320 783
rect 3466 783 3472 784
rect 2690 778 2696 779
rect 3466 779 3467 783
rect 3471 779 3472 783
rect 3618 783 3619 787
rect 3623 783 3624 787
rect 3618 782 3624 783
rect 3642 787 3648 788
rect 3642 783 3643 787
rect 3647 783 3648 787
rect 3642 782 3648 783
rect 3466 778 3472 779
rect 2046 774 2052 775
rect 2334 776 2340 777
rect 2006 771 2012 772
rect 1454 768 1460 769
rect 1454 764 1455 768
rect 1459 764 1460 768
rect 2006 767 2007 771
rect 2011 767 2012 771
rect 2006 766 2012 767
rect 1454 763 1460 764
rect 1456 735 1458 763
rect 2008 735 2010 766
rect 2048 743 2050 774
rect 2334 772 2335 776
rect 2339 772 2340 776
rect 2334 771 2340 772
rect 2470 776 2476 777
rect 2470 772 2471 776
rect 2475 772 2476 776
rect 2470 771 2476 772
rect 2614 776 2620 777
rect 2614 772 2615 776
rect 2619 772 2620 776
rect 2614 771 2620 772
rect 2336 743 2338 771
rect 2472 743 2474 771
rect 2616 743 2618 771
rect 2047 742 2051 743
rect 2047 737 2051 738
rect 2071 742 2075 743
rect 2071 737 2075 738
rect 2183 742 2187 743
rect 2183 737 2187 738
rect 2335 742 2339 743
rect 2335 737 2339 738
rect 2471 742 2475 743
rect 2471 737 2475 738
rect 2487 742 2491 743
rect 2487 737 2491 738
rect 2615 742 2619 743
rect 2615 737 2619 738
rect 2639 742 2643 743
rect 2639 737 2643 738
rect 1455 734 1459 735
rect 1455 729 1459 730
rect 1607 734 1611 735
rect 1607 729 1611 730
rect 1767 734 1771 735
rect 1767 729 1771 730
rect 1903 734 1907 735
rect 1903 729 1907 730
rect 2007 734 2011 735
rect 2007 729 2011 730
rect 1456 705 1458 729
rect 1608 705 1610 729
rect 1768 705 1770 729
rect 1904 705 1906 729
rect 1454 704 1460 705
rect 1454 700 1455 704
rect 1459 700 1460 704
rect 1454 699 1460 700
rect 1606 704 1612 705
rect 1606 700 1607 704
rect 1611 700 1612 704
rect 1606 699 1612 700
rect 1766 704 1772 705
rect 1766 700 1767 704
rect 1771 700 1772 704
rect 1766 699 1772 700
rect 1902 704 1908 705
rect 1902 700 1903 704
rect 1907 700 1908 704
rect 2008 702 2010 729
rect 2048 710 2050 737
rect 2072 713 2074 737
rect 2184 713 2186 737
rect 2336 713 2338 737
rect 2488 713 2490 737
rect 2640 713 2642 737
rect 2070 712 2076 713
rect 2046 709 2052 710
rect 2046 705 2047 709
rect 2051 705 2052 709
rect 2070 708 2071 712
rect 2075 708 2076 712
rect 2070 707 2076 708
rect 2182 712 2188 713
rect 2182 708 2183 712
rect 2187 708 2188 712
rect 2182 707 2188 708
rect 2334 712 2340 713
rect 2334 708 2335 712
rect 2339 708 2340 712
rect 2334 707 2340 708
rect 2486 712 2492 713
rect 2486 708 2487 712
rect 2491 708 2492 712
rect 2486 707 2492 708
rect 2638 712 2644 713
rect 2638 708 2639 712
rect 2643 708 2644 712
rect 2638 707 2644 708
rect 2046 704 2052 705
rect 2054 703 2060 704
rect 1902 699 1908 700
rect 2006 701 2012 702
rect 2006 697 2007 701
rect 2011 697 2012 701
rect 2054 699 2055 703
rect 2059 699 2060 703
rect 2054 698 2060 699
rect 2154 703 2160 704
rect 2154 699 2155 703
rect 2159 699 2160 703
rect 2154 698 2160 699
rect 2266 703 2272 704
rect 2266 699 2267 703
rect 2271 699 2272 703
rect 2266 698 2272 699
rect 2418 703 2424 704
rect 2418 699 2419 703
rect 2423 699 2424 703
rect 2418 698 2424 699
rect 2570 703 2576 704
rect 2570 699 2571 703
rect 2575 699 2576 703
rect 2570 698 2576 699
rect 2006 696 2012 697
rect 942 695 948 696
rect 942 691 943 695
rect 947 691 948 695
rect 942 690 948 691
rect 1042 695 1048 696
rect 1042 691 1043 695
rect 1047 691 1048 695
rect 1042 690 1048 691
rect 1210 695 1216 696
rect 1210 691 1211 695
rect 1215 691 1216 695
rect 1210 690 1216 691
rect 1370 695 1376 696
rect 1370 691 1371 695
rect 1375 691 1376 695
rect 1370 690 1376 691
rect 1582 695 1588 696
rect 1582 691 1583 695
rect 1587 691 1588 695
rect 1582 690 1588 691
rect 1682 695 1688 696
rect 1682 691 1683 695
rect 1687 691 1688 695
rect 1682 690 1688 691
rect 1698 695 1704 696
rect 1698 691 1699 695
rect 1703 691 1704 695
rect 1698 690 1704 691
rect 1858 695 1864 696
rect 1858 691 1859 695
rect 1863 691 1864 695
rect 1858 690 1864 691
rect 2046 692 2052 693
rect 944 664 946 690
rect 974 685 980 686
rect 974 681 975 685
rect 979 681 980 685
rect 974 680 980 681
rect 890 663 896 664
rect 890 659 891 663
rect 895 659 896 663
rect 546 658 552 659
rect 615 658 619 659
rect 471 653 475 654
rect 112 633 114 653
rect 110 632 116 633
rect 296 632 298 653
rect 370 651 376 652
rect 314 647 320 648
rect 314 643 315 647
rect 319 643 320 647
rect 370 647 371 651
rect 375 647 376 651
rect 370 646 376 647
rect 314 642 320 643
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 294 631 300 632
rect 294 627 295 631
rect 299 627 300 631
rect 294 626 300 627
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 110 610 116 611
rect 294 612 300 613
rect 112 579 114 610
rect 294 608 295 612
rect 299 608 300 612
rect 294 607 300 608
rect 296 579 298 607
rect 111 578 115 579
rect 111 573 115 574
rect 239 578 243 579
rect 239 573 243 574
rect 295 578 299 579
rect 295 573 299 574
rect 112 546 114 573
rect 240 549 242 573
rect 238 548 244 549
rect 110 545 116 546
rect 110 541 111 545
rect 115 541 116 545
rect 238 544 239 548
rect 243 544 244 548
rect 238 543 244 544
rect 110 540 116 541
rect 316 540 318 642
rect 372 624 374 646
rect 448 632 450 653
rect 446 631 452 632
rect 446 627 447 631
rect 451 627 452 631
rect 446 626 452 627
rect 524 624 526 658
rect 615 653 619 654
rect 639 658 643 659
rect 639 653 643 654
rect 783 658 787 659
rect 783 653 787 654
rect 807 658 811 659
rect 890 658 896 659
rect 942 663 948 664
rect 942 659 943 663
rect 947 659 948 663
rect 976 659 978 680
rect 942 658 948 659
rect 951 658 955 659
rect 807 653 811 654
rect 951 653 955 654
rect 975 658 979 659
rect 975 653 979 654
rect 616 632 618 653
rect 698 651 704 652
rect 698 647 699 651
rect 703 647 704 651
rect 698 646 704 647
rect 614 631 620 632
rect 614 627 615 631
rect 619 627 620 631
rect 614 626 620 627
rect 700 624 702 646
rect 784 632 786 653
rect 866 651 872 652
rect 866 647 867 651
rect 871 647 872 651
rect 866 646 872 647
rect 782 631 788 632
rect 782 627 783 631
rect 787 627 788 631
rect 782 626 788 627
rect 868 624 870 646
rect 952 632 954 653
rect 1044 652 1046 690
rect 1134 685 1140 686
rect 1134 681 1135 685
rect 1139 681 1140 685
rect 1134 680 1140 681
rect 1136 659 1138 680
rect 1203 668 1207 669
rect 1212 664 1214 690
rect 1294 685 1300 686
rect 1294 681 1295 685
rect 1299 681 1300 685
rect 1294 680 1300 681
rect 1454 685 1460 686
rect 1454 681 1455 685
rect 1459 681 1460 685
rect 1454 680 1460 681
rect 1202 663 1208 664
rect 1202 659 1203 663
rect 1207 659 1208 663
rect 1111 658 1115 659
rect 1111 653 1115 654
rect 1135 658 1139 659
rect 1202 658 1208 659
rect 1210 663 1216 664
rect 1210 659 1211 663
rect 1215 659 1216 663
rect 1296 659 1298 680
rect 1456 659 1458 680
rect 1584 664 1586 690
rect 1606 685 1612 686
rect 1606 681 1607 685
rect 1611 681 1612 685
rect 1606 680 1612 681
rect 1474 663 1480 664
rect 1474 659 1475 663
rect 1479 659 1480 663
rect 1582 663 1588 664
rect 1582 659 1583 663
rect 1587 659 1588 663
rect 1608 659 1610 680
rect 1684 664 1686 690
rect 1700 669 1702 690
rect 1766 685 1772 686
rect 1766 681 1767 685
rect 1771 681 1772 685
rect 1766 680 1772 681
rect 1699 668 1703 669
rect 1682 663 1688 664
rect 1699 663 1703 664
rect 1682 659 1683 663
rect 1687 659 1688 663
rect 1768 659 1770 680
rect 1210 658 1216 659
rect 1263 658 1267 659
rect 1135 653 1139 654
rect 1263 653 1267 654
rect 1295 658 1299 659
rect 1295 653 1299 654
rect 1399 658 1403 659
rect 1399 653 1403 654
rect 1455 658 1459 659
rect 1474 658 1480 659
rect 1535 658 1539 659
rect 1582 658 1588 659
rect 1607 658 1611 659
rect 1455 653 1459 654
rect 1042 651 1048 652
rect 1042 647 1043 651
rect 1047 647 1048 651
rect 1042 646 1048 647
rect 1112 632 1114 653
rect 1186 651 1192 652
rect 1186 647 1187 651
rect 1191 647 1192 651
rect 1186 646 1192 647
rect 950 631 956 632
rect 950 627 951 631
rect 955 627 956 631
rect 950 626 956 627
rect 1110 631 1116 632
rect 1110 627 1111 631
rect 1115 627 1116 631
rect 1110 626 1116 627
rect 1188 624 1190 646
rect 1264 632 1266 653
rect 1338 651 1344 652
rect 1338 647 1339 651
rect 1343 647 1344 651
rect 1338 646 1344 647
rect 1262 631 1268 632
rect 1262 627 1263 631
rect 1267 627 1268 631
rect 1262 626 1268 627
rect 1340 624 1342 646
rect 1400 632 1402 653
rect 1398 631 1404 632
rect 1398 627 1399 631
rect 1403 627 1404 631
rect 1398 626 1404 627
rect 1476 624 1478 658
rect 1535 653 1539 654
rect 1607 653 1611 654
rect 1663 658 1667 659
rect 1682 658 1688 659
rect 1767 658 1771 659
rect 1663 653 1667 654
rect 1767 653 1771 654
rect 1791 658 1795 659
rect 1791 653 1795 654
rect 1482 643 1488 644
rect 1482 639 1483 643
rect 1487 639 1488 643
rect 1482 638 1488 639
rect 1484 624 1486 638
rect 1536 632 1538 653
rect 1618 651 1624 652
rect 1618 647 1619 651
rect 1623 647 1624 651
rect 1618 646 1624 647
rect 1534 631 1540 632
rect 1534 627 1535 631
rect 1539 627 1540 631
rect 1534 626 1540 627
rect 1620 624 1622 646
rect 1664 632 1666 653
rect 1792 632 1794 653
rect 1860 652 1862 690
rect 2046 688 2047 692
rect 2051 688 2052 692
rect 2046 687 2052 688
rect 1902 685 1908 686
rect 1902 681 1903 685
rect 1907 681 1908 685
rect 1902 680 1908 681
rect 2006 684 2012 685
rect 2006 680 2007 684
rect 2011 680 2012 684
rect 1904 659 1906 680
rect 2006 679 2012 680
rect 2008 659 2010 679
rect 1903 658 1907 659
rect 1903 653 1907 654
rect 2007 658 2011 659
rect 2048 655 2050 687
rect 2056 664 2058 698
rect 2070 693 2076 694
rect 2070 689 2071 693
rect 2075 689 2076 693
rect 2070 688 2076 689
rect 2054 663 2060 664
rect 2054 659 2055 663
rect 2059 659 2060 663
rect 2054 658 2060 659
rect 2072 655 2074 688
rect 2156 672 2158 698
rect 2182 693 2188 694
rect 2182 689 2183 693
rect 2187 689 2188 693
rect 2182 688 2188 689
rect 2154 671 2160 672
rect 2154 667 2155 671
rect 2159 667 2160 671
rect 2154 666 2160 667
rect 2184 655 2186 688
rect 2268 672 2270 698
rect 2334 693 2340 694
rect 2334 689 2335 693
rect 2339 689 2340 693
rect 2334 688 2340 689
rect 2266 671 2272 672
rect 2266 667 2267 671
rect 2271 667 2272 671
rect 2266 666 2272 667
rect 2336 655 2338 688
rect 2420 672 2422 698
rect 2486 693 2492 694
rect 2486 689 2487 693
rect 2491 689 2492 693
rect 2486 688 2492 689
rect 2418 671 2424 672
rect 2418 667 2419 671
rect 2423 667 2424 671
rect 2418 666 2424 667
rect 2488 655 2490 688
rect 2572 672 2574 698
rect 2638 693 2644 694
rect 2638 689 2639 693
rect 2643 689 2644 693
rect 2638 688 2644 689
rect 2570 671 2576 672
rect 2570 667 2571 671
rect 2575 667 2576 671
rect 2570 666 2576 667
rect 2640 655 2642 688
rect 2692 672 2694 778
rect 2766 776 2772 777
rect 2766 772 2767 776
rect 2771 772 2772 776
rect 2766 771 2772 772
rect 2918 776 2924 777
rect 2918 772 2919 776
rect 2923 772 2924 776
rect 2918 771 2924 772
rect 3078 776 3084 777
rect 3078 772 3079 776
rect 3083 772 3084 776
rect 3078 771 3084 772
rect 3238 776 3244 777
rect 3238 772 3239 776
rect 3243 772 3244 776
rect 3238 771 3244 772
rect 3390 776 3396 777
rect 3390 772 3391 776
rect 3395 772 3396 776
rect 3390 771 3396 772
rect 2768 743 2770 771
rect 2920 743 2922 771
rect 3080 743 3082 771
rect 3240 743 3242 771
rect 3392 743 3394 771
rect 2767 742 2771 743
rect 2767 737 2771 738
rect 2807 742 2811 743
rect 2807 737 2811 738
rect 2919 742 2923 743
rect 2919 737 2923 738
rect 2983 742 2987 743
rect 2983 737 2987 738
rect 3079 742 3083 743
rect 3079 737 3083 738
rect 3167 742 3171 743
rect 3167 737 3171 738
rect 3239 742 3243 743
rect 3239 737 3243 738
rect 3367 742 3371 743
rect 3367 737 3371 738
rect 3391 742 3395 743
rect 3391 737 3395 738
rect 2808 713 2810 737
rect 2984 713 2986 737
rect 3168 713 3170 737
rect 3368 713 3370 737
rect 2806 712 2812 713
rect 2806 708 2807 712
rect 2811 708 2812 712
rect 2806 707 2812 708
rect 2982 712 2988 713
rect 2982 708 2983 712
rect 2987 708 2988 712
rect 2982 707 2988 708
rect 3166 712 3172 713
rect 3166 708 3167 712
rect 3171 708 3172 712
rect 3166 707 3172 708
rect 3366 712 3372 713
rect 3366 708 3367 712
rect 3371 708 3372 712
rect 3366 707 3372 708
rect 2882 703 2888 704
rect 2882 699 2883 703
rect 2887 699 2888 703
rect 2882 698 2888 699
rect 3058 703 3064 704
rect 3058 699 3059 703
rect 3063 699 3064 703
rect 3058 698 3064 699
rect 3242 703 3248 704
rect 3242 699 3243 703
rect 3247 699 3248 703
rect 3242 698 3248 699
rect 3318 703 3324 704
rect 3318 699 3319 703
rect 3323 699 3324 703
rect 3318 698 3324 699
rect 3450 703 3456 704
rect 3450 699 3451 703
rect 3455 699 3456 703
rect 3450 698 3456 699
rect 2806 693 2812 694
rect 2806 689 2807 693
rect 2811 689 2812 693
rect 2806 688 2812 689
rect 2690 671 2696 672
rect 2690 667 2691 671
rect 2695 667 2696 671
rect 2690 666 2696 667
rect 2808 655 2810 688
rect 2884 672 2886 698
rect 2982 693 2988 694
rect 2982 689 2983 693
rect 2987 689 2988 693
rect 2982 688 2988 689
rect 2882 671 2888 672
rect 2882 667 2883 671
rect 2887 667 2888 671
rect 2882 666 2888 667
rect 2984 655 2986 688
rect 3060 672 3062 698
rect 3166 693 3172 694
rect 3166 689 3167 693
rect 3171 689 3172 693
rect 3166 688 3172 689
rect 3058 671 3064 672
rect 3058 667 3059 671
rect 3063 667 3064 671
rect 3058 666 3064 667
rect 3168 655 3170 688
rect 2007 653 2011 654
rect 2047 654 2051 655
rect 1818 651 1824 652
rect 1818 647 1819 651
rect 1823 647 1824 651
rect 1818 646 1824 647
rect 1858 651 1864 652
rect 1858 647 1859 651
rect 1863 647 1864 651
rect 1858 646 1864 647
rect 1866 651 1872 652
rect 1866 647 1867 651
rect 1871 647 1872 651
rect 1866 646 1872 647
rect 1662 631 1668 632
rect 1662 627 1663 631
rect 1667 627 1668 631
rect 1662 626 1668 627
rect 1790 631 1796 632
rect 1790 627 1791 631
rect 1795 627 1796 631
rect 1790 626 1796 627
rect 370 623 376 624
rect 370 619 371 623
rect 375 619 376 623
rect 370 618 376 619
rect 522 623 528 624
rect 522 619 523 623
rect 527 619 528 623
rect 698 623 704 624
rect 522 618 528 619
rect 690 619 696 620
rect 690 615 691 619
rect 695 615 696 619
rect 698 619 699 623
rect 703 619 704 623
rect 698 618 704 619
rect 866 623 872 624
rect 866 619 867 623
rect 871 619 872 623
rect 866 618 872 619
rect 1186 623 1192 624
rect 1186 619 1187 623
rect 1191 619 1192 623
rect 1186 618 1192 619
rect 1338 623 1344 624
rect 1338 619 1339 623
rect 1343 619 1344 623
rect 1338 618 1344 619
rect 1474 623 1480 624
rect 1474 619 1475 623
rect 1479 619 1480 623
rect 1474 618 1480 619
rect 1482 623 1488 624
rect 1482 619 1483 623
rect 1487 619 1488 623
rect 1482 618 1488 619
rect 1618 623 1624 624
rect 1618 619 1619 623
rect 1623 619 1624 623
rect 1618 618 1624 619
rect 690 614 696 615
rect 446 612 452 613
rect 446 608 447 612
rect 451 608 452 612
rect 446 607 452 608
rect 614 612 620 613
rect 614 608 615 612
rect 619 608 620 612
rect 614 607 620 608
rect 448 579 450 607
rect 616 579 618 607
rect 415 578 419 579
rect 415 573 419 574
rect 447 578 451 579
rect 447 573 451 574
rect 607 578 611 579
rect 607 573 611 574
rect 615 578 619 579
rect 615 573 619 574
rect 416 549 418 573
rect 608 549 610 573
rect 414 548 420 549
rect 414 544 415 548
rect 419 544 420 548
rect 414 543 420 544
rect 606 548 612 549
rect 606 544 607 548
rect 611 544 612 548
rect 606 543 612 544
rect 314 539 320 540
rect 314 535 315 539
rect 319 535 320 539
rect 314 534 320 535
rect 370 539 376 540
rect 370 535 371 539
rect 375 535 376 539
rect 370 534 376 535
rect 238 529 244 530
rect 110 528 116 529
rect 110 524 111 528
rect 115 524 116 528
rect 238 525 239 529
rect 243 525 244 529
rect 238 524 244 525
rect 110 523 116 524
rect 112 503 114 523
rect 240 503 242 524
rect 372 508 374 534
rect 414 529 420 530
rect 414 525 415 529
rect 419 525 420 529
rect 414 524 420 525
rect 606 529 612 530
rect 606 525 607 529
rect 611 525 612 529
rect 606 524 612 525
rect 370 507 376 508
rect 370 503 371 507
rect 375 503 376 507
rect 416 503 418 524
rect 538 507 544 508
rect 538 503 539 507
rect 543 503 544 507
rect 608 503 610 524
rect 692 508 694 614
rect 782 612 788 613
rect 782 608 783 612
rect 787 608 788 612
rect 782 607 788 608
rect 950 612 956 613
rect 950 608 951 612
rect 955 608 956 612
rect 950 607 956 608
rect 1110 612 1116 613
rect 1110 608 1111 612
rect 1115 608 1116 612
rect 1110 607 1116 608
rect 1262 612 1268 613
rect 1262 608 1263 612
rect 1267 608 1268 612
rect 1262 607 1268 608
rect 1398 612 1404 613
rect 1398 608 1399 612
rect 1403 608 1404 612
rect 1398 607 1404 608
rect 1534 612 1540 613
rect 1534 608 1535 612
rect 1539 608 1540 612
rect 1534 607 1540 608
rect 1662 612 1668 613
rect 1662 608 1663 612
rect 1667 608 1668 612
rect 1662 607 1668 608
rect 1790 612 1796 613
rect 1790 608 1791 612
rect 1795 608 1796 612
rect 1790 607 1796 608
rect 784 579 786 607
rect 952 579 954 607
rect 1112 579 1114 607
rect 1264 579 1266 607
rect 1400 579 1402 607
rect 1536 579 1538 607
rect 1664 579 1666 607
rect 1792 579 1794 607
rect 783 578 787 579
rect 783 573 787 574
rect 799 578 803 579
rect 799 573 803 574
rect 951 578 955 579
rect 951 573 955 574
rect 991 578 995 579
rect 991 573 995 574
rect 1111 578 1115 579
rect 1111 573 1115 574
rect 1175 578 1179 579
rect 1175 573 1179 574
rect 1263 578 1267 579
rect 1263 573 1267 574
rect 1351 578 1355 579
rect 1351 573 1355 574
rect 1399 578 1403 579
rect 1399 573 1403 574
rect 1519 578 1523 579
rect 1519 573 1523 574
rect 1535 578 1539 579
rect 1535 573 1539 574
rect 1663 578 1667 579
rect 1663 573 1667 574
rect 1687 578 1691 579
rect 1687 573 1691 574
rect 1791 578 1795 579
rect 1791 573 1795 574
rect 800 549 802 573
rect 992 549 994 573
rect 1176 549 1178 573
rect 1352 549 1354 573
rect 1520 549 1522 573
rect 1688 549 1690 573
rect 798 548 804 549
rect 798 544 799 548
rect 803 544 804 548
rect 798 543 804 544
rect 990 548 996 549
rect 990 544 991 548
rect 995 544 996 548
rect 990 543 996 544
rect 1174 548 1180 549
rect 1174 544 1175 548
rect 1179 544 1180 548
rect 1174 543 1180 544
rect 1350 548 1356 549
rect 1350 544 1351 548
rect 1355 544 1356 548
rect 1350 543 1356 544
rect 1518 548 1524 549
rect 1518 544 1519 548
rect 1523 544 1524 548
rect 1518 543 1524 544
rect 1686 548 1692 549
rect 1686 544 1687 548
rect 1691 544 1692 548
rect 1686 543 1692 544
rect 1820 540 1822 646
rect 1868 624 1870 646
rect 1904 632 1906 653
rect 1978 647 1984 648
rect 1978 643 1979 647
rect 1983 643 1984 647
rect 1978 642 1984 643
rect 1902 631 1908 632
rect 1902 627 1903 631
rect 1907 627 1908 631
rect 1902 626 1908 627
rect 1980 624 1982 642
rect 2008 633 2010 653
rect 2047 649 2051 650
rect 2071 654 2075 655
rect 2071 649 2075 650
rect 2183 654 2187 655
rect 2183 649 2187 650
rect 2239 654 2243 655
rect 2239 649 2243 650
rect 2335 654 2339 655
rect 2335 649 2339 650
rect 2423 654 2427 655
rect 2423 649 2427 650
rect 2487 654 2491 655
rect 2487 649 2491 650
rect 2623 654 2627 655
rect 2623 649 2627 650
rect 2639 654 2643 655
rect 2639 649 2643 650
rect 2807 654 2811 655
rect 2807 649 2811 650
rect 2839 654 2843 655
rect 2839 649 2843 650
rect 2983 654 2987 655
rect 2983 649 2987 650
rect 3071 654 3075 655
rect 3071 649 3075 650
rect 3167 654 3171 655
rect 3167 649 3171 650
rect 2006 632 2012 633
rect 2006 628 2007 632
rect 2011 628 2012 632
rect 2048 629 2050 649
rect 2006 627 2012 628
rect 2046 628 2052 629
rect 2072 628 2074 649
rect 2146 647 2152 648
rect 2146 643 2147 647
rect 2151 643 2152 647
rect 2146 642 2152 643
rect 2046 624 2047 628
rect 2051 624 2052 628
rect 1866 623 1872 624
rect 1866 619 1867 623
rect 1871 619 1872 623
rect 1866 618 1872 619
rect 1978 623 1984 624
rect 2046 623 2052 624
rect 2070 627 2076 628
rect 2070 623 2071 627
rect 2075 623 2076 627
rect 1978 619 1979 623
rect 1983 619 1984 623
rect 2070 622 2076 623
rect 2148 620 2150 642
rect 2240 628 2242 649
rect 2314 647 2320 648
rect 2314 643 2315 647
rect 2319 643 2320 647
rect 2314 642 2320 643
rect 2238 627 2244 628
rect 2238 623 2239 627
rect 2243 623 2244 627
rect 2238 622 2244 623
rect 2316 620 2318 642
rect 2424 628 2426 649
rect 2624 628 2626 649
rect 2762 647 2768 648
rect 2762 643 2763 647
rect 2767 643 2768 647
rect 2762 642 2768 643
rect 2422 627 2428 628
rect 2422 623 2423 627
rect 2427 623 2428 627
rect 2422 622 2428 623
rect 2622 627 2628 628
rect 2622 623 2623 627
rect 2627 623 2628 627
rect 2622 622 2628 623
rect 2764 620 2766 642
rect 2840 628 2842 649
rect 2922 647 2928 648
rect 2922 643 2923 647
rect 2927 643 2928 647
rect 2922 642 2928 643
rect 2838 627 2844 628
rect 2838 623 2839 627
rect 2843 623 2844 627
rect 2838 622 2844 623
rect 2924 620 2926 642
rect 3072 628 3074 649
rect 3244 648 3246 698
rect 3320 680 3322 698
rect 3366 693 3372 694
rect 3366 689 3367 693
rect 3371 689 3372 693
rect 3366 688 3372 689
rect 3318 679 3324 680
rect 3318 675 3319 679
rect 3323 675 3324 679
rect 3318 674 3324 675
rect 3368 655 3370 688
rect 3452 672 3454 698
rect 3468 676 3470 778
rect 3542 776 3548 777
rect 3542 772 3543 776
rect 3547 772 3548 776
rect 3542 771 3548 772
rect 3702 776 3708 777
rect 3702 772 3703 776
rect 3707 772 3708 776
rect 3702 771 3708 772
rect 3544 743 3546 771
rect 3704 743 3706 771
rect 3543 742 3547 743
rect 3543 737 3547 738
rect 3575 742 3579 743
rect 3575 737 3579 738
rect 3703 742 3707 743
rect 3703 737 3707 738
rect 3576 713 3578 737
rect 3574 712 3580 713
rect 3574 708 3575 712
rect 3579 708 3580 712
rect 3574 707 3580 708
rect 3772 704 3774 810
rect 3840 796 3842 817
rect 3908 816 3910 858
rect 3916 832 3918 938
rect 3942 935 3943 939
rect 3947 935 3948 939
rect 3942 934 3948 935
rect 3944 903 3946 934
rect 3943 902 3947 903
rect 3943 897 3947 898
rect 3944 870 3946 897
rect 3942 869 3948 870
rect 3942 865 3943 869
rect 3947 865 3948 869
rect 3942 864 3948 865
rect 3942 852 3948 853
rect 3942 848 3943 852
rect 3947 848 3948 852
rect 3942 847 3948 848
rect 3914 831 3920 832
rect 3914 827 3915 831
rect 3919 827 3920 831
rect 3914 826 3920 827
rect 3944 823 3946 847
rect 3943 822 3947 823
rect 3943 817 3947 818
rect 3906 815 3912 816
rect 3906 811 3907 815
rect 3911 811 3912 815
rect 3906 810 3912 811
rect 3944 797 3946 817
rect 3942 796 3948 797
rect 3838 795 3844 796
rect 3838 791 3839 795
rect 3843 791 3844 795
rect 3942 792 3943 796
rect 3947 792 3948 796
rect 3942 791 3948 792
rect 3838 790 3844 791
rect 3914 783 3920 784
rect 3914 779 3915 783
rect 3919 779 3920 783
rect 3914 778 3920 779
rect 3942 779 3948 780
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3838 771 3844 772
rect 3840 743 3842 771
rect 3783 742 3787 743
rect 3783 737 3787 738
rect 3839 742 3843 743
rect 3839 737 3843 738
rect 3784 713 3786 737
rect 3782 712 3788 713
rect 3782 708 3783 712
rect 3787 708 3788 712
rect 3782 707 3788 708
rect 3770 703 3776 704
rect 3770 699 3771 703
rect 3775 699 3776 703
rect 3770 698 3776 699
rect 3574 693 3580 694
rect 3574 689 3575 693
rect 3579 689 3580 693
rect 3574 688 3580 689
rect 3782 693 3788 694
rect 3782 689 3783 693
rect 3787 689 3788 693
rect 3782 688 3788 689
rect 3466 675 3472 676
rect 3450 671 3456 672
rect 3450 667 3451 671
rect 3455 667 3456 671
rect 3466 671 3467 675
rect 3471 671 3472 675
rect 3466 670 3472 671
rect 3450 666 3456 667
rect 3576 655 3578 688
rect 3784 655 3786 688
rect 3874 671 3880 672
rect 3874 667 3875 671
rect 3879 667 3880 671
rect 3874 666 3880 667
rect 3319 654 3323 655
rect 3319 649 3323 650
rect 3367 654 3371 655
rect 3367 649 3371 650
rect 3575 654 3579 655
rect 3575 649 3579 650
rect 3783 654 3787 655
rect 3783 649 3787 650
rect 3839 654 3843 655
rect 3839 649 3843 650
rect 3242 647 3248 648
rect 3242 643 3243 647
rect 3247 643 3248 647
rect 3242 642 3248 643
rect 3320 628 3322 649
rect 3394 647 3400 648
rect 3394 643 3395 647
rect 3399 643 3400 647
rect 3394 642 3400 643
rect 3070 627 3076 628
rect 3070 623 3071 627
rect 3075 623 3076 627
rect 3070 622 3076 623
rect 3318 627 3324 628
rect 3318 623 3319 627
rect 3323 623 3324 627
rect 3318 622 3324 623
rect 3396 620 3398 642
rect 3402 639 3408 640
rect 3402 635 3403 639
rect 3407 635 3408 639
rect 3402 634 3408 635
rect 3404 620 3406 634
rect 3576 628 3578 649
rect 3840 628 3842 649
rect 3574 627 3580 628
rect 3574 623 3575 627
rect 3579 623 3580 627
rect 3574 622 3580 623
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3838 622 3844 623
rect 1978 618 1984 619
rect 2146 619 2152 620
rect 2006 615 2012 616
rect 1902 612 1908 613
rect 1902 608 1903 612
rect 1907 608 1908 612
rect 2006 611 2007 615
rect 2011 611 2012 615
rect 2146 615 2147 619
rect 2151 615 2152 619
rect 2146 614 2152 615
rect 2314 619 2320 620
rect 2314 615 2315 619
rect 2319 615 2320 619
rect 2314 614 2320 615
rect 2322 619 2328 620
rect 2322 615 2323 619
rect 2327 615 2328 619
rect 2762 619 2768 620
rect 2322 614 2328 615
rect 2698 615 2704 616
rect 2006 610 2012 611
rect 2046 611 2052 612
rect 1902 607 1908 608
rect 1904 579 1906 607
rect 2008 579 2010 610
rect 2046 607 2047 611
rect 2051 607 2052 611
rect 2046 606 2052 607
rect 2070 608 2076 609
rect 2048 579 2050 606
rect 2070 604 2071 608
rect 2075 604 2076 608
rect 2070 603 2076 604
rect 2238 608 2244 609
rect 2238 604 2239 608
rect 2243 604 2244 608
rect 2238 603 2244 604
rect 2072 579 2074 603
rect 2240 579 2242 603
rect 1863 578 1867 579
rect 1863 573 1867 574
rect 1903 578 1907 579
rect 1903 573 1907 574
rect 2007 578 2011 579
rect 2007 573 2011 574
rect 2047 578 2051 579
rect 2047 573 2051 574
rect 2071 578 2075 579
rect 2071 573 2075 574
rect 2191 578 2195 579
rect 2191 573 2195 574
rect 2239 578 2243 579
rect 2239 573 2243 574
rect 2287 578 2291 579
rect 2287 573 2291 574
rect 1864 549 1866 573
rect 1862 548 1868 549
rect 1862 544 1863 548
rect 1867 544 1868 548
rect 2008 546 2010 573
rect 2048 546 2050 573
rect 2192 549 2194 573
rect 2288 549 2290 573
rect 2190 548 2196 549
rect 1862 543 1868 544
rect 2006 545 2012 546
rect 2006 541 2007 545
rect 2011 541 2012 545
rect 2006 540 2012 541
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2190 544 2191 548
rect 2195 544 2196 548
rect 2190 543 2196 544
rect 2286 548 2292 549
rect 2286 544 2287 548
rect 2291 544 2292 548
rect 2286 543 2292 544
rect 2046 540 2052 541
rect 754 539 760 540
rect 754 535 755 539
rect 759 535 760 539
rect 754 534 760 535
rect 874 539 880 540
rect 874 535 875 539
rect 879 535 880 539
rect 874 534 880 535
rect 882 539 888 540
rect 882 535 883 539
rect 887 535 888 539
rect 882 534 888 535
rect 1250 539 1256 540
rect 1250 535 1251 539
rect 1255 535 1256 539
rect 1250 534 1256 535
rect 1426 539 1432 540
rect 1426 535 1427 539
rect 1431 535 1432 539
rect 1426 534 1432 535
rect 1594 539 1600 540
rect 1594 535 1595 539
rect 1599 535 1600 539
rect 1594 534 1600 535
rect 1762 539 1768 540
rect 1762 535 1763 539
rect 1767 535 1768 539
rect 1762 534 1768 535
rect 1818 539 1824 540
rect 1818 535 1819 539
rect 1823 535 1824 539
rect 1818 534 1824 535
rect 2266 539 2272 540
rect 2266 535 2267 539
rect 2271 535 2272 539
rect 2266 534 2272 535
rect 756 508 758 534
rect 798 529 804 530
rect 798 525 799 529
rect 803 525 804 529
rect 798 524 804 525
rect 690 507 696 508
rect 690 503 691 507
rect 695 503 696 507
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 135 497 139 498
rect 239 502 243 503
rect 239 497 243 498
rect 287 502 291 503
rect 370 502 376 503
rect 415 502 419 503
rect 287 497 291 498
rect 415 497 419 498
rect 463 502 467 503
rect 538 502 544 503
rect 607 502 611 503
rect 463 497 467 498
rect 112 477 114 497
rect 110 476 116 477
rect 136 476 138 497
rect 202 495 208 496
rect 202 491 203 495
rect 207 491 208 495
rect 202 490 208 491
rect 210 495 216 496
rect 210 491 211 495
rect 215 491 216 495
rect 210 490 216 491
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 134 475 140 476
rect 134 471 135 475
rect 139 471 140 475
rect 134 470 140 471
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 110 454 116 455
rect 134 456 140 457
rect 112 423 114 454
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 136 423 138 451
rect 111 422 115 423
rect 111 417 115 418
rect 135 422 139 423
rect 135 417 139 418
rect 112 390 114 417
rect 136 393 138 417
rect 134 392 140 393
rect 110 389 116 390
rect 110 385 111 389
rect 115 385 116 389
rect 134 388 135 392
rect 139 388 140 392
rect 134 387 140 388
rect 110 384 116 385
rect 204 384 206 490
rect 212 468 214 490
rect 288 476 290 497
rect 362 495 368 496
rect 362 491 363 495
rect 367 491 368 495
rect 362 490 368 491
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 364 468 366 490
rect 464 476 466 497
rect 462 475 468 476
rect 462 471 463 475
rect 467 471 468 475
rect 462 470 468 471
rect 540 468 542 502
rect 607 497 611 498
rect 639 502 643 503
rect 690 502 696 503
rect 754 507 760 508
rect 754 503 755 507
rect 759 503 760 507
rect 800 503 802 524
rect 876 508 878 534
rect 874 507 880 508
rect 874 503 875 507
rect 879 503 880 507
rect 754 502 760 503
rect 799 502 803 503
rect 639 497 643 498
rect 799 497 803 498
rect 807 502 811 503
rect 874 502 880 503
rect 807 497 811 498
rect 640 476 642 497
rect 808 476 810 497
rect 884 496 886 534
rect 990 529 996 530
rect 990 525 991 529
rect 995 525 996 529
rect 990 524 996 525
rect 1174 529 1180 530
rect 1174 525 1175 529
rect 1179 525 1180 529
rect 1174 524 1180 525
rect 992 503 994 524
rect 1176 503 1178 524
rect 1252 508 1254 534
rect 1350 529 1356 530
rect 1350 525 1351 529
rect 1355 525 1356 529
rect 1350 524 1356 525
rect 1250 507 1256 508
rect 1250 503 1251 507
rect 1255 503 1256 507
rect 1352 503 1354 524
rect 1428 508 1430 534
rect 1518 529 1524 530
rect 1518 525 1519 529
rect 1523 525 1524 529
rect 1518 524 1524 525
rect 1426 507 1432 508
rect 1426 503 1427 507
rect 1431 503 1432 507
rect 1520 503 1522 524
rect 1596 508 1598 534
rect 1686 529 1692 530
rect 1686 525 1687 529
rect 1691 525 1692 529
rect 1686 524 1692 525
rect 1594 507 1600 508
rect 1594 503 1595 507
rect 1599 503 1600 507
rect 1688 503 1690 524
rect 1764 508 1766 534
rect 1862 529 1868 530
rect 2190 529 2196 530
rect 1862 525 1863 529
rect 1867 525 1868 529
rect 1862 524 1868 525
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 1762 507 1768 508
rect 1762 503 1763 507
rect 1767 503 1768 507
rect 1864 503 1866 524
rect 2006 523 2012 524
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2190 525 2191 529
rect 2195 525 2196 529
rect 2190 524 2196 525
rect 2046 523 2052 524
rect 2008 503 2010 523
rect 2048 503 2050 523
rect 2192 503 2194 524
rect 2268 508 2270 534
rect 2286 529 2292 530
rect 2286 525 2287 529
rect 2291 525 2292 529
rect 2286 524 2292 525
rect 2266 507 2272 508
rect 2266 503 2267 507
rect 2271 503 2272 507
rect 2288 503 2290 524
rect 2324 516 2326 614
rect 2698 611 2699 615
rect 2703 611 2704 615
rect 2762 615 2763 619
rect 2767 615 2768 619
rect 2762 614 2768 615
rect 2922 619 2928 620
rect 2922 615 2923 619
rect 2927 615 2928 619
rect 2922 614 2928 615
rect 3394 619 3400 620
rect 3394 615 3395 619
rect 3399 615 3400 619
rect 3394 614 3400 615
rect 3402 619 3408 620
rect 3402 615 3403 619
rect 3407 615 3408 619
rect 3402 614 3408 615
rect 2698 610 2704 611
rect 2422 608 2428 609
rect 2422 604 2423 608
rect 2427 604 2428 608
rect 2422 603 2428 604
rect 2622 608 2628 609
rect 2622 604 2623 608
rect 2627 604 2628 608
rect 2622 603 2628 604
rect 2424 579 2426 603
rect 2624 579 2626 603
rect 2383 578 2387 579
rect 2383 573 2387 574
rect 2423 578 2427 579
rect 2423 573 2427 574
rect 2479 578 2483 579
rect 2479 573 2483 574
rect 2583 578 2587 579
rect 2583 573 2587 574
rect 2623 578 2627 579
rect 2623 573 2627 574
rect 2384 549 2386 573
rect 2480 549 2482 573
rect 2584 549 2586 573
rect 2382 548 2388 549
rect 2382 544 2383 548
rect 2387 544 2388 548
rect 2382 543 2388 544
rect 2478 548 2484 549
rect 2478 544 2479 548
rect 2483 544 2484 548
rect 2478 543 2484 544
rect 2582 548 2588 549
rect 2582 544 2583 548
rect 2587 544 2588 548
rect 2582 543 2588 544
rect 2362 539 2368 540
rect 2362 535 2363 539
rect 2367 535 2368 539
rect 2362 534 2368 535
rect 2458 539 2464 540
rect 2458 535 2459 539
rect 2463 535 2464 539
rect 2458 534 2464 535
rect 2554 539 2560 540
rect 2554 535 2555 539
rect 2559 535 2560 539
rect 2554 534 2560 535
rect 2562 539 2568 540
rect 2562 535 2563 539
rect 2567 535 2568 539
rect 2562 534 2568 535
rect 2322 515 2328 516
rect 2322 511 2323 515
rect 2327 511 2328 515
rect 2322 510 2328 511
rect 2364 508 2366 534
rect 2382 529 2388 530
rect 2382 525 2383 529
rect 2387 525 2388 529
rect 2382 524 2388 525
rect 2362 507 2368 508
rect 2362 503 2363 507
rect 2367 503 2368 507
rect 2384 503 2386 524
rect 2460 508 2462 534
rect 2478 529 2484 530
rect 2478 525 2479 529
rect 2483 525 2484 529
rect 2478 524 2484 525
rect 2458 507 2464 508
rect 2458 503 2459 507
rect 2463 503 2464 507
rect 2480 503 2482 524
rect 2556 508 2558 534
rect 2554 507 2560 508
rect 2554 503 2555 507
rect 2559 503 2560 507
rect 967 502 971 503
rect 967 497 971 498
rect 991 502 995 503
rect 991 497 995 498
rect 1119 502 1123 503
rect 1119 497 1123 498
rect 1175 502 1179 503
rect 1250 502 1256 503
rect 1271 502 1275 503
rect 1175 497 1179 498
rect 1271 497 1275 498
rect 1351 502 1355 503
rect 1351 497 1355 498
rect 1415 502 1419 503
rect 1426 502 1432 503
rect 1519 502 1523 503
rect 1415 497 1419 498
rect 1519 497 1523 498
rect 1567 502 1571 503
rect 1594 502 1600 503
rect 1687 502 1691 503
rect 1762 502 1768 503
rect 1863 502 1867 503
rect 1567 497 1571 498
rect 1687 497 1691 498
rect 1863 497 1867 498
rect 2007 502 2011 503
rect 2007 497 2011 498
rect 2047 502 2051 503
rect 2047 497 2051 498
rect 2191 502 2195 503
rect 2266 502 2272 503
rect 2287 502 2291 503
rect 2362 502 2368 503
rect 2383 502 2387 503
rect 2191 497 2195 498
rect 2287 497 2291 498
rect 2383 497 2387 498
rect 2431 502 2435 503
rect 2458 502 2464 503
rect 2479 502 2483 503
rect 2431 497 2435 498
rect 2479 497 2483 498
rect 2527 502 2531 503
rect 2554 502 2560 503
rect 2527 497 2531 498
rect 882 495 888 496
rect 882 491 883 495
rect 887 491 888 495
rect 882 490 888 491
rect 968 476 970 497
rect 1102 495 1108 496
rect 1102 491 1103 495
rect 1107 491 1108 495
rect 1102 490 1108 491
rect 638 475 644 476
rect 638 471 639 475
rect 643 471 644 475
rect 638 470 644 471
rect 806 475 812 476
rect 806 471 807 475
rect 811 471 812 475
rect 806 470 812 471
rect 966 475 972 476
rect 966 471 967 475
rect 971 471 972 475
rect 966 470 972 471
rect 1104 468 1106 490
rect 1120 476 1122 497
rect 1194 495 1200 496
rect 1194 491 1195 495
rect 1199 491 1200 495
rect 1194 490 1200 491
rect 1118 475 1124 476
rect 1118 471 1119 475
rect 1123 471 1124 475
rect 1118 470 1124 471
rect 1196 468 1198 490
rect 1272 476 1274 497
rect 1394 495 1400 496
rect 1394 491 1395 495
rect 1399 491 1400 495
rect 1394 490 1400 491
rect 1290 487 1296 488
rect 1290 483 1291 487
rect 1295 483 1296 487
rect 1290 482 1296 483
rect 1270 475 1276 476
rect 1270 471 1271 475
rect 1275 471 1276 475
rect 1270 470 1276 471
rect 210 467 216 468
rect 210 463 211 467
rect 215 463 216 467
rect 210 462 216 463
rect 362 467 368 468
rect 362 463 363 467
rect 367 463 368 467
rect 362 462 368 463
rect 538 467 544 468
rect 538 463 539 467
rect 543 463 544 467
rect 538 462 544 463
rect 546 467 552 468
rect 546 463 547 467
rect 551 463 552 467
rect 546 462 552 463
rect 1102 467 1108 468
rect 1102 463 1103 467
rect 1107 463 1108 467
rect 1102 462 1108 463
rect 1194 467 1200 468
rect 1194 463 1195 467
rect 1199 463 1200 467
rect 1194 462 1200 463
rect 286 456 292 457
rect 286 452 287 456
rect 291 452 292 456
rect 286 451 292 452
rect 462 456 468 457
rect 462 452 463 456
rect 467 452 468 456
rect 462 451 468 452
rect 288 423 290 451
rect 464 423 466 451
rect 279 422 283 423
rect 279 417 283 418
rect 287 422 291 423
rect 287 417 291 418
rect 439 422 443 423
rect 439 417 443 418
rect 463 422 467 423
rect 463 417 467 418
rect 280 393 282 417
rect 440 393 442 417
rect 278 392 284 393
rect 278 388 279 392
rect 283 388 284 392
rect 278 387 284 388
rect 438 392 444 393
rect 438 388 439 392
rect 443 388 444 392
rect 438 387 444 388
rect 202 383 208 384
rect 202 379 203 383
rect 207 379 208 383
rect 202 378 208 379
rect 514 383 520 384
rect 514 379 515 383
rect 519 379 520 383
rect 514 378 520 379
rect 202 375 208 376
rect 134 373 140 374
rect 110 372 116 373
rect 110 368 111 372
rect 115 368 116 372
rect 134 369 135 373
rect 139 369 140 373
rect 202 371 203 375
rect 207 371 208 375
rect 202 370 208 371
rect 278 373 284 374
rect 134 368 140 369
rect 110 367 116 368
rect 112 347 114 367
rect 136 347 138 368
rect 204 352 206 370
rect 278 369 279 373
rect 283 369 284 373
rect 278 368 284 369
rect 438 373 444 374
rect 438 369 439 373
rect 443 369 444 373
rect 438 368 444 369
rect 202 351 208 352
rect 202 347 203 351
rect 207 347 208 351
rect 111 346 115 347
rect 111 341 115 342
rect 135 346 139 347
rect 135 341 139 342
rect 143 346 147 347
rect 202 346 208 347
rect 218 351 224 352
rect 218 347 219 351
rect 223 347 224 351
rect 280 347 282 368
rect 440 347 442 368
rect 516 352 518 378
rect 548 360 550 462
rect 638 456 644 457
rect 638 452 639 456
rect 643 452 644 456
rect 638 451 644 452
rect 806 456 812 457
rect 806 452 807 456
rect 811 452 812 456
rect 806 451 812 452
rect 966 456 972 457
rect 966 452 967 456
rect 971 452 972 456
rect 966 451 972 452
rect 1118 456 1124 457
rect 1118 452 1119 456
rect 1123 452 1124 456
rect 1118 451 1124 452
rect 1270 456 1276 457
rect 1270 452 1271 456
rect 1275 452 1276 456
rect 1270 451 1276 452
rect 640 423 642 451
rect 808 423 810 451
rect 968 423 970 451
rect 1120 423 1122 451
rect 1272 423 1274 451
rect 583 422 587 423
rect 583 417 587 418
rect 639 422 643 423
rect 639 417 643 418
rect 719 422 723 423
rect 719 417 723 418
rect 807 422 811 423
rect 807 417 811 418
rect 847 422 851 423
rect 847 417 851 418
rect 967 422 971 423
rect 967 417 971 418
rect 1087 422 1091 423
rect 1087 417 1091 418
rect 1119 422 1123 423
rect 1119 417 1123 418
rect 1207 422 1211 423
rect 1207 417 1211 418
rect 1271 422 1275 423
rect 1271 417 1275 418
rect 584 393 586 417
rect 720 393 722 417
rect 848 393 850 417
rect 968 393 970 417
rect 1088 393 1090 417
rect 1208 393 1210 417
rect 582 392 588 393
rect 582 388 583 392
rect 587 388 588 392
rect 582 387 588 388
rect 718 392 724 393
rect 718 388 719 392
rect 723 388 724 392
rect 718 387 724 388
rect 846 392 852 393
rect 846 388 847 392
rect 851 388 852 392
rect 846 387 852 388
rect 966 392 972 393
rect 966 388 967 392
rect 971 388 972 392
rect 966 387 972 388
rect 1086 392 1092 393
rect 1086 388 1087 392
rect 1091 388 1092 392
rect 1086 387 1092 388
rect 1206 392 1212 393
rect 1206 388 1207 392
rect 1211 388 1212 392
rect 1206 387 1212 388
rect 1292 384 1294 482
rect 1396 468 1398 490
rect 1416 476 1418 497
rect 1490 495 1496 496
rect 1490 491 1491 495
rect 1495 491 1496 495
rect 1490 490 1496 491
rect 1414 475 1420 476
rect 1414 471 1415 475
rect 1419 471 1420 475
rect 1414 470 1420 471
rect 1492 468 1494 490
rect 1568 476 1570 497
rect 2008 477 2010 497
rect 2048 477 2050 497
rect 2006 476 2012 477
rect 1566 475 1572 476
rect 1566 471 1567 475
rect 1571 471 1572 475
rect 2006 472 2007 476
rect 2011 472 2012 476
rect 2006 471 2012 472
rect 2046 476 2052 477
rect 2432 476 2434 497
rect 2506 495 2512 496
rect 2506 491 2507 495
rect 2511 491 2512 495
rect 2506 490 2512 491
rect 2046 472 2047 476
rect 2051 472 2052 476
rect 2046 471 2052 472
rect 2430 475 2436 476
rect 2430 471 2431 475
rect 2435 471 2436 475
rect 1566 470 1572 471
rect 2430 470 2436 471
rect 2508 468 2510 490
rect 2528 476 2530 497
rect 2564 488 2566 534
rect 2582 529 2588 530
rect 2582 525 2583 529
rect 2587 525 2588 529
rect 2582 524 2588 525
rect 2584 503 2586 524
rect 2700 508 2702 610
rect 2838 608 2844 609
rect 2838 604 2839 608
rect 2843 604 2844 608
rect 2838 603 2844 604
rect 3070 608 3076 609
rect 3070 604 3071 608
rect 3075 604 3076 608
rect 3070 603 3076 604
rect 3318 608 3324 609
rect 3318 604 3319 608
rect 3323 604 3324 608
rect 3318 603 3324 604
rect 3574 608 3580 609
rect 3574 604 3575 608
rect 3579 604 3580 608
rect 3574 603 3580 604
rect 3838 608 3844 609
rect 3838 604 3839 608
rect 3843 604 3844 608
rect 3838 603 3844 604
rect 2840 579 2842 603
rect 3072 579 3074 603
rect 3320 579 3322 603
rect 3576 579 3578 603
rect 3840 579 3842 603
rect 2711 578 2715 579
rect 2711 573 2715 574
rect 2839 578 2843 579
rect 2839 573 2843 574
rect 2871 578 2875 579
rect 2871 573 2875 574
rect 3071 578 3075 579
rect 3071 573 3075 574
rect 3303 578 3307 579
rect 3303 573 3307 574
rect 3319 578 3323 579
rect 3319 573 3323 574
rect 3551 578 3555 579
rect 3551 573 3555 574
rect 3575 578 3579 579
rect 3575 573 3579 574
rect 3807 578 3811 579
rect 3807 573 3811 574
rect 3839 578 3843 579
rect 3839 573 3843 574
rect 2712 549 2714 573
rect 2872 549 2874 573
rect 3072 549 3074 573
rect 3304 549 3306 573
rect 3552 549 3554 573
rect 3808 549 3810 573
rect 2710 548 2716 549
rect 2710 544 2711 548
rect 2715 544 2716 548
rect 2710 543 2716 544
rect 2870 548 2876 549
rect 2870 544 2871 548
rect 2875 544 2876 548
rect 2870 543 2876 544
rect 3070 548 3076 549
rect 3070 544 3071 548
rect 3075 544 3076 548
rect 3070 543 3076 544
rect 3302 548 3308 549
rect 3302 544 3303 548
rect 3307 544 3308 548
rect 3302 543 3308 544
rect 3550 548 3556 549
rect 3550 544 3551 548
rect 3555 544 3556 548
rect 3550 543 3556 544
rect 3806 548 3812 549
rect 3806 544 3807 548
rect 3811 544 3812 548
rect 3806 543 3812 544
rect 3876 540 3878 666
rect 3916 648 3918 778
rect 3942 775 3943 779
rect 3947 775 3948 779
rect 3942 774 3948 775
rect 3944 743 3946 774
rect 3943 742 3947 743
rect 3943 737 3947 738
rect 3944 710 3946 737
rect 3942 709 3948 710
rect 3942 705 3943 709
rect 3947 705 3948 709
rect 3942 704 3948 705
rect 3942 692 3948 693
rect 3942 688 3943 692
rect 3947 688 3948 692
rect 3942 687 3948 688
rect 3944 655 3946 687
rect 3943 654 3947 655
rect 3943 649 3947 650
rect 3914 647 3920 648
rect 3914 643 3915 647
rect 3919 643 3920 647
rect 3914 642 3920 643
rect 3944 629 3946 649
rect 3942 628 3948 629
rect 3942 624 3943 628
rect 3947 624 3948 628
rect 3942 623 3948 624
rect 3914 615 3920 616
rect 3914 611 3915 615
rect 3919 611 3920 615
rect 3914 610 3920 611
rect 3942 611 3948 612
rect 2786 539 2792 540
rect 2786 535 2787 539
rect 2791 535 2792 539
rect 2786 534 2792 535
rect 2946 539 2952 540
rect 2946 535 2947 539
rect 2951 535 2952 539
rect 2946 534 2952 535
rect 3146 539 3152 540
rect 3146 535 3147 539
rect 3151 535 3152 539
rect 3146 534 3152 535
rect 3478 539 3484 540
rect 3478 535 3479 539
rect 3483 535 3484 539
rect 3478 534 3484 535
rect 3626 539 3632 540
rect 3626 535 3627 539
rect 3631 535 3632 539
rect 3626 534 3632 535
rect 3874 539 3880 540
rect 3874 535 3875 539
rect 3879 535 3880 539
rect 3874 534 3880 535
rect 2710 529 2716 530
rect 2710 525 2711 529
rect 2715 525 2716 529
rect 2710 524 2716 525
rect 2698 507 2704 508
rect 2698 503 2699 507
rect 2703 503 2704 507
rect 2712 503 2714 524
rect 2788 508 2790 534
rect 2870 529 2876 530
rect 2870 525 2871 529
rect 2875 525 2876 529
rect 2870 524 2876 525
rect 2786 507 2792 508
rect 2786 503 2787 507
rect 2791 503 2792 507
rect 2872 503 2874 524
rect 2948 508 2950 534
rect 3070 529 3076 530
rect 3070 525 3071 529
rect 3075 525 3076 529
rect 3070 524 3076 525
rect 2946 507 2952 508
rect 2946 503 2947 507
rect 2951 503 2952 507
rect 3072 503 3074 524
rect 3148 508 3150 534
rect 3302 529 3308 530
rect 3302 525 3303 529
rect 3307 525 3308 529
rect 3302 524 3308 525
rect 3146 507 3152 508
rect 3146 503 3147 507
rect 3151 503 3152 507
rect 3304 503 3306 524
rect 3480 508 3482 534
rect 3550 529 3556 530
rect 3550 525 3551 529
rect 3555 525 3556 529
rect 3550 524 3556 525
rect 3478 507 3484 508
rect 3478 503 3479 507
rect 3483 503 3484 507
rect 3552 503 3554 524
rect 2583 502 2587 503
rect 2583 497 2587 498
rect 2623 502 2627 503
rect 2698 502 2704 503
rect 2711 502 2715 503
rect 2623 497 2627 498
rect 2711 497 2715 498
rect 2727 502 2731 503
rect 2786 502 2792 503
rect 2847 502 2851 503
rect 2727 497 2731 498
rect 2847 497 2851 498
rect 2871 502 2875 503
rect 2946 502 2952 503
rect 2999 502 3003 503
rect 2871 497 2875 498
rect 2999 497 3003 498
rect 3071 502 3075 503
rect 3146 502 3152 503
rect 3175 502 3179 503
rect 3071 497 3075 498
rect 3175 497 3179 498
rect 3303 502 3307 503
rect 3303 497 3307 498
rect 3375 502 3379 503
rect 3478 502 3484 503
rect 3551 502 3555 503
rect 3375 497 3379 498
rect 3551 497 3555 498
rect 3591 502 3595 503
rect 3591 497 3595 498
rect 2602 495 2608 496
rect 2602 491 2603 495
rect 2607 491 2608 495
rect 2602 490 2608 491
rect 2562 487 2568 488
rect 2562 483 2563 487
rect 2567 483 2568 487
rect 2562 482 2568 483
rect 2526 475 2532 476
rect 2526 471 2527 475
rect 2531 471 2532 475
rect 2526 470 2532 471
rect 2604 468 2606 490
rect 2624 476 2626 497
rect 2698 495 2704 496
rect 2698 491 2699 495
rect 2703 491 2704 495
rect 2698 490 2704 491
rect 2622 475 2628 476
rect 2622 471 2623 475
rect 2627 471 2628 475
rect 2622 470 2628 471
rect 2700 468 2702 490
rect 2728 476 2730 497
rect 2802 495 2808 496
rect 2802 491 2803 495
rect 2807 491 2808 495
rect 2802 490 2808 491
rect 2726 475 2732 476
rect 2726 471 2727 475
rect 2731 471 2732 475
rect 2726 470 2732 471
rect 2804 468 2806 490
rect 2848 476 2850 497
rect 2922 495 2928 496
rect 2922 491 2923 495
rect 2927 491 2928 495
rect 2922 490 2928 491
rect 2846 475 2852 476
rect 2846 471 2847 475
rect 2851 471 2852 475
rect 2846 470 2852 471
rect 2924 468 2926 490
rect 3000 476 3002 497
rect 3176 476 3178 497
rect 3258 495 3264 496
rect 3258 491 3259 495
rect 3263 491 3264 495
rect 3258 490 3264 491
rect 2998 475 3004 476
rect 2998 471 2999 475
rect 3003 471 3004 475
rect 2998 470 3004 471
rect 3174 475 3180 476
rect 3174 471 3175 475
rect 3179 471 3180 475
rect 3174 470 3180 471
rect 3260 468 3262 490
rect 3376 476 3378 497
rect 3458 495 3464 496
rect 3458 491 3459 495
rect 3463 491 3464 495
rect 3458 490 3464 491
rect 3374 475 3380 476
rect 3374 471 3375 475
rect 3379 471 3380 475
rect 3374 470 3380 471
rect 3460 468 3462 490
rect 3592 476 3594 497
rect 3628 496 3630 534
rect 3806 529 3812 530
rect 3806 525 3807 529
rect 3811 525 3812 529
rect 3806 524 3812 525
rect 3808 503 3810 524
rect 3916 508 3918 610
rect 3942 607 3943 611
rect 3947 607 3948 611
rect 3942 606 3948 607
rect 3944 579 3946 606
rect 3943 578 3947 579
rect 3943 573 3947 574
rect 3944 546 3946 573
rect 3942 545 3948 546
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 3942 523 3948 524
rect 3914 507 3920 508
rect 3914 503 3915 507
rect 3919 503 3920 507
rect 3944 503 3946 523
rect 3807 502 3811 503
rect 3914 502 3920 503
rect 3943 502 3947 503
rect 3807 497 3811 498
rect 3943 497 3947 498
rect 3626 495 3632 496
rect 3626 491 3627 495
rect 3631 491 3632 495
rect 3626 490 3632 491
rect 3808 476 3810 497
rect 3858 495 3864 496
rect 3858 491 3859 495
rect 3863 491 3864 495
rect 3858 490 3864 491
rect 3590 475 3596 476
rect 3590 471 3591 475
rect 3595 471 3596 475
rect 3590 470 3596 471
rect 3806 475 3812 476
rect 3806 471 3807 475
rect 3811 471 3812 475
rect 3806 470 3812 471
rect 1394 467 1400 468
rect 1394 463 1395 467
rect 1399 463 1400 467
rect 1394 462 1400 463
rect 1490 467 1496 468
rect 1490 463 1491 467
rect 1495 463 1496 467
rect 1490 462 1496 463
rect 2506 467 2512 468
rect 2506 463 2507 467
rect 2511 463 2512 467
rect 2506 462 2512 463
rect 2602 467 2608 468
rect 2602 463 2603 467
rect 2607 463 2608 467
rect 2602 462 2608 463
rect 2698 467 2704 468
rect 2698 463 2699 467
rect 2703 463 2704 467
rect 2698 462 2704 463
rect 2802 467 2808 468
rect 2802 463 2803 467
rect 2807 463 2808 467
rect 2802 462 2808 463
rect 2922 467 2928 468
rect 2922 463 2923 467
rect 2927 463 2928 467
rect 2922 462 2928 463
rect 2934 467 2940 468
rect 2934 463 2935 467
rect 2939 463 2940 467
rect 2934 462 2940 463
rect 3082 467 3088 468
rect 3082 463 3083 467
rect 3087 463 3088 467
rect 3082 462 3088 463
rect 3258 467 3264 468
rect 3258 463 3259 467
rect 3263 463 3264 467
rect 3258 462 3264 463
rect 3458 467 3464 468
rect 3458 463 3459 467
rect 3463 463 3464 467
rect 3458 462 3464 463
rect 2006 459 2012 460
rect 1414 456 1420 457
rect 1414 452 1415 456
rect 1419 452 1420 456
rect 1414 451 1420 452
rect 1566 456 1572 457
rect 1566 452 1567 456
rect 1571 452 1572 456
rect 2006 455 2007 459
rect 2011 455 2012 459
rect 2006 454 2012 455
rect 2046 459 2052 460
rect 2046 455 2047 459
rect 2051 455 2052 459
rect 2046 454 2052 455
rect 2430 456 2436 457
rect 1566 451 1572 452
rect 1416 423 1418 451
rect 1568 423 1570 451
rect 2008 423 2010 454
rect 2048 427 2050 454
rect 2430 452 2431 456
rect 2435 452 2436 456
rect 2430 451 2436 452
rect 2526 456 2532 457
rect 2526 452 2527 456
rect 2531 452 2532 456
rect 2526 451 2532 452
rect 2622 456 2628 457
rect 2622 452 2623 456
rect 2627 452 2628 456
rect 2622 451 2628 452
rect 2726 456 2732 457
rect 2726 452 2727 456
rect 2731 452 2732 456
rect 2726 451 2732 452
rect 2846 456 2852 457
rect 2846 452 2847 456
rect 2851 452 2852 456
rect 2846 451 2852 452
rect 2432 427 2434 451
rect 2528 427 2530 451
rect 2624 427 2626 451
rect 2728 427 2730 451
rect 2848 427 2850 451
rect 2047 426 2051 427
rect 1327 422 1331 423
rect 1327 417 1331 418
rect 1415 422 1419 423
rect 1415 417 1419 418
rect 1567 422 1571 423
rect 1567 417 1571 418
rect 2007 422 2011 423
rect 2047 421 2051 422
rect 2431 426 2435 427
rect 2431 421 2435 422
rect 2527 426 2531 427
rect 2527 421 2531 422
rect 2623 426 2627 427
rect 2623 421 2627 422
rect 2719 426 2723 427
rect 2719 421 2723 422
rect 2727 426 2731 427
rect 2727 421 2731 422
rect 2815 426 2819 427
rect 2815 421 2819 422
rect 2847 426 2851 427
rect 2847 421 2851 422
rect 2927 426 2931 427
rect 2927 421 2931 422
rect 2007 417 2011 418
rect 1328 393 1330 417
rect 1326 392 1332 393
rect 1326 388 1327 392
rect 1331 388 1332 392
rect 2008 390 2010 417
rect 2048 394 2050 421
rect 2432 397 2434 421
rect 2528 397 2530 421
rect 2624 397 2626 421
rect 2720 397 2722 421
rect 2816 397 2818 421
rect 2928 397 2930 421
rect 2430 396 2436 397
rect 2046 393 2052 394
rect 1326 387 1332 388
rect 2006 389 2012 390
rect 2006 385 2007 389
rect 2011 385 2012 389
rect 2046 389 2047 393
rect 2051 389 2052 393
rect 2430 392 2431 396
rect 2435 392 2436 396
rect 2430 391 2436 392
rect 2526 396 2532 397
rect 2526 392 2527 396
rect 2531 392 2532 396
rect 2526 391 2532 392
rect 2622 396 2628 397
rect 2622 392 2623 396
rect 2627 392 2628 396
rect 2622 391 2628 392
rect 2718 396 2724 397
rect 2718 392 2719 396
rect 2723 392 2724 396
rect 2718 391 2724 392
rect 2814 396 2820 397
rect 2814 392 2815 396
rect 2819 392 2820 396
rect 2814 391 2820 392
rect 2926 396 2932 397
rect 2926 392 2927 396
rect 2931 392 2932 396
rect 2926 391 2932 392
rect 2046 388 2052 389
rect 2006 384 2012 385
rect 2506 387 2512 388
rect 658 383 664 384
rect 658 379 659 383
rect 663 379 664 383
rect 658 378 664 379
rect 794 383 800 384
rect 794 379 795 383
rect 799 379 800 383
rect 794 378 800 379
rect 922 383 928 384
rect 922 379 923 383
rect 927 379 928 383
rect 922 378 928 379
rect 1042 383 1048 384
rect 1042 379 1043 383
rect 1047 379 1048 383
rect 1042 378 1048 379
rect 1162 383 1168 384
rect 1162 379 1163 383
rect 1167 379 1168 383
rect 1162 378 1168 379
rect 1282 383 1288 384
rect 1282 379 1283 383
rect 1287 379 1288 383
rect 1282 378 1288 379
rect 1290 383 1296 384
rect 1290 379 1291 383
rect 1295 379 1296 383
rect 2506 383 2507 387
rect 2511 383 2512 387
rect 2506 382 2512 383
rect 2602 387 2608 388
rect 2602 383 2603 387
rect 2607 383 2608 387
rect 2602 382 2608 383
rect 2610 387 2616 388
rect 2610 383 2611 387
rect 2615 383 2616 387
rect 2610 382 2616 383
rect 2706 387 2712 388
rect 2706 383 2707 387
rect 2711 383 2712 387
rect 2706 382 2712 383
rect 2802 387 2808 388
rect 2802 383 2803 387
rect 2807 383 2808 387
rect 2802 382 2808 383
rect 1290 378 1296 379
rect 582 373 588 374
rect 582 369 583 373
rect 587 369 588 373
rect 582 368 588 369
rect 546 359 552 360
rect 546 355 547 359
rect 551 355 552 359
rect 546 354 552 355
rect 514 351 520 352
rect 514 347 515 351
rect 519 347 520 351
rect 584 347 586 368
rect 660 352 662 378
rect 718 373 724 374
rect 718 369 719 373
rect 723 369 724 373
rect 718 368 724 369
rect 658 351 664 352
rect 658 347 659 351
rect 663 347 664 351
rect 720 347 722 368
rect 218 346 224 347
rect 279 346 283 347
rect 143 341 147 342
rect 112 321 114 341
rect 110 320 116 321
rect 144 320 146 341
rect 220 320 222 346
rect 279 341 283 342
rect 319 346 323 347
rect 319 341 323 342
rect 439 346 443 347
rect 439 341 443 342
rect 479 346 483 347
rect 514 346 520 347
rect 583 346 587 347
rect 479 341 483 342
rect 583 341 587 342
rect 631 346 635 347
rect 658 346 664 347
rect 719 346 723 347
rect 631 341 635 342
rect 719 341 723 342
rect 775 346 779 347
rect 775 341 779 342
rect 320 320 322 341
rect 480 320 482 341
rect 498 339 504 340
rect 498 335 499 339
rect 503 335 504 339
rect 498 334 504 335
rect 618 339 624 340
rect 618 335 619 339
rect 623 335 624 339
rect 618 334 624 335
rect 110 316 111 320
rect 115 316 116 320
rect 110 315 116 316
rect 142 319 148 320
rect 142 315 143 319
rect 147 315 148 319
rect 142 314 148 315
rect 218 319 224 320
rect 218 315 219 319
rect 223 315 224 319
rect 218 314 224 315
rect 318 319 324 320
rect 318 315 319 319
rect 323 315 324 319
rect 318 314 324 315
rect 478 319 484 320
rect 478 315 479 319
rect 483 315 484 319
rect 478 314 484 315
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 110 298 116 299
rect 142 300 148 301
rect 112 267 114 298
rect 142 296 143 300
rect 147 296 148 300
rect 142 295 148 296
rect 318 300 324 301
rect 318 296 319 300
rect 323 296 324 300
rect 318 295 324 296
rect 478 300 484 301
rect 478 296 479 300
rect 483 296 484 300
rect 478 295 484 296
rect 144 267 146 295
rect 320 267 322 295
rect 480 267 482 295
rect 111 266 115 267
rect 111 261 115 262
rect 143 266 147 267
rect 143 261 147 262
rect 223 266 227 267
rect 223 261 227 262
rect 319 266 323 267
rect 319 261 323 262
rect 391 266 395 267
rect 391 261 395 262
rect 479 266 483 267
rect 479 261 483 262
rect 112 234 114 261
rect 224 237 226 261
rect 392 237 394 261
rect 222 236 228 237
rect 110 233 116 234
rect 110 229 111 233
rect 115 229 116 233
rect 222 232 223 236
rect 227 232 228 236
rect 222 231 228 232
rect 390 236 396 237
rect 390 232 391 236
rect 395 232 396 236
rect 390 231 396 232
rect 110 228 116 229
rect 500 228 502 334
rect 620 312 622 334
rect 632 320 634 341
rect 746 331 752 332
rect 746 327 747 331
rect 751 327 752 331
rect 746 326 752 327
rect 630 319 636 320
rect 630 315 631 319
rect 635 315 636 319
rect 630 314 636 315
rect 748 312 750 326
rect 776 320 778 341
rect 796 340 798 378
rect 846 373 852 374
rect 846 369 847 373
rect 851 369 852 373
rect 846 368 852 369
rect 848 347 850 368
rect 924 352 926 378
rect 966 373 972 374
rect 966 369 967 373
rect 971 369 972 373
rect 966 368 972 369
rect 894 351 900 352
rect 894 347 895 351
rect 899 347 900 351
rect 922 351 928 352
rect 922 347 923 351
rect 927 347 928 351
rect 968 347 970 368
rect 1044 352 1046 378
rect 1086 373 1092 374
rect 1086 369 1087 373
rect 1091 369 1092 373
rect 1086 368 1092 369
rect 1042 351 1048 352
rect 1042 347 1043 351
rect 1047 347 1048 351
rect 1088 347 1090 368
rect 1164 352 1166 378
rect 1206 373 1212 374
rect 1206 369 1207 373
rect 1211 369 1212 373
rect 1206 368 1212 369
rect 1162 351 1168 352
rect 1162 347 1163 351
rect 1167 347 1168 351
rect 1208 347 1210 368
rect 1284 352 1286 378
rect 2430 377 2436 378
rect 2046 376 2052 377
rect 1326 373 1332 374
rect 1326 369 1327 373
rect 1331 369 1332 373
rect 1326 368 1332 369
rect 2006 372 2012 373
rect 2006 368 2007 372
rect 2011 368 2012 372
rect 2046 372 2047 376
rect 2051 372 2052 376
rect 2430 373 2431 377
rect 2435 373 2436 377
rect 2430 372 2436 373
rect 2046 371 2052 372
rect 1282 351 1288 352
rect 1282 347 1283 351
rect 1287 347 1288 351
rect 1328 347 1330 368
rect 2006 367 2012 368
rect 2008 347 2010 367
rect 2048 347 2050 371
rect 2432 347 2434 372
rect 2508 356 2510 382
rect 2526 377 2532 378
rect 2526 373 2527 377
rect 2531 373 2532 377
rect 2526 372 2532 373
rect 2506 355 2512 356
rect 2506 351 2507 355
rect 2511 351 2512 355
rect 2506 350 2512 351
rect 2528 347 2530 372
rect 2604 348 2606 382
rect 2612 364 2614 382
rect 2622 377 2628 378
rect 2622 373 2623 377
rect 2627 373 2628 377
rect 2622 372 2628 373
rect 2610 363 2616 364
rect 2610 359 2611 363
rect 2615 359 2616 363
rect 2610 358 2616 359
rect 2602 347 2608 348
rect 2624 347 2626 372
rect 2708 356 2710 382
rect 2718 377 2724 378
rect 2718 373 2719 377
rect 2723 373 2724 377
rect 2718 372 2724 373
rect 2706 355 2712 356
rect 2706 351 2707 355
rect 2711 351 2712 355
rect 2706 350 2712 351
rect 2720 347 2722 372
rect 2804 356 2806 382
rect 2814 377 2820 378
rect 2814 373 2815 377
rect 2819 373 2820 377
rect 2814 372 2820 373
rect 2926 377 2932 378
rect 2926 373 2927 377
rect 2931 373 2932 377
rect 2926 372 2932 373
rect 2802 355 2808 356
rect 2802 351 2803 355
rect 2807 351 2808 355
rect 2802 350 2808 351
rect 2816 347 2818 372
rect 2928 347 2930 372
rect 2936 356 2938 462
rect 2998 456 3004 457
rect 2998 452 2999 456
rect 3003 452 3004 456
rect 2998 451 3004 452
rect 3000 427 3002 451
rect 2999 426 3003 427
rect 2999 421 3003 422
rect 3063 426 3067 427
rect 3063 421 3067 422
rect 3064 397 3066 421
rect 3062 396 3068 397
rect 3062 392 3063 396
rect 3067 392 3068 396
rect 3062 391 3068 392
rect 3002 387 3008 388
rect 3002 383 3003 387
rect 3007 383 3008 387
rect 3002 382 3008 383
rect 3004 356 3006 382
rect 3062 377 3068 378
rect 3062 373 3063 377
rect 3067 373 3068 377
rect 3062 372 3068 373
rect 2934 355 2940 356
rect 2934 351 2935 355
rect 2939 351 2940 355
rect 2934 350 2940 351
rect 3002 355 3008 356
rect 3002 351 3003 355
rect 3007 351 3008 355
rect 3002 350 3008 351
rect 3064 347 3066 372
rect 3084 364 3086 462
rect 3174 456 3180 457
rect 3174 452 3175 456
rect 3179 452 3180 456
rect 3174 451 3180 452
rect 3374 456 3380 457
rect 3374 452 3375 456
rect 3379 452 3380 456
rect 3374 451 3380 452
rect 3590 456 3596 457
rect 3590 452 3591 456
rect 3595 452 3596 456
rect 3590 451 3596 452
rect 3806 456 3812 457
rect 3806 452 3807 456
rect 3811 452 3812 456
rect 3806 451 3812 452
rect 3176 427 3178 451
rect 3376 427 3378 451
rect 3592 427 3594 451
rect 3808 427 3810 451
rect 3175 426 3179 427
rect 3175 421 3179 422
rect 3223 426 3227 427
rect 3223 421 3227 422
rect 3375 426 3379 427
rect 3375 421 3379 422
rect 3399 426 3403 427
rect 3399 421 3403 422
rect 3591 426 3595 427
rect 3591 421 3595 422
rect 3783 426 3787 427
rect 3783 421 3787 422
rect 3807 426 3811 427
rect 3807 421 3811 422
rect 3224 397 3226 421
rect 3400 397 3402 421
rect 3592 397 3594 421
rect 3784 397 3786 421
rect 3222 396 3228 397
rect 3222 392 3223 396
rect 3227 392 3228 396
rect 3222 391 3228 392
rect 3398 396 3404 397
rect 3398 392 3399 396
rect 3403 392 3404 396
rect 3398 391 3404 392
rect 3590 396 3596 397
rect 3590 392 3591 396
rect 3595 392 3596 396
rect 3590 391 3596 392
rect 3782 396 3788 397
rect 3782 392 3783 396
rect 3787 392 3788 396
rect 3782 391 3788 392
rect 3860 388 3862 490
rect 3944 477 3946 497
rect 3942 476 3948 477
rect 3942 472 3943 476
rect 3947 472 3948 476
rect 3942 471 3948 472
rect 3882 463 3888 464
rect 3882 459 3883 463
rect 3887 459 3888 463
rect 3882 458 3888 459
rect 3942 459 3948 460
rect 3138 387 3144 388
rect 3138 383 3139 387
rect 3143 383 3144 387
rect 3138 382 3144 383
rect 3298 387 3304 388
rect 3298 383 3299 387
rect 3303 383 3304 387
rect 3298 382 3304 383
rect 3474 387 3480 388
rect 3474 383 3475 387
rect 3479 383 3480 387
rect 3474 382 3480 383
rect 3498 387 3504 388
rect 3498 383 3499 387
rect 3503 383 3504 387
rect 3498 382 3504 383
rect 3858 387 3864 388
rect 3858 383 3859 387
rect 3863 383 3864 387
rect 3858 382 3864 383
rect 3082 363 3088 364
rect 3082 359 3083 363
rect 3087 359 3088 363
rect 3082 358 3088 359
rect 3140 356 3142 382
rect 3222 377 3228 378
rect 3222 373 3223 377
rect 3227 373 3228 377
rect 3222 372 3228 373
rect 3138 355 3144 356
rect 3138 351 3139 355
rect 3143 351 3144 355
rect 3138 350 3144 351
rect 3224 347 3226 372
rect 3300 356 3302 382
rect 3398 377 3404 378
rect 3398 373 3399 377
rect 3403 373 3404 377
rect 3398 372 3404 373
rect 3298 355 3304 356
rect 3298 351 3299 355
rect 3303 351 3304 355
rect 3298 350 3304 351
rect 3400 347 3402 372
rect 3476 356 3478 382
rect 3474 355 3480 356
rect 3474 351 3475 355
rect 3479 351 3480 355
rect 3474 350 3480 351
rect 3500 348 3502 382
rect 3590 377 3596 378
rect 3590 373 3591 377
rect 3595 373 3596 377
rect 3590 372 3596 373
rect 3782 377 3788 378
rect 3782 373 3783 377
rect 3787 373 3788 377
rect 3782 372 3788 373
rect 3498 347 3504 348
rect 3592 347 3594 372
rect 3730 355 3736 356
rect 3730 351 3731 355
rect 3735 351 3736 355
rect 3730 350 3736 351
rect 847 346 851 347
rect 894 346 900 347
rect 903 346 907 347
rect 922 346 928 347
rect 967 346 971 347
rect 847 341 851 342
rect 794 339 800 340
rect 794 335 795 339
rect 799 335 800 339
rect 794 334 800 335
rect 774 319 780 320
rect 774 315 775 319
rect 779 315 780 319
rect 774 314 780 315
rect 896 312 898 346
rect 903 341 907 342
rect 967 341 971 342
rect 1031 346 1035 347
rect 1042 346 1048 347
rect 1087 346 1091 347
rect 1031 341 1035 342
rect 1087 341 1091 342
rect 1151 346 1155 347
rect 1162 346 1168 347
rect 1207 346 1211 347
rect 1151 341 1155 342
rect 1207 341 1211 342
rect 1271 346 1275 347
rect 1282 346 1288 347
rect 1327 346 1331 347
rect 1271 341 1275 342
rect 1327 341 1331 342
rect 1391 346 1395 347
rect 1391 341 1395 342
rect 2007 346 2011 347
rect 2007 341 2011 342
rect 2047 346 2051 347
rect 2047 341 2051 342
rect 2191 346 2195 347
rect 2191 341 2195 342
rect 2327 346 2331 347
rect 2327 341 2331 342
rect 2431 346 2435 347
rect 2431 341 2435 342
rect 2471 346 2475 347
rect 2471 341 2475 342
rect 2527 346 2531 347
rect 2602 343 2603 347
rect 2607 343 2608 347
rect 2602 342 2608 343
rect 2623 346 2627 347
rect 2527 341 2531 342
rect 2623 341 2627 342
rect 2719 346 2723 347
rect 2719 341 2723 342
rect 2783 346 2787 347
rect 2783 341 2787 342
rect 2815 346 2819 347
rect 2815 341 2819 342
rect 2927 346 2931 347
rect 2927 341 2931 342
rect 2951 346 2955 347
rect 2951 341 2955 342
rect 3063 346 3067 347
rect 3063 341 3067 342
rect 3119 346 3123 347
rect 3119 341 3123 342
rect 3223 346 3227 347
rect 3223 341 3227 342
rect 3295 346 3299 347
rect 3295 341 3299 342
rect 3399 346 3403 347
rect 3399 341 3403 342
rect 3471 346 3475 347
rect 3498 343 3499 347
rect 3503 343 3504 347
rect 3498 342 3504 343
rect 3591 346 3595 347
rect 3471 341 3475 342
rect 3591 341 3595 342
rect 3655 346 3659 347
rect 3655 341 3659 342
rect 904 320 906 341
rect 986 339 992 340
rect 986 335 987 339
rect 991 335 992 339
rect 986 334 992 335
rect 902 319 908 320
rect 902 315 903 319
rect 907 315 908 319
rect 902 314 908 315
rect 988 312 990 334
rect 1032 320 1034 341
rect 1114 339 1120 340
rect 1114 335 1115 339
rect 1119 335 1120 339
rect 1114 334 1120 335
rect 1030 319 1036 320
rect 1030 315 1031 319
rect 1035 315 1036 319
rect 1030 314 1036 315
rect 1116 312 1118 334
rect 1152 320 1154 341
rect 1234 339 1240 340
rect 1234 335 1235 339
rect 1239 335 1240 339
rect 1234 334 1240 335
rect 1150 319 1156 320
rect 1150 315 1151 319
rect 1155 315 1156 319
rect 1150 314 1156 315
rect 1236 312 1238 334
rect 1272 320 1274 341
rect 1354 339 1360 340
rect 1354 335 1355 339
rect 1359 335 1360 339
rect 1354 334 1360 335
rect 1270 319 1276 320
rect 1270 315 1271 319
rect 1275 315 1276 319
rect 1270 314 1276 315
rect 1356 312 1358 334
rect 1392 320 1394 341
rect 1602 339 1608 340
rect 1602 335 1603 339
rect 1607 335 1608 339
rect 1602 334 1608 335
rect 1390 319 1396 320
rect 1390 315 1391 319
rect 1395 315 1396 319
rect 1390 314 1396 315
rect 618 311 624 312
rect 618 307 619 311
rect 623 307 624 311
rect 746 311 752 312
rect 618 306 624 307
rect 706 307 712 308
rect 706 303 707 307
rect 711 303 712 307
rect 746 307 747 311
rect 751 307 752 311
rect 746 306 752 307
rect 894 311 900 312
rect 894 307 895 311
rect 899 307 900 311
rect 894 306 900 307
rect 986 311 992 312
rect 986 307 987 311
rect 991 307 992 311
rect 986 306 992 307
rect 1114 311 1120 312
rect 1114 307 1115 311
rect 1119 307 1120 311
rect 1114 306 1120 307
rect 1234 311 1240 312
rect 1234 307 1235 311
rect 1239 307 1240 311
rect 1234 306 1240 307
rect 1354 311 1360 312
rect 1354 307 1355 311
rect 1359 307 1360 311
rect 1354 306 1360 307
rect 706 302 712 303
rect 630 300 636 301
rect 630 296 631 300
rect 635 296 636 300
rect 630 295 636 296
rect 632 267 634 295
rect 559 266 563 267
rect 559 261 563 262
rect 631 266 635 267
rect 631 261 635 262
rect 560 237 562 261
rect 558 236 564 237
rect 558 232 559 236
rect 563 232 564 236
rect 558 231 564 232
rect 298 227 304 228
rect 298 223 299 227
rect 303 223 304 227
rect 298 222 304 223
rect 466 227 472 228
rect 466 223 467 227
rect 471 223 472 227
rect 466 222 472 223
rect 498 227 504 228
rect 498 223 499 227
rect 503 223 504 227
rect 498 222 504 223
rect 222 217 228 218
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 222 213 223 217
rect 227 213 228 217
rect 222 212 228 213
rect 110 211 116 212
rect 112 159 114 211
rect 224 159 226 212
rect 300 196 302 222
rect 390 217 396 218
rect 390 213 391 217
rect 395 213 396 217
rect 390 212 396 213
rect 230 195 236 196
rect 230 191 231 195
rect 235 191 236 195
rect 230 190 236 191
rect 298 195 304 196
rect 298 191 299 195
rect 303 191 304 195
rect 298 190 304 191
rect 111 158 115 159
rect 111 153 115 154
rect 151 158 155 159
rect 151 153 155 154
rect 223 158 227 159
rect 223 153 227 154
rect 112 133 114 153
rect 110 132 116 133
rect 152 132 154 153
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 150 131 156 132
rect 150 127 151 131
rect 155 127 156 131
rect 150 126 156 127
rect 232 124 234 190
rect 392 159 394 212
rect 468 196 470 222
rect 558 217 564 218
rect 558 213 559 217
rect 563 213 564 217
rect 558 212 564 213
rect 466 195 472 196
rect 466 191 467 195
rect 471 191 472 195
rect 466 190 472 191
rect 560 159 562 212
rect 708 196 710 302
rect 774 300 780 301
rect 774 296 775 300
rect 779 296 780 300
rect 774 295 780 296
rect 902 300 908 301
rect 902 296 903 300
rect 907 296 908 300
rect 902 295 908 296
rect 1030 300 1036 301
rect 1030 296 1031 300
rect 1035 296 1036 300
rect 1030 295 1036 296
rect 1150 300 1156 301
rect 1150 296 1151 300
rect 1155 296 1156 300
rect 1150 295 1156 296
rect 1270 300 1276 301
rect 1270 296 1271 300
rect 1275 296 1276 300
rect 1270 295 1276 296
rect 1390 300 1396 301
rect 1390 296 1391 300
rect 1395 296 1396 300
rect 1390 295 1396 296
rect 776 267 778 295
rect 904 267 906 295
rect 1032 267 1034 295
rect 1152 267 1154 295
rect 1272 267 1274 295
rect 1392 267 1394 295
rect 735 266 739 267
rect 735 261 739 262
rect 775 266 779 267
rect 775 261 779 262
rect 903 266 907 267
rect 903 261 907 262
rect 1031 266 1035 267
rect 1031 261 1035 262
rect 1063 266 1067 267
rect 1063 261 1067 262
rect 1151 266 1155 267
rect 1151 261 1155 262
rect 1215 266 1219 267
rect 1215 261 1219 262
rect 1271 266 1275 267
rect 1271 261 1275 262
rect 1359 266 1363 267
rect 1359 261 1363 262
rect 1391 266 1395 267
rect 1391 261 1395 262
rect 1511 266 1515 267
rect 1511 261 1515 262
rect 736 237 738 261
rect 904 237 906 261
rect 1064 237 1066 261
rect 1216 237 1218 261
rect 1360 237 1362 261
rect 1512 237 1514 261
rect 734 236 740 237
rect 734 232 735 236
rect 739 232 740 236
rect 734 231 740 232
rect 902 236 908 237
rect 902 232 903 236
rect 907 232 908 236
rect 902 231 908 232
rect 1062 236 1068 237
rect 1062 232 1063 236
rect 1067 232 1068 236
rect 1062 231 1068 232
rect 1214 236 1220 237
rect 1214 232 1215 236
rect 1219 232 1220 236
rect 1214 231 1220 232
rect 1358 236 1364 237
rect 1358 232 1359 236
rect 1363 232 1364 236
rect 1358 231 1364 232
rect 1510 236 1516 237
rect 1510 232 1511 236
rect 1515 232 1516 236
rect 1510 231 1516 232
rect 1604 228 1606 334
rect 2008 321 2010 341
rect 2048 321 2050 341
rect 2006 320 2012 321
rect 2006 316 2007 320
rect 2011 316 2012 320
rect 2006 315 2012 316
rect 2046 320 2052 321
rect 2192 320 2194 341
rect 2314 339 2320 340
rect 2314 335 2315 339
rect 2319 335 2320 339
rect 2314 334 2320 335
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2190 319 2196 320
rect 2190 315 2191 319
rect 2195 315 2196 319
rect 2190 314 2196 315
rect 2316 312 2318 334
rect 2328 320 2330 341
rect 2434 331 2440 332
rect 2434 327 2435 331
rect 2439 327 2440 331
rect 2434 326 2440 327
rect 2326 319 2332 320
rect 2326 315 2327 319
rect 2331 315 2332 319
rect 2326 314 2332 315
rect 2436 312 2438 326
rect 2472 320 2474 341
rect 2624 320 2626 341
rect 2698 339 2704 340
rect 2698 335 2699 339
rect 2703 335 2704 339
rect 2698 334 2704 335
rect 2470 319 2476 320
rect 2470 315 2471 319
rect 2475 315 2476 319
rect 2470 314 2476 315
rect 2622 319 2628 320
rect 2622 315 2623 319
rect 2627 315 2628 319
rect 2622 314 2628 315
rect 2700 312 2702 334
rect 2706 331 2712 332
rect 2706 327 2707 331
rect 2711 327 2712 331
rect 2706 326 2712 327
rect 2708 312 2710 326
rect 2784 320 2786 341
rect 2952 320 2954 341
rect 3026 339 3032 340
rect 3026 335 3027 339
rect 3031 335 3032 339
rect 3026 334 3032 335
rect 2782 319 2788 320
rect 2782 315 2783 319
rect 2787 315 2788 319
rect 2782 314 2788 315
rect 2950 319 2956 320
rect 2950 315 2951 319
rect 2955 315 2956 319
rect 2950 314 2956 315
rect 3028 312 3030 334
rect 3120 320 3122 341
rect 3194 339 3200 340
rect 3194 335 3195 339
rect 3199 335 3200 339
rect 3194 334 3200 335
rect 3118 319 3124 320
rect 3118 315 3119 319
rect 3123 315 3124 319
rect 3118 314 3124 315
rect 3196 312 3198 334
rect 3296 320 3298 341
rect 3370 339 3376 340
rect 3370 335 3371 339
rect 3375 335 3376 339
rect 3370 334 3376 335
rect 3294 319 3300 320
rect 3294 315 3295 319
rect 3299 315 3300 319
rect 3294 314 3300 315
rect 3372 312 3374 334
rect 3472 320 3474 341
rect 3656 320 3658 341
rect 3470 319 3476 320
rect 3470 315 3471 319
rect 3475 315 3476 319
rect 3470 314 3476 315
rect 3654 319 3660 320
rect 3654 315 3655 319
rect 3659 315 3660 319
rect 3654 314 3660 315
rect 3732 312 3734 350
rect 3784 347 3786 372
rect 3783 346 3787 347
rect 3783 341 3787 342
rect 3839 346 3843 347
rect 3839 341 3843 342
rect 3754 339 3760 340
rect 3754 335 3755 339
rect 3759 335 3760 339
rect 3754 334 3760 335
rect 2314 311 2320 312
rect 2314 307 2315 311
rect 2319 307 2320 311
rect 2434 311 2440 312
rect 2314 306 2320 307
rect 2414 307 2420 308
rect 2006 303 2012 304
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 2414 303 2415 307
rect 2419 303 2420 307
rect 2434 307 2435 311
rect 2439 307 2440 311
rect 2434 306 2440 307
rect 2698 311 2704 312
rect 2698 307 2699 311
rect 2703 307 2704 311
rect 2698 306 2704 307
rect 2706 311 2712 312
rect 2706 307 2707 311
rect 2711 307 2712 311
rect 2706 306 2712 307
rect 3026 311 3032 312
rect 3026 307 3027 311
rect 3031 307 3032 311
rect 3026 306 3032 307
rect 3194 311 3200 312
rect 3194 307 3195 311
rect 3199 307 3200 311
rect 3194 306 3200 307
rect 3370 311 3376 312
rect 3370 307 3371 311
rect 3375 307 3376 311
rect 3370 306 3376 307
rect 3410 311 3416 312
rect 3410 307 3411 311
rect 3415 307 3416 311
rect 3410 306 3416 307
rect 3730 311 3736 312
rect 3730 307 3731 311
rect 3735 307 3736 311
rect 3730 306 3736 307
rect 2414 302 2420 303
rect 2046 298 2052 299
rect 2190 300 2196 301
rect 2008 267 2010 298
rect 2048 271 2050 298
rect 2190 296 2191 300
rect 2195 296 2196 300
rect 2190 295 2196 296
rect 2326 300 2332 301
rect 2326 296 2327 300
rect 2331 296 2332 300
rect 2326 295 2332 296
rect 2192 271 2194 295
rect 2328 271 2330 295
rect 2047 270 2051 271
rect 1663 266 1667 267
rect 1663 261 1667 262
rect 2007 266 2011 267
rect 2047 265 2051 266
rect 2071 270 2075 271
rect 2071 265 2075 266
rect 2191 270 2195 271
rect 2191 265 2195 266
rect 2215 270 2219 271
rect 2215 265 2219 266
rect 2327 270 2331 271
rect 2327 265 2331 266
rect 2399 270 2403 271
rect 2399 265 2403 266
rect 2007 261 2011 262
rect 1664 237 1666 261
rect 1662 236 1668 237
rect 1662 232 1663 236
rect 1667 232 1668 236
rect 2008 234 2010 261
rect 2048 238 2050 265
rect 2072 241 2074 265
rect 2216 241 2218 265
rect 2400 241 2402 265
rect 2070 240 2076 241
rect 2046 237 2052 238
rect 1662 231 1668 232
rect 2006 233 2012 234
rect 2006 229 2007 233
rect 2011 229 2012 233
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2214 240 2220 241
rect 2214 236 2215 240
rect 2219 236 2220 240
rect 2214 235 2220 236
rect 2398 240 2404 241
rect 2398 236 2399 240
rect 2403 236 2404 240
rect 2398 235 2404 236
rect 2046 232 2052 233
rect 2006 228 2012 229
rect 2146 231 2152 232
rect 810 227 816 228
rect 810 223 811 227
rect 815 223 816 227
rect 810 222 816 223
rect 1138 227 1144 228
rect 1138 223 1139 227
rect 1143 223 1144 227
rect 1138 222 1144 223
rect 1290 227 1296 228
rect 1290 223 1291 227
rect 1295 223 1296 227
rect 1290 222 1296 223
rect 1434 227 1440 228
rect 1434 223 1435 227
rect 1439 223 1440 227
rect 1434 222 1440 223
rect 1586 227 1592 228
rect 1586 223 1587 227
rect 1591 223 1592 227
rect 1586 222 1592 223
rect 1602 227 1608 228
rect 1602 223 1603 227
rect 1607 223 1608 227
rect 2146 227 2147 231
rect 2151 227 2152 231
rect 2146 226 2152 227
rect 2290 231 2296 232
rect 2290 227 2291 231
rect 2295 227 2296 231
rect 2290 226 2296 227
rect 1602 222 1608 223
rect 734 217 740 218
rect 734 213 735 217
rect 739 213 740 217
rect 734 212 740 213
rect 706 195 712 196
rect 706 191 707 195
rect 711 191 712 195
rect 706 190 712 191
rect 736 159 738 212
rect 812 196 814 222
rect 902 217 908 218
rect 902 213 903 217
rect 907 213 908 217
rect 902 212 908 213
rect 1062 217 1068 218
rect 1062 213 1063 217
rect 1067 213 1068 217
rect 1062 212 1068 213
rect 810 195 816 196
rect 810 191 811 195
rect 815 191 816 195
rect 810 190 816 191
rect 904 159 906 212
rect 1064 159 1066 212
rect 1140 196 1142 222
rect 1214 217 1220 218
rect 1214 213 1215 217
rect 1219 213 1220 217
rect 1214 212 1220 213
rect 1090 195 1096 196
rect 1090 191 1091 195
rect 1095 191 1096 195
rect 1090 190 1096 191
rect 1138 195 1144 196
rect 1138 191 1139 195
rect 1143 191 1144 195
rect 1138 190 1144 191
rect 247 158 251 159
rect 247 153 251 154
rect 343 158 347 159
rect 343 153 347 154
rect 391 158 395 159
rect 391 153 395 154
rect 439 158 443 159
rect 439 153 443 154
rect 535 158 539 159
rect 535 153 539 154
rect 559 158 563 159
rect 559 153 563 154
rect 631 158 635 159
rect 631 153 635 154
rect 727 158 731 159
rect 727 153 731 154
rect 735 158 739 159
rect 735 153 739 154
rect 823 158 827 159
rect 823 153 827 154
rect 903 158 907 159
rect 903 153 907 154
rect 919 158 923 159
rect 919 153 923 154
rect 1015 158 1019 159
rect 1015 153 1019 154
rect 1063 158 1067 159
rect 1063 153 1067 154
rect 248 132 250 153
rect 344 132 346 153
rect 426 151 432 152
rect 426 147 427 151
rect 431 147 432 151
rect 426 146 432 147
rect 246 131 252 132
rect 246 127 247 131
rect 251 127 252 131
rect 246 126 252 127
rect 342 131 348 132
rect 342 127 343 131
rect 347 127 348 131
rect 342 126 348 127
rect 428 124 430 146
rect 440 132 442 153
rect 522 151 528 152
rect 522 147 523 151
rect 527 147 528 151
rect 522 146 528 147
rect 438 131 444 132
rect 438 127 439 131
rect 443 127 444 131
rect 438 126 444 127
rect 524 124 526 146
rect 536 132 538 153
rect 618 151 624 152
rect 618 147 619 151
rect 623 147 624 151
rect 618 146 624 147
rect 534 131 540 132
rect 534 127 535 131
rect 539 127 540 131
rect 534 126 540 127
rect 620 124 622 146
rect 632 132 634 153
rect 714 151 720 152
rect 714 147 715 151
rect 719 147 720 151
rect 714 146 720 147
rect 630 131 636 132
rect 630 127 631 131
rect 635 127 636 131
rect 630 126 636 127
rect 716 124 718 146
rect 728 132 730 153
rect 810 151 816 152
rect 810 147 811 151
rect 815 147 816 151
rect 810 146 816 147
rect 726 131 732 132
rect 726 127 727 131
rect 731 127 732 131
rect 726 126 732 127
rect 812 124 814 146
rect 824 132 826 153
rect 920 132 922 153
rect 994 151 1000 152
rect 994 147 995 151
rect 999 147 1000 151
rect 994 146 1000 147
rect 822 131 828 132
rect 822 127 823 131
rect 827 127 828 131
rect 822 126 828 127
rect 918 131 924 132
rect 918 127 919 131
rect 923 127 924 131
rect 918 126 924 127
rect 996 124 998 146
rect 1016 132 1018 153
rect 1014 131 1020 132
rect 1014 127 1015 131
rect 1019 127 1020 131
rect 1014 126 1020 127
rect 1092 124 1094 190
rect 1216 159 1218 212
rect 1292 196 1294 222
rect 1358 217 1364 218
rect 1358 213 1359 217
rect 1363 213 1364 217
rect 1358 212 1364 213
rect 1290 195 1296 196
rect 1290 191 1291 195
rect 1295 191 1296 195
rect 1290 190 1296 191
rect 1360 159 1362 212
rect 1436 196 1438 222
rect 1510 217 1516 218
rect 1510 213 1511 217
rect 1515 213 1516 217
rect 1510 212 1516 213
rect 1434 195 1440 196
rect 1434 191 1435 195
rect 1439 191 1440 195
rect 1434 190 1440 191
rect 1512 159 1514 212
rect 1588 196 1590 222
rect 2070 221 2076 222
rect 2046 220 2052 221
rect 1662 217 1668 218
rect 1662 213 1663 217
rect 1667 213 1668 217
rect 1662 212 1668 213
rect 2006 216 2012 217
rect 2006 212 2007 216
rect 2011 212 2012 216
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2070 217 2071 221
rect 2075 217 2076 221
rect 2070 216 2076 217
rect 2046 215 2052 216
rect 1586 195 1592 196
rect 1586 191 1587 195
rect 1591 191 1592 195
rect 1586 190 1592 191
rect 1664 159 1666 212
rect 2006 211 2012 212
rect 2008 159 2010 211
rect 2048 171 2050 215
rect 2072 171 2074 216
rect 2148 200 2150 226
rect 2214 221 2220 222
rect 2214 217 2215 221
rect 2219 217 2220 221
rect 2214 216 2220 217
rect 2146 199 2152 200
rect 2146 195 2147 199
rect 2151 195 2152 199
rect 2146 194 2152 195
rect 2216 171 2218 216
rect 2047 170 2051 171
rect 2047 165 2051 166
rect 2071 170 2075 171
rect 2071 165 2075 166
rect 2191 170 2195 171
rect 2191 165 2195 166
rect 2215 170 2219 171
rect 2215 165 2219 166
rect 1111 158 1115 159
rect 1111 153 1115 154
rect 1207 158 1211 159
rect 1207 153 1211 154
rect 1215 158 1219 159
rect 1215 153 1219 154
rect 1303 158 1307 159
rect 1303 153 1307 154
rect 1359 158 1363 159
rect 1359 153 1363 154
rect 1407 158 1411 159
rect 1407 153 1411 154
rect 1511 158 1515 159
rect 1511 153 1515 154
rect 1615 158 1619 159
rect 1615 153 1619 154
rect 1663 158 1667 159
rect 1663 153 1667 154
rect 1711 158 1715 159
rect 1711 153 1715 154
rect 1807 158 1811 159
rect 1807 153 1811 154
rect 1903 158 1907 159
rect 1903 153 1907 154
rect 2007 158 2011 159
rect 2007 153 2011 154
rect 1098 143 1104 144
rect 1098 139 1099 143
rect 1103 139 1104 143
rect 1098 138 1104 139
rect 1100 124 1102 138
rect 1112 132 1114 153
rect 1194 151 1200 152
rect 1194 147 1195 151
rect 1199 147 1200 151
rect 1194 146 1200 147
rect 1110 131 1116 132
rect 1110 127 1111 131
rect 1115 127 1116 131
rect 1110 126 1116 127
rect 1196 124 1198 146
rect 1208 132 1210 153
rect 1290 151 1296 152
rect 1290 147 1291 151
rect 1295 147 1296 151
rect 1290 146 1296 147
rect 1206 131 1212 132
rect 1206 127 1207 131
rect 1211 127 1212 131
rect 1206 126 1212 127
rect 1292 124 1294 146
rect 1304 132 1306 153
rect 1408 132 1410 153
rect 1512 132 1514 153
rect 1616 132 1618 153
rect 1698 151 1704 152
rect 1698 147 1699 151
rect 1703 147 1704 151
rect 1698 146 1704 147
rect 1302 131 1308 132
rect 1302 127 1303 131
rect 1307 127 1308 131
rect 1302 126 1308 127
rect 1406 131 1412 132
rect 1406 127 1407 131
rect 1411 127 1412 131
rect 1406 126 1412 127
rect 1510 131 1516 132
rect 1510 127 1511 131
rect 1515 127 1516 131
rect 1510 126 1516 127
rect 1614 131 1620 132
rect 1614 127 1615 131
rect 1619 127 1620 131
rect 1614 126 1620 127
rect 1700 124 1702 146
rect 1712 132 1714 153
rect 1794 151 1800 152
rect 1794 147 1795 151
rect 1799 147 1800 151
rect 1794 146 1800 147
rect 1710 131 1716 132
rect 1710 127 1711 131
rect 1715 127 1716 131
rect 1710 126 1716 127
rect 1796 124 1798 146
rect 1808 132 1810 153
rect 1890 151 1896 152
rect 1890 147 1891 151
rect 1895 147 1896 151
rect 1890 146 1896 147
rect 1806 131 1812 132
rect 1806 127 1807 131
rect 1811 127 1812 131
rect 1806 126 1812 127
rect 1892 124 1894 146
rect 1904 132 1906 153
rect 2008 133 2010 153
rect 2048 145 2050 165
rect 2046 144 2052 145
rect 2072 144 2074 165
rect 2192 144 2194 165
rect 2292 164 2294 226
rect 2398 221 2404 222
rect 2398 217 2399 221
rect 2403 217 2404 221
rect 2398 216 2404 217
rect 2400 171 2402 216
rect 2416 200 2418 302
rect 2470 300 2476 301
rect 2470 296 2471 300
rect 2475 296 2476 300
rect 2470 295 2476 296
rect 2622 300 2628 301
rect 2622 296 2623 300
rect 2627 296 2628 300
rect 2622 295 2628 296
rect 2782 300 2788 301
rect 2782 296 2783 300
rect 2787 296 2788 300
rect 2782 295 2788 296
rect 2950 300 2956 301
rect 2950 296 2951 300
rect 2955 296 2956 300
rect 2950 295 2956 296
rect 3118 300 3124 301
rect 3118 296 3119 300
rect 3123 296 3124 300
rect 3118 295 3124 296
rect 3294 300 3300 301
rect 3294 296 3295 300
rect 3299 296 3300 300
rect 3294 295 3300 296
rect 2472 271 2474 295
rect 2624 271 2626 295
rect 2784 271 2786 295
rect 2952 271 2954 295
rect 3120 271 3122 295
rect 3296 271 3298 295
rect 2471 270 2475 271
rect 2471 265 2475 266
rect 2591 270 2595 271
rect 2591 265 2595 266
rect 2623 270 2627 271
rect 2623 265 2627 266
rect 2783 270 2787 271
rect 2783 265 2787 266
rect 2791 270 2795 271
rect 2791 265 2795 266
rect 2951 270 2955 271
rect 2951 265 2955 266
rect 2983 270 2987 271
rect 2983 265 2987 266
rect 3119 270 3123 271
rect 3119 265 3123 266
rect 3167 270 3171 271
rect 3167 265 3171 266
rect 3295 270 3299 271
rect 3295 265 3299 266
rect 3343 270 3347 271
rect 3343 265 3347 266
rect 2592 241 2594 265
rect 2792 241 2794 265
rect 2984 241 2986 265
rect 3168 241 3170 265
rect 3344 241 3346 265
rect 2590 240 2596 241
rect 2590 236 2591 240
rect 2595 236 2596 240
rect 2590 235 2596 236
rect 2790 240 2796 241
rect 2790 236 2791 240
rect 2795 236 2796 240
rect 2790 235 2796 236
rect 2982 240 2988 241
rect 2982 236 2983 240
rect 2987 236 2988 240
rect 2982 235 2988 236
rect 3166 240 3172 241
rect 3166 236 3167 240
rect 3171 236 3172 240
rect 3166 235 3172 236
rect 3342 240 3348 241
rect 3342 236 3343 240
rect 3347 236 3348 240
rect 3342 235 3348 236
rect 2474 231 2480 232
rect 2474 227 2475 231
rect 2479 227 2480 231
rect 2474 226 2480 227
rect 2666 231 2672 232
rect 2666 227 2667 231
rect 2671 227 2672 231
rect 2666 226 2672 227
rect 2674 231 2680 232
rect 2674 227 2675 231
rect 2679 227 2680 231
rect 2674 226 2680 227
rect 2874 231 2880 232
rect 2874 227 2875 231
rect 2879 227 2880 231
rect 2874 226 2880 227
rect 3066 231 3072 232
rect 3066 227 3067 231
rect 3071 227 3072 231
rect 3066 226 3072 227
rect 3250 231 3256 232
rect 3250 227 3251 231
rect 3255 227 3256 231
rect 3250 226 3256 227
rect 2476 200 2478 226
rect 2590 221 2596 222
rect 2590 217 2591 221
rect 2595 217 2596 221
rect 2590 216 2596 217
rect 2414 199 2420 200
rect 2414 195 2415 199
rect 2419 195 2420 199
rect 2414 194 2420 195
rect 2474 199 2480 200
rect 2474 195 2475 199
rect 2479 195 2480 199
rect 2474 194 2480 195
rect 2592 171 2594 216
rect 2668 200 2670 226
rect 2676 208 2678 226
rect 2790 221 2796 222
rect 2790 217 2791 221
rect 2795 217 2796 221
rect 2790 216 2796 217
rect 2674 207 2680 208
rect 2674 203 2675 207
rect 2679 203 2680 207
rect 2674 202 2680 203
rect 2666 199 2672 200
rect 2666 195 2667 199
rect 2671 195 2672 199
rect 2666 194 2672 195
rect 2792 171 2794 216
rect 2343 170 2347 171
rect 2343 165 2347 166
rect 2399 170 2403 171
rect 2399 165 2403 166
rect 2495 170 2499 171
rect 2495 165 2499 166
rect 2591 170 2595 171
rect 2591 165 2595 166
rect 2647 170 2651 171
rect 2647 165 2651 166
rect 2791 170 2795 171
rect 2791 165 2795 166
rect 2799 170 2803 171
rect 2799 165 2803 166
rect 2290 163 2296 164
rect 2290 159 2291 163
rect 2295 159 2296 163
rect 2290 158 2296 159
rect 2344 144 2346 165
rect 2418 163 2424 164
rect 2418 159 2419 163
rect 2423 159 2424 163
rect 2418 158 2424 159
rect 2046 140 2047 144
rect 2051 140 2052 144
rect 2046 139 2052 140
rect 2070 143 2076 144
rect 2070 139 2071 143
rect 2075 139 2076 143
rect 2070 138 2076 139
rect 2190 143 2196 144
rect 2190 139 2191 143
rect 2195 139 2196 143
rect 2190 138 2196 139
rect 2342 143 2348 144
rect 2342 139 2343 143
rect 2347 139 2348 143
rect 2342 138 2348 139
rect 2420 136 2422 158
rect 2496 144 2498 165
rect 2570 163 2576 164
rect 2570 159 2571 163
rect 2575 159 2576 163
rect 2570 158 2576 159
rect 2494 143 2500 144
rect 2494 139 2495 143
rect 2499 139 2500 143
rect 2494 138 2500 139
rect 2572 136 2574 158
rect 2578 155 2584 156
rect 2578 151 2579 155
rect 2583 151 2584 155
rect 2578 150 2584 151
rect 2580 136 2582 150
rect 2648 144 2650 165
rect 2800 144 2802 165
rect 2876 164 2878 226
rect 2982 221 2988 222
rect 2982 217 2983 221
rect 2987 217 2988 221
rect 2982 216 2988 217
rect 2984 171 2986 216
rect 3068 200 3070 226
rect 3166 221 3172 222
rect 3166 217 3167 221
rect 3171 217 3172 221
rect 3166 216 3172 217
rect 3066 199 3072 200
rect 3066 195 3067 199
rect 3071 195 3072 199
rect 3066 194 3072 195
rect 3168 171 3170 216
rect 3252 200 3254 226
rect 3342 221 3348 222
rect 3342 217 3343 221
rect 3347 217 3348 221
rect 3342 216 3348 217
rect 3250 199 3256 200
rect 3250 195 3251 199
rect 3255 195 3256 199
rect 3250 194 3256 195
rect 3344 171 3346 216
rect 3412 200 3414 306
rect 3470 300 3476 301
rect 3470 296 3471 300
rect 3475 296 3476 300
rect 3470 295 3476 296
rect 3654 300 3660 301
rect 3654 296 3655 300
rect 3659 296 3660 300
rect 3654 295 3660 296
rect 3472 271 3474 295
rect 3656 271 3658 295
rect 3471 270 3475 271
rect 3471 265 3475 266
rect 3511 270 3515 271
rect 3511 265 3515 266
rect 3655 270 3659 271
rect 3655 265 3659 266
rect 3687 270 3691 271
rect 3687 265 3691 266
rect 3512 241 3514 265
rect 3688 241 3690 265
rect 3510 240 3516 241
rect 3510 236 3511 240
rect 3515 236 3516 240
rect 3510 235 3516 236
rect 3686 240 3692 241
rect 3686 236 3687 240
rect 3691 236 3692 240
rect 3686 235 3692 236
rect 3756 232 3758 334
rect 3840 320 3842 341
rect 3884 340 3886 458
rect 3942 455 3943 459
rect 3947 455 3948 459
rect 3942 454 3948 455
rect 3944 427 3946 454
rect 3943 426 3947 427
rect 3943 421 3947 422
rect 3944 394 3946 421
rect 3942 393 3948 394
rect 3942 389 3943 393
rect 3947 389 3948 393
rect 3942 388 3948 389
rect 3942 376 3948 377
rect 3942 372 3943 376
rect 3947 372 3948 376
rect 3942 371 3948 372
rect 3944 347 3946 371
rect 3943 346 3947 347
rect 3943 341 3947 342
rect 3882 339 3888 340
rect 3882 335 3883 339
rect 3887 335 3888 339
rect 3882 334 3888 335
rect 3944 321 3946 341
rect 3942 320 3948 321
rect 3838 319 3844 320
rect 3838 315 3839 319
rect 3843 315 3844 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3838 314 3844 315
rect 3914 307 3920 308
rect 3914 303 3915 307
rect 3919 303 3920 307
rect 3914 302 3920 303
rect 3942 303 3948 304
rect 3838 300 3844 301
rect 3838 296 3839 300
rect 3843 296 3844 300
rect 3838 295 3844 296
rect 3840 271 3842 295
rect 3839 270 3843 271
rect 3839 265 3843 266
rect 3840 241 3842 265
rect 3838 240 3844 241
rect 3838 236 3839 240
rect 3843 236 3844 240
rect 3838 235 3844 236
rect 3586 231 3592 232
rect 3586 227 3587 231
rect 3591 227 3592 231
rect 3586 226 3592 227
rect 3754 231 3760 232
rect 3754 227 3755 231
rect 3759 227 3760 231
rect 3754 226 3760 227
rect 3906 231 3912 232
rect 3906 227 3907 231
rect 3911 227 3912 231
rect 3906 226 3912 227
rect 3510 221 3516 222
rect 3510 217 3511 221
rect 3515 217 3516 221
rect 3510 216 3516 217
rect 3410 199 3416 200
rect 3410 195 3411 199
rect 3415 195 3416 199
rect 3410 194 3416 195
rect 3512 171 3514 216
rect 3588 200 3590 226
rect 3686 221 3692 222
rect 3686 217 3687 221
rect 3691 217 3692 221
rect 3686 216 3692 217
rect 3838 221 3844 222
rect 3838 217 3839 221
rect 3843 217 3844 221
rect 3838 216 3844 217
rect 3586 199 3592 200
rect 3586 195 3587 199
rect 3591 195 3592 199
rect 3586 194 3592 195
rect 3630 191 3636 192
rect 3630 187 3631 191
rect 3635 187 3636 191
rect 3630 186 3636 187
rect 2943 170 2947 171
rect 2943 165 2947 166
rect 2983 170 2987 171
rect 2983 165 2987 166
rect 3071 170 3075 171
rect 3071 165 3075 166
rect 3167 170 3171 171
rect 3167 165 3171 166
rect 3191 170 3195 171
rect 3191 165 3195 166
rect 3311 170 3315 171
rect 3311 165 3315 166
rect 3343 170 3347 171
rect 3343 165 3347 166
rect 3423 170 3427 171
rect 3423 165 3427 166
rect 3511 170 3515 171
rect 3511 165 3515 166
rect 3527 170 3531 171
rect 3527 165 3531 166
rect 2874 163 2880 164
rect 2874 159 2875 163
rect 2879 159 2880 163
rect 2874 158 2880 159
rect 2918 163 2924 164
rect 2918 159 2919 163
rect 2923 159 2924 163
rect 2918 158 2924 159
rect 2646 143 2652 144
rect 2646 139 2647 143
rect 2651 139 2652 143
rect 2646 138 2652 139
rect 2798 143 2804 144
rect 2798 139 2799 143
rect 2803 139 2804 143
rect 2798 138 2804 139
rect 2920 136 2922 158
rect 2944 144 2946 165
rect 3018 163 3024 164
rect 3018 159 3019 163
rect 3023 159 3024 163
rect 3018 158 3024 159
rect 2942 143 2948 144
rect 2942 139 2943 143
rect 2947 139 2948 143
rect 2942 138 2948 139
rect 3020 136 3022 158
rect 3072 144 3074 165
rect 3146 163 3152 164
rect 3146 159 3147 163
rect 3151 159 3152 163
rect 3146 158 3152 159
rect 3070 143 3076 144
rect 3070 139 3071 143
rect 3075 139 3076 143
rect 3070 138 3076 139
rect 3148 136 3150 158
rect 3192 144 3194 165
rect 3266 163 3272 164
rect 3266 159 3267 163
rect 3271 159 3272 163
rect 3266 158 3272 159
rect 3190 143 3196 144
rect 3190 139 3191 143
rect 3195 139 3196 143
rect 3190 138 3196 139
rect 3268 136 3270 158
rect 3312 144 3314 165
rect 3386 163 3392 164
rect 3386 159 3387 163
rect 3391 159 3392 163
rect 3386 158 3392 159
rect 3310 143 3316 144
rect 3310 139 3311 143
rect 3315 139 3316 143
rect 3310 138 3316 139
rect 3388 136 3390 158
rect 3424 144 3426 165
rect 3498 163 3504 164
rect 3498 159 3499 163
rect 3503 159 3504 163
rect 3498 158 3504 159
rect 3422 143 3428 144
rect 3422 139 3423 143
rect 3427 139 3428 143
rect 3422 138 3428 139
rect 3500 136 3502 158
rect 3528 144 3530 165
rect 3602 163 3608 164
rect 3602 159 3603 163
rect 3607 159 3608 163
rect 3602 158 3608 159
rect 3526 143 3532 144
rect 3526 139 3527 143
rect 3531 139 3532 143
rect 3526 138 3532 139
rect 3604 136 3606 158
rect 3632 136 3634 186
rect 3688 171 3690 216
rect 3840 171 3842 216
rect 3639 170 3643 171
rect 3639 165 3643 166
rect 3687 170 3691 171
rect 3687 165 3691 166
rect 3743 170 3747 171
rect 3743 165 3747 166
rect 3839 170 3843 171
rect 3839 165 3843 166
rect 3640 144 3642 165
rect 3744 144 3746 165
rect 3826 163 3832 164
rect 3826 159 3827 163
rect 3831 159 3832 163
rect 3826 158 3832 159
rect 3638 143 3644 144
rect 3638 139 3639 143
rect 3643 139 3644 143
rect 3638 138 3644 139
rect 3742 143 3748 144
rect 3742 139 3743 143
rect 3747 139 3748 143
rect 3742 138 3748 139
rect 3828 136 3830 158
rect 3840 144 3842 165
rect 3908 164 3910 226
rect 3916 200 3918 302
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3944 271 3946 298
rect 3943 270 3947 271
rect 3943 265 3947 266
rect 3944 238 3946 265
rect 3942 237 3948 238
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 3942 215 3948 216
rect 3914 199 3920 200
rect 3914 195 3915 199
rect 3919 195 3920 199
rect 3914 194 3920 195
rect 3944 171 3946 215
rect 3943 170 3947 171
rect 3943 165 3947 166
rect 3906 163 3912 164
rect 3906 159 3907 163
rect 3911 159 3912 163
rect 3906 158 3912 159
rect 3944 145 3946 165
rect 3942 144 3948 145
rect 3838 143 3844 144
rect 3838 139 3839 143
rect 3843 139 3844 143
rect 3942 140 3943 144
rect 3947 140 3948 144
rect 3942 139 3948 140
rect 3838 138 3844 139
rect 2418 135 2424 136
rect 2006 132 2012 133
rect 1902 131 1908 132
rect 1902 127 1903 131
rect 1907 127 1908 131
rect 2006 128 2007 132
rect 2011 128 2012 132
rect 2418 131 2419 135
rect 2423 131 2424 135
rect 2418 130 2424 131
rect 2570 135 2576 136
rect 2570 131 2571 135
rect 2575 131 2576 135
rect 2570 130 2576 131
rect 2578 135 2584 136
rect 2578 131 2579 135
rect 2583 131 2584 135
rect 2578 130 2584 131
rect 2918 135 2924 136
rect 2918 131 2919 135
rect 2923 131 2924 135
rect 2918 130 2924 131
rect 3018 135 3024 136
rect 3018 131 3019 135
rect 3023 131 3024 135
rect 3018 130 3024 131
rect 3146 135 3152 136
rect 3146 131 3147 135
rect 3151 131 3152 135
rect 3146 130 3152 131
rect 3266 135 3272 136
rect 3266 131 3267 135
rect 3271 131 3272 135
rect 3266 130 3272 131
rect 3386 135 3392 136
rect 3386 131 3387 135
rect 3391 131 3392 135
rect 3386 130 3392 131
rect 3498 135 3504 136
rect 3498 131 3499 135
rect 3503 131 3504 135
rect 3498 130 3504 131
rect 3602 135 3608 136
rect 3602 131 3603 135
rect 3607 131 3608 135
rect 3602 130 3608 131
rect 3630 135 3636 136
rect 3630 131 3631 135
rect 3635 131 3636 135
rect 3630 130 3636 131
rect 3826 135 3832 136
rect 3826 131 3827 135
rect 3831 131 3832 135
rect 3826 130 3832 131
rect 2006 127 2012 128
rect 2046 127 2052 128
rect 1902 126 1908 127
rect 226 123 234 124
rect 226 119 227 123
rect 231 120 234 123
rect 426 123 432 124
rect 231 119 232 120
rect 226 118 232 119
rect 426 119 427 123
rect 431 119 432 123
rect 426 118 432 119
rect 522 123 528 124
rect 522 119 523 123
rect 527 119 528 123
rect 522 118 528 119
rect 618 123 624 124
rect 618 119 619 123
rect 623 119 624 123
rect 618 118 624 119
rect 714 123 720 124
rect 714 119 715 123
rect 719 119 720 123
rect 714 118 720 119
rect 810 123 816 124
rect 810 119 811 123
rect 815 119 816 123
rect 810 118 816 119
rect 994 123 1000 124
rect 994 119 995 123
rect 999 119 1000 123
rect 994 118 1000 119
rect 1090 123 1096 124
rect 1090 119 1091 123
rect 1095 119 1096 123
rect 1090 118 1096 119
rect 1098 123 1104 124
rect 1098 119 1099 123
rect 1103 119 1104 123
rect 1098 118 1104 119
rect 1194 123 1200 124
rect 1194 119 1195 123
rect 1199 119 1200 123
rect 1194 118 1200 119
rect 1290 123 1296 124
rect 1290 119 1291 123
rect 1295 119 1296 123
rect 1290 118 1296 119
rect 1698 123 1704 124
rect 1698 119 1699 123
rect 1703 119 1704 123
rect 1698 118 1704 119
rect 1794 123 1800 124
rect 1794 119 1795 123
rect 1799 119 1800 123
rect 1794 118 1800 119
rect 1890 123 1896 124
rect 1890 119 1891 123
rect 1895 119 1896 123
rect 2046 123 2047 127
rect 2051 123 2052 127
rect 3942 127 3948 128
rect 2046 122 2052 123
rect 2070 124 2076 125
rect 1890 118 1896 119
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 2006 115 2012 116
rect 110 110 116 111
rect 150 112 156 113
rect 112 83 114 110
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 246 112 252 113
rect 246 108 247 112
rect 251 108 252 112
rect 246 107 252 108
rect 342 112 348 113
rect 342 108 343 112
rect 347 108 348 112
rect 342 107 348 108
rect 438 112 444 113
rect 438 108 439 112
rect 443 108 444 112
rect 438 107 444 108
rect 534 112 540 113
rect 534 108 535 112
rect 539 108 540 112
rect 534 107 540 108
rect 630 112 636 113
rect 630 108 631 112
rect 635 108 636 112
rect 630 107 636 108
rect 726 112 732 113
rect 726 108 727 112
rect 731 108 732 112
rect 726 107 732 108
rect 822 112 828 113
rect 822 108 823 112
rect 827 108 828 112
rect 822 107 828 108
rect 918 112 924 113
rect 918 108 919 112
rect 923 108 924 112
rect 918 107 924 108
rect 1014 112 1020 113
rect 1014 108 1015 112
rect 1019 108 1020 112
rect 1014 107 1020 108
rect 1110 112 1116 113
rect 1110 108 1111 112
rect 1115 108 1116 112
rect 1110 107 1116 108
rect 1206 112 1212 113
rect 1206 108 1207 112
rect 1211 108 1212 112
rect 1206 107 1212 108
rect 1302 112 1308 113
rect 1302 108 1303 112
rect 1307 108 1308 112
rect 1302 107 1308 108
rect 1406 112 1412 113
rect 1406 108 1407 112
rect 1411 108 1412 112
rect 1406 107 1412 108
rect 1510 112 1516 113
rect 1510 108 1511 112
rect 1515 108 1516 112
rect 1510 107 1516 108
rect 1614 112 1620 113
rect 1614 108 1615 112
rect 1619 108 1620 112
rect 1614 107 1620 108
rect 1710 112 1716 113
rect 1710 108 1711 112
rect 1715 108 1716 112
rect 1710 107 1716 108
rect 1806 112 1812 113
rect 1806 108 1807 112
rect 1811 108 1812 112
rect 1806 107 1812 108
rect 1902 112 1908 113
rect 1902 108 1903 112
rect 1907 108 1908 112
rect 2006 111 2007 115
rect 2011 111 2012 115
rect 2006 110 2012 111
rect 1902 107 1908 108
rect 152 83 154 107
rect 248 83 250 107
rect 344 83 346 107
rect 440 83 442 107
rect 536 83 538 107
rect 632 83 634 107
rect 728 83 730 107
rect 824 83 826 107
rect 920 83 922 107
rect 1016 83 1018 107
rect 1112 83 1114 107
rect 1208 83 1210 107
rect 1304 83 1306 107
rect 1408 83 1410 107
rect 1512 83 1514 107
rect 1616 83 1618 107
rect 1712 83 1714 107
rect 1808 83 1810 107
rect 1904 83 1906 107
rect 2008 83 2010 110
rect 2048 95 2050 122
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 2190 124 2196 125
rect 2190 120 2191 124
rect 2195 120 2196 124
rect 2190 119 2196 120
rect 2342 124 2348 125
rect 2342 120 2343 124
rect 2347 120 2348 124
rect 2342 119 2348 120
rect 2494 124 2500 125
rect 2494 120 2495 124
rect 2499 120 2500 124
rect 2494 119 2500 120
rect 2646 124 2652 125
rect 2646 120 2647 124
rect 2651 120 2652 124
rect 2646 119 2652 120
rect 2798 124 2804 125
rect 2798 120 2799 124
rect 2803 120 2804 124
rect 2798 119 2804 120
rect 2942 124 2948 125
rect 2942 120 2943 124
rect 2947 120 2948 124
rect 2942 119 2948 120
rect 3070 124 3076 125
rect 3070 120 3071 124
rect 3075 120 3076 124
rect 3070 119 3076 120
rect 3190 124 3196 125
rect 3190 120 3191 124
rect 3195 120 3196 124
rect 3190 119 3196 120
rect 3310 124 3316 125
rect 3310 120 3311 124
rect 3315 120 3316 124
rect 3310 119 3316 120
rect 3422 124 3428 125
rect 3422 120 3423 124
rect 3427 120 3428 124
rect 3422 119 3428 120
rect 3526 124 3532 125
rect 3526 120 3527 124
rect 3531 120 3532 124
rect 3526 119 3532 120
rect 3638 124 3644 125
rect 3638 120 3639 124
rect 3643 120 3644 124
rect 3638 119 3644 120
rect 3742 124 3748 125
rect 3742 120 3743 124
rect 3747 120 3748 124
rect 3742 119 3748 120
rect 3838 124 3844 125
rect 3838 120 3839 124
rect 3843 120 3844 124
rect 3942 123 3943 127
rect 3947 123 3948 127
rect 3942 122 3948 123
rect 3838 119 3844 120
rect 2072 95 2074 119
rect 2192 95 2194 119
rect 2344 95 2346 119
rect 2496 95 2498 119
rect 2648 95 2650 119
rect 2800 95 2802 119
rect 2944 95 2946 119
rect 3072 95 3074 119
rect 3192 95 3194 119
rect 3312 95 3314 119
rect 3424 95 3426 119
rect 3528 95 3530 119
rect 3640 95 3642 119
rect 3744 95 3746 119
rect 3840 95 3842 119
rect 3944 95 3946 122
rect 2047 94 2051 95
rect 2047 89 2051 90
rect 2071 94 2075 95
rect 2071 89 2075 90
rect 2191 94 2195 95
rect 2191 89 2195 90
rect 2343 94 2347 95
rect 2343 89 2347 90
rect 2495 94 2499 95
rect 2495 89 2499 90
rect 2647 94 2651 95
rect 2647 89 2651 90
rect 2799 94 2803 95
rect 2799 89 2803 90
rect 2943 94 2947 95
rect 2943 89 2947 90
rect 3071 94 3075 95
rect 3071 89 3075 90
rect 3191 94 3195 95
rect 3191 89 3195 90
rect 3311 94 3315 95
rect 3311 89 3315 90
rect 3423 94 3427 95
rect 3423 89 3427 90
rect 3527 94 3531 95
rect 3527 89 3531 90
rect 3639 94 3643 95
rect 3639 89 3643 90
rect 3743 94 3747 95
rect 3743 89 3747 90
rect 3839 94 3843 95
rect 3839 89 3843 90
rect 3943 94 3947 95
rect 3943 89 3947 90
rect 111 82 115 83
rect 111 77 115 78
rect 151 82 155 83
rect 151 77 155 78
rect 247 82 251 83
rect 247 77 251 78
rect 343 82 347 83
rect 343 77 347 78
rect 439 82 443 83
rect 439 77 443 78
rect 535 82 539 83
rect 535 77 539 78
rect 631 82 635 83
rect 631 77 635 78
rect 727 82 731 83
rect 727 77 731 78
rect 823 82 827 83
rect 823 77 827 78
rect 919 82 923 83
rect 919 77 923 78
rect 1015 82 1019 83
rect 1015 77 1019 78
rect 1111 82 1115 83
rect 1111 77 1115 78
rect 1207 82 1211 83
rect 1207 77 1211 78
rect 1303 82 1307 83
rect 1303 77 1307 78
rect 1407 82 1411 83
rect 1407 77 1411 78
rect 1511 82 1515 83
rect 1511 77 1515 78
rect 1615 82 1619 83
rect 1615 77 1619 78
rect 1711 82 1715 83
rect 1711 77 1715 78
rect 1807 82 1811 83
rect 1807 77 1811 78
rect 1903 82 1907 83
rect 1903 77 1907 78
rect 2007 82 2011 83
rect 2007 77 2011 78
<< m4c >>
rect 2047 4018 2051 4022
rect 2071 4018 2075 4022
rect 2327 4018 2331 4022
rect 2591 4018 2595 4022
rect 2839 4018 2843 4022
rect 3087 4018 3091 4022
rect 3343 4018 3347 4022
rect 3943 4018 3947 4022
rect 111 3998 115 4002
rect 311 3998 315 4002
rect 511 3998 515 4002
rect 703 3998 707 4002
rect 887 3998 891 4002
rect 1063 3998 1067 4002
rect 1231 3998 1235 4002
rect 1383 3998 1387 4002
rect 1519 3998 1523 4002
rect 1655 3998 1659 4002
rect 1791 3998 1795 4002
rect 1903 3998 1907 4002
rect 2007 3998 2011 4002
rect 111 3922 115 3926
rect 279 3922 283 3926
rect 311 3922 315 3926
rect 111 3838 115 3842
rect 231 3838 235 3842
rect 279 3838 283 3842
rect 415 3922 419 3926
rect 511 3922 515 3926
rect 567 3922 571 3926
rect 703 3922 707 3926
rect 735 3922 739 3926
rect 887 3922 891 3926
rect 911 3922 915 3926
rect 1063 3922 1067 3926
rect 2047 3942 2051 3946
rect 2071 3942 2075 3946
rect 2127 3942 2131 3946
rect 1095 3922 1099 3926
rect 1231 3922 1235 3926
rect 1287 3922 1291 3926
rect 1383 3922 1387 3926
rect 1479 3922 1483 3926
rect 1519 3922 1523 3926
rect 1655 3922 1659 3926
rect 1679 3922 1683 3926
rect 1791 3922 1795 3926
rect 1903 3922 1907 3926
rect 2007 3922 2011 3926
rect 335 3838 339 3842
rect 415 3838 419 3842
rect 439 3838 443 3842
rect 535 3838 539 3842
rect 567 3838 571 3842
rect 631 3838 635 3842
rect 727 3838 731 3842
rect 735 3838 739 3842
rect 831 3838 835 3842
rect 911 3838 915 3842
rect 935 3838 939 3842
rect 1039 3838 1043 3842
rect 111 3762 115 3766
rect 159 3762 163 3766
rect 231 3762 235 3766
rect 335 3762 339 3766
rect 351 3762 355 3766
rect 439 3762 443 3766
rect 535 3762 539 3766
rect 551 3762 555 3766
rect 631 3762 635 3766
rect 727 3762 731 3766
rect 751 3762 755 3766
rect 111 3678 115 3682
rect 151 3678 155 3682
rect 159 3678 163 3682
rect 1095 3838 1099 3842
rect 1151 3838 1155 3842
rect 1263 3838 1267 3842
rect 1287 3838 1291 3842
rect 1383 3838 1387 3842
rect 1479 3838 1483 3842
rect 1503 3838 1507 3842
rect 1631 3838 1635 3842
rect 1679 3838 1683 3842
rect 2271 3942 2275 3946
rect 2327 3942 2331 3946
rect 2439 3942 2443 3946
rect 2591 3942 2595 3946
rect 2615 3942 2619 3946
rect 2799 3942 2803 3946
rect 2839 3942 2843 3946
rect 2983 3942 2987 3946
rect 3087 3942 3091 3946
rect 3175 3942 3179 3946
rect 2047 3866 2051 3870
rect 2127 3866 2131 3870
rect 2263 3866 2267 3870
rect 2271 3866 2275 3870
rect 2375 3866 2379 3870
rect 2439 3866 2443 3870
rect 2495 3866 2499 3870
rect 2615 3866 2619 3870
rect 2631 3866 2635 3870
rect 2775 3866 2779 3870
rect 2799 3866 2803 3870
rect 2007 3838 2011 3842
rect 2047 3774 2051 3778
rect 2071 3774 2075 3778
rect 2183 3774 2187 3778
rect 2263 3774 2267 3778
rect 2327 3774 2331 3778
rect 2375 3774 2379 3778
rect 831 3762 835 3766
rect 935 3762 939 3766
rect 959 3762 963 3766
rect 1039 3762 1043 3766
rect 1151 3762 1155 3766
rect 1167 3762 1171 3766
rect 1263 3762 1267 3766
rect 1383 3762 1387 3766
rect 1503 3762 1507 3766
rect 1607 3762 1611 3766
rect 1631 3762 1635 3766
rect 2007 3762 2011 3766
rect 351 3678 355 3682
rect 383 3678 387 3682
rect 551 3678 555 3682
rect 615 3678 619 3682
rect 751 3678 755 3682
rect 839 3678 843 3682
rect 959 3678 963 3682
rect 1055 3678 1059 3682
rect 1167 3678 1171 3682
rect 1263 3678 1267 3682
rect 111 3598 115 3602
rect 151 3598 155 3602
rect 167 3598 171 3602
rect 359 3598 363 3602
rect 383 3598 387 3602
rect 559 3598 563 3602
rect 615 3598 619 3602
rect 775 3598 779 3602
rect 839 3598 843 3602
rect 991 3598 995 3602
rect 1055 3598 1059 3602
rect 1215 3598 1219 3602
rect 1263 3598 1267 3602
rect 1383 3678 1387 3682
rect 1479 3678 1483 3682
rect 2919 3866 2923 3870
rect 2983 3866 2987 3870
rect 3343 3942 3347 3946
rect 3367 3942 3371 3946
rect 3559 3942 3563 3946
rect 3943 3942 3947 3946
rect 3063 3866 3067 3870
rect 3175 3866 3179 3870
rect 3207 3866 3211 3870
rect 3343 3866 3347 3870
rect 3367 3866 3371 3870
rect 3471 3866 3475 3870
rect 2479 3774 2483 3778
rect 2495 3774 2499 3778
rect 2631 3774 2635 3778
rect 2639 3774 2643 3778
rect 2775 3774 2779 3778
rect 2807 3774 2811 3778
rect 2919 3774 2923 3778
rect 2983 3774 2987 3778
rect 3063 3774 3067 3778
rect 3159 3774 3163 3778
rect 3207 3774 3211 3778
rect 2047 3686 2051 3690
rect 2071 3686 2075 3690
rect 1607 3678 1611 3682
rect 1695 3678 1699 3682
rect 2007 3678 2011 3682
rect 1447 3598 1451 3602
rect 1479 3598 1483 3602
rect 1687 3598 1691 3602
rect 1695 3598 1699 3602
rect 111 3514 115 3518
rect 167 3514 171 3518
rect 295 3514 299 3518
rect 359 3514 363 3518
rect 431 3514 435 3518
rect 559 3514 563 3518
rect 583 3514 587 3518
rect 743 3514 747 3518
rect 775 3514 779 3518
rect 911 3514 915 3518
rect 991 3514 995 3518
rect 1079 3514 1083 3518
rect 1215 3514 1219 3518
rect 1247 3514 1251 3518
rect 1423 3514 1427 3518
rect 1447 3514 1451 3518
rect 1599 3514 1603 3518
rect 1687 3514 1691 3518
rect 2183 3686 2187 3690
rect 2199 3686 2203 3690
rect 2327 3686 2331 3690
rect 2367 3686 2371 3690
rect 2479 3686 2483 3690
rect 2551 3686 2555 3690
rect 2639 3686 2643 3690
rect 2735 3686 2739 3690
rect 2807 3686 2811 3690
rect 2927 3686 2931 3690
rect 2983 3686 2987 3690
rect 3559 3866 3563 3870
rect 3599 3866 3603 3870
rect 3727 3866 3731 3870
rect 3839 3866 3843 3870
rect 3943 3866 3947 3870
rect 3335 3774 3339 3778
rect 3343 3774 3347 3778
rect 3471 3774 3475 3778
rect 3511 3774 3515 3778
rect 3599 3774 3603 3778
rect 3687 3774 3691 3778
rect 3727 3774 3731 3778
rect 3839 3774 3843 3778
rect 3111 3686 3115 3690
rect 3159 3686 3163 3690
rect 3295 3686 3299 3690
rect 3335 3686 3339 3690
rect 3479 3686 3483 3690
rect 3511 3686 3515 3690
rect 2047 3606 2051 3610
rect 2071 3606 2075 3610
rect 2103 3606 2107 3610
rect 2007 3598 2011 3602
rect 2199 3606 2203 3610
rect 2279 3606 2283 3610
rect 2367 3606 2371 3610
rect 2471 3606 2475 3610
rect 2551 3606 2555 3610
rect 2671 3606 2675 3610
rect 2735 3606 2739 3610
rect 2871 3606 2875 3610
rect 2927 3606 2931 3610
rect 3063 3606 3067 3610
rect 3111 3606 3115 3610
rect 2047 3526 2051 3530
rect 2103 3526 2107 3530
rect 2279 3526 2283 3530
rect 2327 3526 2331 3530
rect 2447 3526 2451 3530
rect 2471 3526 2475 3530
rect 2583 3526 2587 3530
rect 1775 3514 1779 3518
rect 2007 3514 2011 3518
rect 111 3418 115 3422
rect 295 3418 299 3422
rect 431 3418 435 3422
rect 495 3418 499 3422
rect 583 3418 587 3422
rect 647 3418 651 3422
rect 743 3418 747 3422
rect 799 3418 803 3422
rect 911 3418 915 3422
rect 959 3418 963 3422
rect 111 3330 115 3334
rect 135 3330 139 3334
rect 295 3330 299 3334
rect 479 3330 483 3334
rect 495 3330 499 3334
rect 1079 3418 1083 3422
rect 1127 3418 1131 3422
rect 1247 3418 1251 3422
rect 1295 3418 1299 3422
rect 1423 3418 1427 3422
rect 1463 3418 1467 3422
rect 1599 3418 1603 3422
rect 1639 3418 1643 3422
rect 2047 3450 2051 3454
rect 2327 3450 2331 3454
rect 2447 3450 2451 3454
rect 2671 3526 2675 3530
rect 2735 3526 2739 3530
rect 2871 3526 2875 3530
rect 2911 3526 2915 3530
rect 3671 3686 3675 3690
rect 3687 3686 3691 3690
rect 3943 3774 3947 3778
rect 3839 3686 3843 3690
rect 3255 3606 3259 3610
rect 3295 3606 3299 3610
rect 3447 3606 3451 3610
rect 3479 3606 3483 3610
rect 3639 3606 3643 3610
rect 3671 3606 3675 3610
rect 3943 3686 3947 3690
rect 3839 3606 3843 3610
rect 3943 3606 3947 3610
rect 3063 3526 3067 3530
rect 3111 3526 3115 3530
rect 3255 3526 3259 3530
rect 3335 3526 3339 3530
rect 3447 3526 3451 3530
rect 3567 3526 3571 3530
rect 3639 3526 3643 3530
rect 3807 3526 3811 3530
rect 3839 3526 3843 3530
rect 2551 3450 2555 3454
rect 2583 3450 2587 3454
rect 2663 3450 2667 3454
rect 2735 3450 2739 3454
rect 2775 3450 2779 3454
rect 2903 3450 2907 3454
rect 2911 3450 2915 3454
rect 3047 3450 3051 3454
rect 3111 3450 3115 3454
rect 3207 3450 3211 3454
rect 3335 3450 3339 3454
rect 3383 3450 3387 3454
rect 3567 3450 3571 3454
rect 1775 3418 1779 3422
rect 1815 3418 1819 3422
rect 2007 3418 2011 3422
rect 647 3330 651 3334
rect 671 3330 675 3334
rect 799 3330 803 3334
rect 863 3330 867 3334
rect 959 3330 963 3334
rect 1055 3330 1059 3334
rect 1127 3330 1131 3334
rect 111 3250 115 3254
rect 135 3250 139 3254
rect 295 3250 299 3254
rect 319 3250 323 3254
rect 479 3250 483 3254
rect 519 3250 523 3254
rect 671 3250 675 3254
rect 719 3250 723 3254
rect 863 3250 867 3254
rect 911 3250 915 3254
rect 111 3166 115 3170
rect 135 3166 139 3170
rect 143 3166 147 3170
rect 319 3166 323 3170
rect 343 3166 347 3170
rect 519 3166 523 3170
rect 543 3166 547 3170
rect 1055 3250 1059 3254
rect 1095 3250 1099 3254
rect 1247 3330 1251 3334
rect 1295 3330 1299 3334
rect 1439 3330 1443 3334
rect 1463 3330 1467 3334
rect 1631 3330 1635 3334
rect 1639 3330 1643 3334
rect 1815 3330 1819 3334
rect 1823 3330 1827 3334
rect 2047 3362 2051 3366
rect 2447 3362 2451 3366
rect 2551 3362 2555 3366
rect 2567 3362 2571 3366
rect 2663 3362 2667 3366
rect 2719 3362 2723 3366
rect 2775 3362 2779 3366
rect 2871 3362 2875 3366
rect 2903 3362 2907 3366
rect 2007 3330 2011 3334
rect 2047 3282 2051 3286
rect 2415 3282 2419 3286
rect 2551 3282 2555 3286
rect 2567 3282 2571 3286
rect 1247 3250 1251 3254
rect 1271 3250 1275 3254
rect 1439 3250 1443 3254
rect 1447 3250 1451 3254
rect 1623 3250 1627 3254
rect 1631 3250 1635 3254
rect 719 3166 723 3170
rect 743 3166 747 3170
rect 911 3166 915 3170
rect 927 3166 931 3170
rect 1095 3166 1099 3170
rect 1103 3166 1107 3170
rect 1263 3166 1267 3170
rect 1271 3166 1275 3170
rect 1423 3166 1427 3170
rect 1447 3166 1451 3170
rect 111 3090 115 3094
rect 143 3090 147 3094
rect 263 3090 267 3094
rect 343 3090 347 3094
rect 439 3090 443 3094
rect 543 3090 547 3094
rect 615 3090 619 3094
rect 743 3090 747 3094
rect 799 3090 803 3094
rect 927 3090 931 3094
rect 975 3090 979 3094
rect 111 2990 115 2994
rect 263 2990 267 2994
rect 343 2990 347 2994
rect 439 2990 443 2994
rect 111 2914 115 2918
rect 207 2914 211 2918
rect 543 2990 547 2994
rect 615 2990 619 2994
rect 655 2990 659 2994
rect 783 2990 787 2994
rect 799 2990 803 2994
rect 1103 3090 1107 3094
rect 1143 3090 1147 3094
rect 1575 3166 1579 3170
rect 1623 3166 1627 3170
rect 1799 3250 1803 3254
rect 1823 3250 1827 3254
rect 2007 3250 2011 3254
rect 3023 3362 3027 3366
rect 3047 3362 3051 3366
rect 3175 3362 3179 3366
rect 3207 3362 3211 3366
rect 3751 3450 3755 3454
rect 3807 3450 3811 3454
rect 3943 3526 3947 3530
rect 3943 3450 3947 3454
rect 3327 3362 3331 3366
rect 3383 3362 3387 3366
rect 3479 3362 3483 3366
rect 3567 3362 3571 3366
rect 3631 3362 3635 3366
rect 3751 3362 3755 3366
rect 3783 3362 3787 3366
rect 2687 3282 2691 3286
rect 2719 3282 2723 3286
rect 2831 3282 2835 3286
rect 2871 3282 2875 3286
rect 2975 3282 2979 3286
rect 3023 3282 3027 3286
rect 3119 3282 3123 3286
rect 3175 3282 3179 3286
rect 3943 3362 3947 3366
rect 3255 3282 3259 3286
rect 3327 3282 3331 3286
rect 3383 3282 3387 3286
rect 3479 3282 3483 3286
rect 3503 3282 3507 3286
rect 3623 3282 3627 3286
rect 3631 3282 3635 3286
rect 3743 3282 3747 3286
rect 3783 3282 3787 3286
rect 3839 3282 3843 3286
rect 3943 3282 3947 3286
rect 2047 3194 2051 3198
rect 2247 3194 2251 3198
rect 2399 3194 2403 3198
rect 2415 3194 2419 3198
rect 2551 3194 2555 3198
rect 2559 3194 2563 3198
rect 1735 3166 1739 3170
rect 1799 3166 1803 3170
rect 2007 3166 2011 3170
rect 2047 3114 2051 3118
rect 2079 3114 2083 3118
rect 2223 3114 2227 3118
rect 2247 3114 2251 3118
rect 1263 3090 1267 3094
rect 1303 3090 1307 3094
rect 1423 3090 1427 3094
rect 1455 3090 1459 3094
rect 1575 3090 1579 3094
rect 1607 3090 1611 3094
rect 1735 3090 1739 3094
rect 1767 3090 1771 3094
rect 2007 3090 2011 3094
rect 2687 3194 2691 3198
rect 2727 3194 2731 3198
rect 2831 3194 2835 3198
rect 2903 3194 2907 3198
rect 2975 3194 2979 3198
rect 3079 3194 3083 3198
rect 3119 3194 3123 3198
rect 3255 3194 3259 3198
rect 3263 3194 3267 3198
rect 3383 3194 3387 3198
rect 3447 3194 3451 3198
rect 3503 3194 3507 3198
rect 3623 3194 3627 3198
rect 3631 3194 3635 3198
rect 3743 3194 3747 3198
rect 3815 3194 3819 3198
rect 3839 3194 3843 3198
rect 2375 3114 2379 3118
rect 2399 3114 2403 3118
rect 2527 3114 2531 3118
rect 2559 3114 2563 3118
rect 2687 3114 2691 3118
rect 2727 3114 2731 3118
rect 2855 3114 2859 3118
rect 2903 3114 2907 3118
rect 3039 3114 3043 3118
rect 3079 3114 3083 3118
rect 3231 3114 3235 3118
rect 3263 3114 3267 3118
rect 3431 3114 3435 3118
rect 3447 3114 3451 3118
rect 3631 3114 3635 3118
rect 2047 3030 2051 3034
rect 2071 3030 2075 3034
rect 2079 3030 2083 3034
rect 2183 3030 2187 3034
rect 2223 3030 2227 3034
rect 935 2990 939 2994
rect 975 2990 979 2994
rect 1103 2990 1107 2994
rect 1143 2990 1147 2994
rect 1295 2990 1299 2994
rect 1303 2990 1307 2994
rect 1455 2990 1459 2994
rect 1495 2990 1499 2994
rect 1607 2990 1611 2994
rect 1711 2990 1715 2994
rect 1767 2990 1771 2994
rect 1903 2990 1907 2994
rect 2007 2990 2011 2994
rect 2047 2950 2051 2954
rect 327 2914 331 2918
rect 343 2914 347 2918
rect 439 2914 443 2918
rect 447 2914 451 2918
rect 543 2914 547 2918
rect 575 2914 579 2918
rect 655 2914 659 2918
rect 703 2914 707 2918
rect 783 2914 787 2918
rect 847 2914 851 2918
rect 935 2914 939 2918
rect 111 2834 115 2838
rect 135 2834 139 2838
rect 207 2834 211 2838
rect 247 2834 251 2838
rect 327 2834 331 2838
rect 399 2834 403 2838
rect 447 2834 451 2838
rect 111 2750 115 2754
rect 135 2750 139 2754
rect 551 2834 555 2838
rect 575 2834 579 2838
rect 703 2834 707 2838
rect 711 2834 715 2838
rect 847 2834 851 2838
rect 879 2834 883 2838
rect 999 2914 1003 2918
rect 1103 2914 1107 2918
rect 1167 2914 1171 2918
rect 1295 2914 1299 2918
rect 1351 2914 1355 2918
rect 1495 2914 1499 2918
rect 1535 2914 1539 2918
rect 1711 2914 1715 2918
rect 1727 2914 1731 2918
rect 2071 2950 2075 2954
rect 2327 3030 2331 3034
rect 2375 3030 2379 3034
rect 2479 3030 2483 3034
rect 2527 3030 2531 3034
rect 2655 3030 2659 3034
rect 2687 3030 2691 3034
rect 2855 3030 2859 3034
rect 3639 3114 3643 3118
rect 3815 3114 3819 3118
rect 3839 3114 3843 3118
rect 3943 3194 3947 3198
rect 3943 3114 3947 3118
rect 3039 3030 3043 3034
rect 3087 3030 3091 3034
rect 3231 3030 3235 3034
rect 3335 3030 3339 3034
rect 3431 3030 3435 3034
rect 3599 3030 3603 3034
rect 3639 3030 3643 3034
rect 3839 3030 3843 3034
rect 2183 2950 2187 2954
rect 2263 2950 2267 2954
rect 2327 2950 2331 2954
rect 2479 2950 2483 2954
rect 2487 2950 2491 2954
rect 2655 2950 2659 2954
rect 2735 2950 2739 2954
rect 2855 2950 2859 2954
rect 2999 2950 3003 2954
rect 3087 2950 3091 2954
rect 3279 2950 3283 2954
rect 3335 2950 3339 2954
rect 3567 2950 3571 2954
rect 1903 2914 1907 2918
rect 2007 2914 2011 2918
rect 999 2834 1003 2838
rect 1047 2834 1051 2838
rect 1167 2834 1171 2838
rect 1223 2834 1227 2838
rect 247 2750 251 2754
rect 255 2750 259 2754
rect 399 2750 403 2754
rect 407 2750 411 2754
rect 551 2750 555 2754
rect 575 2750 579 2754
rect 711 2750 715 2754
rect 743 2750 747 2754
rect 879 2750 883 2754
rect 919 2750 923 2754
rect 1047 2750 1051 2754
rect 1087 2750 1091 2754
rect 111 2674 115 2678
rect 135 2674 139 2678
rect 167 2674 171 2678
rect 255 2674 259 2678
rect 359 2674 363 2678
rect 407 2674 411 2678
rect 559 2674 563 2678
rect 575 2674 579 2678
rect 743 2674 747 2678
rect 759 2674 763 2678
rect 919 2674 923 2678
rect 951 2674 955 2678
rect 1351 2834 1355 2838
rect 1399 2834 1403 2838
rect 1535 2834 1539 2838
rect 1575 2834 1579 2838
rect 1727 2834 1731 2838
rect 1751 2834 1755 2838
rect 1223 2750 1227 2754
rect 1255 2750 1259 2754
rect 1399 2750 1403 2754
rect 1423 2750 1427 2754
rect 1575 2750 1579 2754
rect 1599 2750 1603 2754
rect 2047 2866 2051 2870
rect 2071 2866 2075 2870
rect 2263 2866 2267 2870
rect 1903 2834 1907 2838
rect 2007 2834 2011 2838
rect 3599 2950 3603 2954
rect 3839 2950 3843 2954
rect 3943 3030 3947 3034
rect 3943 2950 3947 2954
rect 2487 2866 2491 2870
rect 2671 2866 2675 2870
rect 2735 2866 2739 2870
rect 2887 2866 2891 2870
rect 2999 2866 3003 2870
rect 3095 2866 3099 2870
rect 3279 2866 3283 2870
rect 3287 2866 3291 2870
rect 3479 2866 3483 2870
rect 3567 2866 3571 2870
rect 3671 2866 3675 2870
rect 3839 2866 3843 2870
rect 3943 2866 3947 2870
rect 2047 2790 2051 2794
rect 2071 2790 2075 2794
rect 2199 2790 2203 2794
rect 2343 2790 2347 2794
rect 2479 2790 2483 2794
rect 2607 2790 2611 2794
rect 2671 2790 2675 2794
rect 1751 2750 1755 2754
rect 1903 2750 1907 2754
rect 2007 2750 2011 2754
rect 1087 2674 1091 2678
rect 1143 2674 1147 2678
rect 1255 2674 1259 2678
rect 1327 2674 1331 2678
rect 111 2582 115 2586
rect 167 2582 171 2586
rect 359 2582 363 2586
rect 559 2582 563 2586
rect 575 2582 579 2586
rect 687 2582 691 2586
rect 759 2582 763 2586
rect 807 2582 811 2586
rect 935 2582 939 2586
rect 951 2582 955 2586
rect 1071 2582 1075 2586
rect 1143 2582 1147 2586
rect 111 2502 115 2506
rect 503 2502 507 2506
rect 575 2502 579 2506
rect 607 2502 611 2506
rect 687 2502 691 2506
rect 2047 2694 2051 2698
rect 2071 2694 2075 2698
rect 2095 2694 2099 2698
rect 1423 2674 1427 2678
rect 1511 2674 1515 2678
rect 1599 2674 1603 2678
rect 1703 2674 1707 2678
rect 2007 2674 2011 2678
rect 1207 2582 1211 2586
rect 1327 2582 1331 2586
rect 1351 2582 1355 2586
rect 1495 2582 1499 2586
rect 1511 2582 1515 2586
rect 1647 2582 1651 2586
rect 1703 2582 1707 2586
rect 719 2502 723 2506
rect 807 2502 811 2506
rect 847 2502 851 2506
rect 935 2502 939 2506
rect 983 2502 987 2506
rect 1071 2502 1075 2506
rect 1127 2502 1131 2506
rect 111 2410 115 2414
rect 503 2410 507 2414
rect 535 2410 539 2414
rect 607 2410 611 2414
rect 1207 2502 1211 2506
rect 1279 2502 1283 2506
rect 1351 2502 1355 2506
rect 2199 2694 2203 2698
rect 2263 2694 2267 2698
rect 2343 2694 2347 2698
rect 2727 2790 2731 2794
rect 2839 2790 2843 2794
rect 2887 2790 2891 2794
rect 2943 2790 2947 2794
rect 3047 2790 3051 2794
rect 3095 2790 3099 2794
rect 3143 2790 3147 2794
rect 3239 2790 3243 2794
rect 3287 2790 3291 2794
rect 3343 2790 3347 2794
rect 3447 2790 3451 2794
rect 3479 2790 3483 2794
rect 3551 2790 3555 2794
rect 3647 2790 3651 2794
rect 3671 2790 3675 2794
rect 3743 2790 3747 2794
rect 3839 2790 3843 2794
rect 3943 2790 3947 2794
rect 2439 2694 2443 2698
rect 2479 2694 2483 2698
rect 2607 2694 2611 2698
rect 2615 2694 2619 2698
rect 2727 2694 2731 2698
rect 2783 2694 2787 2698
rect 2839 2694 2843 2698
rect 2047 2610 2051 2614
rect 2095 2610 2099 2614
rect 2215 2610 2219 2614
rect 2263 2610 2267 2614
rect 2367 2610 2371 2614
rect 2439 2610 2443 2614
rect 2519 2610 2523 2614
rect 2615 2610 2619 2614
rect 2671 2610 2675 2614
rect 1799 2582 1803 2586
rect 2007 2582 2011 2586
rect 1431 2502 1435 2506
rect 1495 2502 1499 2506
rect 2047 2530 2051 2534
rect 2095 2530 2099 2534
rect 2215 2530 2219 2534
rect 2343 2530 2347 2534
rect 1583 2502 1587 2506
rect 1647 2502 1651 2506
rect 1743 2502 1747 2506
rect 1799 2502 1803 2506
rect 1903 2502 1907 2506
rect 2007 2502 2011 2506
rect 671 2410 675 2414
rect 719 2410 723 2414
rect 815 2410 819 2414
rect 847 2410 851 2414
rect 959 2410 963 2414
rect 983 2410 987 2414
rect 1103 2410 1107 2414
rect 1127 2410 1131 2414
rect 1247 2410 1251 2414
rect 1279 2410 1283 2414
rect 1391 2410 1395 2414
rect 1431 2410 1435 2414
rect 1527 2410 1531 2414
rect 1583 2410 1587 2414
rect 1655 2410 1659 2414
rect 1743 2410 1747 2414
rect 1791 2410 1795 2414
rect 1903 2410 1907 2414
rect 111 2330 115 2334
rect 535 2330 539 2334
rect 647 2330 651 2334
rect 671 2330 675 2334
rect 767 2330 771 2334
rect 815 2330 819 2334
rect 111 2250 115 2254
rect 415 2250 419 2254
rect 895 2330 899 2334
rect 959 2330 963 2334
rect 1031 2330 1035 2334
rect 1103 2330 1107 2334
rect 1167 2330 1171 2334
rect 1247 2330 1251 2334
rect 1295 2330 1299 2334
rect 2047 2442 2051 2446
rect 2071 2442 2075 2446
rect 2095 2442 2099 2446
rect 2007 2410 2011 2414
rect 2367 2530 2371 2534
rect 2943 2694 2947 2698
rect 3047 2694 3051 2698
rect 3095 2694 3099 2698
rect 3143 2694 3147 2698
rect 3239 2694 3243 2698
rect 3343 2694 3347 2698
rect 3383 2694 3387 2698
rect 3447 2694 3451 2698
rect 3535 2694 3539 2698
rect 3551 2694 3555 2698
rect 3647 2694 3651 2698
rect 3743 2694 3747 2698
rect 3839 2694 3843 2698
rect 3943 2694 3947 2698
rect 2783 2610 2787 2614
rect 2815 2610 2819 2614
rect 2943 2610 2947 2614
rect 2951 2610 2955 2614
rect 3087 2610 3091 2614
rect 3095 2610 3099 2614
rect 3223 2610 3227 2614
rect 3239 2610 3243 2614
rect 3367 2610 3371 2614
rect 3383 2610 3387 2614
rect 3535 2610 3539 2614
rect 3943 2610 3947 2614
rect 2471 2530 2475 2534
rect 2519 2530 2523 2534
rect 2599 2530 2603 2534
rect 2671 2530 2675 2534
rect 2719 2530 2723 2534
rect 2191 2442 2195 2446
rect 2215 2442 2219 2446
rect 2319 2442 2323 2446
rect 2343 2442 2347 2446
rect 2439 2442 2443 2446
rect 2471 2442 2475 2446
rect 2559 2442 2563 2446
rect 2599 2442 2603 2446
rect 1391 2330 1395 2334
rect 1423 2330 1427 2334
rect 1527 2330 1531 2334
rect 1551 2330 1555 2334
rect 1655 2330 1659 2334
rect 1671 2330 1675 2334
rect 1791 2330 1795 2334
rect 1799 2330 1803 2334
rect 535 2250 539 2254
rect 647 2250 651 2254
rect 671 2250 675 2254
rect 767 2250 771 2254
rect 823 2250 827 2254
rect 895 2250 899 2254
rect 991 2250 995 2254
rect 1031 2250 1035 2254
rect 1167 2250 1171 2254
rect 1175 2250 1179 2254
rect 1295 2250 1299 2254
rect 1367 2250 1371 2254
rect 1423 2250 1427 2254
rect 1551 2250 1555 2254
rect 1567 2250 1571 2254
rect 111 2166 115 2170
rect 135 2166 139 2170
rect 247 2166 251 2170
rect 391 2166 395 2170
rect 415 2166 419 2170
rect 535 2166 539 2170
rect 551 2166 555 2170
rect 671 2166 675 2170
rect 711 2166 715 2170
rect 2047 2362 2051 2366
rect 2071 2362 2075 2366
rect 2167 2362 2171 2366
rect 2191 2362 2195 2366
rect 1903 2330 1907 2334
rect 2007 2330 2011 2334
rect 2815 2530 2819 2534
rect 2839 2530 2843 2534
rect 2951 2530 2955 2534
rect 2967 2530 2971 2534
rect 3087 2530 3091 2534
rect 3095 2530 3099 2534
rect 3223 2530 3227 2534
rect 3367 2530 3371 2534
rect 3943 2530 3947 2534
rect 2679 2442 2683 2446
rect 2719 2442 2723 2446
rect 2791 2442 2795 2446
rect 2839 2442 2843 2446
rect 2911 2442 2915 2446
rect 2967 2442 2971 2446
rect 3031 2442 3035 2446
rect 3095 2442 3099 2446
rect 3151 2442 3155 2446
rect 3223 2442 3227 2446
rect 3943 2442 3947 2446
rect 2319 2362 2323 2366
rect 2359 2362 2363 2366
rect 2047 2286 2051 2290
rect 2071 2286 2075 2290
rect 2167 2286 2171 2290
rect 2287 2286 2291 2290
rect 2439 2362 2443 2366
rect 2535 2362 2539 2366
rect 2559 2362 2563 2366
rect 2679 2362 2683 2366
rect 2703 2362 2707 2366
rect 2791 2362 2795 2366
rect 2871 2362 2875 2366
rect 2911 2362 2915 2366
rect 3031 2362 3035 2366
rect 3151 2362 3155 2366
rect 3199 2362 3203 2366
rect 3943 2362 3947 2366
rect 2359 2286 2363 2290
rect 2423 2286 2427 2290
rect 2535 2286 2539 2290
rect 2559 2286 2563 2290
rect 2703 2286 2707 2290
rect 2839 2286 2843 2290
rect 2871 2286 2875 2290
rect 2983 2286 2987 2290
rect 3031 2286 3035 2290
rect 1671 2250 1675 2254
rect 1767 2250 1771 2254
rect 1799 2250 1803 2254
rect 1903 2250 1907 2254
rect 2007 2250 2011 2254
rect 823 2166 827 2170
rect 871 2166 875 2170
rect 991 2166 995 2170
rect 1031 2166 1035 2170
rect 1175 2166 1179 2170
rect 1191 2166 1195 2170
rect 111 2082 115 2086
rect 135 2082 139 2086
rect 247 2082 251 2086
rect 391 2082 395 2086
rect 399 2082 403 2086
rect 551 2082 555 2086
rect 703 2082 707 2086
rect 711 2082 715 2086
rect 847 2082 851 2086
rect 871 2082 875 2086
rect 1351 2166 1355 2170
rect 1367 2166 1371 2170
rect 1511 2166 1515 2170
rect 1567 2166 1571 2170
rect 1679 2166 1683 2170
rect 2047 2210 2051 2214
rect 2071 2210 2075 2214
rect 1767 2166 1771 2170
rect 2007 2166 2011 2170
rect 2167 2210 2171 2214
rect 2287 2210 2291 2214
rect 2295 2210 2299 2214
rect 3127 2286 3131 2290
rect 3199 2286 3203 2290
rect 3271 2286 3275 2290
rect 3943 2286 3947 2290
rect 2423 2210 2427 2214
rect 2503 2210 2507 2214
rect 2559 2210 2563 2214
rect 2687 2210 2691 2214
rect 2703 2210 2707 2214
rect 2839 2210 2843 2214
rect 2863 2210 2867 2214
rect 2983 2210 2987 2214
rect 3023 2210 3027 2214
rect 3127 2210 3131 2214
rect 3175 2210 3179 2214
rect 2047 2110 2051 2114
rect 2071 2110 2075 2114
rect 2295 2110 2299 2114
rect 2399 2110 2403 2114
rect 2495 2110 2499 2114
rect 2503 2110 2507 2114
rect 2591 2110 2595 2114
rect 2687 2110 2691 2114
rect 991 2082 995 2086
rect 1031 2082 1035 2086
rect 1127 2082 1131 2086
rect 1191 2082 1195 2086
rect 1255 2082 1259 2086
rect 1351 2082 1355 2086
rect 1383 2082 1387 2086
rect 1511 2082 1515 2086
rect 1519 2082 1523 2086
rect 1679 2082 1683 2086
rect 2007 2082 2011 2086
rect 111 1990 115 1994
rect 135 1990 139 1994
rect 231 1990 235 1994
rect 247 1990 251 1994
rect 391 1990 395 1994
rect 399 1990 403 1994
rect 551 1990 555 1994
rect 567 1990 571 1994
rect 703 1990 707 1994
rect 751 1990 755 1994
rect 847 1990 851 1994
rect 2947 2120 2951 2124
rect 2783 2110 2787 2114
rect 2863 2110 2867 2114
rect 2879 2110 2883 2114
rect 3271 2210 3275 2214
rect 3319 2210 3323 2214
rect 3471 2210 3475 2214
rect 3943 2210 3947 2214
rect 3439 2120 3443 2124
rect 2975 2110 2979 2114
rect 3023 2110 3027 2114
rect 3071 2110 3075 2114
rect 3167 2110 3171 2114
rect 3175 2110 3179 2114
rect 3263 2110 3267 2114
rect 3319 2110 3323 2114
rect 3359 2110 3363 2114
rect 3455 2110 3459 2114
rect 3471 2110 3475 2114
rect 3551 2110 3555 2114
rect 3647 2110 3651 2114
rect 3743 2110 3747 2114
rect 3839 2110 3843 2114
rect 3943 2110 3947 2114
rect 2047 2034 2051 2038
rect 2191 2034 2195 2038
rect 2399 2034 2403 2038
rect 2495 2034 2499 2038
rect 2591 2034 2595 2038
rect 2647 2034 2651 2038
rect 2687 2034 2691 2038
rect 2783 2034 2787 2038
rect 2879 2034 2883 2038
rect 2919 2034 2923 2038
rect 2975 2034 2979 2038
rect 3071 2034 3075 2038
rect 3167 2034 3171 2038
rect 3215 2034 3219 2038
rect 3263 2034 3267 2038
rect 3359 2034 3363 2038
rect 3455 2034 3459 2038
rect 3527 2034 3531 2038
rect 3551 2034 3555 2038
rect 3647 2034 3651 2038
rect 3743 2034 3747 2038
rect 3839 2034 3843 2038
rect 943 1990 947 1994
rect 991 1990 995 1994
rect 1127 1990 1131 1994
rect 1135 1990 1139 1994
rect 1255 1990 1259 1994
rect 1335 1990 1339 1994
rect 1383 1990 1387 1994
rect 1519 1990 1523 1994
rect 1543 1990 1547 1994
rect 2007 1990 2011 1994
rect 111 1914 115 1918
rect 1203 1928 1207 1932
rect 231 1914 235 1918
rect 391 1914 395 1918
rect 511 1914 515 1918
rect 567 1914 571 1918
rect 623 1914 627 1918
rect 743 1914 747 1918
rect 751 1914 755 1918
rect 863 1914 867 1918
rect 943 1914 947 1918
rect 983 1914 987 1918
rect 1103 1914 1107 1918
rect 1135 1914 1139 1918
rect 1223 1914 1227 1918
rect 1335 1914 1339 1918
rect 111 1830 115 1834
rect 511 1830 515 1834
rect 615 1830 619 1834
rect 623 1830 627 1834
rect 711 1830 715 1834
rect 743 1830 747 1834
rect 815 1830 819 1834
rect 863 1830 867 1834
rect 927 1830 931 1834
rect 983 1830 987 1834
rect 1039 1830 1043 1834
rect 1103 1830 1107 1834
rect 2047 1946 2051 1950
rect 2071 1946 2075 1950
rect 2191 1946 2195 1950
rect 2239 1946 2243 1950
rect 2399 1946 2403 1950
rect 2447 1946 2451 1950
rect 1459 1928 1463 1932
rect 1455 1914 1459 1918
rect 1543 1914 1547 1918
rect 1575 1914 1579 1918
rect 1695 1914 1699 1918
rect 2007 1914 2011 1918
rect 3943 2034 3947 2038
rect 2647 1946 2651 1950
rect 2671 1946 2675 1950
rect 2895 1946 2899 1950
rect 2919 1946 2923 1950
rect 3127 1946 3131 1950
rect 3215 1946 3219 1950
rect 3359 1946 3363 1950
rect 3527 1946 3531 1950
rect 3591 1946 3595 1950
rect 3831 1946 3835 1950
rect 3839 1946 3843 1950
rect 3943 1946 3947 1950
rect 1159 1830 1163 1834
rect 111 1754 115 1758
rect 367 1754 371 1758
rect 495 1754 499 1758
rect 615 1754 619 1758
rect 1223 1830 1227 1834
rect 1279 1830 1283 1834
rect 1335 1830 1339 1834
rect 1399 1830 1403 1834
rect 1455 1830 1459 1834
rect 1519 1830 1523 1834
rect 1575 1830 1579 1834
rect 1639 1830 1643 1834
rect 1695 1830 1699 1834
rect 2047 1870 2051 1874
rect 2071 1870 2075 1874
rect 2199 1870 2203 1874
rect 2239 1870 2243 1874
rect 2007 1830 2011 1834
rect 2047 1790 2051 1794
rect 639 1754 643 1758
rect 111 1674 115 1678
rect 135 1674 139 1678
rect 247 1674 251 1678
rect 367 1674 371 1678
rect 399 1674 403 1678
rect 711 1754 715 1758
rect 799 1754 803 1758
rect 815 1754 819 1758
rect 927 1754 931 1758
rect 967 1754 971 1758
rect 1039 1754 1043 1758
rect 1143 1754 1147 1758
rect 1159 1754 1163 1758
rect 1279 1754 1283 1758
rect 1327 1754 1331 1758
rect 683 1736 687 1740
rect 919 1736 923 1740
rect 2071 1790 2075 1794
rect 1399 1754 1403 1758
rect 1511 1754 1515 1758
rect 2367 1870 2371 1874
rect 2447 1870 2451 1874
rect 2543 1870 2547 1874
rect 2671 1870 2675 1874
rect 2719 1870 2723 1874
rect 2887 1870 2891 1874
rect 2895 1870 2899 1874
rect 3039 1870 3043 1874
rect 3127 1870 3131 1874
rect 3183 1870 3187 1874
rect 3319 1870 3323 1874
rect 3359 1870 3363 1874
rect 3455 1870 3459 1874
rect 3583 1870 3587 1874
rect 3591 1870 3595 1874
rect 3711 1870 3715 1874
rect 3831 1870 3835 1874
rect 3839 1870 3843 1874
rect 2183 1790 2187 1794
rect 2199 1790 2203 1794
rect 2327 1790 2331 1794
rect 2367 1790 2371 1794
rect 2487 1790 2491 1794
rect 2543 1790 2547 1794
rect 2655 1790 2659 1794
rect 2719 1790 2723 1794
rect 2831 1790 2835 1794
rect 2887 1790 2891 1794
rect 3023 1790 3027 1794
rect 3039 1790 3043 1794
rect 3183 1790 3187 1794
rect 3223 1790 3227 1794
rect 3319 1790 3323 1794
rect 3431 1790 3435 1794
rect 3455 1790 3459 1794
rect 3583 1790 3587 1794
rect 3647 1790 3651 1794
rect 3711 1790 3715 1794
rect 3839 1790 3843 1794
rect 1519 1754 1523 1758
rect 1639 1754 1643 1758
rect 1703 1754 1707 1758
rect 2007 1754 2011 1758
rect 495 1674 499 1678
rect 567 1674 571 1678
rect 639 1674 643 1678
rect 743 1674 747 1678
rect 799 1674 803 1678
rect 935 1674 939 1678
rect 967 1674 971 1678
rect 111 1594 115 1598
rect 135 1594 139 1598
rect 1135 1674 1139 1678
rect 1143 1674 1147 1678
rect 1327 1674 1331 1678
rect 1343 1674 1347 1678
rect 1511 1674 1515 1678
rect 1551 1674 1555 1678
rect 1703 1674 1707 1678
rect 2047 1706 2051 1710
rect 2071 1706 2075 1710
rect 2183 1706 2187 1710
rect 2223 1706 2227 1710
rect 2327 1706 2331 1710
rect 2439 1706 2443 1710
rect 2487 1706 2491 1710
rect 2559 1706 2563 1710
rect 1767 1674 1771 1678
rect 2007 1674 2011 1678
rect 247 1594 251 1598
rect 255 1594 259 1598
rect 399 1594 403 1598
rect 423 1594 427 1598
rect 567 1594 571 1598
rect 615 1594 619 1598
rect 743 1594 747 1598
rect 831 1594 835 1598
rect 935 1594 939 1598
rect 1063 1594 1067 1598
rect 1135 1594 1139 1598
rect 1311 1594 1315 1598
rect 1343 1594 1347 1598
rect 111 1514 115 1518
rect 135 1514 139 1518
rect 239 1514 243 1518
rect 255 1514 259 1518
rect 407 1514 411 1518
rect 423 1514 427 1518
rect 583 1514 587 1518
rect 615 1514 619 1518
rect 775 1514 779 1518
rect 831 1514 835 1518
rect 2655 1706 2659 1710
rect 2687 1706 2691 1710
rect 2823 1706 2827 1710
rect 2831 1706 2835 1710
rect 2967 1706 2971 1710
rect 3023 1706 3027 1710
rect 3127 1706 3131 1710
rect 3223 1706 3227 1710
rect 3303 1706 3307 1710
rect 3431 1706 3435 1710
rect 3487 1706 3491 1710
rect 3647 1706 3651 1710
rect 3671 1706 3675 1710
rect 3943 1870 3947 1874
rect 3943 1790 3947 1794
rect 3839 1706 3843 1710
rect 2047 1626 2051 1630
rect 2223 1626 2227 1630
rect 2327 1626 2331 1630
rect 2391 1626 2395 1630
rect 2439 1626 2443 1630
rect 2503 1626 2507 1630
rect 2559 1626 2563 1630
rect 2615 1626 2619 1630
rect 2687 1626 2691 1630
rect 2735 1626 2739 1630
rect 2823 1626 2827 1630
rect 2855 1626 2859 1630
rect 2967 1626 2971 1630
rect 2975 1626 2979 1630
rect 3095 1626 3099 1630
rect 3127 1626 3131 1630
rect 3215 1626 3219 1630
rect 3303 1626 3307 1630
rect 3335 1626 3339 1630
rect 3455 1626 3459 1630
rect 3487 1626 3491 1630
rect 3671 1626 3675 1630
rect 1551 1594 1555 1598
rect 1567 1594 1571 1598
rect 1767 1594 1771 1598
rect 1831 1594 1835 1598
rect 2007 1594 2011 1598
rect 967 1514 971 1518
rect 1063 1514 1067 1518
rect 1159 1514 1163 1518
rect 1311 1514 1315 1518
rect 1351 1514 1355 1518
rect 1543 1514 1547 1518
rect 1567 1514 1571 1518
rect 1735 1514 1739 1518
rect 2047 1550 2051 1554
rect 2391 1550 2395 1554
rect 2503 1550 2507 1554
rect 2543 1550 2547 1554
rect 2615 1550 2619 1554
rect 2671 1550 2675 1554
rect 2735 1550 2739 1554
rect 2799 1550 2803 1554
rect 1831 1514 1835 1518
rect 1903 1514 1907 1518
rect 2007 1514 2011 1518
rect 111 1430 115 1434
rect 239 1430 243 1434
rect 407 1430 411 1434
rect 463 1430 467 1434
rect 583 1430 587 1434
rect 711 1430 715 1434
rect 775 1430 779 1434
rect 855 1430 859 1434
rect 967 1430 971 1434
rect 1007 1430 1011 1434
rect 1159 1430 1163 1434
rect 1167 1430 1171 1434
rect 1335 1430 1339 1434
rect 1351 1430 1355 1434
rect 111 1354 115 1358
rect 463 1354 467 1358
rect 583 1354 587 1358
rect 655 1354 659 1358
rect 711 1354 715 1358
rect 767 1354 771 1358
rect 855 1354 859 1358
rect 887 1354 891 1358
rect 1007 1354 1011 1358
rect 1015 1354 1019 1358
rect 2855 1550 2859 1554
rect 2935 1550 2939 1554
rect 2975 1550 2979 1554
rect 3071 1550 3075 1554
rect 3095 1550 3099 1554
rect 3207 1550 3211 1554
rect 3215 1550 3219 1554
rect 3335 1550 3339 1554
rect 1511 1430 1515 1434
rect 1543 1430 1547 1434
rect 1687 1430 1691 1434
rect 1735 1430 1739 1434
rect 1871 1430 1875 1434
rect 1903 1430 1907 1434
rect 1143 1354 1147 1358
rect 1167 1354 1171 1358
rect 1279 1354 1283 1358
rect 1335 1354 1339 1358
rect 1415 1354 1419 1358
rect 1511 1354 1515 1358
rect 1559 1354 1563 1358
rect 1687 1354 1691 1358
rect 1703 1354 1707 1358
rect 2047 1462 2051 1466
rect 2519 1462 2523 1466
rect 2543 1462 2547 1466
rect 2631 1462 2635 1466
rect 2671 1462 2675 1466
rect 2759 1462 2763 1466
rect 2799 1462 2803 1466
rect 2895 1462 2899 1466
rect 2935 1462 2939 1466
rect 3031 1462 3035 1466
rect 3071 1462 3075 1466
rect 2007 1430 2011 1434
rect 3455 1550 3459 1554
rect 3463 1550 3467 1554
rect 3591 1550 3595 1554
rect 3727 1550 3731 1554
rect 3943 1706 3947 1710
rect 3839 1626 3843 1630
rect 3839 1550 3843 1554
rect 3175 1462 3179 1466
rect 3207 1462 3211 1466
rect 3311 1462 3315 1466
rect 3335 1462 3339 1466
rect 3447 1462 3451 1466
rect 3463 1462 3467 1466
rect 3583 1462 3587 1466
rect 3591 1462 3595 1466
rect 3719 1462 3723 1466
rect 3727 1462 3731 1466
rect 2047 1386 2051 1390
rect 2399 1386 2403 1390
rect 2519 1386 2523 1390
rect 2535 1386 2539 1390
rect 2631 1386 2635 1390
rect 2679 1386 2683 1390
rect 1847 1354 1851 1358
rect 1871 1354 1875 1358
rect 2007 1354 2011 1358
rect 111 1274 115 1278
rect 439 1274 443 1278
rect 551 1274 555 1278
rect 655 1274 659 1278
rect 671 1274 675 1278
rect 767 1274 771 1278
rect 799 1274 803 1278
rect 887 1274 891 1278
rect 935 1274 939 1278
rect 1015 1274 1019 1278
rect 1079 1274 1083 1278
rect 1143 1274 1147 1278
rect 1231 1274 1235 1278
rect 1279 1274 1283 1278
rect 1391 1274 1395 1278
rect 1415 1274 1419 1278
rect 111 1198 115 1202
rect 167 1198 171 1202
rect 303 1198 307 1202
rect 439 1198 443 1202
rect 463 1198 467 1202
rect 551 1198 555 1202
rect 631 1198 635 1202
rect 671 1198 675 1202
rect 1551 1274 1555 1278
rect 1559 1274 1563 1278
rect 2047 1306 2051 1310
rect 2247 1306 2251 1310
rect 2375 1306 2379 1310
rect 2399 1306 2403 1310
rect 1703 1274 1707 1278
rect 1719 1274 1723 1278
rect 1847 1274 1851 1278
rect 2007 1274 2011 1278
rect 2759 1386 2763 1390
rect 2823 1386 2827 1390
rect 2895 1386 2899 1390
rect 2967 1386 2971 1390
rect 3031 1386 3035 1390
rect 3111 1386 3115 1390
rect 3175 1386 3179 1390
rect 3255 1386 3259 1390
rect 3311 1386 3315 1390
rect 3407 1386 3411 1390
rect 3447 1386 3451 1390
rect 3559 1386 3563 1390
rect 3583 1386 3587 1390
rect 3711 1386 3715 1390
rect 3719 1386 3723 1390
rect 2511 1306 2515 1310
rect 2535 1306 2539 1310
rect 2647 1306 2651 1310
rect 2679 1306 2683 1310
rect 2791 1306 2795 1310
rect 2823 1306 2827 1310
rect 2943 1306 2947 1310
rect 2967 1306 2971 1310
rect 3839 1462 3843 1466
rect 3943 1626 3947 1630
rect 3943 1550 3947 1554
rect 3943 1462 3947 1466
rect 3839 1386 3843 1390
rect 3111 1306 3115 1310
rect 3255 1306 3259 1310
rect 3287 1306 3291 1310
rect 3407 1306 3411 1310
rect 3471 1306 3475 1310
rect 3559 1306 3563 1310
rect 3663 1306 3667 1310
rect 3711 1306 3715 1310
rect 3839 1306 3843 1310
rect 3943 1386 3947 1390
rect 3943 1306 3947 1310
rect 799 1198 803 1202
rect 807 1198 811 1202
rect 935 1198 939 1202
rect 983 1198 987 1202
rect 1079 1198 1083 1202
rect 1159 1198 1163 1202
rect 1231 1198 1235 1202
rect 1335 1198 1339 1202
rect 1391 1198 1395 1202
rect 1511 1198 1515 1202
rect 1551 1198 1555 1202
rect 1695 1198 1699 1202
rect 1719 1198 1723 1202
rect 2047 1226 2051 1230
rect 2071 1226 2075 1230
rect 2183 1226 2187 1230
rect 2247 1226 2251 1230
rect 2303 1226 2307 1230
rect 2007 1198 2011 1202
rect 111 1118 115 1122
rect 135 1118 139 1122
rect 167 1118 171 1122
rect 239 1118 243 1122
rect 303 1118 307 1122
rect 375 1118 379 1122
rect 463 1118 467 1122
rect 527 1118 531 1122
rect 631 1118 635 1122
rect 111 1042 115 1046
rect 135 1042 139 1046
rect 695 1118 699 1122
rect 807 1118 811 1122
rect 863 1118 867 1122
rect 983 1118 987 1122
rect 1039 1118 1043 1122
rect 1159 1118 1163 1122
rect 1215 1118 1219 1122
rect 2047 1146 2051 1150
rect 2071 1146 2075 1150
rect 2183 1146 2187 1150
rect 2199 1146 2203 1150
rect 2375 1226 2379 1230
rect 2431 1226 2435 1230
rect 2511 1226 2515 1230
rect 2559 1226 2563 1230
rect 2647 1226 2651 1230
rect 2711 1226 2715 1230
rect 2791 1226 2795 1230
rect 2887 1226 2891 1230
rect 2943 1226 2947 1230
rect 3087 1226 3091 1230
rect 3111 1226 3115 1230
rect 3287 1226 3291 1230
rect 3311 1226 3315 1230
rect 3471 1226 3475 1230
rect 3543 1226 3547 1230
rect 2303 1146 2307 1150
rect 2351 1146 2355 1150
rect 2431 1146 2435 1150
rect 2511 1146 2515 1150
rect 2559 1146 2563 1150
rect 2679 1146 2683 1150
rect 2711 1146 2715 1150
rect 1335 1118 1339 1122
rect 1391 1118 1395 1122
rect 1511 1118 1515 1122
rect 1567 1118 1571 1122
rect 1695 1118 1699 1122
rect 1743 1118 1747 1122
rect 1903 1118 1907 1122
rect 2007 1118 2011 1122
rect 239 1042 243 1046
rect 287 1042 291 1046
rect 375 1042 379 1046
rect 471 1042 475 1046
rect 527 1042 531 1046
rect 655 1042 659 1046
rect 695 1042 699 1046
rect 839 1042 843 1046
rect 863 1042 867 1046
rect 111 962 115 966
rect 135 962 139 966
rect 1015 1042 1019 1046
rect 1039 1042 1043 1046
rect 1199 1042 1203 1046
rect 1215 1042 1219 1046
rect 1383 1042 1387 1046
rect 1391 1042 1395 1046
rect 3663 1226 3667 1230
rect 3783 1226 3787 1230
rect 3839 1226 3843 1230
rect 3943 1226 3947 1230
rect 2871 1146 2875 1150
rect 2887 1146 2891 1150
rect 3087 1146 3091 1150
rect 3311 1146 3315 1150
rect 3319 1146 3323 1150
rect 3543 1146 3547 1150
rect 3559 1146 3563 1150
rect 2047 1058 2051 1062
rect 2071 1058 2075 1062
rect 1567 1042 1571 1046
rect 1743 1042 1747 1046
rect 1903 1042 1907 1046
rect 2007 1042 2011 1046
rect 287 962 291 966
rect 295 962 299 966
rect 471 962 475 966
rect 639 962 643 966
rect 655 962 659 966
rect 799 962 803 966
rect 839 962 843 966
rect 951 962 955 966
rect 111 886 115 890
rect 135 886 139 890
rect 159 886 163 890
rect 295 886 299 890
rect 319 886 323 890
rect 1015 962 1019 966
rect 1087 962 1091 966
rect 1199 962 1203 966
rect 1223 962 1227 966
rect 1359 962 1363 966
rect 1383 962 1387 966
rect 1495 962 1499 966
rect 1567 962 1571 966
rect 471 886 475 890
rect 615 886 619 890
rect 639 886 643 890
rect 111 810 115 814
rect 159 810 163 814
rect 223 810 227 814
rect 319 810 323 814
rect 383 810 387 814
rect 471 810 475 814
rect 535 810 539 814
rect 111 730 115 734
rect 223 730 227 734
rect 311 730 315 734
rect 383 730 387 734
rect 751 886 755 890
rect 799 886 803 890
rect 879 886 883 890
rect 951 886 955 890
rect 999 886 1003 890
rect 1087 886 1091 890
rect 1111 886 1115 890
rect 1223 886 1227 890
rect 1231 886 1235 890
rect 2199 1058 2203 1062
rect 2263 1058 2267 1062
rect 2351 1058 2355 1062
rect 2487 1058 2491 1062
rect 2511 1058 2515 1062
rect 2679 1058 2683 1062
rect 2703 1058 2707 1062
rect 2871 1058 2875 1062
rect 2919 1058 2923 1062
rect 3087 1058 3091 1062
rect 3119 1058 3123 1062
rect 3311 1058 3315 1062
rect 3319 1058 3323 1062
rect 2047 978 2051 982
rect 2071 978 2075 982
rect 2263 978 2267 982
rect 2303 978 2307 982
rect 2455 978 2459 982
rect 2487 978 2491 982
rect 2615 978 2619 982
rect 2703 978 2707 982
rect 2783 978 2787 982
rect 2919 978 2923 982
rect 2951 978 2955 982
rect 2007 962 2011 966
rect 3495 1058 3499 1062
rect 3559 1058 3563 1062
rect 3679 1058 3683 1062
rect 3783 1146 3787 1150
rect 3807 1146 3811 1150
rect 3943 1146 3947 1150
rect 3807 1058 3811 1062
rect 3839 1058 3843 1062
rect 3111 978 3115 982
rect 3119 978 3123 982
rect 3263 978 3267 982
rect 3311 978 3315 982
rect 3415 978 3419 982
rect 3495 978 3499 982
rect 3943 1058 3947 1062
rect 3559 978 3563 982
rect 3679 978 3683 982
rect 3711 978 3715 982
rect 3839 978 3843 982
rect 2047 898 2051 902
rect 2303 898 2307 902
rect 2455 898 2459 902
rect 2559 898 2563 902
rect 2615 898 2619 902
rect 2679 898 2683 902
rect 2783 898 2787 902
rect 2807 898 2811 902
rect 1351 886 1355 890
rect 1359 886 1363 890
rect 1495 886 1499 890
rect 2007 886 2011 890
rect 615 810 619 814
rect 2943 898 2947 902
rect 2951 898 2955 902
rect 3079 898 3083 902
rect 3111 898 3115 902
rect 3207 898 3211 902
rect 3263 898 3267 902
rect 3335 898 3339 902
rect 3415 898 3419 902
rect 3463 898 3467 902
rect 3559 898 3563 902
rect 3591 898 3595 902
rect 2047 818 2051 822
rect 2335 818 2339 822
rect 2471 818 2475 822
rect 2559 818 2563 822
rect 2615 818 2619 822
rect 2679 818 2683 822
rect 2767 818 2771 822
rect 2807 818 2811 822
rect 2919 818 2923 822
rect 2943 818 2947 822
rect 679 810 683 814
rect 751 810 755 814
rect 815 810 819 814
rect 879 810 883 814
rect 951 810 955 814
rect 999 810 1003 814
rect 1079 810 1083 814
rect 1111 810 1115 814
rect 1199 810 1203 814
rect 1231 810 1235 814
rect 1327 810 1331 814
rect 1351 810 1355 814
rect 1455 810 1459 814
rect 2007 810 2011 814
rect 471 730 475 734
rect 535 730 539 734
rect 639 730 643 734
rect 679 730 683 734
rect 807 730 811 734
rect 815 730 819 734
rect 111 654 115 658
rect 295 654 299 658
rect 311 654 315 658
rect 447 654 451 658
rect 951 730 955 734
rect 975 730 979 734
rect 1079 730 1083 734
rect 1135 730 1139 734
rect 1199 730 1203 734
rect 1295 730 1299 734
rect 1327 730 1331 734
rect 3079 818 3083 822
rect 3711 898 3715 902
rect 3727 898 3731 902
rect 3943 978 3947 982
rect 3839 898 3843 902
rect 3207 818 3211 822
rect 3239 818 3243 822
rect 3335 818 3339 822
rect 3391 818 3395 822
rect 3463 818 3467 822
rect 3543 818 3547 822
rect 3591 818 3595 822
rect 3703 818 3707 822
rect 3727 818 3731 822
rect 3839 818 3843 822
rect 2047 738 2051 742
rect 2071 738 2075 742
rect 2183 738 2187 742
rect 2335 738 2339 742
rect 2471 738 2475 742
rect 2487 738 2491 742
rect 2615 738 2619 742
rect 2639 738 2643 742
rect 1455 730 1459 734
rect 1607 730 1611 734
rect 1767 730 1771 734
rect 1903 730 1907 734
rect 2007 730 2011 734
rect 471 654 475 658
rect 111 574 115 578
rect 239 574 243 578
rect 295 574 299 578
rect 615 654 619 658
rect 639 654 643 658
rect 783 654 787 658
rect 807 654 811 658
rect 951 654 955 658
rect 975 654 979 658
rect 1203 664 1207 668
rect 1111 654 1115 658
rect 1699 664 1703 668
rect 1135 654 1139 658
rect 1263 654 1267 658
rect 1295 654 1299 658
rect 1399 654 1403 658
rect 1455 654 1459 658
rect 1535 654 1539 658
rect 1607 654 1611 658
rect 1663 654 1667 658
rect 1767 654 1771 658
rect 1791 654 1795 658
rect 1903 654 1907 658
rect 2007 654 2011 658
rect 2767 738 2771 742
rect 2807 738 2811 742
rect 2919 738 2923 742
rect 2983 738 2987 742
rect 3079 738 3083 742
rect 3167 738 3171 742
rect 3239 738 3243 742
rect 3367 738 3371 742
rect 3391 738 3395 742
rect 415 574 419 578
rect 447 574 451 578
rect 607 574 611 578
rect 615 574 619 578
rect 783 574 787 578
rect 799 574 803 578
rect 951 574 955 578
rect 991 574 995 578
rect 1111 574 1115 578
rect 1175 574 1179 578
rect 1263 574 1267 578
rect 1351 574 1355 578
rect 1399 574 1403 578
rect 1519 574 1523 578
rect 1535 574 1539 578
rect 1663 574 1667 578
rect 1687 574 1691 578
rect 1791 574 1795 578
rect 2047 650 2051 654
rect 2071 650 2075 654
rect 2183 650 2187 654
rect 2239 650 2243 654
rect 2335 650 2339 654
rect 2423 650 2427 654
rect 2487 650 2491 654
rect 2623 650 2627 654
rect 2639 650 2643 654
rect 2807 650 2811 654
rect 2839 650 2843 654
rect 2983 650 2987 654
rect 3071 650 3075 654
rect 3167 650 3171 654
rect 3543 738 3547 742
rect 3575 738 3579 742
rect 3703 738 3707 742
rect 3943 898 3947 902
rect 3943 818 3947 822
rect 3783 738 3787 742
rect 3839 738 3843 742
rect 3319 650 3323 654
rect 3367 650 3371 654
rect 3575 650 3579 654
rect 3783 650 3787 654
rect 3839 650 3843 654
rect 1863 574 1867 578
rect 1903 574 1907 578
rect 2007 574 2011 578
rect 2047 574 2051 578
rect 2071 574 2075 578
rect 2191 574 2195 578
rect 2239 574 2243 578
rect 2287 574 2291 578
rect 111 498 115 502
rect 135 498 139 502
rect 239 498 243 502
rect 287 498 291 502
rect 415 498 419 502
rect 463 498 467 502
rect 111 418 115 422
rect 135 418 139 422
rect 607 498 611 502
rect 639 498 643 502
rect 799 498 803 502
rect 807 498 811 502
rect 2383 574 2387 578
rect 2423 574 2427 578
rect 2479 574 2483 578
rect 2583 574 2587 578
rect 2623 574 2627 578
rect 967 498 971 502
rect 991 498 995 502
rect 1119 498 1123 502
rect 1175 498 1179 502
rect 1271 498 1275 502
rect 1351 498 1355 502
rect 1415 498 1419 502
rect 1519 498 1523 502
rect 1567 498 1571 502
rect 1687 498 1691 502
rect 1863 498 1867 502
rect 2007 498 2011 502
rect 2047 498 2051 502
rect 2191 498 2195 502
rect 2287 498 2291 502
rect 2383 498 2387 502
rect 2431 498 2435 502
rect 2479 498 2483 502
rect 2527 498 2531 502
rect 279 418 283 422
rect 287 418 291 422
rect 439 418 443 422
rect 463 418 467 422
rect 111 342 115 346
rect 135 342 139 346
rect 583 418 587 422
rect 639 418 643 422
rect 719 418 723 422
rect 807 418 811 422
rect 847 418 851 422
rect 967 418 971 422
rect 1087 418 1091 422
rect 1119 418 1123 422
rect 1207 418 1211 422
rect 1271 418 1275 422
rect 2711 574 2715 578
rect 2839 574 2843 578
rect 2871 574 2875 578
rect 3071 574 3075 578
rect 3303 574 3307 578
rect 3319 574 3323 578
rect 3551 574 3555 578
rect 3575 574 3579 578
rect 3807 574 3811 578
rect 3839 574 3843 578
rect 3943 738 3947 742
rect 3943 650 3947 654
rect 2583 498 2587 502
rect 2623 498 2627 502
rect 2711 498 2715 502
rect 2727 498 2731 502
rect 2847 498 2851 502
rect 2871 498 2875 502
rect 2999 498 3003 502
rect 3071 498 3075 502
rect 3175 498 3179 502
rect 3303 498 3307 502
rect 3375 498 3379 502
rect 3551 498 3555 502
rect 3591 498 3595 502
rect 3943 574 3947 578
rect 3807 498 3811 502
rect 3943 498 3947 502
rect 1327 418 1331 422
rect 1415 418 1419 422
rect 1567 418 1571 422
rect 2007 418 2011 422
rect 2047 422 2051 426
rect 2431 422 2435 426
rect 2527 422 2531 426
rect 2623 422 2627 426
rect 2719 422 2723 426
rect 2727 422 2731 426
rect 2815 422 2819 426
rect 2847 422 2851 426
rect 2927 422 2931 426
rect 143 342 147 346
rect 279 342 283 346
rect 319 342 323 346
rect 439 342 443 346
rect 479 342 483 346
rect 583 342 587 346
rect 631 342 635 346
rect 719 342 723 346
rect 775 342 779 346
rect 111 262 115 266
rect 143 262 147 266
rect 223 262 227 266
rect 319 262 323 266
rect 391 262 395 266
rect 479 262 483 266
rect 2999 422 3003 426
rect 3063 422 3067 426
rect 3175 422 3179 426
rect 3223 422 3227 426
rect 3375 422 3379 426
rect 3399 422 3403 426
rect 3591 422 3595 426
rect 3783 422 3787 426
rect 3807 422 3811 426
rect 847 342 851 346
rect 903 342 907 346
rect 967 342 971 346
rect 1031 342 1035 346
rect 1087 342 1091 346
rect 1151 342 1155 346
rect 1207 342 1211 346
rect 1271 342 1275 346
rect 1327 342 1331 346
rect 1391 342 1395 346
rect 2007 342 2011 346
rect 2047 342 2051 346
rect 2191 342 2195 346
rect 2327 342 2331 346
rect 2431 342 2435 346
rect 2471 342 2475 346
rect 2527 342 2531 346
rect 2623 342 2627 346
rect 2719 342 2723 346
rect 2783 342 2787 346
rect 2815 342 2819 346
rect 2927 342 2931 346
rect 2951 342 2955 346
rect 3063 342 3067 346
rect 3119 342 3123 346
rect 3223 342 3227 346
rect 3295 342 3299 346
rect 3399 342 3403 346
rect 3471 342 3475 346
rect 3591 342 3595 346
rect 3655 342 3659 346
rect 559 262 563 266
rect 631 262 635 266
rect 111 154 115 158
rect 151 154 155 158
rect 223 154 227 158
rect 735 262 739 266
rect 775 262 779 266
rect 903 262 907 266
rect 1031 262 1035 266
rect 1063 262 1067 266
rect 1151 262 1155 266
rect 1215 262 1219 266
rect 1271 262 1275 266
rect 1359 262 1363 266
rect 1391 262 1395 266
rect 1511 262 1515 266
rect 3783 342 3787 346
rect 3839 342 3843 346
rect 1663 262 1667 266
rect 2007 262 2011 266
rect 2047 266 2051 270
rect 2071 266 2075 270
rect 2191 266 2195 270
rect 2215 266 2219 270
rect 2327 266 2331 270
rect 2399 266 2403 270
rect 247 154 251 158
rect 343 154 347 158
rect 391 154 395 158
rect 439 154 443 158
rect 535 154 539 158
rect 559 154 563 158
rect 631 154 635 158
rect 727 154 731 158
rect 735 154 739 158
rect 823 154 827 158
rect 903 154 907 158
rect 919 154 923 158
rect 1015 154 1019 158
rect 1063 154 1067 158
rect 2047 166 2051 170
rect 2071 166 2075 170
rect 2191 166 2195 170
rect 2215 166 2219 170
rect 1111 154 1115 158
rect 1207 154 1211 158
rect 1215 154 1219 158
rect 1303 154 1307 158
rect 1359 154 1363 158
rect 1407 154 1411 158
rect 1511 154 1515 158
rect 1615 154 1619 158
rect 1663 154 1667 158
rect 1711 154 1715 158
rect 1807 154 1811 158
rect 1903 154 1907 158
rect 2007 154 2011 158
rect 2471 266 2475 270
rect 2591 266 2595 270
rect 2623 266 2627 270
rect 2783 266 2787 270
rect 2791 266 2795 270
rect 2951 266 2955 270
rect 2983 266 2987 270
rect 3119 266 3123 270
rect 3167 266 3171 270
rect 3295 266 3299 270
rect 3343 266 3347 270
rect 2343 166 2347 170
rect 2399 166 2403 170
rect 2495 166 2499 170
rect 2591 166 2595 170
rect 2647 166 2651 170
rect 2791 166 2795 170
rect 2799 166 2803 170
rect 3471 266 3475 270
rect 3511 266 3515 270
rect 3655 266 3659 270
rect 3687 266 3691 270
rect 3943 422 3947 426
rect 3943 342 3947 346
rect 3839 266 3843 270
rect 2943 166 2947 170
rect 2983 166 2987 170
rect 3071 166 3075 170
rect 3167 166 3171 170
rect 3191 166 3195 170
rect 3311 166 3315 170
rect 3343 166 3347 170
rect 3423 166 3427 170
rect 3511 166 3515 170
rect 3527 166 3531 170
rect 3639 166 3643 170
rect 3687 166 3691 170
rect 3743 166 3747 170
rect 3839 166 3843 170
rect 3943 266 3947 270
rect 3943 166 3947 170
rect 2047 90 2051 94
rect 2071 90 2075 94
rect 2191 90 2195 94
rect 2343 90 2347 94
rect 2495 90 2499 94
rect 2647 90 2651 94
rect 2799 90 2803 94
rect 2943 90 2947 94
rect 3071 90 3075 94
rect 3191 90 3195 94
rect 3311 90 3315 94
rect 3423 90 3427 94
rect 3527 90 3531 94
rect 3639 90 3643 94
rect 3743 90 3747 94
rect 3839 90 3843 94
rect 3943 90 3947 94
rect 111 78 115 82
rect 151 78 155 82
rect 247 78 251 82
rect 343 78 347 82
rect 439 78 443 82
rect 535 78 539 82
rect 631 78 635 82
rect 727 78 731 82
rect 823 78 827 82
rect 919 78 923 82
rect 1015 78 1019 82
rect 1111 78 1115 82
rect 1207 78 1211 82
rect 1303 78 1307 82
rect 1407 78 1411 82
rect 1511 78 1515 82
rect 1615 78 1619 82
rect 1711 78 1715 82
rect 1807 78 1811 82
rect 1903 78 1907 82
rect 2007 78 2011 82
<< m4 >>
rect 2018 4017 2019 4023
rect 2025 4022 3967 4023
rect 2025 4018 2047 4022
rect 2051 4018 2071 4022
rect 2075 4018 2327 4022
rect 2331 4018 2591 4022
rect 2595 4018 2839 4022
rect 2843 4018 3087 4022
rect 3091 4018 3343 4022
rect 3347 4018 3943 4022
rect 3947 4018 3967 4022
rect 2025 4017 3967 4018
rect 3973 4017 3974 4023
rect 84 3997 85 4003
rect 91 4002 2019 4003
rect 91 3998 111 4002
rect 115 3998 311 4002
rect 315 3998 511 4002
rect 515 3998 703 4002
rect 707 3998 887 4002
rect 891 3998 1063 4002
rect 1067 3998 1231 4002
rect 1235 3998 1383 4002
rect 1387 3998 1519 4002
rect 1523 3998 1655 4002
rect 1659 3998 1791 4002
rect 1795 3998 1903 4002
rect 1907 3998 2007 4002
rect 2011 3998 2019 4002
rect 91 3997 2019 3998
rect 2025 3997 2026 4003
rect 2030 3941 2031 3947
rect 2037 3946 3979 3947
rect 2037 3942 2047 3946
rect 2051 3942 2071 3946
rect 2075 3942 2127 3946
rect 2131 3942 2271 3946
rect 2275 3942 2327 3946
rect 2331 3942 2439 3946
rect 2443 3942 2591 3946
rect 2595 3942 2615 3946
rect 2619 3942 2799 3946
rect 2803 3942 2839 3946
rect 2843 3942 2983 3946
rect 2987 3942 3087 3946
rect 3091 3942 3175 3946
rect 3179 3942 3343 3946
rect 3347 3942 3367 3946
rect 3371 3942 3559 3946
rect 3563 3942 3943 3946
rect 3947 3942 3979 3946
rect 2037 3941 3979 3942
rect 3985 3941 3986 3947
rect 96 3921 97 3927
rect 103 3926 2031 3927
rect 103 3922 111 3926
rect 115 3922 279 3926
rect 283 3922 311 3926
rect 315 3922 415 3926
rect 419 3922 511 3926
rect 515 3922 567 3926
rect 571 3922 703 3926
rect 707 3922 735 3926
rect 739 3922 887 3926
rect 891 3922 911 3926
rect 915 3922 1063 3926
rect 1067 3922 1095 3926
rect 1099 3922 1231 3926
rect 1235 3922 1287 3926
rect 1291 3922 1383 3926
rect 1387 3922 1479 3926
rect 1483 3922 1519 3926
rect 1523 3922 1655 3926
rect 1659 3922 1679 3926
rect 1683 3922 1791 3926
rect 1795 3922 1903 3926
rect 1907 3922 2007 3926
rect 2011 3922 2031 3926
rect 103 3921 2031 3922
rect 2037 3921 2038 3927
rect 2018 3865 2019 3871
rect 2025 3870 3967 3871
rect 2025 3866 2047 3870
rect 2051 3866 2127 3870
rect 2131 3866 2263 3870
rect 2267 3866 2271 3870
rect 2275 3866 2375 3870
rect 2379 3866 2439 3870
rect 2443 3866 2495 3870
rect 2499 3866 2615 3870
rect 2619 3866 2631 3870
rect 2635 3866 2775 3870
rect 2779 3866 2799 3870
rect 2803 3866 2919 3870
rect 2923 3866 2983 3870
rect 2987 3866 3063 3870
rect 3067 3866 3175 3870
rect 3179 3866 3207 3870
rect 3211 3866 3343 3870
rect 3347 3866 3367 3870
rect 3371 3866 3471 3870
rect 3475 3866 3559 3870
rect 3563 3866 3599 3870
rect 3603 3866 3727 3870
rect 3731 3866 3839 3870
rect 3843 3866 3943 3870
rect 3947 3866 3967 3870
rect 2025 3865 3967 3866
rect 3973 3865 3974 3871
rect 84 3837 85 3843
rect 91 3842 2019 3843
rect 91 3838 111 3842
rect 115 3838 231 3842
rect 235 3838 279 3842
rect 283 3838 335 3842
rect 339 3838 415 3842
rect 419 3838 439 3842
rect 443 3838 535 3842
rect 539 3838 567 3842
rect 571 3838 631 3842
rect 635 3838 727 3842
rect 731 3838 735 3842
rect 739 3838 831 3842
rect 835 3838 911 3842
rect 915 3838 935 3842
rect 939 3838 1039 3842
rect 1043 3838 1095 3842
rect 1099 3838 1151 3842
rect 1155 3838 1263 3842
rect 1267 3838 1287 3842
rect 1291 3838 1383 3842
rect 1387 3838 1479 3842
rect 1483 3838 1503 3842
rect 1507 3838 1631 3842
rect 1635 3838 1679 3842
rect 1683 3838 2007 3842
rect 2011 3838 2019 3842
rect 91 3837 2019 3838
rect 2025 3837 2026 3843
rect 2030 3773 2031 3779
rect 2037 3778 3979 3779
rect 2037 3774 2047 3778
rect 2051 3774 2071 3778
rect 2075 3774 2183 3778
rect 2187 3774 2263 3778
rect 2267 3774 2327 3778
rect 2331 3774 2375 3778
rect 2379 3774 2479 3778
rect 2483 3774 2495 3778
rect 2499 3774 2631 3778
rect 2635 3774 2639 3778
rect 2643 3774 2775 3778
rect 2779 3774 2807 3778
rect 2811 3774 2919 3778
rect 2923 3774 2983 3778
rect 2987 3774 3063 3778
rect 3067 3774 3159 3778
rect 3163 3774 3207 3778
rect 3211 3774 3335 3778
rect 3339 3774 3343 3778
rect 3347 3774 3471 3778
rect 3475 3774 3511 3778
rect 3515 3774 3599 3778
rect 3603 3774 3687 3778
rect 3691 3774 3727 3778
rect 3731 3774 3839 3778
rect 3843 3774 3943 3778
rect 3947 3774 3979 3778
rect 2037 3773 3979 3774
rect 3985 3773 3986 3779
rect 96 3761 97 3767
rect 103 3766 2031 3767
rect 103 3762 111 3766
rect 115 3762 159 3766
rect 163 3762 231 3766
rect 235 3762 335 3766
rect 339 3762 351 3766
rect 355 3762 439 3766
rect 443 3762 535 3766
rect 539 3762 551 3766
rect 555 3762 631 3766
rect 635 3762 727 3766
rect 731 3762 751 3766
rect 755 3762 831 3766
rect 835 3762 935 3766
rect 939 3762 959 3766
rect 963 3762 1039 3766
rect 1043 3762 1151 3766
rect 1155 3762 1167 3766
rect 1171 3762 1263 3766
rect 1267 3762 1383 3766
rect 1387 3762 1503 3766
rect 1507 3762 1607 3766
rect 1611 3762 1631 3766
rect 1635 3762 2007 3766
rect 2011 3762 2031 3766
rect 103 3761 2031 3762
rect 2037 3761 2038 3767
rect 2018 3685 2019 3691
rect 2025 3690 3967 3691
rect 2025 3686 2047 3690
rect 2051 3686 2071 3690
rect 2075 3686 2183 3690
rect 2187 3686 2199 3690
rect 2203 3686 2327 3690
rect 2331 3686 2367 3690
rect 2371 3686 2479 3690
rect 2483 3686 2551 3690
rect 2555 3686 2639 3690
rect 2643 3686 2735 3690
rect 2739 3686 2807 3690
rect 2811 3686 2927 3690
rect 2931 3686 2983 3690
rect 2987 3686 3111 3690
rect 3115 3686 3159 3690
rect 3163 3686 3295 3690
rect 3299 3686 3335 3690
rect 3339 3686 3479 3690
rect 3483 3686 3511 3690
rect 3515 3686 3671 3690
rect 3675 3686 3687 3690
rect 3691 3686 3839 3690
rect 3843 3686 3943 3690
rect 3947 3686 3967 3690
rect 2025 3685 3967 3686
rect 3973 3685 3974 3691
rect 2018 3683 2026 3685
rect 84 3677 85 3683
rect 91 3682 2019 3683
rect 91 3678 111 3682
rect 115 3678 151 3682
rect 155 3678 159 3682
rect 163 3678 351 3682
rect 355 3678 383 3682
rect 387 3678 551 3682
rect 555 3678 615 3682
rect 619 3678 751 3682
rect 755 3678 839 3682
rect 843 3678 959 3682
rect 963 3678 1055 3682
rect 1059 3678 1167 3682
rect 1171 3678 1263 3682
rect 1267 3678 1383 3682
rect 1387 3678 1479 3682
rect 1483 3678 1607 3682
rect 1611 3678 1695 3682
rect 1699 3678 2007 3682
rect 2011 3678 2019 3682
rect 91 3677 2019 3678
rect 2025 3677 2026 3683
rect 2030 3605 2031 3611
rect 2037 3610 3979 3611
rect 2037 3606 2047 3610
rect 2051 3606 2071 3610
rect 2075 3606 2103 3610
rect 2107 3606 2199 3610
rect 2203 3606 2279 3610
rect 2283 3606 2367 3610
rect 2371 3606 2471 3610
rect 2475 3606 2551 3610
rect 2555 3606 2671 3610
rect 2675 3606 2735 3610
rect 2739 3606 2871 3610
rect 2875 3606 2927 3610
rect 2931 3606 3063 3610
rect 3067 3606 3111 3610
rect 3115 3606 3255 3610
rect 3259 3606 3295 3610
rect 3299 3606 3447 3610
rect 3451 3606 3479 3610
rect 3483 3606 3639 3610
rect 3643 3606 3671 3610
rect 3675 3606 3839 3610
rect 3843 3606 3943 3610
rect 3947 3606 3979 3610
rect 2037 3605 3979 3606
rect 3985 3605 3986 3611
rect 2030 3603 2038 3605
rect 96 3597 97 3603
rect 103 3602 2031 3603
rect 103 3598 111 3602
rect 115 3598 151 3602
rect 155 3598 167 3602
rect 171 3598 359 3602
rect 363 3598 383 3602
rect 387 3598 559 3602
rect 563 3598 615 3602
rect 619 3598 775 3602
rect 779 3598 839 3602
rect 843 3598 991 3602
rect 995 3598 1055 3602
rect 1059 3598 1215 3602
rect 1219 3598 1263 3602
rect 1267 3598 1447 3602
rect 1451 3598 1479 3602
rect 1483 3598 1687 3602
rect 1691 3598 1695 3602
rect 1699 3598 2007 3602
rect 2011 3598 2031 3602
rect 103 3597 2031 3598
rect 2037 3597 2038 3603
rect 2018 3525 2019 3531
rect 2025 3530 3967 3531
rect 2025 3526 2047 3530
rect 2051 3526 2103 3530
rect 2107 3526 2279 3530
rect 2283 3526 2327 3530
rect 2331 3526 2447 3530
rect 2451 3526 2471 3530
rect 2475 3526 2583 3530
rect 2587 3526 2671 3530
rect 2675 3526 2735 3530
rect 2739 3526 2871 3530
rect 2875 3526 2911 3530
rect 2915 3526 3063 3530
rect 3067 3526 3111 3530
rect 3115 3526 3255 3530
rect 3259 3526 3335 3530
rect 3339 3526 3447 3530
rect 3451 3526 3567 3530
rect 3571 3526 3639 3530
rect 3643 3526 3807 3530
rect 3811 3526 3839 3530
rect 3843 3526 3943 3530
rect 3947 3526 3967 3530
rect 2025 3525 3967 3526
rect 3973 3525 3974 3531
rect 84 3513 85 3519
rect 91 3518 2019 3519
rect 91 3514 111 3518
rect 115 3514 167 3518
rect 171 3514 295 3518
rect 299 3514 359 3518
rect 363 3514 431 3518
rect 435 3514 559 3518
rect 563 3514 583 3518
rect 587 3514 743 3518
rect 747 3514 775 3518
rect 779 3514 911 3518
rect 915 3514 991 3518
rect 995 3514 1079 3518
rect 1083 3514 1215 3518
rect 1219 3514 1247 3518
rect 1251 3514 1423 3518
rect 1427 3514 1447 3518
rect 1451 3514 1599 3518
rect 1603 3514 1687 3518
rect 1691 3514 1775 3518
rect 1779 3514 2007 3518
rect 2011 3514 2019 3518
rect 91 3513 2019 3514
rect 2025 3513 2026 3519
rect 2030 3449 2031 3455
rect 2037 3454 3979 3455
rect 2037 3450 2047 3454
rect 2051 3450 2327 3454
rect 2331 3450 2447 3454
rect 2451 3450 2551 3454
rect 2555 3450 2583 3454
rect 2587 3450 2663 3454
rect 2667 3450 2735 3454
rect 2739 3450 2775 3454
rect 2779 3450 2903 3454
rect 2907 3450 2911 3454
rect 2915 3450 3047 3454
rect 3051 3450 3111 3454
rect 3115 3450 3207 3454
rect 3211 3450 3335 3454
rect 3339 3450 3383 3454
rect 3387 3450 3567 3454
rect 3571 3450 3751 3454
rect 3755 3450 3807 3454
rect 3811 3450 3943 3454
rect 3947 3450 3979 3454
rect 2037 3449 3979 3450
rect 3985 3449 3986 3455
rect 96 3417 97 3423
rect 103 3422 2031 3423
rect 103 3418 111 3422
rect 115 3418 295 3422
rect 299 3418 431 3422
rect 435 3418 495 3422
rect 499 3418 583 3422
rect 587 3418 647 3422
rect 651 3418 743 3422
rect 747 3418 799 3422
rect 803 3418 911 3422
rect 915 3418 959 3422
rect 963 3418 1079 3422
rect 1083 3418 1127 3422
rect 1131 3418 1247 3422
rect 1251 3418 1295 3422
rect 1299 3418 1423 3422
rect 1427 3418 1463 3422
rect 1467 3418 1599 3422
rect 1603 3418 1639 3422
rect 1643 3418 1775 3422
rect 1779 3418 1815 3422
rect 1819 3418 2007 3422
rect 2011 3418 2031 3422
rect 103 3417 2031 3418
rect 2037 3417 2038 3423
rect 2018 3361 2019 3367
rect 2025 3366 3967 3367
rect 2025 3362 2047 3366
rect 2051 3362 2447 3366
rect 2451 3362 2551 3366
rect 2555 3362 2567 3366
rect 2571 3362 2663 3366
rect 2667 3362 2719 3366
rect 2723 3362 2775 3366
rect 2779 3362 2871 3366
rect 2875 3362 2903 3366
rect 2907 3362 3023 3366
rect 3027 3362 3047 3366
rect 3051 3362 3175 3366
rect 3179 3362 3207 3366
rect 3211 3362 3327 3366
rect 3331 3362 3383 3366
rect 3387 3362 3479 3366
rect 3483 3362 3567 3366
rect 3571 3362 3631 3366
rect 3635 3362 3751 3366
rect 3755 3362 3783 3366
rect 3787 3362 3943 3366
rect 3947 3362 3967 3366
rect 2025 3361 3967 3362
rect 3973 3361 3974 3367
rect 84 3329 85 3335
rect 91 3334 2019 3335
rect 91 3330 111 3334
rect 115 3330 135 3334
rect 139 3330 295 3334
rect 299 3330 479 3334
rect 483 3330 495 3334
rect 499 3330 647 3334
rect 651 3330 671 3334
rect 675 3330 799 3334
rect 803 3330 863 3334
rect 867 3330 959 3334
rect 963 3330 1055 3334
rect 1059 3330 1127 3334
rect 1131 3330 1247 3334
rect 1251 3330 1295 3334
rect 1299 3330 1439 3334
rect 1443 3330 1463 3334
rect 1467 3330 1631 3334
rect 1635 3330 1639 3334
rect 1643 3330 1815 3334
rect 1819 3330 1823 3334
rect 1827 3330 2007 3334
rect 2011 3330 2019 3334
rect 91 3329 2019 3330
rect 2025 3329 2026 3335
rect 2030 3281 2031 3287
rect 2037 3286 3979 3287
rect 2037 3282 2047 3286
rect 2051 3282 2415 3286
rect 2419 3282 2551 3286
rect 2555 3282 2567 3286
rect 2571 3282 2687 3286
rect 2691 3282 2719 3286
rect 2723 3282 2831 3286
rect 2835 3282 2871 3286
rect 2875 3282 2975 3286
rect 2979 3282 3023 3286
rect 3027 3282 3119 3286
rect 3123 3282 3175 3286
rect 3179 3282 3255 3286
rect 3259 3282 3327 3286
rect 3331 3282 3383 3286
rect 3387 3282 3479 3286
rect 3483 3282 3503 3286
rect 3507 3282 3623 3286
rect 3627 3282 3631 3286
rect 3635 3282 3743 3286
rect 3747 3282 3783 3286
rect 3787 3282 3839 3286
rect 3843 3282 3943 3286
rect 3947 3282 3979 3286
rect 2037 3281 3979 3282
rect 3985 3281 3986 3287
rect 96 3249 97 3255
rect 103 3254 2031 3255
rect 103 3250 111 3254
rect 115 3250 135 3254
rect 139 3250 295 3254
rect 299 3250 319 3254
rect 323 3250 479 3254
rect 483 3250 519 3254
rect 523 3250 671 3254
rect 675 3250 719 3254
rect 723 3250 863 3254
rect 867 3250 911 3254
rect 915 3250 1055 3254
rect 1059 3250 1095 3254
rect 1099 3250 1247 3254
rect 1251 3250 1271 3254
rect 1275 3250 1439 3254
rect 1443 3250 1447 3254
rect 1451 3250 1623 3254
rect 1627 3250 1631 3254
rect 1635 3250 1799 3254
rect 1803 3250 1823 3254
rect 1827 3250 2007 3254
rect 2011 3250 2031 3254
rect 103 3249 2031 3250
rect 2037 3249 2038 3255
rect 2018 3193 2019 3199
rect 2025 3198 3967 3199
rect 2025 3194 2047 3198
rect 2051 3194 2247 3198
rect 2251 3194 2399 3198
rect 2403 3194 2415 3198
rect 2419 3194 2551 3198
rect 2555 3194 2559 3198
rect 2563 3194 2687 3198
rect 2691 3194 2727 3198
rect 2731 3194 2831 3198
rect 2835 3194 2903 3198
rect 2907 3194 2975 3198
rect 2979 3194 3079 3198
rect 3083 3194 3119 3198
rect 3123 3194 3255 3198
rect 3259 3194 3263 3198
rect 3267 3194 3383 3198
rect 3387 3194 3447 3198
rect 3451 3194 3503 3198
rect 3507 3194 3623 3198
rect 3627 3194 3631 3198
rect 3635 3194 3743 3198
rect 3747 3194 3815 3198
rect 3819 3194 3839 3198
rect 3843 3194 3943 3198
rect 3947 3194 3967 3198
rect 2025 3193 3967 3194
rect 3973 3193 3974 3199
rect 84 3165 85 3171
rect 91 3170 2019 3171
rect 91 3166 111 3170
rect 115 3166 135 3170
rect 139 3166 143 3170
rect 147 3166 319 3170
rect 323 3166 343 3170
rect 347 3166 519 3170
rect 523 3166 543 3170
rect 547 3166 719 3170
rect 723 3166 743 3170
rect 747 3166 911 3170
rect 915 3166 927 3170
rect 931 3166 1095 3170
rect 1099 3166 1103 3170
rect 1107 3166 1263 3170
rect 1267 3166 1271 3170
rect 1275 3166 1423 3170
rect 1427 3166 1447 3170
rect 1451 3166 1575 3170
rect 1579 3166 1623 3170
rect 1627 3166 1735 3170
rect 1739 3166 1799 3170
rect 1803 3166 2007 3170
rect 2011 3166 2019 3170
rect 91 3165 2019 3166
rect 2025 3165 2026 3171
rect 2030 3113 2031 3119
rect 2037 3118 3979 3119
rect 2037 3114 2047 3118
rect 2051 3114 2079 3118
rect 2083 3114 2223 3118
rect 2227 3114 2247 3118
rect 2251 3114 2375 3118
rect 2379 3114 2399 3118
rect 2403 3114 2527 3118
rect 2531 3114 2559 3118
rect 2563 3114 2687 3118
rect 2691 3114 2727 3118
rect 2731 3114 2855 3118
rect 2859 3114 2903 3118
rect 2907 3114 3039 3118
rect 3043 3114 3079 3118
rect 3083 3114 3231 3118
rect 3235 3114 3263 3118
rect 3267 3114 3431 3118
rect 3435 3114 3447 3118
rect 3451 3114 3631 3118
rect 3635 3114 3639 3118
rect 3643 3114 3815 3118
rect 3819 3114 3839 3118
rect 3843 3114 3943 3118
rect 3947 3114 3979 3118
rect 2037 3113 3979 3114
rect 3985 3113 3986 3119
rect 96 3089 97 3095
rect 103 3094 2031 3095
rect 103 3090 111 3094
rect 115 3090 143 3094
rect 147 3090 263 3094
rect 267 3090 343 3094
rect 347 3090 439 3094
rect 443 3090 543 3094
rect 547 3090 615 3094
rect 619 3090 743 3094
rect 747 3090 799 3094
rect 803 3090 927 3094
rect 931 3090 975 3094
rect 979 3090 1103 3094
rect 1107 3090 1143 3094
rect 1147 3090 1263 3094
rect 1267 3090 1303 3094
rect 1307 3090 1423 3094
rect 1427 3090 1455 3094
rect 1459 3090 1575 3094
rect 1579 3090 1607 3094
rect 1611 3090 1735 3094
rect 1739 3090 1767 3094
rect 1771 3090 2007 3094
rect 2011 3090 2031 3094
rect 103 3089 2031 3090
rect 2037 3089 2038 3095
rect 2018 3029 2019 3035
rect 2025 3034 3967 3035
rect 2025 3030 2047 3034
rect 2051 3030 2071 3034
rect 2075 3030 2079 3034
rect 2083 3030 2183 3034
rect 2187 3030 2223 3034
rect 2227 3030 2327 3034
rect 2331 3030 2375 3034
rect 2379 3030 2479 3034
rect 2483 3030 2527 3034
rect 2531 3030 2655 3034
rect 2659 3030 2687 3034
rect 2691 3030 2855 3034
rect 2859 3030 3039 3034
rect 3043 3030 3087 3034
rect 3091 3030 3231 3034
rect 3235 3030 3335 3034
rect 3339 3030 3431 3034
rect 3435 3030 3599 3034
rect 3603 3030 3639 3034
rect 3643 3030 3839 3034
rect 3843 3030 3943 3034
rect 3947 3030 3967 3034
rect 2025 3029 3967 3030
rect 3973 3029 3974 3035
rect 84 2989 85 2995
rect 91 2994 2019 2995
rect 91 2990 111 2994
rect 115 2990 263 2994
rect 267 2990 343 2994
rect 347 2990 439 2994
rect 443 2990 543 2994
rect 547 2990 615 2994
rect 619 2990 655 2994
rect 659 2990 783 2994
rect 787 2990 799 2994
rect 803 2990 935 2994
rect 939 2990 975 2994
rect 979 2990 1103 2994
rect 1107 2990 1143 2994
rect 1147 2990 1295 2994
rect 1299 2990 1303 2994
rect 1307 2990 1455 2994
rect 1459 2990 1495 2994
rect 1499 2990 1607 2994
rect 1611 2990 1711 2994
rect 1715 2990 1767 2994
rect 1771 2990 1903 2994
rect 1907 2990 2007 2994
rect 2011 2990 2019 2994
rect 91 2989 2019 2990
rect 2025 2989 2026 2995
rect 2030 2949 2031 2955
rect 2037 2954 3979 2955
rect 2037 2950 2047 2954
rect 2051 2950 2071 2954
rect 2075 2950 2183 2954
rect 2187 2950 2263 2954
rect 2267 2950 2327 2954
rect 2331 2950 2479 2954
rect 2483 2950 2487 2954
rect 2491 2950 2655 2954
rect 2659 2950 2735 2954
rect 2739 2950 2855 2954
rect 2859 2950 2999 2954
rect 3003 2950 3087 2954
rect 3091 2950 3279 2954
rect 3283 2950 3335 2954
rect 3339 2950 3567 2954
rect 3571 2950 3599 2954
rect 3603 2950 3839 2954
rect 3843 2950 3943 2954
rect 3947 2950 3979 2954
rect 2037 2949 3979 2950
rect 3985 2949 3986 2955
rect 96 2913 97 2919
rect 103 2918 2031 2919
rect 103 2914 111 2918
rect 115 2914 207 2918
rect 211 2914 327 2918
rect 331 2914 343 2918
rect 347 2914 439 2918
rect 443 2914 447 2918
rect 451 2914 543 2918
rect 547 2914 575 2918
rect 579 2914 655 2918
rect 659 2914 703 2918
rect 707 2914 783 2918
rect 787 2914 847 2918
rect 851 2914 935 2918
rect 939 2914 999 2918
rect 1003 2914 1103 2918
rect 1107 2914 1167 2918
rect 1171 2914 1295 2918
rect 1299 2914 1351 2918
rect 1355 2914 1495 2918
rect 1499 2914 1535 2918
rect 1539 2914 1711 2918
rect 1715 2914 1727 2918
rect 1731 2914 1903 2918
rect 1907 2914 2007 2918
rect 2011 2914 2031 2918
rect 103 2913 2031 2914
rect 2037 2913 2038 2919
rect 2018 2865 2019 2871
rect 2025 2870 3967 2871
rect 2025 2866 2047 2870
rect 2051 2866 2071 2870
rect 2075 2866 2263 2870
rect 2267 2866 2487 2870
rect 2491 2866 2671 2870
rect 2675 2866 2735 2870
rect 2739 2866 2887 2870
rect 2891 2866 2999 2870
rect 3003 2866 3095 2870
rect 3099 2866 3279 2870
rect 3283 2866 3287 2870
rect 3291 2866 3479 2870
rect 3483 2866 3567 2870
rect 3571 2866 3671 2870
rect 3675 2866 3839 2870
rect 3843 2866 3943 2870
rect 3947 2866 3967 2870
rect 2025 2865 3967 2866
rect 3973 2865 3974 2871
rect 84 2833 85 2839
rect 91 2838 2019 2839
rect 91 2834 111 2838
rect 115 2834 135 2838
rect 139 2834 207 2838
rect 211 2834 247 2838
rect 251 2834 327 2838
rect 331 2834 399 2838
rect 403 2834 447 2838
rect 451 2834 551 2838
rect 555 2834 575 2838
rect 579 2834 703 2838
rect 707 2834 711 2838
rect 715 2834 847 2838
rect 851 2834 879 2838
rect 883 2834 999 2838
rect 1003 2834 1047 2838
rect 1051 2834 1167 2838
rect 1171 2834 1223 2838
rect 1227 2834 1351 2838
rect 1355 2834 1399 2838
rect 1403 2834 1535 2838
rect 1539 2834 1575 2838
rect 1579 2834 1727 2838
rect 1731 2834 1751 2838
rect 1755 2834 1903 2838
rect 1907 2834 2007 2838
rect 2011 2834 2019 2838
rect 91 2833 2019 2834
rect 2025 2833 2026 2839
rect 2030 2789 2031 2795
rect 2037 2794 3979 2795
rect 2037 2790 2047 2794
rect 2051 2790 2071 2794
rect 2075 2790 2199 2794
rect 2203 2790 2343 2794
rect 2347 2790 2479 2794
rect 2483 2790 2607 2794
rect 2611 2790 2671 2794
rect 2675 2790 2727 2794
rect 2731 2790 2839 2794
rect 2843 2790 2887 2794
rect 2891 2790 2943 2794
rect 2947 2790 3047 2794
rect 3051 2790 3095 2794
rect 3099 2790 3143 2794
rect 3147 2790 3239 2794
rect 3243 2790 3287 2794
rect 3291 2790 3343 2794
rect 3347 2790 3447 2794
rect 3451 2790 3479 2794
rect 3483 2790 3551 2794
rect 3555 2790 3647 2794
rect 3651 2790 3671 2794
rect 3675 2790 3743 2794
rect 3747 2790 3839 2794
rect 3843 2790 3943 2794
rect 3947 2790 3979 2794
rect 2037 2789 3979 2790
rect 3985 2789 3986 2795
rect 96 2749 97 2755
rect 103 2754 2031 2755
rect 103 2750 111 2754
rect 115 2750 135 2754
rect 139 2750 247 2754
rect 251 2750 255 2754
rect 259 2750 399 2754
rect 403 2750 407 2754
rect 411 2750 551 2754
rect 555 2750 575 2754
rect 579 2750 711 2754
rect 715 2750 743 2754
rect 747 2750 879 2754
rect 883 2750 919 2754
rect 923 2750 1047 2754
rect 1051 2750 1087 2754
rect 1091 2750 1223 2754
rect 1227 2750 1255 2754
rect 1259 2750 1399 2754
rect 1403 2750 1423 2754
rect 1427 2750 1575 2754
rect 1579 2750 1599 2754
rect 1603 2750 1751 2754
rect 1755 2750 1903 2754
rect 1907 2750 2007 2754
rect 2011 2750 2031 2754
rect 103 2749 2031 2750
rect 2037 2749 2038 2755
rect 2018 2693 2019 2699
rect 2025 2698 3967 2699
rect 2025 2694 2047 2698
rect 2051 2694 2071 2698
rect 2075 2694 2095 2698
rect 2099 2694 2199 2698
rect 2203 2694 2263 2698
rect 2267 2694 2343 2698
rect 2347 2694 2439 2698
rect 2443 2694 2479 2698
rect 2483 2694 2607 2698
rect 2611 2694 2615 2698
rect 2619 2694 2727 2698
rect 2731 2694 2783 2698
rect 2787 2694 2839 2698
rect 2843 2694 2943 2698
rect 2947 2694 3047 2698
rect 3051 2694 3095 2698
rect 3099 2694 3143 2698
rect 3147 2694 3239 2698
rect 3243 2694 3343 2698
rect 3347 2694 3383 2698
rect 3387 2694 3447 2698
rect 3451 2694 3535 2698
rect 3539 2694 3551 2698
rect 3555 2694 3647 2698
rect 3651 2694 3743 2698
rect 3747 2694 3839 2698
rect 3843 2694 3943 2698
rect 3947 2694 3967 2698
rect 2025 2693 3967 2694
rect 3973 2693 3974 2699
rect 84 2673 85 2679
rect 91 2678 2019 2679
rect 91 2674 111 2678
rect 115 2674 135 2678
rect 139 2674 167 2678
rect 171 2674 255 2678
rect 259 2674 359 2678
rect 363 2674 407 2678
rect 411 2674 559 2678
rect 563 2674 575 2678
rect 579 2674 743 2678
rect 747 2674 759 2678
rect 763 2674 919 2678
rect 923 2674 951 2678
rect 955 2674 1087 2678
rect 1091 2674 1143 2678
rect 1147 2674 1255 2678
rect 1259 2674 1327 2678
rect 1331 2674 1423 2678
rect 1427 2674 1511 2678
rect 1515 2674 1599 2678
rect 1603 2674 1703 2678
rect 1707 2674 2007 2678
rect 2011 2674 2019 2678
rect 91 2673 2019 2674
rect 2025 2673 2026 2679
rect 2030 2609 2031 2615
rect 2037 2614 3979 2615
rect 2037 2610 2047 2614
rect 2051 2610 2095 2614
rect 2099 2610 2215 2614
rect 2219 2610 2263 2614
rect 2267 2610 2367 2614
rect 2371 2610 2439 2614
rect 2443 2610 2519 2614
rect 2523 2610 2615 2614
rect 2619 2610 2671 2614
rect 2675 2610 2783 2614
rect 2787 2610 2815 2614
rect 2819 2610 2943 2614
rect 2947 2610 2951 2614
rect 2955 2610 3087 2614
rect 3091 2610 3095 2614
rect 3099 2610 3223 2614
rect 3227 2610 3239 2614
rect 3243 2610 3367 2614
rect 3371 2610 3383 2614
rect 3387 2610 3535 2614
rect 3539 2610 3943 2614
rect 3947 2610 3979 2614
rect 2037 2609 3979 2610
rect 3985 2609 3986 2615
rect 96 2581 97 2587
rect 103 2586 2031 2587
rect 103 2582 111 2586
rect 115 2582 167 2586
rect 171 2582 359 2586
rect 363 2582 559 2586
rect 563 2582 575 2586
rect 579 2582 687 2586
rect 691 2582 759 2586
rect 763 2582 807 2586
rect 811 2582 935 2586
rect 939 2582 951 2586
rect 955 2582 1071 2586
rect 1075 2582 1143 2586
rect 1147 2582 1207 2586
rect 1211 2582 1327 2586
rect 1331 2582 1351 2586
rect 1355 2582 1495 2586
rect 1499 2582 1511 2586
rect 1515 2582 1647 2586
rect 1651 2582 1703 2586
rect 1707 2582 1799 2586
rect 1803 2582 2007 2586
rect 2011 2582 2031 2586
rect 103 2581 2031 2582
rect 2037 2581 2038 2587
rect 2018 2529 2019 2535
rect 2025 2534 3967 2535
rect 2025 2530 2047 2534
rect 2051 2530 2095 2534
rect 2099 2530 2215 2534
rect 2219 2530 2343 2534
rect 2347 2530 2367 2534
rect 2371 2530 2471 2534
rect 2475 2530 2519 2534
rect 2523 2530 2599 2534
rect 2603 2530 2671 2534
rect 2675 2530 2719 2534
rect 2723 2530 2815 2534
rect 2819 2530 2839 2534
rect 2843 2530 2951 2534
rect 2955 2530 2967 2534
rect 2971 2530 3087 2534
rect 3091 2530 3095 2534
rect 3099 2530 3223 2534
rect 3227 2530 3367 2534
rect 3371 2530 3943 2534
rect 3947 2530 3967 2534
rect 2025 2529 3967 2530
rect 3973 2529 3974 2535
rect 84 2501 85 2507
rect 91 2506 2019 2507
rect 91 2502 111 2506
rect 115 2502 503 2506
rect 507 2502 575 2506
rect 579 2502 607 2506
rect 611 2502 687 2506
rect 691 2502 719 2506
rect 723 2502 807 2506
rect 811 2502 847 2506
rect 851 2502 935 2506
rect 939 2502 983 2506
rect 987 2502 1071 2506
rect 1075 2502 1127 2506
rect 1131 2502 1207 2506
rect 1211 2502 1279 2506
rect 1283 2502 1351 2506
rect 1355 2502 1431 2506
rect 1435 2502 1495 2506
rect 1499 2502 1583 2506
rect 1587 2502 1647 2506
rect 1651 2502 1743 2506
rect 1747 2502 1799 2506
rect 1803 2502 1903 2506
rect 1907 2502 2007 2506
rect 2011 2502 2019 2506
rect 91 2501 2019 2502
rect 2025 2501 2026 2507
rect 2030 2441 2031 2447
rect 2037 2446 3979 2447
rect 2037 2442 2047 2446
rect 2051 2442 2071 2446
rect 2075 2442 2095 2446
rect 2099 2442 2191 2446
rect 2195 2442 2215 2446
rect 2219 2442 2319 2446
rect 2323 2442 2343 2446
rect 2347 2442 2439 2446
rect 2443 2442 2471 2446
rect 2475 2442 2559 2446
rect 2563 2442 2599 2446
rect 2603 2442 2679 2446
rect 2683 2442 2719 2446
rect 2723 2442 2791 2446
rect 2795 2442 2839 2446
rect 2843 2442 2911 2446
rect 2915 2442 2967 2446
rect 2971 2442 3031 2446
rect 3035 2442 3095 2446
rect 3099 2442 3151 2446
rect 3155 2442 3223 2446
rect 3227 2442 3943 2446
rect 3947 2442 3979 2446
rect 2037 2441 3979 2442
rect 3985 2441 3986 2447
rect 96 2409 97 2415
rect 103 2414 2031 2415
rect 103 2410 111 2414
rect 115 2410 503 2414
rect 507 2410 535 2414
rect 539 2410 607 2414
rect 611 2410 671 2414
rect 675 2410 719 2414
rect 723 2410 815 2414
rect 819 2410 847 2414
rect 851 2410 959 2414
rect 963 2410 983 2414
rect 987 2410 1103 2414
rect 1107 2410 1127 2414
rect 1131 2410 1247 2414
rect 1251 2410 1279 2414
rect 1283 2410 1391 2414
rect 1395 2410 1431 2414
rect 1435 2410 1527 2414
rect 1531 2410 1583 2414
rect 1587 2410 1655 2414
rect 1659 2410 1743 2414
rect 1747 2410 1791 2414
rect 1795 2410 1903 2414
rect 1907 2410 2007 2414
rect 2011 2410 2031 2414
rect 103 2409 2031 2410
rect 2037 2409 2038 2415
rect 2018 2361 2019 2367
rect 2025 2366 3967 2367
rect 2025 2362 2047 2366
rect 2051 2362 2071 2366
rect 2075 2362 2167 2366
rect 2171 2362 2191 2366
rect 2195 2362 2319 2366
rect 2323 2362 2359 2366
rect 2363 2362 2439 2366
rect 2443 2362 2535 2366
rect 2539 2362 2559 2366
rect 2563 2362 2679 2366
rect 2683 2362 2703 2366
rect 2707 2362 2791 2366
rect 2795 2362 2871 2366
rect 2875 2362 2911 2366
rect 2915 2362 3031 2366
rect 3035 2362 3151 2366
rect 3155 2362 3199 2366
rect 3203 2362 3943 2366
rect 3947 2362 3967 2366
rect 2025 2361 3967 2362
rect 3973 2361 3974 2367
rect 84 2329 85 2335
rect 91 2334 2019 2335
rect 91 2330 111 2334
rect 115 2330 535 2334
rect 539 2330 647 2334
rect 651 2330 671 2334
rect 675 2330 767 2334
rect 771 2330 815 2334
rect 819 2330 895 2334
rect 899 2330 959 2334
rect 963 2330 1031 2334
rect 1035 2330 1103 2334
rect 1107 2330 1167 2334
rect 1171 2330 1247 2334
rect 1251 2330 1295 2334
rect 1299 2330 1391 2334
rect 1395 2330 1423 2334
rect 1427 2330 1527 2334
rect 1531 2330 1551 2334
rect 1555 2330 1655 2334
rect 1659 2330 1671 2334
rect 1675 2330 1791 2334
rect 1795 2330 1799 2334
rect 1803 2330 1903 2334
rect 1907 2330 2007 2334
rect 2011 2330 2019 2334
rect 91 2329 2019 2330
rect 2025 2329 2026 2335
rect 2030 2285 2031 2291
rect 2037 2290 3979 2291
rect 2037 2286 2047 2290
rect 2051 2286 2071 2290
rect 2075 2286 2167 2290
rect 2171 2286 2287 2290
rect 2291 2286 2359 2290
rect 2363 2286 2423 2290
rect 2427 2286 2535 2290
rect 2539 2286 2559 2290
rect 2563 2286 2703 2290
rect 2707 2286 2839 2290
rect 2843 2286 2871 2290
rect 2875 2286 2983 2290
rect 2987 2286 3031 2290
rect 3035 2286 3127 2290
rect 3131 2286 3199 2290
rect 3203 2286 3271 2290
rect 3275 2286 3943 2290
rect 3947 2286 3979 2290
rect 2037 2285 3979 2286
rect 3985 2285 3986 2291
rect 96 2249 97 2255
rect 103 2254 2031 2255
rect 103 2250 111 2254
rect 115 2250 415 2254
rect 419 2250 535 2254
rect 539 2250 647 2254
rect 651 2250 671 2254
rect 675 2250 767 2254
rect 771 2250 823 2254
rect 827 2250 895 2254
rect 899 2250 991 2254
rect 995 2250 1031 2254
rect 1035 2250 1167 2254
rect 1171 2250 1175 2254
rect 1179 2250 1295 2254
rect 1299 2250 1367 2254
rect 1371 2250 1423 2254
rect 1427 2250 1551 2254
rect 1555 2250 1567 2254
rect 1571 2250 1671 2254
rect 1675 2250 1767 2254
rect 1771 2250 1799 2254
rect 1803 2250 1903 2254
rect 1907 2250 2007 2254
rect 2011 2250 2031 2254
rect 103 2249 2031 2250
rect 2037 2249 2038 2255
rect 2018 2209 2019 2215
rect 2025 2214 3967 2215
rect 2025 2210 2047 2214
rect 2051 2210 2071 2214
rect 2075 2210 2167 2214
rect 2171 2210 2287 2214
rect 2291 2210 2295 2214
rect 2299 2210 2423 2214
rect 2427 2210 2503 2214
rect 2507 2210 2559 2214
rect 2563 2210 2687 2214
rect 2691 2210 2703 2214
rect 2707 2210 2839 2214
rect 2843 2210 2863 2214
rect 2867 2210 2983 2214
rect 2987 2210 3023 2214
rect 3027 2210 3127 2214
rect 3131 2210 3175 2214
rect 3179 2210 3271 2214
rect 3275 2210 3319 2214
rect 3323 2210 3471 2214
rect 3475 2210 3943 2214
rect 3947 2210 3967 2214
rect 2025 2209 3967 2210
rect 3973 2209 3974 2215
rect 84 2165 85 2171
rect 91 2170 2019 2171
rect 91 2166 111 2170
rect 115 2166 135 2170
rect 139 2166 247 2170
rect 251 2166 391 2170
rect 395 2166 415 2170
rect 419 2166 535 2170
rect 539 2166 551 2170
rect 555 2166 671 2170
rect 675 2166 711 2170
rect 715 2166 823 2170
rect 827 2166 871 2170
rect 875 2166 991 2170
rect 995 2166 1031 2170
rect 1035 2166 1175 2170
rect 1179 2166 1191 2170
rect 1195 2166 1351 2170
rect 1355 2166 1367 2170
rect 1371 2166 1511 2170
rect 1515 2166 1567 2170
rect 1571 2166 1679 2170
rect 1683 2166 1767 2170
rect 1771 2166 2007 2170
rect 2011 2166 2019 2170
rect 91 2165 2019 2166
rect 2025 2165 2026 2171
rect 2946 2124 2952 2125
rect 3438 2124 3444 2125
rect 2946 2120 2947 2124
rect 2951 2120 3439 2124
rect 3443 2120 3444 2124
rect 2946 2119 2952 2120
rect 3438 2119 3444 2120
rect 2030 2109 2031 2115
rect 2037 2114 3979 2115
rect 2037 2110 2047 2114
rect 2051 2110 2071 2114
rect 2075 2110 2295 2114
rect 2299 2110 2399 2114
rect 2403 2110 2495 2114
rect 2499 2110 2503 2114
rect 2507 2110 2591 2114
rect 2595 2110 2687 2114
rect 2691 2110 2783 2114
rect 2787 2110 2863 2114
rect 2867 2110 2879 2114
rect 2883 2110 2975 2114
rect 2979 2110 3023 2114
rect 3027 2110 3071 2114
rect 3075 2110 3167 2114
rect 3171 2110 3175 2114
rect 3179 2110 3263 2114
rect 3267 2110 3319 2114
rect 3323 2110 3359 2114
rect 3363 2110 3455 2114
rect 3459 2110 3471 2114
rect 3475 2110 3551 2114
rect 3555 2110 3647 2114
rect 3651 2110 3743 2114
rect 3747 2110 3839 2114
rect 3843 2110 3943 2114
rect 3947 2110 3979 2114
rect 2037 2109 3979 2110
rect 3985 2109 3986 2115
rect 96 2081 97 2087
rect 103 2086 2031 2087
rect 103 2082 111 2086
rect 115 2082 135 2086
rect 139 2082 247 2086
rect 251 2082 391 2086
rect 395 2082 399 2086
rect 403 2082 551 2086
rect 555 2082 703 2086
rect 707 2082 711 2086
rect 715 2082 847 2086
rect 851 2082 871 2086
rect 875 2082 991 2086
rect 995 2082 1031 2086
rect 1035 2082 1127 2086
rect 1131 2082 1191 2086
rect 1195 2082 1255 2086
rect 1259 2082 1351 2086
rect 1355 2082 1383 2086
rect 1387 2082 1511 2086
rect 1515 2082 1519 2086
rect 1523 2082 1679 2086
rect 1683 2082 2007 2086
rect 2011 2082 2031 2086
rect 103 2081 2031 2082
rect 2037 2081 2038 2087
rect 2018 2033 2019 2039
rect 2025 2038 3967 2039
rect 2025 2034 2047 2038
rect 2051 2034 2191 2038
rect 2195 2034 2399 2038
rect 2403 2034 2495 2038
rect 2499 2034 2591 2038
rect 2595 2034 2647 2038
rect 2651 2034 2687 2038
rect 2691 2034 2783 2038
rect 2787 2034 2879 2038
rect 2883 2034 2919 2038
rect 2923 2034 2975 2038
rect 2979 2034 3071 2038
rect 3075 2034 3167 2038
rect 3171 2034 3215 2038
rect 3219 2034 3263 2038
rect 3267 2034 3359 2038
rect 3363 2034 3455 2038
rect 3459 2034 3527 2038
rect 3531 2034 3551 2038
rect 3555 2034 3647 2038
rect 3651 2034 3743 2038
rect 3747 2034 3839 2038
rect 3843 2034 3943 2038
rect 3947 2034 3967 2038
rect 2025 2033 3967 2034
rect 3973 2033 3974 2039
rect 84 1989 85 1995
rect 91 1994 2019 1995
rect 91 1990 111 1994
rect 115 1990 135 1994
rect 139 1990 231 1994
rect 235 1990 247 1994
rect 251 1990 391 1994
rect 395 1990 399 1994
rect 403 1990 551 1994
rect 555 1990 567 1994
rect 571 1990 703 1994
rect 707 1990 751 1994
rect 755 1990 847 1994
rect 851 1990 943 1994
rect 947 1990 991 1994
rect 995 1990 1127 1994
rect 1131 1990 1135 1994
rect 1139 1990 1255 1994
rect 1259 1990 1335 1994
rect 1339 1990 1383 1994
rect 1387 1990 1519 1994
rect 1523 1990 1543 1994
rect 1547 1990 2007 1994
rect 2011 1990 2019 1994
rect 91 1989 2019 1990
rect 2025 1989 2026 1995
rect 2030 1945 2031 1951
rect 2037 1950 3979 1951
rect 2037 1946 2047 1950
rect 2051 1946 2071 1950
rect 2075 1946 2191 1950
rect 2195 1946 2239 1950
rect 2243 1946 2399 1950
rect 2403 1946 2447 1950
rect 2451 1946 2647 1950
rect 2651 1946 2671 1950
rect 2675 1946 2895 1950
rect 2899 1946 2919 1950
rect 2923 1946 3127 1950
rect 3131 1946 3215 1950
rect 3219 1946 3359 1950
rect 3363 1946 3527 1950
rect 3531 1946 3591 1950
rect 3595 1946 3831 1950
rect 3835 1946 3839 1950
rect 3843 1946 3943 1950
rect 3947 1946 3979 1950
rect 2037 1945 3979 1946
rect 3985 1945 3986 1951
rect 1202 1932 1208 1933
rect 1458 1932 1464 1933
rect 1202 1928 1203 1932
rect 1207 1928 1459 1932
rect 1463 1928 1464 1932
rect 1202 1927 1208 1928
rect 1458 1927 1464 1928
rect 96 1913 97 1919
rect 103 1918 2031 1919
rect 103 1914 111 1918
rect 115 1914 231 1918
rect 235 1914 391 1918
rect 395 1914 511 1918
rect 515 1914 567 1918
rect 571 1914 623 1918
rect 627 1914 743 1918
rect 747 1914 751 1918
rect 755 1914 863 1918
rect 867 1914 943 1918
rect 947 1914 983 1918
rect 987 1914 1103 1918
rect 1107 1914 1135 1918
rect 1139 1914 1223 1918
rect 1227 1914 1335 1918
rect 1339 1914 1455 1918
rect 1459 1914 1543 1918
rect 1547 1914 1575 1918
rect 1579 1914 1695 1918
rect 1699 1914 2007 1918
rect 2011 1914 2031 1918
rect 103 1913 2031 1914
rect 2037 1913 2038 1919
rect 2018 1869 2019 1875
rect 2025 1874 3967 1875
rect 2025 1870 2047 1874
rect 2051 1870 2071 1874
rect 2075 1870 2199 1874
rect 2203 1870 2239 1874
rect 2243 1870 2367 1874
rect 2371 1870 2447 1874
rect 2451 1870 2543 1874
rect 2547 1870 2671 1874
rect 2675 1870 2719 1874
rect 2723 1870 2887 1874
rect 2891 1870 2895 1874
rect 2899 1870 3039 1874
rect 3043 1870 3127 1874
rect 3131 1870 3183 1874
rect 3187 1870 3319 1874
rect 3323 1870 3359 1874
rect 3363 1870 3455 1874
rect 3459 1870 3583 1874
rect 3587 1870 3591 1874
rect 3595 1870 3711 1874
rect 3715 1870 3831 1874
rect 3835 1870 3839 1874
rect 3843 1870 3943 1874
rect 3947 1870 3967 1874
rect 2025 1869 3967 1870
rect 3973 1869 3974 1875
rect 84 1829 85 1835
rect 91 1834 2019 1835
rect 91 1830 111 1834
rect 115 1830 511 1834
rect 515 1830 615 1834
rect 619 1830 623 1834
rect 627 1830 711 1834
rect 715 1830 743 1834
rect 747 1830 815 1834
rect 819 1830 863 1834
rect 867 1830 927 1834
rect 931 1830 983 1834
rect 987 1830 1039 1834
rect 1043 1830 1103 1834
rect 1107 1830 1159 1834
rect 1163 1830 1223 1834
rect 1227 1830 1279 1834
rect 1283 1830 1335 1834
rect 1339 1830 1399 1834
rect 1403 1830 1455 1834
rect 1459 1830 1519 1834
rect 1523 1830 1575 1834
rect 1579 1830 1639 1834
rect 1643 1830 1695 1834
rect 1699 1830 2007 1834
rect 2011 1830 2019 1834
rect 91 1829 2019 1830
rect 2025 1829 2026 1835
rect 2030 1789 2031 1795
rect 2037 1794 3979 1795
rect 2037 1790 2047 1794
rect 2051 1790 2071 1794
rect 2075 1790 2183 1794
rect 2187 1790 2199 1794
rect 2203 1790 2327 1794
rect 2331 1790 2367 1794
rect 2371 1790 2487 1794
rect 2491 1790 2543 1794
rect 2547 1790 2655 1794
rect 2659 1790 2719 1794
rect 2723 1790 2831 1794
rect 2835 1790 2887 1794
rect 2891 1790 3023 1794
rect 3027 1790 3039 1794
rect 3043 1790 3183 1794
rect 3187 1790 3223 1794
rect 3227 1790 3319 1794
rect 3323 1790 3431 1794
rect 3435 1790 3455 1794
rect 3459 1790 3583 1794
rect 3587 1790 3647 1794
rect 3651 1790 3711 1794
rect 3715 1790 3839 1794
rect 3843 1790 3943 1794
rect 3947 1790 3979 1794
rect 2037 1789 3979 1790
rect 3985 1789 3986 1795
rect 96 1753 97 1759
rect 103 1758 2031 1759
rect 103 1754 111 1758
rect 115 1754 367 1758
rect 371 1754 495 1758
rect 499 1754 615 1758
rect 619 1754 639 1758
rect 643 1754 711 1758
rect 715 1754 799 1758
rect 803 1754 815 1758
rect 819 1754 927 1758
rect 931 1754 967 1758
rect 971 1754 1039 1758
rect 1043 1754 1143 1758
rect 1147 1754 1159 1758
rect 1163 1754 1279 1758
rect 1283 1754 1327 1758
rect 1331 1754 1399 1758
rect 1403 1754 1511 1758
rect 1515 1754 1519 1758
rect 1523 1754 1639 1758
rect 1643 1754 1703 1758
rect 1707 1754 2007 1758
rect 2011 1754 2031 1758
rect 103 1753 2031 1754
rect 2037 1753 2038 1759
rect 682 1740 688 1741
rect 918 1740 924 1741
rect 682 1736 683 1740
rect 687 1736 919 1740
rect 923 1736 924 1740
rect 682 1735 688 1736
rect 918 1735 924 1736
rect 2018 1705 2019 1711
rect 2025 1710 3967 1711
rect 2025 1706 2047 1710
rect 2051 1706 2071 1710
rect 2075 1706 2183 1710
rect 2187 1706 2223 1710
rect 2227 1706 2327 1710
rect 2331 1706 2439 1710
rect 2443 1706 2487 1710
rect 2491 1706 2559 1710
rect 2563 1706 2655 1710
rect 2659 1706 2687 1710
rect 2691 1706 2823 1710
rect 2827 1706 2831 1710
rect 2835 1706 2967 1710
rect 2971 1706 3023 1710
rect 3027 1706 3127 1710
rect 3131 1706 3223 1710
rect 3227 1706 3303 1710
rect 3307 1706 3431 1710
rect 3435 1706 3487 1710
rect 3491 1706 3647 1710
rect 3651 1706 3671 1710
rect 3675 1706 3839 1710
rect 3843 1706 3943 1710
rect 3947 1706 3967 1710
rect 2025 1705 3967 1706
rect 3973 1705 3974 1711
rect 84 1673 85 1679
rect 91 1678 2019 1679
rect 91 1674 111 1678
rect 115 1674 135 1678
rect 139 1674 247 1678
rect 251 1674 367 1678
rect 371 1674 399 1678
rect 403 1674 495 1678
rect 499 1674 567 1678
rect 571 1674 639 1678
rect 643 1674 743 1678
rect 747 1674 799 1678
rect 803 1674 935 1678
rect 939 1674 967 1678
rect 971 1674 1135 1678
rect 1139 1674 1143 1678
rect 1147 1674 1327 1678
rect 1331 1674 1343 1678
rect 1347 1674 1511 1678
rect 1515 1674 1551 1678
rect 1555 1674 1703 1678
rect 1707 1674 1767 1678
rect 1771 1674 2007 1678
rect 2011 1674 2019 1678
rect 91 1673 2019 1674
rect 2025 1673 2026 1679
rect 2030 1625 2031 1631
rect 2037 1630 3979 1631
rect 2037 1626 2047 1630
rect 2051 1626 2223 1630
rect 2227 1626 2327 1630
rect 2331 1626 2391 1630
rect 2395 1626 2439 1630
rect 2443 1626 2503 1630
rect 2507 1626 2559 1630
rect 2563 1626 2615 1630
rect 2619 1626 2687 1630
rect 2691 1626 2735 1630
rect 2739 1626 2823 1630
rect 2827 1626 2855 1630
rect 2859 1626 2967 1630
rect 2971 1626 2975 1630
rect 2979 1626 3095 1630
rect 3099 1626 3127 1630
rect 3131 1626 3215 1630
rect 3219 1626 3303 1630
rect 3307 1626 3335 1630
rect 3339 1626 3455 1630
rect 3459 1626 3487 1630
rect 3491 1626 3671 1630
rect 3675 1626 3839 1630
rect 3843 1626 3943 1630
rect 3947 1626 3979 1630
rect 2037 1625 3979 1626
rect 3985 1625 3986 1631
rect 96 1593 97 1599
rect 103 1598 2031 1599
rect 103 1594 111 1598
rect 115 1594 135 1598
rect 139 1594 247 1598
rect 251 1594 255 1598
rect 259 1594 399 1598
rect 403 1594 423 1598
rect 427 1594 567 1598
rect 571 1594 615 1598
rect 619 1594 743 1598
rect 747 1594 831 1598
rect 835 1594 935 1598
rect 939 1594 1063 1598
rect 1067 1594 1135 1598
rect 1139 1594 1311 1598
rect 1315 1594 1343 1598
rect 1347 1594 1551 1598
rect 1555 1594 1567 1598
rect 1571 1594 1767 1598
rect 1771 1594 1831 1598
rect 1835 1594 2007 1598
rect 2011 1594 2031 1598
rect 103 1593 2031 1594
rect 2037 1593 2038 1599
rect 2018 1549 2019 1555
rect 2025 1554 3967 1555
rect 2025 1550 2047 1554
rect 2051 1550 2391 1554
rect 2395 1550 2503 1554
rect 2507 1550 2543 1554
rect 2547 1550 2615 1554
rect 2619 1550 2671 1554
rect 2675 1550 2735 1554
rect 2739 1550 2799 1554
rect 2803 1550 2855 1554
rect 2859 1550 2935 1554
rect 2939 1550 2975 1554
rect 2979 1550 3071 1554
rect 3075 1550 3095 1554
rect 3099 1550 3207 1554
rect 3211 1550 3215 1554
rect 3219 1550 3335 1554
rect 3339 1550 3455 1554
rect 3459 1550 3463 1554
rect 3467 1550 3591 1554
rect 3595 1550 3727 1554
rect 3731 1550 3839 1554
rect 3843 1550 3943 1554
rect 3947 1550 3967 1554
rect 2025 1549 3967 1550
rect 3973 1549 3974 1555
rect 84 1513 85 1519
rect 91 1518 2019 1519
rect 91 1514 111 1518
rect 115 1514 135 1518
rect 139 1514 239 1518
rect 243 1514 255 1518
rect 259 1514 407 1518
rect 411 1514 423 1518
rect 427 1514 583 1518
rect 587 1514 615 1518
rect 619 1514 775 1518
rect 779 1514 831 1518
rect 835 1514 967 1518
rect 971 1514 1063 1518
rect 1067 1514 1159 1518
rect 1163 1514 1311 1518
rect 1315 1514 1351 1518
rect 1355 1514 1543 1518
rect 1547 1514 1567 1518
rect 1571 1514 1735 1518
rect 1739 1514 1831 1518
rect 1835 1514 1903 1518
rect 1907 1514 2007 1518
rect 2011 1514 2019 1518
rect 91 1513 2019 1514
rect 2025 1513 2026 1519
rect 2030 1461 2031 1467
rect 2037 1466 3979 1467
rect 2037 1462 2047 1466
rect 2051 1462 2519 1466
rect 2523 1462 2543 1466
rect 2547 1462 2631 1466
rect 2635 1462 2671 1466
rect 2675 1462 2759 1466
rect 2763 1462 2799 1466
rect 2803 1462 2895 1466
rect 2899 1462 2935 1466
rect 2939 1462 3031 1466
rect 3035 1462 3071 1466
rect 3075 1462 3175 1466
rect 3179 1462 3207 1466
rect 3211 1462 3311 1466
rect 3315 1462 3335 1466
rect 3339 1462 3447 1466
rect 3451 1462 3463 1466
rect 3467 1462 3583 1466
rect 3587 1462 3591 1466
rect 3595 1462 3719 1466
rect 3723 1462 3727 1466
rect 3731 1462 3839 1466
rect 3843 1462 3943 1466
rect 3947 1462 3979 1466
rect 2037 1461 3979 1462
rect 3985 1461 3986 1467
rect 96 1429 97 1435
rect 103 1434 2031 1435
rect 103 1430 111 1434
rect 115 1430 239 1434
rect 243 1430 407 1434
rect 411 1430 463 1434
rect 467 1430 583 1434
rect 587 1430 711 1434
rect 715 1430 775 1434
rect 779 1430 855 1434
rect 859 1430 967 1434
rect 971 1430 1007 1434
rect 1011 1430 1159 1434
rect 1163 1430 1167 1434
rect 1171 1430 1335 1434
rect 1339 1430 1351 1434
rect 1355 1430 1511 1434
rect 1515 1430 1543 1434
rect 1547 1430 1687 1434
rect 1691 1430 1735 1434
rect 1739 1430 1871 1434
rect 1875 1430 1903 1434
rect 1907 1430 2007 1434
rect 2011 1430 2031 1434
rect 103 1429 2031 1430
rect 2037 1429 2038 1435
rect 2018 1385 2019 1391
rect 2025 1390 3967 1391
rect 2025 1386 2047 1390
rect 2051 1386 2399 1390
rect 2403 1386 2519 1390
rect 2523 1386 2535 1390
rect 2539 1386 2631 1390
rect 2635 1386 2679 1390
rect 2683 1386 2759 1390
rect 2763 1386 2823 1390
rect 2827 1386 2895 1390
rect 2899 1386 2967 1390
rect 2971 1386 3031 1390
rect 3035 1386 3111 1390
rect 3115 1386 3175 1390
rect 3179 1386 3255 1390
rect 3259 1386 3311 1390
rect 3315 1386 3407 1390
rect 3411 1386 3447 1390
rect 3451 1386 3559 1390
rect 3563 1386 3583 1390
rect 3587 1386 3711 1390
rect 3715 1386 3719 1390
rect 3723 1386 3839 1390
rect 3843 1386 3943 1390
rect 3947 1386 3967 1390
rect 2025 1385 3967 1386
rect 3973 1385 3974 1391
rect 84 1353 85 1359
rect 91 1358 2019 1359
rect 91 1354 111 1358
rect 115 1354 463 1358
rect 467 1354 583 1358
rect 587 1354 655 1358
rect 659 1354 711 1358
rect 715 1354 767 1358
rect 771 1354 855 1358
rect 859 1354 887 1358
rect 891 1354 1007 1358
rect 1011 1354 1015 1358
rect 1019 1354 1143 1358
rect 1147 1354 1167 1358
rect 1171 1354 1279 1358
rect 1283 1354 1335 1358
rect 1339 1354 1415 1358
rect 1419 1354 1511 1358
rect 1515 1354 1559 1358
rect 1563 1354 1687 1358
rect 1691 1354 1703 1358
rect 1707 1354 1847 1358
rect 1851 1354 1871 1358
rect 1875 1354 2007 1358
rect 2011 1354 2019 1358
rect 91 1353 2019 1354
rect 2025 1353 2026 1359
rect 2030 1305 2031 1311
rect 2037 1310 3979 1311
rect 2037 1306 2047 1310
rect 2051 1306 2247 1310
rect 2251 1306 2375 1310
rect 2379 1306 2399 1310
rect 2403 1306 2511 1310
rect 2515 1306 2535 1310
rect 2539 1306 2647 1310
rect 2651 1306 2679 1310
rect 2683 1306 2791 1310
rect 2795 1306 2823 1310
rect 2827 1306 2943 1310
rect 2947 1306 2967 1310
rect 2971 1306 3111 1310
rect 3115 1306 3255 1310
rect 3259 1306 3287 1310
rect 3291 1306 3407 1310
rect 3411 1306 3471 1310
rect 3475 1306 3559 1310
rect 3563 1306 3663 1310
rect 3667 1306 3711 1310
rect 3715 1306 3839 1310
rect 3843 1306 3943 1310
rect 3947 1306 3979 1310
rect 2037 1305 3979 1306
rect 3985 1305 3986 1311
rect 96 1273 97 1279
rect 103 1278 2031 1279
rect 103 1274 111 1278
rect 115 1274 439 1278
rect 443 1274 551 1278
rect 555 1274 655 1278
rect 659 1274 671 1278
rect 675 1274 767 1278
rect 771 1274 799 1278
rect 803 1274 887 1278
rect 891 1274 935 1278
rect 939 1274 1015 1278
rect 1019 1274 1079 1278
rect 1083 1274 1143 1278
rect 1147 1274 1231 1278
rect 1235 1274 1279 1278
rect 1283 1274 1391 1278
rect 1395 1274 1415 1278
rect 1419 1274 1551 1278
rect 1555 1274 1559 1278
rect 1563 1274 1703 1278
rect 1707 1274 1719 1278
rect 1723 1274 1847 1278
rect 1851 1274 2007 1278
rect 2011 1274 2031 1278
rect 103 1273 2031 1274
rect 2037 1273 2038 1279
rect 2018 1225 2019 1231
rect 2025 1230 3967 1231
rect 2025 1226 2047 1230
rect 2051 1226 2071 1230
rect 2075 1226 2183 1230
rect 2187 1226 2247 1230
rect 2251 1226 2303 1230
rect 2307 1226 2375 1230
rect 2379 1226 2431 1230
rect 2435 1226 2511 1230
rect 2515 1226 2559 1230
rect 2563 1226 2647 1230
rect 2651 1226 2711 1230
rect 2715 1226 2791 1230
rect 2795 1226 2887 1230
rect 2891 1226 2943 1230
rect 2947 1226 3087 1230
rect 3091 1226 3111 1230
rect 3115 1226 3287 1230
rect 3291 1226 3311 1230
rect 3315 1226 3471 1230
rect 3475 1226 3543 1230
rect 3547 1226 3663 1230
rect 3667 1226 3783 1230
rect 3787 1226 3839 1230
rect 3843 1226 3943 1230
rect 3947 1226 3967 1230
rect 2025 1225 3967 1226
rect 3973 1225 3974 1231
rect 84 1197 85 1203
rect 91 1202 2019 1203
rect 91 1198 111 1202
rect 115 1198 167 1202
rect 171 1198 303 1202
rect 307 1198 439 1202
rect 443 1198 463 1202
rect 467 1198 551 1202
rect 555 1198 631 1202
rect 635 1198 671 1202
rect 675 1198 799 1202
rect 803 1198 807 1202
rect 811 1198 935 1202
rect 939 1198 983 1202
rect 987 1198 1079 1202
rect 1083 1198 1159 1202
rect 1163 1198 1231 1202
rect 1235 1198 1335 1202
rect 1339 1198 1391 1202
rect 1395 1198 1511 1202
rect 1515 1198 1551 1202
rect 1555 1198 1695 1202
rect 1699 1198 1719 1202
rect 1723 1198 2007 1202
rect 2011 1198 2019 1202
rect 91 1197 2019 1198
rect 2025 1197 2026 1203
rect 2030 1145 2031 1151
rect 2037 1150 3979 1151
rect 2037 1146 2047 1150
rect 2051 1146 2071 1150
rect 2075 1146 2183 1150
rect 2187 1146 2199 1150
rect 2203 1146 2303 1150
rect 2307 1146 2351 1150
rect 2355 1146 2431 1150
rect 2435 1146 2511 1150
rect 2515 1146 2559 1150
rect 2563 1146 2679 1150
rect 2683 1146 2711 1150
rect 2715 1146 2871 1150
rect 2875 1146 2887 1150
rect 2891 1146 3087 1150
rect 3091 1146 3311 1150
rect 3315 1146 3319 1150
rect 3323 1146 3543 1150
rect 3547 1146 3559 1150
rect 3563 1146 3783 1150
rect 3787 1146 3807 1150
rect 3811 1146 3943 1150
rect 3947 1146 3979 1150
rect 2037 1145 3979 1146
rect 3985 1145 3986 1151
rect 96 1117 97 1123
rect 103 1122 2031 1123
rect 103 1118 111 1122
rect 115 1118 135 1122
rect 139 1118 167 1122
rect 171 1118 239 1122
rect 243 1118 303 1122
rect 307 1118 375 1122
rect 379 1118 463 1122
rect 467 1118 527 1122
rect 531 1118 631 1122
rect 635 1118 695 1122
rect 699 1118 807 1122
rect 811 1118 863 1122
rect 867 1118 983 1122
rect 987 1118 1039 1122
rect 1043 1118 1159 1122
rect 1163 1118 1215 1122
rect 1219 1118 1335 1122
rect 1339 1118 1391 1122
rect 1395 1118 1511 1122
rect 1515 1118 1567 1122
rect 1571 1118 1695 1122
rect 1699 1118 1743 1122
rect 1747 1118 1903 1122
rect 1907 1118 2007 1122
rect 2011 1118 2031 1122
rect 103 1117 2031 1118
rect 2037 1117 2038 1123
rect 2018 1057 2019 1063
rect 2025 1062 3967 1063
rect 2025 1058 2047 1062
rect 2051 1058 2071 1062
rect 2075 1058 2199 1062
rect 2203 1058 2263 1062
rect 2267 1058 2351 1062
rect 2355 1058 2487 1062
rect 2491 1058 2511 1062
rect 2515 1058 2679 1062
rect 2683 1058 2703 1062
rect 2707 1058 2871 1062
rect 2875 1058 2919 1062
rect 2923 1058 3087 1062
rect 3091 1058 3119 1062
rect 3123 1058 3311 1062
rect 3315 1058 3319 1062
rect 3323 1058 3495 1062
rect 3499 1058 3559 1062
rect 3563 1058 3679 1062
rect 3683 1058 3807 1062
rect 3811 1058 3839 1062
rect 3843 1058 3943 1062
rect 3947 1058 3967 1062
rect 2025 1057 3967 1058
rect 3973 1057 3974 1063
rect 84 1041 85 1047
rect 91 1046 2019 1047
rect 91 1042 111 1046
rect 115 1042 135 1046
rect 139 1042 239 1046
rect 243 1042 287 1046
rect 291 1042 375 1046
rect 379 1042 471 1046
rect 475 1042 527 1046
rect 531 1042 655 1046
rect 659 1042 695 1046
rect 699 1042 839 1046
rect 843 1042 863 1046
rect 867 1042 1015 1046
rect 1019 1042 1039 1046
rect 1043 1042 1199 1046
rect 1203 1042 1215 1046
rect 1219 1042 1383 1046
rect 1387 1042 1391 1046
rect 1395 1042 1567 1046
rect 1571 1042 1743 1046
rect 1747 1042 1903 1046
rect 1907 1042 2007 1046
rect 2011 1042 2019 1046
rect 91 1041 2019 1042
rect 2025 1041 2026 1047
rect 2030 977 2031 983
rect 2037 982 3979 983
rect 2037 978 2047 982
rect 2051 978 2071 982
rect 2075 978 2263 982
rect 2267 978 2303 982
rect 2307 978 2455 982
rect 2459 978 2487 982
rect 2491 978 2615 982
rect 2619 978 2703 982
rect 2707 978 2783 982
rect 2787 978 2919 982
rect 2923 978 2951 982
rect 2955 978 3111 982
rect 3115 978 3119 982
rect 3123 978 3263 982
rect 3267 978 3311 982
rect 3315 978 3415 982
rect 3419 978 3495 982
rect 3499 978 3559 982
rect 3563 978 3679 982
rect 3683 978 3711 982
rect 3715 978 3839 982
rect 3843 978 3943 982
rect 3947 978 3979 982
rect 2037 977 3979 978
rect 3985 977 3986 983
rect 96 961 97 967
rect 103 966 2031 967
rect 103 962 111 966
rect 115 962 135 966
rect 139 962 287 966
rect 291 962 295 966
rect 299 962 471 966
rect 475 962 639 966
rect 643 962 655 966
rect 659 962 799 966
rect 803 962 839 966
rect 843 962 951 966
rect 955 962 1015 966
rect 1019 962 1087 966
rect 1091 962 1199 966
rect 1203 962 1223 966
rect 1227 962 1359 966
rect 1363 962 1383 966
rect 1387 962 1495 966
rect 1499 962 1567 966
rect 1571 962 2007 966
rect 2011 962 2031 966
rect 103 961 2031 962
rect 2037 961 2038 967
rect 2018 897 2019 903
rect 2025 902 3967 903
rect 2025 898 2047 902
rect 2051 898 2303 902
rect 2307 898 2455 902
rect 2459 898 2559 902
rect 2563 898 2615 902
rect 2619 898 2679 902
rect 2683 898 2783 902
rect 2787 898 2807 902
rect 2811 898 2943 902
rect 2947 898 2951 902
rect 2955 898 3079 902
rect 3083 898 3111 902
rect 3115 898 3207 902
rect 3211 898 3263 902
rect 3267 898 3335 902
rect 3339 898 3415 902
rect 3419 898 3463 902
rect 3467 898 3559 902
rect 3563 898 3591 902
rect 3595 898 3711 902
rect 3715 898 3727 902
rect 3731 898 3839 902
rect 3843 898 3943 902
rect 3947 898 3967 902
rect 2025 897 3967 898
rect 3973 897 3974 903
rect 84 885 85 891
rect 91 890 2019 891
rect 91 886 111 890
rect 115 886 135 890
rect 139 886 159 890
rect 163 886 295 890
rect 299 886 319 890
rect 323 886 471 890
rect 475 886 615 890
rect 619 886 639 890
rect 643 886 751 890
rect 755 886 799 890
rect 803 886 879 890
rect 883 886 951 890
rect 955 886 999 890
rect 1003 886 1087 890
rect 1091 886 1111 890
rect 1115 886 1223 890
rect 1227 886 1231 890
rect 1235 886 1351 890
rect 1355 886 1359 890
rect 1363 886 1495 890
rect 1499 886 2007 890
rect 2011 886 2019 890
rect 91 885 2019 886
rect 2025 885 2026 891
rect 2030 817 2031 823
rect 2037 822 3979 823
rect 2037 818 2047 822
rect 2051 818 2335 822
rect 2339 818 2471 822
rect 2475 818 2559 822
rect 2563 818 2615 822
rect 2619 818 2679 822
rect 2683 818 2767 822
rect 2771 818 2807 822
rect 2811 818 2919 822
rect 2923 818 2943 822
rect 2947 818 3079 822
rect 3083 818 3207 822
rect 3211 818 3239 822
rect 3243 818 3335 822
rect 3339 818 3391 822
rect 3395 818 3463 822
rect 3467 818 3543 822
rect 3547 818 3591 822
rect 3595 818 3703 822
rect 3707 818 3727 822
rect 3731 818 3839 822
rect 3843 818 3943 822
rect 3947 818 3979 822
rect 2037 817 3979 818
rect 3985 817 3986 823
rect 2030 815 2038 817
rect 96 809 97 815
rect 103 814 2031 815
rect 103 810 111 814
rect 115 810 159 814
rect 163 810 223 814
rect 227 810 319 814
rect 323 810 383 814
rect 387 810 471 814
rect 475 810 535 814
rect 539 810 615 814
rect 619 810 679 814
rect 683 810 751 814
rect 755 810 815 814
rect 819 810 879 814
rect 883 810 951 814
rect 955 810 999 814
rect 1003 810 1079 814
rect 1083 810 1111 814
rect 1115 810 1199 814
rect 1203 810 1231 814
rect 1235 810 1327 814
rect 1331 810 1351 814
rect 1355 810 1455 814
rect 1459 810 2007 814
rect 2011 810 2031 814
rect 103 809 2031 810
rect 2037 809 2038 815
rect 2018 737 2019 743
rect 2025 742 3967 743
rect 2025 738 2047 742
rect 2051 738 2071 742
rect 2075 738 2183 742
rect 2187 738 2335 742
rect 2339 738 2471 742
rect 2475 738 2487 742
rect 2491 738 2615 742
rect 2619 738 2639 742
rect 2643 738 2767 742
rect 2771 738 2807 742
rect 2811 738 2919 742
rect 2923 738 2983 742
rect 2987 738 3079 742
rect 3083 738 3167 742
rect 3171 738 3239 742
rect 3243 738 3367 742
rect 3371 738 3391 742
rect 3395 738 3543 742
rect 3547 738 3575 742
rect 3579 738 3703 742
rect 3707 738 3783 742
rect 3787 738 3839 742
rect 3843 738 3943 742
rect 3947 738 3967 742
rect 2025 737 3967 738
rect 3973 737 3974 743
rect 2018 735 2026 737
rect 84 729 85 735
rect 91 734 2019 735
rect 91 730 111 734
rect 115 730 223 734
rect 227 730 311 734
rect 315 730 383 734
rect 387 730 471 734
rect 475 730 535 734
rect 539 730 639 734
rect 643 730 679 734
rect 683 730 807 734
rect 811 730 815 734
rect 819 730 951 734
rect 955 730 975 734
rect 979 730 1079 734
rect 1083 730 1135 734
rect 1139 730 1199 734
rect 1203 730 1295 734
rect 1299 730 1327 734
rect 1331 730 1455 734
rect 1459 730 1607 734
rect 1611 730 1767 734
rect 1771 730 1903 734
rect 1907 730 2007 734
rect 2011 730 2019 734
rect 91 729 2019 730
rect 2025 729 2026 735
rect 1202 668 1208 669
rect 1698 668 1704 669
rect 1202 664 1203 668
rect 1207 664 1699 668
rect 1703 664 1704 668
rect 1202 663 1208 664
rect 1698 663 1704 664
rect 96 653 97 659
rect 103 658 2031 659
rect 103 654 111 658
rect 115 654 295 658
rect 299 654 311 658
rect 315 654 447 658
rect 451 654 471 658
rect 475 654 615 658
rect 619 654 639 658
rect 643 654 783 658
rect 787 654 807 658
rect 811 654 951 658
rect 955 654 975 658
rect 979 654 1111 658
rect 1115 654 1135 658
rect 1139 654 1263 658
rect 1267 654 1295 658
rect 1299 654 1399 658
rect 1403 654 1455 658
rect 1459 654 1535 658
rect 1539 654 1607 658
rect 1611 654 1663 658
rect 1667 654 1767 658
rect 1771 654 1791 658
rect 1795 654 1903 658
rect 1907 654 2007 658
rect 2011 654 2031 658
rect 103 653 2031 654
rect 2037 655 2038 659
rect 2037 654 3986 655
rect 2037 653 2047 654
rect 2030 650 2047 653
rect 2051 650 2071 654
rect 2075 650 2183 654
rect 2187 650 2239 654
rect 2243 650 2335 654
rect 2339 650 2423 654
rect 2427 650 2487 654
rect 2491 650 2623 654
rect 2627 650 2639 654
rect 2643 650 2807 654
rect 2811 650 2839 654
rect 2843 650 2983 654
rect 2987 650 3071 654
rect 3075 650 3167 654
rect 3171 650 3319 654
rect 3323 650 3367 654
rect 3371 650 3575 654
rect 3579 650 3783 654
rect 3787 650 3839 654
rect 3843 650 3943 654
rect 3947 650 3986 654
rect 2030 649 3986 650
rect 84 573 85 579
rect 91 578 2019 579
rect 91 574 111 578
rect 115 574 239 578
rect 243 574 295 578
rect 299 574 415 578
rect 419 574 447 578
rect 451 574 607 578
rect 611 574 615 578
rect 619 574 783 578
rect 787 574 799 578
rect 803 574 951 578
rect 955 574 991 578
rect 995 574 1111 578
rect 1115 574 1175 578
rect 1179 574 1263 578
rect 1267 574 1351 578
rect 1355 574 1399 578
rect 1403 574 1519 578
rect 1523 574 1535 578
rect 1539 574 1663 578
rect 1667 574 1687 578
rect 1691 574 1791 578
rect 1795 574 1863 578
rect 1867 574 1903 578
rect 1907 574 2007 578
rect 2011 574 2019 578
rect 91 573 2019 574
rect 2025 578 3974 579
rect 2025 574 2047 578
rect 2051 574 2071 578
rect 2075 574 2191 578
rect 2195 574 2239 578
rect 2243 574 2287 578
rect 2291 574 2383 578
rect 2387 574 2423 578
rect 2427 574 2479 578
rect 2483 574 2583 578
rect 2587 574 2623 578
rect 2627 574 2711 578
rect 2715 574 2839 578
rect 2843 574 2871 578
rect 2875 574 3071 578
rect 3075 574 3303 578
rect 3307 574 3319 578
rect 3323 574 3551 578
rect 3555 574 3575 578
rect 3579 574 3807 578
rect 3811 574 3839 578
rect 3843 574 3943 578
rect 3947 574 3974 578
rect 2025 573 3974 574
rect 96 497 97 503
rect 103 502 2031 503
rect 103 498 111 502
rect 115 498 135 502
rect 139 498 239 502
rect 243 498 287 502
rect 291 498 415 502
rect 419 498 463 502
rect 467 498 607 502
rect 611 498 639 502
rect 643 498 799 502
rect 803 498 807 502
rect 811 498 967 502
rect 971 498 991 502
rect 995 498 1119 502
rect 1123 498 1175 502
rect 1179 498 1271 502
rect 1275 498 1351 502
rect 1355 498 1415 502
rect 1419 498 1519 502
rect 1523 498 1567 502
rect 1571 498 1687 502
rect 1691 498 1863 502
rect 1867 498 2007 502
rect 2011 498 2031 502
rect 103 497 2031 498
rect 2037 502 3986 503
rect 2037 498 2047 502
rect 2051 498 2191 502
rect 2195 498 2287 502
rect 2291 498 2383 502
rect 2387 498 2431 502
rect 2435 498 2479 502
rect 2483 498 2527 502
rect 2531 498 2583 502
rect 2587 498 2623 502
rect 2627 498 2711 502
rect 2715 498 2727 502
rect 2731 498 2847 502
rect 2851 498 2871 502
rect 2875 498 2999 502
rect 3003 498 3071 502
rect 3075 498 3175 502
rect 3179 498 3303 502
rect 3307 498 3375 502
rect 3379 498 3551 502
rect 3555 498 3591 502
rect 3595 498 3807 502
rect 3811 498 3943 502
rect 3947 498 3986 502
rect 2037 497 3986 498
rect 2018 426 3974 427
rect 2018 423 2047 426
rect 84 417 85 423
rect 91 422 2019 423
rect 91 418 111 422
rect 115 418 135 422
rect 139 418 279 422
rect 283 418 287 422
rect 291 418 439 422
rect 443 418 463 422
rect 467 418 583 422
rect 587 418 639 422
rect 643 418 719 422
rect 723 418 807 422
rect 811 418 847 422
rect 851 418 967 422
rect 971 418 1087 422
rect 1091 418 1119 422
rect 1123 418 1207 422
rect 1211 418 1271 422
rect 1275 418 1327 422
rect 1331 418 1415 422
rect 1419 418 1567 422
rect 1571 418 2007 422
rect 2011 418 2019 422
rect 91 417 2019 418
rect 2025 422 2047 423
rect 2051 422 2431 426
rect 2435 422 2527 426
rect 2531 422 2623 426
rect 2627 422 2719 426
rect 2723 422 2727 426
rect 2731 422 2815 426
rect 2819 422 2847 426
rect 2851 422 2927 426
rect 2931 422 2999 426
rect 3003 422 3063 426
rect 3067 422 3175 426
rect 3179 422 3223 426
rect 3227 422 3375 426
rect 3379 422 3399 426
rect 3403 422 3591 426
rect 3595 422 3783 426
rect 3787 422 3807 426
rect 3811 422 3943 426
rect 3947 422 3974 426
rect 2025 421 3974 422
rect 2025 417 2026 421
rect 96 341 97 347
rect 103 346 2031 347
rect 103 342 111 346
rect 115 342 135 346
rect 139 342 143 346
rect 147 342 279 346
rect 283 342 319 346
rect 323 342 439 346
rect 443 342 479 346
rect 483 342 583 346
rect 587 342 631 346
rect 635 342 719 346
rect 723 342 775 346
rect 779 342 847 346
rect 851 342 903 346
rect 907 342 967 346
rect 971 342 1031 346
rect 1035 342 1087 346
rect 1091 342 1151 346
rect 1155 342 1207 346
rect 1211 342 1271 346
rect 1275 342 1327 346
rect 1331 342 1391 346
rect 1395 342 2007 346
rect 2011 342 2031 346
rect 103 341 2031 342
rect 2037 346 3986 347
rect 2037 342 2047 346
rect 2051 342 2191 346
rect 2195 342 2327 346
rect 2331 342 2431 346
rect 2435 342 2471 346
rect 2475 342 2527 346
rect 2531 342 2623 346
rect 2627 342 2719 346
rect 2723 342 2783 346
rect 2787 342 2815 346
rect 2819 342 2927 346
rect 2931 342 2951 346
rect 2955 342 3063 346
rect 3067 342 3119 346
rect 3123 342 3223 346
rect 3227 342 3295 346
rect 3299 342 3399 346
rect 3403 342 3471 346
rect 3475 342 3591 346
rect 3595 342 3655 346
rect 3659 342 3783 346
rect 3787 342 3839 346
rect 3843 342 3943 346
rect 3947 342 3986 346
rect 2037 341 3986 342
rect 2018 270 3974 271
rect 2018 267 2047 270
rect 84 261 85 267
rect 91 266 2019 267
rect 91 262 111 266
rect 115 262 143 266
rect 147 262 223 266
rect 227 262 319 266
rect 323 262 391 266
rect 395 262 479 266
rect 483 262 559 266
rect 563 262 631 266
rect 635 262 735 266
rect 739 262 775 266
rect 779 262 903 266
rect 907 262 1031 266
rect 1035 262 1063 266
rect 1067 262 1151 266
rect 1155 262 1215 266
rect 1219 262 1271 266
rect 1275 262 1359 266
rect 1363 262 1391 266
rect 1395 262 1511 266
rect 1515 262 1663 266
rect 1667 262 2007 266
rect 2011 262 2019 266
rect 91 261 2019 262
rect 2025 266 2047 267
rect 2051 266 2071 270
rect 2075 266 2191 270
rect 2195 266 2215 270
rect 2219 266 2327 270
rect 2331 266 2399 270
rect 2403 266 2471 270
rect 2475 266 2591 270
rect 2595 266 2623 270
rect 2627 266 2783 270
rect 2787 266 2791 270
rect 2795 266 2951 270
rect 2955 266 2983 270
rect 2987 266 3119 270
rect 3123 266 3167 270
rect 3171 266 3295 270
rect 3299 266 3343 270
rect 3347 266 3471 270
rect 3475 266 3511 270
rect 3515 266 3655 270
rect 3659 266 3687 270
rect 3691 266 3839 270
rect 3843 266 3943 270
rect 3947 266 3974 270
rect 2025 265 3974 266
rect 2025 261 2026 265
rect 2030 165 2031 171
rect 2037 170 3979 171
rect 2037 166 2047 170
rect 2051 166 2071 170
rect 2075 166 2191 170
rect 2195 166 2215 170
rect 2219 166 2343 170
rect 2347 166 2399 170
rect 2403 166 2495 170
rect 2499 166 2591 170
rect 2595 166 2647 170
rect 2651 166 2791 170
rect 2795 166 2799 170
rect 2803 166 2943 170
rect 2947 166 2983 170
rect 2987 166 3071 170
rect 3075 166 3167 170
rect 3171 166 3191 170
rect 3195 166 3311 170
rect 3315 166 3343 170
rect 3347 166 3423 170
rect 3427 166 3511 170
rect 3515 166 3527 170
rect 3531 166 3639 170
rect 3643 166 3687 170
rect 3691 166 3743 170
rect 3747 166 3839 170
rect 3843 166 3943 170
rect 3947 166 3979 170
rect 2037 165 3979 166
rect 3985 165 3986 171
rect 96 153 97 159
rect 103 158 2031 159
rect 103 154 111 158
rect 115 154 151 158
rect 155 154 223 158
rect 227 154 247 158
rect 251 154 343 158
rect 347 154 391 158
rect 395 154 439 158
rect 443 154 535 158
rect 539 154 559 158
rect 563 154 631 158
rect 635 154 727 158
rect 731 154 735 158
rect 739 154 823 158
rect 827 154 903 158
rect 907 154 919 158
rect 923 154 1015 158
rect 1019 154 1063 158
rect 1067 154 1111 158
rect 1115 154 1207 158
rect 1211 154 1215 158
rect 1219 154 1303 158
rect 1307 154 1359 158
rect 1363 154 1407 158
rect 1411 154 1511 158
rect 1515 154 1615 158
rect 1619 154 1663 158
rect 1667 154 1711 158
rect 1715 154 1807 158
rect 1811 154 1903 158
rect 1907 154 2007 158
rect 2011 154 2031 158
rect 103 153 2031 154
rect 2037 153 2038 159
rect 2018 89 2019 95
rect 2025 94 3967 95
rect 2025 90 2047 94
rect 2051 90 2071 94
rect 2075 90 2191 94
rect 2195 90 2343 94
rect 2347 90 2495 94
rect 2499 90 2647 94
rect 2651 90 2799 94
rect 2803 90 2943 94
rect 2947 90 3071 94
rect 3075 90 3191 94
rect 3195 90 3311 94
rect 3315 90 3423 94
rect 3427 90 3527 94
rect 3531 90 3639 94
rect 3643 90 3743 94
rect 3747 90 3839 94
rect 3843 90 3943 94
rect 3947 90 3967 94
rect 2025 89 3967 90
rect 3973 89 3974 95
rect 84 77 85 83
rect 91 82 2019 83
rect 91 78 111 82
rect 115 78 151 82
rect 155 78 247 82
rect 251 78 343 82
rect 347 78 439 82
rect 443 78 535 82
rect 539 78 631 82
rect 635 78 727 82
rect 731 78 823 82
rect 827 78 919 82
rect 923 78 1015 82
rect 1019 78 1111 82
rect 1115 78 1207 82
rect 1211 78 1303 82
rect 1307 78 1407 82
rect 1411 78 1511 82
rect 1515 78 1615 82
rect 1619 78 1711 82
rect 1715 78 1807 82
rect 1811 78 1903 82
rect 1907 78 2007 82
rect 2011 78 2019 82
rect 91 77 2019 78
rect 2025 77 2026 83
<< m5c >>
rect 2019 4017 2025 4023
rect 3967 4017 3973 4023
rect 85 3997 91 4003
rect 2019 3997 2025 4003
rect 2031 3941 2037 3947
rect 3979 3941 3985 3947
rect 97 3921 103 3927
rect 2031 3921 2037 3927
rect 2019 3865 2025 3871
rect 3967 3865 3973 3871
rect 85 3837 91 3843
rect 2019 3837 2025 3843
rect 2031 3773 2037 3779
rect 3979 3773 3985 3779
rect 97 3761 103 3767
rect 2031 3761 2037 3767
rect 2019 3685 2025 3691
rect 3967 3685 3973 3691
rect 85 3677 91 3683
rect 2019 3677 2025 3683
rect 2031 3605 2037 3611
rect 3979 3605 3985 3611
rect 97 3597 103 3603
rect 2031 3597 2037 3603
rect 2019 3525 2025 3531
rect 3967 3525 3973 3531
rect 85 3513 91 3519
rect 2019 3513 2025 3519
rect 2031 3449 2037 3455
rect 3979 3449 3985 3455
rect 97 3417 103 3423
rect 2031 3417 2037 3423
rect 2019 3361 2025 3367
rect 3967 3361 3973 3367
rect 85 3329 91 3335
rect 2019 3329 2025 3335
rect 2031 3281 2037 3287
rect 3979 3281 3985 3287
rect 97 3249 103 3255
rect 2031 3249 2037 3255
rect 2019 3193 2025 3199
rect 3967 3193 3973 3199
rect 85 3165 91 3171
rect 2019 3165 2025 3171
rect 2031 3113 2037 3119
rect 3979 3113 3985 3119
rect 97 3089 103 3095
rect 2031 3089 2037 3095
rect 2019 3029 2025 3035
rect 3967 3029 3973 3035
rect 85 2989 91 2995
rect 2019 2989 2025 2995
rect 2031 2949 2037 2955
rect 3979 2949 3985 2955
rect 97 2913 103 2919
rect 2031 2913 2037 2919
rect 2019 2865 2025 2871
rect 3967 2865 3973 2871
rect 85 2833 91 2839
rect 2019 2833 2025 2839
rect 2031 2789 2037 2795
rect 3979 2789 3985 2795
rect 97 2749 103 2755
rect 2031 2749 2037 2755
rect 2019 2693 2025 2699
rect 3967 2693 3973 2699
rect 85 2673 91 2679
rect 2019 2673 2025 2679
rect 2031 2609 2037 2615
rect 3979 2609 3985 2615
rect 97 2581 103 2587
rect 2031 2581 2037 2587
rect 2019 2529 2025 2535
rect 3967 2529 3973 2535
rect 85 2501 91 2507
rect 2019 2501 2025 2507
rect 2031 2441 2037 2447
rect 3979 2441 3985 2447
rect 97 2409 103 2415
rect 2031 2409 2037 2415
rect 2019 2361 2025 2367
rect 3967 2361 3973 2367
rect 85 2329 91 2335
rect 2019 2329 2025 2335
rect 2031 2285 2037 2291
rect 3979 2285 3985 2291
rect 97 2249 103 2255
rect 2031 2249 2037 2255
rect 2019 2209 2025 2215
rect 3967 2209 3973 2215
rect 85 2165 91 2171
rect 2019 2165 2025 2171
rect 2031 2109 2037 2115
rect 3979 2109 3985 2115
rect 97 2081 103 2087
rect 2031 2081 2037 2087
rect 2019 2033 2025 2039
rect 3967 2033 3973 2039
rect 85 1989 91 1995
rect 2019 1989 2025 1995
rect 2031 1945 2037 1951
rect 3979 1945 3985 1951
rect 97 1913 103 1919
rect 2031 1913 2037 1919
rect 2019 1869 2025 1875
rect 3967 1869 3973 1875
rect 85 1829 91 1835
rect 2019 1829 2025 1835
rect 2031 1789 2037 1795
rect 3979 1789 3985 1795
rect 97 1753 103 1759
rect 2031 1753 2037 1759
rect 2019 1705 2025 1711
rect 3967 1705 3973 1711
rect 85 1673 91 1679
rect 2019 1673 2025 1679
rect 2031 1625 2037 1631
rect 3979 1625 3985 1631
rect 97 1593 103 1599
rect 2031 1593 2037 1599
rect 2019 1549 2025 1555
rect 3967 1549 3973 1555
rect 85 1513 91 1519
rect 2019 1513 2025 1519
rect 2031 1461 2037 1467
rect 3979 1461 3985 1467
rect 97 1429 103 1435
rect 2031 1429 2037 1435
rect 2019 1385 2025 1391
rect 3967 1385 3973 1391
rect 85 1353 91 1359
rect 2019 1353 2025 1359
rect 2031 1305 2037 1311
rect 3979 1305 3985 1311
rect 97 1273 103 1279
rect 2031 1273 2037 1279
rect 2019 1225 2025 1231
rect 3967 1225 3973 1231
rect 85 1197 91 1203
rect 2019 1197 2025 1203
rect 2031 1145 2037 1151
rect 3979 1145 3985 1151
rect 97 1117 103 1123
rect 2031 1117 2037 1123
rect 2019 1057 2025 1063
rect 3967 1057 3973 1063
rect 85 1041 91 1047
rect 2019 1041 2025 1047
rect 2031 977 2037 983
rect 3979 977 3985 983
rect 97 961 103 967
rect 2031 961 2037 967
rect 2019 897 2025 903
rect 3967 897 3973 903
rect 85 885 91 891
rect 2019 885 2025 891
rect 2031 817 2037 823
rect 3979 817 3985 823
rect 97 809 103 815
rect 2031 809 2037 815
rect 2019 737 2025 743
rect 3967 737 3973 743
rect 85 729 91 735
rect 2019 729 2025 735
rect 97 653 103 659
rect 2031 653 2037 659
rect 85 573 91 579
rect 2019 573 2025 579
rect 97 497 103 503
rect 2031 497 2037 503
rect 85 417 91 423
rect 2019 417 2025 423
rect 97 341 103 347
rect 2031 341 2037 347
rect 85 261 91 267
rect 2019 261 2025 267
rect 2031 165 2037 171
rect 3979 165 3985 171
rect 97 153 103 159
rect 2031 153 2037 159
rect 2019 89 2025 95
rect 3967 89 3973 95
rect 85 77 91 83
rect 2019 77 2025 83
<< m5 >>
rect 84 4003 92 4032
rect 84 3997 85 4003
rect 91 3997 92 4003
rect 84 3843 92 3997
rect 84 3837 85 3843
rect 91 3837 92 3843
rect 84 3683 92 3837
rect 84 3677 85 3683
rect 91 3677 92 3683
rect 84 3519 92 3677
rect 84 3513 85 3519
rect 91 3513 92 3519
rect 84 3335 92 3513
rect 84 3329 85 3335
rect 91 3329 92 3335
rect 84 3171 92 3329
rect 84 3165 85 3171
rect 91 3165 92 3171
rect 84 2995 92 3165
rect 84 2989 85 2995
rect 91 2989 92 2995
rect 84 2839 92 2989
rect 84 2833 85 2839
rect 91 2833 92 2839
rect 84 2679 92 2833
rect 84 2673 85 2679
rect 91 2673 92 2679
rect 84 2507 92 2673
rect 84 2501 85 2507
rect 91 2501 92 2507
rect 84 2335 92 2501
rect 84 2329 85 2335
rect 91 2329 92 2335
rect 84 2171 92 2329
rect 84 2165 85 2171
rect 91 2165 92 2171
rect 84 1995 92 2165
rect 84 1989 85 1995
rect 91 1989 92 1995
rect 84 1835 92 1989
rect 84 1829 85 1835
rect 91 1829 92 1835
rect 84 1679 92 1829
rect 84 1673 85 1679
rect 91 1673 92 1679
rect 84 1519 92 1673
rect 84 1513 85 1519
rect 91 1513 92 1519
rect 84 1359 92 1513
rect 84 1353 85 1359
rect 91 1353 92 1359
rect 84 1203 92 1353
rect 84 1197 85 1203
rect 91 1197 92 1203
rect 84 1047 92 1197
rect 84 1041 85 1047
rect 91 1041 92 1047
rect 84 891 92 1041
rect 84 885 85 891
rect 91 885 92 891
rect 84 735 92 885
rect 84 729 85 735
rect 91 729 92 735
rect 84 579 92 729
rect 84 573 85 579
rect 91 573 92 579
rect 84 423 92 573
rect 84 417 85 423
rect 91 417 92 423
rect 84 267 92 417
rect 84 261 85 267
rect 91 261 92 267
rect 84 83 92 261
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 3927 104 4032
rect 96 3921 97 3927
rect 103 3921 104 3927
rect 96 3767 104 3921
rect 96 3761 97 3767
rect 103 3761 104 3767
rect 96 3603 104 3761
rect 96 3597 97 3603
rect 103 3597 104 3603
rect 96 3423 104 3597
rect 96 3417 97 3423
rect 103 3417 104 3423
rect 96 3255 104 3417
rect 96 3249 97 3255
rect 103 3249 104 3255
rect 96 3095 104 3249
rect 96 3089 97 3095
rect 103 3089 104 3095
rect 96 2919 104 3089
rect 96 2913 97 2919
rect 103 2913 104 2919
rect 96 2755 104 2913
rect 96 2749 97 2755
rect 103 2749 104 2755
rect 96 2587 104 2749
rect 96 2581 97 2587
rect 103 2581 104 2587
rect 96 2415 104 2581
rect 96 2409 97 2415
rect 103 2409 104 2415
rect 96 2255 104 2409
rect 96 2249 97 2255
rect 103 2249 104 2255
rect 96 2087 104 2249
rect 96 2081 97 2087
rect 103 2081 104 2087
rect 96 1919 104 2081
rect 96 1913 97 1919
rect 103 1913 104 1919
rect 96 1759 104 1913
rect 96 1753 97 1759
rect 103 1753 104 1759
rect 96 1599 104 1753
rect 96 1593 97 1599
rect 103 1593 104 1599
rect 96 1435 104 1593
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1279 104 1429
rect 96 1273 97 1279
rect 103 1273 104 1279
rect 96 1123 104 1273
rect 96 1117 97 1123
rect 103 1117 104 1123
rect 96 967 104 1117
rect 96 961 97 967
rect 103 961 104 967
rect 96 815 104 961
rect 96 809 97 815
rect 103 809 104 815
rect 96 659 104 809
rect 96 653 97 659
rect 103 653 104 659
rect 96 503 104 653
rect 96 497 97 503
rect 103 497 104 503
rect 96 347 104 497
rect 96 341 97 347
rect 103 341 104 347
rect 96 159 104 341
rect 96 153 97 159
rect 103 153 104 159
rect 96 72 104 153
rect 2018 4023 2026 4032
rect 2018 4017 2019 4023
rect 2025 4017 2026 4023
rect 2018 4003 2026 4017
rect 2018 3997 2019 4003
rect 2025 3997 2026 4003
rect 2018 3871 2026 3997
rect 2018 3865 2019 3871
rect 2025 3865 2026 3871
rect 2018 3843 2026 3865
rect 2018 3837 2019 3843
rect 2025 3837 2026 3843
rect 2018 3691 2026 3837
rect 2018 3685 2019 3691
rect 2025 3685 2026 3691
rect 2018 3683 2026 3685
rect 2018 3677 2019 3683
rect 2025 3677 2026 3683
rect 2018 3531 2026 3677
rect 2018 3525 2019 3531
rect 2025 3525 2026 3531
rect 2018 3519 2026 3525
rect 2018 3513 2019 3519
rect 2025 3513 2026 3519
rect 2018 3367 2026 3513
rect 2018 3361 2019 3367
rect 2025 3361 2026 3367
rect 2018 3335 2026 3361
rect 2018 3329 2019 3335
rect 2025 3329 2026 3335
rect 2018 3199 2026 3329
rect 2018 3193 2019 3199
rect 2025 3193 2026 3199
rect 2018 3171 2026 3193
rect 2018 3165 2019 3171
rect 2025 3165 2026 3171
rect 2018 3035 2026 3165
rect 2018 3029 2019 3035
rect 2025 3029 2026 3035
rect 2018 2995 2026 3029
rect 2018 2989 2019 2995
rect 2025 2989 2026 2995
rect 2018 2871 2026 2989
rect 2018 2865 2019 2871
rect 2025 2865 2026 2871
rect 2018 2839 2026 2865
rect 2018 2833 2019 2839
rect 2025 2833 2026 2839
rect 2018 2699 2026 2833
rect 2018 2693 2019 2699
rect 2025 2693 2026 2699
rect 2018 2679 2026 2693
rect 2018 2673 2019 2679
rect 2025 2673 2026 2679
rect 2018 2535 2026 2673
rect 2018 2529 2019 2535
rect 2025 2529 2026 2535
rect 2018 2507 2026 2529
rect 2018 2501 2019 2507
rect 2025 2501 2026 2507
rect 2018 2367 2026 2501
rect 2018 2361 2019 2367
rect 2025 2361 2026 2367
rect 2018 2335 2026 2361
rect 2018 2329 2019 2335
rect 2025 2329 2026 2335
rect 2018 2215 2026 2329
rect 2018 2209 2019 2215
rect 2025 2209 2026 2215
rect 2018 2171 2026 2209
rect 2018 2165 2019 2171
rect 2025 2165 2026 2171
rect 2018 2039 2026 2165
rect 2018 2033 2019 2039
rect 2025 2033 2026 2039
rect 2018 1995 2026 2033
rect 2018 1989 2019 1995
rect 2025 1989 2026 1995
rect 2018 1875 2026 1989
rect 2018 1869 2019 1875
rect 2025 1869 2026 1875
rect 2018 1835 2026 1869
rect 2018 1829 2019 1835
rect 2025 1829 2026 1835
rect 2018 1711 2026 1829
rect 2018 1705 2019 1711
rect 2025 1705 2026 1711
rect 2018 1679 2026 1705
rect 2018 1673 2019 1679
rect 2025 1673 2026 1679
rect 2018 1555 2026 1673
rect 2018 1549 2019 1555
rect 2025 1549 2026 1555
rect 2018 1519 2026 1549
rect 2018 1513 2019 1519
rect 2025 1513 2026 1519
rect 2018 1391 2026 1513
rect 2018 1385 2019 1391
rect 2025 1385 2026 1391
rect 2018 1359 2026 1385
rect 2018 1353 2019 1359
rect 2025 1353 2026 1359
rect 2018 1231 2026 1353
rect 2018 1225 2019 1231
rect 2025 1225 2026 1231
rect 2018 1203 2026 1225
rect 2018 1197 2019 1203
rect 2025 1197 2026 1203
rect 2018 1063 2026 1197
rect 2018 1057 2019 1063
rect 2025 1057 2026 1063
rect 2018 1047 2026 1057
rect 2018 1041 2019 1047
rect 2025 1041 2026 1047
rect 2018 903 2026 1041
rect 2018 897 2019 903
rect 2025 897 2026 903
rect 2018 891 2026 897
rect 2018 885 2019 891
rect 2025 885 2026 891
rect 2018 743 2026 885
rect 2018 737 2019 743
rect 2025 737 2026 743
rect 2018 735 2026 737
rect 2018 729 2019 735
rect 2025 729 2026 735
rect 2018 579 2026 729
rect 2018 573 2019 579
rect 2025 573 2026 579
rect 2018 423 2026 573
rect 2018 417 2019 423
rect 2025 417 2026 423
rect 2018 267 2026 417
rect 2018 261 2019 267
rect 2025 261 2026 267
rect 2018 95 2026 261
rect 2018 89 2019 95
rect 2025 89 2026 95
rect 2018 83 2026 89
rect 2018 77 2019 83
rect 2025 77 2026 83
rect 2018 72 2026 77
rect 2030 3947 2038 4032
rect 2030 3941 2031 3947
rect 2037 3941 2038 3947
rect 2030 3927 2038 3941
rect 2030 3921 2031 3927
rect 2037 3921 2038 3927
rect 2030 3779 2038 3921
rect 2030 3773 2031 3779
rect 2037 3773 2038 3779
rect 2030 3767 2038 3773
rect 2030 3761 2031 3767
rect 2037 3761 2038 3767
rect 2030 3611 2038 3761
rect 2030 3605 2031 3611
rect 2037 3605 2038 3611
rect 2030 3603 2038 3605
rect 2030 3597 2031 3603
rect 2037 3597 2038 3603
rect 2030 3455 2038 3597
rect 2030 3449 2031 3455
rect 2037 3449 2038 3455
rect 2030 3423 2038 3449
rect 2030 3417 2031 3423
rect 2037 3417 2038 3423
rect 2030 3287 2038 3417
rect 2030 3281 2031 3287
rect 2037 3281 2038 3287
rect 2030 3255 2038 3281
rect 2030 3249 2031 3255
rect 2037 3249 2038 3255
rect 2030 3119 2038 3249
rect 2030 3113 2031 3119
rect 2037 3113 2038 3119
rect 2030 3095 2038 3113
rect 2030 3089 2031 3095
rect 2037 3089 2038 3095
rect 2030 2955 2038 3089
rect 2030 2949 2031 2955
rect 2037 2949 2038 2955
rect 2030 2919 2038 2949
rect 2030 2913 2031 2919
rect 2037 2913 2038 2919
rect 2030 2795 2038 2913
rect 2030 2789 2031 2795
rect 2037 2789 2038 2795
rect 2030 2755 2038 2789
rect 2030 2749 2031 2755
rect 2037 2749 2038 2755
rect 2030 2615 2038 2749
rect 2030 2609 2031 2615
rect 2037 2609 2038 2615
rect 2030 2587 2038 2609
rect 2030 2581 2031 2587
rect 2037 2581 2038 2587
rect 2030 2447 2038 2581
rect 2030 2441 2031 2447
rect 2037 2441 2038 2447
rect 2030 2415 2038 2441
rect 2030 2409 2031 2415
rect 2037 2409 2038 2415
rect 2030 2291 2038 2409
rect 2030 2285 2031 2291
rect 2037 2285 2038 2291
rect 2030 2255 2038 2285
rect 2030 2249 2031 2255
rect 2037 2249 2038 2255
rect 2030 2115 2038 2249
rect 2030 2109 2031 2115
rect 2037 2109 2038 2115
rect 2030 2087 2038 2109
rect 2030 2081 2031 2087
rect 2037 2081 2038 2087
rect 2030 1951 2038 2081
rect 2030 1945 2031 1951
rect 2037 1945 2038 1951
rect 2030 1919 2038 1945
rect 2030 1913 2031 1919
rect 2037 1913 2038 1919
rect 2030 1795 2038 1913
rect 2030 1789 2031 1795
rect 2037 1789 2038 1795
rect 2030 1759 2038 1789
rect 2030 1753 2031 1759
rect 2037 1753 2038 1759
rect 2030 1631 2038 1753
rect 2030 1625 2031 1631
rect 2037 1625 2038 1631
rect 2030 1599 2038 1625
rect 2030 1593 2031 1599
rect 2037 1593 2038 1599
rect 2030 1467 2038 1593
rect 2030 1461 2031 1467
rect 2037 1461 2038 1467
rect 2030 1435 2038 1461
rect 2030 1429 2031 1435
rect 2037 1429 2038 1435
rect 2030 1311 2038 1429
rect 2030 1305 2031 1311
rect 2037 1305 2038 1311
rect 2030 1279 2038 1305
rect 2030 1273 2031 1279
rect 2037 1273 2038 1279
rect 2030 1151 2038 1273
rect 2030 1145 2031 1151
rect 2037 1145 2038 1151
rect 2030 1123 2038 1145
rect 2030 1117 2031 1123
rect 2037 1117 2038 1123
rect 2030 983 2038 1117
rect 2030 977 2031 983
rect 2037 977 2038 983
rect 2030 967 2038 977
rect 2030 961 2031 967
rect 2037 961 2038 967
rect 2030 823 2038 961
rect 2030 817 2031 823
rect 2037 817 2038 823
rect 2030 815 2038 817
rect 2030 809 2031 815
rect 2037 809 2038 815
rect 2030 659 2038 809
rect 2030 653 2031 659
rect 2037 653 2038 659
rect 2030 503 2038 653
rect 2030 497 2031 503
rect 2037 497 2038 503
rect 2030 347 2038 497
rect 2030 341 2031 347
rect 2037 341 2038 347
rect 2030 171 2038 341
rect 2030 165 2031 171
rect 2037 165 2038 171
rect 2030 159 2038 165
rect 2030 153 2031 159
rect 2037 153 2038 159
rect 2030 72 2038 153
rect 3966 4023 3974 4032
rect 3966 4017 3967 4023
rect 3973 4017 3974 4023
rect 3966 3871 3974 4017
rect 3966 3865 3967 3871
rect 3973 3865 3974 3871
rect 3966 3691 3974 3865
rect 3966 3685 3967 3691
rect 3973 3685 3974 3691
rect 3966 3531 3974 3685
rect 3966 3525 3967 3531
rect 3973 3525 3974 3531
rect 3966 3367 3974 3525
rect 3966 3361 3967 3367
rect 3973 3361 3974 3367
rect 3966 3199 3974 3361
rect 3966 3193 3967 3199
rect 3973 3193 3974 3199
rect 3966 3035 3974 3193
rect 3966 3029 3967 3035
rect 3973 3029 3974 3035
rect 3966 2871 3974 3029
rect 3966 2865 3967 2871
rect 3973 2865 3974 2871
rect 3966 2699 3974 2865
rect 3966 2693 3967 2699
rect 3973 2693 3974 2699
rect 3966 2535 3974 2693
rect 3966 2529 3967 2535
rect 3973 2529 3974 2535
rect 3966 2367 3974 2529
rect 3966 2361 3967 2367
rect 3973 2361 3974 2367
rect 3966 2215 3974 2361
rect 3966 2209 3967 2215
rect 3973 2209 3974 2215
rect 3966 2039 3974 2209
rect 3966 2033 3967 2039
rect 3973 2033 3974 2039
rect 3966 1875 3974 2033
rect 3966 1869 3967 1875
rect 3973 1869 3974 1875
rect 3966 1711 3974 1869
rect 3966 1705 3967 1711
rect 3973 1705 3974 1711
rect 3966 1555 3974 1705
rect 3966 1549 3967 1555
rect 3973 1549 3974 1555
rect 3966 1391 3974 1549
rect 3966 1385 3967 1391
rect 3973 1385 3974 1391
rect 3966 1231 3974 1385
rect 3966 1225 3967 1231
rect 3973 1225 3974 1231
rect 3966 1063 3974 1225
rect 3966 1057 3967 1063
rect 3973 1057 3974 1063
rect 3966 903 3974 1057
rect 3966 897 3967 903
rect 3973 897 3974 903
rect 3966 743 3974 897
rect 3966 737 3967 743
rect 3973 737 3974 743
rect 3966 95 3974 737
rect 3966 89 3967 95
rect 3973 89 3974 95
rect 3966 72 3974 89
rect 3978 3947 3986 4032
rect 3978 3941 3979 3947
rect 3985 3941 3986 3947
rect 3978 3779 3986 3941
rect 3978 3773 3979 3779
rect 3985 3773 3986 3779
rect 3978 3611 3986 3773
rect 3978 3605 3979 3611
rect 3985 3605 3986 3611
rect 3978 3455 3986 3605
rect 3978 3449 3979 3455
rect 3985 3449 3986 3455
rect 3978 3287 3986 3449
rect 3978 3281 3979 3287
rect 3985 3281 3986 3287
rect 3978 3119 3986 3281
rect 3978 3113 3979 3119
rect 3985 3113 3986 3119
rect 3978 2955 3986 3113
rect 3978 2949 3979 2955
rect 3985 2949 3986 2955
rect 3978 2795 3986 2949
rect 3978 2789 3979 2795
rect 3985 2789 3986 2795
rect 3978 2615 3986 2789
rect 3978 2609 3979 2615
rect 3985 2609 3986 2615
rect 3978 2447 3986 2609
rect 3978 2441 3979 2447
rect 3985 2441 3986 2447
rect 3978 2291 3986 2441
rect 3978 2285 3979 2291
rect 3985 2285 3986 2291
rect 3978 2115 3986 2285
rect 3978 2109 3979 2115
rect 3985 2109 3986 2115
rect 3978 1951 3986 2109
rect 3978 1945 3979 1951
rect 3985 1945 3986 1951
rect 3978 1795 3986 1945
rect 3978 1789 3979 1795
rect 3985 1789 3986 1795
rect 3978 1631 3986 1789
rect 3978 1625 3979 1631
rect 3985 1625 3986 1631
rect 3978 1467 3986 1625
rect 3978 1461 3979 1467
rect 3985 1461 3986 1467
rect 3978 1311 3986 1461
rect 3978 1305 3979 1311
rect 3985 1305 3986 1311
rect 3978 1151 3986 1305
rect 3978 1145 3979 1151
rect 3985 1145 3986 1151
rect 3978 983 3986 1145
rect 3978 977 3979 983
rect 3985 977 3986 983
rect 3978 823 3986 977
rect 3978 817 3979 823
rect 3985 817 3986 823
rect 3978 171 3986 817
rect 3978 165 3979 171
rect 3985 165 3986 171
rect 3978 72 3986 165
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__191
timestamp 1731220350
transform 1 0 3936 0 -1 3992
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220350
transform 1 0 2040 0 -1 3992
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220350
transform 1 0 3936 0 1 3896
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220350
transform 1 0 2040 0 1 3896
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220350
transform 1 0 3936 0 -1 3840
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220350
transform 1 0 2040 0 -1 3840
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220350
transform 1 0 3936 0 1 3728
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220350
transform 1 0 2040 0 1 3728
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220350
transform 1 0 3936 0 -1 3660
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220350
transform 1 0 2040 0 -1 3660
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220350
transform 1 0 3936 0 1 3560
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220350
transform 1 0 2040 0 1 3560
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220350
transform 1 0 3936 0 -1 3500
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220350
transform 1 0 2040 0 -1 3500
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220350
transform 1 0 3936 0 1 3404
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220350
transform 1 0 2040 0 1 3404
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220350
transform 1 0 3936 0 -1 3336
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220350
transform 1 0 2040 0 -1 3336
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220350
transform 1 0 3936 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220350
transform 1 0 2040 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220350
transform 1 0 3936 0 -1 3168
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220350
transform 1 0 2040 0 -1 3168
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220350
transform 1 0 3936 0 1 3068
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220350
transform 1 0 2040 0 1 3068
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220350
transform 1 0 3936 0 -1 3004
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220350
transform 1 0 2040 0 -1 3004
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220350
transform 1 0 3936 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220350
transform 1 0 2040 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220350
transform 1 0 3936 0 -1 2840
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220350
transform 1 0 2040 0 -1 2840
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220350
transform 1 0 3936 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220350
transform 1 0 2040 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220350
transform 1 0 3936 0 -1 2668
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220350
transform 1 0 2040 0 -1 2668
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220350
transform 1 0 3936 0 1 2564
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220350
transform 1 0 2040 0 1 2564
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220350
transform 1 0 3936 0 -1 2504
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220350
transform 1 0 2040 0 -1 2504
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220350
transform 1 0 3936 0 1 2396
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220350
transform 1 0 2040 0 1 2396
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220350
transform 1 0 3936 0 -1 2336
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220350
transform 1 0 2040 0 -1 2336
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220350
transform 1 0 3936 0 1 2240
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220350
transform 1 0 2040 0 1 2240
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220350
transform 1 0 3936 0 -1 2184
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220350
transform 1 0 2040 0 -1 2184
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220350
transform 1 0 3936 0 1 2064
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220350
transform 1 0 2040 0 1 2064
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220350
transform 1 0 3936 0 -1 2008
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220350
transform 1 0 2040 0 -1 2008
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220350
transform 1 0 3936 0 1 1900
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220350
transform 1 0 2040 0 1 1900
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220350
transform 1 0 3936 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220350
transform 1 0 2040 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220350
transform 1 0 3936 0 1 1744
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220350
transform 1 0 2040 0 1 1744
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220350
transform 1 0 3936 0 -1 1680
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220350
transform 1 0 2040 0 -1 1680
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220350
transform 1 0 3936 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220350
transform 1 0 2040 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220350
transform 1 0 3936 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220350
transform 1 0 2040 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220350
transform 1 0 3936 0 1 1416
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220350
transform 1 0 2040 0 1 1416
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220350
transform 1 0 3936 0 -1 1360
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220350
transform 1 0 2040 0 -1 1360
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220350
transform 1 0 3936 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220350
transform 1 0 2040 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220350
transform 1 0 3936 0 -1 1200
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220350
transform 1 0 2040 0 -1 1200
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220350
transform 1 0 3936 0 1 1100
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220350
transform 1 0 2040 0 1 1100
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220350
transform 1 0 3936 0 -1 1032
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220350
transform 1 0 2040 0 -1 1032
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220350
transform 1 0 3936 0 1 932
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220350
transform 1 0 2040 0 1 932
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220350
transform 1 0 3936 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220350
transform 1 0 2040 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220350
transform 1 0 3936 0 1 772
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220350
transform 1 0 2040 0 1 772
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220350
transform 1 0 3936 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220350
transform 1 0 2040 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220350
transform 1 0 3936 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220350
transform 1 0 2040 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220350
transform 1 0 3936 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220350
transform 1 0 2040 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220350
transform 1 0 3936 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220350
transform 1 0 2040 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220350
transform 1 0 3936 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220350
transform 1 0 2040 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220350
transform 1 0 3936 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220350
transform 1 0 2040 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220350
transform 1 0 3936 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220350
transform 1 0 2040 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220350
transform 1 0 3936 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220350
transform 1 0 2040 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220350
transform 1 0 2000 0 -1 3972
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220350
transform 1 0 104 0 -1 3972
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220350
transform 1 0 2000 0 1 3876
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220350
transform 1 0 104 0 1 3876
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220350
transform 1 0 2000 0 -1 3812
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220350
transform 1 0 104 0 -1 3812
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220350
transform 1 0 2000 0 1 3716
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220350
transform 1 0 104 0 1 3716
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220350
transform 1 0 2000 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220350
transform 1 0 104 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220350
transform 1 0 2000 0 1 3552
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220350
transform 1 0 104 0 1 3552
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220350
transform 1 0 2000 0 -1 3488
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220350
transform 1 0 104 0 -1 3488
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220350
transform 1 0 2000 0 1 3372
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220350
transform 1 0 104 0 1 3372
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220350
transform 1 0 2000 0 -1 3304
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220350
transform 1 0 104 0 -1 3304
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220350
transform 1 0 2000 0 1 3204
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220350
transform 1 0 104 0 1 3204
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220350
transform 1 0 2000 0 -1 3140
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220350
transform 1 0 104 0 -1 3140
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220350
transform 1 0 2000 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220350
transform 1 0 104 0 1 3044
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220350
transform 1 0 2000 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220350
transform 1 0 104 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220350
transform 1 0 2000 0 1 2868
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220350
transform 1 0 104 0 1 2868
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220350
transform 1 0 2000 0 -1 2808
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220350
transform 1 0 104 0 -1 2808
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220350
transform 1 0 2000 0 1 2704
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220350
transform 1 0 104 0 1 2704
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220350
transform 1 0 2000 0 -1 2648
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220350
transform 1 0 104 0 -1 2648
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220350
transform 1 0 2000 0 1 2536
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220350
transform 1 0 104 0 1 2536
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220350
transform 1 0 2000 0 -1 2476
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220350
transform 1 0 104 0 -1 2476
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220350
transform 1 0 2000 0 1 2364
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220350
transform 1 0 104 0 1 2364
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220350
transform 1 0 2000 0 -1 2304
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220350
transform 1 0 104 0 -1 2304
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220350
transform 1 0 2000 0 1 2204
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220350
transform 1 0 104 0 1 2204
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220350
transform 1 0 2000 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220350
transform 1 0 104 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220350
transform 1 0 2000 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220350
transform 1 0 104 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220350
transform 1 0 2000 0 -1 1964
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220350
transform 1 0 104 0 -1 1964
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220350
transform 1 0 2000 0 1 1868
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220350
transform 1 0 104 0 1 1868
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220350
transform 1 0 2000 0 -1 1804
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220350
transform 1 0 104 0 -1 1804
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220350
transform 1 0 2000 0 1 1708
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220350
transform 1 0 104 0 1 1708
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220350
transform 1 0 2000 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220350
transform 1 0 104 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220350
transform 1 0 2000 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220350
transform 1 0 104 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220350
transform 1 0 2000 0 -1 1488
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220350
transform 1 0 104 0 -1 1488
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220350
transform 1 0 2000 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220350
transform 1 0 104 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220350
transform 1 0 2000 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220350
transform 1 0 104 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220350
transform 1 0 2000 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220350
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220350
transform 1 0 2000 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220350
transform 1 0 104 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220350
transform 1 0 2000 0 1 1072
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220350
transform 1 0 104 0 1 1072
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220350
transform 1 0 2000 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220350
transform 1 0 104 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220350
transform 1 0 2000 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220350
transform 1 0 104 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220350
transform 1 0 2000 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220350
transform 1 0 104 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220350
transform 1 0 2000 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220350
transform 1 0 104 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220350
transform 1 0 2000 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220350
transform 1 0 104 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220350
transform 1 0 2000 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220350
transform 1 0 104 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220350
transform 1 0 2000 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220350
transform 1 0 104 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220350
transform 1 0 2000 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220350
transform 1 0 104 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220350
transform 1 0 2000 0 -1 392
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220350
transform 1 0 104 0 -1 392
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220350
transform 1 0 2000 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220350
transform 1 0 104 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220350
transform 1 0 2000 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220350
transform 1 0 104 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220350
transform 1 0 2000 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220350
transform 1 0 104 0 1 108
box 7 3 12 24
use _0_0cell_0_0gcelem3x0  tst_5999_6
timestamp 1731220350
transform 1 0 3736 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5998_6
timestamp 1731220350
transform 1 0 3832 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5997_6
timestamp 1731220350
transform 1 0 3832 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5996_6
timestamp 1731220350
transform 1 0 3832 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5995_6
timestamp 1731220350
transform 1 0 3800 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5994_6
timestamp 1731220350
transform 1 0 3776 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5993_6
timestamp 1731220350
transform 1 0 3648 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5992_6
timestamp 1731220350
transform 1 0 3680 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5991_6
timestamp 1731220350
transform 1 0 3504 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5990_6
timestamp 1731220350
transform 1 0 3632 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5989_6
timestamp 1731220350
transform 1 0 3520 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5988_6
timestamp 1731220350
transform 1 0 3416 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5987_6
timestamp 1731220350
transform 1 0 3304 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5986_6
timestamp 1731220350
transform 1 0 3184 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5985_6
timestamp 1731220350
transform 1 0 3064 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5984_6
timestamp 1731220350
transform 1 0 2936 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5983_6
timestamp 1731220350
transform 1 0 2792 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5982_6
timestamp 1731220350
transform 1 0 2976 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5981_6
timestamp 1731220350
transform 1 0 3160 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5980_6
timestamp 1731220350
transform 1 0 3336 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5979_6
timestamp 1731220350
transform 1 0 3464 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5978_6
timestamp 1731220350
transform 1 0 3288 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5977_6
timestamp 1731220350
transform 1 0 3112 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5976_6
timestamp 1731220350
transform 1 0 2944 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5975_6
timestamp 1731220350
transform 1 0 3584 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5974_6
timestamp 1731220350
transform 1 0 3392 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5973_6
timestamp 1731220350
transform 1 0 3216 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5972_6
timestamp 1731220350
transform 1 0 3056 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5971_6
timestamp 1731220350
transform 1 0 2920 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5970_6
timestamp 1731220350
transform 1 0 3168 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5969_6
timestamp 1731220350
transform 1 0 3368 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5968_6
timestamp 1731220350
transform 1 0 3584 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5967_6
timestamp 1731220350
transform 1 0 3544 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5966_6
timestamp 1731220350
transform 1 0 3296 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5965_6
timestamp 1731220350
transform 1 0 3064 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5964_6
timestamp 1731220350
transform 1 0 2864 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5963_6
timestamp 1731220350
transform 1 0 2704 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5962_6
timestamp 1731220350
transform 1 0 2616 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5961_6
timestamp 1731220350
transform 1 0 2832 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5960_6
timestamp 1731220350
transform 1 0 3064 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5959_6
timestamp 1731220350
transform 1 0 3568 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5958_6
timestamp 1731220350
transform 1 0 3312 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5957_6
timestamp 1731220350
transform 1 0 3160 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5956_6
timestamp 1731220350
transform 1 0 2976 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5955_6
timestamp 1731220350
transform 1 0 2800 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5954_6
timestamp 1731220350
transform 1 0 3360 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5953_6
timestamp 1731220350
transform 1 0 3568 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5952_6
timestamp 1731220350
transform 1 0 3384 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5951_6
timestamp 1731220350
transform 1 0 3232 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5950_6
timestamp 1731220350
transform 1 0 3072 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5949_6
timestamp 1731220350
transform 1 0 3200 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5948_6
timestamp 1731220350
transform 1 0 3328 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5947_6
timestamp 1731220350
transform 1 0 3456 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5946_6
timestamp 1731220350
transform 1 0 3704 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5945_6
timestamp 1731220350
transform 1 0 3720 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5944_6
timestamp 1731220350
transform 1 0 3584 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5943_6
timestamp 1731220350
transform 1 0 3536 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5942_6
timestamp 1731220350
transform 1 0 3696 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5941_6
timestamp 1731220350
transform 1 0 3776 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5940_6
timestamp 1731220350
transform 1 0 3800 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5939_6
timestamp 1731220350
transform 1 0 3832 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5938_6
timestamp 1731220350
transform 1 0 3832 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5937_6
timestamp 1731220350
transform 1 0 3832 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5936_6
timestamp 1731220350
transform 1 0 3832 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5935_6
timestamp 1731220350
transform 1 0 3832 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5934_6
timestamp 1731220350
transform 1 0 3800 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5933_6
timestamp 1731220350
transform 1 0 3776 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5932_6
timestamp 1731220350
transform 1 0 3672 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5931_6
timestamp 1731220350
transform 1 0 3488 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5930_6
timestamp 1731220350
transform 1 0 3552 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5929_6
timestamp 1731220350
transform 1 0 3408 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5928_6
timestamp 1731220350
transform 1 0 3256 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5927_6
timestamp 1731220350
transform 1 0 3104 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5926_6
timestamp 1731220350
transform 1 0 2912 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5925_6
timestamp 1731220350
transform 1 0 3112 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5924_6
timestamp 1731220350
transform 1 0 3304 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5923_6
timestamp 1731220350
transform 1 0 3552 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5922_6
timestamp 1731220350
transform 1 0 3312 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5921_6
timestamp 1731220350
transform 1 0 3080 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5920_6
timestamp 1731220350
transform 1 0 2864 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5919_6
timestamp 1731220350
transform 1 0 2672 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5918_6
timestamp 1731220350
transform 1 0 2704 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5917_6
timestamp 1731220350
transform 1 0 2880 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5916_6
timestamp 1731220350
transform 1 0 3080 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5915_6
timestamp 1731220350
transform 1 0 3304 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5914_6
timestamp 1731220350
transform 1 0 3536 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5913_6
timestamp 1731220350
transform 1 0 3656 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5912_6
timestamp 1731220350
transform 1 0 3464 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5911_6
timestamp 1731220350
transform 1 0 3280 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5910_6
timestamp 1731220350
transform 1 0 3104 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5909_6
timestamp 1731220350
transform 1 0 2936 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5908_6
timestamp 1731220350
transform 1 0 3104 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5907_6
timestamp 1731220350
transform 1 0 3248 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5906_6
timestamp 1731220350
transform 1 0 3400 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5905_6
timestamp 1731220350
transform 1 0 3704 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5904_6
timestamp 1731220350
transform 1 0 3552 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5903_6
timestamp 1731220350
transform 1 0 3440 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5902_6
timestamp 1731220350
transform 1 0 3304 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5901_6
timestamp 1731220350
transform 1 0 3576 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5900_6
timestamp 1731220350
transform 1 0 3712 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5899_6
timestamp 1731220350
transform 1 0 3584 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5898_6
timestamp 1731220350
transform 1 0 3456 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5897_6
timestamp 1731220350
transform 1 0 3328 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5896_6
timestamp 1731220350
transform 1 0 3200 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5895_6
timestamp 1731220350
transform 1 0 3448 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5894_6
timestamp 1731220350
transform 1 0 3328 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5893_6
timestamp 1731220350
transform 1 0 3208 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5892_6
timestamp 1731220350
transform 1 0 3088 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5891_6
timestamp 1731220350
transform 1 0 2968 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5890_6
timestamp 1731220350
transform 1 0 3480 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5889_6
timestamp 1731220350
transform 1 0 3296 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5888_6
timestamp 1731220350
transform 1 0 3120 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5887_6
timestamp 1731220350
transform 1 0 2960 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5886_6
timestamp 1731220350
transform 1 0 2816 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5885_6
timestamp 1731220350
transform 1 0 2824 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5884_6
timestamp 1731220350
transform 1 0 3016 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5883_6
timestamp 1731220350
transform 1 0 3216 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5882_6
timestamp 1731220350
transform 1 0 3424 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5881_6
timestamp 1731220350
transform 1 0 3448 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5880_6
timestamp 1731220350
transform 1 0 3312 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5879_6
timestamp 1731220350
transform 1 0 3176 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5878_6
timestamp 1731220350
transform 1 0 3032 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5877_6
timestamp 1731220350
transform 1 0 2880 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5876_6
timestamp 1731220350
transform 1 0 3120 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5875_6
timestamp 1731220350
transform 1 0 3352 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5874_6
timestamp 1731220350
transform 1 0 3584 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5873_6
timestamp 1731220350
transform 1 0 3576 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5872_6
timestamp 1731220350
transform 1 0 3704 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5871_6
timestamp 1731220350
transform 1 0 3640 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5870_6
timestamp 1731220350
transform 1 0 3664 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5869_6
timestamp 1731220350
transform 1 0 3720 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5868_6
timestamp 1731220350
transform 1 0 3832 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5867_6
timestamp 1731220350
transform 1 0 3832 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5866_6
timestamp 1731220350
transform 1 0 3832 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5865_6
timestamp 1731220350
transform 1 0 3832 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5864_6
timestamp 1731220350
transform 1 0 3832 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5863_6
timestamp 1731220350
transform 1 0 3832 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5862_6
timestamp 1731220350
transform 1 0 3832 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5861_6
timestamp 1731220350
transform 1 0 3824 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5860_6
timestamp 1731220350
transform 1 0 3520 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5859_6
timestamp 1731220350
transform 1 0 3832 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5858_6
timestamp 1731220350
transform 1 0 3832 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5857_6
timestamp 1731220350
transform 1 0 3736 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5856_6
timestamp 1731220350
transform 1 0 3640 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5855_6
timestamp 1731220350
transform 1 0 3544 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5854_6
timestamp 1731220350
transform 1 0 3448 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5853_6
timestamp 1731220350
transform 1 0 3352 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5852_6
timestamp 1731220350
transform 1 0 3256 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5851_6
timestamp 1731220350
transform 1 0 3160 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5850_6
timestamp 1731220350
transform 1 0 3064 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5849_6
timestamp 1731220350
transform 1 0 2968 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5848_6
timestamp 1731220350
transform 1 0 2872 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5847_6
timestamp 1731220350
transform 1 0 3464 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5846_6
timestamp 1731220350
transform 1 0 3312 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5845_6
timestamp 1731220350
transform 1 0 3168 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5844_6
timestamp 1731220350
transform 1 0 3016 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5843_6
timestamp 1731220350
transform 1 0 2856 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5842_6
timestamp 1731220350
transform 1 0 3264 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5841_6
timestamp 1731220350
transform 1 0 3120 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5840_6
timestamp 1731220350
transform 1 0 2976 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5839_6
timestamp 1731220350
transform 1 0 2832 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5838_6
timestamp 1731220350
transform 1 0 3192 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5837_6
timestamp 1731220350
transform 1 0 3024 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5836_6
timestamp 1731220350
transform 1 0 2864 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5835_6
timestamp 1731220350
transform 1 0 2696 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5834_6
timestamp 1731220350
transform 1 0 2528 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5833_6
timestamp 1731220350
transform 1 0 2672 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5832_6
timestamp 1731220350
transform 1 0 2784 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5831_6
timestamp 1731220350
transform 1 0 2904 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5830_6
timestamp 1731220350
transform 1 0 3024 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5829_6
timestamp 1731220350
transform 1 0 3144 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5828_6
timestamp 1731220350
transform 1 0 3216 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5827_6
timestamp 1731220350
transform 1 0 3088 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5826_6
timestamp 1731220350
transform 1 0 2960 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5825_6
timestamp 1731220350
transform 1 0 2832 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5824_6
timestamp 1731220350
transform 1 0 2712 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5823_6
timestamp 1731220350
transform 1 0 2808 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5822_6
timestamp 1731220350
transform 1 0 2944 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5821_6
timestamp 1731220350
transform 1 0 3080 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5820_6
timestamp 1731220350
transform 1 0 3216 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5819_6
timestamp 1731220350
transform 1 0 3360 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5818_6
timestamp 1731220350
transform 1 0 3528 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5817_6
timestamp 1731220350
transform 1 0 3376 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5816_6
timestamp 1731220350
transform 1 0 3232 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5815_6
timestamp 1731220350
transform 1 0 3088 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5814_6
timestamp 1731220350
transform 1 0 2936 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5813_6
timestamp 1731220350
transform 1 0 2832 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5812_6
timestamp 1731220350
transform 1 0 2720 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5811_6
timestamp 1731220350
transform 1 0 2936 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5810_6
timestamp 1731220350
transform 1 0 3040 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5809_6
timestamp 1731220350
transform 1 0 3136 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5808_6
timestamp 1731220350
transform 1 0 3232 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5807_6
timestamp 1731220350
transform 1 0 3280 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5806_6
timestamp 1731220350
transform 1 0 3472 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5805_6
timestamp 1731220350
transform 1 0 3440 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5804_6
timestamp 1731220350
transform 1 0 3336 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5803_6
timestamp 1731220350
transform 1 0 3544 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5802_6
timestamp 1731220350
transform 1 0 3640 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5801_6
timestamp 1731220350
transform 1 0 3832 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5800_6
timestamp 1731220350
transform 1 0 3736 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5799_6
timestamp 1731220350
transform 1 0 3664 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5798_6
timestamp 1731220350
transform 1 0 3832 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5797_6
timestamp 1731220350
transform 1 0 3832 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5796_6
timestamp 1731220350
transform 1 0 3832 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5795_6
timestamp 1731220350
transform 1 0 3832 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5794_6
timestamp 1731220350
transform 1 0 3808 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5793_6
timestamp 1731220350
transform 1 0 3832 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5792_6
timestamp 1731220350
transform 1 0 3736 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5791_6
timestamp 1731220350
transform 1 0 3616 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5790_6
timestamp 1731220350
transform 1 0 3496 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5789_6
timestamp 1731220350
transform 1 0 3376 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5788_6
timestamp 1731220350
transform 1 0 3472 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5787_6
timestamp 1731220350
transform 1 0 3624 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5786_6
timestamp 1731220350
transform 1 0 3776 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5785_6
timestamp 1731220350
transform 1 0 3744 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5784_6
timestamp 1731220350
transform 1 0 3800 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5783_6
timestamp 1731220350
transform 1 0 3832 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5782_6
timestamp 1731220350
transform 1 0 3832 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5781_6
timestamp 1731220350
transform 1 0 3832 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5780_6
timestamp 1731220350
transform 1 0 3832 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5779_6
timestamp 1731220350
transform 1 0 3720 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5778_6
timestamp 1731220350
transform 1 0 3592 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5777_6
timestamp 1731220350
transform 1 0 3680 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5776_6
timestamp 1731220350
transform 1 0 3664 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5775_6
timestamp 1731220350
transform 1 0 3632 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5774_6
timestamp 1731220350
transform 1 0 3440 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5773_6
timestamp 1731220350
transform 1 0 3248 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5772_6
timestamp 1731220350
transform 1 0 3104 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5771_6
timestamp 1731220350
transform 1 0 3288 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5770_6
timestamp 1731220350
transform 1 0 3472 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5769_6
timestamp 1731220350
transform 1 0 3504 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5768_6
timestamp 1731220350
transform 1 0 3328 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5767_6
timestamp 1731220350
transform 1 0 3152 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5766_6
timestamp 1731220350
transform 1 0 3200 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5765_6
timestamp 1731220350
transform 1 0 3336 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5764_6
timestamp 1731220350
transform 1 0 3464 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5763_6
timestamp 1731220350
transform 1 0 3552 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5762_6
timestamp 1731220350
transform 1 0 3360 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5761_6
timestamp 1731220350
transform 1 0 3168 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5760_6
timestamp 1731220350
transform 1 0 3336 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5759_6
timestamp 1731220350
transform 1 0 3080 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5758_6
timestamp 1731220350
transform 1 0 2832 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5757_6
timestamp 1731220350
transform 1 0 2584 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5756_6
timestamp 1731220350
transform 1 0 2976 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5755_6
timestamp 1731220350
transform 1 0 3056 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5754_6
timestamp 1731220350
transform 1 0 2912 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5753_6
timestamp 1731220350
transform 1 0 2800 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5752_6
timestamp 1731220350
transform 1 0 2976 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5751_6
timestamp 1731220350
transform 1 0 2920 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5750_6
timestamp 1731220350
transform 1 0 3056 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5749_6
timestamp 1731220350
transform 1 0 2864 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5748_6
timestamp 1731220350
transform 1 0 2904 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5747_6
timestamp 1731220350
transform 1 0 3104 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5746_6
timestamp 1731220350
transform 1 0 3328 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5745_6
timestamp 1731220350
transform 1 0 3560 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5744_6
timestamp 1731220350
transform 1 0 3560 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5743_6
timestamp 1731220350
transform 1 0 3376 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5742_6
timestamp 1731220350
transform 1 0 3200 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5741_6
timestamp 1731220350
transform 1 0 3040 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5740_6
timestamp 1731220350
transform 1 0 3320 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5739_6
timestamp 1731220350
transform 1 0 3168 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5738_6
timestamp 1731220350
transform 1 0 3112 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5737_6
timestamp 1731220350
transform 1 0 3248 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5736_6
timestamp 1731220350
transform 1 0 3624 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5735_6
timestamp 1731220350
transform 1 0 3440 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5734_6
timestamp 1731220350
transform 1 0 3256 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5733_6
timestamp 1731220350
transform 1 0 3072 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5732_6
timestamp 1731220350
transform 1 0 3632 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5731_6
timestamp 1731220350
transform 1 0 3424 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5730_6
timestamp 1731220350
transform 1 0 3224 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5729_6
timestamp 1731220350
transform 1 0 3032 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5728_6
timestamp 1731220350
transform 1 0 2848 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5727_6
timestamp 1731220350
transform 1 0 3592 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5726_6
timestamp 1731220350
transform 1 0 3328 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5725_6
timestamp 1731220350
transform 1 0 3080 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5724_6
timestamp 1731220350
transform 1 0 2848 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5723_6
timestamp 1731220350
transform 1 0 3560 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5722_6
timestamp 1731220350
transform 1 0 3272 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5721_6
timestamp 1731220350
transform 1 0 2992 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5720_6
timestamp 1731220350
transform 1 0 2728 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5719_6
timestamp 1731220350
transform 1 0 2480 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5718_6
timestamp 1731220350
transform 1 0 2256 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5717_6
timestamp 1731220350
transform 1 0 3088 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5716_6
timestamp 1731220350
transform 1 0 2880 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5715_6
timestamp 1731220350
transform 1 0 2664 0 -1 2868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5714_6
timestamp 1731220350
transform 1 0 2600 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5713_6
timestamp 1731220350
transform 1 0 2472 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5712_6
timestamp 1731220350
transform 1 0 2336 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5711_6
timestamp 1731220350
transform 1 0 2432 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5710_6
timestamp 1731220350
transform 1 0 2608 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5709_6
timestamp 1731220350
transform 1 0 2776 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5708_6
timestamp 1731220350
transform 1 0 2664 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5707_6
timestamp 1731220350
transform 1 0 2512 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5706_6
timestamp 1731220350
transform 1 0 2360 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5705_6
timestamp 1731220350
transform 1 0 2336 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5704_6
timestamp 1731220350
transform 1 0 2208 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5703_6
timestamp 1731220350
transform 1 0 2088 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5702_6
timestamp 1731220350
transform 1 0 2064 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5701_6
timestamp 1731220350
transform 1 0 2312 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5700_6
timestamp 1731220350
transform 1 0 2184 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5699_6
timestamp 1731220350
transform 1 0 2160 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5698_6
timestamp 1731220350
transform 1 0 2696 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5697_6
timestamp 1731220350
transform 1 0 2552 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5696_6
timestamp 1731220350
transform 1 0 2416 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5695_6
timestamp 1731220350
transform 1 0 2064 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5694_6
timestamp 1731220350
transform 1 0 2160 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5693_6
timestamp 1731220350
transform 1 0 2064 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5692_6
timestamp 1731220350
transform 1 0 1896 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5691_6
timestamp 1731220350
transform 1 0 1792 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5690_6
timestamp 1731220350
transform 1 0 1784 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5689_6
timestamp 1731220350
transform 1 0 1648 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5688_6
timestamp 1731220350
transform 1 0 1896 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5687_6
timestamp 1731220350
transform 1 0 1896 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5686_6
timestamp 1731220350
transform 1 0 1736 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5685_6
timestamp 1731220350
transform 1 0 1576 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5684_6
timestamp 1731220350
transform 1 0 1488 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5683_6
timestamp 1731220350
transform 1 0 1640 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5682_6
timestamp 1731220350
transform 1 0 1792 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5681_6
timestamp 1731220350
transform 1 0 1696 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5680_6
timestamp 1731220350
transform 1 0 1504 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5679_6
timestamp 1731220350
transform 1 0 1320 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5678_6
timestamp 1731220350
transform 1 0 1248 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5677_6
timestamp 1731220350
transform 1 0 1416 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5676_6
timestamp 1731220350
transform 1 0 1592 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5675_6
timestamp 1731220350
transform 1 0 1568 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5674_6
timestamp 1731220350
transform 1 0 1392 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5673_6
timestamp 1731220350
transform 1 0 1216 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5672_6
timestamp 1731220350
transform 1 0 1160 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5671_6
timestamp 1731220350
transform 1 0 1344 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5670_6
timestamp 1731220350
transform 1 0 1528 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5669_6
timestamp 1731220350
transform 1 0 1488 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5668_6
timestamp 1731220350
transform 1 0 1288 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5667_6
timestamp 1731220350
transform 1 0 1096 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5666_6
timestamp 1731220350
transform 1 0 928 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5665_6
timestamp 1731220350
transform 1 0 992 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5664_6
timestamp 1731220350
transform 1 0 840 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5663_6
timestamp 1731220350
transform 1 0 872 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5662_6
timestamp 1731220350
transform 1 0 1040 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5661_6
timestamp 1731220350
transform 1 0 1080 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5660_6
timestamp 1731220350
transform 1 0 912 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5659_6
timestamp 1731220350
transform 1 0 944 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5658_6
timestamp 1731220350
transform 1 0 1136 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5657_6
timestamp 1731220350
transform 1 0 1200 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5656_6
timestamp 1731220350
transform 1 0 1344 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5655_6
timestamp 1731220350
transform 1 0 1272 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5654_6
timestamp 1731220350
transform 1 0 1424 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5653_6
timestamp 1731220350
transform 1 0 1520 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5652_6
timestamp 1731220350
transform 1 0 1384 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5651_6
timestamp 1731220350
transform 1 0 1240 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5650_6
timestamp 1731220350
transform 1 0 1416 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5649_6
timestamp 1731220350
transform 1 0 1288 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5648_6
timestamp 1731220350
transform 1 0 1544 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5647_6
timestamp 1731220350
transform 1 0 1664 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5646_6
timestamp 1731220350
transform 1 0 1560 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5645_6
timestamp 1731220350
transform 1 0 1760 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5644_6
timestamp 1731220350
transform 1 0 1672 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5643_6
timestamp 1731220350
transform 1 0 1504 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5642_6
timestamp 1731220350
transform 1 0 1344 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5641_6
timestamp 1731220350
transform 1 0 1512 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5640_6
timestamp 1731220350
transform 1 0 1376 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5639_6
timestamp 1731220350
transform 1 0 1248 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5638_6
timestamp 1731220350
transform 1 0 1120 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5637_6
timestamp 1731220350
transform 1 0 984 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5636_6
timestamp 1731220350
transform 1 0 840 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5635_6
timestamp 1731220350
transform 1 0 864 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5634_6
timestamp 1731220350
transform 1 0 1024 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5633_6
timestamp 1731220350
transform 1 0 1184 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5632_6
timestamp 1731220350
transform 1 0 1360 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5631_6
timestamp 1731220350
transform 1 0 1168 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5630_6
timestamp 1731220350
transform 1 0 984 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5629_6
timestamp 1731220350
transform 1 0 816 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5628_6
timestamp 1731220350
transform 1 0 1160 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5627_6
timestamp 1731220350
transform 1 0 1024 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5626_6
timestamp 1731220350
transform 1 0 888 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5625_6
timestamp 1731220350
transform 1 0 760 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5624_6
timestamp 1731220350
transform 1 0 808 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5623_6
timestamp 1731220350
transform 1 0 1096 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5622_6
timestamp 1731220350
transform 1 0 952 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5621_6
timestamp 1731220350
transform 1 0 840 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5620_6
timestamp 1731220350
transform 1 0 976 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5619_6
timestamp 1731220350
transform 1 0 1120 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5618_6
timestamp 1731220350
transform 1 0 1064 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5617_6
timestamp 1731220350
transform 1 0 928 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5616_6
timestamp 1731220350
transform 1 0 800 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5615_6
timestamp 1731220350
transform 1 0 680 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5614_6
timestamp 1731220350
transform 1 0 568 0 1 2508
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5613_6
timestamp 1731220350
transform 1 0 712 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5612_6
timestamp 1731220350
transform 1 0 600 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5611_6
timestamp 1731220350
transform 1 0 496 0 -1 2504
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5610_6
timestamp 1731220350
transform 1 0 528 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5609_6
timestamp 1731220350
transform 1 0 664 0 1 2336
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5608_6
timestamp 1731220350
transform 1 0 640 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5607_6
timestamp 1731220350
transform 1 0 528 0 -1 2332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5606_6
timestamp 1731220350
transform 1 0 408 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5605_6
timestamp 1731220350
transform 1 0 528 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5604_6
timestamp 1731220350
transform 1 0 664 0 1 2176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5603_6
timestamp 1731220350
transform 1 0 704 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5602_6
timestamp 1731220350
transform 1 0 544 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5601_6
timestamp 1731220350
transform 1 0 384 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5600_6
timestamp 1731220350
transform 1 0 240 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5599_6
timestamp 1731220350
transform 1 0 128 0 -1 2168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5598_6
timestamp 1731220350
transform 1 0 128 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5597_6
timestamp 1731220350
transform 1 0 240 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5596_6
timestamp 1731220350
transform 1 0 392 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5595_6
timestamp 1731220350
transform 1 0 544 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5594_6
timestamp 1731220350
transform 1 0 696 0 1 2008
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5593_6
timestamp 1731220350
transform 1 0 936 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5592_6
timestamp 1731220350
transform 1 0 744 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5591_6
timestamp 1731220350
transform 1 0 560 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5590_6
timestamp 1731220350
transform 1 0 384 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5589_6
timestamp 1731220350
transform 1 0 224 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5588_6
timestamp 1731220350
transform 1 0 504 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5587_6
timestamp 1731220350
transform 1 0 616 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5586_6
timestamp 1731220350
transform 1 0 736 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5585_6
timestamp 1731220350
transform 1 0 856 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5584_6
timestamp 1731220350
transform 1 0 976 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5583_6
timestamp 1731220350
transform 1 0 1032 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5582_6
timestamp 1731220350
transform 1 0 920 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5581_6
timestamp 1731220350
transform 1 0 808 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5580_6
timestamp 1731220350
transform 1 0 704 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5579_6
timestamp 1731220350
transform 1 0 608 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5578_6
timestamp 1731220350
transform 1 0 960 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5577_6
timestamp 1731220350
transform 1 0 792 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5576_6
timestamp 1731220350
transform 1 0 632 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5575_6
timestamp 1731220350
transform 1 0 488 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5574_6
timestamp 1731220350
transform 1 0 360 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5573_6
timestamp 1731220350
transform 1 0 736 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5572_6
timestamp 1731220350
transform 1 0 560 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5571_6
timestamp 1731220350
transform 1 0 392 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5570_6
timestamp 1731220350
transform 1 0 240 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5569_6
timestamp 1731220350
transform 1 0 128 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5568_6
timestamp 1731220350
transform 1 0 128 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5567_6
timestamp 1731220350
transform 1 0 248 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5566_6
timestamp 1731220350
transform 1 0 416 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5565_6
timestamp 1731220350
transform 1 0 608 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5564_6
timestamp 1731220350
transform 1 0 824 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5563_6
timestamp 1731220350
transform 1 0 768 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5562_6
timestamp 1731220350
transform 1 0 576 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5561_6
timestamp 1731220350
transform 1 0 400 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5560_6
timestamp 1731220350
transform 1 0 232 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5559_6
timestamp 1731220350
transform 1 0 456 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5558_6
timestamp 1731220350
transform 1 0 576 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5557_6
timestamp 1731220350
transform 1 0 704 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5556_6
timestamp 1731220350
transform 1 0 848 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5555_6
timestamp 1731220350
transform 1 0 1000 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5554_6
timestamp 1731220350
transform 1 0 1136 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5553_6
timestamp 1731220350
transform 1 0 1008 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5552_6
timestamp 1731220350
transform 1 0 880 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5551_6
timestamp 1731220350
transform 1 0 760 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5550_6
timestamp 1731220350
transform 1 0 648 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5549_6
timestamp 1731220350
transform 1 0 928 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5548_6
timestamp 1731220350
transform 1 0 792 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5547_6
timestamp 1731220350
transform 1 0 664 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5546_6
timestamp 1731220350
transform 1 0 544 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5545_6
timestamp 1731220350
transform 1 0 432 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5544_6
timestamp 1731220350
transform 1 0 800 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5543_6
timestamp 1731220350
transform 1 0 624 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5542_6
timestamp 1731220350
transform 1 0 456 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5541_6
timestamp 1731220350
transform 1 0 296 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5540_6
timestamp 1731220350
transform 1 0 160 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5539_6
timestamp 1731220350
transform 1 0 688 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5538_6
timestamp 1731220350
transform 1 0 520 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5537_6
timestamp 1731220350
transform 1 0 368 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5536_6
timestamp 1731220350
transform 1 0 232 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5535_6
timestamp 1731220350
transform 1 0 128 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5534_6
timestamp 1731220350
transform 1 0 648 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5533_6
timestamp 1731220350
transform 1 0 464 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5532_6
timestamp 1731220350
transform 1 0 280 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5531_6
timestamp 1731220350
transform 1 0 128 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5530_6
timestamp 1731220350
transform 1 0 128 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5529_6
timestamp 1731220350
transform 1 0 288 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5528_6
timestamp 1731220350
transform 1 0 464 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5527_6
timestamp 1731220350
transform 1 0 312 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5526_6
timestamp 1731220350
transform 1 0 152 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5525_6
timestamp 1731220350
transform 1 0 216 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5524_6
timestamp 1731220350
transform 1 0 376 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5523_6
timestamp 1731220350
transform 1 0 304 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5522_6
timestamp 1731220350
transform 1 0 632 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5521_6
timestamp 1731220350
transform 1 0 464 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5520_6
timestamp 1731220350
transform 1 0 440 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5519_6
timestamp 1731220350
transform 1 0 288 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5518_6
timestamp 1731220350
transform 1 0 232 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5517_6
timestamp 1731220350
transform 1 0 408 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5516_6
timestamp 1731220350
transform 1 0 456 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5515_6
timestamp 1731220350
transform 1 0 280 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5514_6
timestamp 1731220350
transform 1 0 128 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5513_6
timestamp 1731220350
transform 1 0 128 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5512_6
timestamp 1731220350
transform 1 0 272 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5511_6
timestamp 1731220350
transform 1 0 136 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5510_6
timestamp 1731220350
transform 1 0 312 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5509_6
timestamp 1731220350
transform 1 0 552 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5508_6
timestamp 1731220350
transform 1 0 384 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5507_6
timestamp 1731220350
transform 1 0 216 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5506_6
timestamp 1731220350
transform 1 0 144 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5505_6
timestamp 1731220350
transform 1 0 240 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5504_6
timestamp 1731220350
transform 1 0 336 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5503_6
timestamp 1731220350
transform 1 0 432 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5502_6
timestamp 1731220350
transform 1 0 528 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5501_6
timestamp 1731220350
transform 1 0 624 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5500_6
timestamp 1731220350
transform 1 0 720 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5499_6
timestamp 1731220350
transform 1 0 816 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5498_6
timestamp 1731220350
transform 1 0 896 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5497_6
timestamp 1731220350
transform 1 0 728 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5496_6
timestamp 1731220350
transform 1 0 624 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5495_6
timestamp 1731220350
transform 1 0 472 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5494_6
timestamp 1731220350
transform 1 0 768 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5493_6
timestamp 1731220350
transform 1 0 712 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5492_6
timestamp 1731220350
transform 1 0 576 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5491_6
timestamp 1731220350
transform 1 0 432 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5490_6
timestamp 1731220350
transform 1 0 632 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5489_6
timestamp 1731220350
transform 1 0 800 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5488_6
timestamp 1731220350
transform 1 0 984 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5487_6
timestamp 1731220350
transform 1 0 792 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5486_6
timestamp 1731220350
transform 1 0 600 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5485_6
timestamp 1731220350
transform 1 0 608 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5484_6
timestamp 1731220350
transform 1 0 776 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5483_6
timestamp 1731220350
transform 1 0 944 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5482_6
timestamp 1731220350
transform 1 0 968 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5481_6
timestamp 1731220350
transform 1 0 800 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5480_6
timestamp 1731220350
transform 1 0 808 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5479_6
timestamp 1731220350
transform 1 0 672 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5478_6
timestamp 1731220350
transform 1 0 528 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5477_6
timestamp 1731220350
transform 1 0 464 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5476_6
timestamp 1731220350
transform 1 0 608 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5475_6
timestamp 1731220350
transform 1 0 744 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5474_6
timestamp 1731220350
transform 1 0 632 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5473_6
timestamp 1731220350
transform 1 0 792 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5472_6
timestamp 1731220350
transform 1 0 944 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5471_6
timestamp 1731220350
transform 1 0 1008 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5470_6
timestamp 1731220350
transform 1 0 832 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5469_6
timestamp 1731220350
transform 1 0 856 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5468_6
timestamp 1731220350
transform 1 0 1032 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5467_6
timestamp 1731220350
transform 1 0 1208 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5466_6
timestamp 1731220350
transform 1 0 1152 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5465_6
timestamp 1731220350
transform 1 0 976 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5464_6
timestamp 1731220350
transform 1 0 1072 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5463_6
timestamp 1731220350
transform 1 0 1224 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5462_6
timestamp 1731220350
transform 1 0 1384 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5461_6
timestamp 1731220350
transform 1 0 1408 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5460_6
timestamp 1731220350
transform 1 0 1272 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5459_6
timestamp 1731220350
transform 1 0 1160 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5458_6
timestamp 1731220350
transform 1 0 1328 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5457_6
timestamp 1731220350
transform 1 0 1504 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5456_6
timestamp 1731220350
transform 1 0 1344 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5455_6
timestamp 1731220350
transform 1 0 1152 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5454_6
timestamp 1731220350
transform 1 0 960 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5453_6
timestamp 1731220350
transform 1 0 1056 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5452_6
timestamp 1731220350
transform 1 0 1304 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5451_6
timestamp 1731220350
transform 1 0 1336 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5450_6
timestamp 1731220350
transform 1 0 1128 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5449_6
timestamp 1731220350
transform 1 0 928 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5448_6
timestamp 1731220350
transform 1 0 1136 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5447_6
timestamp 1731220350
transform 1 0 1320 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5446_6
timestamp 1731220350
transform 1 0 1392 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5445_6
timestamp 1731220350
transform 1 0 1272 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5444_6
timestamp 1731220350
transform 1 0 1152 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5443_6
timestamp 1731220350
transform 1 0 1096 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5442_6
timestamp 1731220350
transform 1 0 1216 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5441_6
timestamp 1731220350
transform 1 0 1328 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5440_6
timestamp 1731220350
transform 1 0 1328 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5439_6
timestamp 1731220350
transform 1 0 1128 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5438_6
timestamp 1731220350
transform 1 0 1536 0 -1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5437_6
timestamp 1731220350
transform 1 0 1448 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5436_6
timestamp 1731220350
transform 1 0 1568 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5435_6
timestamp 1731220350
transform 1 0 1688 0 1 1840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5434_6
timestamp 1731220350
transform 1 0 1632 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5433_6
timestamp 1731220350
transform 1 0 1512 0 -1 1832
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5432_6
timestamp 1731220350
transform 1 0 1504 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5431_6
timestamp 1731220350
transform 1 0 1696 0 1 1680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5430_6
timestamp 1731220350
transform 1 0 1760 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5429_6
timestamp 1731220350
transform 1 0 1544 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5428_6
timestamp 1731220350
transform 1 0 1560 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5427_6
timestamp 1731220350
transform 1 0 1824 0 1 1520
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5426_6
timestamp 1731220350
transform 1 0 1728 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5425_6
timestamp 1731220350
transform 1 0 1536 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5424_6
timestamp 1731220350
transform 1 0 1896 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5423_6
timestamp 1731220350
transform 1 0 1864 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5422_6
timestamp 1731220350
transform 1 0 1680 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5421_6
timestamp 1731220350
transform 1 0 1840 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5420_6
timestamp 1731220350
transform 1 0 1696 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5419_6
timestamp 1731220350
transform 1 0 1552 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5418_6
timestamp 1731220350
transform 1 0 1544 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5417_6
timestamp 1731220350
transform 1 0 1712 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5416_6
timestamp 1731220350
transform 1 0 1688 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5415_6
timestamp 1731220350
transform 1 0 1504 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5414_6
timestamp 1731220350
transform 1 0 1328 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5413_6
timestamp 1731220350
transform 1 0 1560 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5412_6
timestamp 1731220350
transform 1 0 1384 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5411_6
timestamp 1731220350
transform 1 0 1376 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5410_6
timestamp 1731220350
transform 1 0 1192 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5409_6
timestamp 1731220350
transform 1 0 1560 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5408_6
timestamp 1731220350
transform 1 0 1488 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5407_6
timestamp 1731220350
transform 1 0 1352 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5406_6
timestamp 1731220350
transform 1 0 1216 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5405_6
timestamp 1731220350
transform 1 0 1080 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5404_6
timestamp 1731220350
transform 1 0 1344 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5403_6
timestamp 1731220350
transform 1 0 1224 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5402_6
timestamp 1731220350
transform 1 0 1104 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5401_6
timestamp 1731220350
transform 1 0 992 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5400_6
timestamp 1731220350
transform 1 0 872 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5399_6
timestamp 1731220350
transform 1 0 944 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5398_6
timestamp 1731220350
transform 1 0 1072 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5397_6
timestamp 1731220350
transform 1 0 1192 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5396_6
timestamp 1731220350
transform 1 0 1448 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5395_6
timestamp 1731220350
transform 1 0 1320 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5394_6
timestamp 1731220350
transform 1 0 1288 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5393_6
timestamp 1731220350
transform 1 0 1128 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5392_6
timestamp 1731220350
transform 1 0 1760 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5391_6
timestamp 1731220350
transform 1 0 1600 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5390_6
timestamp 1731220350
transform 1 0 1448 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5389_6
timestamp 1731220350
transform 1 0 1392 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5388_6
timestamp 1731220350
transform 1 0 1256 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5387_6
timestamp 1731220350
transform 1 0 1104 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5386_6
timestamp 1731220350
transform 1 0 1528 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5385_6
timestamp 1731220350
transform 1 0 1656 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5384_6
timestamp 1731220350
transform 1 0 1856 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5383_6
timestamp 1731220350
transform 1 0 1680 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5382_6
timestamp 1731220350
transform 1 0 1512 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5381_6
timestamp 1731220350
transform 1 0 1344 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5380_6
timestamp 1731220350
transform 1 0 1168 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5379_6
timestamp 1731220350
transform 1 0 1560 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5378_6
timestamp 1731220350
transform 1 0 1408 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5377_6
timestamp 1731220350
transform 1 0 1264 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5376_6
timestamp 1731220350
transform 1 0 1112 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5375_6
timestamp 1731220350
transform 1 0 960 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5374_6
timestamp 1731220350
transform 1 0 1320 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5373_6
timestamp 1731220350
transform 1 0 1200 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5372_6
timestamp 1731220350
transform 1 0 1080 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5371_6
timestamp 1731220350
transform 1 0 960 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5370_6
timestamp 1731220350
transform 1 0 840 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5369_6
timestamp 1731220350
transform 1 0 896 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5368_6
timestamp 1731220350
transform 1 0 1024 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5367_6
timestamp 1731220350
transform 1 0 1144 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5366_6
timestamp 1731220350
transform 1 0 1264 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5365_6
timestamp 1731220350
transform 1 0 1384 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5364_6
timestamp 1731220350
transform 1 0 1656 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5363_6
timestamp 1731220350
transform 1 0 1504 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5362_6
timestamp 1731220350
transform 1 0 1352 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5361_6
timestamp 1731220350
transform 1 0 1208 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5360_6
timestamp 1731220350
transform 1 0 1056 0 -1 264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5359_6
timestamp 1731220350
transform 1 0 1008 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5358_6
timestamp 1731220350
transform 1 0 912 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5357_6
timestamp 1731220350
transform 1 0 1104 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5356_6
timestamp 1731220350
transform 1 0 1200 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5355_6
timestamp 1731220350
transform 1 0 1296 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5354_6
timestamp 1731220350
transform 1 0 1400 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5353_6
timestamp 1731220350
transform 1 0 1504 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5352_6
timestamp 1731220350
transform 1 0 1608 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5351_6
timestamp 1731220350
transform 1 0 1704 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5350_6
timestamp 1731220350
transform 1 0 1800 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5349_6
timestamp 1731220350
transform 1 0 1896 0 1 80
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5348_6
timestamp 1731220350
transform 1 0 2064 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5347_6
timestamp 1731220350
transform 1 0 2184 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5346_6
timestamp 1731220350
transform 1 0 2640 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5345_6
timestamp 1731220350
transform 1 0 2488 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5344_6
timestamp 1731220350
transform 1 0 2336 0 1 92
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5343_6
timestamp 1731220350
transform 1 0 2208 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5342_6
timestamp 1731220350
transform 1 0 2064 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5341_6
timestamp 1731220350
transform 1 0 2784 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5340_6
timestamp 1731220350
transform 1 0 2584 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5339_6
timestamp 1731220350
transform 1 0 2392 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5338_6
timestamp 1731220350
transform 1 0 2320 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5337_6
timestamp 1731220350
transform 1 0 2184 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5336_6
timestamp 1731220350
transform 1 0 2464 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5335_6
timestamp 1731220350
transform 1 0 2776 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5334_6
timestamp 1731220350
transform 1 0 2616 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5333_6
timestamp 1731220350
transform 1 0 2520 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5332_6
timestamp 1731220350
transform 1 0 2424 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5331_6
timestamp 1731220350
transform 1 0 2616 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5330_6
timestamp 1731220350
transform 1 0 2712 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5329_6
timestamp 1731220350
transform 1 0 2808 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5328_6
timestamp 1731220350
transform 1 0 2992 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5327_6
timestamp 1731220350
transform 1 0 2840 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5326_6
timestamp 1731220350
transform 1 0 2720 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5325_6
timestamp 1731220350
transform 1 0 2616 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5324_6
timestamp 1731220350
transform 1 0 2520 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5323_6
timestamp 1731220350
transform 1 0 2424 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5322_6
timestamp 1731220350
transform 1 0 2576 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5321_6
timestamp 1731220350
transform 1 0 2472 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5320_6
timestamp 1731220350
transform 1 0 2376 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5319_6
timestamp 1731220350
transform 1 0 2280 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5318_6
timestamp 1731220350
transform 1 0 2184 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5317_6
timestamp 1731220350
transform 1 0 2416 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5316_6
timestamp 1731220350
transform 1 0 2232 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5315_6
timestamp 1731220350
transform 1 0 2064 0 1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5314_6
timestamp 1731220350
transform 1 0 1896 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5313_6
timestamp 1731220350
transform 1 0 1784 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5312_6
timestamp 1731220350
transform 1 0 1896 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5311_6
timestamp 1731220350
transform 1 0 2064 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5310_6
timestamp 1731220350
transform 1 0 2176 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5309_6
timestamp 1731220350
transform 1 0 2328 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5308_6
timestamp 1731220350
transform 1 0 2480 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5307_6
timestamp 1731220350
transform 1 0 2632 0 -1 740
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5306_6
timestamp 1731220350
transform 1 0 2608 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5305_6
timestamp 1731220350
transform 1 0 2464 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5304_6
timestamp 1731220350
transform 1 0 2328 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5303_6
timestamp 1731220350
transform 1 0 2760 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5302_6
timestamp 1731220350
transform 1 0 2912 0 1 744
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5301_6
timestamp 1731220350
transform 1 0 3072 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5300_6
timestamp 1731220350
transform 1 0 2936 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5299_6
timestamp 1731220350
transform 1 0 2800 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5298_6
timestamp 1731220350
transform 1 0 2672 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5297_6
timestamp 1731220350
transform 1 0 2552 0 -1 900
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5296_6
timestamp 1731220350
transform 1 0 2944 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5295_6
timestamp 1731220350
transform 1 0 2776 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5294_6
timestamp 1731220350
transform 1 0 2608 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5293_6
timestamp 1731220350
transform 1 0 2448 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5292_6
timestamp 1731220350
transform 1 0 2296 0 1 904
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5291_6
timestamp 1731220350
transform 1 0 2696 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5290_6
timestamp 1731220350
transform 1 0 2480 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5289_6
timestamp 1731220350
transform 1 0 2256 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5288_6
timestamp 1731220350
transform 1 0 2064 0 -1 1060
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5287_6
timestamp 1731220350
transform 1 0 1896 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5286_6
timestamp 1731220350
transform 1 0 1736 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5285_6
timestamp 1731220350
transform 1 0 2064 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5284_6
timestamp 1731220350
transform 1 0 2504 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5283_6
timestamp 1731220350
transform 1 0 2344 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5282_6
timestamp 1731220350
transform 1 0 2192 0 1 1072
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5281_6
timestamp 1731220350
transform 1 0 2176 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5280_6
timestamp 1731220350
transform 1 0 2064 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5279_6
timestamp 1731220350
transform 1 0 2552 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5278_6
timestamp 1731220350
transform 1 0 2424 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5277_6
timestamp 1731220350
transform 1 0 2296 0 -1 1228
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5276_6
timestamp 1731220350
transform 1 0 2240 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5275_6
timestamp 1731220350
transform 1 0 2368 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5274_6
timestamp 1731220350
transform 1 0 2784 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5273_6
timestamp 1731220350
transform 1 0 2640 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5272_6
timestamp 1731220350
transform 1 0 2504 0 1 1232
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5271_6
timestamp 1731220350
transform 1 0 2392 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5270_6
timestamp 1731220350
transform 1 0 2528 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5269_6
timestamp 1731220350
transform 1 0 2960 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5268_6
timestamp 1731220350
transform 1 0 2816 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5267_6
timestamp 1731220350
transform 1 0 2672 0 -1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5266_6
timestamp 1731220350
transform 1 0 2624 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5265_6
timestamp 1731220350
transform 1 0 2512 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5264_6
timestamp 1731220350
transform 1 0 2752 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5263_6
timestamp 1731220350
transform 1 0 2888 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5262_6
timestamp 1731220350
transform 1 0 3024 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5261_6
timestamp 1731220350
transform 1 0 3168 0 1 1388
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5260_6
timestamp 1731220350
transform 1 0 3064 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5259_6
timestamp 1731220350
transform 1 0 2928 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5258_6
timestamp 1731220350
transform 1 0 2792 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5257_6
timestamp 1731220350
transform 1 0 2664 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5256_6
timestamp 1731220350
transform 1 0 2536 0 -1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5255_6
timestamp 1731220350
transform 1 0 2848 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5254_6
timestamp 1731220350
transform 1 0 2728 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5253_6
timestamp 1731220350
transform 1 0 2608 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5252_6
timestamp 1731220350
transform 1 0 2496 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5251_6
timestamp 1731220350
transform 1 0 2384 0 1 1552
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5250_6
timestamp 1731220350
transform 1 0 2680 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5249_6
timestamp 1731220350
transform 1 0 2552 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5248_6
timestamp 1731220350
transform 1 0 2432 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5247_6
timestamp 1731220350
transform 1 0 2320 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5246_6
timestamp 1731220350
transform 1 0 2216 0 -1 1708
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5245_6
timestamp 1731220350
transform 1 0 2648 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5244_6
timestamp 1731220350
transform 1 0 2480 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5243_6
timestamp 1731220350
transform 1 0 2320 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5242_6
timestamp 1731220350
transform 1 0 2176 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5241_6
timestamp 1731220350
transform 1 0 2064 0 1 1716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5240_6
timestamp 1731220350
transform 1 0 2064 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5239_6
timestamp 1731220350
transform 1 0 2192 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5238_6
timestamp 1731220350
transform 1 0 2712 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5237_6
timestamp 1731220350
transform 1 0 2536 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5236_6
timestamp 1731220350
transform 1 0 2360 0 -1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5235_6
timestamp 1731220350
transform 1 0 2232 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5234_6
timestamp 1731220350
transform 1 0 2064 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5233_6
timestamp 1731220350
transform 1 0 2888 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5232_6
timestamp 1731220350
transform 1 0 2664 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5231_6
timestamp 1731220350
transform 1 0 2440 0 1 1872
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5230_6
timestamp 1731220350
transform 1 0 2392 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5229_6
timestamp 1731220350
transform 1 0 2184 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5228_6
timestamp 1731220350
transform 1 0 2640 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5227_6
timestamp 1731220350
transform 1 0 3208 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5226_6
timestamp 1731220350
transform 1 0 2912 0 -1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5225_6
timestamp 1731220350
transform 1 0 2776 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5224_6
timestamp 1731220350
transform 1 0 2584 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5223_6
timestamp 1731220350
transform 1 0 2488 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5222_6
timestamp 1731220350
transform 1 0 2392 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5221_6
timestamp 1731220350
transform 1 0 2680 0 1 2036
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5220_6
timestamp 1731220350
transform 1 0 2680 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5219_6
timestamp 1731220350
transform 1 0 2496 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5218_6
timestamp 1731220350
transform 1 0 2288 0 -1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5217_6
timestamp 1731220350
transform 1 0 2280 0 1 2212
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5216_6
timestamp 1731220350
transform 1 0 2352 0 -1 2364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5215_6
timestamp 1731220350
transform 1 0 2432 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5214_6
timestamp 1731220350
transform 1 0 2552 0 1 2368
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5213_6
timestamp 1731220350
transform 1 0 2592 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5212_6
timestamp 1731220350
transform 1 0 2464 0 -1 2532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5211_6
timestamp 1731220350
transform 1 0 2208 0 1 2536
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5210_6
timestamp 1731220350
transform 1 0 2256 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5209_6
timestamp 1731220350
transform 1 0 2088 0 -1 2696
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5208_6
timestamp 1731220350
transform 1 0 2192 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5207_6
timestamp 1731220350
transform 1 0 2064 0 1 2716
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5206_6
timestamp 1731220350
transform 1 0 1896 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5205_6
timestamp 1731220350
transform 1 0 1744 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5204_6
timestamp 1731220350
transform 1 0 1896 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5203_6
timestamp 1731220350
transform 1 0 1720 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5202_6
timestamp 1731220350
transform 1 0 1704 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5201_6
timestamp 1731220350
transform 1 0 1896 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5200_6
timestamp 1731220350
transform 1 0 2064 0 1 2876
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5199_6
timestamp 1731220350
transform 1 0 2064 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5198_6
timestamp 1731220350
transform 1 0 2176 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5197_6
timestamp 1731220350
transform 1 0 2648 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5196_6
timestamp 1731220350
transform 1 0 2472 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5195_6
timestamp 1731220350
transform 1 0 2320 0 -1 3032
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5194_6
timestamp 1731220350
transform 1 0 2216 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5193_6
timestamp 1731220350
transform 1 0 2072 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5192_6
timestamp 1731220350
transform 1 0 2680 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5191_6
timestamp 1731220350
transform 1 0 2520 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5190_6
timestamp 1731220350
transform 1 0 2368 0 1 3040
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5189_6
timestamp 1731220350
transform 1 0 2240 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5188_6
timestamp 1731220350
transform 1 0 2392 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5187_6
timestamp 1731220350
transform 1 0 2896 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5186_6
timestamp 1731220350
transform 1 0 2720 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5185_6
timestamp 1731220350
transform 1 0 2552 0 -1 3196
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5184_6
timestamp 1731220350
transform 1 0 2544 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5183_6
timestamp 1731220350
transform 1 0 2408 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5182_6
timestamp 1731220350
transform 1 0 2968 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5181_6
timestamp 1731220350
transform 1 0 2824 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5180_6
timestamp 1731220350
transform 1 0 2680 0 1 3208
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5179_6
timestamp 1731220350
transform 1 0 2560 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5178_6
timestamp 1731220350
transform 1 0 2712 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5177_6
timestamp 1731220350
transform 1 0 2864 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5176_6
timestamp 1731220350
transform 1 0 3016 0 -1 3364
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5175_6
timestamp 1731220350
transform 1 0 2896 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5174_6
timestamp 1731220350
transform 1 0 2768 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5173_6
timestamp 1731220350
transform 1 0 2656 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5172_6
timestamp 1731220350
transform 1 0 2544 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5171_6
timestamp 1731220350
transform 1 0 2440 0 1 3376
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5170_6
timestamp 1731220350
transform 1 0 2728 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5169_6
timestamp 1731220350
transform 1 0 2576 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5168_6
timestamp 1731220350
transform 1 0 2440 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5167_6
timestamp 1731220350
transform 1 0 2320 0 -1 3528
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5166_6
timestamp 1731220350
transform 1 0 2664 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5165_6
timestamp 1731220350
transform 1 0 2464 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5164_6
timestamp 1731220350
transform 1 0 2272 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5163_6
timestamp 1731220350
transform 1 0 2096 0 1 3532
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5162_6
timestamp 1731220350
transform 1 0 2728 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5161_6
timestamp 1731220350
transform 1 0 2544 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5160_6
timestamp 1731220350
transform 1 0 2360 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5159_6
timestamp 1731220350
transform 1 0 2192 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5158_6
timestamp 1731220350
transform 1 0 2064 0 -1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5157_6
timestamp 1731220350
transform 1 0 2064 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5156_6
timestamp 1731220350
transform 1 0 2176 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5155_6
timestamp 1731220350
transform 1 0 2320 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5154_6
timestamp 1731220350
transform 1 0 2632 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5153_6
timestamp 1731220350
transform 1 0 2472 0 1 3700
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5152_6
timestamp 1731220350
transform 1 0 2368 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5151_6
timestamp 1731220350
transform 1 0 2256 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5150_6
timestamp 1731220350
transform 1 0 2488 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5149_6
timestamp 1731220350
transform 1 0 2624 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5148_6
timestamp 1731220350
transform 1 0 2768 0 -1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5147_6
timestamp 1731220350
transform 1 0 2792 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5146_6
timestamp 1731220350
transform 1 0 2608 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5145_6
timestamp 1731220350
transform 1 0 2432 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5144_6
timestamp 1731220350
transform 1 0 2264 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5143_6
timestamp 1731220350
transform 1 0 2120 0 1 3868
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5142_6
timestamp 1731220350
transform 1 0 2320 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5141_6
timestamp 1731220350
transform 1 0 2064 0 -1 4020
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5140_6
timestamp 1731220350
transform 1 0 1896 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5139_6
timestamp 1731220350
transform 1 0 1784 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5138_6
timestamp 1731220350
transform 1 0 1648 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5137_6
timestamp 1731220350
transform 1 0 1512 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5136_6
timestamp 1731220350
transform 1 0 1376 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5135_6
timestamp 1731220350
transform 1 0 1224 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5134_6
timestamp 1731220350
transform 1 0 1056 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5133_6
timestamp 1731220350
transform 1 0 1280 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5132_6
timestamp 1731220350
transform 1 0 1472 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5131_6
timestamp 1731220350
transform 1 0 1672 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5130_6
timestamp 1731220350
transform 1 0 1624 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5129_6
timestamp 1731220350
transform 1 0 1496 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5128_6
timestamp 1731220350
transform 1 0 1600 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5127_6
timestamp 1731220350
transform 1 0 1472 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5126_6
timestamp 1731220350
transform 1 0 1688 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5125_6
timestamp 1731220350
transform 1 0 1680 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5124_6
timestamp 1731220350
transform 1 0 1768 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5123_6
timestamp 1731220350
transform 1 0 1592 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5122_6
timestamp 1731220350
transform 1 0 1632 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5121_6
timestamp 1731220350
transform 1 0 1808 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5120_6
timestamp 1731220350
transform 1 0 1816 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5119_6
timestamp 1731220350
transform 1 0 1624 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5118_6
timestamp 1731220350
transform 1 0 1792 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5117_6
timestamp 1731220350
transform 1 0 1616 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5116_6
timestamp 1731220350
transform 1 0 1568 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5115_6
timestamp 1731220350
transform 1 0 1728 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5114_6
timestamp 1731220350
transform 1 0 1760 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5113_6
timestamp 1731220350
transform 1 0 1600 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5112_6
timestamp 1731220350
transform 1 0 1448 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5111_6
timestamp 1731220350
transform 1 0 1296 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5110_6
timestamp 1731220350
transform 1 0 1136 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5109_6
timestamp 1731220350
transform 1 0 1096 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5108_6
timestamp 1731220350
transform 1 0 1256 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5107_6
timestamp 1731220350
transform 1 0 1416 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5106_6
timestamp 1731220350
transform 1 0 1440 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5105_6
timestamp 1731220350
transform 1 0 1264 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5104_6
timestamp 1731220350
transform 1 0 1088 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5103_6
timestamp 1731220350
transform 1 0 1048 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5102_6
timestamp 1731220350
transform 1 0 1432 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5101_6
timestamp 1731220350
transform 1 0 1240 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5100_6
timestamp 1731220350
transform 1 0 1120 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_599_6
timestamp 1731220350
transform 1 0 1288 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_598_6
timestamp 1731220350
transform 1 0 1456 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_597_6
timestamp 1731220350
transform 1 0 1416 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_596_6
timestamp 1731220350
transform 1 0 1240 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_595_6
timestamp 1731220350
transform 1 0 1072 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_594_6
timestamp 1731220350
transform 1 0 984 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_593_6
timestamp 1731220350
transform 1 0 1208 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_592_6
timestamp 1731220350
transform 1 0 1440 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_591_6
timestamp 1731220350
transform 1 0 1256 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_590_6
timestamp 1731220350
transform 1 0 1048 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_589_6
timestamp 1731220350
transform 1 0 832 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_588_6
timestamp 1731220350
transform 1 0 1376 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_587_6
timestamp 1731220350
transform 1 0 1160 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_586_6
timestamp 1731220350
transform 1 0 952 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_585_6
timestamp 1731220350
transform 1 0 744 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_584_6
timestamp 1731220350
transform 1 0 1376 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_583_6
timestamp 1731220350
transform 1 0 1256 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_582_6
timestamp 1731220350
transform 1 0 1144 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_581_6
timestamp 1731220350
transform 1 0 1032 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_580_6
timestamp 1731220350
transform 1 0 928 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_579_6
timestamp 1731220350
transform 1 0 824 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_578_6
timestamp 1731220350
transform 1 0 720 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_577_6
timestamp 1731220350
transform 1 0 624 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_576_6
timestamp 1731220350
transform 1 0 528 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_575_6
timestamp 1731220350
transform 1 0 432 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_574_6
timestamp 1731220350
transform 1 0 1088 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_573_6
timestamp 1731220350
transform 1 0 904 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_572_6
timestamp 1731220350
transform 1 0 728 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_571_6
timestamp 1731220350
transform 1 0 560 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_570_6
timestamp 1731220350
transform 1 0 880 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_569_6
timestamp 1731220350
transform 1 0 696 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_568_6
timestamp 1731220350
transform 1 0 504 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_567_6
timestamp 1731220350
transform 1 0 304 0 -1 4000
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_566_6
timestamp 1731220350
transform 1 0 408 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_565_6
timestamp 1731220350
transform 1 0 272 0 1 3848
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_564_6
timestamp 1731220350
transform 1 0 224 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_563_6
timestamp 1731220350
transform 1 0 328 0 -1 3840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_562_6
timestamp 1731220350
transform 1 0 544 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_561_6
timestamp 1731220350
transform 1 0 344 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_560_6
timestamp 1731220350
transform 1 0 152 0 1 3688
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_559_6
timestamp 1731220350
transform 1 0 144 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_558_6
timestamp 1731220350
transform 1 0 376 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_557_6
timestamp 1731220350
transform 1 0 608 0 -1 3680
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_556_6
timestamp 1731220350
transform 1 0 768 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_555_6
timestamp 1731220350
transform 1 0 552 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_554_6
timestamp 1731220350
transform 1 0 352 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_553_6
timestamp 1731220350
transform 1 0 160 0 1 3524
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_552_6
timestamp 1731220350
transform 1 0 288 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_551_6
timestamp 1731220350
transform 1 0 424 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_550_6
timestamp 1731220350
transform 1 0 576 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_549_6
timestamp 1731220350
transform 1 0 736 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_548_6
timestamp 1731220350
transform 1 0 904 0 -1 3516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_547_6
timestamp 1731220350
transform 1 0 952 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_546_6
timestamp 1731220350
transform 1 0 792 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_545_6
timestamp 1731220350
transform 1 0 640 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_544_6
timestamp 1731220350
transform 1 0 488 0 1 3344
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_543_6
timestamp 1731220350
transform 1 0 664 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_542_6
timestamp 1731220350
transform 1 0 856 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_541_6
timestamp 1731220350
transform 1 0 904 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_540_6
timestamp 1731220350
transform 1 0 712 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_539_6
timestamp 1731220350
transform 1 0 512 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_538_6
timestamp 1731220350
transform 1 0 736 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_537_6
timestamp 1731220350
transform 1 0 920 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_536_6
timestamp 1731220350
transform 1 0 968 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_535_6
timestamp 1731220350
transform 1 0 792 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_534_6
timestamp 1731220350
transform 1 0 776 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_533_6
timestamp 1731220350
transform 1 0 648 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_532_6
timestamp 1731220350
transform 1 0 536 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_531_6
timestamp 1731220350
transform 1 0 568 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_530_6
timestamp 1731220350
transform 1 0 696 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_529_6
timestamp 1731220350
transform 1 0 704 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_528_6
timestamp 1731220350
transform 1 0 544 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_527_6
timestamp 1731220350
transform 1 0 568 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_526_6
timestamp 1731220350
transform 1 0 736 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_525_6
timestamp 1731220350
transform 1 0 752 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_524_6
timestamp 1731220350
transform 1 0 552 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_523_6
timestamp 1731220350
transform 1 0 352 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_522_6
timestamp 1731220350
transform 1 0 160 0 -1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_521_6
timestamp 1731220350
transform 1 0 400 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_520_6
timestamp 1731220350
transform 1 0 248 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_519_6
timestamp 1731220350
transform 1 0 128 0 1 2676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_518_6
timestamp 1731220350
transform 1 0 128 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_517_6
timestamp 1731220350
transform 1 0 240 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_516_6
timestamp 1731220350
transform 1 0 392 0 -1 2836
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_515_6
timestamp 1731220350
transform 1 0 440 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_514_6
timestamp 1731220350
transform 1 0 320 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_513_6
timestamp 1731220350
transform 1 0 200 0 1 2840
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_512_6
timestamp 1731220350
transform 1 0 336 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_511_6
timestamp 1731220350
transform 1 0 432 0 -1 2992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_510_6
timestamp 1731220350
transform 1 0 432 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_59_6
timestamp 1731220350
transform 1 0 256 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_58_6
timestamp 1731220350
transform 1 0 608 0 1 3016
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_57_6
timestamp 1731220350
transform 1 0 536 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_56_6
timestamp 1731220350
transform 1 0 336 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_55_6
timestamp 1731220350
transform 1 0 136 0 -1 3168
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_54_6
timestamp 1731220350
transform 1 0 128 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_53_6
timestamp 1731220350
transform 1 0 312 0 1 3176
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_52_6
timestamp 1731220350
transform 1 0 472 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_51_6
timestamp 1731220350
transform 1 0 288 0 -1 3332
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_50_6
timestamp 1731220350
transform 1 0 128 0 -1 3332
box 8 5 92 72
<< end >>
