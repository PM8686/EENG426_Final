magic
tech sky130l
timestamp 1730743878
<< m2c >>
rect 111 757 115 761
rect 151 756 155 760
rect 191 756 195 760
rect 231 756 235 760
rect 271 756 275 760
rect 280 755 284 759
rect 311 756 315 760
rect 351 756 355 760
rect 391 756 395 760
rect 431 756 435 760
rect 687 757 691 761
rect 111 739 115 743
rect 687 739 691 743
rect 144 735 148 739
rect 160 735 164 739
rect 200 735 204 739
rect 224 735 228 739
rect 240 735 244 739
rect 304 735 308 739
rect 320 735 324 739
rect 360 735 364 739
rect 400 735 404 739
rect 440 735 444 739
rect 184 731 188 735
rect 264 731 268 735
rect 344 731 348 735
rect 384 731 388 735
rect 144 723 148 727
rect 184 719 188 723
rect 224 719 228 723
rect 264 719 268 723
rect 304 719 308 723
rect 344 719 348 723
rect 111 713 115 717
rect 160 715 164 719
rect 200 715 204 719
rect 240 715 244 719
rect 280 715 284 719
rect 320 715 324 719
rect 687 713 691 717
rect 360 703 364 707
rect 111 695 115 699
rect 151 696 155 700
rect 191 696 195 700
rect 231 696 235 700
rect 271 696 275 700
rect 311 696 315 700
rect 351 696 355 700
rect 687 695 691 699
rect 111 645 115 649
rect 151 644 155 648
rect 191 644 195 648
rect 231 644 235 648
rect 271 644 275 648
rect 311 644 315 648
rect 351 644 355 648
rect 687 645 691 649
rect 111 627 115 631
rect 687 627 691 631
rect 144 623 148 627
rect 160 623 164 627
rect 184 623 188 627
rect 200 623 204 627
rect 224 623 228 627
rect 240 623 244 627
rect 264 623 268 627
rect 280 623 284 627
rect 304 623 308 627
rect 320 623 324 627
rect 344 623 348 627
rect 360 623 364 627
rect 144 603 148 607
rect 184 599 188 603
rect 224 599 228 603
rect 264 599 268 603
rect 304 599 308 603
rect 111 593 115 597
rect 160 595 164 599
rect 200 595 204 599
rect 240 595 244 599
rect 280 595 284 599
rect 687 593 691 597
rect 320 583 324 587
rect 111 575 115 579
rect 151 576 155 580
rect 191 576 195 580
rect 231 576 235 580
rect 271 576 275 580
rect 311 576 315 580
rect 687 575 691 579
rect 111 529 115 533
rect 151 528 155 532
rect 191 528 195 532
rect 231 528 235 532
rect 271 528 275 532
rect 311 528 315 532
rect 351 528 355 532
rect 687 529 691 533
rect 111 511 115 515
rect 687 511 691 515
rect 144 507 148 511
rect 160 507 164 511
rect 184 507 188 511
rect 200 507 204 511
rect 224 507 228 511
rect 240 507 244 511
rect 264 507 268 511
rect 280 507 284 511
rect 304 507 308 511
rect 320 507 324 511
rect 344 507 348 511
rect 360 507 364 511
rect 144 491 148 495
rect 184 487 188 491
rect 224 487 228 491
rect 264 487 268 491
rect 304 487 308 491
rect 344 487 348 491
rect 384 487 388 491
rect 111 481 115 485
rect 160 483 164 487
rect 200 483 204 487
rect 240 483 244 487
rect 280 483 284 487
rect 320 483 324 487
rect 360 483 364 487
rect 687 481 691 485
rect 400 471 404 475
rect 111 463 115 467
rect 151 464 155 468
rect 191 464 195 468
rect 231 464 235 468
rect 271 464 275 468
rect 311 464 315 468
rect 351 464 355 468
rect 391 464 395 468
rect 687 463 691 467
rect 111 413 115 417
rect 279 412 283 416
rect 319 412 323 416
rect 359 412 363 416
rect 407 412 411 416
rect 455 412 459 416
rect 503 412 507 416
rect 551 412 555 416
rect 607 412 611 416
rect 655 412 659 416
rect 687 413 691 417
rect 111 395 115 399
rect 687 395 691 399
rect 288 391 292 395
rect 312 391 316 395
rect 328 391 332 395
rect 352 391 356 395
rect 368 391 372 395
rect 400 391 404 395
rect 416 391 420 395
rect 448 391 452 395
rect 464 391 468 395
rect 496 391 500 395
rect 512 391 516 395
rect 560 391 564 395
rect 600 391 604 395
rect 616 391 620 395
rect 648 391 652 395
rect 664 391 668 395
rect 272 387 276 391
rect 544 387 548 391
rect 208 379 212 383
rect 408 379 412 383
rect 648 379 652 383
rect 248 375 252 379
rect 288 375 292 379
rect 328 375 332 379
rect 368 375 372 379
rect 448 375 452 379
rect 488 375 492 379
rect 528 375 532 379
rect 568 375 572 379
rect 608 375 612 379
rect 111 369 115 373
rect 224 371 228 375
rect 464 371 468 375
rect 504 371 508 375
rect 544 371 548 375
rect 687 369 691 373
rect 344 359 348 363
rect 384 359 388 363
rect 424 359 428 363
rect 624 359 628 363
rect 664 359 668 363
rect 111 351 115 355
rect 215 352 219 356
rect 255 352 259 356
rect 264 351 268 355
rect 295 352 299 356
rect 304 351 308 355
rect 335 352 339 356
rect 375 352 379 356
rect 415 352 419 356
rect 455 352 459 356
rect 495 352 499 356
rect 535 352 539 356
rect 575 352 579 356
rect 584 351 588 355
rect 615 352 619 356
rect 655 352 659 356
rect 687 351 691 355
rect 111 305 115 309
rect 223 304 227 308
rect 263 304 267 308
rect 311 304 315 308
rect 367 304 371 308
rect 423 304 427 308
rect 479 304 483 308
rect 488 303 492 307
rect 543 304 547 308
rect 607 304 611 308
rect 655 304 659 308
rect 687 305 691 309
rect 111 287 115 291
rect 687 287 691 291
rect 232 283 236 287
rect 256 283 260 287
rect 272 283 276 287
rect 304 283 308 287
rect 320 283 324 287
rect 360 283 364 287
rect 376 283 380 287
rect 416 283 420 287
rect 432 283 436 287
rect 552 283 556 287
rect 600 283 604 287
rect 616 283 620 287
rect 648 283 652 287
rect 664 283 668 287
rect 216 279 220 283
rect 472 279 476 283
rect 536 279 540 283
rect 280 267 284 271
rect 648 267 652 271
rect 152 263 156 267
rect 216 263 220 267
rect 344 263 348 267
rect 408 263 412 267
rect 472 263 476 267
rect 536 263 540 267
rect 600 263 604 267
rect 111 257 115 261
rect 296 259 300 263
rect 424 259 428 263
rect 488 259 492 263
rect 687 257 691 261
rect 232 247 236 251
rect 360 247 364 251
rect 552 247 556 251
rect 616 247 620 251
rect 664 247 668 251
rect 111 239 115 243
rect 159 240 163 244
rect 168 239 172 243
rect 223 240 227 244
rect 287 240 291 244
rect 351 240 355 244
rect 415 240 419 244
rect 479 240 483 244
rect 543 240 547 244
rect 607 240 611 244
rect 655 240 659 244
rect 687 239 691 243
rect 111 189 115 193
rect 167 188 171 192
rect 215 188 219 192
rect 271 188 275 192
rect 327 188 331 192
rect 383 188 387 192
rect 392 187 396 191
rect 439 188 443 192
rect 495 188 499 192
rect 551 188 555 192
rect 615 188 619 192
rect 655 188 659 192
rect 687 189 691 193
rect 111 171 115 175
rect 687 171 691 175
rect 176 167 180 171
rect 208 167 212 171
rect 224 167 228 171
rect 264 167 268 171
rect 280 167 284 171
rect 320 167 324 171
rect 336 167 340 171
rect 376 167 380 171
rect 448 167 452 171
rect 504 167 508 171
rect 544 167 548 171
rect 560 167 564 171
rect 608 167 612 171
rect 624 167 628 171
rect 648 167 652 171
rect 664 167 668 171
rect 160 163 164 167
rect 431 163 435 167
rect 488 163 492 167
rect 160 151 164 155
rect 648 151 652 155
rect 200 147 204 151
rect 240 147 244 151
rect 280 147 284 151
rect 320 147 324 151
rect 360 147 364 151
rect 400 147 404 151
rect 440 147 444 151
rect 480 147 484 151
rect 528 147 532 151
rect 568 147 572 151
rect 608 147 612 151
rect 111 141 115 145
rect 176 143 180 147
rect 216 143 220 147
rect 256 143 260 147
rect 296 143 300 147
rect 336 143 340 147
rect 376 143 380 147
rect 416 143 420 147
rect 456 143 460 147
rect 496 143 500 147
rect 687 141 691 145
rect 544 131 548 135
rect 624 131 628 135
rect 664 131 668 135
rect 111 123 115 127
rect 167 124 171 128
rect 207 124 211 128
rect 247 124 251 128
rect 287 124 291 128
rect 327 124 331 128
rect 367 124 371 128
rect 407 124 411 128
rect 447 124 451 128
rect 487 124 491 128
rect 535 124 539 128
rect 575 124 579 128
rect 615 124 619 128
rect 655 124 659 128
rect 687 123 691 127
<< m2 >>
rect 222 779 228 780
rect 222 775 223 779
rect 227 778 228 779
rect 278 779 284 780
rect 278 778 279 779
rect 227 776 279 778
rect 227 775 228 776
rect 222 774 228 775
rect 278 775 279 776
rect 283 775 284 779
rect 278 774 284 775
rect 110 761 116 762
rect 686 761 692 762
rect 110 757 111 761
rect 115 757 116 761
rect 110 756 116 757
rect 150 760 156 761
rect 150 756 151 760
rect 155 756 156 760
rect 150 755 156 756
rect 190 760 196 761
rect 190 756 191 760
rect 195 756 196 760
rect 190 755 196 756
rect 230 760 236 761
rect 230 756 231 760
rect 235 756 236 760
rect 230 755 236 756
rect 270 760 276 761
rect 310 760 316 761
rect 270 756 271 760
rect 275 756 276 760
rect 270 755 276 756
rect 278 759 285 760
rect 278 755 279 759
rect 284 755 285 759
rect 310 756 311 760
rect 315 756 316 760
rect 310 755 316 756
rect 350 760 356 761
rect 350 756 351 760
rect 355 756 356 760
rect 350 755 356 756
rect 390 760 396 761
rect 390 756 391 760
rect 395 756 396 760
rect 390 755 396 756
rect 430 760 436 761
rect 430 756 431 760
rect 435 756 436 760
rect 686 757 687 761
rect 691 757 692 761
rect 686 756 692 757
rect 430 755 436 756
rect 278 754 285 755
rect 134 745 140 746
rect 110 743 116 744
rect 110 739 111 743
rect 115 739 116 743
rect 134 741 135 745
rect 139 741 140 745
rect 134 740 140 741
rect 174 745 180 746
rect 174 741 175 745
rect 179 741 180 745
rect 174 740 180 741
rect 214 745 220 746
rect 214 741 215 745
rect 219 741 220 745
rect 214 740 220 741
rect 254 745 260 746
rect 254 741 255 745
rect 259 741 260 745
rect 254 740 260 741
rect 294 745 300 746
rect 294 741 295 745
rect 299 741 300 745
rect 294 740 300 741
rect 334 745 340 746
rect 334 741 335 745
rect 339 741 340 745
rect 334 740 340 741
rect 374 745 380 746
rect 374 741 375 745
rect 379 741 380 745
rect 374 740 380 741
rect 414 745 420 746
rect 414 741 415 745
rect 419 741 420 745
rect 414 740 420 741
rect 686 743 692 744
rect 110 738 116 739
rect 142 739 149 740
rect 142 735 143 739
rect 148 735 149 739
rect 159 739 165 740
rect 159 738 160 739
rect 142 734 149 735
rect 152 736 160 738
rect 143 727 149 728
rect 143 723 144 727
rect 148 726 149 727
rect 152 726 154 736
rect 159 735 160 736
rect 164 735 165 739
rect 198 739 205 740
rect 159 734 165 735
rect 183 735 189 736
rect 183 731 184 735
rect 188 734 189 735
rect 198 735 199 739
rect 204 735 205 739
rect 198 734 205 735
rect 222 739 229 740
rect 222 735 223 739
rect 228 735 229 739
rect 239 739 245 740
rect 239 738 240 739
rect 222 734 229 735
rect 232 736 240 738
rect 188 732 194 734
rect 188 731 189 732
rect 183 730 189 731
rect 192 730 194 732
rect 232 730 234 736
rect 239 735 240 736
rect 244 735 245 739
rect 303 739 312 740
rect 239 734 245 735
rect 263 735 269 736
rect 263 731 264 735
rect 268 734 269 735
rect 303 735 304 739
rect 311 735 312 739
rect 303 734 312 735
rect 319 739 325 740
rect 319 735 320 739
rect 324 735 325 739
rect 354 739 365 740
rect 319 734 325 735
rect 343 735 349 736
rect 268 732 275 734
rect 268 731 269 732
rect 263 730 269 731
rect 273 730 275 732
rect 319 730 321 734
rect 343 731 344 735
rect 348 734 349 735
rect 354 735 355 739
rect 359 735 360 739
rect 364 735 365 739
rect 398 739 405 740
rect 354 734 365 735
rect 383 735 389 736
rect 348 731 350 734
rect 343 730 350 731
rect 383 731 384 735
rect 388 734 389 735
rect 398 735 399 739
rect 404 735 405 739
rect 439 739 445 740
rect 439 738 440 739
rect 398 734 405 735
rect 408 736 440 738
rect 388 732 394 734
rect 388 731 389 732
rect 383 730 389 731
rect 392 730 394 732
rect 408 730 410 736
rect 439 735 440 736
rect 444 735 445 739
rect 686 739 687 743
rect 691 739 692 743
rect 686 738 692 739
rect 439 734 445 735
rect 192 728 234 730
rect 273 728 321 730
rect 348 728 354 730
rect 392 728 410 730
rect 148 724 154 726
rect 148 723 149 724
rect 143 722 149 723
rect 183 723 189 724
rect 183 722 184 723
rect 168 720 184 722
rect 159 719 165 720
rect 110 717 116 718
rect 110 713 111 717
rect 115 713 116 717
rect 110 712 116 713
rect 134 715 140 716
rect 134 711 135 715
rect 139 711 140 715
rect 159 715 160 719
rect 164 718 165 719
rect 168 718 170 720
rect 183 719 184 720
rect 188 719 189 723
rect 223 723 229 724
rect 223 722 224 723
rect 208 720 224 722
rect 183 718 189 719
rect 199 719 205 720
rect 164 716 170 718
rect 164 715 165 716
rect 159 714 165 715
rect 174 715 180 716
rect 134 710 140 711
rect 174 711 175 715
rect 179 711 180 715
rect 199 715 200 719
rect 204 718 205 719
rect 208 718 210 720
rect 223 719 224 720
rect 228 719 229 723
rect 263 723 269 724
rect 263 722 264 723
rect 248 720 264 722
rect 223 718 229 719
rect 239 719 245 720
rect 204 716 210 718
rect 204 715 205 716
rect 199 714 205 715
rect 214 715 220 716
rect 174 710 180 711
rect 214 711 215 715
rect 219 711 220 715
rect 239 715 240 719
rect 244 718 245 719
rect 248 718 250 720
rect 263 719 264 720
rect 268 719 269 723
rect 303 723 309 724
rect 303 722 304 723
rect 288 720 304 722
rect 263 718 269 719
rect 279 719 285 720
rect 244 716 250 718
rect 244 715 245 716
rect 239 714 245 715
rect 254 715 260 716
rect 214 710 220 711
rect 254 711 255 715
rect 259 711 260 715
rect 279 715 280 719
rect 284 718 285 719
rect 288 718 290 720
rect 303 719 304 720
rect 308 719 309 723
rect 343 723 349 724
rect 343 722 344 723
rect 321 720 344 722
rect 303 718 309 719
rect 319 719 325 720
rect 284 716 290 718
rect 284 715 285 716
rect 279 714 285 715
rect 294 715 300 716
rect 254 710 260 711
rect 294 711 295 715
rect 299 711 300 715
rect 319 715 320 719
rect 324 715 325 719
rect 343 719 344 720
rect 348 719 349 723
rect 352 722 354 728
rect 398 723 404 724
rect 398 722 399 723
rect 352 720 399 722
rect 343 718 349 719
rect 398 719 399 720
rect 403 719 404 723
rect 398 718 404 719
rect 686 717 692 718
rect 319 714 325 715
rect 334 715 340 716
rect 294 710 300 711
rect 334 711 335 715
rect 339 711 340 715
rect 686 713 687 717
rect 691 713 692 717
rect 686 712 692 713
rect 334 710 340 711
rect 359 707 365 708
rect 359 706 360 707
rect 144 704 360 706
rect 142 703 148 704
rect 110 699 116 700
rect 110 695 111 699
rect 115 695 116 699
rect 142 699 143 703
rect 147 699 148 703
rect 359 703 360 704
rect 364 703 365 707
rect 359 702 365 703
rect 142 698 148 699
rect 150 700 156 701
rect 150 696 151 700
rect 155 696 156 700
rect 150 695 156 696
rect 190 700 196 701
rect 190 696 191 700
rect 195 696 196 700
rect 190 695 196 696
rect 230 700 236 701
rect 230 696 231 700
rect 235 696 236 700
rect 230 695 236 696
rect 270 700 276 701
rect 270 696 271 700
rect 275 696 276 700
rect 270 695 276 696
rect 310 700 316 701
rect 310 696 311 700
rect 315 696 316 700
rect 310 695 316 696
rect 350 700 356 701
rect 350 696 351 700
rect 355 696 356 700
rect 350 695 356 696
rect 686 699 692 700
rect 686 695 687 699
rect 691 695 692 699
rect 110 694 116 695
rect 686 694 692 695
rect 110 649 116 650
rect 686 649 692 650
rect 110 645 111 649
rect 115 645 116 649
rect 110 644 116 645
rect 150 648 156 649
rect 150 644 151 648
rect 155 644 156 648
rect 150 643 156 644
rect 190 648 196 649
rect 190 644 191 648
rect 195 644 196 648
rect 190 643 196 644
rect 230 648 236 649
rect 230 644 231 648
rect 235 644 236 648
rect 230 643 236 644
rect 270 648 276 649
rect 270 644 271 648
rect 275 644 276 648
rect 270 643 276 644
rect 310 648 316 649
rect 310 644 311 648
rect 315 644 316 648
rect 310 643 316 644
rect 350 648 356 649
rect 350 644 351 648
rect 355 644 356 648
rect 686 645 687 649
rect 691 645 692 649
rect 686 644 692 645
rect 350 643 356 644
rect 134 633 140 634
rect 110 631 116 632
rect 110 627 111 631
rect 115 627 116 631
rect 134 629 135 633
rect 139 629 140 633
rect 134 628 140 629
rect 174 633 180 634
rect 174 629 175 633
rect 179 629 180 633
rect 174 628 180 629
rect 214 633 220 634
rect 214 629 215 633
rect 219 629 220 633
rect 214 628 220 629
rect 254 633 260 634
rect 254 629 255 633
rect 259 629 260 633
rect 254 628 260 629
rect 294 633 300 634
rect 294 629 295 633
rect 299 629 300 633
rect 294 628 300 629
rect 334 633 340 634
rect 334 629 335 633
rect 339 629 340 633
rect 334 628 340 629
rect 686 631 692 632
rect 110 626 116 627
rect 142 627 149 628
rect 142 623 143 627
rect 148 623 149 627
rect 142 622 149 623
rect 159 627 165 628
rect 159 623 160 627
rect 164 626 165 627
rect 183 627 189 628
rect 183 626 184 627
rect 164 624 184 626
rect 164 623 165 624
rect 159 622 165 623
rect 183 623 184 624
rect 188 623 189 627
rect 183 622 189 623
rect 199 627 205 628
rect 199 623 200 627
rect 204 626 205 627
rect 223 627 229 628
rect 223 626 224 627
rect 204 624 224 626
rect 204 623 205 624
rect 199 622 205 623
rect 223 623 224 624
rect 228 623 229 627
rect 223 622 229 623
rect 239 627 245 628
rect 239 623 240 627
rect 244 626 245 627
rect 263 627 269 628
rect 263 626 264 627
rect 244 624 264 626
rect 244 623 245 624
rect 239 622 245 623
rect 263 623 264 624
rect 268 623 269 627
rect 263 622 269 623
rect 279 627 285 628
rect 279 623 280 627
rect 284 626 285 627
rect 303 627 309 628
rect 303 626 304 627
rect 284 624 304 626
rect 284 623 285 624
rect 279 622 285 623
rect 303 623 304 624
rect 308 623 309 627
rect 303 622 309 623
rect 319 627 325 628
rect 319 623 320 627
rect 324 626 325 627
rect 343 627 349 628
rect 343 626 344 627
rect 324 624 344 626
rect 324 623 325 624
rect 319 622 325 623
rect 343 623 344 624
rect 348 623 349 627
rect 343 622 349 623
rect 359 627 365 628
rect 359 623 360 627
rect 364 623 365 627
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 359 622 365 623
rect 361 610 363 622
rect 176 608 363 610
rect 143 607 149 608
rect 143 603 144 607
rect 148 606 149 607
rect 176 606 178 608
rect 148 604 178 606
rect 148 603 149 604
rect 143 602 149 603
rect 183 603 189 604
rect 183 602 184 603
rect 168 600 184 602
rect 159 599 165 600
rect 110 597 116 598
rect 110 593 111 597
rect 115 593 116 597
rect 110 592 116 593
rect 134 595 140 596
rect 134 591 135 595
rect 139 591 140 595
rect 159 595 160 599
rect 164 598 165 599
rect 168 598 170 600
rect 183 599 184 600
rect 188 599 189 603
rect 223 603 229 604
rect 223 602 224 603
rect 208 600 224 602
rect 183 598 189 599
rect 199 599 205 600
rect 164 596 170 598
rect 164 595 165 596
rect 159 594 165 595
rect 174 595 180 596
rect 134 590 140 591
rect 174 591 175 595
rect 179 591 180 595
rect 199 595 200 599
rect 204 598 205 599
rect 208 598 210 600
rect 223 599 224 600
rect 228 599 229 603
rect 263 603 269 604
rect 263 602 264 603
rect 248 600 264 602
rect 223 598 229 599
rect 239 599 245 600
rect 204 596 210 598
rect 204 595 205 596
rect 199 594 205 595
rect 214 595 220 596
rect 174 590 180 591
rect 214 591 215 595
rect 219 591 220 595
rect 239 595 240 599
rect 244 598 245 599
rect 248 598 250 600
rect 263 599 264 600
rect 268 599 269 603
rect 303 603 309 604
rect 303 602 304 603
rect 288 600 304 602
rect 263 598 269 599
rect 279 599 285 600
rect 244 596 250 598
rect 244 595 245 596
rect 239 594 245 595
rect 254 595 260 596
rect 214 590 220 591
rect 254 591 255 595
rect 259 591 260 595
rect 279 595 280 599
rect 284 598 285 599
rect 288 598 290 600
rect 303 599 304 600
rect 308 599 309 603
rect 303 598 309 599
rect 284 596 290 598
rect 686 597 692 598
rect 284 595 285 596
rect 279 594 285 595
rect 294 595 300 596
rect 254 590 260 591
rect 294 591 295 595
rect 299 591 300 595
rect 686 593 687 597
rect 691 593 692 597
rect 686 592 692 593
rect 294 590 300 591
rect 319 587 325 588
rect 319 586 320 587
rect 144 584 320 586
rect 142 583 148 584
rect 110 579 116 580
rect 110 575 111 579
rect 115 575 116 579
rect 142 579 143 583
rect 147 579 148 583
rect 319 583 320 584
rect 324 583 325 587
rect 319 582 325 583
rect 142 578 148 579
rect 150 580 156 581
rect 150 576 151 580
rect 155 576 156 580
rect 150 575 156 576
rect 190 580 196 581
rect 190 576 191 580
rect 195 576 196 580
rect 190 575 196 576
rect 230 580 236 581
rect 230 576 231 580
rect 235 576 236 580
rect 230 575 236 576
rect 270 580 276 581
rect 270 576 271 580
rect 275 576 276 580
rect 270 575 276 576
rect 310 580 316 581
rect 310 576 311 580
rect 315 576 316 580
rect 310 575 316 576
rect 686 579 692 580
rect 686 575 687 579
rect 691 575 692 579
rect 110 574 116 575
rect 686 574 692 575
rect 110 533 116 534
rect 686 533 692 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 150 532 156 533
rect 150 528 151 532
rect 155 528 156 532
rect 150 527 156 528
rect 190 532 196 533
rect 190 528 191 532
rect 195 528 196 532
rect 190 527 196 528
rect 230 532 236 533
rect 230 528 231 532
rect 235 528 236 532
rect 230 527 236 528
rect 270 532 276 533
rect 270 528 271 532
rect 275 528 276 532
rect 270 527 276 528
rect 310 532 316 533
rect 310 528 311 532
rect 315 528 316 532
rect 310 527 316 528
rect 350 532 356 533
rect 350 528 351 532
rect 355 528 356 532
rect 686 529 687 533
rect 691 529 692 533
rect 686 528 692 529
rect 350 527 356 528
rect 134 517 140 518
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 134 513 135 517
rect 139 513 140 517
rect 134 512 140 513
rect 174 517 180 518
rect 174 513 175 517
rect 179 513 180 517
rect 174 512 180 513
rect 214 517 220 518
rect 214 513 215 517
rect 219 513 220 517
rect 214 512 220 513
rect 254 517 260 518
rect 254 513 255 517
rect 259 513 260 517
rect 254 512 260 513
rect 294 517 300 518
rect 294 513 295 517
rect 299 513 300 517
rect 294 512 300 513
rect 334 517 340 518
rect 334 513 335 517
rect 339 513 340 517
rect 334 512 340 513
rect 686 515 692 516
rect 110 510 116 511
rect 142 511 149 512
rect 142 507 143 511
rect 148 507 149 511
rect 142 506 149 507
rect 159 511 165 512
rect 159 507 160 511
rect 164 510 165 511
rect 183 511 189 512
rect 183 510 184 511
rect 164 508 184 510
rect 164 507 165 508
rect 159 506 165 507
rect 183 507 184 508
rect 188 507 189 511
rect 183 506 189 507
rect 199 511 205 512
rect 199 507 200 511
rect 204 510 205 511
rect 223 511 229 512
rect 223 510 224 511
rect 204 508 224 510
rect 204 507 205 508
rect 199 506 205 507
rect 223 507 224 508
rect 228 507 229 511
rect 223 506 229 507
rect 239 511 245 512
rect 239 507 240 511
rect 244 510 245 511
rect 263 511 269 512
rect 263 510 264 511
rect 244 508 264 510
rect 244 507 245 508
rect 239 506 245 507
rect 263 507 264 508
rect 268 507 269 511
rect 263 506 269 507
rect 279 511 285 512
rect 279 507 280 511
rect 284 510 285 511
rect 303 511 309 512
rect 303 510 304 511
rect 284 508 304 510
rect 284 507 285 508
rect 279 506 285 507
rect 303 507 304 508
rect 308 507 309 511
rect 303 506 309 507
rect 319 511 325 512
rect 319 507 320 511
rect 324 510 325 511
rect 343 511 349 512
rect 343 510 344 511
rect 324 508 344 510
rect 324 507 325 508
rect 319 506 325 507
rect 343 507 344 508
rect 348 507 349 511
rect 343 506 349 507
rect 359 511 365 512
rect 359 507 360 511
rect 364 507 365 511
rect 686 511 687 515
rect 691 511 692 515
rect 686 510 692 511
rect 359 506 365 507
rect 361 498 363 506
rect 176 496 363 498
rect 143 495 149 496
rect 143 491 144 495
rect 148 494 149 495
rect 176 494 178 496
rect 148 492 178 494
rect 148 491 149 492
rect 143 490 149 491
rect 183 491 189 492
rect 183 490 184 491
rect 168 488 184 490
rect 159 487 165 488
rect 110 485 116 486
rect 110 481 111 485
rect 115 481 116 485
rect 110 480 116 481
rect 134 483 140 484
rect 134 479 135 483
rect 139 479 140 483
rect 159 483 160 487
rect 164 486 165 487
rect 168 486 170 488
rect 183 487 184 488
rect 188 487 189 491
rect 223 491 229 492
rect 223 490 224 491
rect 208 488 224 490
rect 183 486 189 487
rect 199 487 205 488
rect 164 484 170 486
rect 164 483 165 484
rect 159 482 165 483
rect 174 483 180 484
rect 134 478 140 479
rect 174 479 175 483
rect 179 479 180 483
rect 199 483 200 487
rect 204 486 205 487
rect 208 486 210 488
rect 223 487 224 488
rect 228 487 229 491
rect 263 491 269 492
rect 263 490 264 491
rect 248 488 264 490
rect 223 486 229 487
rect 239 487 245 488
rect 204 484 210 486
rect 204 483 205 484
rect 199 482 205 483
rect 214 483 220 484
rect 174 478 180 479
rect 214 479 215 483
rect 219 479 220 483
rect 239 483 240 487
rect 244 486 245 487
rect 248 486 250 488
rect 263 487 264 488
rect 268 487 269 491
rect 303 491 309 492
rect 303 490 304 491
rect 288 488 304 490
rect 263 486 269 487
rect 279 487 285 488
rect 244 484 250 486
rect 244 483 245 484
rect 239 482 245 483
rect 254 483 260 484
rect 214 478 220 479
rect 254 479 255 483
rect 259 479 260 483
rect 279 483 280 487
rect 284 486 285 487
rect 288 486 290 488
rect 303 487 304 488
rect 308 487 309 491
rect 343 491 349 492
rect 343 490 344 491
rect 321 488 344 490
rect 303 486 309 487
rect 319 487 325 488
rect 284 484 290 486
rect 284 483 285 484
rect 279 482 285 483
rect 294 483 300 484
rect 254 478 260 479
rect 294 479 295 483
rect 299 479 300 483
rect 319 483 320 487
rect 324 483 325 487
rect 343 487 344 488
rect 348 487 349 491
rect 383 491 389 492
rect 383 490 384 491
rect 361 488 384 490
rect 343 486 349 487
rect 359 487 365 488
rect 319 482 325 483
rect 334 483 340 484
rect 294 478 300 479
rect 334 479 335 483
rect 339 479 340 483
rect 359 483 360 487
rect 364 483 365 487
rect 383 487 384 488
rect 388 487 389 491
rect 383 486 389 487
rect 686 485 692 486
rect 359 482 365 483
rect 374 483 380 484
rect 334 478 340 479
rect 374 479 375 483
rect 379 479 380 483
rect 686 481 687 485
rect 691 481 692 485
rect 686 480 692 481
rect 374 478 380 479
rect 286 475 292 476
rect 286 471 287 475
rect 291 474 292 475
rect 399 475 405 476
rect 399 474 400 475
rect 291 472 400 474
rect 291 471 292 472
rect 286 470 292 471
rect 399 471 400 472
rect 404 471 405 475
rect 399 470 405 471
rect 150 468 156 469
rect 110 467 116 468
rect 110 463 111 467
rect 115 463 116 467
rect 150 464 151 468
rect 155 464 156 468
rect 150 463 156 464
rect 190 468 196 469
rect 190 464 191 468
rect 195 464 196 468
rect 190 463 196 464
rect 230 468 236 469
rect 230 464 231 468
rect 235 464 236 468
rect 230 463 236 464
rect 270 468 276 469
rect 270 464 271 468
rect 275 464 276 468
rect 270 463 276 464
rect 310 468 316 469
rect 310 464 311 468
rect 315 464 316 468
rect 310 463 316 464
rect 350 468 356 469
rect 350 464 351 468
rect 355 464 356 468
rect 350 463 356 464
rect 390 468 396 469
rect 390 464 391 468
rect 395 464 396 468
rect 390 463 396 464
rect 686 467 692 468
rect 686 463 687 467
rect 691 463 692 467
rect 110 462 116 463
rect 686 462 692 463
rect 110 417 116 418
rect 686 417 692 418
rect 110 413 111 417
rect 115 413 116 417
rect 110 412 116 413
rect 278 416 284 417
rect 278 412 279 416
rect 283 412 284 416
rect 278 411 284 412
rect 318 416 324 417
rect 318 412 319 416
rect 323 412 324 416
rect 318 411 324 412
rect 358 416 364 417
rect 358 412 359 416
rect 363 412 364 416
rect 358 411 364 412
rect 406 416 412 417
rect 406 412 407 416
rect 411 412 412 416
rect 406 411 412 412
rect 454 416 460 417
rect 454 412 455 416
rect 459 412 460 416
rect 454 411 460 412
rect 502 416 508 417
rect 502 412 503 416
rect 507 412 508 416
rect 502 411 508 412
rect 550 416 556 417
rect 550 412 551 416
rect 555 412 556 416
rect 550 411 556 412
rect 606 416 612 417
rect 606 412 607 416
rect 611 412 612 416
rect 606 411 612 412
rect 654 416 660 417
rect 654 412 655 416
rect 659 412 660 416
rect 686 413 687 417
rect 691 413 692 417
rect 686 412 692 413
rect 654 411 660 412
rect 262 401 268 402
rect 110 399 116 400
rect 110 395 111 399
rect 115 395 116 399
rect 262 397 263 401
rect 267 397 268 401
rect 262 396 268 397
rect 302 401 308 402
rect 302 397 303 401
rect 307 397 308 401
rect 302 396 308 397
rect 342 401 348 402
rect 342 397 343 401
rect 347 397 348 401
rect 342 396 348 397
rect 390 401 396 402
rect 390 397 391 401
rect 395 397 396 401
rect 390 396 396 397
rect 438 401 444 402
rect 438 397 439 401
rect 443 397 444 401
rect 438 396 444 397
rect 486 401 492 402
rect 486 397 487 401
rect 491 397 492 401
rect 486 396 492 397
rect 534 401 540 402
rect 534 397 535 401
rect 539 397 540 401
rect 534 396 540 397
rect 590 401 596 402
rect 590 397 591 401
rect 595 397 596 401
rect 590 396 596 397
rect 638 401 644 402
rect 638 397 639 401
rect 643 397 644 401
rect 638 396 644 397
rect 686 399 692 400
rect 110 394 116 395
rect 287 395 293 396
rect 271 391 277 392
rect 271 387 272 391
rect 276 387 277 391
rect 287 391 288 395
rect 292 394 293 395
rect 311 395 317 396
rect 311 394 312 395
rect 292 392 312 394
rect 292 391 293 392
rect 287 390 293 391
rect 311 391 312 392
rect 316 391 317 395
rect 311 390 317 391
rect 327 395 333 396
rect 327 391 328 395
rect 332 394 333 395
rect 351 395 357 396
rect 351 394 352 395
rect 332 392 352 394
rect 332 391 333 392
rect 327 390 333 391
rect 351 391 352 392
rect 356 391 357 395
rect 351 390 357 391
rect 367 395 373 396
rect 367 391 368 395
rect 372 394 373 395
rect 399 395 405 396
rect 399 394 400 395
rect 372 392 400 394
rect 372 391 373 392
rect 367 390 373 391
rect 399 391 400 392
rect 404 391 405 395
rect 399 390 405 391
rect 415 395 421 396
rect 415 391 416 395
rect 420 394 421 395
rect 447 395 453 396
rect 447 394 448 395
rect 420 392 448 394
rect 420 391 421 392
rect 415 390 421 391
rect 447 391 448 392
rect 452 391 453 395
rect 447 390 453 391
rect 463 395 469 396
rect 463 391 464 395
rect 468 394 469 395
rect 495 395 501 396
rect 495 394 496 395
rect 468 392 496 394
rect 468 391 469 392
rect 463 390 469 391
rect 495 391 496 392
rect 500 391 501 395
rect 511 395 517 396
rect 511 394 512 395
rect 495 390 501 391
rect 504 392 512 394
rect 271 386 277 387
rect 286 387 292 388
rect 286 386 287 387
rect 273 384 287 386
rect 207 383 213 384
rect 207 379 208 383
rect 212 382 213 383
rect 222 383 228 384
rect 222 382 223 383
rect 212 380 223 382
rect 212 379 213 380
rect 207 378 213 379
rect 222 379 223 380
rect 227 379 228 383
rect 286 383 287 384
rect 291 383 292 387
rect 504 386 506 392
rect 511 391 512 392
rect 516 391 517 395
rect 559 395 565 396
rect 511 390 517 391
rect 543 391 549 392
rect 543 387 544 391
rect 548 387 549 391
rect 559 391 560 395
rect 564 394 565 395
rect 599 395 605 396
rect 599 394 600 395
rect 564 392 600 394
rect 564 391 565 392
rect 559 390 565 391
rect 599 391 600 392
rect 604 391 605 395
rect 599 390 605 391
rect 615 395 621 396
rect 615 391 616 395
rect 620 394 621 395
rect 647 395 653 396
rect 647 394 648 395
rect 620 392 648 394
rect 620 391 621 392
rect 615 390 621 391
rect 647 391 648 392
rect 652 391 653 395
rect 647 390 653 391
rect 663 395 669 396
rect 663 391 664 395
rect 668 391 669 395
rect 686 395 687 399
rect 691 395 692 399
rect 686 394 692 395
rect 663 390 669 391
rect 543 386 549 387
rect 440 384 506 386
rect 286 382 292 383
rect 407 383 413 384
rect 222 378 228 379
rect 247 379 253 380
rect 247 378 248 379
rect 233 376 248 378
rect 223 375 229 376
rect 110 373 116 374
rect 110 369 111 373
rect 115 369 116 373
rect 110 368 116 369
rect 198 371 204 372
rect 198 367 199 371
rect 203 367 204 371
rect 223 371 224 375
rect 228 374 229 375
rect 233 374 235 376
rect 247 375 248 376
rect 252 375 253 379
rect 247 374 253 375
rect 287 379 293 380
rect 287 375 288 379
rect 292 378 293 379
rect 327 379 333 380
rect 292 376 307 378
rect 292 375 293 376
rect 287 374 293 375
rect 228 372 235 374
rect 228 371 229 372
rect 223 370 229 371
rect 238 371 244 372
rect 198 366 204 367
rect 238 367 239 371
rect 243 367 244 371
rect 238 366 244 367
rect 278 371 284 372
rect 278 367 279 371
rect 283 367 284 371
rect 278 366 284 367
rect 305 366 307 376
rect 327 375 328 379
rect 332 378 333 379
rect 367 379 373 380
rect 332 376 354 378
rect 332 375 333 376
rect 327 374 333 375
rect 318 371 324 372
rect 318 367 319 371
rect 323 367 324 371
rect 318 366 324 367
rect 305 364 310 366
rect 222 363 228 364
rect 222 359 223 363
rect 227 362 228 363
rect 308 362 310 364
rect 343 363 349 364
rect 343 362 344 363
rect 227 360 306 362
rect 308 360 344 362
rect 227 359 228 360
rect 222 358 228 359
rect 214 356 220 357
rect 110 355 116 356
rect 110 351 111 355
rect 115 351 116 355
rect 214 352 215 356
rect 219 352 220 356
rect 214 351 220 352
rect 254 356 260 357
rect 294 356 300 357
rect 304 356 306 360
rect 343 359 344 360
rect 348 359 349 363
rect 352 362 354 376
rect 367 375 368 379
rect 372 378 373 379
rect 407 379 408 383
rect 412 382 413 383
rect 440 382 442 384
rect 412 380 442 382
rect 412 379 413 380
rect 407 378 413 379
rect 446 379 453 380
rect 372 376 394 378
rect 372 375 373 376
rect 367 374 373 375
rect 358 371 364 372
rect 358 367 359 371
rect 363 367 364 371
rect 358 366 364 367
rect 383 363 389 364
rect 383 362 384 363
rect 352 360 384 362
rect 343 358 349 359
rect 383 359 384 360
rect 388 359 389 363
rect 392 362 394 376
rect 446 375 447 379
rect 452 375 453 379
rect 487 379 493 380
rect 487 378 488 379
rect 472 376 488 378
rect 446 374 453 375
rect 463 375 469 376
rect 398 371 404 372
rect 398 367 399 371
rect 403 367 404 371
rect 398 366 404 367
rect 438 371 444 372
rect 438 367 439 371
rect 443 367 444 371
rect 463 371 464 375
rect 468 374 469 375
rect 472 374 474 376
rect 487 375 488 376
rect 492 375 493 379
rect 527 379 533 380
rect 527 378 528 379
rect 512 376 528 378
rect 487 374 493 375
rect 503 375 509 376
rect 468 372 474 374
rect 468 371 469 372
rect 463 370 469 371
rect 478 371 484 372
rect 438 366 444 367
rect 478 367 479 371
rect 483 367 484 371
rect 503 371 504 375
rect 508 374 509 375
rect 512 374 514 376
rect 527 375 528 376
rect 532 375 533 379
rect 544 376 546 386
rect 647 383 653 384
rect 567 379 573 380
rect 527 374 533 375
rect 543 375 549 376
rect 508 372 514 374
rect 508 371 509 372
rect 503 370 509 371
rect 518 371 524 372
rect 478 366 484 367
rect 518 367 519 371
rect 523 367 524 371
rect 543 371 544 375
rect 548 371 549 375
rect 567 375 568 379
rect 572 378 573 379
rect 607 379 613 380
rect 572 376 594 378
rect 572 375 573 376
rect 567 374 573 375
rect 543 370 549 371
rect 558 371 564 372
rect 518 366 524 367
rect 558 367 559 371
rect 563 367 564 371
rect 558 366 564 367
rect 423 363 429 364
rect 423 362 424 363
rect 392 360 424 362
rect 383 358 389 359
rect 423 359 424 360
rect 428 359 429 363
rect 592 362 594 376
rect 607 375 608 379
rect 612 378 613 379
rect 647 379 648 383
rect 652 382 653 383
rect 665 382 667 390
rect 652 380 667 382
rect 652 379 653 380
rect 647 378 653 379
rect 612 376 634 378
rect 612 375 613 376
rect 607 374 613 375
rect 598 371 604 372
rect 598 367 599 371
rect 603 367 604 371
rect 598 366 604 367
rect 623 363 629 364
rect 623 362 624 363
rect 592 360 624 362
rect 423 358 429 359
rect 623 359 624 360
rect 628 359 629 363
rect 632 362 634 376
rect 686 373 692 374
rect 638 371 644 372
rect 638 367 639 371
rect 643 367 644 371
rect 686 369 687 373
rect 691 369 692 373
rect 686 368 692 369
rect 638 366 644 367
rect 663 363 669 364
rect 663 362 664 363
rect 632 360 664 362
rect 623 358 629 359
rect 663 359 664 360
rect 668 359 669 363
rect 663 358 669 359
rect 334 356 340 357
rect 254 352 255 356
rect 259 352 260 356
rect 254 351 260 352
rect 263 355 269 356
rect 263 351 264 355
rect 268 354 269 355
rect 286 355 292 356
rect 286 354 287 355
rect 268 352 287 354
rect 268 351 269 352
rect 110 350 116 351
rect 263 350 269 351
rect 286 351 287 352
rect 291 351 292 355
rect 294 352 295 356
rect 299 352 300 356
rect 294 351 300 352
rect 303 355 309 356
rect 303 351 304 355
rect 308 351 309 355
rect 334 352 335 356
rect 339 352 340 356
rect 334 351 340 352
rect 374 356 380 357
rect 374 352 375 356
rect 379 352 380 356
rect 374 351 380 352
rect 414 356 420 357
rect 414 352 415 356
rect 419 352 420 356
rect 414 351 420 352
rect 454 356 460 357
rect 454 352 455 356
rect 459 352 460 356
rect 454 351 460 352
rect 494 356 500 357
rect 494 352 495 356
rect 499 352 500 356
rect 494 351 500 352
rect 534 356 540 357
rect 534 352 535 356
rect 539 352 540 356
rect 534 351 540 352
rect 574 356 580 357
rect 614 356 620 357
rect 574 352 575 356
rect 579 352 580 356
rect 574 351 580 352
rect 583 355 589 356
rect 583 351 584 355
rect 588 354 589 355
rect 598 355 604 356
rect 598 354 599 355
rect 588 352 599 354
rect 588 351 589 352
rect 286 350 292 351
rect 303 350 309 351
rect 583 350 589 351
rect 598 351 599 352
rect 603 351 604 355
rect 614 352 615 356
rect 619 352 620 356
rect 614 351 620 352
rect 654 356 660 357
rect 654 352 655 356
rect 659 352 660 356
rect 654 351 660 352
rect 686 355 692 356
rect 686 351 687 355
rect 691 351 692 355
rect 598 350 604 351
rect 686 350 692 351
rect 446 339 452 340
rect 446 335 447 339
rect 451 338 452 339
rect 486 339 492 340
rect 486 338 487 339
rect 451 336 487 338
rect 451 335 452 336
rect 446 334 452 335
rect 486 335 487 336
rect 491 335 492 339
rect 486 334 492 335
rect 110 309 116 310
rect 686 309 692 310
rect 110 305 111 309
rect 115 305 116 309
rect 110 304 116 305
rect 222 308 228 309
rect 222 304 223 308
rect 227 304 228 308
rect 222 303 228 304
rect 262 308 268 309
rect 262 304 263 308
rect 267 304 268 308
rect 262 303 268 304
rect 310 308 316 309
rect 310 304 311 308
rect 315 304 316 308
rect 310 303 316 304
rect 366 308 372 309
rect 366 304 367 308
rect 371 304 372 308
rect 366 303 372 304
rect 422 308 428 309
rect 422 304 423 308
rect 427 304 428 308
rect 422 303 428 304
rect 478 308 484 309
rect 542 308 548 309
rect 478 304 479 308
rect 483 304 484 308
rect 478 303 484 304
rect 486 307 493 308
rect 486 303 487 307
rect 492 303 493 307
rect 542 304 543 308
rect 547 304 548 308
rect 542 303 548 304
rect 606 308 612 309
rect 606 304 607 308
rect 611 304 612 308
rect 606 303 612 304
rect 654 308 660 309
rect 654 304 655 308
rect 659 304 660 308
rect 686 305 687 309
rect 691 305 692 309
rect 686 304 692 305
rect 654 303 660 304
rect 486 302 493 303
rect 206 293 212 294
rect 110 291 116 292
rect 110 287 111 291
rect 115 287 116 291
rect 206 289 207 293
rect 211 289 212 293
rect 206 288 212 289
rect 246 293 252 294
rect 246 289 247 293
rect 251 289 252 293
rect 246 288 252 289
rect 294 293 300 294
rect 294 289 295 293
rect 299 289 300 293
rect 294 288 300 289
rect 350 293 356 294
rect 350 289 351 293
rect 355 289 356 293
rect 350 288 356 289
rect 406 293 412 294
rect 406 289 407 293
rect 411 289 412 293
rect 406 288 412 289
rect 462 293 468 294
rect 462 289 463 293
rect 467 289 468 293
rect 462 288 468 289
rect 526 293 532 294
rect 526 289 527 293
rect 531 289 532 293
rect 526 288 532 289
rect 590 293 596 294
rect 590 289 591 293
rect 595 289 596 293
rect 590 288 596 289
rect 638 293 644 294
rect 638 289 639 293
rect 643 289 644 293
rect 638 288 644 289
rect 686 291 692 292
rect 110 286 116 287
rect 231 287 237 288
rect 215 283 221 284
rect 215 279 216 283
rect 220 282 221 283
rect 231 283 232 287
rect 236 286 237 287
rect 255 287 261 288
rect 255 286 256 287
rect 236 284 256 286
rect 236 283 237 284
rect 231 282 237 283
rect 255 283 256 284
rect 260 283 261 287
rect 255 282 261 283
rect 271 287 280 288
rect 271 283 272 287
rect 279 283 280 287
rect 271 282 280 283
rect 286 287 292 288
rect 286 283 287 287
rect 291 286 292 287
rect 303 287 309 288
rect 303 286 304 287
rect 291 284 304 286
rect 291 283 292 284
rect 286 282 292 283
rect 303 283 304 284
rect 308 283 309 287
rect 303 282 309 283
rect 319 287 325 288
rect 319 283 320 287
rect 324 286 325 287
rect 359 287 365 288
rect 359 286 360 287
rect 324 284 360 286
rect 324 283 325 284
rect 319 282 325 283
rect 359 283 360 284
rect 364 283 365 287
rect 359 282 365 283
rect 375 287 381 288
rect 375 283 376 287
rect 380 286 381 287
rect 415 287 421 288
rect 415 286 416 287
rect 380 284 416 286
rect 380 283 381 284
rect 375 282 381 283
rect 415 283 416 284
rect 420 283 421 287
rect 431 287 437 288
rect 431 286 432 287
rect 415 282 421 283
rect 424 284 432 286
rect 220 280 226 282
rect 220 279 221 280
rect 215 278 221 279
rect 224 278 226 280
rect 424 278 426 284
rect 431 283 432 284
rect 436 283 437 287
rect 551 287 557 288
rect 551 286 552 287
rect 544 284 552 286
rect 431 282 437 283
rect 471 283 477 284
rect 471 279 472 283
rect 476 282 477 283
rect 490 283 496 284
rect 476 280 486 282
rect 476 279 477 280
rect 471 278 477 279
rect 224 276 426 278
rect 484 274 486 280
rect 490 279 491 283
rect 495 282 496 283
rect 535 283 541 284
rect 535 282 536 283
rect 495 280 536 282
rect 495 279 496 280
rect 490 278 496 279
rect 535 279 536 280
rect 540 279 541 283
rect 535 278 541 279
rect 544 274 546 284
rect 551 283 552 284
rect 556 283 557 287
rect 551 282 557 283
rect 598 287 605 288
rect 598 283 599 287
rect 604 283 605 287
rect 598 282 605 283
rect 615 287 621 288
rect 615 283 616 287
rect 620 286 621 287
rect 647 287 653 288
rect 647 286 648 287
rect 620 284 648 286
rect 620 283 621 284
rect 615 282 621 283
rect 647 283 648 284
rect 652 283 653 287
rect 663 287 669 288
rect 663 286 664 287
rect 647 282 653 283
rect 656 284 664 286
rect 484 272 546 274
rect 278 271 285 272
rect 151 267 157 268
rect 151 263 152 267
rect 156 266 157 267
rect 215 267 221 268
rect 156 264 194 266
rect 156 263 157 264
rect 151 262 157 263
rect 110 261 116 262
rect 110 257 111 261
rect 115 257 116 261
rect 110 256 116 257
rect 142 259 148 260
rect 142 255 143 259
rect 147 255 148 259
rect 142 254 148 255
rect 192 250 194 264
rect 215 263 216 267
rect 220 266 221 267
rect 278 267 279 271
rect 284 267 285 271
rect 647 271 653 272
rect 278 266 285 267
rect 343 267 349 268
rect 343 266 344 267
rect 220 264 266 266
rect 319 264 344 266
rect 220 263 221 264
rect 215 262 221 263
rect 206 259 212 260
rect 206 255 207 259
rect 211 255 212 259
rect 206 254 212 255
rect 231 251 237 252
rect 231 250 232 251
rect 192 248 232 250
rect 231 247 232 248
rect 236 247 237 251
rect 264 250 266 264
rect 295 263 301 264
rect 270 259 276 260
rect 270 255 271 259
rect 275 255 276 259
rect 295 259 296 263
rect 300 262 301 263
rect 319 262 321 264
rect 343 263 344 264
rect 348 263 349 267
rect 343 262 349 263
rect 390 267 396 268
rect 390 263 391 267
rect 395 266 396 267
rect 407 267 413 268
rect 407 266 408 267
rect 395 264 408 266
rect 395 263 396 264
rect 390 262 396 263
rect 407 263 408 264
rect 412 263 413 267
rect 471 267 477 268
rect 471 266 472 267
rect 448 264 472 266
rect 407 262 413 263
rect 423 263 429 264
rect 300 260 321 262
rect 300 259 301 260
rect 295 258 301 259
rect 334 259 340 260
rect 270 254 276 255
rect 334 255 335 259
rect 339 255 340 259
rect 334 254 340 255
rect 398 259 404 260
rect 398 255 399 259
rect 403 255 404 259
rect 423 259 424 263
rect 428 262 429 263
rect 448 262 450 264
rect 471 263 472 264
rect 476 263 477 267
rect 535 267 541 268
rect 471 262 477 263
rect 487 263 496 264
rect 428 260 450 262
rect 428 259 429 260
rect 423 258 429 259
rect 462 259 468 260
rect 398 254 404 255
rect 462 255 463 259
rect 467 255 468 259
rect 487 259 488 263
rect 495 259 496 263
rect 535 263 536 267
rect 540 266 541 267
rect 599 267 605 268
rect 540 264 578 266
rect 540 263 541 264
rect 535 262 541 263
rect 487 258 496 259
rect 526 259 532 260
rect 462 254 468 255
rect 526 255 527 259
rect 531 255 532 259
rect 526 254 532 255
rect 359 251 365 252
rect 359 250 360 251
rect 264 248 360 250
rect 231 246 237 247
rect 359 247 360 248
rect 364 247 365 251
rect 551 251 557 252
rect 551 250 552 251
rect 528 248 552 250
rect 359 246 365 247
rect 526 247 532 248
rect 158 244 164 245
rect 222 244 228 245
rect 110 243 116 244
rect 110 239 111 243
rect 115 239 116 243
rect 158 240 159 244
rect 163 240 164 244
rect 158 239 164 240
rect 167 243 173 244
rect 167 239 168 243
rect 172 242 173 243
rect 178 243 184 244
rect 178 242 179 243
rect 172 240 179 242
rect 172 239 173 240
rect 110 238 116 239
rect 167 238 173 239
rect 178 239 179 240
rect 183 239 184 243
rect 222 240 223 244
rect 227 240 228 244
rect 222 239 228 240
rect 286 244 292 245
rect 286 240 287 244
rect 291 240 292 244
rect 286 239 292 240
rect 350 244 356 245
rect 350 240 351 244
rect 355 240 356 244
rect 350 239 356 240
rect 414 244 420 245
rect 414 240 415 244
rect 419 240 420 244
rect 414 239 420 240
rect 478 244 484 245
rect 478 240 479 244
rect 483 240 484 244
rect 526 243 527 247
rect 531 243 532 247
rect 551 247 552 248
rect 556 247 557 251
rect 576 250 578 264
rect 599 263 600 267
rect 604 266 605 267
rect 647 267 648 271
rect 652 270 653 271
rect 656 270 658 284
rect 663 283 664 284
rect 668 283 669 287
rect 686 287 687 291
rect 691 287 692 291
rect 686 286 692 287
rect 663 282 669 283
rect 652 268 658 270
rect 652 267 653 268
rect 647 266 653 267
rect 604 264 634 266
rect 604 263 605 264
rect 599 262 605 263
rect 590 259 596 260
rect 590 255 591 259
rect 595 255 596 259
rect 590 254 596 255
rect 615 251 621 252
rect 615 250 616 251
rect 576 248 616 250
rect 551 246 557 247
rect 615 247 616 248
rect 620 247 621 251
rect 632 250 634 264
rect 686 261 692 262
rect 638 259 644 260
rect 638 255 639 259
rect 643 255 644 259
rect 686 257 687 261
rect 691 257 692 261
rect 686 256 692 257
rect 638 254 644 255
rect 663 251 669 252
rect 663 250 664 251
rect 632 248 664 250
rect 615 246 621 247
rect 663 247 664 248
rect 668 247 669 251
rect 663 246 669 247
rect 526 242 532 243
rect 542 244 548 245
rect 478 239 484 240
rect 542 240 543 244
rect 547 240 548 244
rect 542 239 548 240
rect 606 244 612 245
rect 606 240 607 244
rect 611 240 612 244
rect 606 239 612 240
rect 654 244 660 245
rect 654 240 655 244
rect 659 240 660 244
rect 654 239 660 240
rect 686 243 692 244
rect 686 239 687 243
rect 691 239 692 243
rect 178 238 184 239
rect 686 238 692 239
rect 110 193 116 194
rect 686 193 692 194
rect 110 189 111 193
rect 115 189 116 193
rect 110 188 116 189
rect 166 192 172 193
rect 166 188 167 192
rect 171 188 172 192
rect 166 187 172 188
rect 214 192 220 193
rect 214 188 215 192
rect 219 188 220 192
rect 214 187 220 188
rect 270 192 276 193
rect 270 188 271 192
rect 275 188 276 192
rect 270 187 276 188
rect 326 192 332 193
rect 326 188 327 192
rect 331 188 332 192
rect 326 187 332 188
rect 382 192 388 193
rect 438 192 444 193
rect 382 188 383 192
rect 387 188 388 192
rect 382 187 388 188
rect 390 191 397 192
rect 390 187 391 191
rect 396 187 397 191
rect 438 188 439 192
rect 443 188 444 192
rect 438 187 444 188
rect 494 192 500 193
rect 494 188 495 192
rect 499 188 500 192
rect 494 187 500 188
rect 550 192 556 193
rect 550 188 551 192
rect 555 188 556 192
rect 550 187 556 188
rect 614 192 620 193
rect 614 188 615 192
rect 619 188 620 192
rect 614 187 620 188
rect 654 192 660 193
rect 654 188 655 192
rect 659 188 660 192
rect 686 189 687 193
rect 691 189 692 193
rect 686 188 692 189
rect 654 187 660 188
rect 390 186 397 187
rect 150 177 156 178
rect 110 175 116 176
rect 110 171 111 175
rect 115 171 116 175
rect 150 173 151 177
rect 155 173 156 177
rect 150 172 156 173
rect 198 177 204 178
rect 198 173 199 177
rect 203 173 204 177
rect 198 172 204 173
rect 254 177 260 178
rect 254 173 255 177
rect 259 173 260 177
rect 254 172 260 173
rect 310 177 316 178
rect 310 173 311 177
rect 315 173 316 177
rect 310 172 316 173
rect 366 177 372 178
rect 366 173 367 177
rect 371 173 372 177
rect 366 172 372 173
rect 422 177 428 178
rect 422 173 423 177
rect 427 173 428 177
rect 422 172 428 173
rect 478 177 484 178
rect 478 173 479 177
rect 483 173 484 177
rect 478 172 484 173
rect 534 177 540 178
rect 534 173 535 177
rect 539 173 540 177
rect 534 172 540 173
rect 598 177 604 178
rect 598 173 599 177
rect 603 173 604 177
rect 598 172 604 173
rect 638 177 644 178
rect 638 173 639 177
rect 643 173 644 177
rect 638 172 644 173
rect 686 175 692 176
rect 110 170 116 171
rect 175 171 181 172
rect 159 167 165 168
rect 159 163 160 167
rect 164 166 165 167
rect 175 167 176 171
rect 180 170 181 171
rect 207 171 213 172
rect 207 170 208 171
rect 180 168 208 170
rect 180 167 181 168
rect 175 166 181 167
rect 207 167 208 168
rect 212 167 213 171
rect 207 166 213 167
rect 223 171 229 172
rect 223 167 224 171
rect 228 170 229 171
rect 263 171 269 172
rect 263 170 264 171
rect 228 168 264 170
rect 228 167 229 168
rect 223 166 229 167
rect 263 167 264 168
rect 268 167 269 171
rect 263 166 269 167
rect 279 171 285 172
rect 279 167 280 171
rect 284 170 285 171
rect 319 171 325 172
rect 319 170 320 171
rect 284 168 320 170
rect 284 167 285 168
rect 279 166 285 167
rect 319 167 320 168
rect 324 167 325 171
rect 335 171 341 172
rect 335 170 336 171
rect 319 166 325 167
rect 328 168 336 170
rect 164 163 166 166
rect 159 162 166 163
rect 178 163 184 164
rect 178 162 179 163
rect 164 160 179 162
rect 178 159 179 160
rect 183 159 184 163
rect 178 158 184 159
rect 328 158 330 168
rect 335 167 336 168
rect 340 167 341 171
rect 335 166 341 167
rect 375 171 384 172
rect 375 167 376 171
rect 383 167 384 171
rect 446 171 453 172
rect 375 166 384 167
rect 430 167 436 168
rect 430 163 431 167
rect 435 166 436 167
rect 446 167 447 171
rect 452 167 453 171
rect 503 171 509 172
rect 503 170 504 171
rect 496 168 504 170
rect 446 166 453 167
rect 486 167 493 168
rect 435 164 442 166
rect 435 163 436 164
rect 430 162 436 163
rect 192 156 330 158
rect 440 158 442 164
rect 486 163 487 167
rect 492 163 493 167
rect 486 162 493 163
rect 496 158 498 168
rect 503 167 504 168
rect 508 167 509 171
rect 503 166 509 167
rect 526 171 532 172
rect 526 167 527 171
rect 531 170 532 171
rect 543 171 549 172
rect 543 170 544 171
rect 531 168 544 170
rect 531 167 532 168
rect 526 166 532 167
rect 543 167 544 168
rect 548 167 549 171
rect 543 166 549 167
rect 559 171 565 172
rect 559 167 560 171
rect 564 170 565 171
rect 607 171 613 172
rect 607 170 608 171
rect 564 168 608 170
rect 564 167 565 168
rect 559 166 565 167
rect 607 167 608 168
rect 612 167 613 171
rect 607 166 613 167
rect 623 171 629 172
rect 623 167 624 171
rect 628 170 629 171
rect 647 171 653 172
rect 647 170 648 171
rect 628 168 648 170
rect 628 167 629 168
rect 623 166 629 167
rect 647 167 648 168
rect 652 167 653 171
rect 663 171 669 172
rect 663 170 664 171
rect 647 166 653 167
rect 656 168 664 170
rect 440 156 498 158
rect 159 155 165 156
rect 159 151 160 155
rect 164 154 165 155
rect 192 154 194 156
rect 164 152 194 154
rect 647 155 653 156
rect 164 151 165 152
rect 159 150 165 151
rect 199 151 205 152
rect 199 150 200 151
rect 184 148 200 150
rect 175 147 181 148
rect 110 145 116 146
rect 110 141 111 145
rect 115 141 116 145
rect 110 140 116 141
rect 150 143 156 144
rect 150 139 151 143
rect 155 139 156 143
rect 175 143 176 147
rect 180 146 181 147
rect 184 146 186 148
rect 199 147 200 148
rect 204 147 205 151
rect 239 151 245 152
rect 239 150 240 151
rect 224 148 240 150
rect 199 146 205 147
rect 215 147 221 148
rect 180 144 186 146
rect 180 143 181 144
rect 175 142 181 143
rect 190 143 196 144
rect 150 138 156 139
rect 190 139 191 143
rect 195 139 196 143
rect 215 143 216 147
rect 220 146 221 147
rect 224 146 226 148
rect 239 147 240 148
rect 244 147 245 151
rect 279 151 285 152
rect 279 150 280 151
rect 264 148 280 150
rect 239 146 245 147
rect 255 147 261 148
rect 220 144 226 146
rect 220 143 221 144
rect 215 142 221 143
rect 230 143 236 144
rect 190 138 196 139
rect 230 139 231 143
rect 235 139 236 143
rect 255 143 256 147
rect 260 146 261 147
rect 264 146 266 148
rect 279 147 280 148
rect 284 147 285 151
rect 319 151 325 152
rect 319 150 320 151
rect 304 148 320 150
rect 279 146 285 147
rect 295 147 301 148
rect 260 144 266 146
rect 260 143 261 144
rect 255 142 261 143
rect 270 143 276 144
rect 230 138 236 139
rect 270 139 271 143
rect 275 139 276 143
rect 295 143 296 147
rect 300 146 301 147
rect 304 146 306 148
rect 319 147 320 148
rect 324 147 325 151
rect 359 151 365 152
rect 359 150 360 151
rect 344 148 360 150
rect 319 146 325 147
rect 335 147 341 148
rect 300 144 306 146
rect 300 143 301 144
rect 295 142 301 143
rect 310 143 316 144
rect 270 138 276 139
rect 310 139 311 143
rect 315 139 316 143
rect 335 143 336 147
rect 340 146 341 147
rect 344 146 346 148
rect 359 147 360 148
rect 364 147 365 151
rect 399 151 405 152
rect 399 150 400 151
rect 384 148 400 150
rect 359 146 365 147
rect 375 147 381 148
rect 340 144 346 146
rect 340 143 341 144
rect 335 142 341 143
rect 350 143 356 144
rect 310 138 316 139
rect 350 139 351 143
rect 355 139 356 143
rect 375 143 376 147
rect 380 146 381 147
rect 384 146 386 148
rect 399 147 400 148
rect 404 147 405 151
rect 439 151 445 152
rect 439 150 440 151
rect 424 148 440 150
rect 399 146 405 147
rect 415 147 421 148
rect 380 144 386 146
rect 380 143 381 144
rect 375 142 381 143
rect 390 143 396 144
rect 350 138 356 139
rect 390 139 391 143
rect 395 139 396 143
rect 415 143 416 147
rect 420 146 421 147
rect 424 146 426 148
rect 439 147 440 148
rect 444 147 445 151
rect 479 151 485 152
rect 479 150 480 151
rect 464 148 480 150
rect 439 146 445 147
rect 455 147 461 148
rect 420 144 426 146
rect 420 143 421 144
rect 415 142 421 143
rect 430 143 436 144
rect 390 138 396 139
rect 430 139 431 143
rect 435 139 436 143
rect 455 143 456 147
rect 460 146 461 147
rect 464 146 466 148
rect 479 147 480 148
rect 484 147 485 151
rect 527 151 533 152
rect 527 150 528 151
rect 512 148 528 150
rect 479 146 485 147
rect 495 147 501 148
rect 460 144 466 146
rect 460 143 461 144
rect 455 142 461 143
rect 470 143 476 144
rect 430 138 436 139
rect 470 139 471 143
rect 475 139 476 143
rect 495 143 496 147
rect 500 146 501 147
rect 512 146 514 148
rect 527 147 528 148
rect 532 147 533 151
rect 527 146 533 147
rect 567 151 573 152
rect 567 147 568 151
rect 572 150 573 151
rect 607 151 613 152
rect 572 148 594 150
rect 572 147 573 148
rect 567 146 573 147
rect 500 144 514 146
rect 500 143 501 144
rect 495 142 501 143
rect 518 143 524 144
rect 470 138 476 139
rect 518 139 519 143
rect 523 139 524 143
rect 518 138 524 139
rect 558 143 564 144
rect 558 139 559 143
rect 563 139 564 143
rect 558 138 564 139
rect 494 135 500 136
rect 494 131 495 135
rect 499 134 500 135
rect 543 135 549 136
rect 543 134 544 135
rect 499 132 544 134
rect 499 131 500 132
rect 494 130 500 131
rect 543 131 544 132
rect 548 131 549 135
rect 592 134 594 148
rect 607 147 608 151
rect 612 150 613 151
rect 647 151 648 155
rect 652 154 653 155
rect 656 154 658 168
rect 663 167 664 168
rect 668 167 669 171
rect 686 171 687 175
rect 691 171 692 175
rect 686 170 692 171
rect 663 166 669 167
rect 652 152 658 154
rect 652 151 653 152
rect 647 150 653 151
rect 612 148 634 150
rect 612 147 613 148
rect 607 146 613 147
rect 598 143 604 144
rect 598 139 599 143
rect 603 139 604 143
rect 598 138 604 139
rect 623 135 629 136
rect 623 134 624 135
rect 592 132 624 134
rect 543 130 549 131
rect 623 131 624 132
rect 628 131 629 135
rect 632 134 634 148
rect 686 145 692 146
rect 638 143 644 144
rect 638 139 639 143
rect 643 139 644 143
rect 686 141 687 145
rect 691 141 692 145
rect 686 140 692 141
rect 638 138 644 139
rect 663 135 669 136
rect 663 134 664 135
rect 632 132 664 134
rect 623 130 629 131
rect 663 131 664 132
rect 668 131 669 135
rect 663 130 669 131
rect 166 128 172 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 166 124 167 128
rect 171 124 172 128
rect 166 123 172 124
rect 206 128 212 129
rect 206 124 207 128
rect 211 124 212 128
rect 206 123 212 124
rect 246 128 252 129
rect 246 124 247 128
rect 251 124 252 128
rect 246 123 252 124
rect 286 128 292 129
rect 286 124 287 128
rect 291 124 292 128
rect 286 123 292 124
rect 326 128 332 129
rect 326 124 327 128
rect 331 124 332 128
rect 326 123 332 124
rect 366 128 372 129
rect 366 124 367 128
rect 371 124 372 128
rect 366 123 372 124
rect 406 128 412 129
rect 406 124 407 128
rect 411 124 412 128
rect 406 123 412 124
rect 446 128 452 129
rect 446 124 447 128
rect 451 124 452 128
rect 446 123 452 124
rect 486 128 492 129
rect 486 124 487 128
rect 491 124 492 128
rect 486 123 492 124
rect 534 128 540 129
rect 534 124 535 128
rect 539 124 540 128
rect 534 123 540 124
rect 574 128 580 129
rect 574 124 575 128
rect 579 124 580 128
rect 574 123 580 124
rect 614 128 620 129
rect 614 124 615 128
rect 619 124 620 128
rect 614 123 620 124
rect 654 128 660 129
rect 654 124 655 128
rect 659 124 660 128
rect 654 123 660 124
rect 686 127 692 128
rect 686 123 687 127
rect 691 123 692 127
rect 110 122 116 123
rect 686 122 692 123
<< m3c >>
rect 223 775 227 779
rect 279 775 283 779
rect 111 757 115 761
rect 151 756 155 760
rect 191 756 195 760
rect 231 756 235 760
rect 271 756 275 760
rect 279 755 280 759
rect 280 755 283 759
rect 311 756 315 760
rect 351 756 355 760
rect 391 756 395 760
rect 431 756 435 760
rect 687 757 691 761
rect 111 739 115 743
rect 135 741 139 745
rect 175 741 179 745
rect 215 741 219 745
rect 255 741 259 745
rect 295 741 299 745
rect 335 741 339 745
rect 375 741 379 745
rect 415 741 419 745
rect 143 735 144 739
rect 144 735 147 739
rect 199 735 200 739
rect 200 735 203 739
rect 223 735 224 739
rect 224 735 227 739
rect 307 735 308 739
rect 308 735 311 739
rect 355 735 359 739
rect 399 735 400 739
rect 400 735 403 739
rect 687 739 691 743
rect 111 713 115 717
rect 135 711 139 715
rect 175 711 179 715
rect 215 711 219 715
rect 255 711 259 715
rect 295 711 299 715
rect 399 719 403 723
rect 335 711 339 715
rect 687 713 691 717
rect 111 695 115 699
rect 143 699 147 703
rect 151 696 155 700
rect 191 696 195 700
rect 231 696 235 700
rect 271 696 275 700
rect 311 696 315 700
rect 351 696 355 700
rect 687 695 691 699
rect 111 645 115 649
rect 151 644 155 648
rect 191 644 195 648
rect 231 644 235 648
rect 271 644 275 648
rect 311 644 315 648
rect 351 644 355 648
rect 687 645 691 649
rect 111 627 115 631
rect 135 629 139 633
rect 175 629 179 633
rect 215 629 219 633
rect 255 629 259 633
rect 295 629 299 633
rect 335 629 339 633
rect 143 623 144 627
rect 144 623 147 627
rect 687 627 691 631
rect 111 593 115 597
rect 135 591 139 595
rect 175 591 179 595
rect 215 591 219 595
rect 255 591 259 595
rect 295 591 299 595
rect 687 593 691 597
rect 111 575 115 579
rect 143 579 147 583
rect 151 576 155 580
rect 191 576 195 580
rect 231 576 235 580
rect 271 576 275 580
rect 311 576 315 580
rect 687 575 691 579
rect 111 529 115 533
rect 151 528 155 532
rect 191 528 195 532
rect 231 528 235 532
rect 271 528 275 532
rect 311 528 315 532
rect 351 528 355 532
rect 687 529 691 533
rect 111 511 115 515
rect 135 513 139 517
rect 175 513 179 517
rect 215 513 219 517
rect 255 513 259 517
rect 295 513 299 517
rect 335 513 339 517
rect 143 507 144 511
rect 144 507 147 511
rect 687 511 691 515
rect 111 481 115 485
rect 135 479 139 483
rect 175 479 179 483
rect 215 479 219 483
rect 255 479 259 483
rect 295 479 299 483
rect 335 479 339 483
rect 375 479 379 483
rect 687 481 691 485
rect 287 471 291 475
rect 111 463 115 467
rect 151 464 155 468
rect 191 464 195 468
rect 231 464 235 468
rect 271 464 275 468
rect 311 464 315 468
rect 351 464 355 468
rect 391 464 395 468
rect 687 463 691 467
rect 111 413 115 417
rect 279 412 283 416
rect 319 412 323 416
rect 359 412 363 416
rect 407 412 411 416
rect 455 412 459 416
rect 503 412 507 416
rect 551 412 555 416
rect 607 412 611 416
rect 655 412 659 416
rect 687 413 691 417
rect 111 395 115 399
rect 263 397 267 401
rect 303 397 307 401
rect 343 397 347 401
rect 391 397 395 401
rect 439 397 443 401
rect 487 397 491 401
rect 535 397 539 401
rect 591 397 595 401
rect 639 397 643 401
rect 223 379 227 383
rect 287 383 291 387
rect 687 395 691 399
rect 111 369 115 373
rect 199 367 203 371
rect 239 367 243 371
rect 279 367 283 371
rect 319 367 323 371
rect 223 359 227 363
rect 111 351 115 355
rect 215 352 219 356
rect 359 367 363 371
rect 447 375 448 379
rect 448 375 451 379
rect 399 367 403 371
rect 439 367 443 371
rect 479 367 483 371
rect 519 367 523 371
rect 559 367 563 371
rect 599 367 603 371
rect 639 367 643 371
rect 687 369 691 373
rect 255 352 259 356
rect 287 351 291 355
rect 295 352 299 356
rect 335 352 339 356
rect 375 352 379 356
rect 415 352 419 356
rect 455 352 459 356
rect 495 352 499 356
rect 535 352 539 356
rect 575 352 579 356
rect 599 351 603 355
rect 615 352 619 356
rect 655 352 659 356
rect 687 351 691 355
rect 447 335 451 339
rect 487 335 491 339
rect 111 305 115 309
rect 223 304 227 308
rect 263 304 267 308
rect 311 304 315 308
rect 367 304 371 308
rect 423 304 427 308
rect 479 304 483 308
rect 487 303 488 307
rect 488 303 491 307
rect 543 304 547 308
rect 607 304 611 308
rect 655 304 659 308
rect 687 305 691 309
rect 111 287 115 291
rect 207 289 211 293
rect 247 289 251 293
rect 295 289 299 293
rect 351 289 355 293
rect 407 289 411 293
rect 463 289 467 293
rect 527 289 531 293
rect 591 289 595 293
rect 639 289 643 293
rect 275 283 276 287
rect 276 283 279 287
rect 287 283 291 287
rect 491 279 495 283
rect 599 283 600 287
rect 600 283 603 287
rect 111 257 115 261
rect 143 255 147 259
rect 279 267 280 271
rect 280 267 283 271
rect 207 255 211 259
rect 271 255 275 259
rect 391 263 395 267
rect 335 255 339 259
rect 399 255 403 259
rect 463 255 467 259
rect 491 259 492 263
rect 492 259 495 263
rect 527 255 531 259
rect 111 239 115 243
rect 159 240 163 244
rect 179 239 183 243
rect 223 240 227 244
rect 287 240 291 244
rect 351 240 355 244
rect 415 240 419 244
rect 479 240 483 244
rect 527 243 531 247
rect 687 287 691 291
rect 591 255 595 259
rect 639 255 643 259
rect 687 257 691 261
rect 543 240 547 244
rect 607 240 611 244
rect 655 240 659 244
rect 687 239 691 243
rect 111 189 115 193
rect 167 188 171 192
rect 215 188 219 192
rect 271 188 275 192
rect 327 188 331 192
rect 383 188 387 192
rect 391 187 392 191
rect 392 187 395 191
rect 439 188 443 192
rect 495 188 499 192
rect 551 188 555 192
rect 615 188 619 192
rect 655 188 659 192
rect 687 189 691 193
rect 111 171 115 175
rect 151 173 155 177
rect 199 173 203 177
rect 255 173 259 177
rect 311 173 315 177
rect 367 173 371 177
rect 423 173 427 177
rect 479 173 483 177
rect 535 173 539 177
rect 599 173 603 177
rect 639 173 643 177
rect 179 159 183 163
rect 379 167 380 171
rect 380 167 383 171
rect 447 167 448 171
rect 448 167 451 171
rect 487 163 488 167
rect 488 163 491 167
rect 527 167 531 171
rect 111 141 115 145
rect 151 139 155 143
rect 191 139 195 143
rect 231 139 235 143
rect 271 139 275 143
rect 311 139 315 143
rect 351 139 355 143
rect 391 139 395 143
rect 431 139 435 143
rect 471 139 475 143
rect 519 139 523 143
rect 559 139 563 143
rect 495 131 499 135
rect 687 171 691 175
rect 599 139 603 143
rect 639 139 643 143
rect 687 141 691 145
rect 111 123 115 127
rect 167 124 171 128
rect 207 124 211 128
rect 247 124 251 128
rect 287 124 291 128
rect 327 124 331 128
rect 367 124 371 128
rect 407 124 411 128
rect 447 124 451 128
rect 487 124 491 128
rect 535 124 539 128
rect 575 124 579 128
rect 615 124 619 128
rect 655 124 659 128
rect 687 123 691 127
<< m3 >>
rect 111 782 115 783
rect 111 777 115 778
rect 151 782 155 783
rect 151 777 155 778
rect 191 782 195 783
rect 231 782 235 783
rect 191 777 195 778
rect 222 779 228 780
rect 112 762 114 777
rect 110 761 116 762
rect 152 761 154 777
rect 192 761 194 777
rect 222 775 223 779
rect 227 775 228 779
rect 231 777 235 778
rect 271 782 275 783
rect 311 782 315 783
rect 271 777 275 778
rect 278 779 284 780
rect 222 774 228 775
rect 110 757 111 761
rect 115 757 116 761
rect 110 756 116 757
rect 150 760 156 761
rect 150 756 151 760
rect 155 756 156 760
rect 150 755 156 756
rect 190 760 196 761
rect 190 756 191 760
rect 195 756 196 760
rect 190 755 196 756
rect 134 745 140 746
rect 110 743 116 744
rect 110 739 111 743
rect 115 739 116 743
rect 134 741 135 745
rect 139 741 140 745
rect 174 745 180 746
rect 174 741 175 745
rect 179 741 180 745
rect 214 745 220 746
rect 214 741 215 745
rect 219 741 220 745
rect 134 740 140 741
rect 143 740 147 741
rect 174 740 180 741
rect 199 740 203 741
rect 214 740 220 741
rect 224 740 226 774
rect 232 761 234 777
rect 272 761 274 777
rect 278 775 279 779
rect 283 775 284 779
rect 311 777 315 778
rect 351 782 355 783
rect 351 777 355 778
rect 391 782 395 783
rect 391 777 395 778
rect 431 782 435 783
rect 431 777 435 778
rect 687 782 691 783
rect 687 777 691 778
rect 278 774 284 775
rect 230 760 236 761
rect 230 756 231 760
rect 235 756 236 760
rect 230 755 236 756
rect 270 760 276 761
rect 280 760 282 774
rect 312 761 314 777
rect 352 761 354 777
rect 392 761 394 777
rect 432 761 434 777
rect 688 762 690 777
rect 686 761 692 762
rect 310 760 316 761
rect 270 756 271 760
rect 275 756 276 760
rect 270 755 276 756
rect 278 759 284 760
rect 278 755 279 759
rect 283 755 284 759
rect 310 756 311 760
rect 315 756 316 760
rect 310 755 316 756
rect 350 760 356 761
rect 350 756 351 760
rect 355 756 356 760
rect 350 755 356 756
rect 390 760 396 761
rect 390 756 391 760
rect 395 756 396 760
rect 390 755 396 756
rect 430 760 436 761
rect 430 756 431 760
rect 435 756 436 760
rect 686 757 687 761
rect 691 757 692 761
rect 686 756 692 757
rect 430 755 436 756
rect 278 754 284 755
rect 254 745 260 746
rect 254 741 255 745
rect 259 741 260 745
rect 254 740 260 741
rect 294 745 300 746
rect 294 741 295 745
rect 299 741 300 745
rect 334 745 340 746
rect 334 741 335 745
rect 339 741 340 745
rect 374 745 380 746
rect 374 741 375 745
rect 379 741 380 745
rect 294 740 300 741
rect 307 740 311 741
rect 334 740 340 741
rect 355 740 359 741
rect 374 740 380 741
rect 414 745 420 746
rect 414 741 415 745
rect 419 741 420 745
rect 414 740 420 741
rect 686 743 692 744
rect 110 738 116 739
rect 112 731 114 738
rect 136 731 138 740
rect 142 735 143 740
rect 147 735 148 740
rect 142 734 148 735
rect 176 731 178 740
rect 198 735 199 740
rect 203 735 204 740
rect 198 734 204 735
rect 216 731 218 740
rect 222 739 228 740
rect 222 735 223 739
rect 227 735 228 739
rect 222 734 228 735
rect 256 731 258 740
rect 296 731 298 740
rect 306 735 307 740
rect 311 735 312 740
rect 306 734 312 735
rect 336 731 338 740
rect 354 735 355 740
rect 359 735 360 740
rect 354 734 360 735
rect 376 731 378 740
rect 398 739 404 740
rect 398 735 399 739
rect 403 735 404 739
rect 398 734 404 735
rect 111 730 115 731
rect 111 725 115 726
rect 135 730 139 731
rect 135 725 139 726
rect 175 730 179 731
rect 175 725 179 726
rect 215 730 219 731
rect 215 725 219 726
rect 255 730 259 731
rect 255 725 259 726
rect 295 730 299 731
rect 295 725 299 726
rect 335 730 339 731
rect 335 725 339 726
rect 375 730 379 731
rect 375 725 379 726
rect 112 718 114 725
rect 110 717 116 718
rect 110 713 111 717
rect 115 713 116 717
rect 136 716 138 725
rect 176 716 178 725
rect 216 716 218 725
rect 256 716 258 725
rect 296 716 298 725
rect 336 716 338 725
rect 400 724 402 734
rect 416 731 418 740
rect 686 739 687 743
rect 691 739 692 743
rect 686 738 692 739
rect 688 731 690 738
rect 415 730 419 731
rect 415 725 419 726
rect 687 730 691 731
rect 687 725 691 726
rect 398 723 404 724
rect 398 719 399 723
rect 403 719 404 723
rect 398 718 404 719
rect 688 718 690 725
rect 686 717 692 718
rect 110 712 116 713
rect 134 715 140 716
rect 134 711 135 715
rect 139 711 140 715
rect 134 710 140 711
rect 174 715 180 716
rect 174 711 175 715
rect 179 711 180 715
rect 174 710 180 711
rect 214 715 220 716
rect 214 711 215 715
rect 219 711 220 715
rect 214 710 220 711
rect 254 715 260 716
rect 254 711 255 715
rect 259 711 260 715
rect 254 710 260 711
rect 294 715 300 716
rect 294 711 295 715
rect 299 711 300 715
rect 294 710 300 711
rect 334 715 340 716
rect 334 711 335 715
rect 339 711 340 715
rect 686 713 687 717
rect 691 713 692 717
rect 686 712 692 713
rect 334 710 340 711
rect 142 703 148 704
rect 110 699 116 700
rect 110 695 111 699
rect 115 695 116 699
rect 142 699 143 703
rect 147 699 148 703
rect 142 698 148 699
rect 150 700 156 701
rect 110 694 116 695
rect 112 671 114 694
rect 111 670 115 671
rect 111 665 115 666
rect 112 650 114 665
rect 110 649 116 650
rect 110 645 111 649
rect 115 645 116 649
rect 110 644 116 645
rect 134 633 140 634
rect 110 631 116 632
rect 110 627 111 631
rect 115 627 116 631
rect 134 629 135 633
rect 139 629 140 633
rect 134 628 140 629
rect 144 628 146 698
rect 150 696 151 700
rect 155 696 156 700
rect 150 695 156 696
rect 190 700 196 701
rect 190 696 191 700
rect 195 696 196 700
rect 190 695 196 696
rect 230 700 236 701
rect 230 696 231 700
rect 235 696 236 700
rect 230 695 236 696
rect 270 700 276 701
rect 270 696 271 700
rect 275 696 276 700
rect 270 695 276 696
rect 310 700 316 701
rect 310 696 311 700
rect 315 696 316 700
rect 310 695 316 696
rect 350 700 356 701
rect 350 696 351 700
rect 355 696 356 700
rect 350 695 356 696
rect 686 699 692 700
rect 686 695 687 699
rect 691 695 692 699
rect 152 671 154 695
rect 192 671 194 695
rect 232 671 234 695
rect 272 671 274 695
rect 312 671 314 695
rect 352 671 354 695
rect 686 694 692 695
rect 688 671 690 694
rect 151 670 155 671
rect 151 665 155 666
rect 191 670 195 671
rect 191 665 195 666
rect 231 670 235 671
rect 231 665 235 666
rect 271 670 275 671
rect 271 665 275 666
rect 311 670 315 671
rect 311 665 315 666
rect 351 670 355 671
rect 351 665 355 666
rect 687 670 691 671
rect 687 665 691 666
rect 152 649 154 665
rect 192 649 194 665
rect 232 649 234 665
rect 272 649 274 665
rect 312 649 314 665
rect 352 649 354 665
rect 688 650 690 665
rect 686 649 692 650
rect 150 648 156 649
rect 150 644 151 648
rect 155 644 156 648
rect 150 643 156 644
rect 190 648 196 649
rect 190 644 191 648
rect 195 644 196 648
rect 190 643 196 644
rect 230 648 236 649
rect 230 644 231 648
rect 235 644 236 648
rect 230 643 236 644
rect 270 648 276 649
rect 270 644 271 648
rect 275 644 276 648
rect 270 643 276 644
rect 310 648 316 649
rect 310 644 311 648
rect 315 644 316 648
rect 310 643 316 644
rect 350 648 356 649
rect 350 644 351 648
rect 355 644 356 648
rect 686 645 687 649
rect 691 645 692 649
rect 686 644 692 645
rect 350 643 356 644
rect 174 633 180 634
rect 174 629 175 633
rect 179 629 180 633
rect 174 628 180 629
rect 214 633 220 634
rect 214 629 215 633
rect 219 629 220 633
rect 214 628 220 629
rect 254 633 260 634
rect 254 629 255 633
rect 259 629 260 633
rect 254 628 260 629
rect 294 633 300 634
rect 294 629 295 633
rect 299 629 300 633
rect 294 628 300 629
rect 334 633 340 634
rect 334 629 335 633
rect 339 629 340 633
rect 334 628 340 629
rect 686 631 692 632
rect 110 626 116 627
rect 112 611 114 626
rect 136 611 138 628
rect 142 627 148 628
rect 142 623 143 627
rect 147 623 148 627
rect 142 622 148 623
rect 176 611 178 628
rect 216 611 218 628
rect 256 611 258 628
rect 296 611 298 628
rect 336 611 338 628
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 688 611 690 626
rect 111 610 115 611
rect 111 605 115 606
rect 135 610 139 611
rect 135 605 139 606
rect 175 610 179 611
rect 175 605 179 606
rect 215 610 219 611
rect 215 605 219 606
rect 255 610 259 611
rect 255 605 259 606
rect 295 610 299 611
rect 295 605 299 606
rect 335 610 339 611
rect 335 605 339 606
rect 687 610 691 611
rect 687 605 691 606
rect 112 598 114 605
rect 110 597 116 598
rect 110 593 111 597
rect 115 593 116 597
rect 136 596 138 605
rect 176 596 178 605
rect 216 596 218 605
rect 256 596 258 605
rect 296 596 298 605
rect 688 598 690 605
rect 686 597 692 598
rect 110 592 116 593
rect 134 595 140 596
rect 134 591 135 595
rect 139 591 140 595
rect 134 590 140 591
rect 174 595 180 596
rect 174 591 175 595
rect 179 591 180 595
rect 174 590 180 591
rect 214 595 220 596
rect 214 591 215 595
rect 219 591 220 595
rect 214 590 220 591
rect 254 595 260 596
rect 254 591 255 595
rect 259 591 260 595
rect 254 590 260 591
rect 294 595 300 596
rect 294 591 295 595
rect 299 591 300 595
rect 686 593 687 597
rect 691 593 692 597
rect 686 592 692 593
rect 294 590 300 591
rect 142 583 148 584
rect 110 579 116 580
rect 110 575 111 579
rect 115 575 116 579
rect 142 579 143 583
rect 147 579 148 583
rect 142 578 148 579
rect 150 580 156 581
rect 110 574 116 575
rect 112 555 114 574
rect 111 554 115 555
rect 111 549 115 550
rect 112 534 114 549
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 134 517 140 518
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 134 513 135 517
rect 139 513 140 517
rect 134 512 140 513
rect 144 512 146 578
rect 150 576 151 580
rect 155 576 156 580
rect 150 575 156 576
rect 190 580 196 581
rect 190 576 191 580
rect 195 576 196 580
rect 190 575 196 576
rect 230 580 236 581
rect 230 576 231 580
rect 235 576 236 580
rect 230 575 236 576
rect 270 580 276 581
rect 270 576 271 580
rect 275 576 276 580
rect 270 575 276 576
rect 310 580 316 581
rect 310 576 311 580
rect 315 576 316 580
rect 310 575 316 576
rect 686 579 692 580
rect 686 575 687 579
rect 691 575 692 579
rect 152 555 154 575
rect 192 555 194 575
rect 232 555 234 575
rect 272 555 274 575
rect 312 555 314 575
rect 686 574 692 575
rect 688 555 690 574
rect 151 554 155 555
rect 151 549 155 550
rect 191 554 195 555
rect 191 549 195 550
rect 231 554 235 555
rect 231 549 235 550
rect 271 554 275 555
rect 271 549 275 550
rect 311 554 315 555
rect 311 549 315 550
rect 351 554 355 555
rect 351 549 355 550
rect 687 554 691 555
rect 687 549 691 550
rect 152 533 154 549
rect 192 533 194 549
rect 232 533 234 549
rect 272 533 274 549
rect 312 533 314 549
rect 352 533 354 549
rect 688 534 690 549
rect 686 533 692 534
rect 150 532 156 533
rect 150 528 151 532
rect 155 528 156 532
rect 150 527 156 528
rect 190 532 196 533
rect 190 528 191 532
rect 195 528 196 532
rect 190 527 196 528
rect 230 532 236 533
rect 230 528 231 532
rect 235 528 236 532
rect 230 527 236 528
rect 270 532 276 533
rect 270 528 271 532
rect 275 528 276 532
rect 270 527 276 528
rect 310 532 316 533
rect 310 528 311 532
rect 315 528 316 532
rect 310 527 316 528
rect 350 532 356 533
rect 350 528 351 532
rect 355 528 356 532
rect 686 529 687 533
rect 691 529 692 533
rect 686 528 692 529
rect 350 527 356 528
rect 174 517 180 518
rect 174 513 175 517
rect 179 513 180 517
rect 174 512 180 513
rect 214 517 220 518
rect 214 513 215 517
rect 219 513 220 517
rect 214 512 220 513
rect 254 517 260 518
rect 254 513 255 517
rect 259 513 260 517
rect 254 512 260 513
rect 294 517 300 518
rect 294 513 295 517
rect 299 513 300 517
rect 294 512 300 513
rect 334 517 340 518
rect 334 513 335 517
rect 339 513 340 517
rect 334 512 340 513
rect 686 515 692 516
rect 110 510 116 511
rect 112 499 114 510
rect 136 499 138 512
rect 142 511 148 512
rect 142 507 143 511
rect 147 507 148 511
rect 142 506 148 507
rect 176 499 178 512
rect 216 499 218 512
rect 256 499 258 512
rect 296 499 298 512
rect 336 499 338 512
rect 686 511 687 515
rect 691 511 692 515
rect 686 510 692 511
rect 688 499 690 510
rect 111 498 115 499
rect 111 493 115 494
rect 135 498 139 499
rect 135 493 139 494
rect 175 498 179 499
rect 175 493 179 494
rect 215 498 219 499
rect 215 493 219 494
rect 255 498 259 499
rect 255 493 259 494
rect 295 498 299 499
rect 295 493 299 494
rect 335 498 339 499
rect 335 493 339 494
rect 375 498 379 499
rect 375 493 379 494
rect 687 498 691 499
rect 687 493 691 494
rect 112 486 114 493
rect 110 485 116 486
rect 110 481 111 485
rect 115 481 116 485
rect 136 484 138 493
rect 176 484 178 493
rect 216 484 218 493
rect 256 484 258 493
rect 296 484 298 493
rect 336 484 338 493
rect 376 484 378 493
rect 688 486 690 493
rect 686 485 692 486
rect 110 480 116 481
rect 134 483 140 484
rect 134 479 135 483
rect 139 479 140 483
rect 134 478 140 479
rect 174 483 180 484
rect 174 479 175 483
rect 179 479 180 483
rect 174 478 180 479
rect 214 483 220 484
rect 214 479 215 483
rect 219 479 220 483
rect 214 478 220 479
rect 254 483 260 484
rect 254 479 255 483
rect 259 479 260 483
rect 254 478 260 479
rect 294 483 300 484
rect 294 479 295 483
rect 299 479 300 483
rect 294 478 300 479
rect 334 483 340 484
rect 334 479 335 483
rect 339 479 340 483
rect 334 478 340 479
rect 374 483 380 484
rect 374 479 375 483
rect 379 479 380 483
rect 686 481 687 485
rect 691 481 692 485
rect 686 480 692 481
rect 374 478 380 479
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 150 468 156 469
rect 110 467 116 468
rect 110 463 111 467
rect 115 463 116 467
rect 150 464 151 468
rect 155 464 156 468
rect 150 463 156 464
rect 190 468 196 469
rect 190 464 191 468
rect 195 464 196 468
rect 190 463 196 464
rect 230 468 236 469
rect 230 464 231 468
rect 235 464 236 468
rect 230 463 236 464
rect 270 468 276 469
rect 270 464 271 468
rect 275 464 276 468
rect 270 463 276 464
rect 110 462 116 463
rect 112 439 114 462
rect 152 439 154 463
rect 192 439 194 463
rect 232 439 234 463
rect 272 439 274 463
rect 111 438 115 439
rect 111 433 115 434
rect 151 438 155 439
rect 151 433 155 434
rect 191 438 195 439
rect 191 433 195 434
rect 231 438 235 439
rect 231 433 235 434
rect 271 438 275 439
rect 271 433 275 434
rect 279 438 283 439
rect 279 433 283 434
rect 112 418 114 433
rect 110 417 116 418
rect 280 417 282 433
rect 110 413 111 417
rect 115 413 116 417
rect 110 412 116 413
rect 278 416 284 417
rect 278 412 279 416
rect 283 412 284 416
rect 278 411 284 412
rect 262 401 268 402
rect 110 399 116 400
rect 110 395 111 399
rect 115 395 116 399
rect 262 397 263 401
rect 267 397 268 401
rect 262 396 268 397
rect 110 394 116 395
rect 112 387 114 394
rect 264 387 266 396
rect 288 388 290 470
rect 310 468 316 469
rect 310 464 311 468
rect 315 464 316 468
rect 310 463 316 464
rect 350 468 356 469
rect 350 464 351 468
rect 355 464 356 468
rect 350 463 356 464
rect 390 468 396 469
rect 390 464 391 468
rect 395 464 396 468
rect 390 463 396 464
rect 686 467 692 468
rect 686 463 687 467
rect 691 463 692 467
rect 312 439 314 463
rect 352 439 354 463
rect 392 439 394 463
rect 686 462 692 463
rect 688 439 690 462
rect 311 438 315 439
rect 311 433 315 434
rect 319 438 323 439
rect 319 433 323 434
rect 351 438 355 439
rect 351 433 355 434
rect 359 438 363 439
rect 359 433 363 434
rect 391 438 395 439
rect 391 433 395 434
rect 407 438 411 439
rect 407 433 411 434
rect 455 438 459 439
rect 455 433 459 434
rect 503 438 507 439
rect 503 433 507 434
rect 551 438 555 439
rect 551 433 555 434
rect 607 438 611 439
rect 607 433 611 434
rect 655 438 659 439
rect 655 433 659 434
rect 687 438 691 439
rect 687 433 691 434
rect 320 417 322 433
rect 360 417 362 433
rect 408 417 410 433
rect 456 417 458 433
rect 504 417 506 433
rect 552 417 554 433
rect 608 417 610 433
rect 656 417 658 433
rect 688 418 690 433
rect 686 417 692 418
rect 318 416 324 417
rect 318 412 319 416
rect 323 412 324 416
rect 318 411 324 412
rect 358 416 364 417
rect 358 412 359 416
rect 363 412 364 416
rect 358 411 364 412
rect 406 416 412 417
rect 406 412 407 416
rect 411 412 412 416
rect 406 411 412 412
rect 454 416 460 417
rect 454 412 455 416
rect 459 412 460 416
rect 454 411 460 412
rect 502 416 508 417
rect 502 412 503 416
rect 507 412 508 416
rect 502 411 508 412
rect 550 416 556 417
rect 550 412 551 416
rect 555 412 556 416
rect 550 411 556 412
rect 606 416 612 417
rect 606 412 607 416
rect 611 412 612 416
rect 606 411 612 412
rect 654 416 660 417
rect 654 412 655 416
rect 659 412 660 416
rect 686 413 687 417
rect 691 413 692 417
rect 686 412 692 413
rect 654 411 660 412
rect 302 401 308 402
rect 302 397 303 401
rect 307 397 308 401
rect 302 396 308 397
rect 342 401 348 402
rect 342 397 343 401
rect 347 397 348 401
rect 342 396 348 397
rect 390 401 396 402
rect 390 397 391 401
rect 395 397 396 401
rect 390 396 396 397
rect 438 401 444 402
rect 438 397 439 401
rect 443 397 444 401
rect 438 396 444 397
rect 486 401 492 402
rect 486 397 487 401
rect 491 397 492 401
rect 486 396 492 397
rect 534 401 540 402
rect 534 397 535 401
rect 539 397 540 401
rect 534 396 540 397
rect 590 401 596 402
rect 590 397 591 401
rect 595 397 596 401
rect 590 396 596 397
rect 638 401 644 402
rect 638 397 639 401
rect 643 397 644 401
rect 638 396 644 397
rect 686 399 692 400
rect 286 387 292 388
rect 304 387 306 396
rect 344 387 346 396
rect 392 387 394 396
rect 440 387 442 396
rect 488 387 490 396
rect 536 387 538 396
rect 592 387 594 396
rect 640 387 642 396
rect 686 395 687 399
rect 691 395 692 399
rect 686 394 692 395
rect 688 387 690 394
rect 111 386 115 387
rect 111 381 115 382
rect 199 386 203 387
rect 239 386 243 387
rect 199 381 203 382
rect 222 383 228 384
rect 112 374 114 381
rect 110 373 116 374
rect 110 369 111 373
rect 115 369 116 373
rect 200 372 202 381
rect 222 379 223 383
rect 227 379 228 383
rect 239 381 243 382
rect 263 386 267 387
rect 263 381 267 382
rect 279 386 283 387
rect 286 383 287 387
rect 291 383 292 387
rect 286 382 292 383
rect 303 386 307 387
rect 279 381 283 382
rect 303 381 307 382
rect 319 386 323 387
rect 319 381 323 382
rect 343 386 347 387
rect 343 381 347 382
rect 359 386 363 387
rect 359 381 363 382
rect 391 386 395 387
rect 391 381 395 382
rect 399 386 403 387
rect 399 381 403 382
rect 439 386 443 387
rect 439 381 443 382
rect 479 386 483 387
rect 479 381 483 382
rect 487 386 491 387
rect 487 381 491 382
rect 519 386 523 387
rect 519 381 523 382
rect 535 386 539 387
rect 535 381 539 382
rect 559 386 563 387
rect 559 381 563 382
rect 591 386 595 387
rect 591 381 595 382
rect 599 386 603 387
rect 599 381 603 382
rect 639 386 643 387
rect 639 381 643 382
rect 687 386 691 387
rect 687 381 691 382
rect 222 378 228 379
rect 110 368 116 369
rect 198 371 204 372
rect 198 367 199 371
rect 203 367 204 371
rect 198 366 204 367
rect 224 364 226 378
rect 240 372 242 381
rect 280 372 282 381
rect 320 372 322 381
rect 360 372 362 381
rect 400 372 402 381
rect 440 372 442 381
rect 446 379 452 380
rect 446 375 447 379
rect 451 375 452 379
rect 446 374 452 375
rect 238 371 244 372
rect 238 367 239 371
rect 243 367 244 371
rect 238 366 244 367
rect 278 371 284 372
rect 278 367 279 371
rect 283 367 284 371
rect 278 366 284 367
rect 318 371 324 372
rect 318 367 319 371
rect 323 367 324 371
rect 318 366 324 367
rect 358 371 364 372
rect 358 367 359 371
rect 363 367 364 371
rect 358 366 364 367
rect 398 371 404 372
rect 398 367 399 371
rect 403 367 404 371
rect 398 366 404 367
rect 438 371 444 372
rect 438 367 439 371
rect 443 367 444 371
rect 438 366 444 367
rect 222 363 228 364
rect 222 359 223 363
rect 227 359 228 363
rect 222 358 228 359
rect 214 356 220 357
rect 110 355 116 356
rect 110 351 111 355
rect 115 351 116 355
rect 214 352 215 356
rect 219 352 220 356
rect 214 351 220 352
rect 254 356 260 357
rect 294 356 300 357
rect 254 352 255 356
rect 259 352 260 356
rect 254 351 260 352
rect 286 355 292 356
rect 286 351 287 355
rect 291 351 292 355
rect 294 352 295 356
rect 299 352 300 356
rect 294 351 300 352
rect 334 356 340 357
rect 334 352 335 356
rect 339 352 340 356
rect 334 351 340 352
rect 374 356 380 357
rect 374 352 375 356
rect 379 352 380 356
rect 374 351 380 352
rect 414 356 420 357
rect 414 352 415 356
rect 419 352 420 356
rect 414 351 420 352
rect 110 350 116 351
rect 112 331 114 350
rect 216 331 218 351
rect 256 331 258 351
rect 286 350 292 351
rect 111 330 115 331
rect 111 325 115 326
rect 215 330 219 331
rect 215 325 219 326
rect 223 330 227 331
rect 223 325 227 326
rect 255 330 259 331
rect 255 325 259 326
rect 263 330 267 331
rect 263 325 267 326
rect 112 310 114 325
rect 110 309 116 310
rect 224 309 226 325
rect 264 309 266 325
rect 110 305 111 309
rect 115 305 116 309
rect 110 304 116 305
rect 222 308 228 309
rect 222 304 223 308
rect 227 304 228 308
rect 222 303 228 304
rect 262 308 268 309
rect 262 304 263 308
rect 267 304 268 308
rect 262 303 268 304
rect 206 293 212 294
rect 110 291 116 292
rect 110 287 111 291
rect 115 287 116 291
rect 206 289 207 293
rect 211 289 212 293
rect 206 288 212 289
rect 246 293 252 294
rect 246 289 247 293
rect 251 289 252 293
rect 246 288 252 289
rect 288 288 290 350
rect 296 331 298 351
rect 336 331 338 351
rect 376 331 378 351
rect 416 331 418 351
rect 448 340 450 374
rect 480 372 482 381
rect 520 372 522 381
rect 560 372 562 381
rect 600 372 602 381
rect 640 372 642 381
rect 688 374 690 381
rect 686 373 692 374
rect 478 371 484 372
rect 478 367 479 371
rect 483 367 484 371
rect 478 366 484 367
rect 518 371 524 372
rect 518 367 519 371
rect 523 367 524 371
rect 518 366 524 367
rect 558 371 564 372
rect 558 367 559 371
rect 563 367 564 371
rect 558 366 564 367
rect 598 371 604 372
rect 598 367 599 371
rect 603 367 604 371
rect 598 366 604 367
rect 638 371 644 372
rect 638 367 639 371
rect 643 367 644 371
rect 686 369 687 373
rect 691 369 692 373
rect 686 368 692 369
rect 638 366 644 367
rect 454 356 460 357
rect 454 352 455 356
rect 459 352 460 356
rect 454 351 460 352
rect 494 356 500 357
rect 494 352 495 356
rect 499 352 500 356
rect 494 351 500 352
rect 534 356 540 357
rect 534 352 535 356
rect 539 352 540 356
rect 534 351 540 352
rect 574 356 580 357
rect 614 356 620 357
rect 574 352 575 356
rect 579 352 580 356
rect 574 351 580 352
rect 598 355 604 356
rect 598 351 599 355
rect 603 351 604 355
rect 614 352 615 356
rect 619 352 620 356
rect 614 351 620 352
rect 654 356 660 357
rect 654 352 655 356
rect 659 352 660 356
rect 654 351 660 352
rect 686 355 692 356
rect 686 351 687 355
rect 691 351 692 355
rect 446 339 452 340
rect 446 335 447 339
rect 451 335 452 339
rect 446 334 452 335
rect 456 331 458 351
rect 486 339 492 340
rect 486 335 487 339
rect 491 335 492 339
rect 486 334 492 335
rect 295 330 299 331
rect 295 325 299 326
rect 311 330 315 331
rect 311 325 315 326
rect 335 330 339 331
rect 335 325 339 326
rect 367 330 371 331
rect 367 325 371 326
rect 375 330 379 331
rect 375 325 379 326
rect 415 330 419 331
rect 415 325 419 326
rect 423 330 427 331
rect 423 325 427 326
rect 455 330 459 331
rect 455 325 459 326
rect 479 330 483 331
rect 479 325 483 326
rect 312 309 314 325
rect 368 309 370 325
rect 424 309 426 325
rect 480 309 482 325
rect 310 308 316 309
rect 310 304 311 308
rect 315 304 316 308
rect 310 303 316 304
rect 366 308 372 309
rect 366 304 367 308
rect 371 304 372 308
rect 366 303 372 304
rect 422 308 428 309
rect 422 304 423 308
rect 427 304 428 308
rect 422 303 428 304
rect 478 308 484 309
rect 488 308 490 334
rect 496 331 498 351
rect 536 331 538 351
rect 576 331 578 351
rect 598 350 604 351
rect 495 330 499 331
rect 495 325 499 326
rect 535 330 539 331
rect 535 325 539 326
rect 543 330 547 331
rect 543 325 547 326
rect 575 330 579 331
rect 575 325 579 326
rect 544 309 546 325
rect 542 308 548 309
rect 478 304 479 308
rect 483 304 484 308
rect 478 303 484 304
rect 486 307 492 308
rect 486 303 487 307
rect 491 303 492 307
rect 542 304 543 308
rect 547 304 548 308
rect 542 303 548 304
rect 486 302 492 303
rect 294 293 300 294
rect 294 289 295 293
rect 299 289 300 293
rect 294 288 300 289
rect 350 293 356 294
rect 350 289 351 293
rect 355 289 356 293
rect 350 288 356 289
rect 406 293 412 294
rect 406 289 407 293
rect 411 289 412 293
rect 406 288 412 289
rect 462 293 468 294
rect 462 289 463 293
rect 467 289 468 293
rect 462 288 468 289
rect 526 293 532 294
rect 526 289 527 293
rect 531 289 532 293
rect 526 288 532 289
rect 590 293 596 294
rect 590 289 591 293
rect 595 289 596 293
rect 590 288 596 289
rect 600 288 602 350
rect 616 331 618 351
rect 656 331 658 351
rect 686 350 692 351
rect 688 331 690 350
rect 607 330 611 331
rect 607 325 611 326
rect 615 330 619 331
rect 615 325 619 326
rect 655 330 659 331
rect 655 325 659 326
rect 687 330 691 331
rect 687 325 691 326
rect 608 309 610 325
rect 656 309 658 325
rect 688 310 690 325
rect 686 309 692 310
rect 606 308 612 309
rect 606 304 607 308
rect 611 304 612 308
rect 606 303 612 304
rect 654 308 660 309
rect 654 304 655 308
rect 659 304 660 308
rect 686 305 687 309
rect 691 305 692 309
rect 686 304 692 305
rect 654 303 660 304
rect 638 293 644 294
rect 638 289 639 293
rect 643 289 644 293
rect 638 288 644 289
rect 686 291 692 292
rect 110 286 116 287
rect 112 275 114 286
rect 208 275 210 288
rect 248 275 250 288
rect 274 287 280 288
rect 274 283 275 287
rect 279 283 280 287
rect 286 287 292 288
rect 286 283 287 287
rect 291 283 292 287
rect 274 282 282 283
rect 286 282 292 283
rect 276 281 282 282
rect 111 274 115 275
rect 111 269 115 270
rect 143 274 147 275
rect 143 269 147 270
rect 207 274 211 275
rect 207 269 211 270
rect 247 274 251 275
rect 247 269 251 270
rect 271 274 275 275
rect 280 272 282 281
rect 296 275 298 288
rect 352 275 354 288
rect 408 275 410 288
rect 464 275 466 288
rect 490 283 496 284
rect 490 279 491 283
rect 495 279 496 283
rect 490 278 496 279
rect 295 274 299 275
rect 271 269 275 270
rect 278 271 284 272
rect 112 262 114 269
rect 110 261 116 262
rect 110 257 111 261
rect 115 257 116 261
rect 144 260 146 269
rect 208 260 210 269
rect 272 260 274 269
rect 278 267 279 271
rect 283 267 284 271
rect 295 269 299 270
rect 335 274 339 275
rect 335 269 339 270
rect 351 274 355 275
rect 351 269 355 270
rect 399 274 403 275
rect 399 269 403 270
rect 407 274 411 275
rect 407 269 411 270
rect 463 274 467 275
rect 463 269 467 270
rect 278 266 284 267
rect 336 260 338 269
rect 390 267 396 268
rect 390 263 391 267
rect 395 263 396 267
rect 390 262 396 263
rect 110 256 116 257
rect 142 259 148 260
rect 142 255 143 259
rect 147 255 148 259
rect 142 254 148 255
rect 206 259 212 260
rect 206 255 207 259
rect 211 255 212 259
rect 206 254 212 255
rect 270 259 276 260
rect 270 255 271 259
rect 275 255 276 259
rect 270 254 276 255
rect 334 259 340 260
rect 334 255 335 259
rect 339 255 340 259
rect 334 254 340 255
rect 158 244 164 245
rect 222 244 228 245
rect 110 243 116 244
rect 110 239 111 243
rect 115 239 116 243
rect 158 240 159 244
rect 163 240 164 244
rect 158 239 164 240
rect 178 243 184 244
rect 178 239 179 243
rect 183 239 184 243
rect 222 240 223 244
rect 227 240 228 244
rect 222 239 228 240
rect 286 244 292 245
rect 286 240 287 244
rect 291 240 292 244
rect 286 239 292 240
rect 350 244 356 245
rect 350 240 351 244
rect 355 240 356 244
rect 350 239 356 240
rect 110 238 116 239
rect 112 215 114 238
rect 160 215 162 239
rect 178 238 184 239
rect 111 214 115 215
rect 111 209 115 210
rect 159 214 163 215
rect 159 209 163 210
rect 167 214 171 215
rect 167 209 171 210
rect 112 194 114 209
rect 110 193 116 194
rect 168 193 170 209
rect 110 189 111 193
rect 115 189 116 193
rect 110 188 116 189
rect 166 192 172 193
rect 166 188 167 192
rect 171 188 172 192
rect 166 187 172 188
rect 150 177 156 178
rect 110 175 116 176
rect 110 171 111 175
rect 115 171 116 175
rect 150 173 151 177
rect 155 173 156 177
rect 150 172 156 173
rect 110 170 116 171
rect 112 159 114 170
rect 152 159 154 172
rect 180 164 182 238
rect 224 215 226 239
rect 288 215 290 239
rect 352 215 354 239
rect 215 214 219 215
rect 215 209 219 210
rect 223 214 227 215
rect 223 209 227 210
rect 271 214 275 215
rect 271 209 275 210
rect 287 214 291 215
rect 287 209 291 210
rect 327 214 331 215
rect 327 209 331 210
rect 351 214 355 215
rect 351 209 355 210
rect 383 214 387 215
rect 383 209 387 210
rect 216 193 218 209
rect 272 193 274 209
rect 328 193 330 209
rect 384 193 386 209
rect 214 192 220 193
rect 214 188 215 192
rect 219 188 220 192
rect 214 187 220 188
rect 270 192 276 193
rect 270 188 271 192
rect 275 188 276 192
rect 270 187 276 188
rect 326 192 332 193
rect 326 188 327 192
rect 331 188 332 192
rect 326 187 332 188
rect 382 192 388 193
rect 392 192 394 262
rect 400 260 402 269
rect 464 260 466 269
rect 492 264 494 278
rect 528 275 530 288
rect 592 275 594 288
rect 598 287 604 288
rect 598 283 599 287
rect 603 283 604 287
rect 598 282 604 283
rect 640 275 642 288
rect 686 287 687 291
rect 691 287 692 291
rect 686 286 692 287
rect 688 275 690 286
rect 527 274 531 275
rect 527 269 531 270
rect 591 274 595 275
rect 591 269 595 270
rect 639 274 643 275
rect 639 269 643 270
rect 687 274 691 275
rect 687 269 691 270
rect 490 263 496 264
rect 398 259 404 260
rect 398 255 399 259
rect 403 255 404 259
rect 398 254 404 255
rect 462 259 468 260
rect 462 255 463 259
rect 467 255 468 259
rect 490 259 491 263
rect 495 259 496 263
rect 528 260 530 269
rect 592 260 594 269
rect 640 260 642 269
rect 688 262 690 269
rect 686 261 692 262
rect 490 258 496 259
rect 526 259 532 260
rect 462 254 468 255
rect 526 255 527 259
rect 531 255 532 259
rect 526 254 532 255
rect 590 259 596 260
rect 590 255 591 259
rect 595 255 596 259
rect 590 254 596 255
rect 638 259 644 260
rect 638 255 639 259
rect 643 255 644 259
rect 686 257 687 261
rect 691 257 692 261
rect 686 256 692 257
rect 638 254 644 255
rect 526 247 532 248
rect 414 244 420 245
rect 414 240 415 244
rect 419 240 420 244
rect 414 239 420 240
rect 478 244 484 245
rect 478 240 479 244
rect 483 240 484 244
rect 526 243 527 247
rect 531 243 532 247
rect 526 242 532 243
rect 542 244 548 245
rect 478 239 484 240
rect 416 215 418 239
rect 480 215 482 239
rect 415 214 419 215
rect 415 209 419 210
rect 439 214 443 215
rect 439 209 443 210
rect 479 214 483 215
rect 479 209 483 210
rect 495 214 499 215
rect 495 209 499 210
rect 440 193 442 209
rect 496 193 498 209
rect 438 192 444 193
rect 382 188 383 192
rect 387 188 388 192
rect 382 187 388 188
rect 390 191 396 192
rect 390 187 391 191
rect 395 187 396 191
rect 438 188 439 192
rect 443 188 444 192
rect 438 187 444 188
rect 494 192 500 193
rect 494 188 495 192
rect 499 188 500 192
rect 494 187 500 188
rect 390 186 396 187
rect 198 177 204 178
rect 198 173 199 177
rect 203 173 204 177
rect 198 172 204 173
rect 254 177 260 178
rect 254 173 255 177
rect 259 173 260 177
rect 254 172 260 173
rect 310 177 316 178
rect 310 173 311 177
rect 315 173 316 177
rect 310 172 316 173
rect 366 177 372 178
rect 366 173 367 177
rect 371 173 372 177
rect 422 177 428 178
rect 422 173 423 177
rect 427 173 428 177
rect 478 177 484 178
rect 478 173 479 177
rect 483 173 484 177
rect 366 172 372 173
rect 379 172 383 173
rect 422 172 428 173
rect 447 172 451 173
rect 478 172 484 173
rect 528 172 530 242
rect 542 240 543 244
rect 547 240 548 244
rect 542 239 548 240
rect 606 244 612 245
rect 606 240 607 244
rect 611 240 612 244
rect 606 239 612 240
rect 654 244 660 245
rect 654 240 655 244
rect 659 240 660 244
rect 654 239 660 240
rect 686 243 692 244
rect 686 239 687 243
rect 691 239 692 243
rect 544 215 546 239
rect 608 215 610 239
rect 656 215 658 239
rect 686 238 692 239
rect 688 215 690 238
rect 543 214 547 215
rect 543 209 547 210
rect 551 214 555 215
rect 551 209 555 210
rect 607 214 611 215
rect 607 209 611 210
rect 615 214 619 215
rect 615 209 619 210
rect 655 214 659 215
rect 655 209 659 210
rect 687 214 691 215
rect 687 209 691 210
rect 552 193 554 209
rect 616 193 618 209
rect 656 193 658 209
rect 688 194 690 209
rect 686 193 692 194
rect 550 192 556 193
rect 550 188 551 192
rect 555 188 556 192
rect 550 187 556 188
rect 614 192 620 193
rect 614 188 615 192
rect 619 188 620 192
rect 614 187 620 188
rect 654 192 660 193
rect 654 188 655 192
rect 659 188 660 192
rect 686 189 687 193
rect 691 189 692 193
rect 686 188 692 189
rect 654 187 660 188
rect 534 177 540 178
rect 534 173 535 177
rect 539 173 540 177
rect 534 172 540 173
rect 598 177 604 178
rect 598 173 599 177
rect 603 173 604 177
rect 598 172 604 173
rect 638 177 644 178
rect 638 173 639 177
rect 643 173 644 177
rect 638 172 644 173
rect 686 175 692 176
rect 178 163 184 164
rect 178 159 179 163
rect 183 159 184 163
rect 200 159 202 172
rect 256 159 258 172
rect 312 159 314 172
rect 368 159 370 172
rect 378 167 379 172
rect 383 167 384 172
rect 378 166 384 167
rect 424 159 426 172
rect 446 167 447 172
rect 451 167 452 172
rect 446 166 452 167
rect 480 159 482 172
rect 526 171 532 172
rect 486 167 492 168
rect 486 163 487 167
rect 491 163 492 167
rect 526 167 527 171
rect 531 167 532 171
rect 526 166 532 167
rect 486 162 492 163
rect 111 158 115 159
rect 111 153 115 154
rect 151 158 155 159
rect 178 158 184 159
rect 191 158 195 159
rect 151 153 155 154
rect 191 153 195 154
rect 199 158 203 159
rect 199 153 203 154
rect 231 158 235 159
rect 231 153 235 154
rect 255 158 259 159
rect 255 153 259 154
rect 271 158 275 159
rect 271 153 275 154
rect 311 158 315 159
rect 311 153 315 154
rect 351 158 355 159
rect 351 153 355 154
rect 367 158 371 159
rect 367 153 371 154
rect 391 158 395 159
rect 391 153 395 154
rect 423 158 427 159
rect 423 153 427 154
rect 431 158 435 159
rect 431 153 435 154
rect 471 158 475 159
rect 471 153 475 154
rect 479 158 483 159
rect 479 153 483 154
rect 112 146 114 153
rect 110 145 116 146
rect 110 141 111 145
rect 115 141 116 145
rect 152 144 154 153
rect 192 144 194 153
rect 232 144 234 153
rect 272 144 274 153
rect 312 144 314 153
rect 352 144 354 153
rect 392 144 394 153
rect 432 144 434 153
rect 472 144 474 153
rect 488 147 490 162
rect 536 159 538 172
rect 600 159 602 172
rect 640 159 642 172
rect 686 171 687 175
rect 691 171 692 175
rect 686 170 692 171
rect 688 159 690 170
rect 519 158 523 159
rect 519 153 523 154
rect 535 158 539 159
rect 535 153 539 154
rect 559 158 563 159
rect 559 153 563 154
rect 599 158 603 159
rect 599 153 603 154
rect 639 158 643 159
rect 639 153 643 154
rect 687 158 691 159
rect 687 153 691 154
rect 488 145 498 147
rect 110 140 116 141
rect 150 143 156 144
rect 150 139 151 143
rect 155 139 156 143
rect 150 138 156 139
rect 190 143 196 144
rect 190 139 191 143
rect 195 139 196 143
rect 190 138 196 139
rect 230 143 236 144
rect 230 139 231 143
rect 235 139 236 143
rect 230 138 236 139
rect 270 143 276 144
rect 270 139 271 143
rect 275 139 276 143
rect 270 138 276 139
rect 310 143 316 144
rect 310 139 311 143
rect 315 139 316 143
rect 310 138 316 139
rect 350 143 356 144
rect 350 139 351 143
rect 355 139 356 143
rect 350 138 356 139
rect 390 143 396 144
rect 390 139 391 143
rect 395 139 396 143
rect 390 138 396 139
rect 430 143 436 144
rect 430 139 431 143
rect 435 139 436 143
rect 430 138 436 139
rect 470 143 476 144
rect 470 139 471 143
rect 475 139 476 143
rect 470 138 476 139
rect 496 136 498 145
rect 520 144 522 153
rect 560 144 562 153
rect 600 144 602 153
rect 640 144 642 153
rect 688 146 690 153
rect 686 145 692 146
rect 518 143 524 144
rect 518 139 519 143
rect 523 139 524 143
rect 518 138 524 139
rect 558 143 564 144
rect 558 139 559 143
rect 563 139 564 143
rect 558 138 564 139
rect 598 143 604 144
rect 598 139 599 143
rect 603 139 604 143
rect 598 138 604 139
rect 638 143 644 144
rect 638 139 639 143
rect 643 139 644 143
rect 686 141 687 145
rect 691 141 692 145
rect 686 140 692 141
rect 638 138 644 139
rect 494 135 500 136
rect 494 131 495 135
rect 499 131 500 135
rect 494 130 500 131
rect 166 128 172 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 166 124 167 128
rect 171 124 172 128
rect 166 123 172 124
rect 206 128 212 129
rect 206 124 207 128
rect 211 124 212 128
rect 206 123 212 124
rect 246 128 252 129
rect 246 124 247 128
rect 251 124 252 128
rect 246 123 252 124
rect 286 128 292 129
rect 286 124 287 128
rect 291 124 292 128
rect 286 123 292 124
rect 326 128 332 129
rect 326 124 327 128
rect 331 124 332 128
rect 326 123 332 124
rect 366 128 372 129
rect 366 124 367 128
rect 371 124 372 128
rect 366 123 372 124
rect 406 128 412 129
rect 406 124 407 128
rect 411 124 412 128
rect 406 123 412 124
rect 446 128 452 129
rect 446 124 447 128
rect 451 124 452 128
rect 446 123 452 124
rect 486 128 492 129
rect 486 124 487 128
rect 491 124 492 128
rect 486 123 492 124
rect 534 128 540 129
rect 534 124 535 128
rect 539 124 540 128
rect 534 123 540 124
rect 574 128 580 129
rect 574 124 575 128
rect 579 124 580 128
rect 574 123 580 124
rect 614 128 620 129
rect 614 124 615 128
rect 619 124 620 128
rect 614 123 620 124
rect 654 128 660 129
rect 654 124 655 128
rect 659 124 660 128
rect 654 123 660 124
rect 686 127 692 128
rect 686 123 687 127
rect 691 123 692 127
rect 110 122 116 123
rect 112 107 114 122
rect 168 107 170 123
rect 208 107 210 123
rect 248 107 250 123
rect 288 107 290 123
rect 328 107 330 123
rect 368 107 370 123
rect 408 107 410 123
rect 448 107 450 123
rect 488 107 490 123
rect 536 107 538 123
rect 576 107 578 123
rect 616 107 618 123
rect 656 107 658 123
rect 686 122 692 123
rect 688 107 690 122
rect 111 106 115 107
rect 111 101 115 102
rect 167 106 171 107
rect 167 101 171 102
rect 207 106 211 107
rect 207 101 211 102
rect 247 106 251 107
rect 247 101 251 102
rect 287 106 291 107
rect 287 101 291 102
rect 327 106 331 107
rect 327 101 331 102
rect 367 106 371 107
rect 367 101 371 102
rect 407 106 411 107
rect 407 101 411 102
rect 447 106 451 107
rect 447 101 451 102
rect 487 106 491 107
rect 487 101 491 102
rect 535 106 539 107
rect 535 101 539 102
rect 575 106 579 107
rect 575 101 579 102
rect 615 106 619 107
rect 615 101 619 102
rect 655 106 659 107
rect 655 101 659 102
rect 687 106 691 107
rect 687 101 691 102
<< m4c >>
rect 111 778 115 782
rect 151 778 155 782
rect 191 778 195 782
rect 231 778 235 782
rect 271 778 275 782
rect 311 778 315 782
rect 351 778 355 782
rect 391 778 395 782
rect 431 778 435 782
rect 687 778 691 782
rect 143 739 147 740
rect 143 736 147 739
rect 199 739 203 740
rect 199 736 203 739
rect 307 739 311 740
rect 307 736 311 739
rect 355 739 359 740
rect 355 736 359 739
rect 111 726 115 730
rect 135 726 139 730
rect 175 726 179 730
rect 215 726 219 730
rect 255 726 259 730
rect 295 726 299 730
rect 335 726 339 730
rect 375 726 379 730
rect 415 726 419 730
rect 687 726 691 730
rect 111 666 115 670
rect 151 666 155 670
rect 191 666 195 670
rect 231 666 235 670
rect 271 666 275 670
rect 311 666 315 670
rect 351 666 355 670
rect 687 666 691 670
rect 111 606 115 610
rect 135 606 139 610
rect 175 606 179 610
rect 215 606 219 610
rect 255 606 259 610
rect 295 606 299 610
rect 335 606 339 610
rect 687 606 691 610
rect 111 550 115 554
rect 151 550 155 554
rect 191 550 195 554
rect 231 550 235 554
rect 271 550 275 554
rect 311 550 315 554
rect 351 550 355 554
rect 687 550 691 554
rect 111 494 115 498
rect 135 494 139 498
rect 175 494 179 498
rect 215 494 219 498
rect 255 494 259 498
rect 295 494 299 498
rect 335 494 339 498
rect 375 494 379 498
rect 687 494 691 498
rect 111 434 115 438
rect 151 434 155 438
rect 191 434 195 438
rect 231 434 235 438
rect 271 434 275 438
rect 279 434 283 438
rect 311 434 315 438
rect 319 434 323 438
rect 351 434 355 438
rect 359 434 363 438
rect 391 434 395 438
rect 407 434 411 438
rect 455 434 459 438
rect 503 434 507 438
rect 551 434 555 438
rect 607 434 611 438
rect 655 434 659 438
rect 687 434 691 438
rect 111 382 115 386
rect 199 382 203 386
rect 239 382 243 386
rect 263 382 267 386
rect 279 382 283 386
rect 303 382 307 386
rect 319 382 323 386
rect 343 382 347 386
rect 359 382 363 386
rect 391 382 395 386
rect 399 382 403 386
rect 439 382 443 386
rect 479 382 483 386
rect 487 382 491 386
rect 519 382 523 386
rect 535 382 539 386
rect 559 382 563 386
rect 591 382 595 386
rect 599 382 603 386
rect 639 382 643 386
rect 687 382 691 386
rect 111 326 115 330
rect 215 326 219 330
rect 223 326 227 330
rect 255 326 259 330
rect 263 326 267 330
rect 295 326 299 330
rect 311 326 315 330
rect 335 326 339 330
rect 367 326 371 330
rect 375 326 379 330
rect 415 326 419 330
rect 423 326 427 330
rect 455 326 459 330
rect 479 326 483 330
rect 495 326 499 330
rect 535 326 539 330
rect 543 326 547 330
rect 575 326 579 330
rect 607 326 611 330
rect 615 326 619 330
rect 655 326 659 330
rect 687 326 691 330
rect 111 270 115 274
rect 143 270 147 274
rect 207 270 211 274
rect 247 270 251 274
rect 271 270 275 274
rect 295 270 299 274
rect 335 270 339 274
rect 351 270 355 274
rect 399 270 403 274
rect 407 270 411 274
rect 463 270 467 274
rect 111 210 115 214
rect 159 210 163 214
rect 167 210 171 214
rect 215 210 219 214
rect 223 210 227 214
rect 271 210 275 214
rect 287 210 291 214
rect 327 210 331 214
rect 351 210 355 214
rect 383 210 387 214
rect 527 270 531 274
rect 591 270 595 274
rect 639 270 643 274
rect 687 270 691 274
rect 415 210 419 214
rect 439 210 443 214
rect 479 210 483 214
rect 495 210 499 214
rect 543 210 547 214
rect 551 210 555 214
rect 607 210 611 214
rect 615 210 619 214
rect 655 210 659 214
rect 687 210 691 214
rect 379 171 383 172
rect 379 168 383 171
rect 447 171 451 172
rect 447 168 451 171
rect 111 154 115 158
rect 151 154 155 158
rect 191 154 195 158
rect 199 154 203 158
rect 231 154 235 158
rect 255 154 259 158
rect 271 154 275 158
rect 311 154 315 158
rect 351 154 355 158
rect 367 154 371 158
rect 391 154 395 158
rect 423 154 427 158
rect 431 154 435 158
rect 471 154 475 158
rect 479 154 483 158
rect 519 154 523 158
rect 535 154 539 158
rect 559 154 563 158
rect 599 154 603 158
rect 639 154 643 158
rect 687 154 691 158
rect 111 102 115 106
rect 167 102 171 106
rect 207 102 211 106
rect 247 102 251 106
rect 287 102 291 106
rect 327 102 331 106
rect 367 102 371 106
rect 407 102 411 106
rect 447 102 451 106
rect 487 102 491 106
rect 535 102 539 106
rect 575 102 579 106
rect 615 102 619 106
rect 655 102 659 106
rect 687 102 691 106
<< m4 >>
rect 84 777 85 783
rect 91 782 711 783
rect 91 778 111 782
rect 115 778 151 782
rect 155 778 191 782
rect 195 778 231 782
rect 235 778 271 782
rect 275 778 311 782
rect 315 778 351 782
rect 355 778 391 782
rect 395 778 431 782
rect 435 778 687 782
rect 691 778 711 782
rect 91 777 711 778
rect 717 777 718 783
rect 142 740 148 741
rect 198 740 204 741
rect 142 736 143 740
rect 147 736 199 740
rect 203 736 204 740
rect 142 735 148 736
rect 198 735 204 736
rect 306 740 312 741
rect 354 740 360 741
rect 306 736 307 740
rect 311 736 355 740
rect 359 736 360 740
rect 306 735 312 736
rect 354 735 360 736
rect 96 725 97 731
rect 103 730 723 731
rect 103 726 111 730
rect 115 726 135 730
rect 139 726 175 730
rect 179 726 215 730
rect 219 726 255 730
rect 259 726 295 730
rect 299 726 335 730
rect 339 726 375 730
rect 379 726 415 730
rect 419 726 687 730
rect 691 726 723 730
rect 103 725 723 726
rect 729 725 730 731
rect 84 665 85 671
rect 91 670 711 671
rect 91 666 111 670
rect 115 666 151 670
rect 155 666 191 670
rect 195 666 231 670
rect 235 666 271 670
rect 275 666 311 670
rect 315 666 351 670
rect 355 666 687 670
rect 691 666 711 670
rect 91 665 711 666
rect 717 665 718 671
rect 96 605 97 611
rect 103 610 723 611
rect 103 606 111 610
rect 115 606 135 610
rect 139 606 175 610
rect 179 606 215 610
rect 219 606 255 610
rect 259 606 295 610
rect 299 606 335 610
rect 339 606 687 610
rect 691 606 723 610
rect 103 605 723 606
rect 729 605 730 611
rect 84 549 85 555
rect 91 554 711 555
rect 91 550 111 554
rect 115 550 151 554
rect 155 550 191 554
rect 195 550 231 554
rect 235 550 271 554
rect 275 550 311 554
rect 315 550 351 554
rect 355 550 687 554
rect 691 550 711 554
rect 91 549 711 550
rect 717 549 718 555
rect 96 493 97 499
rect 103 498 723 499
rect 103 494 111 498
rect 115 494 135 498
rect 139 494 175 498
rect 179 494 215 498
rect 219 494 255 498
rect 259 494 295 498
rect 299 494 335 498
rect 339 494 375 498
rect 379 494 687 498
rect 691 494 723 498
rect 103 493 723 494
rect 729 493 730 499
rect 84 433 85 439
rect 91 438 711 439
rect 91 434 111 438
rect 115 434 151 438
rect 155 434 191 438
rect 195 434 231 438
rect 235 434 271 438
rect 275 434 279 438
rect 283 434 311 438
rect 315 434 319 438
rect 323 434 351 438
rect 355 434 359 438
rect 363 434 391 438
rect 395 434 407 438
rect 411 434 455 438
rect 459 434 503 438
rect 507 434 551 438
rect 555 434 607 438
rect 611 434 655 438
rect 659 434 687 438
rect 691 434 711 438
rect 91 433 711 434
rect 717 433 718 439
rect 96 381 97 387
rect 103 386 723 387
rect 103 382 111 386
rect 115 382 199 386
rect 203 382 239 386
rect 243 382 263 386
rect 267 382 279 386
rect 283 382 303 386
rect 307 382 319 386
rect 323 382 343 386
rect 347 382 359 386
rect 363 382 391 386
rect 395 382 399 386
rect 403 382 439 386
rect 443 382 479 386
rect 483 382 487 386
rect 491 382 519 386
rect 523 382 535 386
rect 539 382 559 386
rect 563 382 591 386
rect 595 382 599 386
rect 603 382 639 386
rect 643 382 687 386
rect 691 382 723 386
rect 103 381 723 382
rect 729 381 730 387
rect 84 325 85 331
rect 91 330 711 331
rect 91 326 111 330
rect 115 326 215 330
rect 219 326 223 330
rect 227 326 255 330
rect 259 326 263 330
rect 267 326 295 330
rect 299 326 311 330
rect 315 326 335 330
rect 339 326 367 330
rect 371 326 375 330
rect 379 326 415 330
rect 419 326 423 330
rect 427 326 455 330
rect 459 326 479 330
rect 483 326 495 330
rect 499 326 535 330
rect 539 326 543 330
rect 547 326 575 330
rect 579 326 607 330
rect 611 326 615 330
rect 619 326 655 330
rect 659 326 687 330
rect 691 326 711 330
rect 91 325 711 326
rect 717 325 718 331
rect 96 269 97 275
rect 103 274 723 275
rect 103 270 111 274
rect 115 270 143 274
rect 147 270 207 274
rect 211 270 247 274
rect 251 270 271 274
rect 275 270 295 274
rect 299 270 335 274
rect 339 270 351 274
rect 355 270 399 274
rect 403 270 407 274
rect 411 270 463 274
rect 467 270 527 274
rect 531 270 591 274
rect 595 270 639 274
rect 643 270 687 274
rect 691 270 723 274
rect 103 269 723 270
rect 729 269 730 275
rect 84 209 85 215
rect 91 214 711 215
rect 91 210 111 214
rect 115 210 159 214
rect 163 210 167 214
rect 171 210 215 214
rect 219 210 223 214
rect 227 210 271 214
rect 275 210 287 214
rect 291 210 327 214
rect 331 210 351 214
rect 355 210 383 214
rect 387 210 415 214
rect 419 210 439 214
rect 443 210 479 214
rect 483 210 495 214
rect 499 210 543 214
rect 547 210 551 214
rect 555 210 607 214
rect 611 210 615 214
rect 619 210 655 214
rect 659 210 687 214
rect 691 210 711 214
rect 91 209 711 210
rect 717 209 718 215
rect 378 172 384 173
rect 446 172 452 173
rect 378 168 379 172
rect 383 168 447 172
rect 451 168 452 172
rect 378 167 384 168
rect 446 167 452 168
rect 96 153 97 159
rect 103 158 723 159
rect 103 154 111 158
rect 115 154 151 158
rect 155 154 191 158
rect 195 154 199 158
rect 203 154 231 158
rect 235 154 255 158
rect 259 154 271 158
rect 275 154 311 158
rect 315 154 351 158
rect 355 154 367 158
rect 371 154 391 158
rect 395 154 423 158
rect 427 154 431 158
rect 435 154 471 158
rect 475 154 479 158
rect 483 154 519 158
rect 523 154 535 158
rect 539 154 559 158
rect 563 154 599 158
rect 603 154 639 158
rect 643 154 687 158
rect 691 154 723 158
rect 103 153 723 154
rect 729 153 730 159
rect 84 101 85 107
rect 91 106 711 107
rect 91 102 111 106
rect 115 102 167 106
rect 171 102 207 106
rect 211 102 247 106
rect 251 102 287 106
rect 291 102 327 106
rect 331 102 367 106
rect 371 102 407 106
rect 411 102 447 106
rect 451 102 487 106
rect 491 102 535 106
rect 539 102 575 106
rect 579 102 615 106
rect 619 102 655 106
rect 659 102 687 106
rect 691 102 711 106
rect 91 101 711 102
rect 717 101 718 107
<< m5c >>
rect 85 777 91 783
rect 711 777 717 783
rect 97 725 103 731
rect 723 725 729 731
rect 85 665 91 671
rect 711 665 717 671
rect 97 605 103 611
rect 723 605 729 611
rect 85 549 91 555
rect 711 549 717 555
rect 97 493 103 499
rect 723 493 729 499
rect 85 433 91 439
rect 711 433 717 439
rect 97 381 103 387
rect 723 381 729 387
rect 85 325 91 331
rect 711 325 717 331
rect 97 269 103 275
rect 723 269 729 275
rect 85 209 91 215
rect 711 209 717 215
rect 97 153 103 159
rect 723 153 729 159
rect 85 101 91 107
rect 711 101 717 107
<< m5 >>
rect 84 783 92 792
rect 84 777 85 783
rect 91 777 92 783
rect 84 671 92 777
rect 84 665 85 671
rect 91 665 92 671
rect 84 555 92 665
rect 84 549 85 555
rect 91 549 92 555
rect 84 439 92 549
rect 84 433 85 439
rect 91 433 92 439
rect 84 331 92 433
rect 84 325 85 331
rect 91 325 92 331
rect 84 215 92 325
rect 84 209 85 215
rect 91 209 92 215
rect 84 107 92 209
rect 84 101 85 107
rect 91 101 92 107
rect 84 72 92 101
rect 96 731 104 792
rect 96 725 97 731
rect 103 725 104 731
rect 96 611 104 725
rect 96 605 97 611
rect 103 605 104 611
rect 96 499 104 605
rect 96 493 97 499
rect 103 493 104 499
rect 96 387 104 493
rect 96 381 97 387
rect 103 381 104 387
rect 96 275 104 381
rect 96 269 97 275
rect 103 269 104 275
rect 96 159 104 269
rect 96 153 97 159
rect 103 153 104 159
rect 96 72 104 153
rect 710 783 718 792
rect 710 777 711 783
rect 717 777 718 783
rect 710 671 718 777
rect 710 665 711 671
rect 717 665 718 671
rect 710 555 718 665
rect 710 549 711 555
rect 717 549 718 555
rect 710 439 718 549
rect 710 433 711 439
rect 717 433 718 439
rect 710 331 718 433
rect 710 325 711 331
rect 717 325 718 331
rect 710 215 718 325
rect 710 209 711 215
rect 717 209 718 215
rect 710 107 718 209
rect 710 101 711 107
rect 717 101 718 107
rect 710 72 718 101
rect 722 731 730 792
rect 722 725 723 731
rect 729 725 730 731
rect 722 611 730 725
rect 722 605 723 611
rect 729 605 730 611
rect 722 499 730 605
rect 722 493 723 499
rect 729 493 730 499
rect 722 387 730 493
rect 722 381 723 387
rect 729 381 730 387
rect 722 275 730 381
rect 722 269 723 275
rect 729 269 730 275
rect 722 159 730 269
rect 722 153 723 159
rect 729 153 730 159
rect 722 72 730 153
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0AND2X1  and_563_6
timestamp 1730743878
transform 1 0 144 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_563_6
timestamp 1730743878
transform 1 0 144 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_564_6
timestamp 1730743878
transform 1 0 184 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_564_6
timestamp 1730743878
transform 1 0 184 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_565_6
timestamp 1730743878
transform 1 0 224 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_565_6
timestamp 1730743878
transform 1 0 224 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_566_6
timestamp 1730743878
transform 1 0 264 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_566_6
timestamp 1730743878
transform 1 0 264 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_567_6
timestamp 1730743878
transform 1 0 304 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_567_6
timestamp 1730743878
transform 1 0 304 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_568_6
timestamp 1730743878
transform 1 0 344 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_568_6
timestamp 1730743878
transform 1 0 344 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_569_6
timestamp 1730743878
transform 1 0 384 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_569_6
timestamp 1730743878
transform 1 0 384 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_570_6
timestamp 1730743878
transform 1 0 424 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_570_6
timestamp 1730743878
transform 1 0 424 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_571_6
timestamp 1730743878
transform 1 0 464 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_571_6
timestamp 1730743878
transform 1 0 464 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_572_6
timestamp 1730743878
transform 1 0 512 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_572_6
timestamp 1730743878
transform 1 0 512 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_599_6
timestamp 1730743878
transform 1 0 552 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_599_6
timestamp 1730743878
transform 1 0 552 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_598_6
timestamp 1730743878
transform 1 0 592 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_598_6
timestamp 1730743878
transform 1 0 592 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_597_6
timestamp 1730743878
transform 1 0 632 0 1 104
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_597_6
timestamp 1730743878
transform 1 0 632 0 1 104
box 8 4 36 49
use welltap_svt  __well_tap__0
timestamp 1730743878
transform 1 0 104 0 1 120
box 8 4 12 24
use welltap_svt  __well_tap__0
timestamp 1730743878
transform 1 0 104 0 1 120
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_559_6
timestamp 1730743878
transform 1 0 144 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_559_6
timestamp 1730743878
transform 1 0 144 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_560_6
timestamp 1730743878
transform 1 0 192 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_560_6
timestamp 1730743878
transform 1 0 192 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_561_6
timestamp 1730743878
transform 1 0 248 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_561_6
timestamp 1730743878
transform 1 0 248 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_562_6
timestamp 1730743878
transform 1 0 304 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_562_6
timestamp 1730743878
transform 1 0 304 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_575_6
timestamp 1730743878
transform 1 0 360 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_575_6
timestamp 1730743878
transform 1 0 360 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_574_6
timestamp 1730743878
transform 1 0 416 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_574_6
timestamp 1730743878
transform 1 0 416 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_573_6
timestamp 1730743878
transform 1 0 472 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_573_6
timestamp 1730743878
transform 1 0 472 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_594_6
timestamp 1730743878
transform 1 0 528 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_594_6
timestamp 1730743878
transform 1 0 528 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_595_6
timestamp 1730743878
transform 1 0 592 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_595_6
timestamp 1730743878
transform 1 0 592 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_596_6
timestamp 1730743878
transform 1 0 632 0 -1 212
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_596_6
timestamp 1730743878
transform 1 0 632 0 -1 212
box 8 4 36 49
use welltap_svt  __well_tap__1
timestamp 1730743878
transform 1 0 680 0 1 120
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730743878
transform 1 0 680 0 1 120
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730743878
transform 1 0 104 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730743878
transform 1 0 104 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730743878
transform 1 0 680 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730743878
transform 1 0 680 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730743878
transform 1 0 104 0 1 236
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730743878
transform 1 0 104 0 1 236
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_558_6
timestamp 1730743878
transform 1 0 136 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_558_6
timestamp 1730743878
transform 1 0 136 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_557_6
timestamp 1730743878
transform 1 0 200 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_557_6
timestamp 1730743878
transform 1 0 200 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_555_6
timestamp 1730743878
transform 1 0 264 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_555_6
timestamp 1730743878
transform 1 0 264 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_556_6
timestamp 1730743878
transform 1 0 328 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_556_6
timestamp 1730743878
transform 1 0 328 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_576_6
timestamp 1730743878
transform 1 0 392 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_576_6
timestamp 1730743878
transform 1 0 392 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_577_6
timestamp 1730743878
transform 1 0 456 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_577_6
timestamp 1730743878
transform 1 0 456 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_593_6
timestamp 1730743878
transform 1 0 520 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_593_6
timestamp 1730743878
transform 1 0 520 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_592_6
timestamp 1730743878
transform 1 0 584 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_592_6
timestamp 1730743878
transform 1 0 584 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_591_6
timestamp 1730743878
transform 1 0 632 0 1 220
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_591_6
timestamp 1730743878
transform 1 0 632 0 1 220
box 8 4 36 49
use welltap_svt  __well_tap__5
timestamp 1730743878
transform 1 0 680 0 1 236
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730743878
transform 1 0 680 0 1 236
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730743878
transform 1 0 104 0 -1 312
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730743878
transform 1 0 104 0 -1 312
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_553_6
timestamp 1730743878
transform 1 0 200 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_553_6
timestamp 1730743878
transform 1 0 200 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_554_6
timestamp 1730743878
transform 1 0 240 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_554_6
timestamp 1730743878
transform 1 0 240 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_550_6
timestamp 1730743878
transform 1 0 288 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_550_6
timestamp 1730743878
transform 1 0 288 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_551_6
timestamp 1730743878
transform 1 0 344 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_551_6
timestamp 1730743878
transform 1 0 344 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_552_6
timestamp 1730743878
transform 1 0 400 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_552_6
timestamp 1730743878
transform 1 0 400 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_579_6
timestamp 1730743878
transform 1 0 456 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_579_6
timestamp 1730743878
transform 1 0 456 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_578_6
timestamp 1730743878
transform 1 0 520 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_578_6
timestamp 1730743878
transform 1 0 520 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_589_6
timestamp 1730743878
transform 1 0 584 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_589_6
timestamp 1730743878
transform 1 0 584 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_590_6
timestamp 1730743878
transform 1 0 632 0 -1 328
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_590_6
timestamp 1730743878
transform 1 0 632 0 -1 328
box 8 4 36 49
use welltap_svt  __well_tap__7
timestamp 1730743878
transform 1 0 680 0 -1 312
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730743878
transform 1 0 680 0 -1 312
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_548_6
timestamp 1730743878
transform 1 0 192 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_548_6
timestamp 1730743878
transform 1 0 192 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_549_6
timestamp 1730743878
transform 1 0 232 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_549_6
timestamp 1730743878
transform 1 0 232 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_547_6
timestamp 1730743878
transform 1 0 272 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_547_6
timestamp 1730743878
transform 1 0 272 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_546_6
timestamp 1730743878
transform 1 0 312 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_546_6
timestamp 1730743878
transform 1 0 312 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_545_6
timestamp 1730743878
transform 1 0 352 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_545_6
timestamp 1730743878
transform 1 0 352 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_544_6
timestamp 1730743878
transform 1 0 392 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_544_6
timestamp 1730743878
transform 1 0 392 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_580_6
timestamp 1730743878
transform 1 0 432 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_580_6
timestamp 1730743878
transform 1 0 432 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_581_6
timestamp 1730743878
transform 1 0 472 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_581_6
timestamp 1730743878
transform 1 0 472 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_582_6
timestamp 1730743878
transform 1 0 512 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_582_6
timestamp 1730743878
transform 1 0 512 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_588_6
timestamp 1730743878
transform 1 0 552 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_588_6
timestamp 1730743878
transform 1 0 552 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_587_6
timestamp 1730743878
transform 1 0 592 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_587_6
timestamp 1730743878
transform 1 0 592 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_586_6
timestamp 1730743878
transform 1 0 632 0 1 332
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_586_6
timestamp 1730743878
transform 1 0 632 0 1 332
box 8 4 36 49
use welltap_svt  __well_tap__8
timestamp 1730743878
transform 1 0 104 0 1 348
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730743878
transform 1 0 104 0 1 348
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_538_6
timestamp 1730743878
transform 1 0 256 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_538_6
timestamp 1730743878
transform 1 0 256 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_539_6
timestamp 1730743878
transform 1 0 296 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_539_6
timestamp 1730743878
transform 1 0 296 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_540_6
timestamp 1730743878
transform 1 0 336 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_540_6
timestamp 1730743878
transform 1 0 336 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_541_6
timestamp 1730743878
transform 1 0 384 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_541_6
timestamp 1730743878
transform 1 0 384 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_542_6
timestamp 1730743878
transform 1 0 432 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_542_6
timestamp 1730743878
transform 1 0 432 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_543_6
timestamp 1730743878
transform 1 0 480 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_543_6
timestamp 1730743878
transform 1 0 480 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_583_6
timestamp 1730743878
transform 1 0 528 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_583_6
timestamp 1730743878
transform 1 0 528 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_584_6
timestamp 1730743878
transform 1 0 584 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_584_6
timestamp 1730743878
transform 1 0 584 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_585_6
timestamp 1730743878
transform 1 0 632 0 -1 436
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_585_6
timestamp 1730743878
transform 1 0 632 0 -1 436
box 8 4 36 49
use welltap_svt  __well_tap__9
timestamp 1730743878
transform 1 0 680 0 1 348
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730743878
transform 1 0 680 0 1 348
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730743878
transform 1 0 104 0 -1 420
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730743878
transform 1 0 104 0 -1 420
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730743878
transform 1 0 680 0 -1 420
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730743878
transform 1 0 680 0 -1 420
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730743878
transform 1 0 104 0 1 460
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730743878
transform 1 0 104 0 1 460
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_531_6
timestamp 1730743878
transform 1 0 128 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_531_6
timestamp 1730743878
transform 1 0 128 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_532_6
timestamp 1730743878
transform 1 0 168 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_532_6
timestamp 1730743878
transform 1 0 168 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_533_6
timestamp 1730743878
transform 1 0 208 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_533_6
timestamp 1730743878
transform 1 0 208 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_534_6
timestamp 1730743878
transform 1 0 248 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_534_6
timestamp 1730743878
transform 1 0 248 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_535_6
timestamp 1730743878
transform 1 0 288 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_535_6
timestamp 1730743878
transform 1 0 288 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_536_6
timestamp 1730743878
transform 1 0 328 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_536_6
timestamp 1730743878
transform 1 0 328 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_537_6
timestamp 1730743878
transform 1 0 368 0 1 444
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_537_6
timestamp 1730743878
transform 1 0 368 0 1 444
box 8 4 36 49
use welltap_svt  __well_tap__13
timestamp 1730743878
transform 1 0 680 0 1 460
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730743878
transform 1 0 680 0 1 460
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730743878
transform 1 0 104 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730743878
transform 1 0 104 0 -1 536
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_525_6
timestamp 1730743878
transform 1 0 128 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_525_6
timestamp 1730743878
transform 1 0 128 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_526_6
timestamp 1730743878
transform 1 0 168 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_526_6
timestamp 1730743878
transform 1 0 168 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_527_6
timestamp 1730743878
transform 1 0 208 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_527_6
timestamp 1730743878
transform 1 0 208 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_528_6
timestamp 1730743878
transform 1 0 248 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_528_6
timestamp 1730743878
transform 1 0 248 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_529_6
timestamp 1730743878
transform 1 0 288 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_529_6
timestamp 1730743878
transform 1 0 288 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_530_6
timestamp 1730743878
transform 1 0 328 0 -1 552
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_530_6
timestamp 1730743878
transform 1 0 328 0 -1 552
box 8 4 36 49
use welltap_svt  __well_tap__15
timestamp 1730743878
transform 1 0 680 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730743878
transform 1 0 680 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730743878
transform 1 0 104 0 1 572
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730743878
transform 1 0 104 0 1 572
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_520_6
timestamp 1730743878
transform 1 0 128 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_520_6
timestamp 1730743878
transform 1 0 128 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_521_6
timestamp 1730743878
transform 1 0 168 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_521_6
timestamp 1730743878
transform 1 0 168 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_522_6
timestamp 1730743878
transform 1 0 208 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_522_6
timestamp 1730743878
transform 1 0 208 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_523_6
timestamp 1730743878
transform 1 0 248 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_523_6
timestamp 1730743878
transform 1 0 248 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_524_6
timestamp 1730743878
transform 1 0 288 0 1 556
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_524_6
timestamp 1730743878
transform 1 0 288 0 1 556
box 8 4 36 49
use welltap_svt  __well_tap__17
timestamp 1730743878
transform 1 0 680 0 1 572
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730743878
transform 1 0 680 0 1 572
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_514_6
timestamp 1730743878
transform 1 0 128 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_514_6
timestamp 1730743878
transform 1 0 128 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_515_6
timestamp 1730743878
transform 1 0 168 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_515_6
timestamp 1730743878
transform 1 0 168 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_516_6
timestamp 1730743878
transform 1 0 208 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_516_6
timestamp 1730743878
transform 1 0 208 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_517_6
timestamp 1730743878
transform 1 0 248 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_517_6
timestamp 1730743878
transform 1 0 248 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_518_6
timestamp 1730743878
transform 1 0 288 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_518_6
timestamp 1730743878
transform 1 0 288 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_519_6
timestamp 1730743878
transform 1 0 328 0 -1 668
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_519_6
timestamp 1730743878
transform 1 0 328 0 -1 668
box 8 4 36 49
use welltap_svt  __well_tap__18
timestamp 1730743878
transform 1 0 104 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730743878
transform 1 0 104 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730743878
transform 1 0 680 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730743878
transform 1 0 680 0 -1 652
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730743878
transform 1 0 104 0 1 692
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730743878
transform 1 0 104 0 1 692
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_58_6
timestamp 1730743878
transform 1 0 128 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_58_6
timestamp 1730743878
transform 1 0 128 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_59_6
timestamp 1730743878
transform 1 0 168 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_59_6
timestamp 1730743878
transform 1 0 168 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_510_6
timestamp 1730743878
transform 1 0 208 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_510_6
timestamp 1730743878
transform 1 0 208 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_511_6
timestamp 1730743878
transform 1 0 248 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_511_6
timestamp 1730743878
transform 1 0 248 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_512_6
timestamp 1730743878
transform 1 0 288 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_512_6
timestamp 1730743878
transform 1 0 288 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_513_6
timestamp 1730743878
transform 1 0 328 0 1 676
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_513_6
timestamp 1730743878
transform 1 0 328 0 1 676
box 8 4 36 49
use welltap_svt  __well_tap__21
timestamp 1730743878
transform 1 0 680 0 1 692
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730743878
transform 1 0 680 0 1 692
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730743878
transform 1 0 104 0 -1 764
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730743878
transform 1 0 104 0 -1 764
box 8 4 12 24
use _0_0std_0_0cells_0_0AND2X1  and_57_6
timestamp 1730743878
transform 1 0 128 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_57_6
timestamp 1730743878
transform 1 0 128 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_56_6
timestamp 1730743878
transform 1 0 168 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_56_6
timestamp 1730743878
transform 1 0 168 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_55_6
timestamp 1730743878
transform 1 0 208 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_55_6
timestamp 1730743878
transform 1 0 208 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_54_6
timestamp 1730743878
transform 1 0 248 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_54_6
timestamp 1730743878
transform 1 0 248 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_53_6
timestamp 1730743878
transform 1 0 288 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_53_6
timestamp 1730743878
transform 1 0 288 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_52_6
timestamp 1730743878
transform 1 0 328 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_52_6
timestamp 1730743878
transform 1 0 328 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_51_6
timestamp 1730743878
transform 1 0 368 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_51_6
timestamp 1730743878
transform 1 0 368 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_50_6
timestamp 1730743878
transform 1 0 408 0 -1 780
box 8 4 36 49
use _0_0std_0_0cells_0_0AND2X1  and_50_6
timestamp 1730743878
transform 1 0 408 0 -1 780
box 8 4 36 49
use welltap_svt  __well_tap__23
timestamp 1730743878
transform 1 0 680 0 -1 764
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730743878
transform 1 0 680 0 -1 764
box 8 4 12 24
<< end >>
