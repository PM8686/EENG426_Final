magic
tech sky130l
timestamp 1731220618
<< m2 >>
rect 1686 2212 1692 2213
rect 134 2208 140 2209
rect 110 2205 116 2206
rect 110 2201 111 2205
rect 115 2201 116 2205
rect 134 2204 135 2208
rect 139 2204 140 2208
rect 134 2203 140 2204
rect 174 2208 180 2209
rect 174 2204 175 2208
rect 179 2204 180 2208
rect 174 2203 180 2204
rect 214 2208 220 2209
rect 214 2204 215 2208
rect 219 2204 220 2208
rect 214 2203 220 2204
rect 254 2208 260 2209
rect 254 2204 255 2208
rect 259 2204 260 2208
rect 254 2203 260 2204
rect 318 2208 324 2209
rect 318 2204 319 2208
rect 323 2204 324 2208
rect 318 2203 324 2204
rect 382 2208 388 2209
rect 382 2204 383 2208
rect 387 2204 388 2208
rect 382 2203 388 2204
rect 446 2208 452 2209
rect 446 2204 447 2208
rect 451 2204 452 2208
rect 446 2203 452 2204
rect 510 2208 516 2209
rect 510 2204 511 2208
rect 515 2204 516 2208
rect 510 2203 516 2204
rect 574 2208 580 2209
rect 574 2204 575 2208
rect 579 2204 580 2208
rect 574 2203 580 2204
rect 630 2208 636 2209
rect 630 2204 631 2208
rect 635 2204 636 2208
rect 630 2203 636 2204
rect 686 2208 692 2209
rect 686 2204 687 2208
rect 691 2204 692 2208
rect 686 2203 692 2204
rect 734 2208 740 2209
rect 734 2204 735 2208
rect 739 2204 740 2208
rect 734 2203 740 2204
rect 790 2208 796 2209
rect 790 2204 791 2208
rect 795 2204 796 2208
rect 790 2203 796 2204
rect 846 2208 852 2209
rect 846 2204 847 2208
rect 851 2204 852 2208
rect 846 2203 852 2204
rect 902 2208 908 2209
rect 902 2204 903 2208
rect 907 2204 908 2208
rect 1686 2208 1687 2212
rect 1691 2208 1692 2212
rect 1686 2207 1692 2208
rect 1726 2212 1732 2213
rect 1726 2208 1727 2212
rect 1731 2208 1732 2212
rect 1726 2207 1732 2208
rect 1766 2212 1772 2213
rect 1766 2208 1767 2212
rect 1771 2208 1772 2212
rect 1766 2207 1772 2208
rect 1806 2212 1812 2213
rect 1806 2208 1807 2212
rect 1811 2208 1812 2212
rect 1806 2207 1812 2208
rect 902 2203 908 2204
rect 1094 2205 1100 2206
rect 110 2200 116 2201
rect 1094 2201 1095 2205
rect 1099 2201 1100 2205
rect 1094 2200 1100 2201
rect 1134 2204 1140 2205
rect 1134 2200 1135 2204
rect 1139 2200 1140 2204
rect 1134 2199 1140 2200
rect 2118 2204 2124 2205
rect 2118 2200 2119 2204
rect 2123 2200 2124 2204
rect 2118 2199 2124 2200
rect 110 2188 116 2189
rect 110 2184 111 2188
rect 115 2184 116 2188
rect 110 2183 116 2184
rect 1094 2188 1100 2189
rect 1094 2184 1095 2188
rect 1099 2184 1100 2188
rect 1094 2183 1100 2184
rect 1134 2187 1140 2188
rect 1134 2183 1135 2187
rect 1139 2183 1140 2187
rect 2118 2187 2124 2188
rect 1134 2182 1140 2183
rect 1686 2184 1692 2185
rect 134 2180 140 2181
rect 134 2176 135 2180
rect 139 2176 140 2180
rect 134 2175 140 2176
rect 174 2180 180 2181
rect 174 2176 175 2180
rect 179 2176 180 2180
rect 174 2175 180 2176
rect 214 2180 220 2181
rect 214 2176 215 2180
rect 219 2176 220 2180
rect 214 2175 220 2176
rect 254 2180 260 2181
rect 254 2176 255 2180
rect 259 2176 260 2180
rect 254 2175 260 2176
rect 318 2180 324 2181
rect 318 2176 319 2180
rect 323 2176 324 2180
rect 318 2175 324 2176
rect 382 2180 388 2181
rect 382 2176 383 2180
rect 387 2176 388 2180
rect 382 2175 388 2176
rect 446 2180 452 2181
rect 446 2176 447 2180
rect 451 2176 452 2180
rect 446 2175 452 2176
rect 510 2180 516 2181
rect 510 2176 511 2180
rect 515 2176 516 2180
rect 510 2175 516 2176
rect 574 2180 580 2181
rect 574 2176 575 2180
rect 579 2176 580 2180
rect 574 2175 580 2176
rect 630 2180 636 2181
rect 630 2176 631 2180
rect 635 2176 636 2180
rect 630 2175 636 2176
rect 686 2180 692 2181
rect 686 2176 687 2180
rect 691 2176 692 2180
rect 686 2175 692 2176
rect 734 2180 740 2181
rect 734 2176 735 2180
rect 739 2176 740 2180
rect 734 2175 740 2176
rect 790 2180 796 2181
rect 790 2176 791 2180
rect 795 2176 796 2180
rect 790 2175 796 2176
rect 846 2180 852 2181
rect 846 2176 847 2180
rect 851 2176 852 2180
rect 846 2175 852 2176
rect 902 2180 908 2181
rect 902 2176 903 2180
rect 907 2176 908 2180
rect 1686 2180 1687 2184
rect 1691 2180 1692 2184
rect 1686 2179 1692 2180
rect 1726 2184 1732 2185
rect 1726 2180 1727 2184
rect 1731 2180 1732 2184
rect 1726 2179 1732 2180
rect 1766 2184 1772 2185
rect 1766 2180 1767 2184
rect 1771 2180 1772 2184
rect 1766 2179 1772 2180
rect 1806 2184 1812 2185
rect 1806 2180 1807 2184
rect 1811 2180 1812 2184
rect 2118 2183 2119 2187
rect 2123 2183 2124 2187
rect 2118 2182 2124 2183
rect 1806 2179 1812 2180
rect 902 2175 908 2176
rect 1158 2172 1164 2173
rect 1134 2169 1140 2170
rect 1134 2165 1135 2169
rect 1139 2165 1140 2169
rect 1158 2168 1159 2172
rect 1163 2168 1164 2172
rect 1158 2167 1164 2168
rect 1198 2172 1204 2173
rect 1198 2168 1199 2172
rect 1203 2168 1204 2172
rect 1198 2167 1204 2168
rect 1238 2172 1244 2173
rect 1238 2168 1239 2172
rect 1243 2168 1244 2172
rect 1238 2167 1244 2168
rect 1278 2172 1284 2173
rect 1278 2168 1279 2172
rect 1283 2168 1284 2172
rect 1278 2167 1284 2168
rect 1334 2172 1340 2173
rect 1334 2168 1335 2172
rect 1339 2168 1340 2172
rect 1334 2167 1340 2168
rect 1390 2172 1396 2173
rect 1390 2168 1391 2172
rect 1395 2168 1396 2172
rect 1390 2167 1396 2168
rect 1454 2172 1460 2173
rect 1454 2168 1455 2172
rect 1459 2168 1460 2172
rect 1454 2167 1460 2168
rect 1526 2172 1532 2173
rect 1526 2168 1527 2172
rect 1531 2168 1532 2172
rect 1526 2167 1532 2168
rect 1590 2172 1596 2173
rect 1590 2168 1591 2172
rect 1595 2168 1596 2172
rect 1590 2167 1596 2168
rect 1662 2172 1668 2173
rect 1662 2168 1663 2172
rect 1667 2168 1668 2172
rect 1662 2167 1668 2168
rect 1734 2172 1740 2173
rect 1734 2168 1735 2172
rect 1739 2168 1740 2172
rect 1734 2167 1740 2168
rect 1806 2172 1812 2173
rect 1806 2168 1807 2172
rect 1811 2168 1812 2172
rect 1806 2167 1812 2168
rect 1878 2172 1884 2173
rect 1878 2168 1879 2172
rect 1883 2168 1884 2172
rect 1878 2167 1884 2168
rect 2118 2169 2124 2170
rect 1134 2164 1140 2165
rect 2118 2165 2119 2169
rect 2123 2165 2124 2169
rect 2118 2164 2124 2165
rect 1134 2152 1140 2153
rect 1134 2148 1135 2152
rect 1139 2148 1140 2152
rect 1134 2147 1140 2148
rect 2118 2152 2124 2153
rect 2118 2148 2119 2152
rect 2123 2148 2124 2152
rect 2118 2147 2124 2148
rect 1158 2144 1164 2145
rect 1158 2140 1159 2144
rect 1163 2140 1164 2144
rect 1158 2139 1164 2140
rect 1198 2144 1204 2145
rect 1198 2140 1199 2144
rect 1203 2140 1204 2144
rect 1198 2139 1204 2140
rect 1238 2144 1244 2145
rect 1238 2140 1239 2144
rect 1243 2140 1244 2144
rect 1238 2139 1244 2140
rect 1278 2144 1284 2145
rect 1278 2140 1279 2144
rect 1283 2140 1284 2144
rect 1278 2139 1284 2140
rect 1334 2144 1340 2145
rect 1334 2140 1335 2144
rect 1339 2140 1340 2144
rect 1334 2139 1340 2140
rect 1390 2144 1396 2145
rect 1390 2140 1391 2144
rect 1395 2140 1396 2144
rect 1390 2139 1396 2140
rect 1454 2144 1460 2145
rect 1454 2140 1455 2144
rect 1459 2140 1460 2144
rect 1454 2139 1460 2140
rect 1526 2144 1532 2145
rect 1526 2140 1527 2144
rect 1531 2140 1532 2144
rect 1526 2139 1532 2140
rect 1590 2144 1596 2145
rect 1590 2140 1591 2144
rect 1595 2140 1596 2144
rect 1590 2139 1596 2140
rect 1662 2144 1668 2145
rect 1662 2140 1663 2144
rect 1667 2140 1668 2144
rect 1662 2139 1668 2140
rect 1734 2144 1740 2145
rect 1734 2140 1735 2144
rect 1739 2140 1740 2144
rect 1734 2139 1740 2140
rect 1806 2144 1812 2145
rect 1806 2140 1807 2144
rect 1811 2140 1812 2144
rect 1806 2139 1812 2140
rect 1878 2144 1884 2145
rect 1878 2140 1879 2144
rect 1883 2140 1884 2144
rect 1878 2139 1884 2140
rect 230 2136 236 2137
rect 230 2132 231 2136
rect 235 2132 236 2136
rect 230 2131 236 2132
rect 270 2136 276 2137
rect 270 2132 271 2136
rect 275 2132 276 2136
rect 270 2131 276 2132
rect 310 2136 316 2137
rect 310 2132 311 2136
rect 315 2132 316 2136
rect 310 2131 316 2132
rect 358 2136 364 2137
rect 358 2132 359 2136
rect 363 2132 364 2136
rect 358 2131 364 2132
rect 422 2136 428 2137
rect 422 2132 423 2136
rect 427 2132 428 2136
rect 422 2131 428 2132
rect 486 2136 492 2137
rect 486 2132 487 2136
rect 491 2132 492 2136
rect 486 2131 492 2132
rect 558 2136 564 2137
rect 558 2132 559 2136
rect 563 2132 564 2136
rect 558 2131 564 2132
rect 638 2136 644 2137
rect 638 2132 639 2136
rect 643 2132 644 2136
rect 638 2131 644 2132
rect 718 2136 724 2137
rect 718 2132 719 2136
rect 723 2132 724 2136
rect 718 2131 724 2132
rect 798 2136 804 2137
rect 798 2132 799 2136
rect 803 2132 804 2136
rect 798 2131 804 2132
rect 878 2136 884 2137
rect 878 2132 879 2136
rect 883 2132 884 2136
rect 878 2131 884 2132
rect 966 2136 972 2137
rect 966 2132 967 2136
rect 971 2132 972 2136
rect 966 2131 972 2132
rect 110 2128 116 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 1094 2128 1100 2129
rect 1094 2124 1095 2128
rect 1099 2124 1100 2128
rect 1094 2123 1100 2124
rect 110 2111 116 2112
rect 110 2107 111 2111
rect 115 2107 116 2111
rect 1094 2111 1100 2112
rect 110 2106 116 2107
rect 230 2108 236 2109
rect 230 2104 231 2108
rect 235 2104 236 2108
rect 230 2103 236 2104
rect 270 2108 276 2109
rect 270 2104 271 2108
rect 275 2104 276 2108
rect 270 2103 276 2104
rect 310 2108 316 2109
rect 310 2104 311 2108
rect 315 2104 316 2108
rect 310 2103 316 2104
rect 358 2108 364 2109
rect 358 2104 359 2108
rect 363 2104 364 2108
rect 358 2103 364 2104
rect 422 2108 428 2109
rect 422 2104 423 2108
rect 427 2104 428 2108
rect 422 2103 428 2104
rect 486 2108 492 2109
rect 486 2104 487 2108
rect 491 2104 492 2108
rect 486 2103 492 2104
rect 558 2108 564 2109
rect 558 2104 559 2108
rect 563 2104 564 2108
rect 558 2103 564 2104
rect 638 2108 644 2109
rect 638 2104 639 2108
rect 643 2104 644 2108
rect 638 2103 644 2104
rect 718 2108 724 2109
rect 718 2104 719 2108
rect 723 2104 724 2108
rect 718 2103 724 2104
rect 798 2108 804 2109
rect 798 2104 799 2108
rect 803 2104 804 2108
rect 798 2103 804 2104
rect 878 2108 884 2109
rect 878 2104 879 2108
rect 883 2104 884 2108
rect 878 2103 884 2104
rect 966 2108 972 2109
rect 966 2104 967 2108
rect 971 2104 972 2108
rect 1094 2107 1095 2111
rect 1099 2107 1100 2111
rect 1094 2106 1100 2107
rect 1158 2108 1164 2109
rect 966 2103 972 2104
rect 1158 2104 1159 2108
rect 1163 2104 1164 2108
rect 1158 2103 1164 2104
rect 1198 2108 1204 2109
rect 1198 2104 1199 2108
rect 1203 2104 1204 2108
rect 1198 2103 1204 2104
rect 1238 2108 1244 2109
rect 1238 2104 1239 2108
rect 1243 2104 1244 2108
rect 1238 2103 1244 2104
rect 1294 2108 1300 2109
rect 1294 2104 1295 2108
rect 1299 2104 1300 2108
rect 1294 2103 1300 2104
rect 1366 2108 1372 2109
rect 1366 2104 1367 2108
rect 1371 2104 1372 2108
rect 1366 2103 1372 2104
rect 1438 2108 1444 2109
rect 1438 2104 1439 2108
rect 1443 2104 1444 2108
rect 1438 2103 1444 2104
rect 1518 2108 1524 2109
rect 1518 2104 1519 2108
rect 1523 2104 1524 2108
rect 1518 2103 1524 2104
rect 1598 2108 1604 2109
rect 1598 2104 1599 2108
rect 1603 2104 1604 2108
rect 1598 2103 1604 2104
rect 1678 2108 1684 2109
rect 1678 2104 1679 2108
rect 1683 2104 1684 2108
rect 1678 2103 1684 2104
rect 1750 2108 1756 2109
rect 1750 2104 1751 2108
rect 1755 2104 1756 2108
rect 1750 2103 1756 2104
rect 1822 2108 1828 2109
rect 1822 2104 1823 2108
rect 1827 2104 1828 2108
rect 1822 2103 1828 2104
rect 1886 2108 1892 2109
rect 1886 2104 1887 2108
rect 1891 2104 1892 2108
rect 1886 2103 1892 2104
rect 1950 2108 1956 2109
rect 1950 2104 1951 2108
rect 1955 2104 1956 2108
rect 1950 2103 1956 2104
rect 2022 2108 2028 2109
rect 2022 2104 2023 2108
rect 2027 2104 2028 2108
rect 2022 2103 2028 2104
rect 2070 2108 2076 2109
rect 2070 2104 2071 2108
rect 2075 2104 2076 2108
rect 2070 2103 2076 2104
rect 1134 2100 1140 2101
rect 1134 2096 1135 2100
rect 1139 2096 1140 2100
rect 1134 2095 1140 2096
rect 2118 2100 2124 2101
rect 2118 2096 2119 2100
rect 2123 2096 2124 2100
rect 2118 2095 2124 2096
rect 302 2092 308 2093
rect 110 2089 116 2090
rect 110 2085 111 2089
rect 115 2085 116 2089
rect 302 2088 303 2092
rect 307 2088 308 2092
rect 302 2087 308 2088
rect 350 2092 356 2093
rect 350 2088 351 2092
rect 355 2088 356 2092
rect 350 2087 356 2088
rect 406 2092 412 2093
rect 406 2088 407 2092
rect 411 2088 412 2092
rect 406 2087 412 2088
rect 470 2092 476 2093
rect 470 2088 471 2092
rect 475 2088 476 2092
rect 470 2087 476 2088
rect 542 2092 548 2093
rect 542 2088 543 2092
rect 547 2088 548 2092
rect 542 2087 548 2088
rect 622 2092 628 2093
rect 622 2088 623 2092
rect 627 2088 628 2092
rect 622 2087 628 2088
rect 702 2092 708 2093
rect 702 2088 703 2092
rect 707 2088 708 2092
rect 702 2087 708 2088
rect 782 2092 788 2093
rect 782 2088 783 2092
rect 787 2088 788 2092
rect 782 2087 788 2088
rect 862 2092 868 2093
rect 862 2088 863 2092
rect 867 2088 868 2092
rect 862 2087 868 2088
rect 950 2092 956 2093
rect 950 2088 951 2092
rect 955 2088 956 2092
rect 950 2087 956 2088
rect 1038 2092 1044 2093
rect 1038 2088 1039 2092
rect 1043 2088 1044 2092
rect 1038 2087 1044 2088
rect 1094 2089 1100 2090
rect 110 2084 116 2085
rect 1094 2085 1095 2089
rect 1099 2085 1100 2089
rect 1094 2084 1100 2085
rect 1134 2083 1140 2084
rect 1134 2079 1135 2083
rect 1139 2079 1140 2083
rect 2118 2083 2124 2084
rect 1134 2078 1140 2079
rect 1158 2080 1164 2081
rect 1158 2076 1159 2080
rect 1163 2076 1164 2080
rect 1158 2075 1164 2076
rect 1198 2080 1204 2081
rect 1198 2076 1199 2080
rect 1203 2076 1204 2080
rect 1198 2075 1204 2076
rect 1238 2080 1244 2081
rect 1238 2076 1239 2080
rect 1243 2076 1244 2080
rect 1238 2075 1244 2076
rect 1294 2080 1300 2081
rect 1294 2076 1295 2080
rect 1299 2076 1300 2080
rect 1294 2075 1300 2076
rect 1366 2080 1372 2081
rect 1366 2076 1367 2080
rect 1371 2076 1372 2080
rect 1366 2075 1372 2076
rect 1438 2080 1444 2081
rect 1438 2076 1439 2080
rect 1443 2076 1444 2080
rect 1438 2075 1444 2076
rect 1518 2080 1524 2081
rect 1518 2076 1519 2080
rect 1523 2076 1524 2080
rect 1518 2075 1524 2076
rect 1598 2080 1604 2081
rect 1598 2076 1599 2080
rect 1603 2076 1604 2080
rect 1598 2075 1604 2076
rect 1678 2080 1684 2081
rect 1678 2076 1679 2080
rect 1683 2076 1684 2080
rect 1678 2075 1684 2076
rect 1750 2080 1756 2081
rect 1750 2076 1751 2080
rect 1755 2076 1756 2080
rect 1750 2075 1756 2076
rect 1822 2080 1828 2081
rect 1822 2076 1823 2080
rect 1827 2076 1828 2080
rect 1822 2075 1828 2076
rect 1886 2080 1892 2081
rect 1886 2076 1887 2080
rect 1891 2076 1892 2080
rect 1886 2075 1892 2076
rect 1950 2080 1956 2081
rect 1950 2076 1951 2080
rect 1955 2076 1956 2080
rect 1950 2075 1956 2076
rect 2022 2080 2028 2081
rect 2022 2076 2023 2080
rect 2027 2076 2028 2080
rect 2022 2075 2028 2076
rect 2070 2080 2076 2081
rect 2070 2076 2071 2080
rect 2075 2076 2076 2080
rect 2118 2079 2119 2083
rect 2123 2079 2124 2083
rect 2118 2078 2124 2079
rect 2070 2075 2076 2076
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 1094 2072 1100 2073
rect 1094 2068 1095 2072
rect 1099 2068 1100 2072
rect 1094 2067 1100 2068
rect 1158 2068 1164 2069
rect 1134 2065 1140 2066
rect 302 2064 308 2065
rect 302 2060 303 2064
rect 307 2060 308 2064
rect 302 2059 308 2060
rect 350 2064 356 2065
rect 350 2060 351 2064
rect 355 2060 356 2064
rect 350 2059 356 2060
rect 406 2064 412 2065
rect 406 2060 407 2064
rect 411 2060 412 2064
rect 406 2059 412 2060
rect 470 2064 476 2065
rect 470 2060 471 2064
rect 475 2060 476 2064
rect 470 2059 476 2060
rect 542 2064 548 2065
rect 542 2060 543 2064
rect 547 2060 548 2064
rect 542 2059 548 2060
rect 622 2064 628 2065
rect 622 2060 623 2064
rect 627 2060 628 2064
rect 622 2059 628 2060
rect 702 2064 708 2065
rect 702 2060 703 2064
rect 707 2060 708 2064
rect 702 2059 708 2060
rect 782 2064 788 2065
rect 782 2060 783 2064
rect 787 2060 788 2064
rect 782 2059 788 2060
rect 862 2064 868 2065
rect 862 2060 863 2064
rect 867 2060 868 2064
rect 862 2059 868 2060
rect 950 2064 956 2065
rect 950 2060 951 2064
rect 955 2060 956 2064
rect 950 2059 956 2060
rect 1038 2064 1044 2065
rect 1038 2060 1039 2064
rect 1043 2060 1044 2064
rect 1134 2061 1135 2065
rect 1139 2061 1140 2065
rect 1158 2064 1159 2068
rect 1163 2064 1164 2068
rect 1158 2063 1164 2064
rect 1214 2068 1220 2069
rect 1214 2064 1215 2068
rect 1219 2064 1220 2068
rect 1214 2063 1220 2064
rect 1302 2068 1308 2069
rect 1302 2064 1303 2068
rect 1307 2064 1308 2068
rect 1302 2063 1308 2064
rect 1398 2068 1404 2069
rect 1398 2064 1399 2068
rect 1403 2064 1404 2068
rect 1398 2063 1404 2064
rect 1494 2068 1500 2069
rect 1494 2064 1495 2068
rect 1499 2064 1500 2068
rect 1494 2063 1500 2064
rect 1590 2068 1596 2069
rect 1590 2064 1591 2068
rect 1595 2064 1596 2068
rect 1590 2063 1596 2064
rect 1678 2068 1684 2069
rect 1678 2064 1679 2068
rect 1683 2064 1684 2068
rect 1678 2063 1684 2064
rect 1758 2068 1764 2069
rect 1758 2064 1759 2068
rect 1763 2064 1764 2068
rect 1758 2063 1764 2064
rect 1830 2068 1836 2069
rect 1830 2064 1831 2068
rect 1835 2064 1836 2068
rect 1830 2063 1836 2064
rect 1894 2068 1900 2069
rect 1894 2064 1895 2068
rect 1899 2064 1900 2068
rect 1894 2063 1900 2064
rect 1958 2068 1964 2069
rect 1958 2064 1959 2068
rect 1963 2064 1964 2068
rect 1958 2063 1964 2064
rect 2022 2068 2028 2069
rect 2022 2064 2023 2068
rect 2027 2064 2028 2068
rect 2022 2063 2028 2064
rect 2070 2068 2076 2069
rect 2070 2064 2071 2068
rect 2075 2064 2076 2068
rect 2070 2063 2076 2064
rect 2118 2065 2124 2066
rect 1134 2060 1140 2061
rect 2118 2061 2119 2065
rect 2123 2061 2124 2065
rect 2118 2060 2124 2061
rect 1038 2059 1044 2060
rect 1134 2048 1140 2049
rect 1134 2044 1135 2048
rect 1139 2044 1140 2048
rect 1134 2043 1140 2044
rect 2118 2048 2124 2049
rect 2118 2044 2119 2048
rect 2123 2044 2124 2048
rect 2118 2043 2124 2044
rect 1158 2040 1164 2041
rect 1158 2036 1159 2040
rect 1163 2036 1164 2040
rect 1158 2035 1164 2036
rect 1214 2040 1220 2041
rect 1214 2036 1215 2040
rect 1219 2036 1220 2040
rect 1214 2035 1220 2036
rect 1302 2040 1308 2041
rect 1302 2036 1303 2040
rect 1307 2036 1308 2040
rect 1302 2035 1308 2036
rect 1398 2040 1404 2041
rect 1398 2036 1399 2040
rect 1403 2036 1404 2040
rect 1398 2035 1404 2036
rect 1494 2040 1500 2041
rect 1494 2036 1495 2040
rect 1499 2036 1500 2040
rect 1494 2035 1500 2036
rect 1590 2040 1596 2041
rect 1590 2036 1591 2040
rect 1595 2036 1596 2040
rect 1590 2035 1596 2036
rect 1678 2040 1684 2041
rect 1678 2036 1679 2040
rect 1683 2036 1684 2040
rect 1678 2035 1684 2036
rect 1758 2040 1764 2041
rect 1758 2036 1759 2040
rect 1763 2036 1764 2040
rect 1758 2035 1764 2036
rect 1830 2040 1836 2041
rect 1830 2036 1831 2040
rect 1835 2036 1836 2040
rect 1830 2035 1836 2036
rect 1894 2040 1900 2041
rect 1894 2036 1895 2040
rect 1899 2036 1900 2040
rect 1894 2035 1900 2036
rect 1958 2040 1964 2041
rect 1958 2036 1959 2040
rect 1963 2036 1964 2040
rect 1958 2035 1964 2036
rect 2022 2040 2028 2041
rect 2022 2036 2023 2040
rect 2027 2036 2028 2040
rect 2022 2035 2028 2036
rect 2070 2040 2076 2041
rect 2070 2036 2071 2040
rect 2075 2036 2076 2040
rect 2070 2035 2076 2036
rect 182 2024 188 2025
rect 182 2020 183 2024
rect 187 2020 188 2024
rect 182 2019 188 2020
rect 278 2024 284 2025
rect 278 2020 279 2024
rect 283 2020 284 2024
rect 278 2019 284 2020
rect 374 2024 380 2025
rect 374 2020 375 2024
rect 379 2020 380 2024
rect 374 2019 380 2020
rect 462 2024 468 2025
rect 462 2020 463 2024
rect 467 2020 468 2024
rect 462 2019 468 2020
rect 542 2024 548 2025
rect 542 2020 543 2024
rect 547 2020 548 2024
rect 542 2019 548 2020
rect 622 2024 628 2025
rect 622 2020 623 2024
rect 627 2020 628 2024
rect 622 2019 628 2020
rect 694 2024 700 2025
rect 694 2020 695 2024
rect 699 2020 700 2024
rect 694 2019 700 2020
rect 758 2024 764 2025
rect 758 2020 759 2024
rect 763 2020 764 2024
rect 758 2019 764 2020
rect 814 2024 820 2025
rect 814 2020 815 2024
rect 819 2020 820 2024
rect 814 2019 820 2020
rect 862 2024 868 2025
rect 862 2020 863 2024
rect 867 2020 868 2024
rect 862 2019 868 2020
rect 910 2024 916 2025
rect 910 2020 911 2024
rect 915 2020 916 2024
rect 910 2019 916 2020
rect 958 2024 964 2025
rect 958 2020 959 2024
rect 963 2020 964 2024
rect 958 2019 964 2020
rect 1006 2024 1012 2025
rect 1006 2020 1007 2024
rect 1011 2020 1012 2024
rect 1006 2019 1012 2020
rect 1046 2024 1052 2025
rect 1046 2020 1047 2024
rect 1051 2020 1052 2024
rect 1046 2019 1052 2020
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 110 2011 116 2012
rect 1094 2016 1100 2017
rect 1094 2012 1095 2016
rect 1099 2012 1100 2016
rect 1094 2011 1100 2012
rect 1158 2004 1164 2005
rect 1158 2000 1159 2004
rect 1163 2000 1164 2004
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 1094 1999 1100 2000
rect 1158 1999 1164 2000
rect 1238 2004 1244 2005
rect 1238 2000 1239 2004
rect 1243 2000 1244 2004
rect 1238 1999 1244 2000
rect 1350 2004 1356 2005
rect 1350 2000 1351 2004
rect 1355 2000 1356 2004
rect 1350 1999 1356 2000
rect 1454 2004 1460 2005
rect 1454 2000 1455 2004
rect 1459 2000 1460 2004
rect 1454 1999 1460 2000
rect 1558 2004 1564 2005
rect 1558 2000 1559 2004
rect 1563 2000 1564 2004
rect 1558 1999 1564 2000
rect 1654 2004 1660 2005
rect 1654 2000 1655 2004
rect 1659 2000 1660 2004
rect 1654 1999 1660 2000
rect 1742 2004 1748 2005
rect 1742 2000 1743 2004
rect 1747 2000 1748 2004
rect 1742 1999 1748 2000
rect 1822 2004 1828 2005
rect 1822 2000 1823 2004
rect 1827 2000 1828 2004
rect 1822 1999 1828 2000
rect 1894 2004 1900 2005
rect 1894 2000 1895 2004
rect 1899 2000 1900 2004
rect 1894 1999 1900 2000
rect 1958 2004 1964 2005
rect 1958 2000 1959 2004
rect 1963 2000 1964 2004
rect 1958 1999 1964 2000
rect 2022 2004 2028 2005
rect 2022 2000 2023 2004
rect 2027 2000 2028 2004
rect 2022 1999 2028 2000
rect 2070 2004 2076 2005
rect 2070 2000 2071 2004
rect 2075 2000 2076 2004
rect 2070 1999 2076 2000
rect 110 1994 116 1995
rect 182 1996 188 1997
rect 182 1992 183 1996
rect 187 1992 188 1996
rect 182 1991 188 1992
rect 278 1996 284 1997
rect 278 1992 279 1996
rect 283 1992 284 1996
rect 278 1991 284 1992
rect 374 1996 380 1997
rect 374 1992 375 1996
rect 379 1992 380 1996
rect 374 1991 380 1992
rect 462 1996 468 1997
rect 462 1992 463 1996
rect 467 1992 468 1996
rect 462 1991 468 1992
rect 542 1996 548 1997
rect 542 1992 543 1996
rect 547 1992 548 1996
rect 542 1991 548 1992
rect 622 1996 628 1997
rect 622 1992 623 1996
rect 627 1992 628 1996
rect 622 1991 628 1992
rect 694 1996 700 1997
rect 694 1992 695 1996
rect 699 1992 700 1996
rect 694 1991 700 1992
rect 758 1996 764 1997
rect 758 1992 759 1996
rect 763 1992 764 1996
rect 758 1991 764 1992
rect 814 1996 820 1997
rect 814 1992 815 1996
rect 819 1992 820 1996
rect 814 1991 820 1992
rect 862 1996 868 1997
rect 862 1992 863 1996
rect 867 1992 868 1996
rect 862 1991 868 1992
rect 910 1996 916 1997
rect 910 1992 911 1996
rect 915 1992 916 1996
rect 910 1991 916 1992
rect 958 1996 964 1997
rect 958 1992 959 1996
rect 963 1992 964 1996
rect 958 1991 964 1992
rect 1006 1996 1012 1997
rect 1006 1992 1007 1996
rect 1011 1992 1012 1996
rect 1006 1991 1012 1992
rect 1046 1996 1052 1997
rect 1046 1992 1047 1996
rect 1051 1992 1052 1996
rect 1094 1995 1095 1999
rect 1099 1995 1100 1999
rect 1094 1994 1100 1995
rect 1134 1996 1140 1997
rect 1046 1991 1052 1992
rect 1134 1992 1135 1996
rect 1139 1992 1140 1996
rect 1134 1991 1140 1992
rect 2118 1996 2124 1997
rect 2118 1992 2119 1996
rect 2123 1992 2124 1996
rect 2118 1991 2124 1992
rect 158 1984 164 1985
rect 110 1981 116 1982
rect 110 1977 111 1981
rect 115 1977 116 1981
rect 158 1980 159 1984
rect 163 1980 164 1984
rect 158 1979 164 1980
rect 230 1984 236 1985
rect 230 1980 231 1984
rect 235 1980 236 1984
rect 230 1979 236 1980
rect 302 1984 308 1985
rect 302 1980 303 1984
rect 307 1980 308 1984
rect 302 1979 308 1980
rect 374 1984 380 1985
rect 374 1980 375 1984
rect 379 1980 380 1984
rect 374 1979 380 1980
rect 446 1984 452 1985
rect 446 1980 447 1984
rect 451 1980 452 1984
rect 446 1979 452 1980
rect 526 1984 532 1985
rect 526 1980 527 1984
rect 531 1980 532 1984
rect 526 1979 532 1980
rect 606 1984 612 1985
rect 606 1980 607 1984
rect 611 1980 612 1984
rect 606 1979 612 1980
rect 686 1984 692 1985
rect 686 1980 687 1984
rect 691 1980 692 1984
rect 686 1979 692 1980
rect 758 1984 764 1985
rect 758 1980 759 1984
rect 763 1980 764 1984
rect 758 1979 764 1980
rect 830 1984 836 1985
rect 830 1980 831 1984
rect 835 1980 836 1984
rect 830 1979 836 1980
rect 910 1984 916 1985
rect 910 1980 911 1984
rect 915 1980 916 1984
rect 910 1979 916 1980
rect 990 1984 996 1985
rect 990 1980 991 1984
rect 995 1980 996 1984
rect 990 1979 996 1980
rect 1094 1981 1100 1982
rect 110 1976 116 1977
rect 1094 1977 1095 1981
rect 1099 1977 1100 1981
rect 1094 1976 1100 1977
rect 1134 1979 1140 1980
rect 1134 1975 1135 1979
rect 1139 1975 1140 1979
rect 2118 1979 2124 1980
rect 1134 1974 1140 1975
rect 1158 1976 1164 1977
rect 1158 1972 1159 1976
rect 1163 1972 1164 1976
rect 1158 1971 1164 1972
rect 1238 1976 1244 1977
rect 1238 1972 1239 1976
rect 1243 1972 1244 1976
rect 1238 1971 1244 1972
rect 1350 1976 1356 1977
rect 1350 1972 1351 1976
rect 1355 1972 1356 1976
rect 1350 1971 1356 1972
rect 1454 1976 1460 1977
rect 1454 1972 1455 1976
rect 1459 1972 1460 1976
rect 1454 1971 1460 1972
rect 1558 1976 1564 1977
rect 1558 1972 1559 1976
rect 1563 1972 1564 1976
rect 1558 1971 1564 1972
rect 1654 1976 1660 1977
rect 1654 1972 1655 1976
rect 1659 1972 1660 1976
rect 1654 1971 1660 1972
rect 1742 1976 1748 1977
rect 1742 1972 1743 1976
rect 1747 1972 1748 1976
rect 1742 1971 1748 1972
rect 1822 1976 1828 1977
rect 1822 1972 1823 1976
rect 1827 1972 1828 1976
rect 1822 1971 1828 1972
rect 1894 1976 1900 1977
rect 1894 1972 1895 1976
rect 1899 1972 1900 1976
rect 1894 1971 1900 1972
rect 1958 1976 1964 1977
rect 1958 1972 1959 1976
rect 1963 1972 1964 1976
rect 1958 1971 1964 1972
rect 2022 1976 2028 1977
rect 2022 1972 2023 1976
rect 2027 1972 2028 1976
rect 2022 1971 2028 1972
rect 2070 1976 2076 1977
rect 2070 1972 2071 1976
rect 2075 1972 2076 1976
rect 2118 1975 2119 1979
rect 2123 1975 2124 1979
rect 2118 1974 2124 1975
rect 2070 1971 2076 1972
rect 110 1964 116 1965
rect 110 1960 111 1964
rect 115 1960 116 1964
rect 110 1959 116 1960
rect 1094 1964 1100 1965
rect 1094 1960 1095 1964
rect 1099 1960 1100 1964
rect 1094 1959 1100 1960
rect 158 1956 164 1957
rect 158 1952 159 1956
rect 163 1952 164 1956
rect 158 1951 164 1952
rect 230 1956 236 1957
rect 230 1952 231 1956
rect 235 1952 236 1956
rect 230 1951 236 1952
rect 302 1956 308 1957
rect 302 1952 303 1956
rect 307 1952 308 1956
rect 302 1951 308 1952
rect 374 1956 380 1957
rect 374 1952 375 1956
rect 379 1952 380 1956
rect 374 1951 380 1952
rect 446 1956 452 1957
rect 446 1952 447 1956
rect 451 1952 452 1956
rect 446 1951 452 1952
rect 526 1956 532 1957
rect 526 1952 527 1956
rect 531 1952 532 1956
rect 526 1951 532 1952
rect 606 1956 612 1957
rect 606 1952 607 1956
rect 611 1952 612 1956
rect 606 1951 612 1952
rect 686 1956 692 1957
rect 686 1952 687 1956
rect 691 1952 692 1956
rect 686 1951 692 1952
rect 758 1956 764 1957
rect 758 1952 759 1956
rect 763 1952 764 1956
rect 758 1951 764 1952
rect 830 1956 836 1957
rect 830 1952 831 1956
rect 835 1952 836 1956
rect 830 1951 836 1952
rect 910 1956 916 1957
rect 910 1952 911 1956
rect 915 1952 916 1956
rect 910 1951 916 1952
rect 990 1956 996 1957
rect 990 1952 991 1956
rect 995 1952 996 1956
rect 990 1951 996 1952
rect 1358 1952 1364 1953
rect 1134 1949 1140 1950
rect 1134 1945 1135 1949
rect 1139 1945 1140 1949
rect 1358 1948 1359 1952
rect 1363 1948 1364 1952
rect 1358 1947 1364 1948
rect 1422 1952 1428 1953
rect 1422 1948 1423 1952
rect 1427 1948 1428 1952
rect 1422 1947 1428 1948
rect 1486 1952 1492 1953
rect 1486 1948 1487 1952
rect 1491 1948 1492 1952
rect 1486 1947 1492 1948
rect 1558 1952 1564 1953
rect 1558 1948 1559 1952
rect 1563 1948 1564 1952
rect 1558 1947 1564 1948
rect 1630 1952 1636 1953
rect 1630 1948 1631 1952
rect 1635 1948 1636 1952
rect 1630 1947 1636 1948
rect 1702 1952 1708 1953
rect 1702 1948 1703 1952
rect 1707 1948 1708 1952
rect 1702 1947 1708 1948
rect 1774 1952 1780 1953
rect 1774 1948 1775 1952
rect 1779 1948 1780 1952
rect 1774 1947 1780 1948
rect 1846 1952 1852 1953
rect 1846 1948 1847 1952
rect 1851 1948 1852 1952
rect 1846 1947 1852 1948
rect 1926 1952 1932 1953
rect 1926 1948 1927 1952
rect 1931 1948 1932 1952
rect 1926 1947 1932 1948
rect 2006 1952 2012 1953
rect 2006 1948 2007 1952
rect 2011 1948 2012 1952
rect 2006 1947 2012 1948
rect 2070 1952 2076 1953
rect 2070 1948 2071 1952
rect 2075 1948 2076 1952
rect 2070 1947 2076 1948
rect 2118 1949 2124 1950
rect 1134 1944 1140 1945
rect 2118 1945 2119 1949
rect 2123 1945 2124 1949
rect 2118 1944 2124 1945
rect 1134 1932 1140 1933
rect 1134 1928 1135 1932
rect 1139 1928 1140 1932
rect 1134 1927 1140 1928
rect 2118 1932 2124 1933
rect 2118 1928 2119 1932
rect 2123 1928 2124 1932
rect 2118 1927 2124 1928
rect 1358 1924 1364 1925
rect 1358 1920 1359 1924
rect 1363 1920 1364 1924
rect 1358 1919 1364 1920
rect 1422 1924 1428 1925
rect 1422 1920 1423 1924
rect 1427 1920 1428 1924
rect 1422 1919 1428 1920
rect 1486 1924 1492 1925
rect 1486 1920 1487 1924
rect 1491 1920 1492 1924
rect 1486 1919 1492 1920
rect 1558 1924 1564 1925
rect 1558 1920 1559 1924
rect 1563 1920 1564 1924
rect 1558 1919 1564 1920
rect 1630 1924 1636 1925
rect 1630 1920 1631 1924
rect 1635 1920 1636 1924
rect 1630 1919 1636 1920
rect 1702 1924 1708 1925
rect 1702 1920 1703 1924
rect 1707 1920 1708 1924
rect 1702 1919 1708 1920
rect 1774 1924 1780 1925
rect 1774 1920 1775 1924
rect 1779 1920 1780 1924
rect 1774 1919 1780 1920
rect 1846 1924 1852 1925
rect 1846 1920 1847 1924
rect 1851 1920 1852 1924
rect 1846 1919 1852 1920
rect 1926 1924 1932 1925
rect 1926 1920 1927 1924
rect 1931 1920 1932 1924
rect 1926 1919 1932 1920
rect 2006 1924 2012 1925
rect 2006 1920 2007 1924
rect 2011 1920 2012 1924
rect 2006 1919 2012 1920
rect 2070 1924 2076 1925
rect 2070 1920 2071 1924
rect 2075 1920 2076 1924
rect 2070 1919 2076 1920
rect 134 1916 140 1917
rect 134 1912 135 1916
rect 139 1912 140 1916
rect 134 1911 140 1912
rect 174 1916 180 1917
rect 174 1912 175 1916
rect 179 1912 180 1916
rect 174 1911 180 1912
rect 230 1916 236 1917
rect 230 1912 231 1916
rect 235 1912 236 1916
rect 230 1911 236 1912
rect 294 1916 300 1917
rect 294 1912 295 1916
rect 299 1912 300 1916
rect 294 1911 300 1912
rect 366 1916 372 1917
rect 366 1912 367 1916
rect 371 1912 372 1916
rect 366 1911 372 1912
rect 446 1916 452 1917
rect 446 1912 447 1916
rect 451 1912 452 1916
rect 446 1911 452 1912
rect 526 1916 532 1917
rect 526 1912 527 1916
rect 531 1912 532 1916
rect 526 1911 532 1912
rect 614 1916 620 1917
rect 614 1912 615 1916
rect 619 1912 620 1916
rect 614 1911 620 1912
rect 702 1916 708 1917
rect 702 1912 703 1916
rect 707 1912 708 1916
rect 702 1911 708 1912
rect 790 1916 796 1917
rect 790 1912 791 1916
rect 795 1912 796 1916
rect 790 1911 796 1912
rect 878 1916 884 1917
rect 878 1912 879 1916
rect 883 1912 884 1916
rect 878 1911 884 1912
rect 110 1908 116 1909
rect 110 1904 111 1908
rect 115 1904 116 1908
rect 110 1903 116 1904
rect 1094 1908 1100 1909
rect 1094 1904 1095 1908
rect 1099 1904 1100 1908
rect 1094 1903 1100 1904
rect 110 1891 116 1892
rect 110 1887 111 1891
rect 115 1887 116 1891
rect 1094 1891 1100 1892
rect 110 1886 116 1887
rect 134 1888 140 1889
rect 134 1884 135 1888
rect 139 1884 140 1888
rect 134 1883 140 1884
rect 174 1888 180 1889
rect 174 1884 175 1888
rect 179 1884 180 1888
rect 174 1883 180 1884
rect 230 1888 236 1889
rect 230 1884 231 1888
rect 235 1884 236 1888
rect 230 1883 236 1884
rect 294 1888 300 1889
rect 294 1884 295 1888
rect 299 1884 300 1888
rect 294 1883 300 1884
rect 366 1888 372 1889
rect 366 1884 367 1888
rect 371 1884 372 1888
rect 366 1883 372 1884
rect 446 1888 452 1889
rect 446 1884 447 1888
rect 451 1884 452 1888
rect 446 1883 452 1884
rect 526 1888 532 1889
rect 526 1884 527 1888
rect 531 1884 532 1888
rect 526 1883 532 1884
rect 614 1888 620 1889
rect 614 1884 615 1888
rect 619 1884 620 1888
rect 614 1883 620 1884
rect 702 1888 708 1889
rect 702 1884 703 1888
rect 707 1884 708 1888
rect 702 1883 708 1884
rect 790 1888 796 1889
rect 790 1884 791 1888
rect 795 1884 796 1888
rect 790 1883 796 1884
rect 878 1888 884 1889
rect 878 1884 879 1888
rect 883 1884 884 1888
rect 1094 1887 1095 1891
rect 1099 1887 1100 1891
rect 1094 1886 1100 1887
rect 1230 1888 1236 1889
rect 878 1883 884 1884
rect 1230 1884 1231 1888
rect 1235 1884 1236 1888
rect 1230 1883 1236 1884
rect 1270 1888 1276 1889
rect 1270 1884 1271 1888
rect 1275 1884 1276 1888
rect 1270 1883 1276 1884
rect 1318 1888 1324 1889
rect 1318 1884 1319 1888
rect 1323 1884 1324 1888
rect 1318 1883 1324 1884
rect 1374 1888 1380 1889
rect 1374 1884 1375 1888
rect 1379 1884 1380 1888
rect 1374 1883 1380 1884
rect 1438 1888 1444 1889
rect 1438 1884 1439 1888
rect 1443 1884 1444 1888
rect 1438 1883 1444 1884
rect 1502 1888 1508 1889
rect 1502 1884 1503 1888
rect 1507 1884 1508 1888
rect 1502 1883 1508 1884
rect 1574 1888 1580 1889
rect 1574 1884 1575 1888
rect 1579 1884 1580 1888
rect 1574 1883 1580 1884
rect 1654 1888 1660 1889
rect 1654 1884 1655 1888
rect 1659 1884 1660 1888
rect 1654 1883 1660 1884
rect 1750 1888 1756 1889
rect 1750 1884 1751 1888
rect 1755 1884 1756 1888
rect 1750 1883 1756 1884
rect 1862 1888 1868 1889
rect 1862 1884 1863 1888
rect 1867 1884 1868 1888
rect 1862 1883 1868 1884
rect 1974 1888 1980 1889
rect 1974 1884 1975 1888
rect 1979 1884 1980 1888
rect 1974 1883 1980 1884
rect 2070 1888 2076 1889
rect 2070 1884 2071 1888
rect 2075 1884 2076 1888
rect 2070 1883 2076 1884
rect 1134 1880 1140 1881
rect 1134 1876 1135 1880
rect 1139 1876 1140 1880
rect 1134 1875 1140 1876
rect 2118 1880 2124 1881
rect 2118 1876 2119 1880
rect 2123 1876 2124 1880
rect 2118 1875 2124 1876
rect 134 1872 140 1873
rect 110 1869 116 1870
rect 110 1865 111 1869
rect 115 1865 116 1869
rect 134 1868 135 1872
rect 139 1868 140 1872
rect 134 1867 140 1868
rect 174 1872 180 1873
rect 174 1868 175 1872
rect 179 1868 180 1872
rect 174 1867 180 1868
rect 222 1872 228 1873
rect 222 1868 223 1872
rect 227 1868 228 1872
rect 222 1867 228 1868
rect 286 1872 292 1873
rect 286 1868 287 1872
rect 291 1868 292 1872
rect 286 1867 292 1868
rect 358 1872 364 1873
rect 358 1868 359 1872
rect 363 1868 364 1872
rect 358 1867 364 1868
rect 430 1872 436 1873
rect 430 1868 431 1872
rect 435 1868 436 1872
rect 430 1867 436 1868
rect 502 1872 508 1873
rect 502 1868 503 1872
rect 507 1868 508 1872
rect 502 1867 508 1868
rect 566 1872 572 1873
rect 566 1868 567 1872
rect 571 1868 572 1872
rect 566 1867 572 1868
rect 630 1872 636 1873
rect 630 1868 631 1872
rect 635 1868 636 1872
rect 630 1867 636 1868
rect 694 1872 700 1873
rect 694 1868 695 1872
rect 699 1868 700 1872
rect 694 1867 700 1868
rect 758 1872 764 1873
rect 758 1868 759 1872
rect 763 1868 764 1872
rect 758 1867 764 1868
rect 830 1872 836 1873
rect 830 1868 831 1872
rect 835 1868 836 1872
rect 830 1867 836 1868
rect 1094 1869 1100 1870
rect 110 1864 116 1865
rect 1094 1865 1095 1869
rect 1099 1865 1100 1869
rect 1094 1864 1100 1865
rect 1134 1863 1140 1864
rect 1134 1859 1135 1863
rect 1139 1859 1140 1863
rect 2118 1863 2124 1864
rect 1134 1858 1140 1859
rect 1230 1860 1236 1861
rect 1230 1856 1231 1860
rect 1235 1856 1236 1860
rect 1230 1855 1236 1856
rect 1270 1860 1276 1861
rect 1270 1856 1271 1860
rect 1275 1856 1276 1860
rect 1270 1855 1276 1856
rect 1318 1860 1324 1861
rect 1318 1856 1319 1860
rect 1323 1856 1324 1860
rect 1318 1855 1324 1856
rect 1374 1860 1380 1861
rect 1374 1856 1375 1860
rect 1379 1856 1380 1860
rect 1374 1855 1380 1856
rect 1438 1860 1444 1861
rect 1438 1856 1439 1860
rect 1443 1856 1444 1860
rect 1438 1855 1444 1856
rect 1502 1860 1508 1861
rect 1502 1856 1503 1860
rect 1507 1856 1508 1860
rect 1502 1855 1508 1856
rect 1574 1860 1580 1861
rect 1574 1856 1575 1860
rect 1579 1856 1580 1860
rect 1574 1855 1580 1856
rect 1654 1860 1660 1861
rect 1654 1856 1655 1860
rect 1659 1856 1660 1860
rect 1654 1855 1660 1856
rect 1750 1860 1756 1861
rect 1750 1856 1751 1860
rect 1755 1856 1756 1860
rect 1750 1855 1756 1856
rect 1862 1860 1868 1861
rect 1862 1856 1863 1860
rect 1867 1856 1868 1860
rect 1862 1855 1868 1856
rect 1974 1860 1980 1861
rect 1974 1856 1975 1860
rect 1979 1856 1980 1860
rect 1974 1855 1980 1856
rect 2070 1860 2076 1861
rect 2070 1856 2071 1860
rect 2075 1856 2076 1860
rect 2118 1859 2119 1863
rect 2123 1859 2124 1863
rect 2118 1858 2124 1859
rect 2070 1855 2076 1856
rect 110 1852 116 1853
rect 110 1848 111 1852
rect 115 1848 116 1852
rect 110 1847 116 1848
rect 1094 1852 1100 1853
rect 1094 1848 1095 1852
rect 1099 1848 1100 1852
rect 1094 1847 1100 1848
rect 134 1844 140 1845
rect 134 1840 135 1844
rect 139 1840 140 1844
rect 134 1839 140 1840
rect 174 1844 180 1845
rect 174 1840 175 1844
rect 179 1840 180 1844
rect 174 1839 180 1840
rect 222 1844 228 1845
rect 222 1840 223 1844
rect 227 1840 228 1844
rect 222 1839 228 1840
rect 286 1844 292 1845
rect 286 1840 287 1844
rect 291 1840 292 1844
rect 286 1839 292 1840
rect 358 1844 364 1845
rect 358 1840 359 1844
rect 363 1840 364 1844
rect 358 1839 364 1840
rect 430 1844 436 1845
rect 430 1840 431 1844
rect 435 1840 436 1844
rect 430 1839 436 1840
rect 502 1844 508 1845
rect 502 1840 503 1844
rect 507 1840 508 1844
rect 502 1839 508 1840
rect 566 1844 572 1845
rect 566 1840 567 1844
rect 571 1840 572 1844
rect 566 1839 572 1840
rect 630 1844 636 1845
rect 630 1840 631 1844
rect 635 1840 636 1844
rect 630 1839 636 1840
rect 694 1844 700 1845
rect 694 1840 695 1844
rect 699 1840 700 1844
rect 694 1839 700 1840
rect 758 1844 764 1845
rect 758 1840 759 1844
rect 763 1840 764 1844
rect 758 1839 764 1840
rect 830 1844 836 1845
rect 830 1840 831 1844
rect 835 1840 836 1844
rect 1158 1844 1164 1845
rect 830 1839 836 1840
rect 1134 1841 1140 1842
rect 1134 1837 1135 1841
rect 1139 1837 1140 1841
rect 1158 1840 1159 1844
rect 1163 1840 1164 1844
rect 1158 1839 1164 1840
rect 1198 1844 1204 1845
rect 1198 1840 1199 1844
rect 1203 1840 1204 1844
rect 1198 1839 1204 1840
rect 1238 1844 1244 1845
rect 1238 1840 1239 1844
rect 1243 1840 1244 1844
rect 1238 1839 1244 1840
rect 1302 1844 1308 1845
rect 1302 1840 1303 1844
rect 1307 1840 1308 1844
rect 1302 1839 1308 1840
rect 1366 1844 1372 1845
rect 1366 1840 1367 1844
rect 1371 1840 1372 1844
rect 1366 1839 1372 1840
rect 1430 1844 1436 1845
rect 1430 1840 1431 1844
rect 1435 1840 1436 1844
rect 1430 1839 1436 1840
rect 1502 1844 1508 1845
rect 1502 1840 1503 1844
rect 1507 1840 1508 1844
rect 1502 1839 1508 1840
rect 1582 1844 1588 1845
rect 1582 1840 1583 1844
rect 1587 1840 1588 1844
rect 1582 1839 1588 1840
rect 1670 1844 1676 1845
rect 1670 1840 1671 1844
rect 1675 1840 1676 1844
rect 1670 1839 1676 1840
rect 1766 1844 1772 1845
rect 1766 1840 1767 1844
rect 1771 1840 1772 1844
rect 1766 1839 1772 1840
rect 1870 1844 1876 1845
rect 1870 1840 1871 1844
rect 1875 1840 1876 1844
rect 1870 1839 1876 1840
rect 1982 1844 1988 1845
rect 1982 1840 1983 1844
rect 1987 1840 1988 1844
rect 1982 1839 1988 1840
rect 2070 1844 2076 1845
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2070 1839 2076 1840
rect 2118 1841 2124 1842
rect 1134 1836 1140 1837
rect 2118 1837 2119 1841
rect 2123 1837 2124 1841
rect 2118 1836 2124 1837
rect 1134 1824 1140 1825
rect 1134 1820 1135 1824
rect 1139 1820 1140 1824
rect 1134 1819 1140 1820
rect 2118 1824 2124 1825
rect 2118 1820 2119 1824
rect 2123 1820 2124 1824
rect 2118 1819 2124 1820
rect 1158 1816 1164 1817
rect 1158 1812 1159 1816
rect 1163 1812 1164 1816
rect 1158 1811 1164 1812
rect 1198 1816 1204 1817
rect 1198 1812 1199 1816
rect 1203 1812 1204 1816
rect 1198 1811 1204 1812
rect 1238 1816 1244 1817
rect 1238 1812 1239 1816
rect 1243 1812 1244 1816
rect 1238 1811 1244 1812
rect 1302 1816 1308 1817
rect 1302 1812 1303 1816
rect 1307 1812 1308 1816
rect 1302 1811 1308 1812
rect 1366 1816 1372 1817
rect 1366 1812 1367 1816
rect 1371 1812 1372 1816
rect 1366 1811 1372 1812
rect 1430 1816 1436 1817
rect 1430 1812 1431 1816
rect 1435 1812 1436 1816
rect 1430 1811 1436 1812
rect 1502 1816 1508 1817
rect 1502 1812 1503 1816
rect 1507 1812 1508 1816
rect 1502 1811 1508 1812
rect 1582 1816 1588 1817
rect 1582 1812 1583 1816
rect 1587 1812 1588 1816
rect 1582 1811 1588 1812
rect 1670 1816 1676 1817
rect 1670 1812 1671 1816
rect 1675 1812 1676 1816
rect 1670 1811 1676 1812
rect 1766 1816 1772 1817
rect 1766 1812 1767 1816
rect 1771 1812 1772 1816
rect 1766 1811 1772 1812
rect 1870 1816 1876 1817
rect 1870 1812 1871 1816
rect 1875 1812 1876 1816
rect 1870 1811 1876 1812
rect 1982 1816 1988 1817
rect 1982 1812 1983 1816
rect 1987 1812 1988 1816
rect 1982 1811 1988 1812
rect 2070 1816 2076 1817
rect 2070 1812 2071 1816
rect 2075 1812 2076 1816
rect 2070 1811 2076 1812
rect 134 1804 140 1805
rect 134 1800 135 1804
rect 139 1800 140 1804
rect 134 1799 140 1800
rect 182 1804 188 1805
rect 182 1800 183 1804
rect 187 1800 188 1804
rect 182 1799 188 1800
rect 262 1804 268 1805
rect 262 1800 263 1804
rect 267 1800 268 1804
rect 262 1799 268 1800
rect 350 1804 356 1805
rect 350 1800 351 1804
rect 355 1800 356 1804
rect 350 1799 356 1800
rect 438 1804 444 1805
rect 438 1800 439 1804
rect 443 1800 444 1804
rect 438 1799 444 1800
rect 526 1804 532 1805
rect 526 1800 527 1804
rect 531 1800 532 1804
rect 526 1799 532 1800
rect 606 1804 612 1805
rect 606 1800 607 1804
rect 611 1800 612 1804
rect 606 1799 612 1800
rect 686 1804 692 1805
rect 686 1800 687 1804
rect 691 1800 692 1804
rect 686 1799 692 1800
rect 766 1804 772 1805
rect 766 1800 767 1804
rect 771 1800 772 1804
rect 766 1799 772 1800
rect 838 1804 844 1805
rect 838 1800 839 1804
rect 843 1800 844 1804
rect 838 1799 844 1800
rect 910 1804 916 1805
rect 910 1800 911 1804
rect 915 1800 916 1804
rect 910 1799 916 1800
rect 990 1804 996 1805
rect 990 1800 991 1804
rect 995 1800 996 1804
rect 990 1799 996 1800
rect 1046 1804 1052 1805
rect 1046 1800 1047 1804
rect 1051 1800 1052 1804
rect 1046 1799 1052 1800
rect 110 1796 116 1797
rect 110 1792 111 1796
rect 115 1792 116 1796
rect 110 1791 116 1792
rect 1094 1796 1100 1797
rect 1094 1792 1095 1796
rect 1099 1792 1100 1796
rect 1094 1791 1100 1792
rect 110 1779 116 1780
rect 110 1775 111 1779
rect 115 1775 116 1779
rect 1094 1779 1100 1780
rect 110 1774 116 1775
rect 134 1776 140 1777
rect 134 1772 135 1776
rect 139 1772 140 1776
rect 134 1771 140 1772
rect 182 1776 188 1777
rect 182 1772 183 1776
rect 187 1772 188 1776
rect 182 1771 188 1772
rect 262 1776 268 1777
rect 262 1772 263 1776
rect 267 1772 268 1776
rect 262 1771 268 1772
rect 350 1776 356 1777
rect 350 1772 351 1776
rect 355 1772 356 1776
rect 350 1771 356 1772
rect 438 1776 444 1777
rect 438 1772 439 1776
rect 443 1772 444 1776
rect 438 1771 444 1772
rect 526 1776 532 1777
rect 526 1772 527 1776
rect 531 1772 532 1776
rect 526 1771 532 1772
rect 606 1776 612 1777
rect 606 1772 607 1776
rect 611 1772 612 1776
rect 606 1771 612 1772
rect 686 1776 692 1777
rect 686 1772 687 1776
rect 691 1772 692 1776
rect 686 1771 692 1772
rect 766 1776 772 1777
rect 766 1772 767 1776
rect 771 1772 772 1776
rect 766 1771 772 1772
rect 838 1776 844 1777
rect 838 1772 839 1776
rect 843 1772 844 1776
rect 838 1771 844 1772
rect 910 1776 916 1777
rect 910 1772 911 1776
rect 915 1772 916 1776
rect 910 1771 916 1772
rect 990 1776 996 1777
rect 990 1772 991 1776
rect 995 1772 996 1776
rect 990 1771 996 1772
rect 1046 1776 1052 1777
rect 1046 1772 1047 1776
rect 1051 1772 1052 1776
rect 1094 1775 1095 1779
rect 1099 1775 1100 1779
rect 1094 1774 1100 1775
rect 1046 1771 1052 1772
rect 1310 1772 1316 1773
rect 1310 1768 1311 1772
rect 1315 1768 1316 1772
rect 1310 1767 1316 1768
rect 1350 1772 1356 1773
rect 1350 1768 1351 1772
rect 1355 1768 1356 1772
rect 1350 1767 1356 1768
rect 1390 1772 1396 1773
rect 1390 1768 1391 1772
rect 1395 1768 1396 1772
rect 1390 1767 1396 1768
rect 1430 1772 1436 1773
rect 1430 1768 1431 1772
rect 1435 1768 1436 1772
rect 1430 1767 1436 1768
rect 1470 1772 1476 1773
rect 1470 1768 1471 1772
rect 1475 1768 1476 1772
rect 1470 1767 1476 1768
rect 1510 1772 1516 1773
rect 1510 1768 1511 1772
rect 1515 1768 1516 1772
rect 1510 1767 1516 1768
rect 1550 1772 1556 1773
rect 1550 1768 1551 1772
rect 1555 1768 1556 1772
rect 1550 1767 1556 1768
rect 1606 1772 1612 1773
rect 1606 1768 1607 1772
rect 1611 1768 1612 1772
rect 1606 1767 1612 1768
rect 1678 1772 1684 1773
rect 1678 1768 1679 1772
rect 1683 1768 1684 1772
rect 1678 1767 1684 1768
rect 1766 1772 1772 1773
rect 1766 1768 1767 1772
rect 1771 1768 1772 1772
rect 1766 1767 1772 1768
rect 1870 1772 1876 1773
rect 1870 1768 1871 1772
rect 1875 1768 1876 1772
rect 1870 1767 1876 1768
rect 1982 1772 1988 1773
rect 1982 1768 1983 1772
rect 1987 1768 1988 1772
rect 1982 1767 1988 1768
rect 2070 1772 2076 1773
rect 2070 1768 2071 1772
rect 2075 1768 2076 1772
rect 2070 1767 2076 1768
rect 1134 1764 1140 1765
rect 1134 1760 1135 1764
rect 1139 1760 1140 1764
rect 1134 1759 1140 1760
rect 2118 1764 2124 1765
rect 2118 1760 2119 1764
rect 2123 1760 2124 1764
rect 2118 1759 2124 1760
rect 134 1756 140 1757
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 134 1752 135 1756
rect 139 1752 140 1756
rect 134 1751 140 1752
rect 198 1756 204 1757
rect 198 1752 199 1756
rect 203 1752 204 1756
rect 198 1751 204 1752
rect 294 1756 300 1757
rect 294 1752 295 1756
rect 299 1752 300 1756
rect 294 1751 300 1752
rect 398 1756 404 1757
rect 398 1752 399 1756
rect 403 1752 404 1756
rect 398 1751 404 1752
rect 494 1756 500 1757
rect 494 1752 495 1756
rect 499 1752 500 1756
rect 494 1751 500 1752
rect 590 1756 596 1757
rect 590 1752 591 1756
rect 595 1752 596 1756
rect 590 1751 596 1752
rect 670 1756 676 1757
rect 670 1752 671 1756
rect 675 1752 676 1756
rect 670 1751 676 1752
rect 750 1756 756 1757
rect 750 1752 751 1756
rect 755 1752 756 1756
rect 750 1751 756 1752
rect 822 1756 828 1757
rect 822 1752 823 1756
rect 827 1752 828 1756
rect 822 1751 828 1752
rect 886 1756 892 1757
rect 886 1752 887 1756
rect 891 1752 892 1756
rect 886 1751 892 1752
rect 958 1756 964 1757
rect 958 1752 959 1756
rect 963 1752 964 1756
rect 958 1751 964 1752
rect 1030 1756 1036 1757
rect 1030 1752 1031 1756
rect 1035 1752 1036 1756
rect 1030 1751 1036 1752
rect 1094 1753 1100 1754
rect 110 1748 116 1749
rect 1094 1749 1095 1753
rect 1099 1749 1100 1753
rect 1094 1748 1100 1749
rect 1134 1747 1140 1748
rect 1134 1743 1135 1747
rect 1139 1743 1140 1747
rect 2118 1747 2124 1748
rect 1134 1742 1140 1743
rect 1310 1744 1316 1745
rect 1310 1740 1311 1744
rect 1315 1740 1316 1744
rect 1310 1739 1316 1740
rect 1350 1744 1356 1745
rect 1350 1740 1351 1744
rect 1355 1740 1356 1744
rect 1350 1739 1356 1740
rect 1390 1744 1396 1745
rect 1390 1740 1391 1744
rect 1395 1740 1396 1744
rect 1390 1739 1396 1740
rect 1430 1744 1436 1745
rect 1430 1740 1431 1744
rect 1435 1740 1436 1744
rect 1430 1739 1436 1740
rect 1470 1744 1476 1745
rect 1470 1740 1471 1744
rect 1475 1740 1476 1744
rect 1470 1739 1476 1740
rect 1510 1744 1516 1745
rect 1510 1740 1511 1744
rect 1515 1740 1516 1744
rect 1510 1739 1516 1740
rect 1550 1744 1556 1745
rect 1550 1740 1551 1744
rect 1555 1740 1556 1744
rect 1550 1739 1556 1740
rect 1606 1744 1612 1745
rect 1606 1740 1607 1744
rect 1611 1740 1612 1744
rect 1606 1739 1612 1740
rect 1678 1744 1684 1745
rect 1678 1740 1679 1744
rect 1683 1740 1684 1744
rect 1678 1739 1684 1740
rect 1766 1744 1772 1745
rect 1766 1740 1767 1744
rect 1771 1740 1772 1744
rect 1766 1739 1772 1740
rect 1870 1744 1876 1745
rect 1870 1740 1871 1744
rect 1875 1740 1876 1744
rect 1870 1739 1876 1740
rect 1982 1744 1988 1745
rect 1982 1740 1983 1744
rect 1987 1740 1988 1744
rect 1982 1739 1988 1740
rect 2070 1744 2076 1745
rect 2070 1740 2071 1744
rect 2075 1740 2076 1744
rect 2118 1743 2119 1747
rect 2123 1743 2124 1747
rect 2118 1742 2124 1743
rect 2070 1739 2076 1740
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 1094 1736 1100 1737
rect 1094 1732 1095 1736
rect 1099 1732 1100 1736
rect 1094 1731 1100 1732
rect 134 1728 140 1729
rect 134 1724 135 1728
rect 139 1724 140 1728
rect 134 1723 140 1724
rect 198 1728 204 1729
rect 198 1724 199 1728
rect 203 1724 204 1728
rect 198 1723 204 1724
rect 294 1728 300 1729
rect 294 1724 295 1728
rect 299 1724 300 1728
rect 294 1723 300 1724
rect 398 1728 404 1729
rect 398 1724 399 1728
rect 403 1724 404 1728
rect 398 1723 404 1724
rect 494 1728 500 1729
rect 494 1724 495 1728
rect 499 1724 500 1728
rect 494 1723 500 1724
rect 590 1728 596 1729
rect 590 1724 591 1728
rect 595 1724 596 1728
rect 590 1723 596 1724
rect 670 1728 676 1729
rect 670 1724 671 1728
rect 675 1724 676 1728
rect 670 1723 676 1724
rect 750 1728 756 1729
rect 750 1724 751 1728
rect 755 1724 756 1728
rect 750 1723 756 1724
rect 822 1728 828 1729
rect 822 1724 823 1728
rect 827 1724 828 1728
rect 822 1723 828 1724
rect 886 1728 892 1729
rect 886 1724 887 1728
rect 891 1724 892 1728
rect 886 1723 892 1724
rect 958 1728 964 1729
rect 958 1724 959 1728
rect 963 1724 964 1728
rect 958 1723 964 1724
rect 1030 1728 1036 1729
rect 1030 1724 1031 1728
rect 1035 1724 1036 1728
rect 1262 1728 1268 1729
rect 1030 1723 1036 1724
rect 1134 1725 1140 1726
rect 1134 1721 1135 1725
rect 1139 1721 1140 1725
rect 1262 1724 1263 1728
rect 1267 1724 1268 1728
rect 1262 1723 1268 1724
rect 1318 1728 1324 1729
rect 1318 1724 1319 1728
rect 1323 1724 1324 1728
rect 1318 1723 1324 1724
rect 1382 1728 1388 1729
rect 1382 1724 1383 1728
rect 1387 1724 1388 1728
rect 1382 1723 1388 1724
rect 1454 1728 1460 1729
rect 1454 1724 1455 1728
rect 1459 1724 1460 1728
rect 1454 1723 1460 1724
rect 1534 1728 1540 1729
rect 1534 1724 1535 1728
rect 1539 1724 1540 1728
rect 1534 1723 1540 1724
rect 1614 1728 1620 1729
rect 1614 1724 1615 1728
rect 1619 1724 1620 1728
rect 1614 1723 1620 1724
rect 1686 1728 1692 1729
rect 1686 1724 1687 1728
rect 1691 1724 1692 1728
rect 1686 1723 1692 1724
rect 1758 1728 1764 1729
rect 1758 1724 1759 1728
rect 1763 1724 1764 1728
rect 1758 1723 1764 1724
rect 1830 1728 1836 1729
rect 1830 1724 1831 1728
rect 1835 1724 1836 1728
rect 1830 1723 1836 1724
rect 1894 1728 1900 1729
rect 1894 1724 1895 1728
rect 1899 1724 1900 1728
rect 1894 1723 1900 1724
rect 1958 1728 1964 1729
rect 1958 1724 1959 1728
rect 1963 1724 1964 1728
rect 1958 1723 1964 1724
rect 2022 1728 2028 1729
rect 2022 1724 2023 1728
rect 2027 1724 2028 1728
rect 2022 1723 2028 1724
rect 2070 1728 2076 1729
rect 2070 1724 2071 1728
rect 2075 1724 2076 1728
rect 2070 1723 2076 1724
rect 2118 1725 2124 1726
rect 1134 1720 1140 1721
rect 2118 1721 2119 1725
rect 2123 1721 2124 1725
rect 2118 1720 2124 1721
rect 1134 1708 1140 1709
rect 1134 1704 1135 1708
rect 1139 1704 1140 1708
rect 1134 1703 1140 1704
rect 2118 1708 2124 1709
rect 2118 1704 2119 1708
rect 2123 1704 2124 1708
rect 2118 1703 2124 1704
rect 1262 1700 1268 1701
rect 1262 1696 1263 1700
rect 1267 1696 1268 1700
rect 1262 1695 1268 1696
rect 1318 1700 1324 1701
rect 1318 1696 1319 1700
rect 1323 1696 1324 1700
rect 1318 1695 1324 1696
rect 1382 1700 1388 1701
rect 1382 1696 1383 1700
rect 1387 1696 1388 1700
rect 1382 1695 1388 1696
rect 1454 1700 1460 1701
rect 1454 1696 1455 1700
rect 1459 1696 1460 1700
rect 1454 1695 1460 1696
rect 1534 1700 1540 1701
rect 1534 1696 1535 1700
rect 1539 1696 1540 1700
rect 1534 1695 1540 1696
rect 1614 1700 1620 1701
rect 1614 1696 1615 1700
rect 1619 1696 1620 1700
rect 1614 1695 1620 1696
rect 1686 1700 1692 1701
rect 1686 1696 1687 1700
rect 1691 1696 1692 1700
rect 1686 1695 1692 1696
rect 1758 1700 1764 1701
rect 1758 1696 1759 1700
rect 1763 1696 1764 1700
rect 1758 1695 1764 1696
rect 1830 1700 1836 1701
rect 1830 1696 1831 1700
rect 1835 1696 1836 1700
rect 1830 1695 1836 1696
rect 1894 1700 1900 1701
rect 1894 1696 1895 1700
rect 1899 1696 1900 1700
rect 1894 1695 1900 1696
rect 1958 1700 1964 1701
rect 1958 1696 1959 1700
rect 1963 1696 1964 1700
rect 1958 1695 1964 1696
rect 2022 1700 2028 1701
rect 2022 1696 2023 1700
rect 2027 1696 2028 1700
rect 2022 1695 2028 1696
rect 2070 1700 2076 1701
rect 2070 1696 2071 1700
rect 2075 1696 2076 1700
rect 2070 1695 2076 1696
rect 150 1688 156 1689
rect 150 1684 151 1688
rect 155 1684 156 1688
rect 150 1683 156 1684
rect 222 1688 228 1689
rect 222 1684 223 1688
rect 227 1684 228 1688
rect 222 1683 228 1684
rect 302 1688 308 1689
rect 302 1684 303 1688
rect 307 1684 308 1688
rect 302 1683 308 1684
rect 382 1688 388 1689
rect 382 1684 383 1688
rect 387 1684 388 1688
rect 382 1683 388 1684
rect 462 1688 468 1689
rect 462 1684 463 1688
rect 467 1684 468 1688
rect 462 1683 468 1684
rect 534 1688 540 1689
rect 534 1684 535 1688
rect 539 1684 540 1688
rect 534 1683 540 1684
rect 606 1688 612 1689
rect 606 1684 607 1688
rect 611 1684 612 1688
rect 606 1683 612 1684
rect 670 1688 676 1689
rect 670 1684 671 1688
rect 675 1684 676 1688
rect 670 1683 676 1684
rect 734 1688 740 1689
rect 734 1684 735 1688
rect 739 1684 740 1688
rect 734 1683 740 1684
rect 806 1688 812 1689
rect 806 1684 807 1688
rect 811 1684 812 1688
rect 806 1683 812 1684
rect 878 1688 884 1689
rect 878 1684 879 1688
rect 883 1684 884 1688
rect 878 1683 884 1684
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 1094 1680 1100 1681
rect 1094 1676 1095 1680
rect 1099 1676 1100 1680
rect 1094 1675 1100 1676
rect 1166 1664 1172 1665
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 1094 1663 1100 1664
rect 110 1658 116 1659
rect 150 1660 156 1661
rect 150 1656 151 1660
rect 155 1656 156 1660
rect 150 1655 156 1656
rect 222 1660 228 1661
rect 222 1656 223 1660
rect 227 1656 228 1660
rect 222 1655 228 1656
rect 302 1660 308 1661
rect 302 1656 303 1660
rect 307 1656 308 1660
rect 302 1655 308 1656
rect 382 1660 388 1661
rect 382 1656 383 1660
rect 387 1656 388 1660
rect 382 1655 388 1656
rect 462 1660 468 1661
rect 462 1656 463 1660
rect 467 1656 468 1660
rect 462 1655 468 1656
rect 534 1660 540 1661
rect 534 1656 535 1660
rect 539 1656 540 1660
rect 534 1655 540 1656
rect 606 1660 612 1661
rect 606 1656 607 1660
rect 611 1656 612 1660
rect 606 1655 612 1656
rect 670 1660 676 1661
rect 670 1656 671 1660
rect 675 1656 676 1660
rect 670 1655 676 1656
rect 734 1660 740 1661
rect 734 1656 735 1660
rect 739 1656 740 1660
rect 734 1655 740 1656
rect 806 1660 812 1661
rect 806 1656 807 1660
rect 811 1656 812 1660
rect 806 1655 812 1656
rect 878 1660 884 1661
rect 878 1656 879 1660
rect 883 1656 884 1660
rect 1094 1659 1095 1663
rect 1099 1659 1100 1663
rect 1166 1660 1167 1664
rect 1171 1660 1172 1664
rect 1166 1659 1172 1660
rect 1246 1664 1252 1665
rect 1246 1660 1247 1664
rect 1251 1660 1252 1664
rect 1246 1659 1252 1660
rect 1334 1664 1340 1665
rect 1334 1660 1335 1664
rect 1339 1660 1340 1664
rect 1334 1659 1340 1660
rect 1422 1664 1428 1665
rect 1422 1660 1423 1664
rect 1427 1660 1428 1664
rect 1422 1659 1428 1660
rect 1510 1664 1516 1665
rect 1510 1660 1511 1664
rect 1515 1660 1516 1664
rect 1510 1659 1516 1660
rect 1598 1664 1604 1665
rect 1598 1660 1599 1664
rect 1603 1660 1604 1664
rect 1598 1659 1604 1660
rect 1678 1664 1684 1665
rect 1678 1660 1679 1664
rect 1683 1660 1684 1664
rect 1678 1659 1684 1660
rect 1750 1664 1756 1665
rect 1750 1660 1751 1664
rect 1755 1660 1756 1664
rect 1750 1659 1756 1660
rect 1814 1664 1820 1665
rect 1814 1660 1815 1664
rect 1819 1660 1820 1664
rect 1814 1659 1820 1660
rect 1870 1664 1876 1665
rect 1870 1660 1871 1664
rect 1875 1660 1876 1664
rect 1870 1659 1876 1660
rect 1926 1664 1932 1665
rect 1926 1660 1927 1664
rect 1931 1660 1932 1664
rect 1926 1659 1932 1660
rect 1982 1664 1988 1665
rect 1982 1660 1983 1664
rect 1987 1660 1988 1664
rect 1982 1659 1988 1660
rect 2030 1664 2036 1665
rect 2030 1660 2031 1664
rect 2035 1660 2036 1664
rect 2030 1659 2036 1660
rect 2070 1664 2076 1665
rect 2070 1660 2071 1664
rect 2075 1660 2076 1664
rect 2070 1659 2076 1660
rect 1094 1658 1100 1659
rect 878 1655 884 1656
rect 1134 1656 1140 1657
rect 1134 1652 1135 1656
rect 1139 1652 1140 1656
rect 1134 1651 1140 1652
rect 2118 1656 2124 1657
rect 2118 1652 2119 1656
rect 2123 1652 2124 1656
rect 2118 1651 2124 1652
rect 174 1644 180 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 174 1640 175 1644
rect 179 1640 180 1644
rect 174 1639 180 1640
rect 214 1644 220 1645
rect 214 1640 215 1644
rect 219 1640 220 1644
rect 214 1639 220 1640
rect 254 1644 260 1645
rect 254 1640 255 1644
rect 259 1640 260 1644
rect 254 1639 260 1640
rect 302 1644 308 1645
rect 302 1640 303 1644
rect 307 1640 308 1644
rect 302 1639 308 1640
rect 358 1644 364 1645
rect 358 1640 359 1644
rect 363 1640 364 1644
rect 358 1639 364 1640
rect 406 1644 412 1645
rect 406 1640 407 1644
rect 411 1640 412 1644
rect 406 1639 412 1640
rect 454 1644 460 1645
rect 454 1640 455 1644
rect 459 1640 460 1644
rect 454 1639 460 1640
rect 502 1644 508 1645
rect 502 1640 503 1644
rect 507 1640 508 1644
rect 502 1639 508 1640
rect 550 1644 556 1645
rect 550 1640 551 1644
rect 555 1640 556 1644
rect 550 1639 556 1640
rect 606 1644 612 1645
rect 606 1640 607 1644
rect 611 1640 612 1644
rect 606 1639 612 1640
rect 662 1644 668 1645
rect 662 1640 663 1644
rect 667 1640 668 1644
rect 662 1639 668 1640
rect 718 1644 724 1645
rect 718 1640 719 1644
rect 723 1640 724 1644
rect 718 1639 724 1640
rect 1094 1641 1100 1642
rect 110 1636 116 1637
rect 1094 1637 1095 1641
rect 1099 1637 1100 1641
rect 1094 1636 1100 1637
rect 1134 1639 1140 1640
rect 1134 1635 1135 1639
rect 1139 1635 1140 1639
rect 2118 1639 2124 1640
rect 1134 1634 1140 1635
rect 1166 1636 1172 1637
rect 1166 1632 1167 1636
rect 1171 1632 1172 1636
rect 1166 1631 1172 1632
rect 1246 1636 1252 1637
rect 1246 1632 1247 1636
rect 1251 1632 1252 1636
rect 1246 1631 1252 1632
rect 1334 1636 1340 1637
rect 1334 1632 1335 1636
rect 1339 1632 1340 1636
rect 1334 1631 1340 1632
rect 1422 1636 1428 1637
rect 1422 1632 1423 1636
rect 1427 1632 1428 1636
rect 1422 1631 1428 1632
rect 1510 1636 1516 1637
rect 1510 1632 1511 1636
rect 1515 1632 1516 1636
rect 1510 1631 1516 1632
rect 1598 1636 1604 1637
rect 1598 1632 1599 1636
rect 1603 1632 1604 1636
rect 1598 1631 1604 1632
rect 1678 1636 1684 1637
rect 1678 1632 1679 1636
rect 1683 1632 1684 1636
rect 1678 1631 1684 1632
rect 1750 1636 1756 1637
rect 1750 1632 1751 1636
rect 1755 1632 1756 1636
rect 1750 1631 1756 1632
rect 1814 1636 1820 1637
rect 1814 1632 1815 1636
rect 1819 1632 1820 1636
rect 1814 1631 1820 1632
rect 1870 1636 1876 1637
rect 1870 1632 1871 1636
rect 1875 1632 1876 1636
rect 1870 1631 1876 1632
rect 1926 1636 1932 1637
rect 1926 1632 1927 1636
rect 1931 1632 1932 1636
rect 1926 1631 1932 1632
rect 1982 1636 1988 1637
rect 1982 1632 1983 1636
rect 1987 1632 1988 1636
rect 1982 1631 1988 1632
rect 2030 1636 2036 1637
rect 2030 1632 2031 1636
rect 2035 1632 2036 1636
rect 2030 1631 2036 1632
rect 2070 1636 2076 1637
rect 2070 1632 2071 1636
rect 2075 1632 2076 1636
rect 2118 1635 2119 1639
rect 2123 1635 2124 1639
rect 2118 1634 2124 1635
rect 2070 1631 2076 1632
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 1094 1624 1100 1625
rect 1094 1620 1095 1624
rect 1099 1620 1100 1624
rect 1094 1619 1100 1620
rect 1158 1620 1164 1621
rect 1134 1617 1140 1618
rect 174 1616 180 1617
rect 174 1612 175 1616
rect 179 1612 180 1616
rect 174 1611 180 1612
rect 214 1616 220 1617
rect 214 1612 215 1616
rect 219 1612 220 1616
rect 214 1611 220 1612
rect 254 1616 260 1617
rect 254 1612 255 1616
rect 259 1612 260 1616
rect 254 1611 260 1612
rect 302 1616 308 1617
rect 302 1612 303 1616
rect 307 1612 308 1616
rect 302 1611 308 1612
rect 358 1616 364 1617
rect 358 1612 359 1616
rect 363 1612 364 1616
rect 358 1611 364 1612
rect 406 1616 412 1617
rect 406 1612 407 1616
rect 411 1612 412 1616
rect 406 1611 412 1612
rect 454 1616 460 1617
rect 454 1612 455 1616
rect 459 1612 460 1616
rect 454 1611 460 1612
rect 502 1616 508 1617
rect 502 1612 503 1616
rect 507 1612 508 1616
rect 502 1611 508 1612
rect 550 1616 556 1617
rect 550 1612 551 1616
rect 555 1612 556 1616
rect 550 1611 556 1612
rect 606 1616 612 1617
rect 606 1612 607 1616
rect 611 1612 612 1616
rect 606 1611 612 1612
rect 662 1616 668 1617
rect 662 1612 663 1616
rect 667 1612 668 1616
rect 662 1611 668 1612
rect 718 1616 724 1617
rect 718 1612 719 1616
rect 723 1612 724 1616
rect 1134 1613 1135 1617
rect 1139 1613 1140 1617
rect 1158 1616 1159 1620
rect 1163 1616 1164 1620
rect 1158 1615 1164 1616
rect 1198 1620 1204 1621
rect 1198 1616 1199 1620
rect 1203 1616 1204 1620
rect 1198 1615 1204 1616
rect 1246 1620 1252 1621
rect 1246 1616 1247 1620
rect 1251 1616 1252 1620
rect 1246 1615 1252 1616
rect 1318 1620 1324 1621
rect 1318 1616 1319 1620
rect 1323 1616 1324 1620
rect 1318 1615 1324 1616
rect 1390 1620 1396 1621
rect 1390 1616 1391 1620
rect 1395 1616 1396 1620
rect 1390 1615 1396 1616
rect 1462 1620 1468 1621
rect 1462 1616 1463 1620
rect 1467 1616 1468 1620
rect 1462 1615 1468 1616
rect 1534 1620 1540 1621
rect 1534 1616 1535 1620
rect 1539 1616 1540 1620
rect 1534 1615 1540 1616
rect 1606 1620 1612 1621
rect 1606 1616 1607 1620
rect 1611 1616 1612 1620
rect 1606 1615 1612 1616
rect 1678 1620 1684 1621
rect 1678 1616 1679 1620
rect 1683 1616 1684 1620
rect 1678 1615 1684 1616
rect 1750 1620 1756 1621
rect 1750 1616 1751 1620
rect 1755 1616 1756 1620
rect 1750 1615 1756 1616
rect 1830 1620 1836 1621
rect 1830 1616 1831 1620
rect 1835 1616 1836 1620
rect 1830 1615 1836 1616
rect 2118 1617 2124 1618
rect 1134 1612 1140 1613
rect 2118 1613 2119 1617
rect 2123 1613 2124 1617
rect 2118 1612 2124 1613
rect 718 1611 724 1612
rect 1134 1600 1140 1601
rect 1134 1596 1135 1600
rect 1139 1596 1140 1600
rect 1134 1595 1140 1596
rect 2118 1600 2124 1601
rect 2118 1596 2119 1600
rect 2123 1596 2124 1600
rect 2118 1595 2124 1596
rect 1158 1592 1164 1593
rect 1158 1588 1159 1592
rect 1163 1588 1164 1592
rect 1158 1587 1164 1588
rect 1198 1592 1204 1593
rect 1198 1588 1199 1592
rect 1203 1588 1204 1592
rect 1198 1587 1204 1588
rect 1246 1592 1252 1593
rect 1246 1588 1247 1592
rect 1251 1588 1252 1592
rect 1246 1587 1252 1588
rect 1318 1592 1324 1593
rect 1318 1588 1319 1592
rect 1323 1588 1324 1592
rect 1318 1587 1324 1588
rect 1390 1592 1396 1593
rect 1390 1588 1391 1592
rect 1395 1588 1396 1592
rect 1390 1587 1396 1588
rect 1462 1592 1468 1593
rect 1462 1588 1463 1592
rect 1467 1588 1468 1592
rect 1462 1587 1468 1588
rect 1534 1592 1540 1593
rect 1534 1588 1535 1592
rect 1539 1588 1540 1592
rect 1534 1587 1540 1588
rect 1606 1592 1612 1593
rect 1606 1588 1607 1592
rect 1611 1588 1612 1592
rect 1606 1587 1612 1588
rect 1678 1592 1684 1593
rect 1678 1588 1679 1592
rect 1683 1588 1684 1592
rect 1678 1587 1684 1588
rect 1750 1592 1756 1593
rect 1750 1588 1751 1592
rect 1755 1588 1756 1592
rect 1750 1587 1756 1588
rect 1830 1592 1836 1593
rect 1830 1588 1831 1592
rect 1835 1588 1836 1592
rect 1830 1587 1836 1588
rect 142 1572 148 1573
rect 142 1568 143 1572
rect 147 1568 148 1572
rect 142 1567 148 1568
rect 182 1572 188 1573
rect 182 1568 183 1572
rect 187 1568 188 1572
rect 182 1567 188 1568
rect 230 1572 236 1573
rect 230 1568 231 1572
rect 235 1568 236 1572
rect 230 1567 236 1568
rect 286 1572 292 1573
rect 286 1568 287 1572
rect 291 1568 292 1572
rect 286 1567 292 1568
rect 350 1572 356 1573
rect 350 1568 351 1572
rect 355 1568 356 1572
rect 350 1567 356 1568
rect 414 1572 420 1573
rect 414 1568 415 1572
rect 419 1568 420 1572
rect 414 1567 420 1568
rect 478 1572 484 1573
rect 478 1568 479 1572
rect 483 1568 484 1572
rect 478 1567 484 1568
rect 542 1572 548 1573
rect 542 1568 543 1572
rect 547 1568 548 1572
rect 542 1567 548 1568
rect 606 1572 612 1573
rect 606 1568 607 1572
rect 611 1568 612 1572
rect 606 1567 612 1568
rect 662 1572 668 1573
rect 662 1568 663 1572
rect 667 1568 668 1572
rect 662 1567 668 1568
rect 726 1572 732 1573
rect 726 1568 727 1572
rect 731 1568 732 1572
rect 726 1567 732 1568
rect 790 1572 796 1573
rect 790 1568 791 1572
rect 795 1568 796 1572
rect 790 1567 796 1568
rect 854 1572 860 1573
rect 854 1568 855 1572
rect 859 1568 860 1572
rect 854 1567 860 1568
rect 110 1564 116 1565
rect 110 1560 111 1564
rect 115 1560 116 1564
rect 110 1559 116 1560
rect 1094 1564 1100 1565
rect 1094 1560 1095 1564
rect 1099 1560 1100 1564
rect 1094 1559 1100 1560
rect 1238 1556 1244 1557
rect 1238 1552 1239 1556
rect 1243 1552 1244 1556
rect 1238 1551 1244 1552
rect 1278 1556 1284 1557
rect 1278 1552 1279 1556
rect 1283 1552 1284 1556
rect 1278 1551 1284 1552
rect 1326 1556 1332 1557
rect 1326 1552 1327 1556
rect 1331 1552 1332 1556
rect 1326 1551 1332 1552
rect 1374 1556 1380 1557
rect 1374 1552 1375 1556
rect 1379 1552 1380 1556
rect 1374 1551 1380 1552
rect 1422 1556 1428 1557
rect 1422 1552 1423 1556
rect 1427 1552 1428 1556
rect 1422 1551 1428 1552
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1518 1556 1524 1557
rect 1518 1552 1519 1556
rect 1523 1552 1524 1556
rect 1518 1551 1524 1552
rect 1566 1556 1572 1557
rect 1566 1552 1567 1556
rect 1571 1552 1572 1556
rect 1566 1551 1572 1552
rect 1622 1556 1628 1557
rect 1622 1552 1623 1556
rect 1627 1552 1628 1556
rect 1622 1551 1628 1552
rect 1678 1556 1684 1557
rect 1678 1552 1679 1556
rect 1683 1552 1684 1556
rect 1678 1551 1684 1552
rect 1734 1556 1740 1557
rect 1734 1552 1735 1556
rect 1739 1552 1740 1556
rect 1734 1551 1740 1552
rect 1134 1548 1140 1549
rect 110 1547 116 1548
rect 110 1543 111 1547
rect 115 1543 116 1547
rect 1094 1547 1100 1548
rect 110 1542 116 1543
rect 142 1544 148 1545
rect 142 1540 143 1544
rect 147 1540 148 1544
rect 142 1539 148 1540
rect 182 1544 188 1545
rect 182 1540 183 1544
rect 187 1540 188 1544
rect 182 1539 188 1540
rect 230 1544 236 1545
rect 230 1540 231 1544
rect 235 1540 236 1544
rect 230 1539 236 1540
rect 286 1544 292 1545
rect 286 1540 287 1544
rect 291 1540 292 1544
rect 286 1539 292 1540
rect 350 1544 356 1545
rect 350 1540 351 1544
rect 355 1540 356 1544
rect 350 1539 356 1540
rect 414 1544 420 1545
rect 414 1540 415 1544
rect 419 1540 420 1544
rect 414 1539 420 1540
rect 478 1544 484 1545
rect 478 1540 479 1544
rect 483 1540 484 1544
rect 478 1539 484 1540
rect 542 1544 548 1545
rect 542 1540 543 1544
rect 547 1540 548 1544
rect 542 1539 548 1540
rect 606 1544 612 1545
rect 606 1540 607 1544
rect 611 1540 612 1544
rect 606 1539 612 1540
rect 662 1544 668 1545
rect 662 1540 663 1544
rect 667 1540 668 1544
rect 662 1539 668 1540
rect 726 1544 732 1545
rect 726 1540 727 1544
rect 731 1540 732 1544
rect 726 1539 732 1540
rect 790 1544 796 1545
rect 790 1540 791 1544
rect 795 1540 796 1544
rect 790 1539 796 1540
rect 854 1544 860 1545
rect 854 1540 855 1544
rect 859 1540 860 1544
rect 1094 1543 1095 1547
rect 1099 1543 1100 1547
rect 1134 1544 1135 1548
rect 1139 1544 1140 1548
rect 1134 1543 1140 1544
rect 2118 1548 2124 1549
rect 2118 1544 2119 1548
rect 2123 1544 2124 1548
rect 2118 1543 2124 1544
rect 1094 1542 1100 1543
rect 854 1539 860 1540
rect 1134 1531 1140 1532
rect 1134 1527 1135 1531
rect 1139 1527 1140 1531
rect 2118 1531 2124 1532
rect 1134 1526 1140 1527
rect 1238 1528 1244 1529
rect 134 1524 140 1525
rect 110 1521 116 1522
rect 110 1517 111 1521
rect 115 1517 116 1521
rect 134 1520 135 1524
rect 139 1520 140 1524
rect 134 1519 140 1520
rect 174 1524 180 1525
rect 174 1520 175 1524
rect 179 1520 180 1524
rect 174 1519 180 1520
rect 214 1524 220 1525
rect 214 1520 215 1524
rect 219 1520 220 1524
rect 214 1519 220 1520
rect 254 1524 260 1525
rect 254 1520 255 1524
rect 259 1520 260 1524
rect 254 1519 260 1520
rect 294 1524 300 1525
rect 294 1520 295 1524
rect 299 1520 300 1524
rect 294 1519 300 1520
rect 334 1524 340 1525
rect 334 1520 335 1524
rect 339 1520 340 1524
rect 334 1519 340 1520
rect 374 1524 380 1525
rect 374 1520 375 1524
rect 379 1520 380 1524
rect 374 1519 380 1520
rect 414 1524 420 1525
rect 414 1520 415 1524
rect 419 1520 420 1524
rect 414 1519 420 1520
rect 454 1524 460 1525
rect 454 1520 455 1524
rect 459 1520 460 1524
rect 454 1519 460 1520
rect 494 1524 500 1525
rect 494 1520 495 1524
rect 499 1520 500 1524
rect 494 1519 500 1520
rect 534 1524 540 1525
rect 534 1520 535 1524
rect 539 1520 540 1524
rect 534 1519 540 1520
rect 574 1524 580 1525
rect 574 1520 575 1524
rect 579 1520 580 1524
rect 574 1519 580 1520
rect 614 1524 620 1525
rect 614 1520 615 1524
rect 619 1520 620 1524
rect 614 1519 620 1520
rect 654 1524 660 1525
rect 654 1520 655 1524
rect 659 1520 660 1524
rect 654 1519 660 1520
rect 694 1524 700 1525
rect 694 1520 695 1524
rect 699 1520 700 1524
rect 694 1519 700 1520
rect 734 1524 740 1525
rect 734 1520 735 1524
rect 739 1520 740 1524
rect 734 1519 740 1520
rect 774 1524 780 1525
rect 774 1520 775 1524
rect 779 1520 780 1524
rect 774 1519 780 1520
rect 830 1524 836 1525
rect 830 1520 831 1524
rect 835 1520 836 1524
rect 830 1519 836 1520
rect 886 1524 892 1525
rect 886 1520 887 1524
rect 891 1520 892 1524
rect 1238 1524 1239 1528
rect 1243 1524 1244 1528
rect 1238 1523 1244 1524
rect 1278 1528 1284 1529
rect 1278 1524 1279 1528
rect 1283 1524 1284 1528
rect 1278 1523 1284 1524
rect 1326 1528 1332 1529
rect 1326 1524 1327 1528
rect 1331 1524 1332 1528
rect 1326 1523 1332 1524
rect 1374 1528 1380 1529
rect 1374 1524 1375 1528
rect 1379 1524 1380 1528
rect 1374 1523 1380 1524
rect 1422 1528 1428 1529
rect 1422 1524 1423 1528
rect 1427 1524 1428 1528
rect 1422 1523 1428 1524
rect 1470 1528 1476 1529
rect 1470 1524 1471 1528
rect 1475 1524 1476 1528
rect 1470 1523 1476 1524
rect 1518 1528 1524 1529
rect 1518 1524 1519 1528
rect 1523 1524 1524 1528
rect 1518 1523 1524 1524
rect 1566 1528 1572 1529
rect 1566 1524 1567 1528
rect 1571 1524 1572 1528
rect 1566 1523 1572 1524
rect 1622 1528 1628 1529
rect 1622 1524 1623 1528
rect 1627 1524 1628 1528
rect 1622 1523 1628 1524
rect 1678 1528 1684 1529
rect 1678 1524 1679 1528
rect 1683 1524 1684 1528
rect 1678 1523 1684 1524
rect 1734 1528 1740 1529
rect 1734 1524 1735 1528
rect 1739 1524 1740 1528
rect 2118 1527 2119 1531
rect 2123 1527 2124 1531
rect 2118 1526 2124 1527
rect 1734 1523 1740 1524
rect 886 1519 892 1520
rect 1094 1521 1100 1522
rect 110 1516 116 1517
rect 1094 1517 1095 1521
rect 1099 1517 1100 1521
rect 1094 1516 1100 1517
rect 1318 1512 1324 1513
rect 1134 1509 1140 1510
rect 1134 1505 1135 1509
rect 1139 1505 1140 1509
rect 1318 1508 1319 1512
rect 1323 1508 1324 1512
rect 1318 1507 1324 1508
rect 1358 1512 1364 1513
rect 1358 1508 1359 1512
rect 1363 1508 1364 1512
rect 1358 1507 1364 1508
rect 1398 1512 1404 1513
rect 1398 1508 1399 1512
rect 1403 1508 1404 1512
rect 1398 1507 1404 1508
rect 1438 1512 1444 1513
rect 1438 1508 1439 1512
rect 1443 1508 1444 1512
rect 1438 1507 1444 1508
rect 1478 1512 1484 1513
rect 1478 1508 1479 1512
rect 1483 1508 1484 1512
rect 1478 1507 1484 1508
rect 1518 1512 1524 1513
rect 1518 1508 1519 1512
rect 1523 1508 1524 1512
rect 1518 1507 1524 1508
rect 1558 1512 1564 1513
rect 1558 1508 1559 1512
rect 1563 1508 1564 1512
rect 1558 1507 1564 1508
rect 1606 1512 1612 1513
rect 1606 1508 1607 1512
rect 1611 1508 1612 1512
rect 1606 1507 1612 1508
rect 1662 1512 1668 1513
rect 1662 1508 1663 1512
rect 1667 1508 1668 1512
rect 1662 1507 1668 1508
rect 1734 1512 1740 1513
rect 1734 1508 1735 1512
rect 1739 1508 1740 1512
rect 1734 1507 1740 1508
rect 1814 1512 1820 1513
rect 1814 1508 1815 1512
rect 1819 1508 1820 1512
rect 1814 1507 1820 1508
rect 1902 1512 1908 1513
rect 1902 1508 1903 1512
rect 1907 1508 1908 1512
rect 1902 1507 1908 1508
rect 1990 1512 1996 1513
rect 1990 1508 1991 1512
rect 1995 1508 1996 1512
rect 1990 1507 1996 1508
rect 2070 1512 2076 1513
rect 2070 1508 2071 1512
rect 2075 1508 2076 1512
rect 2070 1507 2076 1508
rect 2118 1509 2124 1510
rect 110 1504 116 1505
rect 110 1500 111 1504
rect 115 1500 116 1504
rect 110 1499 116 1500
rect 1094 1504 1100 1505
rect 1134 1504 1140 1505
rect 2118 1505 2119 1509
rect 2123 1505 2124 1509
rect 2118 1504 2124 1505
rect 1094 1500 1095 1504
rect 1099 1500 1100 1504
rect 1094 1499 1100 1500
rect 134 1496 140 1497
rect 134 1492 135 1496
rect 139 1492 140 1496
rect 134 1491 140 1492
rect 174 1496 180 1497
rect 174 1492 175 1496
rect 179 1492 180 1496
rect 174 1491 180 1492
rect 214 1496 220 1497
rect 214 1492 215 1496
rect 219 1492 220 1496
rect 214 1491 220 1492
rect 254 1496 260 1497
rect 254 1492 255 1496
rect 259 1492 260 1496
rect 254 1491 260 1492
rect 294 1496 300 1497
rect 294 1492 295 1496
rect 299 1492 300 1496
rect 294 1491 300 1492
rect 334 1496 340 1497
rect 334 1492 335 1496
rect 339 1492 340 1496
rect 334 1491 340 1492
rect 374 1496 380 1497
rect 374 1492 375 1496
rect 379 1492 380 1496
rect 374 1491 380 1492
rect 414 1496 420 1497
rect 414 1492 415 1496
rect 419 1492 420 1496
rect 414 1491 420 1492
rect 454 1496 460 1497
rect 454 1492 455 1496
rect 459 1492 460 1496
rect 454 1491 460 1492
rect 494 1496 500 1497
rect 494 1492 495 1496
rect 499 1492 500 1496
rect 494 1491 500 1492
rect 534 1496 540 1497
rect 534 1492 535 1496
rect 539 1492 540 1496
rect 534 1491 540 1492
rect 574 1496 580 1497
rect 574 1492 575 1496
rect 579 1492 580 1496
rect 574 1491 580 1492
rect 614 1496 620 1497
rect 614 1492 615 1496
rect 619 1492 620 1496
rect 614 1491 620 1492
rect 654 1496 660 1497
rect 654 1492 655 1496
rect 659 1492 660 1496
rect 654 1491 660 1492
rect 694 1496 700 1497
rect 694 1492 695 1496
rect 699 1492 700 1496
rect 694 1491 700 1492
rect 734 1496 740 1497
rect 734 1492 735 1496
rect 739 1492 740 1496
rect 734 1491 740 1492
rect 774 1496 780 1497
rect 774 1492 775 1496
rect 779 1492 780 1496
rect 774 1491 780 1492
rect 830 1496 836 1497
rect 830 1492 831 1496
rect 835 1492 836 1496
rect 830 1491 836 1492
rect 886 1496 892 1497
rect 886 1492 887 1496
rect 891 1492 892 1496
rect 886 1491 892 1492
rect 1134 1492 1140 1493
rect 1134 1488 1135 1492
rect 1139 1488 1140 1492
rect 1134 1487 1140 1488
rect 2118 1492 2124 1493
rect 2118 1488 2119 1492
rect 2123 1488 2124 1492
rect 2118 1487 2124 1488
rect 1318 1484 1324 1485
rect 1318 1480 1319 1484
rect 1323 1480 1324 1484
rect 1318 1479 1324 1480
rect 1358 1484 1364 1485
rect 1358 1480 1359 1484
rect 1363 1480 1364 1484
rect 1358 1479 1364 1480
rect 1398 1484 1404 1485
rect 1398 1480 1399 1484
rect 1403 1480 1404 1484
rect 1398 1479 1404 1480
rect 1438 1484 1444 1485
rect 1438 1480 1439 1484
rect 1443 1480 1444 1484
rect 1438 1479 1444 1480
rect 1478 1484 1484 1485
rect 1478 1480 1479 1484
rect 1483 1480 1484 1484
rect 1478 1479 1484 1480
rect 1518 1484 1524 1485
rect 1518 1480 1519 1484
rect 1523 1480 1524 1484
rect 1518 1479 1524 1480
rect 1558 1484 1564 1485
rect 1558 1480 1559 1484
rect 1563 1480 1564 1484
rect 1558 1479 1564 1480
rect 1606 1484 1612 1485
rect 1606 1480 1607 1484
rect 1611 1480 1612 1484
rect 1606 1479 1612 1480
rect 1662 1484 1668 1485
rect 1662 1480 1663 1484
rect 1667 1480 1668 1484
rect 1662 1479 1668 1480
rect 1734 1484 1740 1485
rect 1734 1480 1735 1484
rect 1739 1480 1740 1484
rect 1734 1479 1740 1480
rect 1814 1484 1820 1485
rect 1814 1480 1815 1484
rect 1819 1480 1820 1484
rect 1814 1479 1820 1480
rect 1902 1484 1908 1485
rect 1902 1480 1903 1484
rect 1907 1480 1908 1484
rect 1902 1479 1908 1480
rect 1990 1484 1996 1485
rect 1990 1480 1991 1484
rect 1995 1480 1996 1484
rect 1990 1479 1996 1480
rect 2070 1484 2076 1485
rect 2070 1480 2071 1484
rect 2075 1480 2076 1484
rect 2070 1479 2076 1480
rect 518 1452 524 1453
rect 518 1448 519 1452
rect 523 1448 524 1452
rect 518 1447 524 1448
rect 558 1452 564 1453
rect 558 1448 559 1452
rect 563 1448 564 1452
rect 558 1447 564 1448
rect 598 1452 604 1453
rect 598 1448 599 1452
rect 603 1448 604 1452
rect 598 1447 604 1448
rect 646 1452 652 1453
rect 646 1448 647 1452
rect 651 1448 652 1452
rect 646 1447 652 1448
rect 694 1452 700 1453
rect 694 1448 695 1452
rect 699 1448 700 1452
rect 694 1447 700 1448
rect 750 1452 756 1453
rect 750 1448 751 1452
rect 755 1448 756 1452
rect 750 1447 756 1448
rect 806 1452 812 1453
rect 806 1448 807 1452
rect 811 1448 812 1452
rect 806 1447 812 1448
rect 870 1452 876 1453
rect 870 1448 871 1452
rect 875 1448 876 1452
rect 870 1447 876 1448
rect 934 1452 940 1453
rect 934 1448 935 1452
rect 939 1448 940 1452
rect 934 1447 940 1448
rect 1230 1448 1236 1449
rect 110 1444 116 1445
rect 110 1440 111 1444
rect 115 1440 116 1444
rect 110 1439 116 1440
rect 1094 1444 1100 1445
rect 1094 1440 1095 1444
rect 1099 1440 1100 1444
rect 1230 1444 1231 1448
rect 1235 1444 1236 1448
rect 1230 1443 1236 1444
rect 1278 1448 1284 1449
rect 1278 1444 1279 1448
rect 1283 1444 1284 1448
rect 1278 1443 1284 1444
rect 1334 1448 1340 1449
rect 1334 1444 1335 1448
rect 1339 1444 1340 1448
rect 1334 1443 1340 1444
rect 1390 1448 1396 1449
rect 1390 1444 1391 1448
rect 1395 1444 1396 1448
rect 1390 1443 1396 1444
rect 1454 1448 1460 1449
rect 1454 1444 1455 1448
rect 1459 1444 1460 1448
rect 1454 1443 1460 1444
rect 1518 1448 1524 1449
rect 1518 1444 1519 1448
rect 1523 1444 1524 1448
rect 1518 1443 1524 1444
rect 1582 1448 1588 1449
rect 1582 1444 1583 1448
rect 1587 1444 1588 1448
rect 1582 1443 1588 1444
rect 1646 1448 1652 1449
rect 1646 1444 1647 1448
rect 1651 1444 1652 1448
rect 1646 1443 1652 1444
rect 1718 1448 1724 1449
rect 1718 1444 1719 1448
rect 1723 1444 1724 1448
rect 1718 1443 1724 1444
rect 1806 1448 1812 1449
rect 1806 1444 1807 1448
rect 1811 1444 1812 1448
rect 1806 1443 1812 1444
rect 1894 1448 1900 1449
rect 1894 1444 1895 1448
rect 1899 1444 1900 1448
rect 1894 1443 1900 1444
rect 1990 1448 1996 1449
rect 1990 1444 1991 1448
rect 1995 1444 1996 1448
rect 1990 1443 1996 1444
rect 2070 1448 2076 1449
rect 2070 1444 2071 1448
rect 2075 1444 2076 1448
rect 2070 1443 2076 1444
rect 1094 1439 1100 1440
rect 1134 1440 1140 1441
rect 1134 1436 1135 1440
rect 1139 1436 1140 1440
rect 1134 1435 1140 1436
rect 2118 1440 2124 1441
rect 2118 1436 2119 1440
rect 2123 1436 2124 1440
rect 2118 1435 2124 1436
rect 110 1427 116 1428
rect 110 1423 111 1427
rect 115 1423 116 1427
rect 1094 1427 1100 1428
rect 110 1422 116 1423
rect 518 1424 524 1425
rect 518 1420 519 1424
rect 523 1420 524 1424
rect 518 1419 524 1420
rect 558 1424 564 1425
rect 558 1420 559 1424
rect 563 1420 564 1424
rect 558 1419 564 1420
rect 598 1424 604 1425
rect 598 1420 599 1424
rect 603 1420 604 1424
rect 598 1419 604 1420
rect 646 1424 652 1425
rect 646 1420 647 1424
rect 651 1420 652 1424
rect 646 1419 652 1420
rect 694 1424 700 1425
rect 694 1420 695 1424
rect 699 1420 700 1424
rect 694 1419 700 1420
rect 750 1424 756 1425
rect 750 1420 751 1424
rect 755 1420 756 1424
rect 750 1419 756 1420
rect 806 1424 812 1425
rect 806 1420 807 1424
rect 811 1420 812 1424
rect 806 1419 812 1420
rect 870 1424 876 1425
rect 870 1420 871 1424
rect 875 1420 876 1424
rect 870 1419 876 1420
rect 934 1424 940 1425
rect 934 1420 935 1424
rect 939 1420 940 1424
rect 1094 1423 1095 1427
rect 1099 1423 1100 1427
rect 1094 1422 1100 1423
rect 1134 1423 1140 1424
rect 934 1419 940 1420
rect 1134 1419 1135 1423
rect 1139 1419 1140 1423
rect 2118 1423 2124 1424
rect 1134 1418 1140 1419
rect 1230 1420 1236 1421
rect 1230 1416 1231 1420
rect 1235 1416 1236 1420
rect 1230 1415 1236 1416
rect 1278 1420 1284 1421
rect 1278 1416 1279 1420
rect 1283 1416 1284 1420
rect 1278 1415 1284 1416
rect 1334 1420 1340 1421
rect 1334 1416 1335 1420
rect 1339 1416 1340 1420
rect 1334 1415 1340 1416
rect 1390 1420 1396 1421
rect 1390 1416 1391 1420
rect 1395 1416 1396 1420
rect 1390 1415 1396 1416
rect 1454 1420 1460 1421
rect 1454 1416 1455 1420
rect 1459 1416 1460 1420
rect 1454 1415 1460 1416
rect 1518 1420 1524 1421
rect 1518 1416 1519 1420
rect 1523 1416 1524 1420
rect 1518 1415 1524 1416
rect 1582 1420 1588 1421
rect 1582 1416 1583 1420
rect 1587 1416 1588 1420
rect 1582 1415 1588 1416
rect 1646 1420 1652 1421
rect 1646 1416 1647 1420
rect 1651 1416 1652 1420
rect 1646 1415 1652 1416
rect 1718 1420 1724 1421
rect 1718 1416 1719 1420
rect 1723 1416 1724 1420
rect 1718 1415 1724 1416
rect 1806 1420 1812 1421
rect 1806 1416 1807 1420
rect 1811 1416 1812 1420
rect 1806 1415 1812 1416
rect 1894 1420 1900 1421
rect 1894 1416 1895 1420
rect 1899 1416 1900 1420
rect 1894 1415 1900 1416
rect 1990 1420 1996 1421
rect 1990 1416 1991 1420
rect 1995 1416 1996 1420
rect 1990 1415 1996 1416
rect 2070 1420 2076 1421
rect 2070 1416 2071 1420
rect 2075 1416 2076 1420
rect 2118 1419 2119 1423
rect 2123 1419 2124 1423
rect 2118 1418 2124 1419
rect 2070 1415 2076 1416
rect 430 1408 436 1409
rect 110 1405 116 1406
rect 110 1401 111 1405
rect 115 1401 116 1405
rect 430 1404 431 1408
rect 435 1404 436 1408
rect 430 1403 436 1404
rect 470 1408 476 1409
rect 470 1404 471 1408
rect 475 1404 476 1408
rect 470 1403 476 1404
rect 518 1408 524 1409
rect 518 1404 519 1408
rect 523 1404 524 1408
rect 518 1403 524 1404
rect 574 1408 580 1409
rect 574 1404 575 1408
rect 579 1404 580 1408
rect 574 1403 580 1404
rect 630 1408 636 1409
rect 630 1404 631 1408
rect 635 1404 636 1408
rect 630 1403 636 1404
rect 694 1408 700 1409
rect 694 1404 695 1408
rect 699 1404 700 1408
rect 694 1403 700 1404
rect 758 1408 764 1409
rect 758 1404 759 1408
rect 763 1404 764 1408
rect 758 1403 764 1404
rect 822 1408 828 1409
rect 822 1404 823 1408
rect 827 1404 828 1408
rect 822 1403 828 1404
rect 894 1408 900 1409
rect 894 1404 895 1408
rect 899 1404 900 1408
rect 894 1403 900 1404
rect 966 1408 972 1409
rect 966 1404 967 1408
rect 971 1404 972 1408
rect 966 1403 972 1404
rect 1094 1405 1100 1406
rect 110 1400 116 1401
rect 1094 1401 1095 1405
rect 1099 1401 1100 1405
rect 1158 1404 1164 1405
rect 1094 1400 1100 1401
rect 1134 1401 1140 1402
rect 1134 1397 1135 1401
rect 1139 1397 1140 1401
rect 1158 1400 1159 1404
rect 1163 1400 1164 1404
rect 1158 1399 1164 1400
rect 1198 1404 1204 1405
rect 1198 1400 1199 1404
rect 1203 1400 1204 1404
rect 1198 1399 1204 1400
rect 1262 1404 1268 1405
rect 1262 1400 1263 1404
rect 1267 1400 1268 1404
rect 1262 1399 1268 1400
rect 1350 1404 1356 1405
rect 1350 1400 1351 1404
rect 1355 1400 1356 1404
rect 1350 1399 1356 1400
rect 1446 1404 1452 1405
rect 1446 1400 1447 1404
rect 1451 1400 1452 1404
rect 1446 1399 1452 1400
rect 1542 1404 1548 1405
rect 1542 1400 1543 1404
rect 1547 1400 1548 1404
rect 1542 1399 1548 1400
rect 1630 1404 1636 1405
rect 1630 1400 1631 1404
rect 1635 1400 1636 1404
rect 1630 1399 1636 1400
rect 1718 1404 1724 1405
rect 1718 1400 1719 1404
rect 1723 1400 1724 1404
rect 1718 1399 1724 1400
rect 1798 1404 1804 1405
rect 1798 1400 1799 1404
rect 1803 1400 1804 1404
rect 1798 1399 1804 1400
rect 1870 1404 1876 1405
rect 1870 1400 1871 1404
rect 1875 1400 1876 1404
rect 1870 1399 1876 1400
rect 1942 1404 1948 1405
rect 1942 1400 1943 1404
rect 1947 1400 1948 1404
rect 1942 1399 1948 1400
rect 2014 1404 2020 1405
rect 2014 1400 2015 1404
rect 2019 1400 2020 1404
rect 2014 1399 2020 1400
rect 2070 1404 2076 1405
rect 2070 1400 2071 1404
rect 2075 1400 2076 1404
rect 2070 1399 2076 1400
rect 2118 1401 2124 1402
rect 1134 1396 1140 1397
rect 2118 1397 2119 1401
rect 2123 1397 2124 1401
rect 2118 1396 2124 1397
rect 110 1388 116 1389
rect 110 1384 111 1388
rect 115 1384 116 1388
rect 110 1383 116 1384
rect 1094 1388 1100 1389
rect 1094 1384 1095 1388
rect 1099 1384 1100 1388
rect 1094 1383 1100 1384
rect 1134 1384 1140 1385
rect 430 1380 436 1381
rect 430 1376 431 1380
rect 435 1376 436 1380
rect 430 1375 436 1376
rect 470 1380 476 1381
rect 470 1376 471 1380
rect 475 1376 476 1380
rect 470 1375 476 1376
rect 518 1380 524 1381
rect 518 1376 519 1380
rect 523 1376 524 1380
rect 518 1375 524 1376
rect 574 1380 580 1381
rect 574 1376 575 1380
rect 579 1376 580 1380
rect 574 1375 580 1376
rect 630 1380 636 1381
rect 630 1376 631 1380
rect 635 1376 636 1380
rect 630 1375 636 1376
rect 694 1380 700 1381
rect 694 1376 695 1380
rect 699 1376 700 1380
rect 694 1375 700 1376
rect 758 1380 764 1381
rect 758 1376 759 1380
rect 763 1376 764 1380
rect 758 1375 764 1376
rect 822 1380 828 1381
rect 822 1376 823 1380
rect 827 1376 828 1380
rect 822 1375 828 1376
rect 894 1380 900 1381
rect 894 1376 895 1380
rect 899 1376 900 1380
rect 894 1375 900 1376
rect 966 1380 972 1381
rect 966 1376 967 1380
rect 971 1376 972 1380
rect 1134 1380 1135 1384
rect 1139 1380 1140 1384
rect 1134 1379 1140 1380
rect 2118 1384 2124 1385
rect 2118 1380 2119 1384
rect 2123 1380 2124 1384
rect 2118 1379 2124 1380
rect 966 1375 972 1376
rect 1158 1376 1164 1377
rect 1158 1372 1159 1376
rect 1163 1372 1164 1376
rect 1158 1371 1164 1372
rect 1198 1376 1204 1377
rect 1198 1372 1199 1376
rect 1203 1372 1204 1376
rect 1198 1371 1204 1372
rect 1262 1376 1268 1377
rect 1262 1372 1263 1376
rect 1267 1372 1268 1376
rect 1262 1371 1268 1372
rect 1350 1376 1356 1377
rect 1350 1372 1351 1376
rect 1355 1372 1356 1376
rect 1350 1371 1356 1372
rect 1446 1376 1452 1377
rect 1446 1372 1447 1376
rect 1451 1372 1452 1376
rect 1446 1371 1452 1372
rect 1542 1376 1548 1377
rect 1542 1372 1543 1376
rect 1547 1372 1548 1376
rect 1542 1371 1548 1372
rect 1630 1376 1636 1377
rect 1630 1372 1631 1376
rect 1635 1372 1636 1376
rect 1630 1371 1636 1372
rect 1718 1376 1724 1377
rect 1718 1372 1719 1376
rect 1723 1372 1724 1376
rect 1718 1371 1724 1372
rect 1798 1376 1804 1377
rect 1798 1372 1799 1376
rect 1803 1372 1804 1376
rect 1798 1371 1804 1372
rect 1870 1376 1876 1377
rect 1870 1372 1871 1376
rect 1875 1372 1876 1376
rect 1870 1371 1876 1372
rect 1942 1376 1948 1377
rect 1942 1372 1943 1376
rect 1947 1372 1948 1376
rect 1942 1371 1948 1372
rect 2014 1376 2020 1377
rect 2014 1372 2015 1376
rect 2019 1372 2020 1376
rect 2014 1371 2020 1372
rect 2070 1376 2076 1377
rect 2070 1372 2071 1376
rect 2075 1372 2076 1376
rect 2070 1371 2076 1372
rect 374 1344 380 1345
rect 374 1340 375 1344
rect 379 1340 380 1344
rect 374 1339 380 1340
rect 422 1344 428 1345
rect 422 1340 423 1344
rect 427 1340 428 1344
rect 422 1339 428 1340
rect 478 1344 484 1345
rect 478 1340 479 1344
rect 483 1340 484 1344
rect 478 1339 484 1340
rect 542 1344 548 1345
rect 542 1340 543 1344
rect 547 1340 548 1344
rect 542 1339 548 1340
rect 606 1344 612 1345
rect 606 1340 607 1344
rect 611 1340 612 1344
rect 606 1339 612 1340
rect 670 1344 676 1345
rect 670 1340 671 1344
rect 675 1340 676 1344
rect 670 1339 676 1340
rect 734 1344 740 1345
rect 734 1340 735 1344
rect 739 1340 740 1344
rect 734 1339 740 1340
rect 798 1344 804 1345
rect 798 1340 799 1344
rect 803 1340 804 1344
rect 798 1339 804 1340
rect 862 1344 868 1345
rect 862 1340 863 1344
rect 867 1340 868 1344
rect 862 1339 868 1340
rect 926 1344 932 1345
rect 926 1340 927 1344
rect 931 1340 932 1344
rect 926 1339 932 1340
rect 998 1344 1004 1345
rect 998 1340 999 1344
rect 1003 1340 1004 1344
rect 998 1339 1004 1340
rect 1046 1344 1052 1345
rect 1046 1340 1047 1344
rect 1051 1340 1052 1344
rect 1046 1339 1052 1340
rect 110 1336 116 1337
rect 110 1332 111 1336
rect 115 1332 116 1336
rect 110 1331 116 1332
rect 1094 1336 1100 1337
rect 1094 1332 1095 1336
rect 1099 1332 1100 1336
rect 1094 1331 1100 1332
rect 1158 1336 1164 1337
rect 1158 1332 1159 1336
rect 1163 1332 1164 1336
rect 1158 1331 1164 1332
rect 1254 1336 1260 1337
rect 1254 1332 1255 1336
rect 1259 1332 1260 1336
rect 1254 1331 1260 1332
rect 1374 1336 1380 1337
rect 1374 1332 1375 1336
rect 1379 1332 1380 1336
rect 1374 1331 1380 1332
rect 1486 1336 1492 1337
rect 1486 1332 1487 1336
rect 1491 1332 1492 1336
rect 1486 1331 1492 1332
rect 1590 1336 1596 1337
rect 1590 1332 1591 1336
rect 1595 1332 1596 1336
rect 1590 1331 1596 1332
rect 1678 1336 1684 1337
rect 1678 1332 1679 1336
rect 1683 1332 1684 1336
rect 1678 1331 1684 1332
rect 1758 1336 1764 1337
rect 1758 1332 1759 1336
rect 1763 1332 1764 1336
rect 1758 1331 1764 1332
rect 1830 1336 1836 1337
rect 1830 1332 1831 1336
rect 1835 1332 1836 1336
rect 1830 1331 1836 1332
rect 1902 1336 1908 1337
rect 1902 1332 1903 1336
rect 1907 1332 1908 1336
rect 1902 1331 1908 1332
rect 1966 1336 1972 1337
rect 1966 1332 1967 1336
rect 1971 1332 1972 1336
rect 1966 1331 1972 1332
rect 2030 1336 2036 1337
rect 2030 1332 2031 1336
rect 2035 1332 2036 1336
rect 2030 1331 2036 1332
rect 2070 1336 2076 1337
rect 2070 1332 2071 1336
rect 2075 1332 2076 1336
rect 2070 1331 2076 1332
rect 1134 1328 1140 1329
rect 1134 1324 1135 1328
rect 1139 1324 1140 1328
rect 1134 1323 1140 1324
rect 2118 1328 2124 1329
rect 2118 1324 2119 1328
rect 2123 1324 2124 1328
rect 2118 1323 2124 1324
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 1094 1319 1100 1320
rect 110 1314 116 1315
rect 374 1316 380 1317
rect 374 1312 375 1316
rect 379 1312 380 1316
rect 374 1311 380 1312
rect 422 1316 428 1317
rect 422 1312 423 1316
rect 427 1312 428 1316
rect 422 1311 428 1312
rect 478 1316 484 1317
rect 478 1312 479 1316
rect 483 1312 484 1316
rect 478 1311 484 1312
rect 542 1316 548 1317
rect 542 1312 543 1316
rect 547 1312 548 1316
rect 542 1311 548 1312
rect 606 1316 612 1317
rect 606 1312 607 1316
rect 611 1312 612 1316
rect 606 1311 612 1312
rect 670 1316 676 1317
rect 670 1312 671 1316
rect 675 1312 676 1316
rect 670 1311 676 1312
rect 734 1316 740 1317
rect 734 1312 735 1316
rect 739 1312 740 1316
rect 734 1311 740 1312
rect 798 1316 804 1317
rect 798 1312 799 1316
rect 803 1312 804 1316
rect 798 1311 804 1312
rect 862 1316 868 1317
rect 862 1312 863 1316
rect 867 1312 868 1316
rect 862 1311 868 1312
rect 926 1316 932 1317
rect 926 1312 927 1316
rect 931 1312 932 1316
rect 926 1311 932 1312
rect 998 1316 1004 1317
rect 998 1312 999 1316
rect 1003 1312 1004 1316
rect 998 1311 1004 1312
rect 1046 1316 1052 1317
rect 1046 1312 1047 1316
rect 1051 1312 1052 1316
rect 1094 1315 1095 1319
rect 1099 1315 1100 1319
rect 1094 1314 1100 1315
rect 1046 1311 1052 1312
rect 1134 1311 1140 1312
rect 1134 1307 1135 1311
rect 1139 1307 1140 1311
rect 2118 1311 2124 1312
rect 1134 1306 1140 1307
rect 1158 1308 1164 1309
rect 334 1304 340 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 334 1300 335 1304
rect 339 1300 340 1304
rect 334 1299 340 1300
rect 390 1304 396 1305
rect 390 1300 391 1304
rect 395 1300 396 1304
rect 390 1299 396 1300
rect 454 1304 460 1305
rect 454 1300 455 1304
rect 459 1300 460 1304
rect 454 1299 460 1300
rect 526 1304 532 1305
rect 526 1300 527 1304
rect 531 1300 532 1304
rect 526 1299 532 1300
rect 598 1304 604 1305
rect 598 1300 599 1304
rect 603 1300 604 1304
rect 598 1299 604 1300
rect 670 1304 676 1305
rect 670 1300 671 1304
rect 675 1300 676 1304
rect 670 1299 676 1300
rect 742 1304 748 1305
rect 742 1300 743 1304
rect 747 1300 748 1304
rect 742 1299 748 1300
rect 822 1304 828 1305
rect 822 1300 823 1304
rect 827 1300 828 1304
rect 822 1299 828 1300
rect 902 1304 908 1305
rect 902 1300 903 1304
rect 907 1300 908 1304
rect 902 1299 908 1300
rect 982 1304 988 1305
rect 982 1300 983 1304
rect 987 1300 988 1304
rect 982 1299 988 1300
rect 1046 1304 1052 1305
rect 1046 1300 1047 1304
rect 1051 1300 1052 1304
rect 1158 1304 1159 1308
rect 1163 1304 1164 1308
rect 1158 1303 1164 1304
rect 1254 1308 1260 1309
rect 1254 1304 1255 1308
rect 1259 1304 1260 1308
rect 1254 1303 1260 1304
rect 1374 1308 1380 1309
rect 1374 1304 1375 1308
rect 1379 1304 1380 1308
rect 1374 1303 1380 1304
rect 1486 1308 1492 1309
rect 1486 1304 1487 1308
rect 1491 1304 1492 1308
rect 1486 1303 1492 1304
rect 1590 1308 1596 1309
rect 1590 1304 1591 1308
rect 1595 1304 1596 1308
rect 1590 1303 1596 1304
rect 1678 1308 1684 1309
rect 1678 1304 1679 1308
rect 1683 1304 1684 1308
rect 1678 1303 1684 1304
rect 1758 1308 1764 1309
rect 1758 1304 1759 1308
rect 1763 1304 1764 1308
rect 1758 1303 1764 1304
rect 1830 1308 1836 1309
rect 1830 1304 1831 1308
rect 1835 1304 1836 1308
rect 1830 1303 1836 1304
rect 1902 1308 1908 1309
rect 1902 1304 1903 1308
rect 1907 1304 1908 1308
rect 1902 1303 1908 1304
rect 1966 1308 1972 1309
rect 1966 1304 1967 1308
rect 1971 1304 1972 1308
rect 1966 1303 1972 1304
rect 2030 1308 2036 1309
rect 2030 1304 2031 1308
rect 2035 1304 2036 1308
rect 2030 1303 2036 1304
rect 2070 1308 2076 1309
rect 2070 1304 2071 1308
rect 2075 1304 2076 1308
rect 2118 1307 2119 1311
rect 2123 1307 2124 1311
rect 2118 1306 2124 1307
rect 2070 1303 2076 1304
rect 1046 1299 1052 1300
rect 1094 1301 1100 1302
rect 110 1296 116 1297
rect 1094 1297 1095 1301
rect 1099 1297 1100 1301
rect 1094 1296 1100 1297
rect 1158 1292 1164 1293
rect 1134 1289 1140 1290
rect 1134 1285 1135 1289
rect 1139 1285 1140 1289
rect 1158 1288 1159 1292
rect 1163 1288 1164 1292
rect 1158 1287 1164 1288
rect 1198 1292 1204 1293
rect 1198 1288 1199 1292
rect 1203 1288 1204 1292
rect 1198 1287 1204 1288
rect 1246 1292 1252 1293
rect 1246 1288 1247 1292
rect 1251 1288 1252 1292
rect 1246 1287 1252 1288
rect 1318 1292 1324 1293
rect 1318 1288 1319 1292
rect 1323 1288 1324 1292
rect 1318 1287 1324 1288
rect 1398 1292 1404 1293
rect 1398 1288 1399 1292
rect 1403 1288 1404 1292
rect 1398 1287 1404 1288
rect 1478 1292 1484 1293
rect 1478 1288 1479 1292
rect 1483 1288 1484 1292
rect 1478 1287 1484 1288
rect 1558 1292 1564 1293
rect 1558 1288 1559 1292
rect 1563 1288 1564 1292
rect 1558 1287 1564 1288
rect 1638 1292 1644 1293
rect 1638 1288 1639 1292
rect 1643 1288 1644 1292
rect 1638 1287 1644 1288
rect 1718 1292 1724 1293
rect 1718 1288 1719 1292
rect 1723 1288 1724 1292
rect 1718 1287 1724 1288
rect 1798 1292 1804 1293
rect 1798 1288 1799 1292
rect 1803 1288 1804 1292
rect 1798 1287 1804 1288
rect 1878 1292 1884 1293
rect 1878 1288 1879 1292
rect 1883 1288 1884 1292
rect 1878 1287 1884 1288
rect 1966 1292 1972 1293
rect 1966 1288 1967 1292
rect 1971 1288 1972 1292
rect 1966 1287 1972 1288
rect 2054 1292 2060 1293
rect 2054 1288 2055 1292
rect 2059 1288 2060 1292
rect 2054 1287 2060 1288
rect 2118 1289 2124 1290
rect 110 1284 116 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 110 1279 116 1280
rect 1094 1284 1100 1285
rect 1134 1284 1140 1285
rect 2118 1285 2119 1289
rect 2123 1285 2124 1289
rect 2118 1284 2124 1285
rect 1094 1280 1095 1284
rect 1099 1280 1100 1284
rect 1094 1279 1100 1280
rect 334 1276 340 1277
rect 334 1272 335 1276
rect 339 1272 340 1276
rect 334 1271 340 1272
rect 390 1276 396 1277
rect 390 1272 391 1276
rect 395 1272 396 1276
rect 390 1271 396 1272
rect 454 1276 460 1277
rect 454 1272 455 1276
rect 459 1272 460 1276
rect 454 1271 460 1272
rect 526 1276 532 1277
rect 526 1272 527 1276
rect 531 1272 532 1276
rect 526 1271 532 1272
rect 598 1276 604 1277
rect 598 1272 599 1276
rect 603 1272 604 1276
rect 598 1271 604 1272
rect 670 1276 676 1277
rect 670 1272 671 1276
rect 675 1272 676 1276
rect 670 1271 676 1272
rect 742 1276 748 1277
rect 742 1272 743 1276
rect 747 1272 748 1276
rect 742 1271 748 1272
rect 822 1276 828 1277
rect 822 1272 823 1276
rect 827 1272 828 1276
rect 822 1271 828 1272
rect 902 1276 908 1277
rect 902 1272 903 1276
rect 907 1272 908 1276
rect 902 1271 908 1272
rect 982 1276 988 1277
rect 982 1272 983 1276
rect 987 1272 988 1276
rect 982 1271 988 1272
rect 1046 1276 1052 1277
rect 1046 1272 1047 1276
rect 1051 1272 1052 1276
rect 1046 1271 1052 1272
rect 1134 1272 1140 1273
rect 1134 1268 1135 1272
rect 1139 1268 1140 1272
rect 1134 1267 1140 1268
rect 2118 1272 2124 1273
rect 2118 1268 2119 1272
rect 2123 1268 2124 1272
rect 2118 1267 2124 1268
rect 1158 1264 1164 1265
rect 1158 1260 1159 1264
rect 1163 1260 1164 1264
rect 1158 1259 1164 1260
rect 1198 1264 1204 1265
rect 1198 1260 1199 1264
rect 1203 1260 1204 1264
rect 1198 1259 1204 1260
rect 1246 1264 1252 1265
rect 1246 1260 1247 1264
rect 1251 1260 1252 1264
rect 1246 1259 1252 1260
rect 1318 1264 1324 1265
rect 1318 1260 1319 1264
rect 1323 1260 1324 1264
rect 1318 1259 1324 1260
rect 1398 1264 1404 1265
rect 1398 1260 1399 1264
rect 1403 1260 1404 1264
rect 1398 1259 1404 1260
rect 1478 1264 1484 1265
rect 1478 1260 1479 1264
rect 1483 1260 1484 1264
rect 1478 1259 1484 1260
rect 1558 1264 1564 1265
rect 1558 1260 1559 1264
rect 1563 1260 1564 1264
rect 1558 1259 1564 1260
rect 1638 1264 1644 1265
rect 1638 1260 1639 1264
rect 1643 1260 1644 1264
rect 1638 1259 1644 1260
rect 1718 1264 1724 1265
rect 1718 1260 1719 1264
rect 1723 1260 1724 1264
rect 1718 1259 1724 1260
rect 1798 1264 1804 1265
rect 1798 1260 1799 1264
rect 1803 1260 1804 1264
rect 1798 1259 1804 1260
rect 1878 1264 1884 1265
rect 1878 1260 1879 1264
rect 1883 1260 1884 1264
rect 1878 1259 1884 1260
rect 1966 1264 1972 1265
rect 1966 1260 1967 1264
rect 1971 1260 1972 1264
rect 1966 1259 1972 1260
rect 2054 1264 2060 1265
rect 2054 1260 2055 1264
rect 2059 1260 2060 1264
rect 2054 1259 2060 1260
rect 262 1236 268 1237
rect 262 1232 263 1236
rect 267 1232 268 1236
rect 262 1231 268 1232
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 358 1236 364 1237
rect 358 1232 359 1236
rect 363 1232 364 1236
rect 358 1231 364 1232
rect 414 1236 420 1237
rect 414 1232 415 1236
rect 419 1232 420 1236
rect 414 1231 420 1232
rect 478 1236 484 1237
rect 478 1232 479 1236
rect 483 1232 484 1236
rect 478 1231 484 1232
rect 542 1236 548 1237
rect 542 1232 543 1236
rect 547 1232 548 1236
rect 542 1231 548 1232
rect 606 1236 612 1237
rect 606 1232 607 1236
rect 611 1232 612 1236
rect 606 1231 612 1232
rect 670 1236 676 1237
rect 670 1232 671 1236
rect 675 1232 676 1236
rect 670 1231 676 1232
rect 734 1236 740 1237
rect 734 1232 735 1236
rect 739 1232 740 1236
rect 734 1231 740 1232
rect 798 1236 804 1237
rect 798 1232 799 1236
rect 803 1232 804 1236
rect 798 1231 804 1232
rect 862 1236 868 1237
rect 862 1232 863 1236
rect 867 1232 868 1236
rect 862 1231 868 1232
rect 926 1236 932 1237
rect 926 1232 927 1236
rect 931 1232 932 1236
rect 926 1231 932 1232
rect 110 1228 116 1229
rect 110 1224 111 1228
rect 115 1224 116 1228
rect 110 1223 116 1224
rect 1094 1228 1100 1229
rect 1094 1224 1095 1228
rect 1099 1224 1100 1228
rect 1094 1223 1100 1224
rect 1158 1224 1164 1225
rect 1158 1220 1159 1224
rect 1163 1220 1164 1224
rect 1158 1219 1164 1220
rect 1198 1224 1204 1225
rect 1198 1220 1199 1224
rect 1203 1220 1204 1224
rect 1198 1219 1204 1220
rect 1238 1224 1244 1225
rect 1238 1220 1239 1224
rect 1243 1220 1244 1224
rect 1238 1219 1244 1220
rect 1278 1224 1284 1225
rect 1278 1220 1279 1224
rect 1283 1220 1284 1224
rect 1278 1219 1284 1220
rect 1326 1224 1332 1225
rect 1326 1220 1327 1224
rect 1331 1220 1332 1224
rect 1326 1219 1332 1220
rect 1374 1224 1380 1225
rect 1374 1220 1375 1224
rect 1379 1220 1380 1224
rect 1374 1219 1380 1220
rect 1422 1224 1428 1225
rect 1422 1220 1423 1224
rect 1427 1220 1428 1224
rect 1422 1219 1428 1220
rect 1470 1224 1476 1225
rect 1470 1220 1471 1224
rect 1475 1220 1476 1224
rect 1470 1219 1476 1220
rect 1534 1224 1540 1225
rect 1534 1220 1535 1224
rect 1539 1220 1540 1224
rect 1534 1219 1540 1220
rect 1614 1224 1620 1225
rect 1614 1220 1615 1224
rect 1619 1220 1620 1224
rect 1614 1219 1620 1220
rect 1718 1224 1724 1225
rect 1718 1220 1719 1224
rect 1723 1220 1724 1224
rect 1718 1219 1724 1220
rect 1838 1224 1844 1225
rect 1838 1220 1839 1224
rect 1843 1220 1844 1224
rect 1838 1219 1844 1220
rect 1966 1224 1972 1225
rect 1966 1220 1967 1224
rect 1971 1220 1972 1224
rect 1966 1219 1972 1220
rect 2070 1224 2076 1225
rect 2070 1220 2071 1224
rect 2075 1220 2076 1224
rect 2070 1219 2076 1220
rect 1134 1216 1140 1217
rect 1134 1212 1135 1216
rect 1139 1212 1140 1216
rect 110 1211 116 1212
rect 110 1207 111 1211
rect 115 1207 116 1211
rect 1094 1211 1100 1212
rect 1134 1211 1140 1212
rect 2118 1216 2124 1217
rect 2118 1212 2119 1216
rect 2123 1212 2124 1216
rect 2118 1211 2124 1212
rect 110 1206 116 1207
rect 262 1208 268 1209
rect 262 1204 263 1208
rect 267 1204 268 1208
rect 262 1203 268 1204
rect 310 1208 316 1209
rect 310 1204 311 1208
rect 315 1204 316 1208
rect 310 1203 316 1204
rect 358 1208 364 1209
rect 358 1204 359 1208
rect 363 1204 364 1208
rect 358 1203 364 1204
rect 414 1208 420 1209
rect 414 1204 415 1208
rect 419 1204 420 1208
rect 414 1203 420 1204
rect 478 1208 484 1209
rect 478 1204 479 1208
rect 483 1204 484 1208
rect 478 1203 484 1204
rect 542 1208 548 1209
rect 542 1204 543 1208
rect 547 1204 548 1208
rect 542 1203 548 1204
rect 606 1208 612 1209
rect 606 1204 607 1208
rect 611 1204 612 1208
rect 606 1203 612 1204
rect 670 1208 676 1209
rect 670 1204 671 1208
rect 675 1204 676 1208
rect 670 1203 676 1204
rect 734 1208 740 1209
rect 734 1204 735 1208
rect 739 1204 740 1208
rect 734 1203 740 1204
rect 798 1208 804 1209
rect 798 1204 799 1208
rect 803 1204 804 1208
rect 798 1203 804 1204
rect 862 1208 868 1209
rect 862 1204 863 1208
rect 867 1204 868 1208
rect 862 1203 868 1204
rect 926 1208 932 1209
rect 926 1204 927 1208
rect 931 1204 932 1208
rect 1094 1207 1095 1211
rect 1099 1207 1100 1211
rect 1094 1206 1100 1207
rect 926 1203 932 1204
rect 1134 1199 1140 1200
rect 222 1196 228 1197
rect 110 1193 116 1194
rect 110 1189 111 1193
rect 115 1189 116 1193
rect 222 1192 223 1196
rect 227 1192 228 1196
rect 222 1191 228 1192
rect 278 1196 284 1197
rect 278 1192 279 1196
rect 283 1192 284 1196
rect 278 1191 284 1192
rect 342 1196 348 1197
rect 342 1192 343 1196
rect 347 1192 348 1196
rect 342 1191 348 1192
rect 406 1196 412 1197
rect 406 1192 407 1196
rect 411 1192 412 1196
rect 406 1191 412 1192
rect 478 1196 484 1197
rect 478 1192 479 1196
rect 483 1192 484 1196
rect 478 1191 484 1192
rect 550 1196 556 1197
rect 550 1192 551 1196
rect 555 1192 556 1196
rect 550 1191 556 1192
rect 630 1196 636 1197
rect 630 1192 631 1196
rect 635 1192 636 1196
rect 630 1191 636 1192
rect 710 1196 716 1197
rect 710 1192 711 1196
rect 715 1192 716 1196
rect 710 1191 716 1192
rect 790 1196 796 1197
rect 790 1192 791 1196
rect 795 1192 796 1196
rect 790 1191 796 1192
rect 870 1196 876 1197
rect 870 1192 871 1196
rect 875 1192 876 1196
rect 870 1191 876 1192
rect 958 1196 964 1197
rect 958 1192 959 1196
rect 963 1192 964 1196
rect 1134 1195 1135 1199
rect 1139 1195 1140 1199
rect 2118 1199 2124 1200
rect 1134 1194 1140 1195
rect 1158 1196 1164 1197
rect 958 1191 964 1192
rect 1094 1193 1100 1194
rect 110 1188 116 1189
rect 1094 1189 1095 1193
rect 1099 1189 1100 1193
rect 1158 1192 1159 1196
rect 1163 1192 1164 1196
rect 1158 1191 1164 1192
rect 1198 1196 1204 1197
rect 1198 1192 1199 1196
rect 1203 1192 1204 1196
rect 1198 1191 1204 1192
rect 1238 1196 1244 1197
rect 1238 1192 1239 1196
rect 1243 1192 1244 1196
rect 1238 1191 1244 1192
rect 1278 1196 1284 1197
rect 1278 1192 1279 1196
rect 1283 1192 1284 1196
rect 1278 1191 1284 1192
rect 1326 1196 1332 1197
rect 1326 1192 1327 1196
rect 1331 1192 1332 1196
rect 1326 1191 1332 1192
rect 1374 1196 1380 1197
rect 1374 1192 1375 1196
rect 1379 1192 1380 1196
rect 1374 1191 1380 1192
rect 1422 1196 1428 1197
rect 1422 1192 1423 1196
rect 1427 1192 1428 1196
rect 1422 1191 1428 1192
rect 1470 1196 1476 1197
rect 1470 1192 1471 1196
rect 1475 1192 1476 1196
rect 1470 1191 1476 1192
rect 1534 1196 1540 1197
rect 1534 1192 1535 1196
rect 1539 1192 1540 1196
rect 1534 1191 1540 1192
rect 1614 1196 1620 1197
rect 1614 1192 1615 1196
rect 1619 1192 1620 1196
rect 1614 1191 1620 1192
rect 1718 1196 1724 1197
rect 1718 1192 1719 1196
rect 1723 1192 1724 1196
rect 1718 1191 1724 1192
rect 1838 1196 1844 1197
rect 1838 1192 1839 1196
rect 1843 1192 1844 1196
rect 1838 1191 1844 1192
rect 1966 1196 1972 1197
rect 1966 1192 1967 1196
rect 1971 1192 1972 1196
rect 1966 1191 1972 1192
rect 2070 1196 2076 1197
rect 2070 1192 2071 1196
rect 2075 1192 2076 1196
rect 2118 1195 2119 1199
rect 2123 1195 2124 1199
rect 2118 1194 2124 1195
rect 2070 1191 2076 1192
rect 1094 1188 1100 1189
rect 1286 1184 1292 1185
rect 1134 1181 1140 1182
rect 1134 1177 1135 1181
rect 1139 1177 1140 1181
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1286 1179 1292 1180
rect 1326 1184 1332 1185
rect 1326 1180 1327 1184
rect 1331 1180 1332 1184
rect 1326 1179 1332 1180
rect 1366 1184 1372 1185
rect 1366 1180 1367 1184
rect 1371 1180 1372 1184
rect 1366 1179 1372 1180
rect 1414 1184 1420 1185
rect 1414 1180 1415 1184
rect 1419 1180 1420 1184
rect 1414 1179 1420 1180
rect 1470 1184 1476 1185
rect 1470 1180 1471 1184
rect 1475 1180 1476 1184
rect 1470 1179 1476 1180
rect 1526 1184 1532 1185
rect 1526 1180 1527 1184
rect 1531 1180 1532 1184
rect 1526 1179 1532 1180
rect 1582 1184 1588 1185
rect 1582 1180 1583 1184
rect 1587 1180 1588 1184
rect 1582 1179 1588 1180
rect 1638 1184 1644 1185
rect 1638 1180 1639 1184
rect 1643 1180 1644 1184
rect 1638 1179 1644 1180
rect 1702 1184 1708 1185
rect 1702 1180 1703 1184
rect 1707 1180 1708 1184
rect 1702 1179 1708 1180
rect 1766 1184 1772 1185
rect 1766 1180 1767 1184
rect 1771 1180 1772 1184
rect 1766 1179 1772 1180
rect 1838 1184 1844 1185
rect 1838 1180 1839 1184
rect 1843 1180 1844 1184
rect 1838 1179 1844 1180
rect 1918 1184 1924 1185
rect 1918 1180 1919 1184
rect 1923 1180 1924 1184
rect 1918 1179 1924 1180
rect 2006 1184 2012 1185
rect 2006 1180 2007 1184
rect 2011 1180 2012 1184
rect 2006 1179 2012 1180
rect 2070 1184 2076 1185
rect 2070 1180 2071 1184
rect 2075 1180 2076 1184
rect 2070 1179 2076 1180
rect 2118 1181 2124 1182
rect 110 1176 116 1177
rect 110 1172 111 1176
rect 115 1172 116 1176
rect 110 1171 116 1172
rect 1094 1176 1100 1177
rect 1134 1176 1140 1177
rect 2118 1177 2119 1181
rect 2123 1177 2124 1181
rect 2118 1176 2124 1177
rect 1094 1172 1095 1176
rect 1099 1172 1100 1176
rect 1094 1171 1100 1172
rect 222 1168 228 1169
rect 222 1164 223 1168
rect 227 1164 228 1168
rect 222 1163 228 1164
rect 278 1168 284 1169
rect 278 1164 279 1168
rect 283 1164 284 1168
rect 278 1163 284 1164
rect 342 1168 348 1169
rect 342 1164 343 1168
rect 347 1164 348 1168
rect 342 1163 348 1164
rect 406 1168 412 1169
rect 406 1164 407 1168
rect 411 1164 412 1168
rect 406 1163 412 1164
rect 478 1168 484 1169
rect 478 1164 479 1168
rect 483 1164 484 1168
rect 478 1163 484 1164
rect 550 1168 556 1169
rect 550 1164 551 1168
rect 555 1164 556 1168
rect 550 1163 556 1164
rect 630 1168 636 1169
rect 630 1164 631 1168
rect 635 1164 636 1168
rect 630 1163 636 1164
rect 710 1168 716 1169
rect 710 1164 711 1168
rect 715 1164 716 1168
rect 710 1163 716 1164
rect 790 1168 796 1169
rect 790 1164 791 1168
rect 795 1164 796 1168
rect 790 1163 796 1164
rect 870 1168 876 1169
rect 870 1164 871 1168
rect 875 1164 876 1168
rect 870 1163 876 1164
rect 958 1168 964 1169
rect 958 1164 959 1168
rect 963 1164 964 1168
rect 958 1163 964 1164
rect 1134 1164 1140 1165
rect 1134 1160 1135 1164
rect 1139 1160 1140 1164
rect 1134 1159 1140 1160
rect 2118 1164 2124 1165
rect 2118 1160 2119 1164
rect 2123 1160 2124 1164
rect 2118 1159 2124 1160
rect 1286 1156 1292 1157
rect 1286 1152 1287 1156
rect 1291 1152 1292 1156
rect 1286 1151 1292 1152
rect 1326 1156 1332 1157
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1326 1151 1332 1152
rect 1366 1156 1372 1157
rect 1366 1152 1367 1156
rect 1371 1152 1372 1156
rect 1366 1151 1372 1152
rect 1414 1156 1420 1157
rect 1414 1152 1415 1156
rect 1419 1152 1420 1156
rect 1414 1151 1420 1152
rect 1470 1156 1476 1157
rect 1470 1152 1471 1156
rect 1475 1152 1476 1156
rect 1470 1151 1476 1152
rect 1526 1156 1532 1157
rect 1526 1152 1527 1156
rect 1531 1152 1532 1156
rect 1526 1151 1532 1152
rect 1582 1156 1588 1157
rect 1582 1152 1583 1156
rect 1587 1152 1588 1156
rect 1582 1151 1588 1152
rect 1638 1156 1644 1157
rect 1638 1152 1639 1156
rect 1643 1152 1644 1156
rect 1638 1151 1644 1152
rect 1702 1156 1708 1157
rect 1702 1152 1703 1156
rect 1707 1152 1708 1156
rect 1702 1151 1708 1152
rect 1766 1156 1772 1157
rect 1766 1152 1767 1156
rect 1771 1152 1772 1156
rect 1766 1151 1772 1152
rect 1838 1156 1844 1157
rect 1838 1152 1839 1156
rect 1843 1152 1844 1156
rect 1838 1151 1844 1152
rect 1918 1156 1924 1157
rect 1918 1152 1919 1156
rect 1923 1152 1924 1156
rect 1918 1151 1924 1152
rect 2006 1156 2012 1157
rect 2006 1152 2007 1156
rect 2011 1152 2012 1156
rect 2006 1151 2012 1152
rect 2070 1156 2076 1157
rect 2070 1152 2071 1156
rect 2075 1152 2076 1156
rect 2070 1151 2076 1152
rect 158 1132 164 1133
rect 158 1128 159 1132
rect 163 1128 164 1132
rect 158 1127 164 1128
rect 198 1132 204 1133
rect 198 1128 199 1132
rect 203 1128 204 1132
rect 198 1127 204 1128
rect 246 1132 252 1133
rect 246 1128 247 1132
rect 251 1128 252 1132
rect 246 1127 252 1128
rect 302 1132 308 1133
rect 302 1128 303 1132
rect 307 1128 308 1132
rect 302 1127 308 1128
rect 366 1132 372 1133
rect 366 1128 367 1132
rect 371 1128 372 1132
rect 366 1127 372 1128
rect 438 1132 444 1133
rect 438 1128 439 1132
rect 443 1128 444 1132
rect 438 1127 444 1128
rect 510 1132 516 1133
rect 510 1128 511 1132
rect 515 1128 516 1132
rect 510 1127 516 1128
rect 590 1132 596 1133
rect 590 1128 591 1132
rect 595 1128 596 1132
rect 590 1127 596 1128
rect 678 1132 684 1133
rect 678 1128 679 1132
rect 683 1128 684 1132
rect 678 1127 684 1128
rect 774 1132 780 1133
rect 774 1128 775 1132
rect 779 1128 780 1132
rect 774 1127 780 1128
rect 878 1132 884 1133
rect 878 1128 879 1132
rect 883 1128 884 1132
rect 878 1127 884 1128
rect 990 1132 996 1133
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 110 1124 116 1125
rect 110 1120 111 1124
rect 115 1120 116 1124
rect 110 1119 116 1120
rect 1094 1124 1100 1125
rect 1094 1120 1095 1124
rect 1099 1120 1100 1124
rect 1094 1119 1100 1120
rect 1382 1112 1388 1113
rect 1382 1108 1383 1112
rect 1387 1108 1388 1112
rect 110 1107 116 1108
rect 110 1103 111 1107
rect 115 1103 116 1107
rect 1094 1107 1100 1108
rect 1382 1107 1388 1108
rect 1422 1112 1428 1113
rect 1422 1108 1423 1112
rect 1427 1108 1428 1112
rect 1422 1107 1428 1108
rect 1470 1112 1476 1113
rect 1470 1108 1471 1112
rect 1475 1108 1476 1112
rect 1470 1107 1476 1108
rect 1526 1112 1532 1113
rect 1526 1108 1527 1112
rect 1531 1108 1532 1112
rect 1526 1107 1532 1108
rect 1590 1112 1596 1113
rect 1590 1108 1591 1112
rect 1595 1108 1596 1112
rect 1590 1107 1596 1108
rect 1654 1112 1660 1113
rect 1654 1108 1655 1112
rect 1659 1108 1660 1112
rect 1654 1107 1660 1108
rect 1710 1112 1716 1113
rect 1710 1108 1711 1112
rect 1715 1108 1716 1112
rect 1710 1107 1716 1108
rect 1766 1112 1772 1113
rect 1766 1108 1767 1112
rect 1771 1108 1772 1112
rect 1766 1107 1772 1108
rect 1822 1112 1828 1113
rect 1822 1108 1823 1112
rect 1827 1108 1828 1112
rect 1822 1107 1828 1108
rect 1870 1112 1876 1113
rect 1870 1108 1871 1112
rect 1875 1108 1876 1112
rect 1870 1107 1876 1108
rect 1926 1112 1932 1113
rect 1926 1108 1927 1112
rect 1931 1108 1932 1112
rect 1926 1107 1932 1108
rect 1982 1112 1988 1113
rect 1982 1108 1983 1112
rect 1987 1108 1988 1112
rect 1982 1107 1988 1108
rect 2030 1112 2036 1113
rect 2030 1108 2031 1112
rect 2035 1108 2036 1112
rect 2030 1107 2036 1108
rect 2070 1112 2076 1113
rect 2070 1108 2071 1112
rect 2075 1108 2076 1112
rect 2070 1107 2076 1108
rect 110 1102 116 1103
rect 158 1104 164 1105
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 198 1104 204 1105
rect 198 1100 199 1104
rect 203 1100 204 1104
rect 198 1099 204 1100
rect 246 1104 252 1105
rect 246 1100 247 1104
rect 251 1100 252 1104
rect 246 1099 252 1100
rect 302 1104 308 1105
rect 302 1100 303 1104
rect 307 1100 308 1104
rect 302 1099 308 1100
rect 366 1104 372 1105
rect 366 1100 367 1104
rect 371 1100 372 1104
rect 366 1099 372 1100
rect 438 1104 444 1105
rect 438 1100 439 1104
rect 443 1100 444 1104
rect 438 1099 444 1100
rect 510 1104 516 1105
rect 510 1100 511 1104
rect 515 1100 516 1104
rect 510 1099 516 1100
rect 590 1104 596 1105
rect 590 1100 591 1104
rect 595 1100 596 1104
rect 590 1099 596 1100
rect 678 1104 684 1105
rect 678 1100 679 1104
rect 683 1100 684 1104
rect 678 1099 684 1100
rect 774 1104 780 1105
rect 774 1100 775 1104
rect 779 1100 780 1104
rect 774 1099 780 1100
rect 878 1104 884 1105
rect 878 1100 879 1104
rect 883 1100 884 1104
rect 878 1099 884 1100
rect 990 1104 996 1105
rect 990 1100 991 1104
rect 995 1100 996 1104
rect 1094 1103 1095 1107
rect 1099 1103 1100 1107
rect 1094 1102 1100 1103
rect 1134 1104 1140 1105
rect 990 1099 996 1100
rect 1134 1100 1135 1104
rect 1139 1100 1140 1104
rect 1134 1099 1140 1100
rect 2118 1104 2124 1105
rect 2118 1100 2119 1104
rect 2123 1100 2124 1104
rect 2118 1099 2124 1100
rect 1134 1087 1140 1088
rect 198 1084 204 1085
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 198 1080 199 1084
rect 203 1080 204 1084
rect 198 1079 204 1080
rect 246 1084 252 1085
rect 246 1080 247 1084
rect 251 1080 252 1084
rect 246 1079 252 1080
rect 302 1084 308 1085
rect 302 1080 303 1084
rect 307 1080 308 1084
rect 302 1079 308 1080
rect 366 1084 372 1085
rect 366 1080 367 1084
rect 371 1080 372 1084
rect 366 1079 372 1080
rect 430 1084 436 1085
rect 430 1080 431 1084
rect 435 1080 436 1084
rect 430 1079 436 1080
rect 502 1084 508 1085
rect 502 1080 503 1084
rect 507 1080 508 1084
rect 502 1079 508 1080
rect 574 1084 580 1085
rect 574 1080 575 1084
rect 579 1080 580 1084
rect 574 1079 580 1080
rect 646 1084 652 1085
rect 646 1080 647 1084
rect 651 1080 652 1084
rect 646 1079 652 1080
rect 718 1084 724 1085
rect 718 1080 719 1084
rect 723 1080 724 1084
rect 718 1079 724 1080
rect 782 1084 788 1085
rect 782 1080 783 1084
rect 787 1080 788 1084
rect 782 1079 788 1080
rect 838 1084 844 1085
rect 838 1080 839 1084
rect 843 1080 844 1084
rect 838 1079 844 1080
rect 894 1084 900 1085
rect 894 1080 895 1084
rect 899 1080 900 1084
rect 894 1079 900 1080
rect 950 1084 956 1085
rect 950 1080 951 1084
rect 955 1080 956 1084
rect 950 1079 956 1080
rect 1006 1084 1012 1085
rect 1006 1080 1007 1084
rect 1011 1080 1012 1084
rect 1006 1079 1012 1080
rect 1046 1084 1052 1085
rect 1046 1080 1047 1084
rect 1051 1080 1052 1084
rect 1134 1083 1135 1087
rect 1139 1083 1140 1087
rect 2118 1087 2124 1088
rect 1134 1082 1140 1083
rect 1382 1084 1388 1085
rect 1046 1079 1052 1080
rect 1094 1081 1100 1082
rect 110 1076 116 1077
rect 1094 1077 1095 1081
rect 1099 1077 1100 1081
rect 1382 1080 1383 1084
rect 1387 1080 1388 1084
rect 1382 1079 1388 1080
rect 1422 1084 1428 1085
rect 1422 1080 1423 1084
rect 1427 1080 1428 1084
rect 1422 1079 1428 1080
rect 1470 1084 1476 1085
rect 1470 1080 1471 1084
rect 1475 1080 1476 1084
rect 1470 1079 1476 1080
rect 1526 1084 1532 1085
rect 1526 1080 1527 1084
rect 1531 1080 1532 1084
rect 1526 1079 1532 1080
rect 1590 1084 1596 1085
rect 1590 1080 1591 1084
rect 1595 1080 1596 1084
rect 1590 1079 1596 1080
rect 1654 1084 1660 1085
rect 1654 1080 1655 1084
rect 1659 1080 1660 1084
rect 1654 1079 1660 1080
rect 1710 1084 1716 1085
rect 1710 1080 1711 1084
rect 1715 1080 1716 1084
rect 1710 1079 1716 1080
rect 1766 1084 1772 1085
rect 1766 1080 1767 1084
rect 1771 1080 1772 1084
rect 1766 1079 1772 1080
rect 1822 1084 1828 1085
rect 1822 1080 1823 1084
rect 1827 1080 1828 1084
rect 1822 1079 1828 1080
rect 1870 1084 1876 1085
rect 1870 1080 1871 1084
rect 1875 1080 1876 1084
rect 1870 1079 1876 1080
rect 1926 1084 1932 1085
rect 1926 1080 1927 1084
rect 1931 1080 1932 1084
rect 1926 1079 1932 1080
rect 1982 1084 1988 1085
rect 1982 1080 1983 1084
rect 1987 1080 1988 1084
rect 1982 1079 1988 1080
rect 2030 1084 2036 1085
rect 2030 1080 2031 1084
rect 2035 1080 2036 1084
rect 2030 1079 2036 1080
rect 2070 1084 2076 1085
rect 2070 1080 2071 1084
rect 2075 1080 2076 1084
rect 2118 1083 2119 1087
rect 2123 1083 2124 1087
rect 2118 1082 2124 1083
rect 2070 1079 2076 1080
rect 1094 1076 1100 1077
rect 1158 1072 1164 1073
rect 1134 1069 1140 1070
rect 1134 1065 1135 1069
rect 1139 1065 1140 1069
rect 1158 1068 1159 1072
rect 1163 1068 1164 1072
rect 1158 1067 1164 1068
rect 1246 1072 1252 1073
rect 1246 1068 1247 1072
rect 1251 1068 1252 1072
rect 1246 1067 1252 1068
rect 1358 1072 1364 1073
rect 1358 1068 1359 1072
rect 1363 1068 1364 1072
rect 1358 1067 1364 1068
rect 1470 1072 1476 1073
rect 1470 1068 1471 1072
rect 1475 1068 1476 1072
rect 1470 1067 1476 1068
rect 1574 1072 1580 1073
rect 1574 1068 1575 1072
rect 1579 1068 1580 1072
rect 1574 1067 1580 1068
rect 1670 1072 1676 1073
rect 1670 1068 1671 1072
rect 1675 1068 1676 1072
rect 1670 1067 1676 1068
rect 1758 1072 1764 1073
rect 1758 1068 1759 1072
rect 1763 1068 1764 1072
rect 1758 1067 1764 1068
rect 1846 1072 1852 1073
rect 1846 1068 1847 1072
rect 1851 1068 1852 1072
rect 1846 1067 1852 1068
rect 1926 1072 1932 1073
rect 1926 1068 1927 1072
rect 1931 1068 1932 1072
rect 1926 1067 1932 1068
rect 2006 1072 2012 1073
rect 2006 1068 2007 1072
rect 2011 1068 2012 1072
rect 2006 1067 2012 1068
rect 2070 1072 2076 1073
rect 2070 1068 2071 1072
rect 2075 1068 2076 1072
rect 2070 1067 2076 1068
rect 2118 1069 2124 1070
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 110 1059 116 1060
rect 1094 1064 1100 1065
rect 1134 1064 1140 1065
rect 2118 1065 2119 1069
rect 2123 1065 2124 1069
rect 2118 1064 2124 1065
rect 1094 1060 1095 1064
rect 1099 1060 1100 1064
rect 1094 1059 1100 1060
rect 198 1056 204 1057
rect 198 1052 199 1056
rect 203 1052 204 1056
rect 198 1051 204 1052
rect 246 1056 252 1057
rect 246 1052 247 1056
rect 251 1052 252 1056
rect 246 1051 252 1052
rect 302 1056 308 1057
rect 302 1052 303 1056
rect 307 1052 308 1056
rect 302 1051 308 1052
rect 366 1056 372 1057
rect 366 1052 367 1056
rect 371 1052 372 1056
rect 366 1051 372 1052
rect 430 1056 436 1057
rect 430 1052 431 1056
rect 435 1052 436 1056
rect 430 1051 436 1052
rect 502 1056 508 1057
rect 502 1052 503 1056
rect 507 1052 508 1056
rect 502 1051 508 1052
rect 574 1056 580 1057
rect 574 1052 575 1056
rect 579 1052 580 1056
rect 574 1051 580 1052
rect 646 1056 652 1057
rect 646 1052 647 1056
rect 651 1052 652 1056
rect 646 1051 652 1052
rect 718 1056 724 1057
rect 718 1052 719 1056
rect 723 1052 724 1056
rect 718 1051 724 1052
rect 782 1056 788 1057
rect 782 1052 783 1056
rect 787 1052 788 1056
rect 782 1051 788 1052
rect 838 1056 844 1057
rect 838 1052 839 1056
rect 843 1052 844 1056
rect 838 1051 844 1052
rect 894 1056 900 1057
rect 894 1052 895 1056
rect 899 1052 900 1056
rect 894 1051 900 1052
rect 950 1056 956 1057
rect 950 1052 951 1056
rect 955 1052 956 1056
rect 950 1051 956 1052
rect 1006 1056 1012 1057
rect 1006 1052 1007 1056
rect 1011 1052 1012 1056
rect 1006 1051 1012 1052
rect 1046 1056 1052 1057
rect 1046 1052 1047 1056
rect 1051 1052 1052 1056
rect 1046 1051 1052 1052
rect 1134 1052 1140 1053
rect 1134 1048 1135 1052
rect 1139 1048 1140 1052
rect 1134 1047 1140 1048
rect 2118 1052 2124 1053
rect 2118 1048 2119 1052
rect 2123 1048 2124 1052
rect 2118 1047 2124 1048
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1246 1044 1252 1045
rect 1246 1040 1247 1044
rect 1251 1040 1252 1044
rect 1246 1039 1252 1040
rect 1358 1044 1364 1045
rect 1358 1040 1359 1044
rect 1363 1040 1364 1044
rect 1358 1039 1364 1040
rect 1470 1044 1476 1045
rect 1470 1040 1471 1044
rect 1475 1040 1476 1044
rect 1470 1039 1476 1040
rect 1574 1044 1580 1045
rect 1574 1040 1575 1044
rect 1579 1040 1580 1044
rect 1574 1039 1580 1040
rect 1670 1044 1676 1045
rect 1670 1040 1671 1044
rect 1675 1040 1676 1044
rect 1670 1039 1676 1040
rect 1758 1044 1764 1045
rect 1758 1040 1759 1044
rect 1763 1040 1764 1044
rect 1758 1039 1764 1040
rect 1846 1044 1852 1045
rect 1846 1040 1847 1044
rect 1851 1040 1852 1044
rect 1846 1039 1852 1040
rect 1926 1044 1932 1045
rect 1926 1040 1927 1044
rect 1931 1040 1932 1044
rect 1926 1039 1932 1040
rect 2006 1044 2012 1045
rect 2006 1040 2007 1044
rect 2011 1040 2012 1044
rect 2006 1039 2012 1040
rect 2070 1044 2076 1045
rect 2070 1040 2071 1044
rect 2075 1040 2076 1044
rect 2070 1039 2076 1040
rect 222 1016 228 1017
rect 222 1012 223 1016
rect 227 1012 228 1016
rect 222 1011 228 1012
rect 270 1016 276 1017
rect 270 1012 271 1016
rect 275 1012 276 1016
rect 270 1011 276 1012
rect 334 1016 340 1017
rect 334 1012 335 1016
rect 339 1012 340 1016
rect 334 1011 340 1012
rect 406 1016 412 1017
rect 406 1012 407 1016
rect 411 1012 412 1016
rect 406 1011 412 1012
rect 478 1016 484 1017
rect 478 1012 479 1016
rect 483 1012 484 1016
rect 478 1011 484 1012
rect 558 1016 564 1017
rect 558 1012 559 1016
rect 563 1012 564 1016
rect 558 1011 564 1012
rect 630 1016 636 1017
rect 630 1012 631 1016
rect 635 1012 636 1016
rect 630 1011 636 1012
rect 702 1016 708 1017
rect 702 1012 703 1016
rect 707 1012 708 1016
rect 702 1011 708 1012
rect 774 1016 780 1017
rect 774 1012 775 1016
rect 779 1012 780 1016
rect 774 1011 780 1012
rect 838 1016 844 1017
rect 838 1012 839 1016
rect 843 1012 844 1016
rect 838 1011 844 1012
rect 902 1016 908 1017
rect 902 1012 903 1016
rect 907 1012 908 1016
rect 902 1011 908 1012
rect 966 1016 972 1017
rect 966 1012 967 1016
rect 971 1012 972 1016
rect 966 1011 972 1012
rect 1038 1016 1044 1017
rect 1038 1012 1039 1016
rect 1043 1012 1044 1016
rect 1038 1011 1044 1012
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 1094 1008 1100 1009
rect 1094 1004 1095 1008
rect 1099 1004 1100 1008
rect 1094 1003 1100 1004
rect 1158 1008 1164 1009
rect 1158 1004 1159 1008
rect 1163 1004 1164 1008
rect 1158 1003 1164 1004
rect 1230 1008 1236 1009
rect 1230 1004 1231 1008
rect 1235 1004 1236 1008
rect 1230 1003 1236 1004
rect 1302 1008 1308 1009
rect 1302 1004 1303 1008
rect 1307 1004 1308 1008
rect 1302 1003 1308 1004
rect 1382 1008 1388 1009
rect 1382 1004 1383 1008
rect 1387 1004 1388 1008
rect 1382 1003 1388 1004
rect 1462 1008 1468 1009
rect 1462 1004 1463 1008
rect 1467 1004 1468 1008
rect 1462 1003 1468 1004
rect 1542 1008 1548 1009
rect 1542 1004 1543 1008
rect 1547 1004 1548 1008
rect 1542 1003 1548 1004
rect 1622 1008 1628 1009
rect 1622 1004 1623 1008
rect 1627 1004 1628 1008
rect 1622 1003 1628 1004
rect 1694 1008 1700 1009
rect 1694 1004 1695 1008
rect 1699 1004 1700 1008
rect 1694 1003 1700 1004
rect 1758 1008 1764 1009
rect 1758 1004 1759 1008
rect 1763 1004 1764 1008
rect 1758 1003 1764 1004
rect 1822 1008 1828 1009
rect 1822 1004 1823 1008
rect 1827 1004 1828 1008
rect 1822 1003 1828 1004
rect 1886 1008 1892 1009
rect 1886 1004 1887 1008
rect 1891 1004 1892 1008
rect 1886 1003 1892 1004
rect 1950 1008 1956 1009
rect 1950 1004 1951 1008
rect 1955 1004 1956 1008
rect 1950 1003 1956 1004
rect 1134 1000 1140 1001
rect 1134 996 1135 1000
rect 1139 996 1140 1000
rect 1134 995 1140 996
rect 2118 1000 2124 1001
rect 2118 996 2119 1000
rect 2123 996 2124 1000
rect 2118 995 2124 996
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1094 991 1100 992
rect 110 986 116 987
rect 222 988 228 989
rect 222 984 223 988
rect 227 984 228 988
rect 222 983 228 984
rect 270 988 276 989
rect 270 984 271 988
rect 275 984 276 988
rect 270 983 276 984
rect 334 988 340 989
rect 334 984 335 988
rect 339 984 340 988
rect 334 983 340 984
rect 406 988 412 989
rect 406 984 407 988
rect 411 984 412 988
rect 406 983 412 984
rect 478 988 484 989
rect 478 984 479 988
rect 483 984 484 988
rect 478 983 484 984
rect 558 988 564 989
rect 558 984 559 988
rect 563 984 564 988
rect 558 983 564 984
rect 630 988 636 989
rect 630 984 631 988
rect 635 984 636 988
rect 630 983 636 984
rect 702 988 708 989
rect 702 984 703 988
rect 707 984 708 988
rect 702 983 708 984
rect 774 988 780 989
rect 774 984 775 988
rect 779 984 780 988
rect 774 983 780 984
rect 838 988 844 989
rect 838 984 839 988
rect 843 984 844 988
rect 838 983 844 984
rect 902 988 908 989
rect 902 984 903 988
rect 907 984 908 988
rect 902 983 908 984
rect 966 988 972 989
rect 966 984 967 988
rect 971 984 972 988
rect 966 983 972 984
rect 1038 988 1044 989
rect 1038 984 1039 988
rect 1043 984 1044 988
rect 1094 987 1095 991
rect 1099 987 1100 991
rect 1094 986 1100 987
rect 1038 983 1044 984
rect 1134 983 1140 984
rect 1134 979 1135 983
rect 1139 979 1140 983
rect 2118 983 2124 984
rect 1134 978 1140 979
rect 1158 980 1164 981
rect 1158 976 1159 980
rect 1163 976 1164 980
rect 1158 975 1164 976
rect 1230 980 1236 981
rect 1230 976 1231 980
rect 1235 976 1236 980
rect 1230 975 1236 976
rect 1302 980 1308 981
rect 1302 976 1303 980
rect 1307 976 1308 980
rect 1302 975 1308 976
rect 1382 980 1388 981
rect 1382 976 1383 980
rect 1387 976 1388 980
rect 1382 975 1388 976
rect 1462 980 1468 981
rect 1462 976 1463 980
rect 1467 976 1468 980
rect 1462 975 1468 976
rect 1542 980 1548 981
rect 1542 976 1543 980
rect 1547 976 1548 980
rect 1542 975 1548 976
rect 1622 980 1628 981
rect 1622 976 1623 980
rect 1627 976 1628 980
rect 1622 975 1628 976
rect 1694 980 1700 981
rect 1694 976 1695 980
rect 1699 976 1700 980
rect 1694 975 1700 976
rect 1758 980 1764 981
rect 1758 976 1759 980
rect 1763 976 1764 980
rect 1758 975 1764 976
rect 1822 980 1828 981
rect 1822 976 1823 980
rect 1827 976 1828 980
rect 1822 975 1828 976
rect 1886 980 1892 981
rect 1886 976 1887 980
rect 1891 976 1892 980
rect 1886 975 1892 976
rect 1950 980 1956 981
rect 1950 976 1951 980
rect 1955 976 1956 980
rect 2118 979 2119 983
rect 2123 979 2124 983
rect 2118 978 2124 979
rect 1950 975 1956 976
rect 150 972 156 973
rect 110 969 116 970
rect 110 965 111 969
rect 115 965 116 969
rect 150 968 151 972
rect 155 968 156 972
rect 150 967 156 968
rect 214 972 220 973
rect 214 968 215 972
rect 219 968 220 972
rect 214 967 220 968
rect 286 972 292 973
rect 286 968 287 972
rect 291 968 292 972
rect 286 967 292 968
rect 366 972 372 973
rect 366 968 367 972
rect 371 968 372 972
rect 366 967 372 968
rect 446 972 452 973
rect 446 968 447 972
rect 451 968 452 972
rect 446 967 452 968
rect 526 972 532 973
rect 526 968 527 972
rect 531 968 532 972
rect 526 967 532 968
rect 598 972 604 973
rect 598 968 599 972
rect 603 968 604 972
rect 598 967 604 968
rect 670 972 676 973
rect 670 968 671 972
rect 675 968 676 972
rect 670 967 676 968
rect 734 972 740 973
rect 734 968 735 972
rect 739 968 740 972
rect 734 967 740 968
rect 798 972 804 973
rect 798 968 799 972
rect 803 968 804 972
rect 798 967 804 968
rect 862 972 868 973
rect 862 968 863 972
rect 867 968 868 972
rect 862 967 868 968
rect 926 972 932 973
rect 926 968 927 972
rect 931 968 932 972
rect 926 967 932 968
rect 990 972 996 973
rect 990 968 991 972
rect 995 968 996 972
rect 990 967 996 968
rect 1046 972 1052 973
rect 1046 968 1047 972
rect 1051 968 1052 972
rect 1046 967 1052 968
rect 1094 969 1100 970
rect 110 964 116 965
rect 1094 965 1095 969
rect 1099 965 1100 969
rect 1238 968 1244 969
rect 1094 964 1100 965
rect 1134 965 1140 966
rect 1134 961 1135 965
rect 1139 961 1140 965
rect 1238 964 1239 968
rect 1243 964 1244 968
rect 1238 963 1244 964
rect 1302 968 1308 969
rect 1302 964 1303 968
rect 1307 964 1308 968
rect 1302 963 1308 964
rect 1374 968 1380 969
rect 1374 964 1375 968
rect 1379 964 1380 968
rect 1374 963 1380 964
rect 1438 968 1444 969
rect 1438 964 1439 968
rect 1443 964 1444 968
rect 1438 963 1444 964
rect 1510 968 1516 969
rect 1510 964 1511 968
rect 1515 964 1516 968
rect 1510 963 1516 964
rect 1582 968 1588 969
rect 1582 964 1583 968
rect 1587 964 1588 968
rect 1582 963 1588 964
rect 1654 968 1660 969
rect 1654 964 1655 968
rect 1659 964 1660 968
rect 1654 963 1660 964
rect 1726 968 1732 969
rect 1726 964 1727 968
rect 1731 964 1732 968
rect 1726 963 1732 964
rect 1798 968 1804 969
rect 1798 964 1799 968
rect 1803 964 1804 968
rect 1798 963 1804 964
rect 1870 968 1876 969
rect 1870 964 1871 968
rect 1875 964 1876 968
rect 1870 963 1876 964
rect 1942 968 1948 969
rect 1942 964 1943 968
rect 1947 964 1948 968
rect 1942 963 1948 964
rect 2014 968 2020 969
rect 2014 964 2015 968
rect 2019 964 2020 968
rect 2014 963 2020 964
rect 2070 968 2076 969
rect 2070 964 2071 968
rect 2075 964 2076 968
rect 2070 963 2076 964
rect 2118 965 2124 966
rect 1134 960 1140 961
rect 2118 961 2119 965
rect 2123 961 2124 965
rect 2118 960 2124 961
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 110 947 116 948
rect 1094 952 1100 953
rect 1094 948 1095 952
rect 1099 948 1100 952
rect 1094 947 1100 948
rect 1134 948 1140 949
rect 150 944 156 945
rect 150 940 151 944
rect 155 940 156 944
rect 150 939 156 940
rect 214 944 220 945
rect 214 940 215 944
rect 219 940 220 944
rect 214 939 220 940
rect 286 944 292 945
rect 286 940 287 944
rect 291 940 292 944
rect 286 939 292 940
rect 366 944 372 945
rect 366 940 367 944
rect 371 940 372 944
rect 366 939 372 940
rect 446 944 452 945
rect 446 940 447 944
rect 451 940 452 944
rect 446 939 452 940
rect 526 944 532 945
rect 526 940 527 944
rect 531 940 532 944
rect 526 939 532 940
rect 598 944 604 945
rect 598 940 599 944
rect 603 940 604 944
rect 598 939 604 940
rect 670 944 676 945
rect 670 940 671 944
rect 675 940 676 944
rect 670 939 676 940
rect 734 944 740 945
rect 734 940 735 944
rect 739 940 740 944
rect 734 939 740 940
rect 798 944 804 945
rect 798 940 799 944
rect 803 940 804 944
rect 798 939 804 940
rect 862 944 868 945
rect 862 940 863 944
rect 867 940 868 944
rect 862 939 868 940
rect 926 944 932 945
rect 926 940 927 944
rect 931 940 932 944
rect 926 939 932 940
rect 990 944 996 945
rect 990 940 991 944
rect 995 940 996 944
rect 990 939 996 940
rect 1046 944 1052 945
rect 1046 940 1047 944
rect 1051 940 1052 944
rect 1134 944 1135 948
rect 1139 944 1140 948
rect 1134 943 1140 944
rect 2118 948 2124 949
rect 2118 944 2119 948
rect 2123 944 2124 948
rect 2118 943 2124 944
rect 1046 939 1052 940
rect 1238 940 1244 941
rect 1238 936 1239 940
rect 1243 936 1244 940
rect 1238 935 1244 936
rect 1302 940 1308 941
rect 1302 936 1303 940
rect 1307 936 1308 940
rect 1302 935 1308 936
rect 1374 940 1380 941
rect 1374 936 1375 940
rect 1379 936 1380 940
rect 1374 935 1380 936
rect 1438 940 1444 941
rect 1438 936 1439 940
rect 1443 936 1444 940
rect 1438 935 1444 936
rect 1510 940 1516 941
rect 1510 936 1511 940
rect 1515 936 1516 940
rect 1510 935 1516 936
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1654 940 1660 941
rect 1654 936 1655 940
rect 1659 936 1660 940
rect 1654 935 1660 936
rect 1726 940 1732 941
rect 1726 936 1727 940
rect 1731 936 1732 940
rect 1726 935 1732 936
rect 1798 940 1804 941
rect 1798 936 1799 940
rect 1803 936 1804 940
rect 1798 935 1804 936
rect 1870 940 1876 941
rect 1870 936 1871 940
rect 1875 936 1876 940
rect 1870 935 1876 936
rect 1942 940 1948 941
rect 1942 936 1943 940
rect 1947 936 1948 940
rect 1942 935 1948 936
rect 2014 940 2020 941
rect 2014 936 2015 940
rect 2019 936 2020 940
rect 2014 935 2020 936
rect 2070 940 2076 941
rect 2070 936 2071 940
rect 2075 936 2076 940
rect 2070 935 2076 936
rect 134 908 140 909
rect 134 904 135 908
rect 139 904 140 908
rect 134 903 140 904
rect 182 908 188 909
rect 182 904 183 908
rect 187 904 188 908
rect 182 903 188 904
rect 254 908 260 909
rect 254 904 255 908
rect 259 904 260 908
rect 254 903 260 904
rect 326 908 332 909
rect 326 904 327 908
rect 331 904 332 908
rect 326 903 332 904
rect 398 908 404 909
rect 398 904 399 908
rect 403 904 404 908
rect 398 903 404 904
rect 462 908 468 909
rect 462 904 463 908
rect 467 904 468 908
rect 462 903 468 904
rect 526 908 532 909
rect 526 904 527 908
rect 531 904 532 908
rect 526 903 532 904
rect 598 908 604 909
rect 598 904 599 908
rect 603 904 604 908
rect 598 903 604 904
rect 670 908 676 909
rect 670 904 671 908
rect 675 904 676 908
rect 670 903 676 904
rect 742 908 748 909
rect 742 904 743 908
rect 747 904 748 908
rect 742 903 748 904
rect 814 908 820 909
rect 814 904 815 908
rect 819 904 820 908
rect 814 903 820 904
rect 894 908 900 909
rect 894 904 895 908
rect 899 904 900 908
rect 894 903 900 904
rect 982 908 988 909
rect 982 904 983 908
rect 987 904 988 908
rect 982 903 988 904
rect 1046 908 1052 909
rect 1046 904 1047 908
rect 1051 904 1052 908
rect 1046 903 1052 904
rect 110 900 116 901
rect 110 896 111 900
rect 115 896 116 900
rect 110 895 116 896
rect 1094 900 1100 901
rect 1094 896 1095 900
rect 1099 896 1100 900
rect 1094 895 1100 896
rect 1286 900 1292 901
rect 1286 896 1287 900
rect 1291 896 1292 900
rect 1286 895 1292 896
rect 1326 900 1332 901
rect 1326 896 1327 900
rect 1331 896 1332 900
rect 1326 895 1332 896
rect 1374 900 1380 901
rect 1374 896 1375 900
rect 1379 896 1380 900
rect 1374 895 1380 896
rect 1422 900 1428 901
rect 1422 896 1423 900
rect 1427 896 1428 900
rect 1422 895 1428 896
rect 1478 900 1484 901
rect 1478 896 1479 900
rect 1483 896 1484 900
rect 1478 895 1484 896
rect 1550 900 1556 901
rect 1550 896 1551 900
rect 1555 896 1556 900
rect 1550 895 1556 896
rect 1622 900 1628 901
rect 1622 896 1623 900
rect 1627 896 1628 900
rect 1622 895 1628 896
rect 1702 900 1708 901
rect 1702 896 1703 900
rect 1707 896 1708 900
rect 1702 895 1708 896
rect 1790 900 1796 901
rect 1790 896 1791 900
rect 1795 896 1796 900
rect 1790 895 1796 896
rect 1878 900 1884 901
rect 1878 896 1879 900
rect 1883 896 1884 900
rect 1878 895 1884 896
rect 1966 900 1972 901
rect 1966 896 1967 900
rect 1971 896 1972 900
rect 1966 895 1972 896
rect 2062 900 2068 901
rect 2062 896 2063 900
rect 2067 896 2068 900
rect 2062 895 2068 896
rect 1134 892 1140 893
rect 1134 888 1135 892
rect 1139 888 1140 892
rect 1134 887 1140 888
rect 2118 892 2124 893
rect 2118 888 2119 892
rect 2123 888 2124 892
rect 2118 887 2124 888
rect 110 883 116 884
rect 110 879 111 883
rect 115 879 116 883
rect 1094 883 1100 884
rect 110 878 116 879
rect 134 880 140 881
rect 134 876 135 880
rect 139 876 140 880
rect 134 875 140 876
rect 182 880 188 881
rect 182 876 183 880
rect 187 876 188 880
rect 182 875 188 876
rect 254 880 260 881
rect 254 876 255 880
rect 259 876 260 880
rect 254 875 260 876
rect 326 880 332 881
rect 326 876 327 880
rect 331 876 332 880
rect 326 875 332 876
rect 398 880 404 881
rect 398 876 399 880
rect 403 876 404 880
rect 398 875 404 876
rect 462 880 468 881
rect 462 876 463 880
rect 467 876 468 880
rect 462 875 468 876
rect 526 880 532 881
rect 526 876 527 880
rect 531 876 532 880
rect 526 875 532 876
rect 598 880 604 881
rect 598 876 599 880
rect 603 876 604 880
rect 598 875 604 876
rect 670 880 676 881
rect 670 876 671 880
rect 675 876 676 880
rect 670 875 676 876
rect 742 880 748 881
rect 742 876 743 880
rect 747 876 748 880
rect 742 875 748 876
rect 814 880 820 881
rect 814 876 815 880
rect 819 876 820 880
rect 814 875 820 876
rect 894 880 900 881
rect 894 876 895 880
rect 899 876 900 880
rect 894 875 900 876
rect 982 880 988 881
rect 982 876 983 880
rect 987 876 988 880
rect 982 875 988 876
rect 1046 880 1052 881
rect 1046 876 1047 880
rect 1051 876 1052 880
rect 1094 879 1095 883
rect 1099 879 1100 883
rect 1094 878 1100 879
rect 1046 875 1052 876
rect 1134 875 1140 876
rect 1134 871 1135 875
rect 1139 871 1140 875
rect 2118 875 2124 876
rect 1134 870 1140 871
rect 1286 872 1292 873
rect 1286 868 1287 872
rect 1291 868 1292 872
rect 1286 867 1292 868
rect 1326 872 1332 873
rect 1326 868 1327 872
rect 1331 868 1332 872
rect 1326 867 1332 868
rect 1374 872 1380 873
rect 1374 868 1375 872
rect 1379 868 1380 872
rect 1374 867 1380 868
rect 1422 872 1428 873
rect 1422 868 1423 872
rect 1427 868 1428 872
rect 1422 867 1428 868
rect 1478 872 1484 873
rect 1478 868 1479 872
rect 1483 868 1484 872
rect 1478 867 1484 868
rect 1550 872 1556 873
rect 1550 868 1551 872
rect 1555 868 1556 872
rect 1550 867 1556 868
rect 1622 872 1628 873
rect 1622 868 1623 872
rect 1627 868 1628 872
rect 1622 867 1628 868
rect 1702 872 1708 873
rect 1702 868 1703 872
rect 1707 868 1708 872
rect 1702 867 1708 868
rect 1790 872 1796 873
rect 1790 868 1791 872
rect 1795 868 1796 872
rect 1790 867 1796 868
rect 1878 872 1884 873
rect 1878 868 1879 872
rect 1883 868 1884 872
rect 1878 867 1884 868
rect 1966 872 1972 873
rect 1966 868 1967 872
rect 1971 868 1972 872
rect 1966 867 1972 868
rect 2062 872 2068 873
rect 2062 868 2063 872
rect 2067 868 2068 872
rect 2118 871 2119 875
rect 2123 871 2124 875
rect 2118 870 2124 871
rect 2062 867 2068 868
rect 134 864 140 865
rect 110 861 116 862
rect 110 857 111 861
rect 115 857 116 861
rect 134 860 135 864
rect 139 860 140 864
rect 134 859 140 860
rect 174 864 180 865
rect 174 860 175 864
rect 179 860 180 864
rect 174 859 180 860
rect 214 864 220 865
rect 214 860 215 864
rect 219 860 220 864
rect 214 859 220 860
rect 278 864 284 865
rect 278 860 279 864
rect 283 860 284 864
rect 278 859 284 860
rect 342 864 348 865
rect 342 860 343 864
rect 347 860 348 864
rect 342 859 348 860
rect 398 864 404 865
rect 398 860 399 864
rect 403 860 404 864
rect 398 859 404 860
rect 462 864 468 865
rect 462 860 463 864
rect 467 860 468 864
rect 462 859 468 860
rect 534 864 540 865
rect 534 860 535 864
rect 539 860 540 864
rect 534 859 540 860
rect 614 864 620 865
rect 614 860 615 864
rect 619 860 620 864
rect 614 859 620 860
rect 710 864 716 865
rect 710 860 711 864
rect 715 860 716 864
rect 710 859 716 860
rect 822 864 828 865
rect 822 860 823 864
rect 827 860 828 864
rect 822 859 828 860
rect 942 864 948 865
rect 942 860 943 864
rect 947 860 948 864
rect 942 859 948 860
rect 1046 864 1052 865
rect 1046 860 1047 864
rect 1051 860 1052 864
rect 1046 859 1052 860
rect 1094 861 1100 862
rect 110 856 116 857
rect 1094 857 1095 861
rect 1099 857 1100 861
rect 1158 860 1164 861
rect 1094 856 1100 857
rect 1134 857 1140 858
rect 1134 853 1135 857
rect 1139 853 1140 857
rect 1158 856 1159 860
rect 1163 856 1164 860
rect 1158 855 1164 856
rect 1198 860 1204 861
rect 1198 856 1199 860
rect 1203 856 1204 860
rect 1198 855 1204 856
rect 1262 860 1268 861
rect 1262 856 1263 860
rect 1267 856 1268 860
rect 1262 855 1268 856
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1398 860 1404 861
rect 1398 856 1399 860
rect 1403 856 1404 860
rect 1398 855 1404 856
rect 1470 860 1476 861
rect 1470 856 1471 860
rect 1475 856 1476 860
rect 1470 855 1476 856
rect 1542 860 1548 861
rect 1542 856 1543 860
rect 1547 856 1548 860
rect 1542 855 1548 856
rect 1622 860 1628 861
rect 1622 856 1623 860
rect 1627 856 1628 860
rect 1622 855 1628 856
rect 1702 860 1708 861
rect 1702 856 1703 860
rect 1707 856 1708 860
rect 1702 855 1708 856
rect 1774 860 1780 861
rect 1774 856 1775 860
rect 1779 856 1780 860
rect 1774 855 1780 856
rect 1854 860 1860 861
rect 1854 856 1855 860
rect 1859 856 1860 860
rect 1854 855 1860 856
rect 1934 860 1940 861
rect 1934 856 1935 860
rect 1939 856 1940 860
rect 1934 855 1940 856
rect 2014 860 2020 861
rect 2014 856 2015 860
rect 2019 856 2020 860
rect 2014 855 2020 856
rect 2070 860 2076 861
rect 2070 856 2071 860
rect 2075 856 2076 860
rect 2070 855 2076 856
rect 2118 857 2124 858
rect 1134 852 1140 853
rect 2118 853 2119 857
rect 2123 853 2124 857
rect 2118 852 2124 853
rect 110 844 116 845
rect 110 840 111 844
rect 115 840 116 844
rect 110 839 116 840
rect 1094 844 1100 845
rect 1094 840 1095 844
rect 1099 840 1100 844
rect 1094 839 1100 840
rect 1134 840 1140 841
rect 134 836 140 837
rect 134 832 135 836
rect 139 832 140 836
rect 134 831 140 832
rect 174 836 180 837
rect 174 832 175 836
rect 179 832 180 836
rect 174 831 180 832
rect 214 836 220 837
rect 214 832 215 836
rect 219 832 220 836
rect 214 831 220 832
rect 278 836 284 837
rect 278 832 279 836
rect 283 832 284 836
rect 278 831 284 832
rect 342 836 348 837
rect 342 832 343 836
rect 347 832 348 836
rect 342 831 348 832
rect 398 836 404 837
rect 398 832 399 836
rect 403 832 404 836
rect 398 831 404 832
rect 462 836 468 837
rect 462 832 463 836
rect 467 832 468 836
rect 462 831 468 832
rect 534 836 540 837
rect 534 832 535 836
rect 539 832 540 836
rect 534 831 540 832
rect 614 836 620 837
rect 614 832 615 836
rect 619 832 620 836
rect 614 831 620 832
rect 710 836 716 837
rect 710 832 711 836
rect 715 832 716 836
rect 710 831 716 832
rect 822 836 828 837
rect 822 832 823 836
rect 827 832 828 836
rect 822 831 828 832
rect 942 836 948 837
rect 942 832 943 836
rect 947 832 948 836
rect 942 831 948 832
rect 1046 836 1052 837
rect 1046 832 1047 836
rect 1051 832 1052 836
rect 1134 836 1135 840
rect 1139 836 1140 840
rect 1134 835 1140 836
rect 2118 840 2124 841
rect 2118 836 2119 840
rect 2123 836 2124 840
rect 2118 835 2124 836
rect 1046 831 1052 832
rect 1158 832 1164 833
rect 1158 828 1159 832
rect 1163 828 1164 832
rect 1158 827 1164 828
rect 1198 832 1204 833
rect 1198 828 1199 832
rect 1203 828 1204 832
rect 1198 827 1204 828
rect 1262 832 1268 833
rect 1262 828 1263 832
rect 1267 828 1268 832
rect 1262 827 1268 828
rect 1326 832 1332 833
rect 1326 828 1327 832
rect 1331 828 1332 832
rect 1326 827 1332 828
rect 1398 832 1404 833
rect 1398 828 1399 832
rect 1403 828 1404 832
rect 1398 827 1404 828
rect 1470 832 1476 833
rect 1470 828 1471 832
rect 1475 828 1476 832
rect 1470 827 1476 828
rect 1542 832 1548 833
rect 1542 828 1543 832
rect 1547 828 1548 832
rect 1542 827 1548 828
rect 1622 832 1628 833
rect 1622 828 1623 832
rect 1627 828 1628 832
rect 1622 827 1628 828
rect 1702 832 1708 833
rect 1702 828 1703 832
rect 1707 828 1708 832
rect 1702 827 1708 828
rect 1774 832 1780 833
rect 1774 828 1775 832
rect 1779 828 1780 832
rect 1774 827 1780 828
rect 1854 832 1860 833
rect 1854 828 1855 832
rect 1859 828 1860 832
rect 1854 827 1860 828
rect 1934 832 1940 833
rect 1934 828 1935 832
rect 1939 828 1940 832
rect 1934 827 1940 828
rect 2014 832 2020 833
rect 2014 828 2015 832
rect 2019 828 2020 832
rect 2014 827 2020 828
rect 2070 832 2076 833
rect 2070 828 2071 832
rect 2075 828 2076 832
rect 2070 827 2076 828
rect 134 800 140 801
rect 134 796 135 800
rect 139 796 140 800
rect 134 795 140 796
rect 174 800 180 801
rect 174 796 175 800
rect 179 796 180 800
rect 174 795 180 796
rect 214 800 220 801
rect 214 796 215 800
rect 219 796 220 800
rect 214 795 220 796
rect 278 800 284 801
rect 278 796 279 800
rect 283 796 284 800
rect 278 795 284 796
rect 334 800 340 801
rect 334 796 335 800
rect 339 796 340 800
rect 334 795 340 796
rect 390 800 396 801
rect 390 796 391 800
rect 395 796 396 800
rect 390 795 396 796
rect 454 800 460 801
rect 454 796 455 800
rect 459 796 460 800
rect 454 795 460 796
rect 518 800 524 801
rect 518 796 519 800
rect 523 796 524 800
rect 518 795 524 796
rect 582 800 588 801
rect 582 796 583 800
rect 587 796 588 800
rect 582 795 588 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 734 800 740 801
rect 734 796 735 800
rect 739 796 740 800
rect 734 795 740 796
rect 814 800 820 801
rect 814 796 815 800
rect 819 796 820 800
rect 814 795 820 796
rect 894 800 900 801
rect 894 796 895 800
rect 899 796 900 800
rect 894 795 900 796
rect 982 800 988 801
rect 982 796 983 800
rect 987 796 988 800
rect 982 795 988 796
rect 1046 800 1052 801
rect 1046 796 1047 800
rect 1051 796 1052 800
rect 1046 795 1052 796
rect 110 792 116 793
rect 110 788 111 792
rect 115 788 116 792
rect 110 787 116 788
rect 1094 792 1100 793
rect 1094 788 1095 792
rect 1099 788 1100 792
rect 1094 787 1100 788
rect 1158 788 1164 789
rect 1158 784 1159 788
rect 1163 784 1164 788
rect 1158 783 1164 784
rect 1238 788 1244 789
rect 1238 784 1239 788
rect 1243 784 1244 788
rect 1238 783 1244 784
rect 1342 788 1348 789
rect 1342 784 1343 788
rect 1347 784 1348 788
rect 1342 783 1348 784
rect 1446 788 1452 789
rect 1446 784 1447 788
rect 1451 784 1452 788
rect 1446 783 1452 784
rect 1550 788 1556 789
rect 1550 784 1551 788
rect 1555 784 1556 788
rect 1550 783 1556 784
rect 1654 788 1660 789
rect 1654 784 1655 788
rect 1659 784 1660 788
rect 1654 783 1660 784
rect 1750 788 1756 789
rect 1750 784 1751 788
rect 1755 784 1756 788
rect 1750 783 1756 784
rect 1838 788 1844 789
rect 1838 784 1839 788
rect 1843 784 1844 788
rect 1838 783 1844 784
rect 1918 788 1924 789
rect 1918 784 1919 788
rect 1923 784 1924 788
rect 1918 783 1924 784
rect 2006 788 2012 789
rect 2006 784 2007 788
rect 2011 784 2012 788
rect 2006 783 2012 784
rect 2070 788 2076 789
rect 2070 784 2071 788
rect 2075 784 2076 788
rect 2070 783 2076 784
rect 1134 780 1140 781
rect 1134 776 1135 780
rect 1139 776 1140 780
rect 110 775 116 776
rect 110 771 111 775
rect 115 771 116 775
rect 1094 775 1100 776
rect 1134 775 1140 776
rect 2118 780 2124 781
rect 2118 776 2119 780
rect 2123 776 2124 780
rect 2118 775 2124 776
rect 110 770 116 771
rect 134 772 140 773
rect 134 768 135 772
rect 139 768 140 772
rect 134 767 140 768
rect 174 772 180 773
rect 174 768 175 772
rect 179 768 180 772
rect 174 767 180 768
rect 214 772 220 773
rect 214 768 215 772
rect 219 768 220 772
rect 214 767 220 768
rect 278 772 284 773
rect 278 768 279 772
rect 283 768 284 772
rect 278 767 284 768
rect 334 772 340 773
rect 334 768 335 772
rect 339 768 340 772
rect 334 767 340 768
rect 390 772 396 773
rect 390 768 391 772
rect 395 768 396 772
rect 390 767 396 768
rect 454 772 460 773
rect 454 768 455 772
rect 459 768 460 772
rect 454 767 460 768
rect 518 772 524 773
rect 518 768 519 772
rect 523 768 524 772
rect 518 767 524 768
rect 582 772 588 773
rect 582 768 583 772
rect 587 768 588 772
rect 582 767 588 768
rect 654 772 660 773
rect 654 768 655 772
rect 659 768 660 772
rect 654 767 660 768
rect 734 772 740 773
rect 734 768 735 772
rect 739 768 740 772
rect 734 767 740 768
rect 814 772 820 773
rect 814 768 815 772
rect 819 768 820 772
rect 814 767 820 768
rect 894 772 900 773
rect 894 768 895 772
rect 899 768 900 772
rect 894 767 900 768
rect 982 772 988 773
rect 982 768 983 772
rect 987 768 988 772
rect 982 767 988 768
rect 1046 772 1052 773
rect 1046 768 1047 772
rect 1051 768 1052 772
rect 1094 771 1095 775
rect 1099 771 1100 775
rect 1094 770 1100 771
rect 1046 767 1052 768
rect 1134 763 1140 764
rect 134 760 140 761
rect 110 757 116 758
rect 110 753 111 757
rect 115 753 116 757
rect 134 756 135 760
rect 139 756 140 760
rect 134 755 140 756
rect 206 760 212 761
rect 206 756 207 760
rect 211 756 212 760
rect 206 755 212 756
rect 294 760 300 761
rect 294 756 295 760
rect 299 756 300 760
rect 294 755 300 756
rect 374 760 380 761
rect 374 756 375 760
rect 379 756 380 760
rect 374 755 380 756
rect 446 760 452 761
rect 446 756 447 760
rect 451 756 452 760
rect 446 755 452 756
rect 518 760 524 761
rect 518 756 519 760
rect 523 756 524 760
rect 518 755 524 756
rect 582 760 588 761
rect 582 756 583 760
rect 587 756 588 760
rect 582 755 588 756
rect 638 760 644 761
rect 638 756 639 760
rect 643 756 644 760
rect 638 755 644 756
rect 686 760 692 761
rect 686 756 687 760
rect 691 756 692 760
rect 686 755 692 756
rect 742 760 748 761
rect 742 756 743 760
rect 747 756 748 760
rect 742 755 748 756
rect 798 760 804 761
rect 798 756 799 760
rect 803 756 804 760
rect 798 755 804 756
rect 854 760 860 761
rect 854 756 855 760
rect 859 756 860 760
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 2118 763 2124 764
rect 1134 758 1140 759
rect 1158 760 1164 761
rect 854 755 860 756
rect 1094 757 1100 758
rect 110 752 116 753
rect 1094 753 1095 757
rect 1099 753 1100 757
rect 1158 756 1159 760
rect 1163 756 1164 760
rect 1158 755 1164 756
rect 1238 760 1244 761
rect 1238 756 1239 760
rect 1243 756 1244 760
rect 1238 755 1244 756
rect 1342 760 1348 761
rect 1342 756 1343 760
rect 1347 756 1348 760
rect 1342 755 1348 756
rect 1446 760 1452 761
rect 1446 756 1447 760
rect 1451 756 1452 760
rect 1446 755 1452 756
rect 1550 760 1556 761
rect 1550 756 1551 760
rect 1555 756 1556 760
rect 1550 755 1556 756
rect 1654 760 1660 761
rect 1654 756 1655 760
rect 1659 756 1660 760
rect 1654 755 1660 756
rect 1750 760 1756 761
rect 1750 756 1751 760
rect 1755 756 1756 760
rect 1750 755 1756 756
rect 1838 760 1844 761
rect 1838 756 1839 760
rect 1843 756 1844 760
rect 1838 755 1844 756
rect 1918 760 1924 761
rect 1918 756 1919 760
rect 1923 756 1924 760
rect 1918 755 1924 756
rect 2006 760 2012 761
rect 2006 756 2007 760
rect 2011 756 2012 760
rect 2006 755 2012 756
rect 2070 760 2076 761
rect 2070 756 2071 760
rect 2075 756 2076 760
rect 2118 759 2119 763
rect 2123 759 2124 763
rect 2118 758 2124 759
rect 2070 755 2076 756
rect 1094 752 1100 753
rect 1158 748 1164 749
rect 1134 745 1140 746
rect 1134 741 1135 745
rect 1139 741 1140 745
rect 1158 744 1159 748
rect 1163 744 1164 748
rect 1158 743 1164 744
rect 1198 748 1204 749
rect 1198 744 1199 748
rect 1203 744 1204 748
rect 1198 743 1204 744
rect 1238 748 1244 749
rect 1238 744 1239 748
rect 1243 744 1244 748
rect 1238 743 1244 744
rect 1286 748 1292 749
rect 1286 744 1287 748
rect 1291 744 1292 748
rect 1286 743 1292 744
rect 1358 748 1364 749
rect 1358 744 1359 748
rect 1363 744 1364 748
rect 1358 743 1364 744
rect 1438 748 1444 749
rect 1438 744 1439 748
rect 1443 744 1444 748
rect 1438 743 1444 744
rect 1526 748 1532 749
rect 1526 744 1527 748
rect 1531 744 1532 748
rect 1526 743 1532 744
rect 1614 748 1620 749
rect 1614 744 1615 748
rect 1619 744 1620 748
rect 1614 743 1620 744
rect 1710 748 1716 749
rect 1710 744 1711 748
rect 1715 744 1716 748
rect 1710 743 1716 744
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 1806 743 1812 744
rect 1902 748 1908 749
rect 1902 744 1903 748
rect 1907 744 1908 748
rect 1902 743 1908 744
rect 1998 748 2004 749
rect 1998 744 1999 748
rect 2003 744 2004 748
rect 1998 743 2004 744
rect 2070 748 2076 749
rect 2070 744 2071 748
rect 2075 744 2076 748
rect 2070 743 2076 744
rect 2118 745 2124 746
rect 110 740 116 741
rect 110 736 111 740
rect 115 736 116 740
rect 110 735 116 736
rect 1094 740 1100 741
rect 1134 740 1140 741
rect 2118 741 2119 745
rect 2123 741 2124 745
rect 2118 740 2124 741
rect 1094 736 1095 740
rect 1099 736 1100 740
rect 1094 735 1100 736
rect 134 732 140 733
rect 134 728 135 732
rect 139 728 140 732
rect 134 727 140 728
rect 206 732 212 733
rect 206 728 207 732
rect 211 728 212 732
rect 206 727 212 728
rect 294 732 300 733
rect 294 728 295 732
rect 299 728 300 732
rect 294 727 300 728
rect 374 732 380 733
rect 374 728 375 732
rect 379 728 380 732
rect 374 727 380 728
rect 446 732 452 733
rect 446 728 447 732
rect 451 728 452 732
rect 446 727 452 728
rect 518 732 524 733
rect 518 728 519 732
rect 523 728 524 732
rect 518 727 524 728
rect 582 732 588 733
rect 582 728 583 732
rect 587 728 588 732
rect 582 727 588 728
rect 638 732 644 733
rect 638 728 639 732
rect 643 728 644 732
rect 638 727 644 728
rect 686 732 692 733
rect 686 728 687 732
rect 691 728 692 732
rect 686 727 692 728
rect 742 732 748 733
rect 742 728 743 732
rect 747 728 748 732
rect 742 727 748 728
rect 798 732 804 733
rect 798 728 799 732
rect 803 728 804 732
rect 798 727 804 728
rect 854 732 860 733
rect 854 728 855 732
rect 859 728 860 732
rect 854 727 860 728
rect 1134 728 1140 729
rect 1134 724 1135 728
rect 1139 724 1140 728
rect 1134 723 1140 724
rect 2118 728 2124 729
rect 2118 724 2119 728
rect 2123 724 2124 728
rect 2118 723 2124 724
rect 1158 720 1164 721
rect 1158 716 1159 720
rect 1163 716 1164 720
rect 1158 715 1164 716
rect 1198 720 1204 721
rect 1198 716 1199 720
rect 1203 716 1204 720
rect 1198 715 1204 716
rect 1238 720 1244 721
rect 1238 716 1239 720
rect 1243 716 1244 720
rect 1238 715 1244 716
rect 1286 720 1292 721
rect 1286 716 1287 720
rect 1291 716 1292 720
rect 1286 715 1292 716
rect 1358 720 1364 721
rect 1358 716 1359 720
rect 1363 716 1364 720
rect 1358 715 1364 716
rect 1438 720 1444 721
rect 1438 716 1439 720
rect 1443 716 1444 720
rect 1438 715 1444 716
rect 1526 720 1532 721
rect 1526 716 1527 720
rect 1531 716 1532 720
rect 1526 715 1532 716
rect 1614 720 1620 721
rect 1614 716 1615 720
rect 1619 716 1620 720
rect 1614 715 1620 716
rect 1710 720 1716 721
rect 1710 716 1711 720
rect 1715 716 1716 720
rect 1710 715 1716 716
rect 1806 720 1812 721
rect 1806 716 1807 720
rect 1811 716 1812 720
rect 1806 715 1812 716
rect 1902 720 1908 721
rect 1902 716 1903 720
rect 1907 716 1908 720
rect 1902 715 1908 716
rect 1998 720 2004 721
rect 1998 716 1999 720
rect 2003 716 2004 720
rect 1998 715 2004 716
rect 2070 720 2076 721
rect 2070 716 2071 720
rect 2075 716 2076 720
rect 2070 715 2076 716
rect 134 692 140 693
rect 134 688 135 692
rect 139 688 140 692
rect 134 687 140 688
rect 182 692 188 693
rect 182 688 183 692
rect 187 688 188 692
rect 182 687 188 688
rect 246 692 252 693
rect 246 688 247 692
rect 251 688 252 692
rect 246 687 252 688
rect 310 692 316 693
rect 310 688 311 692
rect 315 688 316 692
rect 310 687 316 688
rect 382 692 388 693
rect 382 688 383 692
rect 387 688 388 692
rect 382 687 388 688
rect 454 692 460 693
rect 454 688 455 692
rect 459 688 460 692
rect 454 687 460 688
rect 518 692 524 693
rect 518 688 519 692
rect 523 688 524 692
rect 518 687 524 688
rect 582 692 588 693
rect 582 688 583 692
rect 587 688 588 692
rect 582 687 588 688
rect 646 692 652 693
rect 646 688 647 692
rect 651 688 652 692
rect 646 687 652 688
rect 710 692 716 693
rect 710 688 711 692
rect 715 688 716 692
rect 710 687 716 688
rect 766 692 772 693
rect 766 688 767 692
rect 771 688 772 692
rect 766 687 772 688
rect 822 692 828 693
rect 822 688 823 692
rect 827 688 828 692
rect 822 687 828 688
rect 878 692 884 693
rect 878 688 879 692
rect 883 688 884 692
rect 878 687 884 688
rect 942 692 948 693
rect 942 688 943 692
rect 947 688 948 692
rect 942 687 948 688
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 110 679 116 680
rect 1094 684 1100 685
rect 1094 680 1095 684
rect 1099 680 1100 684
rect 1094 679 1100 680
rect 1238 680 1244 681
rect 1238 676 1239 680
rect 1243 676 1244 680
rect 1238 675 1244 676
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 1334 680 1340 681
rect 1334 676 1335 680
rect 1339 676 1340 680
rect 1334 675 1340 676
rect 1390 680 1396 681
rect 1390 676 1391 680
rect 1395 676 1396 680
rect 1390 675 1396 676
rect 1446 680 1452 681
rect 1446 676 1447 680
rect 1451 676 1452 680
rect 1446 675 1452 676
rect 1510 680 1516 681
rect 1510 676 1511 680
rect 1515 676 1516 680
rect 1510 675 1516 676
rect 1574 680 1580 681
rect 1574 676 1575 680
rect 1579 676 1580 680
rect 1574 675 1580 676
rect 1638 680 1644 681
rect 1638 676 1639 680
rect 1643 676 1644 680
rect 1638 675 1644 676
rect 1702 680 1708 681
rect 1702 676 1703 680
rect 1707 676 1708 680
rect 1702 675 1708 676
rect 1766 680 1772 681
rect 1766 676 1767 680
rect 1771 676 1772 680
rect 1766 675 1772 676
rect 1830 680 1836 681
rect 1830 676 1831 680
rect 1835 676 1836 680
rect 1830 675 1836 676
rect 1894 680 1900 681
rect 1894 676 1895 680
rect 1899 676 1900 680
rect 1894 675 1900 676
rect 1958 680 1964 681
rect 1958 676 1959 680
rect 1963 676 1964 680
rect 1958 675 1964 676
rect 2022 680 2028 681
rect 2022 676 2023 680
rect 2027 676 2028 680
rect 2022 675 2028 676
rect 2070 680 2076 681
rect 2070 676 2071 680
rect 2075 676 2076 680
rect 2070 675 2076 676
rect 1134 672 1140 673
rect 1134 668 1135 672
rect 1139 668 1140 672
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 1094 667 1100 668
rect 1134 667 1140 668
rect 2118 672 2124 673
rect 2118 668 2119 672
rect 2123 668 2124 672
rect 2118 667 2124 668
rect 110 662 116 663
rect 134 664 140 665
rect 134 660 135 664
rect 139 660 140 664
rect 134 659 140 660
rect 182 664 188 665
rect 182 660 183 664
rect 187 660 188 664
rect 182 659 188 660
rect 246 664 252 665
rect 246 660 247 664
rect 251 660 252 664
rect 246 659 252 660
rect 310 664 316 665
rect 310 660 311 664
rect 315 660 316 664
rect 310 659 316 660
rect 382 664 388 665
rect 382 660 383 664
rect 387 660 388 664
rect 382 659 388 660
rect 454 664 460 665
rect 454 660 455 664
rect 459 660 460 664
rect 454 659 460 660
rect 518 664 524 665
rect 518 660 519 664
rect 523 660 524 664
rect 518 659 524 660
rect 582 664 588 665
rect 582 660 583 664
rect 587 660 588 664
rect 582 659 588 660
rect 646 664 652 665
rect 646 660 647 664
rect 651 660 652 664
rect 646 659 652 660
rect 710 664 716 665
rect 710 660 711 664
rect 715 660 716 664
rect 710 659 716 660
rect 766 664 772 665
rect 766 660 767 664
rect 771 660 772 664
rect 766 659 772 660
rect 822 664 828 665
rect 822 660 823 664
rect 827 660 828 664
rect 822 659 828 660
rect 878 664 884 665
rect 878 660 879 664
rect 883 660 884 664
rect 878 659 884 660
rect 942 664 948 665
rect 942 660 943 664
rect 947 660 948 664
rect 1094 663 1095 667
rect 1099 663 1100 667
rect 1094 662 1100 663
rect 942 659 948 660
rect 1134 655 1140 656
rect 1134 651 1135 655
rect 1139 651 1140 655
rect 2118 655 2124 656
rect 1134 650 1140 651
rect 1238 652 1244 653
rect 1238 648 1239 652
rect 1243 648 1244 652
rect 1238 647 1244 648
rect 1286 652 1292 653
rect 1286 648 1287 652
rect 1291 648 1292 652
rect 1286 647 1292 648
rect 1334 652 1340 653
rect 1334 648 1335 652
rect 1339 648 1340 652
rect 1334 647 1340 648
rect 1390 652 1396 653
rect 1390 648 1391 652
rect 1395 648 1396 652
rect 1390 647 1396 648
rect 1446 652 1452 653
rect 1446 648 1447 652
rect 1451 648 1452 652
rect 1446 647 1452 648
rect 1510 652 1516 653
rect 1510 648 1511 652
rect 1515 648 1516 652
rect 1510 647 1516 648
rect 1574 652 1580 653
rect 1574 648 1575 652
rect 1579 648 1580 652
rect 1574 647 1580 648
rect 1638 652 1644 653
rect 1638 648 1639 652
rect 1643 648 1644 652
rect 1638 647 1644 648
rect 1702 652 1708 653
rect 1702 648 1703 652
rect 1707 648 1708 652
rect 1702 647 1708 648
rect 1766 652 1772 653
rect 1766 648 1767 652
rect 1771 648 1772 652
rect 1766 647 1772 648
rect 1830 652 1836 653
rect 1830 648 1831 652
rect 1835 648 1836 652
rect 1830 647 1836 648
rect 1894 652 1900 653
rect 1894 648 1895 652
rect 1899 648 1900 652
rect 1894 647 1900 648
rect 1958 652 1964 653
rect 1958 648 1959 652
rect 1963 648 1964 652
rect 1958 647 1964 648
rect 2022 652 2028 653
rect 2022 648 2023 652
rect 2027 648 2028 652
rect 2022 647 2028 648
rect 2070 652 2076 653
rect 2070 648 2071 652
rect 2075 648 2076 652
rect 2118 651 2119 655
rect 2123 651 2124 655
rect 2118 650 2124 651
rect 2070 647 2076 648
rect 158 644 164 645
rect 110 641 116 642
rect 110 637 111 641
rect 115 637 116 641
rect 158 640 159 644
rect 163 640 164 644
rect 158 639 164 640
rect 214 644 220 645
rect 214 640 215 644
rect 219 640 220 644
rect 214 639 220 640
rect 286 644 292 645
rect 286 640 287 644
rect 291 640 292 644
rect 286 639 292 640
rect 366 644 372 645
rect 366 640 367 644
rect 371 640 372 644
rect 366 639 372 640
rect 454 644 460 645
rect 454 640 455 644
rect 459 640 460 644
rect 454 639 460 640
rect 542 644 548 645
rect 542 640 543 644
rect 547 640 548 644
rect 542 639 548 640
rect 630 644 636 645
rect 630 640 631 644
rect 635 640 636 644
rect 630 639 636 640
rect 718 644 724 645
rect 718 640 719 644
rect 723 640 724 644
rect 718 639 724 640
rect 798 644 804 645
rect 798 640 799 644
rect 803 640 804 644
rect 798 639 804 640
rect 870 644 876 645
rect 870 640 871 644
rect 875 640 876 644
rect 870 639 876 640
rect 950 644 956 645
rect 950 640 951 644
rect 955 640 956 644
rect 950 639 956 640
rect 1030 644 1036 645
rect 1030 640 1031 644
rect 1035 640 1036 644
rect 1030 639 1036 640
rect 1094 641 1100 642
rect 110 636 116 637
rect 1094 637 1095 641
rect 1099 637 1100 641
rect 1278 640 1284 641
rect 1094 636 1100 637
rect 1134 637 1140 638
rect 1134 633 1135 637
rect 1139 633 1140 637
rect 1278 636 1279 640
rect 1283 636 1284 640
rect 1278 635 1284 636
rect 1318 640 1324 641
rect 1318 636 1319 640
rect 1323 636 1324 640
rect 1318 635 1324 636
rect 1366 640 1372 641
rect 1366 636 1367 640
rect 1371 636 1372 640
rect 1366 635 1372 636
rect 1422 640 1428 641
rect 1422 636 1423 640
rect 1427 636 1428 640
rect 1422 635 1428 636
rect 1478 640 1484 641
rect 1478 636 1479 640
rect 1483 636 1484 640
rect 1478 635 1484 636
rect 1534 640 1540 641
rect 1534 636 1535 640
rect 1539 636 1540 640
rect 1534 635 1540 636
rect 1590 640 1596 641
rect 1590 636 1591 640
rect 1595 636 1596 640
rect 1590 635 1596 636
rect 1646 640 1652 641
rect 1646 636 1647 640
rect 1651 636 1652 640
rect 1646 635 1652 636
rect 1718 640 1724 641
rect 1718 636 1719 640
rect 1723 636 1724 640
rect 1718 635 1724 636
rect 1798 640 1804 641
rect 1798 636 1799 640
rect 1803 636 1804 640
rect 1798 635 1804 636
rect 1878 640 1884 641
rect 1878 636 1879 640
rect 1883 636 1884 640
rect 1878 635 1884 636
rect 1966 640 1972 641
rect 1966 636 1967 640
rect 1971 636 1972 640
rect 1966 635 1972 636
rect 2062 640 2068 641
rect 2062 636 2063 640
rect 2067 636 2068 640
rect 2062 635 2068 636
rect 2118 637 2124 638
rect 1134 632 1140 633
rect 2118 633 2119 637
rect 2123 633 2124 637
rect 2118 632 2124 633
rect 110 624 116 625
rect 110 620 111 624
rect 115 620 116 624
rect 110 619 116 620
rect 1094 624 1100 625
rect 1094 620 1095 624
rect 1099 620 1100 624
rect 1094 619 1100 620
rect 1134 620 1140 621
rect 158 616 164 617
rect 158 612 159 616
rect 163 612 164 616
rect 158 611 164 612
rect 214 616 220 617
rect 214 612 215 616
rect 219 612 220 616
rect 214 611 220 612
rect 286 616 292 617
rect 286 612 287 616
rect 291 612 292 616
rect 286 611 292 612
rect 366 616 372 617
rect 366 612 367 616
rect 371 612 372 616
rect 366 611 372 612
rect 454 616 460 617
rect 454 612 455 616
rect 459 612 460 616
rect 454 611 460 612
rect 542 616 548 617
rect 542 612 543 616
rect 547 612 548 616
rect 542 611 548 612
rect 630 616 636 617
rect 630 612 631 616
rect 635 612 636 616
rect 630 611 636 612
rect 718 616 724 617
rect 718 612 719 616
rect 723 612 724 616
rect 718 611 724 612
rect 798 616 804 617
rect 798 612 799 616
rect 803 612 804 616
rect 798 611 804 612
rect 870 616 876 617
rect 870 612 871 616
rect 875 612 876 616
rect 870 611 876 612
rect 950 616 956 617
rect 950 612 951 616
rect 955 612 956 616
rect 950 611 956 612
rect 1030 616 1036 617
rect 1030 612 1031 616
rect 1035 612 1036 616
rect 1134 616 1135 620
rect 1139 616 1140 620
rect 1134 615 1140 616
rect 2118 620 2124 621
rect 2118 616 2119 620
rect 2123 616 2124 620
rect 2118 615 2124 616
rect 1030 611 1036 612
rect 1278 612 1284 613
rect 1278 608 1279 612
rect 1283 608 1284 612
rect 1278 607 1284 608
rect 1318 612 1324 613
rect 1318 608 1319 612
rect 1323 608 1324 612
rect 1318 607 1324 608
rect 1366 612 1372 613
rect 1366 608 1367 612
rect 1371 608 1372 612
rect 1366 607 1372 608
rect 1422 612 1428 613
rect 1422 608 1423 612
rect 1427 608 1428 612
rect 1422 607 1428 608
rect 1478 612 1484 613
rect 1478 608 1479 612
rect 1483 608 1484 612
rect 1478 607 1484 608
rect 1534 612 1540 613
rect 1534 608 1535 612
rect 1539 608 1540 612
rect 1534 607 1540 608
rect 1590 612 1596 613
rect 1590 608 1591 612
rect 1595 608 1596 612
rect 1590 607 1596 608
rect 1646 612 1652 613
rect 1646 608 1647 612
rect 1651 608 1652 612
rect 1646 607 1652 608
rect 1718 612 1724 613
rect 1718 608 1719 612
rect 1723 608 1724 612
rect 1718 607 1724 608
rect 1798 612 1804 613
rect 1798 608 1799 612
rect 1803 608 1804 612
rect 1798 607 1804 608
rect 1878 612 1884 613
rect 1878 608 1879 612
rect 1883 608 1884 612
rect 1878 607 1884 608
rect 1966 612 1972 613
rect 1966 608 1967 612
rect 1971 608 1972 612
rect 1966 607 1972 608
rect 2062 612 2068 613
rect 2062 608 2063 612
rect 2067 608 2068 612
rect 2062 607 2068 608
rect 158 576 164 577
rect 158 572 159 576
rect 163 572 164 576
rect 158 571 164 572
rect 206 576 212 577
rect 206 572 207 576
rect 211 572 212 576
rect 206 571 212 572
rect 254 576 260 577
rect 254 572 255 576
rect 259 572 260 576
rect 254 571 260 572
rect 310 576 316 577
rect 310 572 311 576
rect 315 572 316 576
rect 310 571 316 572
rect 382 576 388 577
rect 382 572 383 576
rect 387 572 388 576
rect 382 571 388 572
rect 462 576 468 577
rect 462 572 463 576
rect 467 572 468 576
rect 462 571 468 572
rect 542 576 548 577
rect 542 572 543 576
rect 547 572 548 576
rect 542 571 548 572
rect 622 576 628 577
rect 622 572 623 576
rect 627 572 628 576
rect 622 571 628 572
rect 702 576 708 577
rect 702 572 703 576
rect 707 572 708 576
rect 702 571 708 572
rect 782 576 788 577
rect 782 572 783 576
rect 787 572 788 576
rect 782 571 788 572
rect 854 576 860 577
rect 854 572 855 576
rect 859 572 860 576
rect 854 571 860 572
rect 926 576 932 577
rect 926 572 927 576
rect 931 572 932 576
rect 926 571 932 572
rect 998 576 1004 577
rect 998 572 999 576
rect 1003 572 1004 576
rect 998 571 1004 572
rect 1046 576 1052 577
rect 1046 572 1047 576
rect 1051 572 1052 576
rect 1046 571 1052 572
rect 1334 576 1340 577
rect 1334 572 1335 576
rect 1339 572 1340 576
rect 1334 571 1340 572
rect 1374 576 1380 577
rect 1374 572 1375 576
rect 1379 572 1380 576
rect 1374 571 1380 572
rect 1414 576 1420 577
rect 1414 572 1415 576
rect 1419 572 1420 576
rect 1414 571 1420 572
rect 1462 576 1468 577
rect 1462 572 1463 576
rect 1467 572 1468 576
rect 1462 571 1468 572
rect 1518 576 1524 577
rect 1518 572 1519 576
rect 1523 572 1524 576
rect 1518 571 1524 572
rect 1582 576 1588 577
rect 1582 572 1583 576
rect 1587 572 1588 576
rect 1582 571 1588 572
rect 1654 576 1660 577
rect 1654 572 1655 576
rect 1659 572 1660 576
rect 1654 571 1660 572
rect 1726 576 1732 577
rect 1726 572 1727 576
rect 1731 572 1732 576
rect 1726 571 1732 572
rect 1806 576 1812 577
rect 1806 572 1807 576
rect 1811 572 1812 576
rect 1806 571 1812 572
rect 1886 576 1892 577
rect 1886 572 1887 576
rect 1891 572 1892 576
rect 1886 571 1892 572
rect 1974 576 1980 577
rect 1974 572 1975 576
rect 1979 572 1980 576
rect 1974 571 1980 572
rect 2062 576 2068 577
rect 2062 572 2063 576
rect 2067 572 2068 576
rect 2062 571 2068 572
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 110 563 116 564
rect 1094 568 1100 569
rect 1094 564 1095 568
rect 1099 564 1100 568
rect 1094 563 1100 564
rect 1134 568 1140 569
rect 1134 564 1135 568
rect 1139 564 1140 568
rect 1134 563 1140 564
rect 2118 568 2124 569
rect 2118 564 2119 568
rect 2123 564 2124 568
rect 2118 563 2124 564
rect 110 551 116 552
rect 110 547 111 551
rect 115 547 116 551
rect 1094 551 1100 552
rect 110 546 116 547
rect 158 548 164 549
rect 158 544 159 548
rect 163 544 164 548
rect 158 543 164 544
rect 206 548 212 549
rect 206 544 207 548
rect 211 544 212 548
rect 206 543 212 544
rect 254 548 260 549
rect 254 544 255 548
rect 259 544 260 548
rect 254 543 260 544
rect 310 548 316 549
rect 310 544 311 548
rect 315 544 316 548
rect 310 543 316 544
rect 382 548 388 549
rect 382 544 383 548
rect 387 544 388 548
rect 382 543 388 544
rect 462 548 468 549
rect 462 544 463 548
rect 467 544 468 548
rect 462 543 468 544
rect 542 548 548 549
rect 542 544 543 548
rect 547 544 548 548
rect 542 543 548 544
rect 622 548 628 549
rect 622 544 623 548
rect 627 544 628 548
rect 622 543 628 544
rect 702 548 708 549
rect 702 544 703 548
rect 707 544 708 548
rect 702 543 708 544
rect 782 548 788 549
rect 782 544 783 548
rect 787 544 788 548
rect 782 543 788 544
rect 854 548 860 549
rect 854 544 855 548
rect 859 544 860 548
rect 854 543 860 544
rect 926 548 932 549
rect 926 544 927 548
rect 931 544 932 548
rect 926 543 932 544
rect 998 548 1004 549
rect 998 544 999 548
rect 1003 544 1004 548
rect 998 543 1004 544
rect 1046 548 1052 549
rect 1046 544 1047 548
rect 1051 544 1052 548
rect 1094 547 1095 551
rect 1099 547 1100 551
rect 1094 546 1100 547
rect 1134 551 1140 552
rect 1134 547 1135 551
rect 1139 547 1140 551
rect 2118 551 2124 552
rect 1134 546 1140 547
rect 1334 548 1340 549
rect 1046 543 1052 544
rect 1334 544 1335 548
rect 1339 544 1340 548
rect 1334 543 1340 544
rect 1374 548 1380 549
rect 1374 544 1375 548
rect 1379 544 1380 548
rect 1374 543 1380 544
rect 1414 548 1420 549
rect 1414 544 1415 548
rect 1419 544 1420 548
rect 1414 543 1420 544
rect 1462 548 1468 549
rect 1462 544 1463 548
rect 1467 544 1468 548
rect 1462 543 1468 544
rect 1518 548 1524 549
rect 1518 544 1519 548
rect 1523 544 1524 548
rect 1518 543 1524 544
rect 1582 548 1588 549
rect 1582 544 1583 548
rect 1587 544 1588 548
rect 1582 543 1588 544
rect 1654 548 1660 549
rect 1654 544 1655 548
rect 1659 544 1660 548
rect 1654 543 1660 544
rect 1726 548 1732 549
rect 1726 544 1727 548
rect 1731 544 1732 548
rect 1726 543 1732 544
rect 1806 548 1812 549
rect 1806 544 1807 548
rect 1811 544 1812 548
rect 1806 543 1812 544
rect 1886 548 1892 549
rect 1886 544 1887 548
rect 1891 544 1892 548
rect 1886 543 1892 544
rect 1974 548 1980 549
rect 1974 544 1975 548
rect 1979 544 1980 548
rect 1974 543 1980 544
rect 2062 548 2068 549
rect 2062 544 2063 548
rect 2067 544 2068 548
rect 2118 547 2119 551
rect 2123 547 2124 551
rect 2118 546 2124 547
rect 2062 543 2068 544
rect 1190 532 1196 533
rect 1134 529 1140 530
rect 166 528 172 529
rect 110 525 116 526
rect 110 521 111 525
rect 115 521 116 525
rect 166 524 167 528
rect 171 524 172 528
rect 166 523 172 524
rect 222 528 228 529
rect 222 524 223 528
rect 227 524 228 528
rect 222 523 228 524
rect 286 528 292 529
rect 286 524 287 528
rect 291 524 292 528
rect 286 523 292 524
rect 358 528 364 529
rect 358 524 359 528
rect 363 524 364 528
rect 358 523 364 524
rect 430 528 436 529
rect 430 524 431 528
rect 435 524 436 528
rect 430 523 436 524
rect 510 528 516 529
rect 510 524 511 528
rect 515 524 516 528
rect 510 523 516 524
rect 590 528 596 529
rect 590 524 591 528
rect 595 524 596 528
rect 590 523 596 524
rect 662 528 668 529
rect 662 524 663 528
rect 667 524 668 528
rect 662 523 668 524
rect 734 528 740 529
rect 734 524 735 528
rect 739 524 740 528
rect 734 523 740 524
rect 806 528 812 529
rect 806 524 807 528
rect 811 524 812 528
rect 806 523 812 524
rect 870 528 876 529
rect 870 524 871 528
rect 875 524 876 528
rect 870 523 876 524
rect 934 528 940 529
rect 934 524 935 528
rect 939 524 940 528
rect 934 523 940 524
rect 998 528 1004 529
rect 998 524 999 528
rect 1003 524 1004 528
rect 998 523 1004 524
rect 1046 528 1052 529
rect 1046 524 1047 528
rect 1051 524 1052 528
rect 1046 523 1052 524
rect 1094 525 1100 526
rect 110 520 116 521
rect 1094 521 1095 525
rect 1099 521 1100 525
rect 1134 525 1135 529
rect 1139 525 1140 529
rect 1190 528 1191 532
rect 1195 528 1196 532
rect 1190 527 1196 528
rect 1238 532 1244 533
rect 1238 528 1239 532
rect 1243 528 1244 532
rect 1238 527 1244 528
rect 1286 532 1292 533
rect 1286 528 1287 532
rect 1291 528 1292 532
rect 1286 527 1292 528
rect 1342 532 1348 533
rect 1342 528 1343 532
rect 1347 528 1348 532
rect 1342 527 1348 528
rect 1406 532 1412 533
rect 1406 528 1407 532
rect 1411 528 1412 532
rect 1406 527 1412 528
rect 1478 532 1484 533
rect 1478 528 1479 532
rect 1483 528 1484 532
rect 1478 527 1484 528
rect 1542 532 1548 533
rect 1542 528 1543 532
rect 1547 528 1548 532
rect 1542 527 1548 528
rect 1606 532 1612 533
rect 1606 528 1607 532
rect 1611 528 1612 532
rect 1606 527 1612 528
rect 1670 532 1676 533
rect 1670 528 1671 532
rect 1675 528 1676 532
rect 1670 527 1676 528
rect 1734 532 1740 533
rect 1734 528 1735 532
rect 1739 528 1740 532
rect 1734 527 1740 528
rect 1798 532 1804 533
rect 1798 528 1799 532
rect 1803 528 1804 532
rect 1798 527 1804 528
rect 1862 532 1868 533
rect 1862 528 1863 532
rect 1867 528 1868 532
rect 1862 527 1868 528
rect 1934 532 1940 533
rect 1934 528 1935 532
rect 1939 528 1940 532
rect 1934 527 1940 528
rect 2006 532 2012 533
rect 2006 528 2007 532
rect 2011 528 2012 532
rect 2006 527 2012 528
rect 2070 532 2076 533
rect 2070 528 2071 532
rect 2075 528 2076 532
rect 2070 527 2076 528
rect 2118 529 2124 530
rect 1134 524 1140 525
rect 2118 525 2119 529
rect 2123 525 2124 529
rect 2118 524 2124 525
rect 1094 520 1100 521
rect 1134 512 1140 513
rect 110 508 116 509
rect 110 504 111 508
rect 115 504 116 508
rect 110 503 116 504
rect 1094 508 1100 509
rect 1094 504 1095 508
rect 1099 504 1100 508
rect 1134 508 1135 512
rect 1139 508 1140 512
rect 1134 507 1140 508
rect 2118 512 2124 513
rect 2118 508 2119 512
rect 2123 508 2124 512
rect 2118 507 2124 508
rect 1094 503 1100 504
rect 1190 504 1196 505
rect 166 500 172 501
rect 166 496 167 500
rect 171 496 172 500
rect 166 495 172 496
rect 222 500 228 501
rect 222 496 223 500
rect 227 496 228 500
rect 222 495 228 496
rect 286 500 292 501
rect 286 496 287 500
rect 291 496 292 500
rect 286 495 292 496
rect 358 500 364 501
rect 358 496 359 500
rect 363 496 364 500
rect 358 495 364 496
rect 430 500 436 501
rect 430 496 431 500
rect 435 496 436 500
rect 430 495 436 496
rect 510 500 516 501
rect 510 496 511 500
rect 515 496 516 500
rect 510 495 516 496
rect 590 500 596 501
rect 590 496 591 500
rect 595 496 596 500
rect 590 495 596 496
rect 662 500 668 501
rect 662 496 663 500
rect 667 496 668 500
rect 662 495 668 496
rect 734 500 740 501
rect 734 496 735 500
rect 739 496 740 500
rect 734 495 740 496
rect 806 500 812 501
rect 806 496 807 500
rect 811 496 812 500
rect 806 495 812 496
rect 870 500 876 501
rect 870 496 871 500
rect 875 496 876 500
rect 870 495 876 496
rect 934 500 940 501
rect 934 496 935 500
rect 939 496 940 500
rect 934 495 940 496
rect 998 500 1004 501
rect 998 496 999 500
rect 1003 496 1004 500
rect 998 495 1004 496
rect 1046 500 1052 501
rect 1046 496 1047 500
rect 1051 496 1052 500
rect 1190 500 1191 504
rect 1195 500 1196 504
rect 1190 499 1196 500
rect 1238 504 1244 505
rect 1238 500 1239 504
rect 1243 500 1244 504
rect 1238 499 1244 500
rect 1286 504 1292 505
rect 1286 500 1287 504
rect 1291 500 1292 504
rect 1286 499 1292 500
rect 1342 504 1348 505
rect 1342 500 1343 504
rect 1347 500 1348 504
rect 1342 499 1348 500
rect 1406 504 1412 505
rect 1406 500 1407 504
rect 1411 500 1412 504
rect 1406 499 1412 500
rect 1478 504 1484 505
rect 1478 500 1479 504
rect 1483 500 1484 504
rect 1478 499 1484 500
rect 1542 504 1548 505
rect 1542 500 1543 504
rect 1547 500 1548 504
rect 1542 499 1548 500
rect 1606 504 1612 505
rect 1606 500 1607 504
rect 1611 500 1612 504
rect 1606 499 1612 500
rect 1670 504 1676 505
rect 1670 500 1671 504
rect 1675 500 1676 504
rect 1670 499 1676 500
rect 1734 504 1740 505
rect 1734 500 1735 504
rect 1739 500 1740 504
rect 1734 499 1740 500
rect 1798 504 1804 505
rect 1798 500 1799 504
rect 1803 500 1804 504
rect 1798 499 1804 500
rect 1862 504 1868 505
rect 1862 500 1863 504
rect 1867 500 1868 504
rect 1862 499 1868 500
rect 1934 504 1940 505
rect 1934 500 1935 504
rect 1939 500 1940 504
rect 1934 499 1940 500
rect 2006 504 2012 505
rect 2006 500 2007 504
rect 2011 500 2012 504
rect 2006 499 2012 500
rect 2070 504 2076 505
rect 2070 500 2071 504
rect 2075 500 2076 504
rect 2070 499 2076 500
rect 1046 495 1052 496
rect 1158 468 1164 469
rect 166 464 172 465
rect 166 460 167 464
rect 171 460 172 464
rect 166 459 172 460
rect 230 464 236 465
rect 230 460 231 464
rect 235 460 236 464
rect 230 459 236 460
rect 302 464 308 465
rect 302 460 303 464
rect 307 460 308 464
rect 302 459 308 460
rect 374 464 380 465
rect 374 460 375 464
rect 379 460 380 464
rect 374 459 380 460
rect 454 464 460 465
rect 454 460 455 464
rect 459 460 460 464
rect 454 459 460 460
rect 534 464 540 465
rect 534 460 535 464
rect 539 460 540 464
rect 534 459 540 460
rect 606 464 612 465
rect 606 460 607 464
rect 611 460 612 464
rect 606 459 612 460
rect 678 464 684 465
rect 678 460 679 464
rect 683 460 684 464
rect 678 459 684 460
rect 742 464 748 465
rect 742 460 743 464
rect 747 460 748 464
rect 742 459 748 460
rect 798 464 804 465
rect 798 460 799 464
rect 803 460 804 464
rect 798 459 804 460
rect 854 464 860 465
rect 854 460 855 464
rect 859 460 860 464
rect 854 459 860 460
rect 902 464 908 465
rect 902 460 903 464
rect 907 460 908 464
rect 902 459 908 460
rect 958 464 964 465
rect 958 460 959 464
rect 963 460 964 464
rect 958 459 964 460
rect 1006 464 1012 465
rect 1006 460 1007 464
rect 1011 460 1012 464
rect 1006 459 1012 460
rect 1046 464 1052 465
rect 1046 460 1047 464
rect 1051 460 1052 464
rect 1158 464 1159 468
rect 1163 464 1164 468
rect 1158 463 1164 464
rect 1262 468 1268 469
rect 1262 464 1263 468
rect 1267 464 1268 468
rect 1262 463 1268 464
rect 1382 468 1388 469
rect 1382 464 1383 468
rect 1387 464 1388 468
rect 1382 463 1388 464
rect 1494 468 1500 469
rect 1494 464 1495 468
rect 1499 464 1500 468
rect 1494 463 1500 464
rect 1598 468 1604 469
rect 1598 464 1599 468
rect 1603 464 1604 468
rect 1598 463 1604 464
rect 1702 468 1708 469
rect 1702 464 1703 468
rect 1707 464 1708 468
rect 1702 463 1708 464
rect 1798 468 1804 469
rect 1798 464 1799 468
rect 1803 464 1804 468
rect 1798 463 1804 464
rect 1886 468 1892 469
rect 1886 464 1887 468
rect 1891 464 1892 468
rect 1886 463 1892 464
rect 1982 468 1988 469
rect 1982 464 1983 468
rect 1987 464 1988 468
rect 1982 463 1988 464
rect 2070 468 2076 469
rect 2070 464 2071 468
rect 2075 464 2076 468
rect 2070 463 2076 464
rect 1046 459 1052 460
rect 1134 460 1140 461
rect 110 456 116 457
rect 110 452 111 456
rect 115 452 116 456
rect 110 451 116 452
rect 1094 456 1100 457
rect 1094 452 1095 456
rect 1099 452 1100 456
rect 1134 456 1135 460
rect 1139 456 1140 460
rect 1134 455 1140 456
rect 2118 460 2124 461
rect 2118 456 2119 460
rect 2123 456 2124 460
rect 2118 455 2124 456
rect 1094 451 1100 452
rect 1134 443 1140 444
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 1094 439 1100 440
rect 110 434 116 435
rect 166 436 172 437
rect 166 432 167 436
rect 171 432 172 436
rect 166 431 172 432
rect 230 436 236 437
rect 230 432 231 436
rect 235 432 236 436
rect 230 431 236 432
rect 302 436 308 437
rect 302 432 303 436
rect 307 432 308 436
rect 302 431 308 432
rect 374 436 380 437
rect 374 432 375 436
rect 379 432 380 436
rect 374 431 380 432
rect 454 436 460 437
rect 454 432 455 436
rect 459 432 460 436
rect 454 431 460 432
rect 534 436 540 437
rect 534 432 535 436
rect 539 432 540 436
rect 534 431 540 432
rect 606 436 612 437
rect 606 432 607 436
rect 611 432 612 436
rect 606 431 612 432
rect 678 436 684 437
rect 678 432 679 436
rect 683 432 684 436
rect 678 431 684 432
rect 742 436 748 437
rect 742 432 743 436
rect 747 432 748 436
rect 742 431 748 432
rect 798 436 804 437
rect 798 432 799 436
rect 803 432 804 436
rect 798 431 804 432
rect 854 436 860 437
rect 854 432 855 436
rect 859 432 860 436
rect 854 431 860 432
rect 902 436 908 437
rect 902 432 903 436
rect 907 432 908 436
rect 902 431 908 432
rect 958 436 964 437
rect 958 432 959 436
rect 963 432 964 436
rect 958 431 964 432
rect 1006 436 1012 437
rect 1006 432 1007 436
rect 1011 432 1012 436
rect 1006 431 1012 432
rect 1046 436 1052 437
rect 1046 432 1047 436
rect 1051 432 1052 436
rect 1094 435 1095 439
rect 1099 435 1100 439
rect 1134 439 1135 443
rect 1139 439 1140 443
rect 2118 443 2124 444
rect 1134 438 1140 439
rect 1158 440 1164 441
rect 1158 436 1159 440
rect 1163 436 1164 440
rect 1158 435 1164 436
rect 1262 440 1268 441
rect 1262 436 1263 440
rect 1267 436 1268 440
rect 1262 435 1268 436
rect 1382 440 1388 441
rect 1382 436 1383 440
rect 1387 436 1388 440
rect 1382 435 1388 436
rect 1494 440 1500 441
rect 1494 436 1495 440
rect 1499 436 1500 440
rect 1494 435 1500 436
rect 1598 440 1604 441
rect 1598 436 1599 440
rect 1603 436 1604 440
rect 1598 435 1604 436
rect 1702 440 1708 441
rect 1702 436 1703 440
rect 1707 436 1708 440
rect 1702 435 1708 436
rect 1798 440 1804 441
rect 1798 436 1799 440
rect 1803 436 1804 440
rect 1798 435 1804 436
rect 1886 440 1892 441
rect 1886 436 1887 440
rect 1891 436 1892 440
rect 1886 435 1892 436
rect 1982 440 1988 441
rect 1982 436 1983 440
rect 1987 436 1988 440
rect 1982 435 1988 436
rect 2070 440 2076 441
rect 2070 436 2071 440
rect 2075 436 2076 440
rect 2118 439 2119 443
rect 2123 439 2124 443
rect 2118 438 2124 439
rect 2070 435 2076 436
rect 1094 434 1100 435
rect 1046 431 1052 432
rect 1158 428 1164 429
rect 1134 425 1140 426
rect 150 424 156 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 150 420 151 424
rect 155 420 156 424
rect 150 419 156 420
rect 214 424 220 425
rect 214 420 215 424
rect 219 420 220 424
rect 214 419 220 420
rect 278 424 284 425
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 350 424 356 425
rect 350 420 351 424
rect 355 420 356 424
rect 350 419 356 420
rect 422 424 428 425
rect 422 420 423 424
rect 427 420 428 424
rect 422 419 428 420
rect 486 424 492 425
rect 486 420 487 424
rect 491 420 492 424
rect 486 419 492 420
rect 550 424 556 425
rect 550 420 551 424
rect 555 420 556 424
rect 550 419 556 420
rect 614 424 620 425
rect 614 420 615 424
rect 619 420 620 424
rect 614 419 620 420
rect 670 424 676 425
rect 670 420 671 424
rect 675 420 676 424
rect 670 419 676 420
rect 726 424 732 425
rect 726 420 727 424
rect 731 420 732 424
rect 726 419 732 420
rect 790 424 796 425
rect 790 420 791 424
rect 795 420 796 424
rect 790 419 796 420
rect 854 424 860 425
rect 854 420 855 424
rect 859 420 860 424
rect 854 419 860 420
rect 1094 421 1100 422
rect 110 416 116 417
rect 1094 417 1095 421
rect 1099 417 1100 421
rect 1134 421 1135 425
rect 1139 421 1140 425
rect 1158 424 1159 428
rect 1163 424 1164 428
rect 1158 423 1164 424
rect 1198 428 1204 429
rect 1198 424 1199 428
rect 1203 424 1204 428
rect 1198 423 1204 424
rect 1254 428 1260 429
rect 1254 424 1255 428
rect 1259 424 1260 428
rect 1254 423 1260 424
rect 1334 428 1340 429
rect 1334 424 1335 428
rect 1339 424 1340 428
rect 1334 423 1340 424
rect 1414 428 1420 429
rect 1414 424 1415 428
rect 1419 424 1420 428
rect 1414 423 1420 424
rect 1502 428 1508 429
rect 1502 424 1503 428
rect 1507 424 1508 428
rect 1502 423 1508 424
rect 1590 428 1596 429
rect 1590 424 1591 428
rect 1595 424 1596 428
rect 1590 423 1596 424
rect 1670 428 1676 429
rect 1670 424 1671 428
rect 1675 424 1676 428
rect 1670 423 1676 424
rect 1750 428 1756 429
rect 1750 424 1751 428
rect 1755 424 1756 428
rect 1750 423 1756 424
rect 1822 428 1828 429
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1822 423 1828 424
rect 1886 428 1892 429
rect 1886 424 1887 428
rect 1891 424 1892 428
rect 1886 423 1892 424
rect 1950 428 1956 429
rect 1950 424 1951 428
rect 1955 424 1956 428
rect 1950 423 1956 424
rect 2022 428 2028 429
rect 2022 424 2023 428
rect 2027 424 2028 428
rect 2022 423 2028 424
rect 2070 428 2076 429
rect 2070 424 2071 428
rect 2075 424 2076 428
rect 2070 423 2076 424
rect 2118 425 2124 426
rect 1134 420 1140 421
rect 2118 421 2119 425
rect 2123 421 2124 425
rect 2118 420 2124 421
rect 1094 416 1100 417
rect 1134 408 1140 409
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 1094 404 1100 405
rect 1094 400 1095 404
rect 1099 400 1100 404
rect 1134 404 1135 408
rect 1139 404 1140 408
rect 1134 403 1140 404
rect 2118 408 2124 409
rect 2118 404 2119 408
rect 2123 404 2124 408
rect 2118 403 2124 404
rect 1094 399 1100 400
rect 1158 400 1164 401
rect 150 396 156 397
rect 150 392 151 396
rect 155 392 156 396
rect 150 391 156 392
rect 214 396 220 397
rect 214 392 215 396
rect 219 392 220 396
rect 214 391 220 392
rect 278 396 284 397
rect 278 392 279 396
rect 283 392 284 396
rect 278 391 284 392
rect 350 396 356 397
rect 350 392 351 396
rect 355 392 356 396
rect 350 391 356 392
rect 422 396 428 397
rect 422 392 423 396
rect 427 392 428 396
rect 422 391 428 392
rect 486 396 492 397
rect 486 392 487 396
rect 491 392 492 396
rect 486 391 492 392
rect 550 396 556 397
rect 550 392 551 396
rect 555 392 556 396
rect 550 391 556 392
rect 614 396 620 397
rect 614 392 615 396
rect 619 392 620 396
rect 614 391 620 392
rect 670 396 676 397
rect 670 392 671 396
rect 675 392 676 396
rect 670 391 676 392
rect 726 396 732 397
rect 726 392 727 396
rect 731 392 732 396
rect 726 391 732 392
rect 790 396 796 397
rect 790 392 791 396
rect 795 392 796 396
rect 790 391 796 392
rect 854 396 860 397
rect 854 392 855 396
rect 859 392 860 396
rect 1158 396 1159 400
rect 1163 396 1164 400
rect 1158 395 1164 396
rect 1198 400 1204 401
rect 1198 396 1199 400
rect 1203 396 1204 400
rect 1198 395 1204 396
rect 1254 400 1260 401
rect 1254 396 1255 400
rect 1259 396 1260 400
rect 1254 395 1260 396
rect 1334 400 1340 401
rect 1334 396 1335 400
rect 1339 396 1340 400
rect 1334 395 1340 396
rect 1414 400 1420 401
rect 1414 396 1415 400
rect 1419 396 1420 400
rect 1414 395 1420 396
rect 1502 400 1508 401
rect 1502 396 1503 400
rect 1507 396 1508 400
rect 1502 395 1508 396
rect 1590 400 1596 401
rect 1590 396 1591 400
rect 1595 396 1596 400
rect 1590 395 1596 396
rect 1670 400 1676 401
rect 1670 396 1671 400
rect 1675 396 1676 400
rect 1670 395 1676 396
rect 1750 400 1756 401
rect 1750 396 1751 400
rect 1755 396 1756 400
rect 1750 395 1756 396
rect 1822 400 1828 401
rect 1822 396 1823 400
rect 1827 396 1828 400
rect 1822 395 1828 396
rect 1886 400 1892 401
rect 1886 396 1887 400
rect 1891 396 1892 400
rect 1886 395 1892 396
rect 1950 400 1956 401
rect 1950 396 1951 400
rect 1955 396 1956 400
rect 1950 395 1956 396
rect 2022 400 2028 401
rect 2022 396 2023 400
rect 2027 396 2028 400
rect 2022 395 2028 396
rect 2070 400 2076 401
rect 2070 396 2071 400
rect 2075 396 2076 400
rect 2070 395 2076 396
rect 854 391 860 392
rect 134 360 140 361
rect 134 356 135 360
rect 139 356 140 360
rect 134 355 140 356
rect 174 360 180 361
rect 174 356 175 360
rect 179 356 180 360
rect 174 355 180 356
rect 214 360 220 361
rect 214 356 215 360
rect 219 356 220 360
rect 214 355 220 356
rect 270 360 276 361
rect 270 356 271 360
rect 275 356 276 360
rect 270 355 276 356
rect 334 360 340 361
rect 334 356 335 360
rect 339 356 340 360
rect 334 355 340 356
rect 398 360 404 361
rect 398 356 399 360
rect 403 356 404 360
rect 398 355 404 356
rect 462 360 468 361
rect 462 356 463 360
rect 467 356 468 360
rect 462 355 468 356
rect 518 360 524 361
rect 518 356 519 360
rect 523 356 524 360
rect 518 355 524 356
rect 574 360 580 361
rect 574 356 575 360
rect 579 356 580 360
rect 574 355 580 356
rect 630 360 636 361
rect 630 356 631 360
rect 635 356 636 360
rect 630 355 636 356
rect 686 360 692 361
rect 686 356 687 360
rect 691 356 692 360
rect 686 355 692 356
rect 750 360 756 361
rect 750 356 751 360
rect 755 356 756 360
rect 750 355 756 356
rect 1302 360 1308 361
rect 1302 356 1303 360
rect 1307 356 1308 360
rect 1302 355 1308 356
rect 1342 360 1348 361
rect 1342 356 1343 360
rect 1347 356 1348 360
rect 1342 355 1348 356
rect 1382 360 1388 361
rect 1382 356 1383 360
rect 1387 356 1388 360
rect 1382 355 1388 356
rect 1422 360 1428 361
rect 1422 356 1423 360
rect 1427 356 1428 360
rect 1422 355 1428 356
rect 1462 360 1468 361
rect 1462 356 1463 360
rect 1467 356 1468 360
rect 1462 355 1468 356
rect 1502 360 1508 361
rect 1502 356 1503 360
rect 1507 356 1508 360
rect 1502 355 1508 356
rect 1550 360 1556 361
rect 1550 356 1551 360
rect 1555 356 1556 360
rect 1550 355 1556 356
rect 1614 360 1620 361
rect 1614 356 1615 360
rect 1619 356 1620 360
rect 1614 355 1620 356
rect 1678 360 1684 361
rect 1678 356 1679 360
rect 1683 356 1684 360
rect 1678 355 1684 356
rect 1750 360 1756 361
rect 1750 356 1751 360
rect 1755 356 1756 360
rect 1750 355 1756 356
rect 1830 360 1836 361
rect 1830 356 1831 360
rect 1835 356 1836 360
rect 1830 355 1836 356
rect 1918 360 1924 361
rect 1918 356 1919 360
rect 1923 356 1924 360
rect 1918 355 1924 356
rect 2006 360 2012 361
rect 2006 356 2007 360
rect 2011 356 2012 360
rect 2006 355 2012 356
rect 2070 360 2076 361
rect 2070 356 2071 360
rect 2075 356 2076 360
rect 2070 355 2076 356
rect 110 352 116 353
rect 110 348 111 352
rect 115 348 116 352
rect 110 347 116 348
rect 1094 352 1100 353
rect 1094 348 1095 352
rect 1099 348 1100 352
rect 1094 347 1100 348
rect 1134 352 1140 353
rect 1134 348 1135 352
rect 1139 348 1140 352
rect 1134 347 1140 348
rect 2118 352 2124 353
rect 2118 348 2119 352
rect 2123 348 2124 352
rect 2118 347 2124 348
rect 110 335 116 336
rect 110 331 111 335
rect 115 331 116 335
rect 1094 335 1100 336
rect 110 330 116 331
rect 134 332 140 333
rect 134 328 135 332
rect 139 328 140 332
rect 134 327 140 328
rect 174 332 180 333
rect 174 328 175 332
rect 179 328 180 332
rect 174 327 180 328
rect 214 332 220 333
rect 214 328 215 332
rect 219 328 220 332
rect 214 327 220 328
rect 270 332 276 333
rect 270 328 271 332
rect 275 328 276 332
rect 270 327 276 328
rect 334 332 340 333
rect 334 328 335 332
rect 339 328 340 332
rect 334 327 340 328
rect 398 332 404 333
rect 398 328 399 332
rect 403 328 404 332
rect 398 327 404 328
rect 462 332 468 333
rect 462 328 463 332
rect 467 328 468 332
rect 462 327 468 328
rect 518 332 524 333
rect 518 328 519 332
rect 523 328 524 332
rect 518 327 524 328
rect 574 332 580 333
rect 574 328 575 332
rect 579 328 580 332
rect 574 327 580 328
rect 630 332 636 333
rect 630 328 631 332
rect 635 328 636 332
rect 630 327 636 328
rect 686 332 692 333
rect 686 328 687 332
rect 691 328 692 332
rect 686 327 692 328
rect 750 332 756 333
rect 750 328 751 332
rect 755 328 756 332
rect 1094 331 1095 335
rect 1099 331 1100 335
rect 1094 330 1100 331
rect 1134 335 1140 336
rect 1134 331 1135 335
rect 1139 331 1140 335
rect 2118 335 2124 336
rect 1134 330 1140 331
rect 1302 332 1308 333
rect 750 327 756 328
rect 1302 328 1303 332
rect 1307 328 1308 332
rect 1302 327 1308 328
rect 1342 332 1348 333
rect 1342 328 1343 332
rect 1347 328 1348 332
rect 1342 327 1348 328
rect 1382 332 1388 333
rect 1382 328 1383 332
rect 1387 328 1388 332
rect 1382 327 1388 328
rect 1422 332 1428 333
rect 1422 328 1423 332
rect 1427 328 1428 332
rect 1422 327 1428 328
rect 1462 332 1468 333
rect 1462 328 1463 332
rect 1467 328 1468 332
rect 1462 327 1468 328
rect 1502 332 1508 333
rect 1502 328 1503 332
rect 1507 328 1508 332
rect 1502 327 1508 328
rect 1550 332 1556 333
rect 1550 328 1551 332
rect 1555 328 1556 332
rect 1550 327 1556 328
rect 1614 332 1620 333
rect 1614 328 1615 332
rect 1619 328 1620 332
rect 1614 327 1620 328
rect 1678 332 1684 333
rect 1678 328 1679 332
rect 1683 328 1684 332
rect 1678 327 1684 328
rect 1750 332 1756 333
rect 1750 328 1751 332
rect 1755 328 1756 332
rect 1750 327 1756 328
rect 1830 332 1836 333
rect 1830 328 1831 332
rect 1835 328 1836 332
rect 1830 327 1836 328
rect 1918 332 1924 333
rect 1918 328 1919 332
rect 1923 328 1924 332
rect 1918 327 1924 328
rect 2006 332 2012 333
rect 2006 328 2007 332
rect 2011 328 2012 332
rect 2006 327 2012 328
rect 2070 332 2076 333
rect 2070 328 2071 332
rect 2075 328 2076 332
rect 2118 331 2119 335
rect 2123 331 2124 335
rect 2118 330 2124 331
rect 2070 327 2076 328
rect 134 316 140 317
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 134 312 135 316
rect 139 312 140 316
rect 134 311 140 312
rect 206 316 212 317
rect 206 312 207 316
rect 211 312 212 316
rect 206 311 212 312
rect 294 316 300 317
rect 294 312 295 316
rect 299 312 300 316
rect 294 311 300 312
rect 382 316 388 317
rect 382 312 383 316
rect 387 312 388 316
rect 382 311 388 312
rect 470 316 476 317
rect 470 312 471 316
rect 475 312 476 316
rect 470 311 476 312
rect 550 316 556 317
rect 550 312 551 316
rect 555 312 556 316
rect 550 311 556 312
rect 622 316 628 317
rect 622 312 623 316
rect 627 312 628 316
rect 622 311 628 312
rect 686 316 692 317
rect 686 312 687 316
rect 691 312 692 316
rect 686 311 692 312
rect 750 316 756 317
rect 750 312 751 316
rect 755 312 756 316
rect 750 311 756 312
rect 806 316 812 317
rect 806 312 807 316
rect 811 312 812 316
rect 806 311 812 312
rect 870 316 876 317
rect 870 312 871 316
rect 875 312 876 316
rect 870 311 876 312
rect 934 316 940 317
rect 934 312 935 316
rect 939 312 940 316
rect 1166 316 1172 317
rect 934 311 940 312
rect 1094 313 1100 314
rect 110 308 116 309
rect 1094 309 1095 313
rect 1099 309 1100 313
rect 1094 308 1100 309
rect 1134 313 1140 314
rect 1134 309 1135 313
rect 1139 309 1140 313
rect 1166 312 1167 316
rect 1171 312 1172 316
rect 1166 311 1172 312
rect 1206 316 1212 317
rect 1206 312 1207 316
rect 1211 312 1212 316
rect 1206 311 1212 312
rect 1246 316 1252 317
rect 1246 312 1247 316
rect 1251 312 1252 316
rect 1246 311 1252 312
rect 1294 316 1300 317
rect 1294 312 1295 316
rect 1299 312 1300 316
rect 1294 311 1300 312
rect 1342 316 1348 317
rect 1342 312 1343 316
rect 1347 312 1348 316
rect 1342 311 1348 312
rect 1390 316 1396 317
rect 1390 312 1391 316
rect 1395 312 1396 316
rect 1390 311 1396 312
rect 1438 316 1444 317
rect 1438 312 1439 316
rect 1443 312 1444 316
rect 1438 311 1444 312
rect 1494 316 1500 317
rect 1494 312 1495 316
rect 1499 312 1500 316
rect 1494 311 1500 312
rect 1558 316 1564 317
rect 1558 312 1559 316
rect 1563 312 1564 316
rect 1558 311 1564 312
rect 1622 316 1628 317
rect 1622 312 1623 316
rect 1627 312 1628 316
rect 1622 311 1628 312
rect 1694 316 1700 317
rect 1694 312 1695 316
rect 1699 312 1700 316
rect 1694 311 1700 312
rect 1774 316 1780 317
rect 1774 312 1775 316
rect 1779 312 1780 316
rect 1774 311 1780 312
rect 1854 316 1860 317
rect 1854 312 1855 316
rect 1859 312 1860 316
rect 1854 311 1860 312
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 1934 311 1940 312
rect 2014 316 2020 317
rect 2014 312 2015 316
rect 2019 312 2020 316
rect 2014 311 2020 312
rect 2070 316 2076 317
rect 2070 312 2071 316
rect 2075 312 2076 316
rect 2070 311 2076 312
rect 2118 313 2124 314
rect 1134 308 1140 309
rect 2118 309 2119 313
rect 2123 309 2124 313
rect 2118 308 2124 309
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 1094 296 1100 297
rect 1094 292 1095 296
rect 1099 292 1100 296
rect 1094 291 1100 292
rect 1134 296 1140 297
rect 1134 292 1135 296
rect 1139 292 1140 296
rect 1134 291 1140 292
rect 2118 296 2124 297
rect 2118 292 2119 296
rect 2123 292 2124 296
rect 2118 291 2124 292
rect 134 288 140 289
rect 134 284 135 288
rect 139 284 140 288
rect 134 283 140 284
rect 206 288 212 289
rect 206 284 207 288
rect 211 284 212 288
rect 206 283 212 284
rect 294 288 300 289
rect 294 284 295 288
rect 299 284 300 288
rect 294 283 300 284
rect 382 288 388 289
rect 382 284 383 288
rect 387 284 388 288
rect 382 283 388 284
rect 470 288 476 289
rect 470 284 471 288
rect 475 284 476 288
rect 470 283 476 284
rect 550 288 556 289
rect 550 284 551 288
rect 555 284 556 288
rect 550 283 556 284
rect 622 288 628 289
rect 622 284 623 288
rect 627 284 628 288
rect 622 283 628 284
rect 686 288 692 289
rect 686 284 687 288
rect 691 284 692 288
rect 686 283 692 284
rect 750 288 756 289
rect 750 284 751 288
rect 755 284 756 288
rect 750 283 756 284
rect 806 288 812 289
rect 806 284 807 288
rect 811 284 812 288
rect 806 283 812 284
rect 870 288 876 289
rect 870 284 871 288
rect 875 284 876 288
rect 870 283 876 284
rect 934 288 940 289
rect 934 284 935 288
rect 939 284 940 288
rect 934 283 940 284
rect 1166 288 1172 289
rect 1166 284 1167 288
rect 1171 284 1172 288
rect 1166 283 1172 284
rect 1206 288 1212 289
rect 1206 284 1207 288
rect 1211 284 1212 288
rect 1206 283 1212 284
rect 1246 288 1252 289
rect 1246 284 1247 288
rect 1251 284 1252 288
rect 1246 283 1252 284
rect 1294 288 1300 289
rect 1294 284 1295 288
rect 1299 284 1300 288
rect 1294 283 1300 284
rect 1342 288 1348 289
rect 1342 284 1343 288
rect 1347 284 1348 288
rect 1342 283 1348 284
rect 1390 288 1396 289
rect 1390 284 1391 288
rect 1395 284 1396 288
rect 1390 283 1396 284
rect 1438 288 1444 289
rect 1438 284 1439 288
rect 1443 284 1444 288
rect 1438 283 1444 284
rect 1494 288 1500 289
rect 1494 284 1495 288
rect 1499 284 1500 288
rect 1494 283 1500 284
rect 1558 288 1564 289
rect 1558 284 1559 288
rect 1563 284 1564 288
rect 1558 283 1564 284
rect 1622 288 1628 289
rect 1622 284 1623 288
rect 1627 284 1628 288
rect 1622 283 1628 284
rect 1694 288 1700 289
rect 1694 284 1695 288
rect 1699 284 1700 288
rect 1694 283 1700 284
rect 1774 288 1780 289
rect 1774 284 1775 288
rect 1779 284 1780 288
rect 1774 283 1780 284
rect 1854 288 1860 289
rect 1854 284 1855 288
rect 1859 284 1860 288
rect 1854 283 1860 284
rect 1934 288 1940 289
rect 1934 284 1935 288
rect 1939 284 1940 288
rect 1934 283 1940 284
rect 2014 288 2020 289
rect 2014 284 2015 288
rect 2019 284 2020 288
rect 2014 283 2020 284
rect 2070 288 2076 289
rect 2070 284 2071 288
rect 2075 284 2076 288
rect 2070 283 2076 284
rect 134 252 140 253
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 198 252 204 253
rect 198 248 199 252
rect 203 248 204 252
rect 198 247 204 248
rect 278 252 284 253
rect 278 248 279 252
rect 283 248 284 252
rect 278 247 284 248
rect 358 252 364 253
rect 358 248 359 252
rect 363 248 364 252
rect 358 247 364 248
rect 438 252 444 253
rect 438 248 439 252
rect 443 248 444 252
rect 438 247 444 248
rect 510 252 516 253
rect 510 248 511 252
rect 515 248 516 252
rect 510 247 516 248
rect 582 252 588 253
rect 582 248 583 252
rect 587 248 588 252
rect 582 247 588 248
rect 646 252 652 253
rect 646 248 647 252
rect 651 248 652 252
rect 646 247 652 248
rect 702 252 708 253
rect 702 248 703 252
rect 707 248 708 252
rect 702 247 708 248
rect 758 252 764 253
rect 758 248 759 252
rect 763 248 764 252
rect 758 247 764 248
rect 814 252 820 253
rect 814 248 815 252
rect 819 248 820 252
rect 814 247 820 248
rect 878 252 884 253
rect 878 248 879 252
rect 883 248 884 252
rect 878 247 884 248
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 110 239 116 240
rect 1094 244 1100 245
rect 1094 240 1095 244
rect 1099 240 1100 244
rect 1094 239 1100 240
rect 1158 244 1164 245
rect 1158 240 1159 244
rect 1163 240 1164 244
rect 1158 239 1164 240
rect 1206 244 1212 245
rect 1206 240 1207 244
rect 1211 240 1212 244
rect 1206 239 1212 240
rect 1270 244 1276 245
rect 1270 240 1271 244
rect 1275 240 1276 244
rect 1270 239 1276 240
rect 1326 244 1332 245
rect 1326 240 1327 244
rect 1331 240 1332 244
rect 1326 239 1332 240
rect 1390 244 1396 245
rect 1390 240 1391 244
rect 1395 240 1396 244
rect 1390 239 1396 240
rect 1454 244 1460 245
rect 1454 240 1455 244
rect 1459 240 1460 244
rect 1454 239 1460 240
rect 1526 244 1532 245
rect 1526 240 1527 244
rect 1531 240 1532 244
rect 1526 239 1532 240
rect 1606 244 1612 245
rect 1606 240 1607 244
rect 1611 240 1612 244
rect 1606 239 1612 240
rect 1686 244 1692 245
rect 1686 240 1687 244
rect 1691 240 1692 244
rect 1686 239 1692 240
rect 1766 244 1772 245
rect 1766 240 1767 244
rect 1771 240 1772 244
rect 1766 239 1772 240
rect 1838 244 1844 245
rect 1838 240 1839 244
rect 1843 240 1844 244
rect 1838 239 1844 240
rect 1918 244 1924 245
rect 1918 240 1919 244
rect 1923 240 1924 244
rect 1918 239 1924 240
rect 1998 244 2004 245
rect 1998 240 1999 244
rect 2003 240 2004 244
rect 1998 239 2004 240
rect 2070 244 2076 245
rect 2070 240 2071 244
rect 2075 240 2076 244
rect 2070 239 2076 240
rect 1134 236 1140 237
rect 1134 232 1135 236
rect 1139 232 1140 236
rect 1134 231 1140 232
rect 2118 236 2124 237
rect 2118 232 2119 236
rect 2123 232 2124 236
rect 2118 231 2124 232
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1094 227 1100 228
rect 110 222 116 223
rect 134 224 140 225
rect 134 220 135 224
rect 139 220 140 224
rect 134 219 140 220
rect 198 224 204 225
rect 198 220 199 224
rect 203 220 204 224
rect 198 219 204 220
rect 278 224 284 225
rect 278 220 279 224
rect 283 220 284 224
rect 278 219 284 220
rect 358 224 364 225
rect 358 220 359 224
rect 363 220 364 224
rect 358 219 364 220
rect 438 224 444 225
rect 438 220 439 224
rect 443 220 444 224
rect 438 219 444 220
rect 510 224 516 225
rect 510 220 511 224
rect 515 220 516 224
rect 510 219 516 220
rect 582 224 588 225
rect 582 220 583 224
rect 587 220 588 224
rect 582 219 588 220
rect 646 224 652 225
rect 646 220 647 224
rect 651 220 652 224
rect 646 219 652 220
rect 702 224 708 225
rect 702 220 703 224
rect 707 220 708 224
rect 702 219 708 220
rect 758 224 764 225
rect 758 220 759 224
rect 763 220 764 224
rect 758 219 764 220
rect 814 224 820 225
rect 814 220 815 224
rect 819 220 820 224
rect 814 219 820 220
rect 878 224 884 225
rect 878 220 879 224
rect 883 220 884 224
rect 1094 223 1095 227
rect 1099 223 1100 227
rect 1094 222 1100 223
rect 878 219 884 220
rect 1134 219 1140 220
rect 1134 215 1135 219
rect 1139 215 1140 219
rect 2118 219 2124 220
rect 1134 214 1140 215
rect 1158 216 1164 217
rect 1158 212 1159 216
rect 1163 212 1164 216
rect 1158 211 1164 212
rect 1206 216 1212 217
rect 1206 212 1207 216
rect 1211 212 1212 216
rect 1206 211 1212 212
rect 1270 216 1276 217
rect 1270 212 1271 216
rect 1275 212 1276 216
rect 1270 211 1276 212
rect 1326 216 1332 217
rect 1326 212 1327 216
rect 1331 212 1332 216
rect 1326 211 1332 212
rect 1390 216 1396 217
rect 1390 212 1391 216
rect 1395 212 1396 216
rect 1390 211 1396 212
rect 1454 216 1460 217
rect 1454 212 1455 216
rect 1459 212 1460 216
rect 1454 211 1460 212
rect 1526 216 1532 217
rect 1526 212 1527 216
rect 1531 212 1532 216
rect 1526 211 1532 212
rect 1606 216 1612 217
rect 1606 212 1607 216
rect 1611 212 1612 216
rect 1606 211 1612 212
rect 1686 216 1692 217
rect 1686 212 1687 216
rect 1691 212 1692 216
rect 1686 211 1692 212
rect 1766 216 1772 217
rect 1766 212 1767 216
rect 1771 212 1772 216
rect 1766 211 1772 212
rect 1838 216 1844 217
rect 1838 212 1839 216
rect 1843 212 1844 216
rect 1838 211 1844 212
rect 1918 216 1924 217
rect 1918 212 1919 216
rect 1923 212 1924 216
rect 1918 211 1924 212
rect 1998 216 2004 217
rect 1998 212 1999 216
rect 2003 212 2004 216
rect 1998 211 2004 212
rect 2070 216 2076 217
rect 2070 212 2071 216
rect 2075 212 2076 216
rect 2118 215 2119 219
rect 2123 215 2124 219
rect 2118 214 2124 215
rect 2070 211 2076 212
rect 134 208 140 209
rect 110 205 116 206
rect 110 201 111 205
rect 115 201 116 205
rect 134 204 135 208
rect 139 204 140 208
rect 134 203 140 204
rect 182 208 188 209
rect 182 204 183 208
rect 187 204 188 208
rect 182 203 188 204
rect 230 208 236 209
rect 230 204 231 208
rect 235 204 236 208
rect 230 203 236 204
rect 278 208 284 209
rect 278 204 279 208
rect 283 204 284 208
rect 278 203 284 204
rect 326 208 332 209
rect 326 204 327 208
rect 331 204 332 208
rect 326 203 332 204
rect 374 208 380 209
rect 374 204 375 208
rect 379 204 380 208
rect 374 203 380 204
rect 414 208 420 209
rect 414 204 415 208
rect 419 204 420 208
rect 414 203 420 204
rect 454 208 460 209
rect 454 204 455 208
rect 459 204 460 208
rect 454 203 460 204
rect 502 208 508 209
rect 502 204 503 208
rect 507 204 508 208
rect 502 203 508 204
rect 550 208 556 209
rect 550 204 551 208
rect 555 204 556 208
rect 550 203 556 204
rect 598 208 604 209
rect 598 204 599 208
rect 603 204 604 208
rect 598 203 604 204
rect 646 208 652 209
rect 646 204 647 208
rect 651 204 652 208
rect 646 203 652 204
rect 694 208 700 209
rect 694 204 695 208
rect 699 204 700 208
rect 694 203 700 204
rect 742 208 748 209
rect 742 204 743 208
rect 747 204 748 208
rect 742 203 748 204
rect 1094 205 1100 206
rect 110 200 116 201
rect 1094 201 1095 205
rect 1099 201 1100 205
rect 1158 204 1164 205
rect 1094 200 1100 201
rect 1134 201 1140 202
rect 1134 197 1135 201
rect 1139 197 1140 201
rect 1158 200 1159 204
rect 1163 200 1164 204
rect 1158 199 1164 200
rect 1198 204 1204 205
rect 1198 200 1199 204
rect 1203 200 1204 204
rect 1198 199 1204 200
rect 1262 204 1268 205
rect 1262 200 1263 204
rect 1267 200 1268 204
rect 1262 199 1268 200
rect 1326 204 1332 205
rect 1326 200 1327 204
rect 1331 200 1332 204
rect 1326 199 1332 200
rect 1398 204 1404 205
rect 1398 200 1399 204
rect 1403 200 1404 204
rect 1398 199 1404 200
rect 1470 204 1476 205
rect 1470 200 1471 204
rect 1475 200 1476 204
rect 1470 199 1476 200
rect 1542 204 1548 205
rect 1542 200 1543 204
rect 1547 200 1548 204
rect 1542 199 1548 200
rect 1606 204 1612 205
rect 1606 200 1607 204
rect 1611 200 1612 204
rect 1606 199 1612 200
rect 1670 204 1676 205
rect 1670 200 1671 204
rect 1675 200 1676 204
rect 1670 199 1676 200
rect 1734 204 1740 205
rect 1734 200 1735 204
rect 1739 200 1740 204
rect 1734 199 1740 200
rect 1806 204 1812 205
rect 1806 200 1807 204
rect 1811 200 1812 204
rect 1806 199 1812 200
rect 1878 204 1884 205
rect 1878 200 1879 204
rect 1883 200 1884 204
rect 1878 199 1884 200
rect 1950 204 1956 205
rect 1950 200 1951 204
rect 1955 200 1956 204
rect 1950 199 1956 200
rect 2022 204 2028 205
rect 2022 200 2023 204
rect 2027 200 2028 204
rect 2022 199 2028 200
rect 2070 204 2076 205
rect 2070 200 2071 204
rect 2075 200 2076 204
rect 2070 199 2076 200
rect 2118 201 2124 202
rect 1134 196 1140 197
rect 2118 197 2119 201
rect 2123 197 2124 201
rect 2118 196 2124 197
rect 110 188 116 189
rect 110 184 111 188
rect 115 184 116 188
rect 110 183 116 184
rect 1094 188 1100 189
rect 1094 184 1095 188
rect 1099 184 1100 188
rect 1094 183 1100 184
rect 1134 184 1140 185
rect 134 180 140 181
rect 134 176 135 180
rect 139 176 140 180
rect 134 175 140 176
rect 182 180 188 181
rect 182 176 183 180
rect 187 176 188 180
rect 182 175 188 176
rect 230 180 236 181
rect 230 176 231 180
rect 235 176 236 180
rect 230 175 236 176
rect 278 180 284 181
rect 278 176 279 180
rect 283 176 284 180
rect 278 175 284 176
rect 326 180 332 181
rect 326 176 327 180
rect 331 176 332 180
rect 326 175 332 176
rect 374 180 380 181
rect 374 176 375 180
rect 379 176 380 180
rect 374 175 380 176
rect 414 180 420 181
rect 414 176 415 180
rect 419 176 420 180
rect 414 175 420 176
rect 454 180 460 181
rect 454 176 455 180
rect 459 176 460 180
rect 454 175 460 176
rect 502 180 508 181
rect 502 176 503 180
rect 507 176 508 180
rect 502 175 508 176
rect 550 180 556 181
rect 550 176 551 180
rect 555 176 556 180
rect 550 175 556 176
rect 598 180 604 181
rect 598 176 599 180
rect 603 176 604 180
rect 598 175 604 176
rect 646 180 652 181
rect 646 176 647 180
rect 651 176 652 180
rect 646 175 652 176
rect 694 180 700 181
rect 694 176 695 180
rect 699 176 700 180
rect 694 175 700 176
rect 742 180 748 181
rect 742 176 743 180
rect 747 176 748 180
rect 1134 180 1135 184
rect 1139 180 1140 184
rect 1134 179 1140 180
rect 2118 184 2124 185
rect 2118 180 2119 184
rect 2123 180 2124 184
rect 2118 179 2124 180
rect 742 175 748 176
rect 1158 176 1164 177
rect 1158 172 1159 176
rect 1163 172 1164 176
rect 1158 171 1164 172
rect 1198 176 1204 177
rect 1198 172 1199 176
rect 1203 172 1204 176
rect 1198 171 1204 172
rect 1262 176 1268 177
rect 1262 172 1263 176
rect 1267 172 1268 176
rect 1262 171 1268 172
rect 1326 176 1332 177
rect 1326 172 1327 176
rect 1331 172 1332 176
rect 1326 171 1332 172
rect 1398 176 1404 177
rect 1398 172 1399 176
rect 1403 172 1404 176
rect 1398 171 1404 172
rect 1470 176 1476 177
rect 1470 172 1471 176
rect 1475 172 1476 176
rect 1470 171 1476 172
rect 1542 176 1548 177
rect 1542 172 1543 176
rect 1547 172 1548 176
rect 1542 171 1548 172
rect 1606 176 1612 177
rect 1606 172 1607 176
rect 1611 172 1612 176
rect 1606 171 1612 172
rect 1670 176 1676 177
rect 1670 172 1671 176
rect 1675 172 1676 176
rect 1670 171 1676 172
rect 1734 176 1740 177
rect 1734 172 1735 176
rect 1739 172 1740 176
rect 1734 171 1740 172
rect 1806 176 1812 177
rect 1806 172 1807 176
rect 1811 172 1812 176
rect 1806 171 1812 172
rect 1878 176 1884 177
rect 1878 172 1879 176
rect 1883 172 1884 176
rect 1878 171 1884 172
rect 1950 176 1956 177
rect 1950 172 1951 176
rect 1955 172 1956 176
rect 1950 171 1956 172
rect 2022 176 2028 177
rect 2022 172 2023 176
rect 2027 172 2028 176
rect 2022 171 2028 172
rect 2070 176 2076 177
rect 2070 172 2071 176
rect 2075 172 2076 176
rect 2070 171 2076 172
rect 142 120 148 121
rect 142 116 143 120
rect 147 116 148 120
rect 142 115 148 116
rect 182 120 188 121
rect 182 116 183 120
rect 187 116 188 120
rect 182 115 188 116
rect 222 120 228 121
rect 222 116 223 120
rect 227 116 228 120
rect 222 115 228 116
rect 262 120 268 121
rect 262 116 263 120
rect 267 116 268 120
rect 262 115 268 116
rect 302 120 308 121
rect 302 116 303 120
rect 307 116 308 120
rect 302 115 308 116
rect 342 120 348 121
rect 342 116 343 120
rect 347 116 348 120
rect 342 115 348 116
rect 382 120 388 121
rect 382 116 383 120
rect 387 116 388 120
rect 382 115 388 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 462 120 468 121
rect 462 116 463 120
rect 467 116 468 120
rect 462 115 468 116
rect 502 120 508 121
rect 502 116 503 120
rect 507 116 508 120
rect 502 115 508 116
rect 542 120 548 121
rect 542 116 543 120
rect 547 116 548 120
rect 542 115 548 116
rect 582 120 588 121
rect 582 116 583 120
rect 587 116 588 120
rect 582 115 588 116
rect 622 120 628 121
rect 622 116 623 120
rect 627 116 628 120
rect 622 115 628 116
rect 662 120 668 121
rect 662 116 663 120
rect 667 116 668 120
rect 662 115 668 116
rect 702 120 708 121
rect 702 116 703 120
rect 707 116 708 120
rect 702 115 708 116
rect 742 120 748 121
rect 742 116 743 120
rect 747 116 748 120
rect 742 115 748 116
rect 782 120 788 121
rect 782 116 783 120
rect 787 116 788 120
rect 782 115 788 116
rect 830 120 836 121
rect 830 116 831 120
rect 835 116 836 120
rect 830 115 836 116
rect 878 120 884 121
rect 878 116 879 120
rect 883 116 884 120
rect 878 115 884 116
rect 926 120 932 121
rect 926 116 927 120
rect 931 116 932 120
rect 926 115 932 116
rect 966 120 972 121
rect 966 116 967 120
rect 971 116 972 120
rect 966 115 972 116
rect 1006 120 1012 121
rect 1006 116 1007 120
rect 1011 116 1012 120
rect 1006 115 1012 116
rect 1046 120 1052 121
rect 1046 116 1047 120
rect 1051 116 1052 120
rect 1046 115 1052 116
rect 1158 120 1164 121
rect 1158 116 1159 120
rect 1163 116 1164 120
rect 1158 115 1164 116
rect 1206 120 1212 121
rect 1206 116 1207 120
rect 1211 116 1212 120
rect 1206 115 1212 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1334 120 1340 121
rect 1334 116 1335 120
rect 1339 116 1340 120
rect 1334 115 1340 116
rect 1398 120 1404 121
rect 1398 116 1399 120
rect 1403 116 1404 120
rect 1398 115 1404 116
rect 1454 120 1460 121
rect 1454 116 1455 120
rect 1459 116 1460 120
rect 1454 115 1460 116
rect 1510 120 1516 121
rect 1510 116 1511 120
rect 1515 116 1516 120
rect 1510 115 1516 116
rect 1558 120 1564 121
rect 1558 116 1559 120
rect 1563 116 1564 120
rect 1558 115 1564 116
rect 1606 120 1612 121
rect 1606 116 1607 120
rect 1611 116 1612 120
rect 1606 115 1612 116
rect 1646 120 1652 121
rect 1646 116 1647 120
rect 1651 116 1652 120
rect 1646 115 1652 116
rect 1686 120 1692 121
rect 1686 116 1687 120
rect 1691 116 1692 120
rect 1686 115 1692 116
rect 1726 120 1732 121
rect 1726 116 1727 120
rect 1731 116 1732 120
rect 1726 115 1732 116
rect 1766 120 1772 121
rect 1766 116 1767 120
rect 1771 116 1772 120
rect 1766 115 1772 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1854 120 1860 121
rect 1854 116 1855 120
rect 1859 116 1860 120
rect 1854 115 1860 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 1902 115 1908 116
rect 1950 120 1956 121
rect 1950 116 1951 120
rect 1955 116 1956 120
rect 1950 115 1956 116
rect 1990 120 1996 121
rect 1990 116 1991 120
rect 1995 116 1996 120
rect 1990 115 1996 116
rect 2030 120 2036 121
rect 2030 116 2031 120
rect 2035 116 2036 120
rect 2030 115 2036 116
rect 2070 120 2076 121
rect 2070 116 2071 120
rect 2075 116 2076 120
rect 2070 115 2076 116
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 110 107 116 108
rect 1094 112 1100 113
rect 1094 108 1095 112
rect 1099 108 1100 112
rect 1094 107 1100 108
rect 1134 112 1140 113
rect 1134 108 1135 112
rect 1139 108 1140 112
rect 1134 107 1140 108
rect 2118 112 2124 113
rect 2118 108 2119 112
rect 2123 108 2124 112
rect 2118 107 2124 108
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1094 95 1100 96
rect 110 90 116 91
rect 142 92 148 93
rect 142 88 143 92
rect 147 88 148 92
rect 142 87 148 88
rect 182 92 188 93
rect 182 88 183 92
rect 187 88 188 92
rect 182 87 188 88
rect 222 92 228 93
rect 222 88 223 92
rect 227 88 228 92
rect 222 87 228 88
rect 262 92 268 93
rect 262 88 263 92
rect 267 88 268 92
rect 262 87 268 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 342 92 348 93
rect 342 88 343 92
rect 347 88 348 92
rect 342 87 348 88
rect 382 92 388 93
rect 382 88 383 92
rect 387 88 388 92
rect 382 87 388 88
rect 422 92 428 93
rect 422 88 423 92
rect 427 88 428 92
rect 422 87 428 88
rect 462 92 468 93
rect 462 88 463 92
rect 467 88 468 92
rect 462 87 468 88
rect 502 92 508 93
rect 502 88 503 92
rect 507 88 508 92
rect 502 87 508 88
rect 542 92 548 93
rect 542 88 543 92
rect 547 88 548 92
rect 542 87 548 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 622 92 628 93
rect 622 88 623 92
rect 627 88 628 92
rect 622 87 628 88
rect 662 92 668 93
rect 662 88 663 92
rect 667 88 668 92
rect 662 87 668 88
rect 702 92 708 93
rect 702 88 703 92
rect 707 88 708 92
rect 702 87 708 88
rect 742 92 748 93
rect 742 88 743 92
rect 747 88 748 92
rect 742 87 748 88
rect 782 92 788 93
rect 782 88 783 92
rect 787 88 788 92
rect 782 87 788 88
rect 830 92 836 93
rect 830 88 831 92
rect 835 88 836 92
rect 830 87 836 88
rect 878 92 884 93
rect 878 88 879 92
rect 883 88 884 92
rect 878 87 884 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 966 92 972 93
rect 966 88 967 92
rect 971 88 972 92
rect 966 87 972 88
rect 1006 92 1012 93
rect 1006 88 1007 92
rect 1011 88 1012 92
rect 1006 87 1012 88
rect 1046 92 1052 93
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1094 91 1095 95
rect 1099 91 1100 95
rect 1094 90 1100 91
rect 1134 95 1140 96
rect 1134 91 1135 95
rect 1139 91 1140 95
rect 2118 95 2124 96
rect 1134 90 1140 91
rect 1158 92 1164 93
rect 1046 87 1052 88
rect 1158 88 1159 92
rect 1163 88 1164 92
rect 1158 87 1164 88
rect 1206 92 1212 93
rect 1206 88 1207 92
rect 1211 88 1212 92
rect 1206 87 1212 88
rect 1270 92 1276 93
rect 1270 88 1271 92
rect 1275 88 1276 92
rect 1270 87 1276 88
rect 1334 92 1340 93
rect 1334 88 1335 92
rect 1339 88 1340 92
rect 1334 87 1340 88
rect 1398 92 1404 93
rect 1398 88 1399 92
rect 1403 88 1404 92
rect 1398 87 1404 88
rect 1454 92 1460 93
rect 1454 88 1455 92
rect 1459 88 1460 92
rect 1454 87 1460 88
rect 1510 92 1516 93
rect 1510 88 1511 92
rect 1515 88 1516 92
rect 1510 87 1516 88
rect 1558 92 1564 93
rect 1558 88 1559 92
rect 1563 88 1564 92
rect 1558 87 1564 88
rect 1606 92 1612 93
rect 1606 88 1607 92
rect 1611 88 1612 92
rect 1606 87 1612 88
rect 1646 92 1652 93
rect 1646 88 1647 92
rect 1651 88 1652 92
rect 1646 87 1652 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1726 92 1732 93
rect 1726 88 1727 92
rect 1731 88 1732 92
rect 1726 87 1732 88
rect 1766 92 1772 93
rect 1766 88 1767 92
rect 1771 88 1772 92
rect 1766 87 1772 88
rect 1806 92 1812 93
rect 1806 88 1807 92
rect 1811 88 1812 92
rect 1806 87 1812 88
rect 1854 92 1860 93
rect 1854 88 1855 92
rect 1859 88 1860 92
rect 1854 87 1860 88
rect 1902 92 1908 93
rect 1902 88 1903 92
rect 1907 88 1908 92
rect 1902 87 1908 88
rect 1950 92 1956 93
rect 1950 88 1951 92
rect 1955 88 1956 92
rect 1950 87 1956 88
rect 1990 92 1996 93
rect 1990 88 1991 92
rect 1995 88 1996 92
rect 1990 87 1996 88
rect 2030 92 2036 93
rect 2030 88 2031 92
rect 2035 88 2036 92
rect 2030 87 2036 88
rect 2070 92 2076 93
rect 2070 88 2071 92
rect 2075 88 2076 92
rect 2118 91 2119 95
rect 2123 91 2124 95
rect 2118 90 2124 91
rect 2070 87 2076 88
<< m3c >>
rect 111 2201 115 2205
rect 135 2204 139 2208
rect 175 2204 179 2208
rect 215 2204 219 2208
rect 255 2204 259 2208
rect 319 2204 323 2208
rect 383 2204 387 2208
rect 447 2204 451 2208
rect 511 2204 515 2208
rect 575 2204 579 2208
rect 631 2204 635 2208
rect 687 2204 691 2208
rect 735 2204 739 2208
rect 791 2204 795 2208
rect 847 2204 851 2208
rect 903 2204 907 2208
rect 1687 2208 1691 2212
rect 1727 2208 1731 2212
rect 1767 2208 1771 2212
rect 1807 2208 1811 2212
rect 1095 2201 1099 2205
rect 1135 2200 1139 2204
rect 2119 2200 2123 2204
rect 111 2184 115 2188
rect 1095 2184 1099 2188
rect 1135 2183 1139 2187
rect 135 2176 139 2180
rect 175 2176 179 2180
rect 215 2176 219 2180
rect 255 2176 259 2180
rect 319 2176 323 2180
rect 383 2176 387 2180
rect 447 2176 451 2180
rect 511 2176 515 2180
rect 575 2176 579 2180
rect 631 2176 635 2180
rect 687 2176 691 2180
rect 735 2176 739 2180
rect 791 2176 795 2180
rect 847 2176 851 2180
rect 903 2176 907 2180
rect 1687 2180 1691 2184
rect 1727 2180 1731 2184
rect 1767 2180 1771 2184
rect 1807 2180 1811 2184
rect 2119 2183 2123 2187
rect 1135 2165 1139 2169
rect 1159 2168 1163 2172
rect 1199 2168 1203 2172
rect 1239 2168 1243 2172
rect 1279 2168 1283 2172
rect 1335 2168 1339 2172
rect 1391 2168 1395 2172
rect 1455 2168 1459 2172
rect 1527 2168 1531 2172
rect 1591 2168 1595 2172
rect 1663 2168 1667 2172
rect 1735 2168 1739 2172
rect 1807 2168 1811 2172
rect 1879 2168 1883 2172
rect 2119 2165 2123 2169
rect 1135 2148 1139 2152
rect 2119 2148 2123 2152
rect 1159 2140 1163 2144
rect 1199 2140 1203 2144
rect 1239 2140 1243 2144
rect 1279 2140 1283 2144
rect 1335 2140 1339 2144
rect 1391 2140 1395 2144
rect 1455 2140 1459 2144
rect 1527 2140 1531 2144
rect 1591 2140 1595 2144
rect 1663 2140 1667 2144
rect 1735 2140 1739 2144
rect 1807 2140 1811 2144
rect 1879 2140 1883 2144
rect 231 2132 235 2136
rect 271 2132 275 2136
rect 311 2132 315 2136
rect 359 2132 363 2136
rect 423 2132 427 2136
rect 487 2132 491 2136
rect 559 2132 563 2136
rect 639 2132 643 2136
rect 719 2132 723 2136
rect 799 2132 803 2136
rect 879 2132 883 2136
rect 967 2132 971 2136
rect 111 2124 115 2128
rect 1095 2124 1099 2128
rect 111 2107 115 2111
rect 231 2104 235 2108
rect 271 2104 275 2108
rect 311 2104 315 2108
rect 359 2104 363 2108
rect 423 2104 427 2108
rect 487 2104 491 2108
rect 559 2104 563 2108
rect 639 2104 643 2108
rect 719 2104 723 2108
rect 799 2104 803 2108
rect 879 2104 883 2108
rect 967 2104 971 2108
rect 1095 2107 1099 2111
rect 1159 2104 1163 2108
rect 1199 2104 1203 2108
rect 1239 2104 1243 2108
rect 1295 2104 1299 2108
rect 1367 2104 1371 2108
rect 1439 2104 1443 2108
rect 1519 2104 1523 2108
rect 1599 2104 1603 2108
rect 1679 2104 1683 2108
rect 1751 2104 1755 2108
rect 1823 2104 1827 2108
rect 1887 2104 1891 2108
rect 1951 2104 1955 2108
rect 2023 2104 2027 2108
rect 2071 2104 2075 2108
rect 1135 2096 1139 2100
rect 2119 2096 2123 2100
rect 111 2085 115 2089
rect 303 2088 307 2092
rect 351 2088 355 2092
rect 407 2088 411 2092
rect 471 2088 475 2092
rect 543 2088 547 2092
rect 623 2088 627 2092
rect 703 2088 707 2092
rect 783 2088 787 2092
rect 863 2088 867 2092
rect 951 2088 955 2092
rect 1039 2088 1043 2092
rect 1095 2085 1099 2089
rect 1135 2079 1139 2083
rect 1159 2076 1163 2080
rect 1199 2076 1203 2080
rect 1239 2076 1243 2080
rect 1295 2076 1299 2080
rect 1367 2076 1371 2080
rect 1439 2076 1443 2080
rect 1519 2076 1523 2080
rect 1599 2076 1603 2080
rect 1679 2076 1683 2080
rect 1751 2076 1755 2080
rect 1823 2076 1827 2080
rect 1887 2076 1891 2080
rect 1951 2076 1955 2080
rect 2023 2076 2027 2080
rect 2071 2076 2075 2080
rect 2119 2079 2123 2083
rect 111 2068 115 2072
rect 1095 2068 1099 2072
rect 303 2060 307 2064
rect 351 2060 355 2064
rect 407 2060 411 2064
rect 471 2060 475 2064
rect 543 2060 547 2064
rect 623 2060 627 2064
rect 703 2060 707 2064
rect 783 2060 787 2064
rect 863 2060 867 2064
rect 951 2060 955 2064
rect 1039 2060 1043 2064
rect 1135 2061 1139 2065
rect 1159 2064 1163 2068
rect 1215 2064 1219 2068
rect 1303 2064 1307 2068
rect 1399 2064 1403 2068
rect 1495 2064 1499 2068
rect 1591 2064 1595 2068
rect 1679 2064 1683 2068
rect 1759 2064 1763 2068
rect 1831 2064 1835 2068
rect 1895 2064 1899 2068
rect 1959 2064 1963 2068
rect 2023 2064 2027 2068
rect 2071 2064 2075 2068
rect 2119 2061 2123 2065
rect 1135 2044 1139 2048
rect 2119 2044 2123 2048
rect 1159 2036 1163 2040
rect 1215 2036 1219 2040
rect 1303 2036 1307 2040
rect 1399 2036 1403 2040
rect 1495 2036 1499 2040
rect 1591 2036 1595 2040
rect 1679 2036 1683 2040
rect 1759 2036 1763 2040
rect 1831 2036 1835 2040
rect 1895 2036 1899 2040
rect 1959 2036 1963 2040
rect 2023 2036 2027 2040
rect 2071 2036 2075 2040
rect 183 2020 187 2024
rect 279 2020 283 2024
rect 375 2020 379 2024
rect 463 2020 467 2024
rect 543 2020 547 2024
rect 623 2020 627 2024
rect 695 2020 699 2024
rect 759 2020 763 2024
rect 815 2020 819 2024
rect 863 2020 867 2024
rect 911 2020 915 2024
rect 959 2020 963 2024
rect 1007 2020 1011 2024
rect 1047 2020 1051 2024
rect 111 2012 115 2016
rect 1095 2012 1099 2016
rect 1159 2000 1163 2004
rect 111 1995 115 1999
rect 1239 2000 1243 2004
rect 1351 2000 1355 2004
rect 1455 2000 1459 2004
rect 1559 2000 1563 2004
rect 1655 2000 1659 2004
rect 1743 2000 1747 2004
rect 1823 2000 1827 2004
rect 1895 2000 1899 2004
rect 1959 2000 1963 2004
rect 2023 2000 2027 2004
rect 2071 2000 2075 2004
rect 183 1992 187 1996
rect 279 1992 283 1996
rect 375 1992 379 1996
rect 463 1992 467 1996
rect 543 1992 547 1996
rect 623 1992 627 1996
rect 695 1992 699 1996
rect 759 1992 763 1996
rect 815 1992 819 1996
rect 863 1992 867 1996
rect 911 1992 915 1996
rect 959 1992 963 1996
rect 1007 1992 1011 1996
rect 1047 1992 1051 1996
rect 1095 1995 1099 1999
rect 1135 1992 1139 1996
rect 2119 1992 2123 1996
rect 111 1977 115 1981
rect 159 1980 163 1984
rect 231 1980 235 1984
rect 303 1980 307 1984
rect 375 1980 379 1984
rect 447 1980 451 1984
rect 527 1980 531 1984
rect 607 1980 611 1984
rect 687 1980 691 1984
rect 759 1980 763 1984
rect 831 1980 835 1984
rect 911 1980 915 1984
rect 991 1980 995 1984
rect 1095 1977 1099 1981
rect 1135 1975 1139 1979
rect 1159 1972 1163 1976
rect 1239 1972 1243 1976
rect 1351 1972 1355 1976
rect 1455 1972 1459 1976
rect 1559 1972 1563 1976
rect 1655 1972 1659 1976
rect 1743 1972 1747 1976
rect 1823 1972 1827 1976
rect 1895 1972 1899 1976
rect 1959 1972 1963 1976
rect 2023 1972 2027 1976
rect 2071 1972 2075 1976
rect 2119 1975 2123 1979
rect 111 1960 115 1964
rect 1095 1960 1099 1964
rect 159 1952 163 1956
rect 231 1952 235 1956
rect 303 1952 307 1956
rect 375 1952 379 1956
rect 447 1952 451 1956
rect 527 1952 531 1956
rect 607 1952 611 1956
rect 687 1952 691 1956
rect 759 1952 763 1956
rect 831 1952 835 1956
rect 911 1952 915 1956
rect 991 1952 995 1956
rect 1135 1945 1139 1949
rect 1359 1948 1363 1952
rect 1423 1948 1427 1952
rect 1487 1948 1491 1952
rect 1559 1948 1563 1952
rect 1631 1948 1635 1952
rect 1703 1948 1707 1952
rect 1775 1948 1779 1952
rect 1847 1948 1851 1952
rect 1927 1948 1931 1952
rect 2007 1948 2011 1952
rect 2071 1948 2075 1952
rect 2119 1945 2123 1949
rect 1135 1928 1139 1932
rect 2119 1928 2123 1932
rect 1359 1920 1363 1924
rect 1423 1920 1427 1924
rect 1487 1920 1491 1924
rect 1559 1920 1563 1924
rect 1631 1920 1635 1924
rect 1703 1920 1707 1924
rect 1775 1920 1779 1924
rect 1847 1920 1851 1924
rect 1927 1920 1931 1924
rect 2007 1920 2011 1924
rect 2071 1920 2075 1924
rect 135 1912 139 1916
rect 175 1912 179 1916
rect 231 1912 235 1916
rect 295 1912 299 1916
rect 367 1912 371 1916
rect 447 1912 451 1916
rect 527 1912 531 1916
rect 615 1912 619 1916
rect 703 1912 707 1916
rect 791 1912 795 1916
rect 879 1912 883 1916
rect 111 1904 115 1908
rect 1095 1904 1099 1908
rect 111 1887 115 1891
rect 135 1884 139 1888
rect 175 1884 179 1888
rect 231 1884 235 1888
rect 295 1884 299 1888
rect 367 1884 371 1888
rect 447 1884 451 1888
rect 527 1884 531 1888
rect 615 1884 619 1888
rect 703 1884 707 1888
rect 791 1884 795 1888
rect 879 1884 883 1888
rect 1095 1887 1099 1891
rect 1231 1884 1235 1888
rect 1271 1884 1275 1888
rect 1319 1884 1323 1888
rect 1375 1884 1379 1888
rect 1439 1884 1443 1888
rect 1503 1884 1507 1888
rect 1575 1884 1579 1888
rect 1655 1884 1659 1888
rect 1751 1884 1755 1888
rect 1863 1884 1867 1888
rect 1975 1884 1979 1888
rect 2071 1884 2075 1888
rect 1135 1876 1139 1880
rect 2119 1876 2123 1880
rect 111 1865 115 1869
rect 135 1868 139 1872
rect 175 1868 179 1872
rect 223 1868 227 1872
rect 287 1868 291 1872
rect 359 1868 363 1872
rect 431 1868 435 1872
rect 503 1868 507 1872
rect 567 1868 571 1872
rect 631 1868 635 1872
rect 695 1868 699 1872
rect 759 1868 763 1872
rect 831 1868 835 1872
rect 1095 1865 1099 1869
rect 1135 1859 1139 1863
rect 1231 1856 1235 1860
rect 1271 1856 1275 1860
rect 1319 1856 1323 1860
rect 1375 1856 1379 1860
rect 1439 1856 1443 1860
rect 1503 1856 1507 1860
rect 1575 1856 1579 1860
rect 1655 1856 1659 1860
rect 1751 1856 1755 1860
rect 1863 1856 1867 1860
rect 1975 1856 1979 1860
rect 2071 1856 2075 1860
rect 2119 1859 2123 1863
rect 111 1848 115 1852
rect 1095 1848 1099 1852
rect 135 1840 139 1844
rect 175 1840 179 1844
rect 223 1840 227 1844
rect 287 1840 291 1844
rect 359 1840 363 1844
rect 431 1840 435 1844
rect 503 1840 507 1844
rect 567 1840 571 1844
rect 631 1840 635 1844
rect 695 1840 699 1844
rect 759 1840 763 1844
rect 831 1840 835 1844
rect 1135 1837 1139 1841
rect 1159 1840 1163 1844
rect 1199 1840 1203 1844
rect 1239 1840 1243 1844
rect 1303 1840 1307 1844
rect 1367 1840 1371 1844
rect 1431 1840 1435 1844
rect 1503 1840 1507 1844
rect 1583 1840 1587 1844
rect 1671 1840 1675 1844
rect 1767 1840 1771 1844
rect 1871 1840 1875 1844
rect 1983 1840 1987 1844
rect 2071 1840 2075 1844
rect 2119 1837 2123 1841
rect 1135 1820 1139 1824
rect 2119 1820 2123 1824
rect 1159 1812 1163 1816
rect 1199 1812 1203 1816
rect 1239 1812 1243 1816
rect 1303 1812 1307 1816
rect 1367 1812 1371 1816
rect 1431 1812 1435 1816
rect 1503 1812 1507 1816
rect 1583 1812 1587 1816
rect 1671 1812 1675 1816
rect 1767 1812 1771 1816
rect 1871 1812 1875 1816
rect 1983 1812 1987 1816
rect 2071 1812 2075 1816
rect 135 1800 139 1804
rect 183 1800 187 1804
rect 263 1800 267 1804
rect 351 1800 355 1804
rect 439 1800 443 1804
rect 527 1800 531 1804
rect 607 1800 611 1804
rect 687 1800 691 1804
rect 767 1800 771 1804
rect 839 1800 843 1804
rect 911 1800 915 1804
rect 991 1800 995 1804
rect 1047 1800 1051 1804
rect 111 1792 115 1796
rect 1095 1792 1099 1796
rect 111 1775 115 1779
rect 135 1772 139 1776
rect 183 1772 187 1776
rect 263 1772 267 1776
rect 351 1772 355 1776
rect 439 1772 443 1776
rect 527 1772 531 1776
rect 607 1772 611 1776
rect 687 1772 691 1776
rect 767 1772 771 1776
rect 839 1772 843 1776
rect 911 1772 915 1776
rect 991 1772 995 1776
rect 1047 1772 1051 1776
rect 1095 1775 1099 1779
rect 1311 1768 1315 1772
rect 1351 1768 1355 1772
rect 1391 1768 1395 1772
rect 1431 1768 1435 1772
rect 1471 1768 1475 1772
rect 1511 1768 1515 1772
rect 1551 1768 1555 1772
rect 1607 1768 1611 1772
rect 1679 1768 1683 1772
rect 1767 1768 1771 1772
rect 1871 1768 1875 1772
rect 1983 1768 1987 1772
rect 2071 1768 2075 1772
rect 1135 1760 1139 1764
rect 2119 1760 2123 1764
rect 111 1749 115 1753
rect 135 1752 139 1756
rect 199 1752 203 1756
rect 295 1752 299 1756
rect 399 1752 403 1756
rect 495 1752 499 1756
rect 591 1752 595 1756
rect 671 1752 675 1756
rect 751 1752 755 1756
rect 823 1752 827 1756
rect 887 1752 891 1756
rect 959 1752 963 1756
rect 1031 1752 1035 1756
rect 1095 1749 1099 1753
rect 1135 1743 1139 1747
rect 1311 1740 1315 1744
rect 1351 1740 1355 1744
rect 1391 1740 1395 1744
rect 1431 1740 1435 1744
rect 1471 1740 1475 1744
rect 1511 1740 1515 1744
rect 1551 1740 1555 1744
rect 1607 1740 1611 1744
rect 1679 1740 1683 1744
rect 1767 1740 1771 1744
rect 1871 1740 1875 1744
rect 1983 1740 1987 1744
rect 2071 1740 2075 1744
rect 2119 1743 2123 1747
rect 111 1732 115 1736
rect 1095 1732 1099 1736
rect 135 1724 139 1728
rect 199 1724 203 1728
rect 295 1724 299 1728
rect 399 1724 403 1728
rect 495 1724 499 1728
rect 591 1724 595 1728
rect 671 1724 675 1728
rect 751 1724 755 1728
rect 823 1724 827 1728
rect 887 1724 891 1728
rect 959 1724 963 1728
rect 1031 1724 1035 1728
rect 1135 1721 1139 1725
rect 1263 1724 1267 1728
rect 1319 1724 1323 1728
rect 1383 1724 1387 1728
rect 1455 1724 1459 1728
rect 1535 1724 1539 1728
rect 1615 1724 1619 1728
rect 1687 1724 1691 1728
rect 1759 1724 1763 1728
rect 1831 1724 1835 1728
rect 1895 1724 1899 1728
rect 1959 1724 1963 1728
rect 2023 1724 2027 1728
rect 2071 1724 2075 1728
rect 2119 1721 2123 1725
rect 1135 1704 1139 1708
rect 2119 1704 2123 1708
rect 1263 1696 1267 1700
rect 1319 1696 1323 1700
rect 1383 1696 1387 1700
rect 1455 1696 1459 1700
rect 1535 1696 1539 1700
rect 1615 1696 1619 1700
rect 1687 1696 1691 1700
rect 1759 1696 1763 1700
rect 1831 1696 1835 1700
rect 1895 1696 1899 1700
rect 1959 1696 1963 1700
rect 2023 1696 2027 1700
rect 2071 1696 2075 1700
rect 151 1684 155 1688
rect 223 1684 227 1688
rect 303 1684 307 1688
rect 383 1684 387 1688
rect 463 1684 467 1688
rect 535 1684 539 1688
rect 607 1684 611 1688
rect 671 1684 675 1688
rect 735 1684 739 1688
rect 807 1684 811 1688
rect 879 1684 883 1688
rect 111 1676 115 1680
rect 1095 1676 1099 1680
rect 111 1659 115 1663
rect 151 1656 155 1660
rect 223 1656 227 1660
rect 303 1656 307 1660
rect 383 1656 387 1660
rect 463 1656 467 1660
rect 535 1656 539 1660
rect 607 1656 611 1660
rect 671 1656 675 1660
rect 735 1656 739 1660
rect 807 1656 811 1660
rect 879 1656 883 1660
rect 1095 1659 1099 1663
rect 1167 1660 1171 1664
rect 1247 1660 1251 1664
rect 1335 1660 1339 1664
rect 1423 1660 1427 1664
rect 1511 1660 1515 1664
rect 1599 1660 1603 1664
rect 1679 1660 1683 1664
rect 1751 1660 1755 1664
rect 1815 1660 1819 1664
rect 1871 1660 1875 1664
rect 1927 1660 1931 1664
rect 1983 1660 1987 1664
rect 2031 1660 2035 1664
rect 2071 1660 2075 1664
rect 1135 1652 1139 1656
rect 2119 1652 2123 1656
rect 111 1637 115 1641
rect 175 1640 179 1644
rect 215 1640 219 1644
rect 255 1640 259 1644
rect 303 1640 307 1644
rect 359 1640 363 1644
rect 407 1640 411 1644
rect 455 1640 459 1644
rect 503 1640 507 1644
rect 551 1640 555 1644
rect 607 1640 611 1644
rect 663 1640 667 1644
rect 719 1640 723 1644
rect 1095 1637 1099 1641
rect 1135 1635 1139 1639
rect 1167 1632 1171 1636
rect 1247 1632 1251 1636
rect 1335 1632 1339 1636
rect 1423 1632 1427 1636
rect 1511 1632 1515 1636
rect 1599 1632 1603 1636
rect 1679 1632 1683 1636
rect 1751 1632 1755 1636
rect 1815 1632 1819 1636
rect 1871 1632 1875 1636
rect 1927 1632 1931 1636
rect 1983 1632 1987 1636
rect 2031 1632 2035 1636
rect 2071 1632 2075 1636
rect 2119 1635 2123 1639
rect 111 1620 115 1624
rect 1095 1620 1099 1624
rect 175 1612 179 1616
rect 215 1612 219 1616
rect 255 1612 259 1616
rect 303 1612 307 1616
rect 359 1612 363 1616
rect 407 1612 411 1616
rect 455 1612 459 1616
rect 503 1612 507 1616
rect 551 1612 555 1616
rect 607 1612 611 1616
rect 663 1612 667 1616
rect 719 1612 723 1616
rect 1135 1613 1139 1617
rect 1159 1616 1163 1620
rect 1199 1616 1203 1620
rect 1247 1616 1251 1620
rect 1319 1616 1323 1620
rect 1391 1616 1395 1620
rect 1463 1616 1467 1620
rect 1535 1616 1539 1620
rect 1607 1616 1611 1620
rect 1679 1616 1683 1620
rect 1751 1616 1755 1620
rect 1831 1616 1835 1620
rect 2119 1613 2123 1617
rect 1135 1596 1139 1600
rect 2119 1596 2123 1600
rect 1159 1588 1163 1592
rect 1199 1588 1203 1592
rect 1247 1588 1251 1592
rect 1319 1588 1323 1592
rect 1391 1588 1395 1592
rect 1463 1588 1467 1592
rect 1535 1588 1539 1592
rect 1607 1588 1611 1592
rect 1679 1588 1683 1592
rect 1751 1588 1755 1592
rect 1831 1588 1835 1592
rect 143 1568 147 1572
rect 183 1568 187 1572
rect 231 1568 235 1572
rect 287 1568 291 1572
rect 351 1568 355 1572
rect 415 1568 419 1572
rect 479 1568 483 1572
rect 543 1568 547 1572
rect 607 1568 611 1572
rect 663 1568 667 1572
rect 727 1568 731 1572
rect 791 1568 795 1572
rect 855 1568 859 1572
rect 111 1560 115 1564
rect 1095 1560 1099 1564
rect 1239 1552 1243 1556
rect 1279 1552 1283 1556
rect 1327 1552 1331 1556
rect 1375 1552 1379 1556
rect 1423 1552 1427 1556
rect 1471 1552 1475 1556
rect 1519 1552 1523 1556
rect 1567 1552 1571 1556
rect 1623 1552 1627 1556
rect 1679 1552 1683 1556
rect 1735 1552 1739 1556
rect 111 1543 115 1547
rect 143 1540 147 1544
rect 183 1540 187 1544
rect 231 1540 235 1544
rect 287 1540 291 1544
rect 351 1540 355 1544
rect 415 1540 419 1544
rect 479 1540 483 1544
rect 543 1540 547 1544
rect 607 1540 611 1544
rect 663 1540 667 1544
rect 727 1540 731 1544
rect 791 1540 795 1544
rect 855 1540 859 1544
rect 1095 1543 1099 1547
rect 1135 1544 1139 1548
rect 2119 1544 2123 1548
rect 1135 1527 1139 1531
rect 111 1517 115 1521
rect 135 1520 139 1524
rect 175 1520 179 1524
rect 215 1520 219 1524
rect 255 1520 259 1524
rect 295 1520 299 1524
rect 335 1520 339 1524
rect 375 1520 379 1524
rect 415 1520 419 1524
rect 455 1520 459 1524
rect 495 1520 499 1524
rect 535 1520 539 1524
rect 575 1520 579 1524
rect 615 1520 619 1524
rect 655 1520 659 1524
rect 695 1520 699 1524
rect 735 1520 739 1524
rect 775 1520 779 1524
rect 831 1520 835 1524
rect 887 1520 891 1524
rect 1239 1524 1243 1528
rect 1279 1524 1283 1528
rect 1327 1524 1331 1528
rect 1375 1524 1379 1528
rect 1423 1524 1427 1528
rect 1471 1524 1475 1528
rect 1519 1524 1523 1528
rect 1567 1524 1571 1528
rect 1623 1524 1627 1528
rect 1679 1524 1683 1528
rect 1735 1524 1739 1528
rect 2119 1527 2123 1531
rect 1095 1517 1099 1521
rect 1135 1505 1139 1509
rect 1319 1508 1323 1512
rect 1359 1508 1363 1512
rect 1399 1508 1403 1512
rect 1439 1508 1443 1512
rect 1479 1508 1483 1512
rect 1519 1508 1523 1512
rect 1559 1508 1563 1512
rect 1607 1508 1611 1512
rect 1663 1508 1667 1512
rect 1735 1508 1739 1512
rect 1815 1508 1819 1512
rect 1903 1508 1907 1512
rect 1991 1508 1995 1512
rect 2071 1508 2075 1512
rect 111 1500 115 1504
rect 2119 1505 2123 1509
rect 1095 1500 1099 1504
rect 135 1492 139 1496
rect 175 1492 179 1496
rect 215 1492 219 1496
rect 255 1492 259 1496
rect 295 1492 299 1496
rect 335 1492 339 1496
rect 375 1492 379 1496
rect 415 1492 419 1496
rect 455 1492 459 1496
rect 495 1492 499 1496
rect 535 1492 539 1496
rect 575 1492 579 1496
rect 615 1492 619 1496
rect 655 1492 659 1496
rect 695 1492 699 1496
rect 735 1492 739 1496
rect 775 1492 779 1496
rect 831 1492 835 1496
rect 887 1492 891 1496
rect 1135 1488 1139 1492
rect 2119 1488 2123 1492
rect 1319 1480 1323 1484
rect 1359 1480 1363 1484
rect 1399 1480 1403 1484
rect 1439 1480 1443 1484
rect 1479 1480 1483 1484
rect 1519 1480 1523 1484
rect 1559 1480 1563 1484
rect 1607 1480 1611 1484
rect 1663 1480 1667 1484
rect 1735 1480 1739 1484
rect 1815 1480 1819 1484
rect 1903 1480 1907 1484
rect 1991 1480 1995 1484
rect 2071 1480 2075 1484
rect 519 1448 523 1452
rect 559 1448 563 1452
rect 599 1448 603 1452
rect 647 1448 651 1452
rect 695 1448 699 1452
rect 751 1448 755 1452
rect 807 1448 811 1452
rect 871 1448 875 1452
rect 935 1448 939 1452
rect 111 1440 115 1444
rect 1095 1440 1099 1444
rect 1231 1444 1235 1448
rect 1279 1444 1283 1448
rect 1335 1444 1339 1448
rect 1391 1444 1395 1448
rect 1455 1444 1459 1448
rect 1519 1444 1523 1448
rect 1583 1444 1587 1448
rect 1647 1444 1651 1448
rect 1719 1444 1723 1448
rect 1807 1444 1811 1448
rect 1895 1444 1899 1448
rect 1991 1444 1995 1448
rect 2071 1444 2075 1448
rect 1135 1436 1139 1440
rect 2119 1436 2123 1440
rect 111 1423 115 1427
rect 519 1420 523 1424
rect 559 1420 563 1424
rect 599 1420 603 1424
rect 647 1420 651 1424
rect 695 1420 699 1424
rect 751 1420 755 1424
rect 807 1420 811 1424
rect 871 1420 875 1424
rect 935 1420 939 1424
rect 1095 1423 1099 1427
rect 1135 1419 1139 1423
rect 1231 1416 1235 1420
rect 1279 1416 1283 1420
rect 1335 1416 1339 1420
rect 1391 1416 1395 1420
rect 1455 1416 1459 1420
rect 1519 1416 1523 1420
rect 1583 1416 1587 1420
rect 1647 1416 1651 1420
rect 1719 1416 1723 1420
rect 1807 1416 1811 1420
rect 1895 1416 1899 1420
rect 1991 1416 1995 1420
rect 2071 1416 2075 1420
rect 2119 1419 2123 1423
rect 111 1401 115 1405
rect 431 1404 435 1408
rect 471 1404 475 1408
rect 519 1404 523 1408
rect 575 1404 579 1408
rect 631 1404 635 1408
rect 695 1404 699 1408
rect 759 1404 763 1408
rect 823 1404 827 1408
rect 895 1404 899 1408
rect 967 1404 971 1408
rect 1095 1401 1099 1405
rect 1135 1397 1139 1401
rect 1159 1400 1163 1404
rect 1199 1400 1203 1404
rect 1263 1400 1267 1404
rect 1351 1400 1355 1404
rect 1447 1400 1451 1404
rect 1543 1400 1547 1404
rect 1631 1400 1635 1404
rect 1719 1400 1723 1404
rect 1799 1400 1803 1404
rect 1871 1400 1875 1404
rect 1943 1400 1947 1404
rect 2015 1400 2019 1404
rect 2071 1400 2075 1404
rect 2119 1397 2123 1401
rect 111 1384 115 1388
rect 1095 1384 1099 1388
rect 431 1376 435 1380
rect 471 1376 475 1380
rect 519 1376 523 1380
rect 575 1376 579 1380
rect 631 1376 635 1380
rect 695 1376 699 1380
rect 759 1376 763 1380
rect 823 1376 827 1380
rect 895 1376 899 1380
rect 967 1376 971 1380
rect 1135 1380 1139 1384
rect 2119 1380 2123 1384
rect 1159 1372 1163 1376
rect 1199 1372 1203 1376
rect 1263 1372 1267 1376
rect 1351 1372 1355 1376
rect 1447 1372 1451 1376
rect 1543 1372 1547 1376
rect 1631 1372 1635 1376
rect 1719 1372 1723 1376
rect 1799 1372 1803 1376
rect 1871 1372 1875 1376
rect 1943 1372 1947 1376
rect 2015 1372 2019 1376
rect 2071 1372 2075 1376
rect 375 1340 379 1344
rect 423 1340 427 1344
rect 479 1340 483 1344
rect 543 1340 547 1344
rect 607 1340 611 1344
rect 671 1340 675 1344
rect 735 1340 739 1344
rect 799 1340 803 1344
rect 863 1340 867 1344
rect 927 1340 931 1344
rect 999 1340 1003 1344
rect 1047 1340 1051 1344
rect 111 1332 115 1336
rect 1095 1332 1099 1336
rect 1159 1332 1163 1336
rect 1255 1332 1259 1336
rect 1375 1332 1379 1336
rect 1487 1332 1491 1336
rect 1591 1332 1595 1336
rect 1679 1332 1683 1336
rect 1759 1332 1763 1336
rect 1831 1332 1835 1336
rect 1903 1332 1907 1336
rect 1967 1332 1971 1336
rect 2031 1332 2035 1336
rect 2071 1332 2075 1336
rect 1135 1324 1139 1328
rect 2119 1324 2123 1328
rect 111 1315 115 1319
rect 375 1312 379 1316
rect 423 1312 427 1316
rect 479 1312 483 1316
rect 543 1312 547 1316
rect 607 1312 611 1316
rect 671 1312 675 1316
rect 735 1312 739 1316
rect 799 1312 803 1316
rect 863 1312 867 1316
rect 927 1312 931 1316
rect 999 1312 1003 1316
rect 1047 1312 1051 1316
rect 1095 1315 1099 1319
rect 1135 1307 1139 1311
rect 111 1297 115 1301
rect 335 1300 339 1304
rect 391 1300 395 1304
rect 455 1300 459 1304
rect 527 1300 531 1304
rect 599 1300 603 1304
rect 671 1300 675 1304
rect 743 1300 747 1304
rect 823 1300 827 1304
rect 903 1300 907 1304
rect 983 1300 987 1304
rect 1047 1300 1051 1304
rect 1159 1304 1163 1308
rect 1255 1304 1259 1308
rect 1375 1304 1379 1308
rect 1487 1304 1491 1308
rect 1591 1304 1595 1308
rect 1679 1304 1683 1308
rect 1759 1304 1763 1308
rect 1831 1304 1835 1308
rect 1903 1304 1907 1308
rect 1967 1304 1971 1308
rect 2031 1304 2035 1308
rect 2071 1304 2075 1308
rect 2119 1307 2123 1311
rect 1095 1297 1099 1301
rect 1135 1285 1139 1289
rect 1159 1288 1163 1292
rect 1199 1288 1203 1292
rect 1247 1288 1251 1292
rect 1319 1288 1323 1292
rect 1399 1288 1403 1292
rect 1479 1288 1483 1292
rect 1559 1288 1563 1292
rect 1639 1288 1643 1292
rect 1719 1288 1723 1292
rect 1799 1288 1803 1292
rect 1879 1288 1883 1292
rect 1967 1288 1971 1292
rect 2055 1288 2059 1292
rect 111 1280 115 1284
rect 2119 1285 2123 1289
rect 1095 1280 1099 1284
rect 335 1272 339 1276
rect 391 1272 395 1276
rect 455 1272 459 1276
rect 527 1272 531 1276
rect 599 1272 603 1276
rect 671 1272 675 1276
rect 743 1272 747 1276
rect 823 1272 827 1276
rect 903 1272 907 1276
rect 983 1272 987 1276
rect 1047 1272 1051 1276
rect 1135 1268 1139 1272
rect 2119 1268 2123 1272
rect 1159 1260 1163 1264
rect 1199 1260 1203 1264
rect 1247 1260 1251 1264
rect 1319 1260 1323 1264
rect 1399 1260 1403 1264
rect 1479 1260 1483 1264
rect 1559 1260 1563 1264
rect 1639 1260 1643 1264
rect 1719 1260 1723 1264
rect 1799 1260 1803 1264
rect 1879 1260 1883 1264
rect 1967 1260 1971 1264
rect 2055 1260 2059 1264
rect 263 1232 267 1236
rect 311 1232 315 1236
rect 359 1232 363 1236
rect 415 1232 419 1236
rect 479 1232 483 1236
rect 543 1232 547 1236
rect 607 1232 611 1236
rect 671 1232 675 1236
rect 735 1232 739 1236
rect 799 1232 803 1236
rect 863 1232 867 1236
rect 927 1232 931 1236
rect 111 1224 115 1228
rect 1095 1224 1099 1228
rect 1159 1220 1163 1224
rect 1199 1220 1203 1224
rect 1239 1220 1243 1224
rect 1279 1220 1283 1224
rect 1327 1220 1331 1224
rect 1375 1220 1379 1224
rect 1423 1220 1427 1224
rect 1471 1220 1475 1224
rect 1535 1220 1539 1224
rect 1615 1220 1619 1224
rect 1719 1220 1723 1224
rect 1839 1220 1843 1224
rect 1967 1220 1971 1224
rect 2071 1220 2075 1224
rect 1135 1212 1139 1216
rect 111 1207 115 1211
rect 2119 1212 2123 1216
rect 263 1204 267 1208
rect 311 1204 315 1208
rect 359 1204 363 1208
rect 415 1204 419 1208
rect 479 1204 483 1208
rect 543 1204 547 1208
rect 607 1204 611 1208
rect 671 1204 675 1208
rect 735 1204 739 1208
rect 799 1204 803 1208
rect 863 1204 867 1208
rect 927 1204 931 1208
rect 1095 1207 1099 1211
rect 111 1189 115 1193
rect 223 1192 227 1196
rect 279 1192 283 1196
rect 343 1192 347 1196
rect 407 1192 411 1196
rect 479 1192 483 1196
rect 551 1192 555 1196
rect 631 1192 635 1196
rect 711 1192 715 1196
rect 791 1192 795 1196
rect 871 1192 875 1196
rect 959 1192 963 1196
rect 1135 1195 1139 1199
rect 1095 1189 1099 1193
rect 1159 1192 1163 1196
rect 1199 1192 1203 1196
rect 1239 1192 1243 1196
rect 1279 1192 1283 1196
rect 1327 1192 1331 1196
rect 1375 1192 1379 1196
rect 1423 1192 1427 1196
rect 1471 1192 1475 1196
rect 1535 1192 1539 1196
rect 1615 1192 1619 1196
rect 1719 1192 1723 1196
rect 1839 1192 1843 1196
rect 1967 1192 1971 1196
rect 2071 1192 2075 1196
rect 2119 1195 2123 1199
rect 1135 1177 1139 1181
rect 1287 1180 1291 1184
rect 1327 1180 1331 1184
rect 1367 1180 1371 1184
rect 1415 1180 1419 1184
rect 1471 1180 1475 1184
rect 1527 1180 1531 1184
rect 1583 1180 1587 1184
rect 1639 1180 1643 1184
rect 1703 1180 1707 1184
rect 1767 1180 1771 1184
rect 1839 1180 1843 1184
rect 1919 1180 1923 1184
rect 2007 1180 2011 1184
rect 2071 1180 2075 1184
rect 111 1172 115 1176
rect 2119 1177 2123 1181
rect 1095 1172 1099 1176
rect 223 1164 227 1168
rect 279 1164 283 1168
rect 343 1164 347 1168
rect 407 1164 411 1168
rect 479 1164 483 1168
rect 551 1164 555 1168
rect 631 1164 635 1168
rect 711 1164 715 1168
rect 791 1164 795 1168
rect 871 1164 875 1168
rect 959 1164 963 1168
rect 1135 1160 1139 1164
rect 2119 1160 2123 1164
rect 1287 1152 1291 1156
rect 1327 1152 1331 1156
rect 1367 1152 1371 1156
rect 1415 1152 1419 1156
rect 1471 1152 1475 1156
rect 1527 1152 1531 1156
rect 1583 1152 1587 1156
rect 1639 1152 1643 1156
rect 1703 1152 1707 1156
rect 1767 1152 1771 1156
rect 1839 1152 1843 1156
rect 1919 1152 1923 1156
rect 2007 1152 2011 1156
rect 2071 1152 2075 1156
rect 159 1128 163 1132
rect 199 1128 203 1132
rect 247 1128 251 1132
rect 303 1128 307 1132
rect 367 1128 371 1132
rect 439 1128 443 1132
rect 511 1128 515 1132
rect 591 1128 595 1132
rect 679 1128 683 1132
rect 775 1128 779 1132
rect 879 1128 883 1132
rect 991 1128 995 1132
rect 111 1120 115 1124
rect 1095 1120 1099 1124
rect 1383 1108 1387 1112
rect 111 1103 115 1107
rect 1423 1108 1427 1112
rect 1471 1108 1475 1112
rect 1527 1108 1531 1112
rect 1591 1108 1595 1112
rect 1655 1108 1659 1112
rect 1711 1108 1715 1112
rect 1767 1108 1771 1112
rect 1823 1108 1827 1112
rect 1871 1108 1875 1112
rect 1927 1108 1931 1112
rect 1983 1108 1987 1112
rect 2031 1108 2035 1112
rect 2071 1108 2075 1112
rect 159 1100 163 1104
rect 199 1100 203 1104
rect 247 1100 251 1104
rect 303 1100 307 1104
rect 367 1100 371 1104
rect 439 1100 443 1104
rect 511 1100 515 1104
rect 591 1100 595 1104
rect 679 1100 683 1104
rect 775 1100 779 1104
rect 879 1100 883 1104
rect 991 1100 995 1104
rect 1095 1103 1099 1107
rect 1135 1100 1139 1104
rect 2119 1100 2123 1104
rect 111 1077 115 1081
rect 199 1080 203 1084
rect 247 1080 251 1084
rect 303 1080 307 1084
rect 367 1080 371 1084
rect 431 1080 435 1084
rect 503 1080 507 1084
rect 575 1080 579 1084
rect 647 1080 651 1084
rect 719 1080 723 1084
rect 783 1080 787 1084
rect 839 1080 843 1084
rect 895 1080 899 1084
rect 951 1080 955 1084
rect 1007 1080 1011 1084
rect 1047 1080 1051 1084
rect 1135 1083 1139 1087
rect 1095 1077 1099 1081
rect 1383 1080 1387 1084
rect 1423 1080 1427 1084
rect 1471 1080 1475 1084
rect 1527 1080 1531 1084
rect 1591 1080 1595 1084
rect 1655 1080 1659 1084
rect 1711 1080 1715 1084
rect 1767 1080 1771 1084
rect 1823 1080 1827 1084
rect 1871 1080 1875 1084
rect 1927 1080 1931 1084
rect 1983 1080 1987 1084
rect 2031 1080 2035 1084
rect 2071 1080 2075 1084
rect 2119 1083 2123 1087
rect 1135 1065 1139 1069
rect 1159 1068 1163 1072
rect 1247 1068 1251 1072
rect 1359 1068 1363 1072
rect 1471 1068 1475 1072
rect 1575 1068 1579 1072
rect 1671 1068 1675 1072
rect 1759 1068 1763 1072
rect 1847 1068 1851 1072
rect 1927 1068 1931 1072
rect 2007 1068 2011 1072
rect 2071 1068 2075 1072
rect 111 1060 115 1064
rect 2119 1065 2123 1069
rect 1095 1060 1099 1064
rect 199 1052 203 1056
rect 247 1052 251 1056
rect 303 1052 307 1056
rect 367 1052 371 1056
rect 431 1052 435 1056
rect 503 1052 507 1056
rect 575 1052 579 1056
rect 647 1052 651 1056
rect 719 1052 723 1056
rect 783 1052 787 1056
rect 839 1052 843 1056
rect 895 1052 899 1056
rect 951 1052 955 1056
rect 1007 1052 1011 1056
rect 1047 1052 1051 1056
rect 1135 1048 1139 1052
rect 2119 1048 2123 1052
rect 1159 1040 1163 1044
rect 1247 1040 1251 1044
rect 1359 1040 1363 1044
rect 1471 1040 1475 1044
rect 1575 1040 1579 1044
rect 1671 1040 1675 1044
rect 1759 1040 1763 1044
rect 1847 1040 1851 1044
rect 1927 1040 1931 1044
rect 2007 1040 2011 1044
rect 2071 1040 2075 1044
rect 223 1012 227 1016
rect 271 1012 275 1016
rect 335 1012 339 1016
rect 407 1012 411 1016
rect 479 1012 483 1016
rect 559 1012 563 1016
rect 631 1012 635 1016
rect 703 1012 707 1016
rect 775 1012 779 1016
rect 839 1012 843 1016
rect 903 1012 907 1016
rect 967 1012 971 1016
rect 1039 1012 1043 1016
rect 111 1004 115 1008
rect 1095 1004 1099 1008
rect 1159 1004 1163 1008
rect 1231 1004 1235 1008
rect 1303 1004 1307 1008
rect 1383 1004 1387 1008
rect 1463 1004 1467 1008
rect 1543 1004 1547 1008
rect 1623 1004 1627 1008
rect 1695 1004 1699 1008
rect 1759 1004 1763 1008
rect 1823 1004 1827 1008
rect 1887 1004 1891 1008
rect 1951 1004 1955 1008
rect 1135 996 1139 1000
rect 2119 996 2123 1000
rect 111 987 115 991
rect 223 984 227 988
rect 271 984 275 988
rect 335 984 339 988
rect 407 984 411 988
rect 479 984 483 988
rect 559 984 563 988
rect 631 984 635 988
rect 703 984 707 988
rect 775 984 779 988
rect 839 984 843 988
rect 903 984 907 988
rect 967 984 971 988
rect 1039 984 1043 988
rect 1095 987 1099 991
rect 1135 979 1139 983
rect 1159 976 1163 980
rect 1231 976 1235 980
rect 1303 976 1307 980
rect 1383 976 1387 980
rect 1463 976 1467 980
rect 1543 976 1547 980
rect 1623 976 1627 980
rect 1695 976 1699 980
rect 1759 976 1763 980
rect 1823 976 1827 980
rect 1887 976 1891 980
rect 1951 976 1955 980
rect 2119 979 2123 983
rect 111 965 115 969
rect 151 968 155 972
rect 215 968 219 972
rect 287 968 291 972
rect 367 968 371 972
rect 447 968 451 972
rect 527 968 531 972
rect 599 968 603 972
rect 671 968 675 972
rect 735 968 739 972
rect 799 968 803 972
rect 863 968 867 972
rect 927 968 931 972
rect 991 968 995 972
rect 1047 968 1051 972
rect 1095 965 1099 969
rect 1135 961 1139 965
rect 1239 964 1243 968
rect 1303 964 1307 968
rect 1375 964 1379 968
rect 1439 964 1443 968
rect 1511 964 1515 968
rect 1583 964 1587 968
rect 1655 964 1659 968
rect 1727 964 1731 968
rect 1799 964 1803 968
rect 1871 964 1875 968
rect 1943 964 1947 968
rect 2015 964 2019 968
rect 2071 964 2075 968
rect 2119 961 2123 965
rect 111 948 115 952
rect 1095 948 1099 952
rect 151 940 155 944
rect 215 940 219 944
rect 287 940 291 944
rect 367 940 371 944
rect 447 940 451 944
rect 527 940 531 944
rect 599 940 603 944
rect 671 940 675 944
rect 735 940 739 944
rect 799 940 803 944
rect 863 940 867 944
rect 927 940 931 944
rect 991 940 995 944
rect 1047 940 1051 944
rect 1135 944 1139 948
rect 2119 944 2123 948
rect 1239 936 1243 940
rect 1303 936 1307 940
rect 1375 936 1379 940
rect 1439 936 1443 940
rect 1511 936 1515 940
rect 1583 936 1587 940
rect 1655 936 1659 940
rect 1727 936 1731 940
rect 1799 936 1803 940
rect 1871 936 1875 940
rect 1943 936 1947 940
rect 2015 936 2019 940
rect 2071 936 2075 940
rect 135 904 139 908
rect 183 904 187 908
rect 255 904 259 908
rect 327 904 331 908
rect 399 904 403 908
rect 463 904 467 908
rect 527 904 531 908
rect 599 904 603 908
rect 671 904 675 908
rect 743 904 747 908
rect 815 904 819 908
rect 895 904 899 908
rect 983 904 987 908
rect 1047 904 1051 908
rect 111 896 115 900
rect 1095 896 1099 900
rect 1287 896 1291 900
rect 1327 896 1331 900
rect 1375 896 1379 900
rect 1423 896 1427 900
rect 1479 896 1483 900
rect 1551 896 1555 900
rect 1623 896 1627 900
rect 1703 896 1707 900
rect 1791 896 1795 900
rect 1879 896 1883 900
rect 1967 896 1971 900
rect 2063 896 2067 900
rect 1135 888 1139 892
rect 2119 888 2123 892
rect 111 879 115 883
rect 135 876 139 880
rect 183 876 187 880
rect 255 876 259 880
rect 327 876 331 880
rect 399 876 403 880
rect 463 876 467 880
rect 527 876 531 880
rect 599 876 603 880
rect 671 876 675 880
rect 743 876 747 880
rect 815 876 819 880
rect 895 876 899 880
rect 983 876 987 880
rect 1047 876 1051 880
rect 1095 879 1099 883
rect 1135 871 1139 875
rect 1287 868 1291 872
rect 1327 868 1331 872
rect 1375 868 1379 872
rect 1423 868 1427 872
rect 1479 868 1483 872
rect 1551 868 1555 872
rect 1623 868 1627 872
rect 1703 868 1707 872
rect 1791 868 1795 872
rect 1879 868 1883 872
rect 1967 868 1971 872
rect 2063 868 2067 872
rect 2119 871 2123 875
rect 111 857 115 861
rect 135 860 139 864
rect 175 860 179 864
rect 215 860 219 864
rect 279 860 283 864
rect 343 860 347 864
rect 399 860 403 864
rect 463 860 467 864
rect 535 860 539 864
rect 615 860 619 864
rect 711 860 715 864
rect 823 860 827 864
rect 943 860 947 864
rect 1047 860 1051 864
rect 1095 857 1099 861
rect 1135 853 1139 857
rect 1159 856 1163 860
rect 1199 856 1203 860
rect 1263 856 1267 860
rect 1327 856 1331 860
rect 1399 856 1403 860
rect 1471 856 1475 860
rect 1543 856 1547 860
rect 1623 856 1627 860
rect 1703 856 1707 860
rect 1775 856 1779 860
rect 1855 856 1859 860
rect 1935 856 1939 860
rect 2015 856 2019 860
rect 2071 856 2075 860
rect 2119 853 2123 857
rect 111 840 115 844
rect 1095 840 1099 844
rect 135 832 139 836
rect 175 832 179 836
rect 215 832 219 836
rect 279 832 283 836
rect 343 832 347 836
rect 399 832 403 836
rect 463 832 467 836
rect 535 832 539 836
rect 615 832 619 836
rect 711 832 715 836
rect 823 832 827 836
rect 943 832 947 836
rect 1047 832 1051 836
rect 1135 836 1139 840
rect 2119 836 2123 840
rect 1159 828 1163 832
rect 1199 828 1203 832
rect 1263 828 1267 832
rect 1327 828 1331 832
rect 1399 828 1403 832
rect 1471 828 1475 832
rect 1543 828 1547 832
rect 1623 828 1627 832
rect 1703 828 1707 832
rect 1775 828 1779 832
rect 1855 828 1859 832
rect 1935 828 1939 832
rect 2015 828 2019 832
rect 2071 828 2075 832
rect 135 796 139 800
rect 175 796 179 800
rect 215 796 219 800
rect 279 796 283 800
rect 335 796 339 800
rect 391 796 395 800
rect 455 796 459 800
rect 519 796 523 800
rect 583 796 587 800
rect 655 796 659 800
rect 735 796 739 800
rect 815 796 819 800
rect 895 796 899 800
rect 983 796 987 800
rect 1047 796 1051 800
rect 111 788 115 792
rect 1095 788 1099 792
rect 1159 784 1163 788
rect 1239 784 1243 788
rect 1343 784 1347 788
rect 1447 784 1451 788
rect 1551 784 1555 788
rect 1655 784 1659 788
rect 1751 784 1755 788
rect 1839 784 1843 788
rect 1919 784 1923 788
rect 2007 784 2011 788
rect 2071 784 2075 788
rect 1135 776 1139 780
rect 111 771 115 775
rect 2119 776 2123 780
rect 135 768 139 772
rect 175 768 179 772
rect 215 768 219 772
rect 279 768 283 772
rect 335 768 339 772
rect 391 768 395 772
rect 455 768 459 772
rect 519 768 523 772
rect 583 768 587 772
rect 655 768 659 772
rect 735 768 739 772
rect 815 768 819 772
rect 895 768 899 772
rect 983 768 987 772
rect 1047 768 1051 772
rect 1095 771 1099 775
rect 111 753 115 757
rect 135 756 139 760
rect 207 756 211 760
rect 295 756 299 760
rect 375 756 379 760
rect 447 756 451 760
rect 519 756 523 760
rect 583 756 587 760
rect 639 756 643 760
rect 687 756 691 760
rect 743 756 747 760
rect 799 756 803 760
rect 855 756 859 760
rect 1135 759 1139 763
rect 1095 753 1099 757
rect 1159 756 1163 760
rect 1239 756 1243 760
rect 1343 756 1347 760
rect 1447 756 1451 760
rect 1551 756 1555 760
rect 1655 756 1659 760
rect 1751 756 1755 760
rect 1839 756 1843 760
rect 1919 756 1923 760
rect 2007 756 2011 760
rect 2071 756 2075 760
rect 2119 759 2123 763
rect 1135 741 1139 745
rect 1159 744 1163 748
rect 1199 744 1203 748
rect 1239 744 1243 748
rect 1287 744 1291 748
rect 1359 744 1363 748
rect 1439 744 1443 748
rect 1527 744 1531 748
rect 1615 744 1619 748
rect 1711 744 1715 748
rect 1807 744 1811 748
rect 1903 744 1907 748
rect 1999 744 2003 748
rect 2071 744 2075 748
rect 111 736 115 740
rect 2119 741 2123 745
rect 1095 736 1099 740
rect 135 728 139 732
rect 207 728 211 732
rect 295 728 299 732
rect 375 728 379 732
rect 447 728 451 732
rect 519 728 523 732
rect 583 728 587 732
rect 639 728 643 732
rect 687 728 691 732
rect 743 728 747 732
rect 799 728 803 732
rect 855 728 859 732
rect 1135 724 1139 728
rect 2119 724 2123 728
rect 1159 716 1163 720
rect 1199 716 1203 720
rect 1239 716 1243 720
rect 1287 716 1291 720
rect 1359 716 1363 720
rect 1439 716 1443 720
rect 1527 716 1531 720
rect 1615 716 1619 720
rect 1711 716 1715 720
rect 1807 716 1811 720
rect 1903 716 1907 720
rect 1999 716 2003 720
rect 2071 716 2075 720
rect 135 688 139 692
rect 183 688 187 692
rect 247 688 251 692
rect 311 688 315 692
rect 383 688 387 692
rect 455 688 459 692
rect 519 688 523 692
rect 583 688 587 692
rect 647 688 651 692
rect 711 688 715 692
rect 767 688 771 692
rect 823 688 827 692
rect 879 688 883 692
rect 943 688 947 692
rect 111 680 115 684
rect 1095 680 1099 684
rect 1239 676 1243 680
rect 1287 676 1291 680
rect 1335 676 1339 680
rect 1391 676 1395 680
rect 1447 676 1451 680
rect 1511 676 1515 680
rect 1575 676 1579 680
rect 1639 676 1643 680
rect 1703 676 1707 680
rect 1767 676 1771 680
rect 1831 676 1835 680
rect 1895 676 1899 680
rect 1959 676 1963 680
rect 2023 676 2027 680
rect 2071 676 2075 680
rect 1135 668 1139 672
rect 111 663 115 667
rect 2119 668 2123 672
rect 135 660 139 664
rect 183 660 187 664
rect 247 660 251 664
rect 311 660 315 664
rect 383 660 387 664
rect 455 660 459 664
rect 519 660 523 664
rect 583 660 587 664
rect 647 660 651 664
rect 711 660 715 664
rect 767 660 771 664
rect 823 660 827 664
rect 879 660 883 664
rect 943 660 947 664
rect 1095 663 1099 667
rect 1135 651 1139 655
rect 1239 648 1243 652
rect 1287 648 1291 652
rect 1335 648 1339 652
rect 1391 648 1395 652
rect 1447 648 1451 652
rect 1511 648 1515 652
rect 1575 648 1579 652
rect 1639 648 1643 652
rect 1703 648 1707 652
rect 1767 648 1771 652
rect 1831 648 1835 652
rect 1895 648 1899 652
rect 1959 648 1963 652
rect 2023 648 2027 652
rect 2071 648 2075 652
rect 2119 651 2123 655
rect 111 637 115 641
rect 159 640 163 644
rect 215 640 219 644
rect 287 640 291 644
rect 367 640 371 644
rect 455 640 459 644
rect 543 640 547 644
rect 631 640 635 644
rect 719 640 723 644
rect 799 640 803 644
rect 871 640 875 644
rect 951 640 955 644
rect 1031 640 1035 644
rect 1095 637 1099 641
rect 1135 633 1139 637
rect 1279 636 1283 640
rect 1319 636 1323 640
rect 1367 636 1371 640
rect 1423 636 1427 640
rect 1479 636 1483 640
rect 1535 636 1539 640
rect 1591 636 1595 640
rect 1647 636 1651 640
rect 1719 636 1723 640
rect 1799 636 1803 640
rect 1879 636 1883 640
rect 1967 636 1971 640
rect 2063 636 2067 640
rect 2119 633 2123 637
rect 111 620 115 624
rect 1095 620 1099 624
rect 159 612 163 616
rect 215 612 219 616
rect 287 612 291 616
rect 367 612 371 616
rect 455 612 459 616
rect 543 612 547 616
rect 631 612 635 616
rect 719 612 723 616
rect 799 612 803 616
rect 871 612 875 616
rect 951 612 955 616
rect 1031 612 1035 616
rect 1135 616 1139 620
rect 2119 616 2123 620
rect 1279 608 1283 612
rect 1319 608 1323 612
rect 1367 608 1371 612
rect 1423 608 1427 612
rect 1479 608 1483 612
rect 1535 608 1539 612
rect 1591 608 1595 612
rect 1647 608 1651 612
rect 1719 608 1723 612
rect 1799 608 1803 612
rect 1879 608 1883 612
rect 1967 608 1971 612
rect 2063 608 2067 612
rect 159 572 163 576
rect 207 572 211 576
rect 255 572 259 576
rect 311 572 315 576
rect 383 572 387 576
rect 463 572 467 576
rect 543 572 547 576
rect 623 572 627 576
rect 703 572 707 576
rect 783 572 787 576
rect 855 572 859 576
rect 927 572 931 576
rect 999 572 1003 576
rect 1047 572 1051 576
rect 1335 572 1339 576
rect 1375 572 1379 576
rect 1415 572 1419 576
rect 1463 572 1467 576
rect 1519 572 1523 576
rect 1583 572 1587 576
rect 1655 572 1659 576
rect 1727 572 1731 576
rect 1807 572 1811 576
rect 1887 572 1891 576
rect 1975 572 1979 576
rect 2063 572 2067 576
rect 111 564 115 568
rect 1095 564 1099 568
rect 1135 564 1139 568
rect 2119 564 2123 568
rect 111 547 115 551
rect 159 544 163 548
rect 207 544 211 548
rect 255 544 259 548
rect 311 544 315 548
rect 383 544 387 548
rect 463 544 467 548
rect 543 544 547 548
rect 623 544 627 548
rect 703 544 707 548
rect 783 544 787 548
rect 855 544 859 548
rect 927 544 931 548
rect 999 544 1003 548
rect 1047 544 1051 548
rect 1095 547 1099 551
rect 1135 547 1139 551
rect 1335 544 1339 548
rect 1375 544 1379 548
rect 1415 544 1419 548
rect 1463 544 1467 548
rect 1519 544 1523 548
rect 1583 544 1587 548
rect 1655 544 1659 548
rect 1727 544 1731 548
rect 1807 544 1811 548
rect 1887 544 1891 548
rect 1975 544 1979 548
rect 2063 544 2067 548
rect 2119 547 2123 551
rect 111 521 115 525
rect 167 524 171 528
rect 223 524 227 528
rect 287 524 291 528
rect 359 524 363 528
rect 431 524 435 528
rect 511 524 515 528
rect 591 524 595 528
rect 663 524 667 528
rect 735 524 739 528
rect 807 524 811 528
rect 871 524 875 528
rect 935 524 939 528
rect 999 524 1003 528
rect 1047 524 1051 528
rect 1095 521 1099 525
rect 1135 525 1139 529
rect 1191 528 1195 532
rect 1239 528 1243 532
rect 1287 528 1291 532
rect 1343 528 1347 532
rect 1407 528 1411 532
rect 1479 528 1483 532
rect 1543 528 1547 532
rect 1607 528 1611 532
rect 1671 528 1675 532
rect 1735 528 1739 532
rect 1799 528 1803 532
rect 1863 528 1867 532
rect 1935 528 1939 532
rect 2007 528 2011 532
rect 2071 528 2075 532
rect 2119 525 2123 529
rect 111 504 115 508
rect 1095 504 1099 508
rect 1135 508 1139 512
rect 2119 508 2123 512
rect 167 496 171 500
rect 223 496 227 500
rect 287 496 291 500
rect 359 496 363 500
rect 431 496 435 500
rect 511 496 515 500
rect 591 496 595 500
rect 663 496 667 500
rect 735 496 739 500
rect 807 496 811 500
rect 871 496 875 500
rect 935 496 939 500
rect 999 496 1003 500
rect 1047 496 1051 500
rect 1191 500 1195 504
rect 1239 500 1243 504
rect 1287 500 1291 504
rect 1343 500 1347 504
rect 1407 500 1411 504
rect 1479 500 1483 504
rect 1543 500 1547 504
rect 1607 500 1611 504
rect 1671 500 1675 504
rect 1735 500 1739 504
rect 1799 500 1803 504
rect 1863 500 1867 504
rect 1935 500 1939 504
rect 2007 500 2011 504
rect 2071 500 2075 504
rect 167 460 171 464
rect 231 460 235 464
rect 303 460 307 464
rect 375 460 379 464
rect 455 460 459 464
rect 535 460 539 464
rect 607 460 611 464
rect 679 460 683 464
rect 743 460 747 464
rect 799 460 803 464
rect 855 460 859 464
rect 903 460 907 464
rect 959 460 963 464
rect 1007 460 1011 464
rect 1047 460 1051 464
rect 1159 464 1163 468
rect 1263 464 1267 468
rect 1383 464 1387 468
rect 1495 464 1499 468
rect 1599 464 1603 468
rect 1703 464 1707 468
rect 1799 464 1803 468
rect 1887 464 1891 468
rect 1983 464 1987 468
rect 2071 464 2075 468
rect 111 452 115 456
rect 1095 452 1099 456
rect 1135 456 1139 460
rect 2119 456 2123 460
rect 111 435 115 439
rect 167 432 171 436
rect 231 432 235 436
rect 303 432 307 436
rect 375 432 379 436
rect 455 432 459 436
rect 535 432 539 436
rect 607 432 611 436
rect 679 432 683 436
rect 743 432 747 436
rect 799 432 803 436
rect 855 432 859 436
rect 903 432 907 436
rect 959 432 963 436
rect 1007 432 1011 436
rect 1047 432 1051 436
rect 1095 435 1099 439
rect 1135 439 1139 443
rect 1159 436 1163 440
rect 1263 436 1267 440
rect 1383 436 1387 440
rect 1495 436 1499 440
rect 1599 436 1603 440
rect 1703 436 1707 440
rect 1799 436 1803 440
rect 1887 436 1891 440
rect 1983 436 1987 440
rect 2071 436 2075 440
rect 2119 439 2123 443
rect 111 417 115 421
rect 151 420 155 424
rect 215 420 219 424
rect 279 420 283 424
rect 351 420 355 424
rect 423 420 427 424
rect 487 420 491 424
rect 551 420 555 424
rect 615 420 619 424
rect 671 420 675 424
rect 727 420 731 424
rect 791 420 795 424
rect 855 420 859 424
rect 1095 417 1099 421
rect 1135 421 1139 425
rect 1159 424 1163 428
rect 1199 424 1203 428
rect 1255 424 1259 428
rect 1335 424 1339 428
rect 1415 424 1419 428
rect 1503 424 1507 428
rect 1591 424 1595 428
rect 1671 424 1675 428
rect 1751 424 1755 428
rect 1823 424 1827 428
rect 1887 424 1891 428
rect 1951 424 1955 428
rect 2023 424 2027 428
rect 2071 424 2075 428
rect 2119 421 2123 425
rect 111 400 115 404
rect 1095 400 1099 404
rect 1135 404 1139 408
rect 2119 404 2123 408
rect 151 392 155 396
rect 215 392 219 396
rect 279 392 283 396
rect 351 392 355 396
rect 423 392 427 396
rect 487 392 491 396
rect 551 392 555 396
rect 615 392 619 396
rect 671 392 675 396
rect 727 392 731 396
rect 791 392 795 396
rect 855 392 859 396
rect 1159 396 1163 400
rect 1199 396 1203 400
rect 1255 396 1259 400
rect 1335 396 1339 400
rect 1415 396 1419 400
rect 1503 396 1507 400
rect 1591 396 1595 400
rect 1671 396 1675 400
rect 1751 396 1755 400
rect 1823 396 1827 400
rect 1887 396 1891 400
rect 1951 396 1955 400
rect 2023 396 2027 400
rect 2071 396 2075 400
rect 135 356 139 360
rect 175 356 179 360
rect 215 356 219 360
rect 271 356 275 360
rect 335 356 339 360
rect 399 356 403 360
rect 463 356 467 360
rect 519 356 523 360
rect 575 356 579 360
rect 631 356 635 360
rect 687 356 691 360
rect 751 356 755 360
rect 1303 356 1307 360
rect 1343 356 1347 360
rect 1383 356 1387 360
rect 1423 356 1427 360
rect 1463 356 1467 360
rect 1503 356 1507 360
rect 1551 356 1555 360
rect 1615 356 1619 360
rect 1679 356 1683 360
rect 1751 356 1755 360
rect 1831 356 1835 360
rect 1919 356 1923 360
rect 2007 356 2011 360
rect 2071 356 2075 360
rect 111 348 115 352
rect 1095 348 1099 352
rect 1135 348 1139 352
rect 2119 348 2123 352
rect 111 331 115 335
rect 135 328 139 332
rect 175 328 179 332
rect 215 328 219 332
rect 271 328 275 332
rect 335 328 339 332
rect 399 328 403 332
rect 463 328 467 332
rect 519 328 523 332
rect 575 328 579 332
rect 631 328 635 332
rect 687 328 691 332
rect 751 328 755 332
rect 1095 331 1099 335
rect 1135 331 1139 335
rect 1303 328 1307 332
rect 1343 328 1347 332
rect 1383 328 1387 332
rect 1423 328 1427 332
rect 1463 328 1467 332
rect 1503 328 1507 332
rect 1551 328 1555 332
rect 1615 328 1619 332
rect 1679 328 1683 332
rect 1751 328 1755 332
rect 1831 328 1835 332
rect 1919 328 1923 332
rect 2007 328 2011 332
rect 2071 328 2075 332
rect 2119 331 2123 335
rect 111 309 115 313
rect 135 312 139 316
rect 207 312 211 316
rect 295 312 299 316
rect 383 312 387 316
rect 471 312 475 316
rect 551 312 555 316
rect 623 312 627 316
rect 687 312 691 316
rect 751 312 755 316
rect 807 312 811 316
rect 871 312 875 316
rect 935 312 939 316
rect 1095 309 1099 313
rect 1135 309 1139 313
rect 1167 312 1171 316
rect 1207 312 1211 316
rect 1247 312 1251 316
rect 1295 312 1299 316
rect 1343 312 1347 316
rect 1391 312 1395 316
rect 1439 312 1443 316
rect 1495 312 1499 316
rect 1559 312 1563 316
rect 1623 312 1627 316
rect 1695 312 1699 316
rect 1775 312 1779 316
rect 1855 312 1859 316
rect 1935 312 1939 316
rect 2015 312 2019 316
rect 2071 312 2075 316
rect 2119 309 2123 313
rect 111 292 115 296
rect 1095 292 1099 296
rect 1135 292 1139 296
rect 2119 292 2123 296
rect 135 284 139 288
rect 207 284 211 288
rect 295 284 299 288
rect 383 284 387 288
rect 471 284 475 288
rect 551 284 555 288
rect 623 284 627 288
rect 687 284 691 288
rect 751 284 755 288
rect 807 284 811 288
rect 871 284 875 288
rect 935 284 939 288
rect 1167 284 1171 288
rect 1207 284 1211 288
rect 1247 284 1251 288
rect 1295 284 1299 288
rect 1343 284 1347 288
rect 1391 284 1395 288
rect 1439 284 1443 288
rect 1495 284 1499 288
rect 1559 284 1563 288
rect 1623 284 1627 288
rect 1695 284 1699 288
rect 1775 284 1779 288
rect 1855 284 1859 288
rect 1935 284 1939 288
rect 2015 284 2019 288
rect 2071 284 2075 288
rect 135 248 139 252
rect 199 248 203 252
rect 279 248 283 252
rect 359 248 363 252
rect 439 248 443 252
rect 511 248 515 252
rect 583 248 587 252
rect 647 248 651 252
rect 703 248 707 252
rect 759 248 763 252
rect 815 248 819 252
rect 879 248 883 252
rect 111 240 115 244
rect 1095 240 1099 244
rect 1159 240 1163 244
rect 1207 240 1211 244
rect 1271 240 1275 244
rect 1327 240 1331 244
rect 1391 240 1395 244
rect 1455 240 1459 244
rect 1527 240 1531 244
rect 1607 240 1611 244
rect 1687 240 1691 244
rect 1767 240 1771 244
rect 1839 240 1843 244
rect 1919 240 1923 244
rect 1999 240 2003 244
rect 2071 240 2075 244
rect 1135 232 1139 236
rect 2119 232 2123 236
rect 111 223 115 227
rect 135 220 139 224
rect 199 220 203 224
rect 279 220 283 224
rect 359 220 363 224
rect 439 220 443 224
rect 511 220 515 224
rect 583 220 587 224
rect 647 220 651 224
rect 703 220 707 224
rect 759 220 763 224
rect 815 220 819 224
rect 879 220 883 224
rect 1095 223 1099 227
rect 1135 215 1139 219
rect 1159 212 1163 216
rect 1207 212 1211 216
rect 1271 212 1275 216
rect 1327 212 1331 216
rect 1391 212 1395 216
rect 1455 212 1459 216
rect 1527 212 1531 216
rect 1607 212 1611 216
rect 1687 212 1691 216
rect 1767 212 1771 216
rect 1839 212 1843 216
rect 1919 212 1923 216
rect 1999 212 2003 216
rect 2071 212 2075 216
rect 2119 215 2123 219
rect 111 201 115 205
rect 135 204 139 208
rect 183 204 187 208
rect 231 204 235 208
rect 279 204 283 208
rect 327 204 331 208
rect 375 204 379 208
rect 415 204 419 208
rect 455 204 459 208
rect 503 204 507 208
rect 551 204 555 208
rect 599 204 603 208
rect 647 204 651 208
rect 695 204 699 208
rect 743 204 747 208
rect 1095 201 1099 205
rect 1135 197 1139 201
rect 1159 200 1163 204
rect 1199 200 1203 204
rect 1263 200 1267 204
rect 1327 200 1331 204
rect 1399 200 1403 204
rect 1471 200 1475 204
rect 1543 200 1547 204
rect 1607 200 1611 204
rect 1671 200 1675 204
rect 1735 200 1739 204
rect 1807 200 1811 204
rect 1879 200 1883 204
rect 1951 200 1955 204
rect 2023 200 2027 204
rect 2071 200 2075 204
rect 2119 197 2123 201
rect 111 184 115 188
rect 1095 184 1099 188
rect 135 176 139 180
rect 183 176 187 180
rect 231 176 235 180
rect 279 176 283 180
rect 327 176 331 180
rect 375 176 379 180
rect 415 176 419 180
rect 455 176 459 180
rect 503 176 507 180
rect 551 176 555 180
rect 599 176 603 180
rect 647 176 651 180
rect 695 176 699 180
rect 743 176 747 180
rect 1135 180 1139 184
rect 2119 180 2123 184
rect 1159 172 1163 176
rect 1199 172 1203 176
rect 1263 172 1267 176
rect 1327 172 1331 176
rect 1399 172 1403 176
rect 1471 172 1475 176
rect 1543 172 1547 176
rect 1607 172 1611 176
rect 1671 172 1675 176
rect 1735 172 1739 176
rect 1807 172 1811 176
rect 1879 172 1883 176
rect 1951 172 1955 176
rect 2023 172 2027 176
rect 2071 172 2075 176
rect 143 116 147 120
rect 183 116 187 120
rect 223 116 227 120
rect 263 116 267 120
rect 303 116 307 120
rect 343 116 347 120
rect 383 116 387 120
rect 423 116 427 120
rect 463 116 467 120
rect 503 116 507 120
rect 543 116 547 120
rect 583 116 587 120
rect 623 116 627 120
rect 663 116 667 120
rect 703 116 707 120
rect 743 116 747 120
rect 783 116 787 120
rect 831 116 835 120
rect 879 116 883 120
rect 927 116 931 120
rect 967 116 971 120
rect 1007 116 1011 120
rect 1047 116 1051 120
rect 1159 116 1163 120
rect 1207 116 1211 120
rect 1271 116 1275 120
rect 1335 116 1339 120
rect 1399 116 1403 120
rect 1455 116 1459 120
rect 1511 116 1515 120
rect 1559 116 1563 120
rect 1607 116 1611 120
rect 1647 116 1651 120
rect 1687 116 1691 120
rect 1727 116 1731 120
rect 1767 116 1771 120
rect 1807 116 1811 120
rect 1855 116 1859 120
rect 1903 116 1907 120
rect 1951 116 1955 120
rect 1991 116 1995 120
rect 2031 116 2035 120
rect 2071 116 2075 120
rect 111 108 115 112
rect 1095 108 1099 112
rect 1135 108 1139 112
rect 2119 108 2123 112
rect 111 91 115 95
rect 143 88 147 92
rect 183 88 187 92
rect 223 88 227 92
rect 263 88 267 92
rect 303 88 307 92
rect 343 88 347 92
rect 383 88 387 92
rect 423 88 427 92
rect 463 88 467 92
rect 503 88 507 92
rect 543 88 547 92
rect 583 88 587 92
rect 623 88 627 92
rect 663 88 667 92
rect 703 88 707 92
rect 743 88 747 92
rect 783 88 787 92
rect 831 88 835 92
rect 879 88 883 92
rect 927 88 931 92
rect 967 88 971 92
rect 1007 88 1011 92
rect 1047 88 1051 92
rect 1095 91 1099 95
rect 1135 91 1139 95
rect 1159 88 1163 92
rect 1207 88 1211 92
rect 1271 88 1275 92
rect 1335 88 1339 92
rect 1399 88 1403 92
rect 1455 88 1459 92
rect 1511 88 1515 92
rect 1559 88 1563 92
rect 1607 88 1611 92
rect 1647 88 1651 92
rect 1687 88 1691 92
rect 1727 88 1731 92
rect 1767 88 1771 92
rect 1807 88 1811 92
rect 1855 88 1859 92
rect 1903 88 1907 92
rect 1951 88 1955 92
rect 1991 88 1995 92
rect 2031 88 2035 92
rect 2071 88 2075 92
rect 2119 91 2123 95
<< m3 >>
rect 1135 2230 1139 2231
rect 1135 2225 1139 2226
rect 1687 2230 1691 2231
rect 1687 2225 1691 2226
rect 1727 2230 1731 2231
rect 1727 2225 1731 2226
rect 1767 2230 1771 2231
rect 1767 2225 1771 2226
rect 1807 2230 1811 2231
rect 1807 2225 1811 2226
rect 2119 2230 2123 2231
rect 2119 2225 2123 2226
rect 111 2214 115 2215
rect 111 2209 115 2210
rect 135 2214 139 2215
rect 135 2209 139 2210
rect 175 2214 179 2215
rect 175 2209 179 2210
rect 215 2214 219 2215
rect 215 2209 219 2210
rect 255 2214 259 2215
rect 255 2209 259 2210
rect 319 2214 323 2215
rect 319 2209 323 2210
rect 383 2214 387 2215
rect 383 2209 387 2210
rect 447 2214 451 2215
rect 447 2209 451 2210
rect 511 2214 515 2215
rect 511 2209 515 2210
rect 575 2214 579 2215
rect 575 2209 579 2210
rect 631 2214 635 2215
rect 631 2209 635 2210
rect 687 2214 691 2215
rect 687 2209 691 2210
rect 735 2214 739 2215
rect 735 2209 739 2210
rect 791 2214 795 2215
rect 791 2209 795 2210
rect 847 2214 851 2215
rect 847 2209 851 2210
rect 903 2214 907 2215
rect 903 2209 907 2210
rect 1095 2214 1099 2215
rect 1095 2209 1099 2210
rect 112 2206 114 2209
rect 134 2208 140 2209
rect 110 2205 116 2206
rect 110 2201 111 2205
rect 115 2201 116 2205
rect 134 2204 135 2208
rect 139 2204 140 2208
rect 134 2203 140 2204
rect 174 2208 180 2209
rect 174 2204 175 2208
rect 179 2204 180 2208
rect 174 2203 180 2204
rect 214 2208 220 2209
rect 214 2204 215 2208
rect 219 2204 220 2208
rect 214 2203 220 2204
rect 254 2208 260 2209
rect 254 2204 255 2208
rect 259 2204 260 2208
rect 254 2203 260 2204
rect 318 2208 324 2209
rect 318 2204 319 2208
rect 323 2204 324 2208
rect 318 2203 324 2204
rect 382 2208 388 2209
rect 382 2204 383 2208
rect 387 2204 388 2208
rect 382 2203 388 2204
rect 446 2208 452 2209
rect 446 2204 447 2208
rect 451 2204 452 2208
rect 446 2203 452 2204
rect 510 2208 516 2209
rect 510 2204 511 2208
rect 515 2204 516 2208
rect 510 2203 516 2204
rect 574 2208 580 2209
rect 574 2204 575 2208
rect 579 2204 580 2208
rect 574 2203 580 2204
rect 630 2208 636 2209
rect 630 2204 631 2208
rect 635 2204 636 2208
rect 630 2203 636 2204
rect 686 2208 692 2209
rect 686 2204 687 2208
rect 691 2204 692 2208
rect 686 2203 692 2204
rect 734 2208 740 2209
rect 734 2204 735 2208
rect 739 2204 740 2208
rect 734 2203 740 2204
rect 790 2208 796 2209
rect 790 2204 791 2208
rect 795 2204 796 2208
rect 790 2203 796 2204
rect 846 2208 852 2209
rect 846 2204 847 2208
rect 851 2204 852 2208
rect 846 2203 852 2204
rect 902 2208 908 2209
rect 902 2204 903 2208
rect 907 2204 908 2208
rect 1096 2206 1098 2209
rect 902 2203 908 2204
rect 1094 2205 1100 2206
rect 1136 2205 1138 2225
rect 1688 2213 1690 2225
rect 1728 2213 1730 2225
rect 1768 2213 1770 2225
rect 1808 2213 1810 2225
rect 1686 2212 1692 2213
rect 1686 2208 1687 2212
rect 1691 2208 1692 2212
rect 1686 2207 1692 2208
rect 1726 2212 1732 2213
rect 1726 2208 1727 2212
rect 1731 2208 1732 2212
rect 1726 2207 1732 2208
rect 1766 2212 1772 2213
rect 1766 2208 1767 2212
rect 1771 2208 1772 2212
rect 1766 2207 1772 2208
rect 1806 2212 1812 2213
rect 1806 2208 1807 2212
rect 1811 2208 1812 2212
rect 1806 2207 1812 2208
rect 2120 2205 2122 2225
rect 110 2200 116 2201
rect 1094 2201 1095 2205
rect 1099 2201 1100 2205
rect 1094 2200 1100 2201
rect 1134 2204 1140 2205
rect 1134 2200 1135 2204
rect 1139 2200 1140 2204
rect 1134 2199 1140 2200
rect 2118 2204 2124 2205
rect 2118 2200 2119 2204
rect 2123 2200 2124 2204
rect 2118 2199 2124 2200
rect 110 2188 116 2189
rect 110 2184 111 2188
rect 115 2184 116 2188
rect 110 2183 116 2184
rect 1094 2188 1100 2189
rect 1094 2184 1095 2188
rect 1099 2184 1100 2188
rect 1094 2183 1100 2184
rect 1134 2187 1140 2188
rect 1134 2183 1135 2187
rect 1139 2183 1140 2187
rect 2118 2187 2124 2188
rect 112 2155 114 2183
rect 134 2180 140 2181
rect 134 2176 135 2180
rect 139 2176 140 2180
rect 134 2175 140 2176
rect 174 2180 180 2181
rect 174 2176 175 2180
rect 179 2176 180 2180
rect 174 2175 180 2176
rect 214 2180 220 2181
rect 214 2176 215 2180
rect 219 2176 220 2180
rect 214 2175 220 2176
rect 254 2180 260 2181
rect 254 2176 255 2180
rect 259 2176 260 2180
rect 254 2175 260 2176
rect 318 2180 324 2181
rect 318 2176 319 2180
rect 323 2176 324 2180
rect 318 2175 324 2176
rect 382 2180 388 2181
rect 382 2176 383 2180
rect 387 2176 388 2180
rect 382 2175 388 2176
rect 446 2180 452 2181
rect 446 2176 447 2180
rect 451 2176 452 2180
rect 446 2175 452 2176
rect 510 2180 516 2181
rect 510 2176 511 2180
rect 515 2176 516 2180
rect 510 2175 516 2176
rect 574 2180 580 2181
rect 574 2176 575 2180
rect 579 2176 580 2180
rect 574 2175 580 2176
rect 630 2180 636 2181
rect 630 2176 631 2180
rect 635 2176 636 2180
rect 630 2175 636 2176
rect 686 2180 692 2181
rect 686 2176 687 2180
rect 691 2176 692 2180
rect 686 2175 692 2176
rect 734 2180 740 2181
rect 734 2176 735 2180
rect 739 2176 740 2180
rect 734 2175 740 2176
rect 790 2180 796 2181
rect 790 2176 791 2180
rect 795 2176 796 2180
rect 790 2175 796 2176
rect 846 2180 852 2181
rect 846 2176 847 2180
rect 851 2176 852 2180
rect 846 2175 852 2176
rect 902 2180 908 2181
rect 902 2176 903 2180
rect 907 2176 908 2180
rect 902 2175 908 2176
rect 136 2155 138 2175
rect 176 2155 178 2175
rect 216 2155 218 2175
rect 256 2155 258 2175
rect 320 2155 322 2175
rect 384 2155 386 2175
rect 448 2155 450 2175
rect 512 2155 514 2175
rect 576 2155 578 2175
rect 632 2155 634 2175
rect 688 2155 690 2175
rect 736 2155 738 2175
rect 792 2155 794 2175
rect 848 2155 850 2175
rect 904 2155 906 2175
rect 1096 2155 1098 2183
rect 1134 2182 1140 2183
rect 1686 2184 1692 2185
rect 1136 2179 1138 2182
rect 1686 2180 1687 2184
rect 1691 2180 1692 2184
rect 1686 2179 1692 2180
rect 1726 2184 1732 2185
rect 1726 2180 1727 2184
rect 1731 2180 1732 2184
rect 1726 2179 1732 2180
rect 1766 2184 1772 2185
rect 1766 2180 1767 2184
rect 1771 2180 1772 2184
rect 1766 2179 1772 2180
rect 1806 2184 1812 2185
rect 1806 2180 1807 2184
rect 1811 2180 1812 2184
rect 2118 2183 2119 2187
rect 2123 2183 2124 2187
rect 2118 2182 2124 2183
rect 1806 2179 1812 2180
rect 2120 2179 2122 2182
rect 1135 2178 1139 2179
rect 1135 2173 1139 2174
rect 1159 2178 1163 2179
rect 1159 2173 1163 2174
rect 1199 2178 1203 2179
rect 1199 2173 1203 2174
rect 1239 2178 1243 2179
rect 1239 2173 1243 2174
rect 1279 2178 1283 2179
rect 1279 2173 1283 2174
rect 1335 2178 1339 2179
rect 1335 2173 1339 2174
rect 1391 2178 1395 2179
rect 1391 2173 1395 2174
rect 1455 2178 1459 2179
rect 1455 2173 1459 2174
rect 1527 2178 1531 2179
rect 1527 2173 1531 2174
rect 1591 2178 1595 2179
rect 1591 2173 1595 2174
rect 1663 2178 1667 2179
rect 1663 2173 1667 2174
rect 1687 2178 1691 2179
rect 1687 2173 1691 2174
rect 1727 2178 1731 2179
rect 1727 2173 1731 2174
rect 1735 2178 1739 2179
rect 1735 2173 1739 2174
rect 1767 2178 1771 2179
rect 1767 2173 1771 2174
rect 1807 2178 1811 2179
rect 1807 2173 1811 2174
rect 1879 2178 1883 2179
rect 1879 2173 1883 2174
rect 2119 2178 2123 2179
rect 2119 2173 2123 2174
rect 1136 2170 1138 2173
rect 1158 2172 1164 2173
rect 1134 2169 1140 2170
rect 1134 2165 1135 2169
rect 1139 2165 1140 2169
rect 1158 2168 1159 2172
rect 1163 2168 1164 2172
rect 1158 2167 1164 2168
rect 1198 2172 1204 2173
rect 1198 2168 1199 2172
rect 1203 2168 1204 2172
rect 1198 2167 1204 2168
rect 1238 2172 1244 2173
rect 1238 2168 1239 2172
rect 1243 2168 1244 2172
rect 1238 2167 1244 2168
rect 1278 2172 1284 2173
rect 1278 2168 1279 2172
rect 1283 2168 1284 2172
rect 1278 2167 1284 2168
rect 1334 2172 1340 2173
rect 1334 2168 1335 2172
rect 1339 2168 1340 2172
rect 1334 2167 1340 2168
rect 1390 2172 1396 2173
rect 1390 2168 1391 2172
rect 1395 2168 1396 2172
rect 1390 2167 1396 2168
rect 1454 2172 1460 2173
rect 1454 2168 1455 2172
rect 1459 2168 1460 2172
rect 1454 2167 1460 2168
rect 1526 2172 1532 2173
rect 1526 2168 1527 2172
rect 1531 2168 1532 2172
rect 1526 2167 1532 2168
rect 1590 2172 1596 2173
rect 1590 2168 1591 2172
rect 1595 2168 1596 2172
rect 1590 2167 1596 2168
rect 1662 2172 1668 2173
rect 1662 2168 1663 2172
rect 1667 2168 1668 2172
rect 1662 2167 1668 2168
rect 1734 2172 1740 2173
rect 1734 2168 1735 2172
rect 1739 2168 1740 2172
rect 1734 2167 1740 2168
rect 1806 2172 1812 2173
rect 1806 2168 1807 2172
rect 1811 2168 1812 2172
rect 1806 2167 1812 2168
rect 1878 2172 1884 2173
rect 1878 2168 1879 2172
rect 1883 2168 1884 2172
rect 2120 2170 2122 2173
rect 1878 2167 1884 2168
rect 2118 2169 2124 2170
rect 1134 2164 1140 2165
rect 2118 2165 2119 2169
rect 2123 2165 2124 2169
rect 2118 2164 2124 2165
rect 111 2154 115 2155
rect 111 2149 115 2150
rect 135 2154 139 2155
rect 135 2149 139 2150
rect 175 2154 179 2155
rect 175 2149 179 2150
rect 215 2154 219 2155
rect 215 2149 219 2150
rect 231 2154 235 2155
rect 231 2149 235 2150
rect 255 2154 259 2155
rect 255 2149 259 2150
rect 271 2154 275 2155
rect 271 2149 275 2150
rect 311 2154 315 2155
rect 311 2149 315 2150
rect 319 2154 323 2155
rect 319 2149 323 2150
rect 359 2154 363 2155
rect 359 2149 363 2150
rect 383 2154 387 2155
rect 383 2149 387 2150
rect 423 2154 427 2155
rect 423 2149 427 2150
rect 447 2154 451 2155
rect 447 2149 451 2150
rect 487 2154 491 2155
rect 487 2149 491 2150
rect 511 2154 515 2155
rect 511 2149 515 2150
rect 559 2154 563 2155
rect 559 2149 563 2150
rect 575 2154 579 2155
rect 575 2149 579 2150
rect 631 2154 635 2155
rect 631 2149 635 2150
rect 639 2154 643 2155
rect 639 2149 643 2150
rect 687 2154 691 2155
rect 687 2149 691 2150
rect 719 2154 723 2155
rect 719 2149 723 2150
rect 735 2154 739 2155
rect 735 2149 739 2150
rect 791 2154 795 2155
rect 791 2149 795 2150
rect 799 2154 803 2155
rect 799 2149 803 2150
rect 847 2154 851 2155
rect 847 2149 851 2150
rect 879 2154 883 2155
rect 879 2149 883 2150
rect 903 2154 907 2155
rect 903 2149 907 2150
rect 967 2154 971 2155
rect 967 2149 971 2150
rect 1095 2154 1099 2155
rect 1095 2149 1099 2150
rect 1134 2152 1140 2153
rect 112 2129 114 2149
rect 232 2137 234 2149
rect 272 2137 274 2149
rect 312 2137 314 2149
rect 360 2137 362 2149
rect 424 2137 426 2149
rect 488 2137 490 2149
rect 560 2137 562 2149
rect 640 2137 642 2149
rect 720 2137 722 2149
rect 800 2137 802 2149
rect 880 2137 882 2149
rect 968 2137 970 2149
rect 230 2136 236 2137
rect 230 2132 231 2136
rect 235 2132 236 2136
rect 230 2131 236 2132
rect 270 2136 276 2137
rect 270 2132 271 2136
rect 275 2132 276 2136
rect 270 2131 276 2132
rect 310 2136 316 2137
rect 310 2132 311 2136
rect 315 2132 316 2136
rect 310 2131 316 2132
rect 358 2136 364 2137
rect 358 2132 359 2136
rect 363 2132 364 2136
rect 358 2131 364 2132
rect 422 2136 428 2137
rect 422 2132 423 2136
rect 427 2132 428 2136
rect 422 2131 428 2132
rect 486 2136 492 2137
rect 486 2132 487 2136
rect 491 2132 492 2136
rect 486 2131 492 2132
rect 558 2136 564 2137
rect 558 2132 559 2136
rect 563 2132 564 2136
rect 558 2131 564 2132
rect 638 2136 644 2137
rect 638 2132 639 2136
rect 643 2132 644 2136
rect 638 2131 644 2132
rect 718 2136 724 2137
rect 718 2132 719 2136
rect 723 2132 724 2136
rect 718 2131 724 2132
rect 798 2136 804 2137
rect 798 2132 799 2136
rect 803 2132 804 2136
rect 798 2131 804 2132
rect 878 2136 884 2137
rect 878 2132 879 2136
rect 883 2132 884 2136
rect 878 2131 884 2132
rect 966 2136 972 2137
rect 966 2132 967 2136
rect 971 2132 972 2136
rect 966 2131 972 2132
rect 1096 2129 1098 2149
rect 1134 2148 1135 2152
rect 1139 2148 1140 2152
rect 1134 2147 1140 2148
rect 2118 2152 2124 2153
rect 2118 2148 2119 2152
rect 2123 2148 2124 2152
rect 2118 2147 2124 2148
rect 110 2128 116 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 1094 2128 1100 2129
rect 1094 2124 1095 2128
rect 1099 2124 1100 2128
rect 1136 2127 1138 2147
rect 1158 2144 1164 2145
rect 1158 2140 1159 2144
rect 1163 2140 1164 2144
rect 1158 2139 1164 2140
rect 1198 2144 1204 2145
rect 1198 2140 1199 2144
rect 1203 2140 1204 2144
rect 1198 2139 1204 2140
rect 1238 2144 1244 2145
rect 1238 2140 1239 2144
rect 1243 2140 1244 2144
rect 1238 2139 1244 2140
rect 1278 2144 1284 2145
rect 1278 2140 1279 2144
rect 1283 2140 1284 2144
rect 1278 2139 1284 2140
rect 1334 2144 1340 2145
rect 1334 2140 1335 2144
rect 1339 2140 1340 2144
rect 1334 2139 1340 2140
rect 1390 2144 1396 2145
rect 1390 2140 1391 2144
rect 1395 2140 1396 2144
rect 1390 2139 1396 2140
rect 1454 2144 1460 2145
rect 1454 2140 1455 2144
rect 1459 2140 1460 2144
rect 1454 2139 1460 2140
rect 1526 2144 1532 2145
rect 1526 2140 1527 2144
rect 1531 2140 1532 2144
rect 1526 2139 1532 2140
rect 1590 2144 1596 2145
rect 1590 2140 1591 2144
rect 1595 2140 1596 2144
rect 1590 2139 1596 2140
rect 1662 2144 1668 2145
rect 1662 2140 1663 2144
rect 1667 2140 1668 2144
rect 1662 2139 1668 2140
rect 1734 2144 1740 2145
rect 1734 2140 1735 2144
rect 1739 2140 1740 2144
rect 1734 2139 1740 2140
rect 1806 2144 1812 2145
rect 1806 2140 1807 2144
rect 1811 2140 1812 2144
rect 1806 2139 1812 2140
rect 1878 2144 1884 2145
rect 1878 2140 1879 2144
rect 1883 2140 1884 2144
rect 1878 2139 1884 2140
rect 1160 2127 1162 2139
rect 1200 2127 1202 2139
rect 1240 2127 1242 2139
rect 1280 2127 1282 2139
rect 1336 2127 1338 2139
rect 1392 2127 1394 2139
rect 1456 2127 1458 2139
rect 1528 2127 1530 2139
rect 1592 2127 1594 2139
rect 1664 2127 1666 2139
rect 1736 2127 1738 2139
rect 1808 2127 1810 2139
rect 1880 2127 1882 2139
rect 2120 2127 2122 2147
rect 1094 2123 1100 2124
rect 1135 2126 1139 2127
rect 1135 2121 1139 2122
rect 1159 2126 1163 2127
rect 1159 2121 1163 2122
rect 1199 2126 1203 2127
rect 1199 2121 1203 2122
rect 1239 2126 1243 2127
rect 1239 2121 1243 2122
rect 1279 2126 1283 2127
rect 1279 2121 1283 2122
rect 1295 2126 1299 2127
rect 1295 2121 1299 2122
rect 1335 2126 1339 2127
rect 1335 2121 1339 2122
rect 1367 2126 1371 2127
rect 1367 2121 1371 2122
rect 1391 2126 1395 2127
rect 1391 2121 1395 2122
rect 1439 2126 1443 2127
rect 1439 2121 1443 2122
rect 1455 2126 1459 2127
rect 1455 2121 1459 2122
rect 1519 2126 1523 2127
rect 1519 2121 1523 2122
rect 1527 2126 1531 2127
rect 1527 2121 1531 2122
rect 1591 2126 1595 2127
rect 1591 2121 1595 2122
rect 1599 2126 1603 2127
rect 1599 2121 1603 2122
rect 1663 2126 1667 2127
rect 1663 2121 1667 2122
rect 1679 2126 1683 2127
rect 1679 2121 1683 2122
rect 1735 2126 1739 2127
rect 1735 2121 1739 2122
rect 1751 2126 1755 2127
rect 1751 2121 1755 2122
rect 1807 2126 1811 2127
rect 1807 2121 1811 2122
rect 1823 2126 1827 2127
rect 1823 2121 1827 2122
rect 1879 2126 1883 2127
rect 1879 2121 1883 2122
rect 1887 2126 1891 2127
rect 1887 2121 1891 2122
rect 1951 2126 1955 2127
rect 1951 2121 1955 2122
rect 2023 2126 2027 2127
rect 2023 2121 2027 2122
rect 2071 2126 2075 2127
rect 2071 2121 2075 2122
rect 2119 2126 2123 2127
rect 2119 2121 2123 2122
rect 110 2111 116 2112
rect 110 2107 111 2111
rect 115 2107 116 2111
rect 1094 2111 1100 2112
rect 110 2106 116 2107
rect 230 2108 236 2109
rect 112 2099 114 2106
rect 230 2104 231 2108
rect 235 2104 236 2108
rect 230 2103 236 2104
rect 270 2108 276 2109
rect 270 2104 271 2108
rect 275 2104 276 2108
rect 270 2103 276 2104
rect 310 2108 316 2109
rect 310 2104 311 2108
rect 315 2104 316 2108
rect 310 2103 316 2104
rect 358 2108 364 2109
rect 358 2104 359 2108
rect 363 2104 364 2108
rect 358 2103 364 2104
rect 422 2108 428 2109
rect 422 2104 423 2108
rect 427 2104 428 2108
rect 422 2103 428 2104
rect 486 2108 492 2109
rect 486 2104 487 2108
rect 491 2104 492 2108
rect 486 2103 492 2104
rect 558 2108 564 2109
rect 558 2104 559 2108
rect 563 2104 564 2108
rect 558 2103 564 2104
rect 638 2108 644 2109
rect 638 2104 639 2108
rect 643 2104 644 2108
rect 638 2103 644 2104
rect 718 2108 724 2109
rect 718 2104 719 2108
rect 723 2104 724 2108
rect 718 2103 724 2104
rect 798 2108 804 2109
rect 798 2104 799 2108
rect 803 2104 804 2108
rect 798 2103 804 2104
rect 878 2108 884 2109
rect 878 2104 879 2108
rect 883 2104 884 2108
rect 878 2103 884 2104
rect 966 2108 972 2109
rect 966 2104 967 2108
rect 971 2104 972 2108
rect 1094 2107 1095 2111
rect 1099 2107 1100 2111
rect 1094 2106 1100 2107
rect 966 2103 972 2104
rect 232 2099 234 2103
rect 272 2099 274 2103
rect 312 2099 314 2103
rect 360 2099 362 2103
rect 424 2099 426 2103
rect 488 2099 490 2103
rect 560 2099 562 2103
rect 640 2099 642 2103
rect 720 2099 722 2103
rect 800 2099 802 2103
rect 880 2099 882 2103
rect 968 2099 970 2103
rect 1096 2099 1098 2106
rect 1136 2101 1138 2121
rect 1160 2109 1162 2121
rect 1200 2109 1202 2121
rect 1240 2109 1242 2121
rect 1296 2109 1298 2121
rect 1368 2109 1370 2121
rect 1440 2109 1442 2121
rect 1520 2109 1522 2121
rect 1600 2109 1602 2121
rect 1680 2109 1682 2121
rect 1752 2109 1754 2121
rect 1824 2109 1826 2121
rect 1888 2109 1890 2121
rect 1952 2109 1954 2121
rect 2024 2109 2026 2121
rect 2072 2109 2074 2121
rect 1158 2108 1164 2109
rect 1158 2104 1159 2108
rect 1163 2104 1164 2108
rect 1158 2103 1164 2104
rect 1198 2108 1204 2109
rect 1198 2104 1199 2108
rect 1203 2104 1204 2108
rect 1198 2103 1204 2104
rect 1238 2108 1244 2109
rect 1238 2104 1239 2108
rect 1243 2104 1244 2108
rect 1238 2103 1244 2104
rect 1294 2108 1300 2109
rect 1294 2104 1295 2108
rect 1299 2104 1300 2108
rect 1294 2103 1300 2104
rect 1366 2108 1372 2109
rect 1366 2104 1367 2108
rect 1371 2104 1372 2108
rect 1366 2103 1372 2104
rect 1438 2108 1444 2109
rect 1438 2104 1439 2108
rect 1443 2104 1444 2108
rect 1438 2103 1444 2104
rect 1518 2108 1524 2109
rect 1518 2104 1519 2108
rect 1523 2104 1524 2108
rect 1518 2103 1524 2104
rect 1598 2108 1604 2109
rect 1598 2104 1599 2108
rect 1603 2104 1604 2108
rect 1598 2103 1604 2104
rect 1678 2108 1684 2109
rect 1678 2104 1679 2108
rect 1683 2104 1684 2108
rect 1678 2103 1684 2104
rect 1750 2108 1756 2109
rect 1750 2104 1751 2108
rect 1755 2104 1756 2108
rect 1750 2103 1756 2104
rect 1822 2108 1828 2109
rect 1822 2104 1823 2108
rect 1827 2104 1828 2108
rect 1822 2103 1828 2104
rect 1886 2108 1892 2109
rect 1886 2104 1887 2108
rect 1891 2104 1892 2108
rect 1886 2103 1892 2104
rect 1950 2108 1956 2109
rect 1950 2104 1951 2108
rect 1955 2104 1956 2108
rect 1950 2103 1956 2104
rect 2022 2108 2028 2109
rect 2022 2104 2023 2108
rect 2027 2104 2028 2108
rect 2022 2103 2028 2104
rect 2070 2108 2076 2109
rect 2070 2104 2071 2108
rect 2075 2104 2076 2108
rect 2070 2103 2076 2104
rect 2120 2101 2122 2121
rect 1134 2100 1140 2101
rect 111 2098 115 2099
rect 111 2093 115 2094
rect 231 2098 235 2099
rect 231 2093 235 2094
rect 271 2098 275 2099
rect 271 2093 275 2094
rect 303 2098 307 2099
rect 303 2093 307 2094
rect 311 2098 315 2099
rect 311 2093 315 2094
rect 351 2098 355 2099
rect 351 2093 355 2094
rect 359 2098 363 2099
rect 359 2093 363 2094
rect 407 2098 411 2099
rect 407 2093 411 2094
rect 423 2098 427 2099
rect 423 2093 427 2094
rect 471 2098 475 2099
rect 471 2093 475 2094
rect 487 2098 491 2099
rect 487 2093 491 2094
rect 543 2098 547 2099
rect 543 2093 547 2094
rect 559 2098 563 2099
rect 559 2093 563 2094
rect 623 2098 627 2099
rect 623 2093 627 2094
rect 639 2098 643 2099
rect 639 2093 643 2094
rect 703 2098 707 2099
rect 703 2093 707 2094
rect 719 2098 723 2099
rect 719 2093 723 2094
rect 783 2098 787 2099
rect 783 2093 787 2094
rect 799 2098 803 2099
rect 799 2093 803 2094
rect 863 2098 867 2099
rect 863 2093 867 2094
rect 879 2098 883 2099
rect 879 2093 883 2094
rect 951 2098 955 2099
rect 951 2093 955 2094
rect 967 2098 971 2099
rect 967 2093 971 2094
rect 1039 2098 1043 2099
rect 1039 2093 1043 2094
rect 1095 2098 1099 2099
rect 1134 2096 1135 2100
rect 1139 2096 1140 2100
rect 1134 2095 1140 2096
rect 2118 2100 2124 2101
rect 2118 2096 2119 2100
rect 2123 2096 2124 2100
rect 2118 2095 2124 2096
rect 1095 2093 1099 2094
rect 112 2090 114 2093
rect 302 2092 308 2093
rect 110 2089 116 2090
rect 110 2085 111 2089
rect 115 2085 116 2089
rect 302 2088 303 2092
rect 307 2088 308 2092
rect 302 2087 308 2088
rect 350 2092 356 2093
rect 350 2088 351 2092
rect 355 2088 356 2092
rect 350 2087 356 2088
rect 406 2092 412 2093
rect 406 2088 407 2092
rect 411 2088 412 2092
rect 406 2087 412 2088
rect 470 2092 476 2093
rect 470 2088 471 2092
rect 475 2088 476 2092
rect 470 2087 476 2088
rect 542 2092 548 2093
rect 542 2088 543 2092
rect 547 2088 548 2092
rect 542 2087 548 2088
rect 622 2092 628 2093
rect 622 2088 623 2092
rect 627 2088 628 2092
rect 622 2087 628 2088
rect 702 2092 708 2093
rect 702 2088 703 2092
rect 707 2088 708 2092
rect 702 2087 708 2088
rect 782 2092 788 2093
rect 782 2088 783 2092
rect 787 2088 788 2092
rect 782 2087 788 2088
rect 862 2092 868 2093
rect 862 2088 863 2092
rect 867 2088 868 2092
rect 862 2087 868 2088
rect 950 2092 956 2093
rect 950 2088 951 2092
rect 955 2088 956 2092
rect 950 2087 956 2088
rect 1038 2092 1044 2093
rect 1038 2088 1039 2092
rect 1043 2088 1044 2092
rect 1096 2090 1098 2093
rect 1038 2087 1044 2088
rect 1094 2089 1100 2090
rect 110 2084 116 2085
rect 1094 2085 1095 2089
rect 1099 2085 1100 2089
rect 1094 2084 1100 2085
rect 1134 2083 1140 2084
rect 1134 2079 1135 2083
rect 1139 2079 1140 2083
rect 2118 2083 2124 2084
rect 1134 2078 1140 2079
rect 1158 2080 1164 2081
rect 1136 2075 1138 2078
rect 1158 2076 1159 2080
rect 1163 2076 1164 2080
rect 1158 2075 1164 2076
rect 1198 2080 1204 2081
rect 1198 2076 1199 2080
rect 1203 2076 1204 2080
rect 1198 2075 1204 2076
rect 1238 2080 1244 2081
rect 1238 2076 1239 2080
rect 1243 2076 1244 2080
rect 1238 2075 1244 2076
rect 1294 2080 1300 2081
rect 1294 2076 1295 2080
rect 1299 2076 1300 2080
rect 1294 2075 1300 2076
rect 1366 2080 1372 2081
rect 1366 2076 1367 2080
rect 1371 2076 1372 2080
rect 1366 2075 1372 2076
rect 1438 2080 1444 2081
rect 1438 2076 1439 2080
rect 1443 2076 1444 2080
rect 1438 2075 1444 2076
rect 1518 2080 1524 2081
rect 1518 2076 1519 2080
rect 1523 2076 1524 2080
rect 1518 2075 1524 2076
rect 1598 2080 1604 2081
rect 1598 2076 1599 2080
rect 1603 2076 1604 2080
rect 1598 2075 1604 2076
rect 1678 2080 1684 2081
rect 1678 2076 1679 2080
rect 1683 2076 1684 2080
rect 1678 2075 1684 2076
rect 1750 2080 1756 2081
rect 1750 2076 1751 2080
rect 1755 2076 1756 2080
rect 1750 2075 1756 2076
rect 1822 2080 1828 2081
rect 1822 2076 1823 2080
rect 1827 2076 1828 2080
rect 1822 2075 1828 2076
rect 1886 2080 1892 2081
rect 1886 2076 1887 2080
rect 1891 2076 1892 2080
rect 1886 2075 1892 2076
rect 1950 2080 1956 2081
rect 1950 2076 1951 2080
rect 1955 2076 1956 2080
rect 1950 2075 1956 2076
rect 2022 2080 2028 2081
rect 2022 2076 2023 2080
rect 2027 2076 2028 2080
rect 2022 2075 2028 2076
rect 2070 2080 2076 2081
rect 2070 2076 2071 2080
rect 2075 2076 2076 2080
rect 2118 2079 2119 2083
rect 2123 2079 2124 2083
rect 2118 2078 2124 2079
rect 2070 2075 2076 2076
rect 2120 2075 2122 2078
rect 1135 2074 1139 2075
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 1094 2072 1100 2073
rect 1094 2068 1095 2072
rect 1099 2068 1100 2072
rect 1135 2069 1139 2070
rect 1159 2074 1163 2075
rect 1159 2069 1163 2070
rect 1199 2074 1203 2075
rect 1199 2069 1203 2070
rect 1215 2074 1219 2075
rect 1215 2069 1219 2070
rect 1239 2074 1243 2075
rect 1239 2069 1243 2070
rect 1295 2074 1299 2075
rect 1295 2069 1299 2070
rect 1303 2074 1307 2075
rect 1303 2069 1307 2070
rect 1367 2074 1371 2075
rect 1367 2069 1371 2070
rect 1399 2074 1403 2075
rect 1399 2069 1403 2070
rect 1439 2074 1443 2075
rect 1439 2069 1443 2070
rect 1495 2074 1499 2075
rect 1495 2069 1499 2070
rect 1519 2074 1523 2075
rect 1519 2069 1523 2070
rect 1591 2074 1595 2075
rect 1591 2069 1595 2070
rect 1599 2074 1603 2075
rect 1599 2069 1603 2070
rect 1679 2074 1683 2075
rect 1679 2069 1683 2070
rect 1751 2074 1755 2075
rect 1751 2069 1755 2070
rect 1759 2074 1763 2075
rect 1759 2069 1763 2070
rect 1823 2074 1827 2075
rect 1823 2069 1827 2070
rect 1831 2074 1835 2075
rect 1831 2069 1835 2070
rect 1887 2074 1891 2075
rect 1887 2069 1891 2070
rect 1895 2074 1899 2075
rect 1895 2069 1899 2070
rect 1951 2074 1955 2075
rect 1951 2069 1955 2070
rect 1959 2074 1963 2075
rect 1959 2069 1963 2070
rect 2023 2074 2027 2075
rect 2023 2069 2027 2070
rect 2071 2074 2075 2075
rect 2071 2069 2075 2070
rect 2119 2074 2123 2075
rect 2119 2069 2123 2070
rect 1094 2067 1100 2068
rect 112 2043 114 2067
rect 302 2064 308 2065
rect 302 2060 303 2064
rect 307 2060 308 2064
rect 302 2059 308 2060
rect 350 2064 356 2065
rect 350 2060 351 2064
rect 355 2060 356 2064
rect 350 2059 356 2060
rect 406 2064 412 2065
rect 406 2060 407 2064
rect 411 2060 412 2064
rect 406 2059 412 2060
rect 470 2064 476 2065
rect 470 2060 471 2064
rect 475 2060 476 2064
rect 470 2059 476 2060
rect 542 2064 548 2065
rect 542 2060 543 2064
rect 547 2060 548 2064
rect 542 2059 548 2060
rect 622 2064 628 2065
rect 622 2060 623 2064
rect 627 2060 628 2064
rect 622 2059 628 2060
rect 702 2064 708 2065
rect 702 2060 703 2064
rect 707 2060 708 2064
rect 702 2059 708 2060
rect 782 2064 788 2065
rect 782 2060 783 2064
rect 787 2060 788 2064
rect 782 2059 788 2060
rect 862 2064 868 2065
rect 862 2060 863 2064
rect 867 2060 868 2064
rect 862 2059 868 2060
rect 950 2064 956 2065
rect 950 2060 951 2064
rect 955 2060 956 2064
rect 950 2059 956 2060
rect 1038 2064 1044 2065
rect 1038 2060 1039 2064
rect 1043 2060 1044 2064
rect 1038 2059 1044 2060
rect 304 2043 306 2059
rect 352 2043 354 2059
rect 408 2043 410 2059
rect 472 2043 474 2059
rect 544 2043 546 2059
rect 624 2043 626 2059
rect 704 2043 706 2059
rect 784 2043 786 2059
rect 864 2043 866 2059
rect 952 2043 954 2059
rect 1040 2043 1042 2059
rect 1096 2043 1098 2067
rect 1136 2066 1138 2069
rect 1158 2068 1164 2069
rect 1134 2065 1140 2066
rect 1134 2061 1135 2065
rect 1139 2061 1140 2065
rect 1158 2064 1159 2068
rect 1163 2064 1164 2068
rect 1158 2063 1164 2064
rect 1214 2068 1220 2069
rect 1214 2064 1215 2068
rect 1219 2064 1220 2068
rect 1214 2063 1220 2064
rect 1302 2068 1308 2069
rect 1302 2064 1303 2068
rect 1307 2064 1308 2068
rect 1302 2063 1308 2064
rect 1398 2068 1404 2069
rect 1398 2064 1399 2068
rect 1403 2064 1404 2068
rect 1398 2063 1404 2064
rect 1494 2068 1500 2069
rect 1494 2064 1495 2068
rect 1499 2064 1500 2068
rect 1494 2063 1500 2064
rect 1590 2068 1596 2069
rect 1590 2064 1591 2068
rect 1595 2064 1596 2068
rect 1590 2063 1596 2064
rect 1678 2068 1684 2069
rect 1678 2064 1679 2068
rect 1683 2064 1684 2068
rect 1678 2063 1684 2064
rect 1758 2068 1764 2069
rect 1758 2064 1759 2068
rect 1763 2064 1764 2068
rect 1758 2063 1764 2064
rect 1830 2068 1836 2069
rect 1830 2064 1831 2068
rect 1835 2064 1836 2068
rect 1830 2063 1836 2064
rect 1894 2068 1900 2069
rect 1894 2064 1895 2068
rect 1899 2064 1900 2068
rect 1894 2063 1900 2064
rect 1958 2068 1964 2069
rect 1958 2064 1959 2068
rect 1963 2064 1964 2068
rect 1958 2063 1964 2064
rect 2022 2068 2028 2069
rect 2022 2064 2023 2068
rect 2027 2064 2028 2068
rect 2022 2063 2028 2064
rect 2070 2068 2076 2069
rect 2070 2064 2071 2068
rect 2075 2064 2076 2068
rect 2120 2066 2122 2069
rect 2070 2063 2076 2064
rect 2118 2065 2124 2066
rect 1134 2060 1140 2061
rect 2118 2061 2119 2065
rect 2123 2061 2124 2065
rect 2118 2060 2124 2061
rect 1134 2048 1140 2049
rect 1134 2044 1135 2048
rect 1139 2044 1140 2048
rect 1134 2043 1140 2044
rect 2118 2048 2124 2049
rect 2118 2044 2119 2048
rect 2123 2044 2124 2048
rect 2118 2043 2124 2044
rect 111 2042 115 2043
rect 111 2037 115 2038
rect 183 2042 187 2043
rect 183 2037 187 2038
rect 279 2042 283 2043
rect 279 2037 283 2038
rect 303 2042 307 2043
rect 303 2037 307 2038
rect 351 2042 355 2043
rect 351 2037 355 2038
rect 375 2042 379 2043
rect 375 2037 379 2038
rect 407 2042 411 2043
rect 407 2037 411 2038
rect 463 2042 467 2043
rect 463 2037 467 2038
rect 471 2042 475 2043
rect 471 2037 475 2038
rect 543 2042 547 2043
rect 543 2037 547 2038
rect 623 2042 627 2043
rect 623 2037 627 2038
rect 695 2042 699 2043
rect 695 2037 699 2038
rect 703 2042 707 2043
rect 703 2037 707 2038
rect 759 2042 763 2043
rect 759 2037 763 2038
rect 783 2042 787 2043
rect 783 2037 787 2038
rect 815 2042 819 2043
rect 815 2037 819 2038
rect 863 2042 867 2043
rect 863 2037 867 2038
rect 911 2042 915 2043
rect 911 2037 915 2038
rect 951 2042 955 2043
rect 951 2037 955 2038
rect 959 2042 963 2043
rect 959 2037 963 2038
rect 1007 2042 1011 2043
rect 1007 2037 1011 2038
rect 1039 2042 1043 2043
rect 1039 2037 1043 2038
rect 1047 2042 1051 2043
rect 1047 2037 1051 2038
rect 1095 2042 1099 2043
rect 1095 2037 1099 2038
rect 112 2017 114 2037
rect 184 2025 186 2037
rect 280 2025 282 2037
rect 376 2025 378 2037
rect 464 2025 466 2037
rect 544 2025 546 2037
rect 624 2025 626 2037
rect 696 2025 698 2037
rect 760 2025 762 2037
rect 816 2025 818 2037
rect 864 2025 866 2037
rect 912 2025 914 2037
rect 960 2025 962 2037
rect 1008 2025 1010 2037
rect 1048 2025 1050 2037
rect 182 2024 188 2025
rect 182 2020 183 2024
rect 187 2020 188 2024
rect 182 2019 188 2020
rect 278 2024 284 2025
rect 278 2020 279 2024
rect 283 2020 284 2024
rect 278 2019 284 2020
rect 374 2024 380 2025
rect 374 2020 375 2024
rect 379 2020 380 2024
rect 374 2019 380 2020
rect 462 2024 468 2025
rect 462 2020 463 2024
rect 467 2020 468 2024
rect 462 2019 468 2020
rect 542 2024 548 2025
rect 542 2020 543 2024
rect 547 2020 548 2024
rect 542 2019 548 2020
rect 622 2024 628 2025
rect 622 2020 623 2024
rect 627 2020 628 2024
rect 622 2019 628 2020
rect 694 2024 700 2025
rect 694 2020 695 2024
rect 699 2020 700 2024
rect 694 2019 700 2020
rect 758 2024 764 2025
rect 758 2020 759 2024
rect 763 2020 764 2024
rect 758 2019 764 2020
rect 814 2024 820 2025
rect 814 2020 815 2024
rect 819 2020 820 2024
rect 814 2019 820 2020
rect 862 2024 868 2025
rect 862 2020 863 2024
rect 867 2020 868 2024
rect 862 2019 868 2020
rect 910 2024 916 2025
rect 910 2020 911 2024
rect 915 2020 916 2024
rect 910 2019 916 2020
rect 958 2024 964 2025
rect 958 2020 959 2024
rect 963 2020 964 2024
rect 958 2019 964 2020
rect 1006 2024 1012 2025
rect 1006 2020 1007 2024
rect 1011 2020 1012 2024
rect 1006 2019 1012 2020
rect 1046 2024 1052 2025
rect 1046 2020 1047 2024
rect 1051 2020 1052 2024
rect 1046 2019 1052 2020
rect 1096 2017 1098 2037
rect 1136 2023 1138 2043
rect 1158 2040 1164 2041
rect 1158 2036 1159 2040
rect 1163 2036 1164 2040
rect 1158 2035 1164 2036
rect 1214 2040 1220 2041
rect 1214 2036 1215 2040
rect 1219 2036 1220 2040
rect 1214 2035 1220 2036
rect 1302 2040 1308 2041
rect 1302 2036 1303 2040
rect 1307 2036 1308 2040
rect 1302 2035 1308 2036
rect 1398 2040 1404 2041
rect 1398 2036 1399 2040
rect 1403 2036 1404 2040
rect 1398 2035 1404 2036
rect 1494 2040 1500 2041
rect 1494 2036 1495 2040
rect 1499 2036 1500 2040
rect 1494 2035 1500 2036
rect 1590 2040 1596 2041
rect 1590 2036 1591 2040
rect 1595 2036 1596 2040
rect 1590 2035 1596 2036
rect 1678 2040 1684 2041
rect 1678 2036 1679 2040
rect 1683 2036 1684 2040
rect 1678 2035 1684 2036
rect 1758 2040 1764 2041
rect 1758 2036 1759 2040
rect 1763 2036 1764 2040
rect 1758 2035 1764 2036
rect 1830 2040 1836 2041
rect 1830 2036 1831 2040
rect 1835 2036 1836 2040
rect 1830 2035 1836 2036
rect 1894 2040 1900 2041
rect 1894 2036 1895 2040
rect 1899 2036 1900 2040
rect 1894 2035 1900 2036
rect 1958 2040 1964 2041
rect 1958 2036 1959 2040
rect 1963 2036 1964 2040
rect 1958 2035 1964 2036
rect 2022 2040 2028 2041
rect 2022 2036 2023 2040
rect 2027 2036 2028 2040
rect 2022 2035 2028 2036
rect 2070 2040 2076 2041
rect 2070 2036 2071 2040
rect 2075 2036 2076 2040
rect 2070 2035 2076 2036
rect 1160 2023 1162 2035
rect 1216 2023 1218 2035
rect 1304 2023 1306 2035
rect 1400 2023 1402 2035
rect 1496 2023 1498 2035
rect 1592 2023 1594 2035
rect 1680 2023 1682 2035
rect 1760 2023 1762 2035
rect 1832 2023 1834 2035
rect 1896 2023 1898 2035
rect 1960 2023 1962 2035
rect 2024 2023 2026 2035
rect 2072 2023 2074 2035
rect 2120 2023 2122 2043
rect 1135 2022 1139 2023
rect 1135 2017 1139 2018
rect 1159 2022 1163 2023
rect 1159 2017 1163 2018
rect 1215 2022 1219 2023
rect 1215 2017 1219 2018
rect 1239 2022 1243 2023
rect 1239 2017 1243 2018
rect 1303 2022 1307 2023
rect 1303 2017 1307 2018
rect 1351 2022 1355 2023
rect 1351 2017 1355 2018
rect 1399 2022 1403 2023
rect 1399 2017 1403 2018
rect 1455 2022 1459 2023
rect 1455 2017 1459 2018
rect 1495 2022 1499 2023
rect 1495 2017 1499 2018
rect 1559 2022 1563 2023
rect 1559 2017 1563 2018
rect 1591 2022 1595 2023
rect 1591 2017 1595 2018
rect 1655 2022 1659 2023
rect 1655 2017 1659 2018
rect 1679 2022 1683 2023
rect 1679 2017 1683 2018
rect 1743 2022 1747 2023
rect 1743 2017 1747 2018
rect 1759 2022 1763 2023
rect 1759 2017 1763 2018
rect 1823 2022 1827 2023
rect 1823 2017 1827 2018
rect 1831 2022 1835 2023
rect 1831 2017 1835 2018
rect 1895 2022 1899 2023
rect 1895 2017 1899 2018
rect 1959 2022 1963 2023
rect 1959 2017 1963 2018
rect 2023 2022 2027 2023
rect 2023 2017 2027 2018
rect 2071 2022 2075 2023
rect 2071 2017 2075 2018
rect 2119 2022 2123 2023
rect 2119 2017 2123 2018
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 110 2011 116 2012
rect 1094 2016 1100 2017
rect 1094 2012 1095 2016
rect 1099 2012 1100 2016
rect 1094 2011 1100 2012
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 1094 1999 1100 2000
rect 110 1994 116 1995
rect 182 1996 188 1997
rect 112 1991 114 1994
rect 182 1992 183 1996
rect 187 1992 188 1996
rect 182 1991 188 1992
rect 278 1996 284 1997
rect 278 1992 279 1996
rect 283 1992 284 1996
rect 278 1991 284 1992
rect 374 1996 380 1997
rect 374 1992 375 1996
rect 379 1992 380 1996
rect 374 1991 380 1992
rect 462 1996 468 1997
rect 462 1992 463 1996
rect 467 1992 468 1996
rect 462 1991 468 1992
rect 542 1996 548 1997
rect 542 1992 543 1996
rect 547 1992 548 1996
rect 542 1991 548 1992
rect 622 1996 628 1997
rect 622 1992 623 1996
rect 627 1992 628 1996
rect 622 1991 628 1992
rect 694 1996 700 1997
rect 694 1992 695 1996
rect 699 1992 700 1996
rect 694 1991 700 1992
rect 758 1996 764 1997
rect 758 1992 759 1996
rect 763 1992 764 1996
rect 758 1991 764 1992
rect 814 1996 820 1997
rect 814 1992 815 1996
rect 819 1992 820 1996
rect 814 1991 820 1992
rect 862 1996 868 1997
rect 862 1992 863 1996
rect 867 1992 868 1996
rect 862 1991 868 1992
rect 910 1996 916 1997
rect 910 1992 911 1996
rect 915 1992 916 1996
rect 910 1991 916 1992
rect 958 1996 964 1997
rect 958 1992 959 1996
rect 963 1992 964 1996
rect 958 1991 964 1992
rect 1006 1996 1012 1997
rect 1006 1992 1007 1996
rect 1011 1992 1012 1996
rect 1006 1991 1012 1992
rect 1046 1996 1052 1997
rect 1046 1992 1047 1996
rect 1051 1992 1052 1996
rect 1094 1995 1095 1999
rect 1099 1995 1100 1999
rect 1136 1997 1138 2017
rect 1160 2005 1162 2017
rect 1240 2005 1242 2017
rect 1352 2005 1354 2017
rect 1456 2005 1458 2017
rect 1560 2005 1562 2017
rect 1656 2005 1658 2017
rect 1744 2005 1746 2017
rect 1824 2005 1826 2017
rect 1896 2005 1898 2017
rect 1960 2005 1962 2017
rect 2024 2005 2026 2017
rect 2072 2005 2074 2017
rect 1158 2004 1164 2005
rect 1158 2000 1159 2004
rect 1163 2000 1164 2004
rect 1158 1999 1164 2000
rect 1238 2004 1244 2005
rect 1238 2000 1239 2004
rect 1243 2000 1244 2004
rect 1238 1999 1244 2000
rect 1350 2004 1356 2005
rect 1350 2000 1351 2004
rect 1355 2000 1356 2004
rect 1350 1999 1356 2000
rect 1454 2004 1460 2005
rect 1454 2000 1455 2004
rect 1459 2000 1460 2004
rect 1454 1999 1460 2000
rect 1558 2004 1564 2005
rect 1558 2000 1559 2004
rect 1563 2000 1564 2004
rect 1558 1999 1564 2000
rect 1654 2004 1660 2005
rect 1654 2000 1655 2004
rect 1659 2000 1660 2004
rect 1654 1999 1660 2000
rect 1742 2004 1748 2005
rect 1742 2000 1743 2004
rect 1747 2000 1748 2004
rect 1742 1999 1748 2000
rect 1822 2004 1828 2005
rect 1822 2000 1823 2004
rect 1827 2000 1828 2004
rect 1822 1999 1828 2000
rect 1894 2004 1900 2005
rect 1894 2000 1895 2004
rect 1899 2000 1900 2004
rect 1894 1999 1900 2000
rect 1958 2004 1964 2005
rect 1958 2000 1959 2004
rect 1963 2000 1964 2004
rect 1958 1999 1964 2000
rect 2022 2004 2028 2005
rect 2022 2000 2023 2004
rect 2027 2000 2028 2004
rect 2022 1999 2028 2000
rect 2070 2004 2076 2005
rect 2070 2000 2071 2004
rect 2075 2000 2076 2004
rect 2070 1999 2076 2000
rect 2120 1997 2122 2017
rect 1094 1994 1100 1995
rect 1134 1996 1140 1997
rect 1046 1991 1052 1992
rect 1096 1991 1098 1994
rect 1134 1992 1135 1996
rect 1139 1992 1140 1996
rect 1134 1991 1140 1992
rect 2118 1996 2124 1997
rect 2118 1992 2119 1996
rect 2123 1992 2124 1996
rect 2118 1991 2124 1992
rect 111 1990 115 1991
rect 111 1985 115 1986
rect 159 1990 163 1991
rect 159 1985 163 1986
rect 183 1990 187 1991
rect 183 1985 187 1986
rect 231 1990 235 1991
rect 231 1985 235 1986
rect 279 1990 283 1991
rect 279 1985 283 1986
rect 303 1990 307 1991
rect 303 1985 307 1986
rect 375 1990 379 1991
rect 375 1985 379 1986
rect 447 1990 451 1991
rect 447 1985 451 1986
rect 463 1990 467 1991
rect 463 1985 467 1986
rect 527 1990 531 1991
rect 527 1985 531 1986
rect 543 1990 547 1991
rect 543 1985 547 1986
rect 607 1990 611 1991
rect 607 1985 611 1986
rect 623 1990 627 1991
rect 623 1985 627 1986
rect 687 1990 691 1991
rect 687 1985 691 1986
rect 695 1990 699 1991
rect 695 1985 699 1986
rect 759 1990 763 1991
rect 759 1985 763 1986
rect 815 1990 819 1991
rect 815 1985 819 1986
rect 831 1990 835 1991
rect 831 1985 835 1986
rect 863 1990 867 1991
rect 863 1985 867 1986
rect 911 1990 915 1991
rect 911 1985 915 1986
rect 959 1990 963 1991
rect 959 1985 963 1986
rect 991 1990 995 1991
rect 991 1985 995 1986
rect 1007 1990 1011 1991
rect 1007 1985 1011 1986
rect 1047 1990 1051 1991
rect 1047 1985 1051 1986
rect 1095 1990 1099 1991
rect 1095 1985 1099 1986
rect 112 1982 114 1985
rect 158 1984 164 1985
rect 110 1981 116 1982
rect 110 1977 111 1981
rect 115 1977 116 1981
rect 158 1980 159 1984
rect 163 1980 164 1984
rect 158 1979 164 1980
rect 230 1984 236 1985
rect 230 1980 231 1984
rect 235 1980 236 1984
rect 230 1979 236 1980
rect 302 1984 308 1985
rect 302 1980 303 1984
rect 307 1980 308 1984
rect 302 1979 308 1980
rect 374 1984 380 1985
rect 374 1980 375 1984
rect 379 1980 380 1984
rect 374 1979 380 1980
rect 446 1984 452 1985
rect 446 1980 447 1984
rect 451 1980 452 1984
rect 446 1979 452 1980
rect 526 1984 532 1985
rect 526 1980 527 1984
rect 531 1980 532 1984
rect 526 1979 532 1980
rect 606 1984 612 1985
rect 606 1980 607 1984
rect 611 1980 612 1984
rect 606 1979 612 1980
rect 686 1984 692 1985
rect 686 1980 687 1984
rect 691 1980 692 1984
rect 686 1979 692 1980
rect 758 1984 764 1985
rect 758 1980 759 1984
rect 763 1980 764 1984
rect 758 1979 764 1980
rect 830 1984 836 1985
rect 830 1980 831 1984
rect 835 1980 836 1984
rect 830 1979 836 1980
rect 910 1984 916 1985
rect 910 1980 911 1984
rect 915 1980 916 1984
rect 910 1979 916 1980
rect 990 1984 996 1985
rect 990 1980 991 1984
rect 995 1980 996 1984
rect 1096 1982 1098 1985
rect 990 1979 996 1980
rect 1094 1981 1100 1982
rect 110 1976 116 1977
rect 1094 1977 1095 1981
rect 1099 1977 1100 1981
rect 1094 1976 1100 1977
rect 1134 1979 1140 1980
rect 1134 1975 1135 1979
rect 1139 1975 1140 1979
rect 2118 1979 2124 1980
rect 1134 1974 1140 1975
rect 1158 1976 1164 1977
rect 110 1964 116 1965
rect 110 1960 111 1964
rect 115 1960 116 1964
rect 110 1959 116 1960
rect 1094 1964 1100 1965
rect 1094 1960 1095 1964
rect 1099 1960 1100 1964
rect 1094 1959 1100 1960
rect 1136 1959 1138 1974
rect 1158 1972 1159 1976
rect 1163 1972 1164 1976
rect 1158 1971 1164 1972
rect 1238 1976 1244 1977
rect 1238 1972 1239 1976
rect 1243 1972 1244 1976
rect 1238 1971 1244 1972
rect 1350 1976 1356 1977
rect 1350 1972 1351 1976
rect 1355 1972 1356 1976
rect 1350 1971 1356 1972
rect 1454 1976 1460 1977
rect 1454 1972 1455 1976
rect 1459 1972 1460 1976
rect 1454 1971 1460 1972
rect 1558 1976 1564 1977
rect 1558 1972 1559 1976
rect 1563 1972 1564 1976
rect 1558 1971 1564 1972
rect 1654 1976 1660 1977
rect 1654 1972 1655 1976
rect 1659 1972 1660 1976
rect 1654 1971 1660 1972
rect 1742 1976 1748 1977
rect 1742 1972 1743 1976
rect 1747 1972 1748 1976
rect 1742 1971 1748 1972
rect 1822 1976 1828 1977
rect 1822 1972 1823 1976
rect 1827 1972 1828 1976
rect 1822 1971 1828 1972
rect 1894 1976 1900 1977
rect 1894 1972 1895 1976
rect 1899 1972 1900 1976
rect 1894 1971 1900 1972
rect 1958 1976 1964 1977
rect 1958 1972 1959 1976
rect 1963 1972 1964 1976
rect 1958 1971 1964 1972
rect 2022 1976 2028 1977
rect 2022 1972 2023 1976
rect 2027 1972 2028 1976
rect 2022 1971 2028 1972
rect 2070 1976 2076 1977
rect 2070 1972 2071 1976
rect 2075 1972 2076 1976
rect 2118 1975 2119 1979
rect 2123 1975 2124 1979
rect 2118 1974 2124 1975
rect 2070 1971 2076 1972
rect 1160 1959 1162 1971
rect 1240 1959 1242 1971
rect 1352 1959 1354 1971
rect 1456 1959 1458 1971
rect 1560 1959 1562 1971
rect 1656 1959 1658 1971
rect 1744 1959 1746 1971
rect 1824 1959 1826 1971
rect 1896 1959 1898 1971
rect 1960 1959 1962 1971
rect 2024 1959 2026 1971
rect 2072 1959 2074 1971
rect 2120 1959 2122 1974
rect 112 1935 114 1959
rect 158 1956 164 1957
rect 158 1952 159 1956
rect 163 1952 164 1956
rect 158 1951 164 1952
rect 230 1956 236 1957
rect 230 1952 231 1956
rect 235 1952 236 1956
rect 230 1951 236 1952
rect 302 1956 308 1957
rect 302 1952 303 1956
rect 307 1952 308 1956
rect 302 1951 308 1952
rect 374 1956 380 1957
rect 374 1952 375 1956
rect 379 1952 380 1956
rect 374 1951 380 1952
rect 446 1956 452 1957
rect 446 1952 447 1956
rect 451 1952 452 1956
rect 446 1951 452 1952
rect 526 1956 532 1957
rect 526 1952 527 1956
rect 531 1952 532 1956
rect 526 1951 532 1952
rect 606 1956 612 1957
rect 606 1952 607 1956
rect 611 1952 612 1956
rect 606 1951 612 1952
rect 686 1956 692 1957
rect 686 1952 687 1956
rect 691 1952 692 1956
rect 686 1951 692 1952
rect 758 1956 764 1957
rect 758 1952 759 1956
rect 763 1952 764 1956
rect 758 1951 764 1952
rect 830 1956 836 1957
rect 830 1952 831 1956
rect 835 1952 836 1956
rect 830 1951 836 1952
rect 910 1956 916 1957
rect 910 1952 911 1956
rect 915 1952 916 1956
rect 910 1951 916 1952
rect 990 1956 996 1957
rect 990 1952 991 1956
rect 995 1952 996 1956
rect 990 1951 996 1952
rect 160 1935 162 1951
rect 232 1935 234 1951
rect 304 1935 306 1951
rect 376 1935 378 1951
rect 448 1935 450 1951
rect 528 1935 530 1951
rect 608 1935 610 1951
rect 688 1935 690 1951
rect 760 1935 762 1951
rect 832 1935 834 1951
rect 912 1935 914 1951
rect 992 1935 994 1951
rect 1096 1935 1098 1959
rect 1135 1958 1139 1959
rect 1135 1953 1139 1954
rect 1159 1958 1163 1959
rect 1159 1953 1163 1954
rect 1239 1958 1243 1959
rect 1239 1953 1243 1954
rect 1351 1958 1355 1959
rect 1351 1953 1355 1954
rect 1359 1958 1363 1959
rect 1359 1953 1363 1954
rect 1423 1958 1427 1959
rect 1423 1953 1427 1954
rect 1455 1958 1459 1959
rect 1455 1953 1459 1954
rect 1487 1958 1491 1959
rect 1487 1953 1491 1954
rect 1559 1958 1563 1959
rect 1559 1953 1563 1954
rect 1631 1958 1635 1959
rect 1631 1953 1635 1954
rect 1655 1958 1659 1959
rect 1655 1953 1659 1954
rect 1703 1958 1707 1959
rect 1703 1953 1707 1954
rect 1743 1958 1747 1959
rect 1743 1953 1747 1954
rect 1775 1958 1779 1959
rect 1775 1953 1779 1954
rect 1823 1958 1827 1959
rect 1823 1953 1827 1954
rect 1847 1958 1851 1959
rect 1847 1953 1851 1954
rect 1895 1958 1899 1959
rect 1895 1953 1899 1954
rect 1927 1958 1931 1959
rect 1927 1953 1931 1954
rect 1959 1958 1963 1959
rect 1959 1953 1963 1954
rect 2007 1958 2011 1959
rect 2007 1953 2011 1954
rect 2023 1958 2027 1959
rect 2023 1953 2027 1954
rect 2071 1958 2075 1959
rect 2071 1953 2075 1954
rect 2119 1958 2123 1959
rect 2119 1953 2123 1954
rect 1136 1950 1138 1953
rect 1358 1952 1364 1953
rect 1134 1949 1140 1950
rect 1134 1945 1135 1949
rect 1139 1945 1140 1949
rect 1358 1948 1359 1952
rect 1363 1948 1364 1952
rect 1358 1947 1364 1948
rect 1422 1952 1428 1953
rect 1422 1948 1423 1952
rect 1427 1948 1428 1952
rect 1422 1947 1428 1948
rect 1486 1952 1492 1953
rect 1486 1948 1487 1952
rect 1491 1948 1492 1952
rect 1486 1947 1492 1948
rect 1558 1952 1564 1953
rect 1558 1948 1559 1952
rect 1563 1948 1564 1952
rect 1558 1947 1564 1948
rect 1630 1952 1636 1953
rect 1630 1948 1631 1952
rect 1635 1948 1636 1952
rect 1630 1947 1636 1948
rect 1702 1952 1708 1953
rect 1702 1948 1703 1952
rect 1707 1948 1708 1952
rect 1702 1947 1708 1948
rect 1774 1952 1780 1953
rect 1774 1948 1775 1952
rect 1779 1948 1780 1952
rect 1774 1947 1780 1948
rect 1846 1952 1852 1953
rect 1846 1948 1847 1952
rect 1851 1948 1852 1952
rect 1846 1947 1852 1948
rect 1926 1952 1932 1953
rect 1926 1948 1927 1952
rect 1931 1948 1932 1952
rect 1926 1947 1932 1948
rect 2006 1952 2012 1953
rect 2006 1948 2007 1952
rect 2011 1948 2012 1952
rect 2006 1947 2012 1948
rect 2070 1952 2076 1953
rect 2070 1948 2071 1952
rect 2075 1948 2076 1952
rect 2120 1950 2122 1953
rect 2070 1947 2076 1948
rect 2118 1949 2124 1950
rect 1134 1944 1140 1945
rect 2118 1945 2119 1949
rect 2123 1945 2124 1949
rect 2118 1944 2124 1945
rect 111 1934 115 1935
rect 111 1929 115 1930
rect 135 1934 139 1935
rect 135 1929 139 1930
rect 159 1934 163 1935
rect 159 1929 163 1930
rect 175 1934 179 1935
rect 175 1929 179 1930
rect 231 1934 235 1935
rect 231 1929 235 1930
rect 295 1934 299 1935
rect 295 1929 299 1930
rect 303 1934 307 1935
rect 303 1929 307 1930
rect 367 1934 371 1935
rect 367 1929 371 1930
rect 375 1934 379 1935
rect 375 1929 379 1930
rect 447 1934 451 1935
rect 447 1929 451 1930
rect 527 1934 531 1935
rect 527 1929 531 1930
rect 607 1934 611 1935
rect 607 1929 611 1930
rect 615 1934 619 1935
rect 615 1929 619 1930
rect 687 1934 691 1935
rect 687 1929 691 1930
rect 703 1934 707 1935
rect 703 1929 707 1930
rect 759 1934 763 1935
rect 759 1929 763 1930
rect 791 1934 795 1935
rect 791 1929 795 1930
rect 831 1934 835 1935
rect 831 1929 835 1930
rect 879 1934 883 1935
rect 879 1929 883 1930
rect 911 1934 915 1935
rect 911 1929 915 1930
rect 991 1934 995 1935
rect 991 1929 995 1930
rect 1095 1934 1099 1935
rect 1095 1929 1099 1930
rect 1134 1932 1140 1933
rect 112 1909 114 1929
rect 136 1917 138 1929
rect 176 1917 178 1929
rect 232 1917 234 1929
rect 296 1917 298 1929
rect 368 1917 370 1929
rect 448 1917 450 1929
rect 528 1917 530 1929
rect 616 1917 618 1929
rect 704 1917 706 1929
rect 792 1917 794 1929
rect 880 1917 882 1929
rect 134 1916 140 1917
rect 134 1912 135 1916
rect 139 1912 140 1916
rect 134 1911 140 1912
rect 174 1916 180 1917
rect 174 1912 175 1916
rect 179 1912 180 1916
rect 174 1911 180 1912
rect 230 1916 236 1917
rect 230 1912 231 1916
rect 235 1912 236 1916
rect 230 1911 236 1912
rect 294 1916 300 1917
rect 294 1912 295 1916
rect 299 1912 300 1916
rect 294 1911 300 1912
rect 366 1916 372 1917
rect 366 1912 367 1916
rect 371 1912 372 1916
rect 366 1911 372 1912
rect 446 1916 452 1917
rect 446 1912 447 1916
rect 451 1912 452 1916
rect 446 1911 452 1912
rect 526 1916 532 1917
rect 526 1912 527 1916
rect 531 1912 532 1916
rect 526 1911 532 1912
rect 614 1916 620 1917
rect 614 1912 615 1916
rect 619 1912 620 1916
rect 614 1911 620 1912
rect 702 1916 708 1917
rect 702 1912 703 1916
rect 707 1912 708 1916
rect 702 1911 708 1912
rect 790 1916 796 1917
rect 790 1912 791 1916
rect 795 1912 796 1916
rect 790 1911 796 1912
rect 878 1916 884 1917
rect 878 1912 879 1916
rect 883 1912 884 1916
rect 878 1911 884 1912
rect 1096 1909 1098 1929
rect 1134 1928 1135 1932
rect 1139 1928 1140 1932
rect 1134 1927 1140 1928
rect 2118 1932 2124 1933
rect 2118 1928 2119 1932
rect 2123 1928 2124 1932
rect 2118 1927 2124 1928
rect 110 1908 116 1909
rect 110 1904 111 1908
rect 115 1904 116 1908
rect 110 1903 116 1904
rect 1094 1908 1100 1909
rect 1094 1904 1095 1908
rect 1099 1904 1100 1908
rect 1136 1907 1138 1927
rect 1358 1924 1364 1925
rect 1358 1920 1359 1924
rect 1363 1920 1364 1924
rect 1358 1919 1364 1920
rect 1422 1924 1428 1925
rect 1422 1920 1423 1924
rect 1427 1920 1428 1924
rect 1422 1919 1428 1920
rect 1486 1924 1492 1925
rect 1486 1920 1487 1924
rect 1491 1920 1492 1924
rect 1486 1919 1492 1920
rect 1558 1924 1564 1925
rect 1558 1920 1559 1924
rect 1563 1920 1564 1924
rect 1558 1919 1564 1920
rect 1630 1924 1636 1925
rect 1630 1920 1631 1924
rect 1635 1920 1636 1924
rect 1630 1919 1636 1920
rect 1702 1924 1708 1925
rect 1702 1920 1703 1924
rect 1707 1920 1708 1924
rect 1702 1919 1708 1920
rect 1774 1924 1780 1925
rect 1774 1920 1775 1924
rect 1779 1920 1780 1924
rect 1774 1919 1780 1920
rect 1846 1924 1852 1925
rect 1846 1920 1847 1924
rect 1851 1920 1852 1924
rect 1846 1919 1852 1920
rect 1926 1924 1932 1925
rect 1926 1920 1927 1924
rect 1931 1920 1932 1924
rect 1926 1919 1932 1920
rect 2006 1924 2012 1925
rect 2006 1920 2007 1924
rect 2011 1920 2012 1924
rect 2006 1919 2012 1920
rect 2070 1924 2076 1925
rect 2070 1920 2071 1924
rect 2075 1920 2076 1924
rect 2070 1919 2076 1920
rect 1360 1907 1362 1919
rect 1424 1907 1426 1919
rect 1488 1907 1490 1919
rect 1560 1907 1562 1919
rect 1632 1907 1634 1919
rect 1704 1907 1706 1919
rect 1776 1907 1778 1919
rect 1848 1907 1850 1919
rect 1928 1907 1930 1919
rect 2008 1907 2010 1919
rect 2072 1907 2074 1919
rect 2120 1907 2122 1927
rect 1094 1903 1100 1904
rect 1135 1906 1139 1907
rect 1135 1901 1139 1902
rect 1231 1906 1235 1907
rect 1231 1901 1235 1902
rect 1271 1906 1275 1907
rect 1271 1901 1275 1902
rect 1319 1906 1323 1907
rect 1319 1901 1323 1902
rect 1359 1906 1363 1907
rect 1359 1901 1363 1902
rect 1375 1906 1379 1907
rect 1375 1901 1379 1902
rect 1423 1906 1427 1907
rect 1423 1901 1427 1902
rect 1439 1906 1443 1907
rect 1439 1901 1443 1902
rect 1487 1906 1491 1907
rect 1487 1901 1491 1902
rect 1503 1906 1507 1907
rect 1503 1901 1507 1902
rect 1559 1906 1563 1907
rect 1559 1901 1563 1902
rect 1575 1906 1579 1907
rect 1575 1901 1579 1902
rect 1631 1906 1635 1907
rect 1631 1901 1635 1902
rect 1655 1906 1659 1907
rect 1655 1901 1659 1902
rect 1703 1906 1707 1907
rect 1703 1901 1707 1902
rect 1751 1906 1755 1907
rect 1751 1901 1755 1902
rect 1775 1906 1779 1907
rect 1775 1901 1779 1902
rect 1847 1906 1851 1907
rect 1847 1901 1851 1902
rect 1863 1906 1867 1907
rect 1863 1901 1867 1902
rect 1927 1906 1931 1907
rect 1927 1901 1931 1902
rect 1975 1906 1979 1907
rect 1975 1901 1979 1902
rect 2007 1906 2011 1907
rect 2007 1901 2011 1902
rect 2071 1906 2075 1907
rect 2071 1901 2075 1902
rect 2119 1906 2123 1907
rect 2119 1901 2123 1902
rect 110 1891 116 1892
rect 110 1887 111 1891
rect 115 1887 116 1891
rect 1094 1891 1100 1892
rect 110 1886 116 1887
rect 134 1888 140 1889
rect 112 1879 114 1886
rect 134 1884 135 1888
rect 139 1884 140 1888
rect 134 1883 140 1884
rect 174 1888 180 1889
rect 174 1884 175 1888
rect 179 1884 180 1888
rect 174 1883 180 1884
rect 230 1888 236 1889
rect 230 1884 231 1888
rect 235 1884 236 1888
rect 230 1883 236 1884
rect 294 1888 300 1889
rect 294 1884 295 1888
rect 299 1884 300 1888
rect 294 1883 300 1884
rect 366 1888 372 1889
rect 366 1884 367 1888
rect 371 1884 372 1888
rect 366 1883 372 1884
rect 446 1888 452 1889
rect 446 1884 447 1888
rect 451 1884 452 1888
rect 446 1883 452 1884
rect 526 1888 532 1889
rect 526 1884 527 1888
rect 531 1884 532 1888
rect 526 1883 532 1884
rect 614 1888 620 1889
rect 614 1884 615 1888
rect 619 1884 620 1888
rect 614 1883 620 1884
rect 702 1888 708 1889
rect 702 1884 703 1888
rect 707 1884 708 1888
rect 702 1883 708 1884
rect 790 1888 796 1889
rect 790 1884 791 1888
rect 795 1884 796 1888
rect 790 1883 796 1884
rect 878 1888 884 1889
rect 878 1884 879 1888
rect 883 1884 884 1888
rect 1094 1887 1095 1891
rect 1099 1887 1100 1891
rect 1094 1886 1100 1887
rect 878 1883 884 1884
rect 136 1879 138 1883
rect 176 1879 178 1883
rect 232 1879 234 1883
rect 296 1879 298 1883
rect 368 1879 370 1883
rect 448 1879 450 1883
rect 528 1879 530 1883
rect 616 1879 618 1883
rect 704 1879 706 1883
rect 792 1879 794 1883
rect 880 1879 882 1883
rect 1096 1879 1098 1886
rect 1136 1881 1138 1901
rect 1232 1889 1234 1901
rect 1272 1889 1274 1901
rect 1320 1889 1322 1901
rect 1376 1889 1378 1901
rect 1440 1889 1442 1901
rect 1504 1889 1506 1901
rect 1576 1889 1578 1901
rect 1656 1889 1658 1901
rect 1752 1889 1754 1901
rect 1864 1889 1866 1901
rect 1976 1889 1978 1901
rect 2072 1889 2074 1901
rect 1230 1888 1236 1889
rect 1230 1884 1231 1888
rect 1235 1884 1236 1888
rect 1230 1883 1236 1884
rect 1270 1888 1276 1889
rect 1270 1884 1271 1888
rect 1275 1884 1276 1888
rect 1270 1883 1276 1884
rect 1318 1888 1324 1889
rect 1318 1884 1319 1888
rect 1323 1884 1324 1888
rect 1318 1883 1324 1884
rect 1374 1888 1380 1889
rect 1374 1884 1375 1888
rect 1379 1884 1380 1888
rect 1374 1883 1380 1884
rect 1438 1888 1444 1889
rect 1438 1884 1439 1888
rect 1443 1884 1444 1888
rect 1438 1883 1444 1884
rect 1502 1888 1508 1889
rect 1502 1884 1503 1888
rect 1507 1884 1508 1888
rect 1502 1883 1508 1884
rect 1574 1888 1580 1889
rect 1574 1884 1575 1888
rect 1579 1884 1580 1888
rect 1574 1883 1580 1884
rect 1654 1888 1660 1889
rect 1654 1884 1655 1888
rect 1659 1884 1660 1888
rect 1654 1883 1660 1884
rect 1750 1888 1756 1889
rect 1750 1884 1751 1888
rect 1755 1884 1756 1888
rect 1750 1883 1756 1884
rect 1862 1888 1868 1889
rect 1862 1884 1863 1888
rect 1867 1884 1868 1888
rect 1862 1883 1868 1884
rect 1974 1888 1980 1889
rect 1974 1884 1975 1888
rect 1979 1884 1980 1888
rect 1974 1883 1980 1884
rect 2070 1888 2076 1889
rect 2070 1884 2071 1888
rect 2075 1884 2076 1888
rect 2070 1883 2076 1884
rect 2120 1881 2122 1901
rect 1134 1880 1140 1881
rect 111 1878 115 1879
rect 111 1873 115 1874
rect 135 1878 139 1879
rect 135 1873 139 1874
rect 175 1878 179 1879
rect 175 1873 179 1874
rect 223 1878 227 1879
rect 223 1873 227 1874
rect 231 1878 235 1879
rect 231 1873 235 1874
rect 287 1878 291 1879
rect 287 1873 291 1874
rect 295 1878 299 1879
rect 295 1873 299 1874
rect 359 1878 363 1879
rect 359 1873 363 1874
rect 367 1878 371 1879
rect 367 1873 371 1874
rect 431 1878 435 1879
rect 431 1873 435 1874
rect 447 1878 451 1879
rect 447 1873 451 1874
rect 503 1878 507 1879
rect 503 1873 507 1874
rect 527 1878 531 1879
rect 527 1873 531 1874
rect 567 1878 571 1879
rect 567 1873 571 1874
rect 615 1878 619 1879
rect 615 1873 619 1874
rect 631 1878 635 1879
rect 631 1873 635 1874
rect 695 1878 699 1879
rect 695 1873 699 1874
rect 703 1878 707 1879
rect 703 1873 707 1874
rect 759 1878 763 1879
rect 759 1873 763 1874
rect 791 1878 795 1879
rect 791 1873 795 1874
rect 831 1878 835 1879
rect 831 1873 835 1874
rect 879 1878 883 1879
rect 879 1873 883 1874
rect 1095 1878 1099 1879
rect 1134 1876 1135 1880
rect 1139 1876 1140 1880
rect 1134 1875 1140 1876
rect 2118 1880 2124 1881
rect 2118 1876 2119 1880
rect 2123 1876 2124 1880
rect 2118 1875 2124 1876
rect 1095 1873 1099 1874
rect 112 1870 114 1873
rect 134 1872 140 1873
rect 110 1869 116 1870
rect 110 1865 111 1869
rect 115 1865 116 1869
rect 134 1868 135 1872
rect 139 1868 140 1872
rect 134 1867 140 1868
rect 174 1872 180 1873
rect 174 1868 175 1872
rect 179 1868 180 1872
rect 174 1867 180 1868
rect 222 1872 228 1873
rect 222 1868 223 1872
rect 227 1868 228 1872
rect 222 1867 228 1868
rect 286 1872 292 1873
rect 286 1868 287 1872
rect 291 1868 292 1872
rect 286 1867 292 1868
rect 358 1872 364 1873
rect 358 1868 359 1872
rect 363 1868 364 1872
rect 358 1867 364 1868
rect 430 1872 436 1873
rect 430 1868 431 1872
rect 435 1868 436 1872
rect 430 1867 436 1868
rect 502 1872 508 1873
rect 502 1868 503 1872
rect 507 1868 508 1872
rect 502 1867 508 1868
rect 566 1872 572 1873
rect 566 1868 567 1872
rect 571 1868 572 1872
rect 566 1867 572 1868
rect 630 1872 636 1873
rect 630 1868 631 1872
rect 635 1868 636 1872
rect 630 1867 636 1868
rect 694 1872 700 1873
rect 694 1868 695 1872
rect 699 1868 700 1872
rect 694 1867 700 1868
rect 758 1872 764 1873
rect 758 1868 759 1872
rect 763 1868 764 1872
rect 758 1867 764 1868
rect 830 1872 836 1873
rect 830 1868 831 1872
rect 835 1868 836 1872
rect 1096 1870 1098 1873
rect 830 1867 836 1868
rect 1094 1869 1100 1870
rect 110 1864 116 1865
rect 1094 1865 1095 1869
rect 1099 1865 1100 1869
rect 1094 1864 1100 1865
rect 1134 1863 1140 1864
rect 1134 1859 1135 1863
rect 1139 1859 1140 1863
rect 2118 1863 2124 1864
rect 1134 1858 1140 1859
rect 1230 1860 1236 1861
rect 110 1852 116 1853
rect 110 1848 111 1852
rect 115 1848 116 1852
rect 110 1847 116 1848
rect 1094 1852 1100 1853
rect 1094 1848 1095 1852
rect 1099 1848 1100 1852
rect 1136 1851 1138 1858
rect 1230 1856 1231 1860
rect 1235 1856 1236 1860
rect 1230 1855 1236 1856
rect 1270 1860 1276 1861
rect 1270 1856 1271 1860
rect 1275 1856 1276 1860
rect 1270 1855 1276 1856
rect 1318 1860 1324 1861
rect 1318 1856 1319 1860
rect 1323 1856 1324 1860
rect 1318 1855 1324 1856
rect 1374 1860 1380 1861
rect 1374 1856 1375 1860
rect 1379 1856 1380 1860
rect 1374 1855 1380 1856
rect 1438 1860 1444 1861
rect 1438 1856 1439 1860
rect 1443 1856 1444 1860
rect 1438 1855 1444 1856
rect 1502 1860 1508 1861
rect 1502 1856 1503 1860
rect 1507 1856 1508 1860
rect 1502 1855 1508 1856
rect 1574 1860 1580 1861
rect 1574 1856 1575 1860
rect 1579 1856 1580 1860
rect 1574 1855 1580 1856
rect 1654 1860 1660 1861
rect 1654 1856 1655 1860
rect 1659 1856 1660 1860
rect 1654 1855 1660 1856
rect 1750 1860 1756 1861
rect 1750 1856 1751 1860
rect 1755 1856 1756 1860
rect 1750 1855 1756 1856
rect 1862 1860 1868 1861
rect 1862 1856 1863 1860
rect 1867 1856 1868 1860
rect 1862 1855 1868 1856
rect 1974 1860 1980 1861
rect 1974 1856 1975 1860
rect 1979 1856 1980 1860
rect 1974 1855 1980 1856
rect 2070 1860 2076 1861
rect 2070 1856 2071 1860
rect 2075 1856 2076 1860
rect 2118 1859 2119 1863
rect 2123 1859 2124 1863
rect 2118 1858 2124 1859
rect 2070 1855 2076 1856
rect 1232 1851 1234 1855
rect 1272 1851 1274 1855
rect 1320 1851 1322 1855
rect 1376 1851 1378 1855
rect 1440 1851 1442 1855
rect 1504 1851 1506 1855
rect 1576 1851 1578 1855
rect 1656 1851 1658 1855
rect 1752 1851 1754 1855
rect 1864 1851 1866 1855
rect 1976 1851 1978 1855
rect 2072 1851 2074 1855
rect 2120 1851 2122 1858
rect 1094 1847 1100 1848
rect 1135 1850 1139 1851
rect 112 1823 114 1847
rect 134 1844 140 1845
rect 134 1840 135 1844
rect 139 1840 140 1844
rect 134 1839 140 1840
rect 174 1844 180 1845
rect 174 1840 175 1844
rect 179 1840 180 1844
rect 174 1839 180 1840
rect 222 1844 228 1845
rect 222 1840 223 1844
rect 227 1840 228 1844
rect 222 1839 228 1840
rect 286 1844 292 1845
rect 286 1840 287 1844
rect 291 1840 292 1844
rect 286 1839 292 1840
rect 358 1844 364 1845
rect 358 1840 359 1844
rect 363 1840 364 1844
rect 358 1839 364 1840
rect 430 1844 436 1845
rect 430 1840 431 1844
rect 435 1840 436 1844
rect 430 1839 436 1840
rect 502 1844 508 1845
rect 502 1840 503 1844
rect 507 1840 508 1844
rect 502 1839 508 1840
rect 566 1844 572 1845
rect 566 1840 567 1844
rect 571 1840 572 1844
rect 566 1839 572 1840
rect 630 1844 636 1845
rect 630 1840 631 1844
rect 635 1840 636 1844
rect 630 1839 636 1840
rect 694 1844 700 1845
rect 694 1840 695 1844
rect 699 1840 700 1844
rect 694 1839 700 1840
rect 758 1844 764 1845
rect 758 1840 759 1844
rect 763 1840 764 1844
rect 758 1839 764 1840
rect 830 1844 836 1845
rect 830 1840 831 1844
rect 835 1840 836 1844
rect 830 1839 836 1840
rect 136 1823 138 1839
rect 176 1823 178 1839
rect 224 1823 226 1839
rect 288 1823 290 1839
rect 360 1823 362 1839
rect 432 1823 434 1839
rect 504 1823 506 1839
rect 568 1823 570 1839
rect 632 1823 634 1839
rect 696 1823 698 1839
rect 760 1823 762 1839
rect 832 1823 834 1839
rect 1096 1823 1098 1847
rect 1135 1845 1139 1846
rect 1159 1850 1163 1851
rect 1159 1845 1163 1846
rect 1199 1850 1203 1851
rect 1199 1845 1203 1846
rect 1231 1850 1235 1851
rect 1231 1845 1235 1846
rect 1239 1850 1243 1851
rect 1239 1845 1243 1846
rect 1271 1850 1275 1851
rect 1271 1845 1275 1846
rect 1303 1850 1307 1851
rect 1303 1845 1307 1846
rect 1319 1850 1323 1851
rect 1319 1845 1323 1846
rect 1367 1850 1371 1851
rect 1367 1845 1371 1846
rect 1375 1850 1379 1851
rect 1375 1845 1379 1846
rect 1431 1850 1435 1851
rect 1431 1845 1435 1846
rect 1439 1850 1443 1851
rect 1439 1845 1443 1846
rect 1503 1850 1507 1851
rect 1503 1845 1507 1846
rect 1575 1850 1579 1851
rect 1575 1845 1579 1846
rect 1583 1850 1587 1851
rect 1583 1845 1587 1846
rect 1655 1850 1659 1851
rect 1655 1845 1659 1846
rect 1671 1850 1675 1851
rect 1671 1845 1675 1846
rect 1751 1850 1755 1851
rect 1751 1845 1755 1846
rect 1767 1850 1771 1851
rect 1767 1845 1771 1846
rect 1863 1850 1867 1851
rect 1863 1845 1867 1846
rect 1871 1850 1875 1851
rect 1871 1845 1875 1846
rect 1975 1850 1979 1851
rect 1975 1845 1979 1846
rect 1983 1850 1987 1851
rect 1983 1845 1987 1846
rect 2071 1850 2075 1851
rect 2071 1845 2075 1846
rect 2119 1850 2123 1851
rect 2119 1845 2123 1846
rect 1136 1842 1138 1845
rect 1158 1844 1164 1845
rect 1134 1841 1140 1842
rect 1134 1837 1135 1841
rect 1139 1837 1140 1841
rect 1158 1840 1159 1844
rect 1163 1840 1164 1844
rect 1158 1839 1164 1840
rect 1198 1844 1204 1845
rect 1198 1840 1199 1844
rect 1203 1840 1204 1844
rect 1198 1839 1204 1840
rect 1238 1844 1244 1845
rect 1238 1840 1239 1844
rect 1243 1840 1244 1844
rect 1238 1839 1244 1840
rect 1302 1844 1308 1845
rect 1302 1840 1303 1844
rect 1307 1840 1308 1844
rect 1302 1839 1308 1840
rect 1366 1844 1372 1845
rect 1366 1840 1367 1844
rect 1371 1840 1372 1844
rect 1366 1839 1372 1840
rect 1430 1844 1436 1845
rect 1430 1840 1431 1844
rect 1435 1840 1436 1844
rect 1430 1839 1436 1840
rect 1502 1844 1508 1845
rect 1502 1840 1503 1844
rect 1507 1840 1508 1844
rect 1502 1839 1508 1840
rect 1582 1844 1588 1845
rect 1582 1840 1583 1844
rect 1587 1840 1588 1844
rect 1582 1839 1588 1840
rect 1670 1844 1676 1845
rect 1670 1840 1671 1844
rect 1675 1840 1676 1844
rect 1670 1839 1676 1840
rect 1766 1844 1772 1845
rect 1766 1840 1767 1844
rect 1771 1840 1772 1844
rect 1766 1839 1772 1840
rect 1870 1844 1876 1845
rect 1870 1840 1871 1844
rect 1875 1840 1876 1844
rect 1870 1839 1876 1840
rect 1982 1844 1988 1845
rect 1982 1840 1983 1844
rect 1987 1840 1988 1844
rect 1982 1839 1988 1840
rect 2070 1844 2076 1845
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2120 1842 2122 1845
rect 2070 1839 2076 1840
rect 2118 1841 2124 1842
rect 1134 1836 1140 1837
rect 2118 1837 2119 1841
rect 2123 1837 2124 1841
rect 2118 1836 2124 1837
rect 1134 1824 1140 1825
rect 111 1822 115 1823
rect 111 1817 115 1818
rect 135 1822 139 1823
rect 135 1817 139 1818
rect 175 1822 179 1823
rect 175 1817 179 1818
rect 183 1822 187 1823
rect 183 1817 187 1818
rect 223 1822 227 1823
rect 223 1817 227 1818
rect 263 1822 267 1823
rect 263 1817 267 1818
rect 287 1822 291 1823
rect 287 1817 291 1818
rect 351 1822 355 1823
rect 351 1817 355 1818
rect 359 1822 363 1823
rect 359 1817 363 1818
rect 431 1822 435 1823
rect 431 1817 435 1818
rect 439 1822 443 1823
rect 439 1817 443 1818
rect 503 1822 507 1823
rect 503 1817 507 1818
rect 527 1822 531 1823
rect 527 1817 531 1818
rect 567 1822 571 1823
rect 567 1817 571 1818
rect 607 1822 611 1823
rect 607 1817 611 1818
rect 631 1822 635 1823
rect 631 1817 635 1818
rect 687 1822 691 1823
rect 687 1817 691 1818
rect 695 1822 699 1823
rect 695 1817 699 1818
rect 759 1822 763 1823
rect 759 1817 763 1818
rect 767 1822 771 1823
rect 767 1817 771 1818
rect 831 1822 835 1823
rect 831 1817 835 1818
rect 839 1822 843 1823
rect 839 1817 843 1818
rect 911 1822 915 1823
rect 911 1817 915 1818
rect 991 1822 995 1823
rect 991 1817 995 1818
rect 1047 1822 1051 1823
rect 1047 1817 1051 1818
rect 1095 1822 1099 1823
rect 1134 1820 1135 1824
rect 1139 1820 1140 1824
rect 1134 1819 1140 1820
rect 2118 1824 2124 1825
rect 2118 1820 2119 1824
rect 2123 1820 2124 1824
rect 2118 1819 2124 1820
rect 1095 1817 1099 1818
rect 112 1797 114 1817
rect 136 1805 138 1817
rect 184 1805 186 1817
rect 264 1805 266 1817
rect 352 1805 354 1817
rect 440 1805 442 1817
rect 528 1805 530 1817
rect 608 1805 610 1817
rect 688 1805 690 1817
rect 768 1805 770 1817
rect 840 1805 842 1817
rect 912 1805 914 1817
rect 992 1805 994 1817
rect 1048 1805 1050 1817
rect 134 1804 140 1805
rect 134 1800 135 1804
rect 139 1800 140 1804
rect 134 1799 140 1800
rect 182 1804 188 1805
rect 182 1800 183 1804
rect 187 1800 188 1804
rect 182 1799 188 1800
rect 262 1804 268 1805
rect 262 1800 263 1804
rect 267 1800 268 1804
rect 262 1799 268 1800
rect 350 1804 356 1805
rect 350 1800 351 1804
rect 355 1800 356 1804
rect 350 1799 356 1800
rect 438 1804 444 1805
rect 438 1800 439 1804
rect 443 1800 444 1804
rect 438 1799 444 1800
rect 526 1804 532 1805
rect 526 1800 527 1804
rect 531 1800 532 1804
rect 526 1799 532 1800
rect 606 1804 612 1805
rect 606 1800 607 1804
rect 611 1800 612 1804
rect 606 1799 612 1800
rect 686 1804 692 1805
rect 686 1800 687 1804
rect 691 1800 692 1804
rect 686 1799 692 1800
rect 766 1804 772 1805
rect 766 1800 767 1804
rect 771 1800 772 1804
rect 766 1799 772 1800
rect 838 1804 844 1805
rect 838 1800 839 1804
rect 843 1800 844 1804
rect 838 1799 844 1800
rect 910 1804 916 1805
rect 910 1800 911 1804
rect 915 1800 916 1804
rect 910 1799 916 1800
rect 990 1804 996 1805
rect 990 1800 991 1804
rect 995 1800 996 1804
rect 990 1799 996 1800
rect 1046 1804 1052 1805
rect 1046 1800 1047 1804
rect 1051 1800 1052 1804
rect 1046 1799 1052 1800
rect 1096 1797 1098 1817
rect 110 1796 116 1797
rect 110 1792 111 1796
rect 115 1792 116 1796
rect 110 1791 116 1792
rect 1094 1796 1100 1797
rect 1094 1792 1095 1796
rect 1099 1792 1100 1796
rect 1094 1791 1100 1792
rect 1136 1791 1138 1819
rect 1158 1816 1164 1817
rect 1158 1812 1159 1816
rect 1163 1812 1164 1816
rect 1158 1811 1164 1812
rect 1198 1816 1204 1817
rect 1198 1812 1199 1816
rect 1203 1812 1204 1816
rect 1198 1811 1204 1812
rect 1238 1816 1244 1817
rect 1238 1812 1239 1816
rect 1243 1812 1244 1816
rect 1238 1811 1244 1812
rect 1302 1816 1308 1817
rect 1302 1812 1303 1816
rect 1307 1812 1308 1816
rect 1302 1811 1308 1812
rect 1366 1816 1372 1817
rect 1366 1812 1367 1816
rect 1371 1812 1372 1816
rect 1366 1811 1372 1812
rect 1430 1816 1436 1817
rect 1430 1812 1431 1816
rect 1435 1812 1436 1816
rect 1430 1811 1436 1812
rect 1502 1816 1508 1817
rect 1502 1812 1503 1816
rect 1507 1812 1508 1816
rect 1502 1811 1508 1812
rect 1582 1816 1588 1817
rect 1582 1812 1583 1816
rect 1587 1812 1588 1816
rect 1582 1811 1588 1812
rect 1670 1816 1676 1817
rect 1670 1812 1671 1816
rect 1675 1812 1676 1816
rect 1670 1811 1676 1812
rect 1766 1816 1772 1817
rect 1766 1812 1767 1816
rect 1771 1812 1772 1816
rect 1766 1811 1772 1812
rect 1870 1816 1876 1817
rect 1870 1812 1871 1816
rect 1875 1812 1876 1816
rect 1870 1811 1876 1812
rect 1982 1816 1988 1817
rect 1982 1812 1983 1816
rect 1987 1812 1988 1816
rect 1982 1811 1988 1812
rect 2070 1816 2076 1817
rect 2070 1812 2071 1816
rect 2075 1812 2076 1816
rect 2070 1811 2076 1812
rect 1160 1791 1162 1811
rect 1200 1791 1202 1811
rect 1240 1791 1242 1811
rect 1304 1791 1306 1811
rect 1368 1791 1370 1811
rect 1432 1791 1434 1811
rect 1504 1791 1506 1811
rect 1584 1791 1586 1811
rect 1672 1791 1674 1811
rect 1768 1791 1770 1811
rect 1872 1791 1874 1811
rect 1984 1791 1986 1811
rect 2072 1791 2074 1811
rect 2120 1791 2122 1819
rect 1135 1790 1139 1791
rect 1135 1785 1139 1786
rect 1159 1790 1163 1791
rect 1159 1785 1163 1786
rect 1199 1790 1203 1791
rect 1199 1785 1203 1786
rect 1239 1790 1243 1791
rect 1239 1785 1243 1786
rect 1303 1790 1307 1791
rect 1303 1785 1307 1786
rect 1311 1790 1315 1791
rect 1311 1785 1315 1786
rect 1351 1790 1355 1791
rect 1351 1785 1355 1786
rect 1367 1790 1371 1791
rect 1367 1785 1371 1786
rect 1391 1790 1395 1791
rect 1391 1785 1395 1786
rect 1431 1790 1435 1791
rect 1431 1785 1435 1786
rect 1471 1790 1475 1791
rect 1471 1785 1475 1786
rect 1503 1790 1507 1791
rect 1503 1785 1507 1786
rect 1511 1790 1515 1791
rect 1511 1785 1515 1786
rect 1551 1790 1555 1791
rect 1551 1785 1555 1786
rect 1583 1790 1587 1791
rect 1583 1785 1587 1786
rect 1607 1790 1611 1791
rect 1607 1785 1611 1786
rect 1671 1790 1675 1791
rect 1671 1785 1675 1786
rect 1679 1790 1683 1791
rect 1679 1785 1683 1786
rect 1767 1790 1771 1791
rect 1767 1785 1771 1786
rect 1871 1790 1875 1791
rect 1871 1785 1875 1786
rect 1983 1790 1987 1791
rect 1983 1785 1987 1786
rect 2071 1790 2075 1791
rect 2071 1785 2075 1786
rect 2119 1790 2123 1791
rect 2119 1785 2123 1786
rect 110 1779 116 1780
rect 110 1775 111 1779
rect 115 1775 116 1779
rect 1094 1779 1100 1780
rect 110 1774 116 1775
rect 134 1776 140 1777
rect 112 1763 114 1774
rect 134 1772 135 1776
rect 139 1772 140 1776
rect 134 1771 140 1772
rect 182 1776 188 1777
rect 182 1772 183 1776
rect 187 1772 188 1776
rect 182 1771 188 1772
rect 262 1776 268 1777
rect 262 1772 263 1776
rect 267 1772 268 1776
rect 262 1771 268 1772
rect 350 1776 356 1777
rect 350 1772 351 1776
rect 355 1772 356 1776
rect 350 1771 356 1772
rect 438 1776 444 1777
rect 438 1772 439 1776
rect 443 1772 444 1776
rect 438 1771 444 1772
rect 526 1776 532 1777
rect 526 1772 527 1776
rect 531 1772 532 1776
rect 526 1771 532 1772
rect 606 1776 612 1777
rect 606 1772 607 1776
rect 611 1772 612 1776
rect 606 1771 612 1772
rect 686 1776 692 1777
rect 686 1772 687 1776
rect 691 1772 692 1776
rect 686 1771 692 1772
rect 766 1776 772 1777
rect 766 1772 767 1776
rect 771 1772 772 1776
rect 766 1771 772 1772
rect 838 1776 844 1777
rect 838 1772 839 1776
rect 843 1772 844 1776
rect 838 1771 844 1772
rect 910 1776 916 1777
rect 910 1772 911 1776
rect 915 1772 916 1776
rect 910 1771 916 1772
rect 990 1776 996 1777
rect 990 1772 991 1776
rect 995 1772 996 1776
rect 990 1771 996 1772
rect 1046 1776 1052 1777
rect 1046 1772 1047 1776
rect 1051 1772 1052 1776
rect 1094 1775 1095 1779
rect 1099 1775 1100 1779
rect 1094 1774 1100 1775
rect 1046 1771 1052 1772
rect 136 1763 138 1771
rect 184 1763 186 1771
rect 264 1763 266 1771
rect 352 1763 354 1771
rect 440 1763 442 1771
rect 528 1763 530 1771
rect 608 1763 610 1771
rect 688 1763 690 1771
rect 768 1763 770 1771
rect 840 1763 842 1771
rect 912 1763 914 1771
rect 992 1763 994 1771
rect 1048 1763 1050 1771
rect 1096 1763 1098 1774
rect 1136 1765 1138 1785
rect 1312 1773 1314 1785
rect 1352 1773 1354 1785
rect 1392 1773 1394 1785
rect 1432 1773 1434 1785
rect 1472 1773 1474 1785
rect 1512 1773 1514 1785
rect 1552 1773 1554 1785
rect 1608 1773 1610 1785
rect 1680 1773 1682 1785
rect 1768 1773 1770 1785
rect 1872 1773 1874 1785
rect 1984 1773 1986 1785
rect 2072 1773 2074 1785
rect 1310 1772 1316 1773
rect 1310 1768 1311 1772
rect 1315 1768 1316 1772
rect 1310 1767 1316 1768
rect 1350 1772 1356 1773
rect 1350 1768 1351 1772
rect 1355 1768 1356 1772
rect 1350 1767 1356 1768
rect 1390 1772 1396 1773
rect 1390 1768 1391 1772
rect 1395 1768 1396 1772
rect 1390 1767 1396 1768
rect 1430 1772 1436 1773
rect 1430 1768 1431 1772
rect 1435 1768 1436 1772
rect 1430 1767 1436 1768
rect 1470 1772 1476 1773
rect 1470 1768 1471 1772
rect 1475 1768 1476 1772
rect 1470 1767 1476 1768
rect 1510 1772 1516 1773
rect 1510 1768 1511 1772
rect 1515 1768 1516 1772
rect 1510 1767 1516 1768
rect 1550 1772 1556 1773
rect 1550 1768 1551 1772
rect 1555 1768 1556 1772
rect 1550 1767 1556 1768
rect 1606 1772 1612 1773
rect 1606 1768 1607 1772
rect 1611 1768 1612 1772
rect 1606 1767 1612 1768
rect 1678 1772 1684 1773
rect 1678 1768 1679 1772
rect 1683 1768 1684 1772
rect 1678 1767 1684 1768
rect 1766 1772 1772 1773
rect 1766 1768 1767 1772
rect 1771 1768 1772 1772
rect 1766 1767 1772 1768
rect 1870 1772 1876 1773
rect 1870 1768 1871 1772
rect 1875 1768 1876 1772
rect 1870 1767 1876 1768
rect 1982 1772 1988 1773
rect 1982 1768 1983 1772
rect 1987 1768 1988 1772
rect 1982 1767 1988 1768
rect 2070 1772 2076 1773
rect 2070 1768 2071 1772
rect 2075 1768 2076 1772
rect 2070 1767 2076 1768
rect 2120 1765 2122 1785
rect 1134 1764 1140 1765
rect 111 1762 115 1763
rect 111 1757 115 1758
rect 135 1762 139 1763
rect 135 1757 139 1758
rect 183 1762 187 1763
rect 183 1757 187 1758
rect 199 1762 203 1763
rect 199 1757 203 1758
rect 263 1762 267 1763
rect 263 1757 267 1758
rect 295 1762 299 1763
rect 295 1757 299 1758
rect 351 1762 355 1763
rect 351 1757 355 1758
rect 399 1762 403 1763
rect 399 1757 403 1758
rect 439 1762 443 1763
rect 439 1757 443 1758
rect 495 1762 499 1763
rect 495 1757 499 1758
rect 527 1762 531 1763
rect 527 1757 531 1758
rect 591 1762 595 1763
rect 591 1757 595 1758
rect 607 1762 611 1763
rect 607 1757 611 1758
rect 671 1762 675 1763
rect 671 1757 675 1758
rect 687 1762 691 1763
rect 687 1757 691 1758
rect 751 1762 755 1763
rect 751 1757 755 1758
rect 767 1762 771 1763
rect 767 1757 771 1758
rect 823 1762 827 1763
rect 823 1757 827 1758
rect 839 1762 843 1763
rect 839 1757 843 1758
rect 887 1762 891 1763
rect 887 1757 891 1758
rect 911 1762 915 1763
rect 911 1757 915 1758
rect 959 1762 963 1763
rect 959 1757 963 1758
rect 991 1762 995 1763
rect 991 1757 995 1758
rect 1031 1762 1035 1763
rect 1031 1757 1035 1758
rect 1047 1762 1051 1763
rect 1047 1757 1051 1758
rect 1095 1762 1099 1763
rect 1134 1760 1135 1764
rect 1139 1760 1140 1764
rect 1134 1759 1140 1760
rect 2118 1764 2124 1765
rect 2118 1760 2119 1764
rect 2123 1760 2124 1764
rect 2118 1759 2124 1760
rect 1095 1757 1099 1758
rect 112 1754 114 1757
rect 134 1756 140 1757
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 134 1752 135 1756
rect 139 1752 140 1756
rect 134 1751 140 1752
rect 198 1756 204 1757
rect 198 1752 199 1756
rect 203 1752 204 1756
rect 198 1751 204 1752
rect 294 1756 300 1757
rect 294 1752 295 1756
rect 299 1752 300 1756
rect 294 1751 300 1752
rect 398 1756 404 1757
rect 398 1752 399 1756
rect 403 1752 404 1756
rect 398 1751 404 1752
rect 494 1756 500 1757
rect 494 1752 495 1756
rect 499 1752 500 1756
rect 494 1751 500 1752
rect 590 1756 596 1757
rect 590 1752 591 1756
rect 595 1752 596 1756
rect 590 1751 596 1752
rect 670 1756 676 1757
rect 670 1752 671 1756
rect 675 1752 676 1756
rect 670 1751 676 1752
rect 750 1756 756 1757
rect 750 1752 751 1756
rect 755 1752 756 1756
rect 750 1751 756 1752
rect 822 1756 828 1757
rect 822 1752 823 1756
rect 827 1752 828 1756
rect 822 1751 828 1752
rect 886 1756 892 1757
rect 886 1752 887 1756
rect 891 1752 892 1756
rect 886 1751 892 1752
rect 958 1756 964 1757
rect 958 1752 959 1756
rect 963 1752 964 1756
rect 958 1751 964 1752
rect 1030 1756 1036 1757
rect 1030 1752 1031 1756
rect 1035 1752 1036 1756
rect 1096 1754 1098 1757
rect 1030 1751 1036 1752
rect 1094 1753 1100 1754
rect 110 1748 116 1749
rect 1094 1749 1095 1753
rect 1099 1749 1100 1753
rect 1094 1748 1100 1749
rect 1134 1747 1140 1748
rect 1134 1743 1135 1747
rect 1139 1743 1140 1747
rect 2118 1747 2124 1748
rect 1134 1742 1140 1743
rect 1310 1744 1316 1745
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 1094 1736 1100 1737
rect 1094 1732 1095 1736
rect 1099 1732 1100 1736
rect 1136 1735 1138 1742
rect 1310 1740 1311 1744
rect 1315 1740 1316 1744
rect 1310 1739 1316 1740
rect 1350 1744 1356 1745
rect 1350 1740 1351 1744
rect 1355 1740 1356 1744
rect 1350 1739 1356 1740
rect 1390 1744 1396 1745
rect 1390 1740 1391 1744
rect 1395 1740 1396 1744
rect 1390 1739 1396 1740
rect 1430 1744 1436 1745
rect 1430 1740 1431 1744
rect 1435 1740 1436 1744
rect 1430 1739 1436 1740
rect 1470 1744 1476 1745
rect 1470 1740 1471 1744
rect 1475 1740 1476 1744
rect 1470 1739 1476 1740
rect 1510 1744 1516 1745
rect 1510 1740 1511 1744
rect 1515 1740 1516 1744
rect 1510 1739 1516 1740
rect 1550 1744 1556 1745
rect 1550 1740 1551 1744
rect 1555 1740 1556 1744
rect 1550 1739 1556 1740
rect 1606 1744 1612 1745
rect 1606 1740 1607 1744
rect 1611 1740 1612 1744
rect 1606 1739 1612 1740
rect 1678 1744 1684 1745
rect 1678 1740 1679 1744
rect 1683 1740 1684 1744
rect 1678 1739 1684 1740
rect 1766 1744 1772 1745
rect 1766 1740 1767 1744
rect 1771 1740 1772 1744
rect 1766 1739 1772 1740
rect 1870 1744 1876 1745
rect 1870 1740 1871 1744
rect 1875 1740 1876 1744
rect 1870 1739 1876 1740
rect 1982 1744 1988 1745
rect 1982 1740 1983 1744
rect 1987 1740 1988 1744
rect 1982 1739 1988 1740
rect 2070 1744 2076 1745
rect 2070 1740 2071 1744
rect 2075 1740 2076 1744
rect 2118 1743 2119 1747
rect 2123 1743 2124 1747
rect 2118 1742 2124 1743
rect 2070 1739 2076 1740
rect 1312 1735 1314 1739
rect 1352 1735 1354 1739
rect 1392 1735 1394 1739
rect 1432 1735 1434 1739
rect 1472 1735 1474 1739
rect 1512 1735 1514 1739
rect 1552 1735 1554 1739
rect 1608 1735 1610 1739
rect 1680 1735 1682 1739
rect 1768 1735 1770 1739
rect 1872 1735 1874 1739
rect 1984 1735 1986 1739
rect 2072 1735 2074 1739
rect 2120 1735 2122 1742
rect 1094 1731 1100 1732
rect 1135 1734 1139 1735
rect 112 1707 114 1731
rect 134 1728 140 1729
rect 134 1724 135 1728
rect 139 1724 140 1728
rect 134 1723 140 1724
rect 198 1728 204 1729
rect 198 1724 199 1728
rect 203 1724 204 1728
rect 198 1723 204 1724
rect 294 1728 300 1729
rect 294 1724 295 1728
rect 299 1724 300 1728
rect 294 1723 300 1724
rect 398 1728 404 1729
rect 398 1724 399 1728
rect 403 1724 404 1728
rect 398 1723 404 1724
rect 494 1728 500 1729
rect 494 1724 495 1728
rect 499 1724 500 1728
rect 494 1723 500 1724
rect 590 1728 596 1729
rect 590 1724 591 1728
rect 595 1724 596 1728
rect 590 1723 596 1724
rect 670 1728 676 1729
rect 670 1724 671 1728
rect 675 1724 676 1728
rect 670 1723 676 1724
rect 750 1728 756 1729
rect 750 1724 751 1728
rect 755 1724 756 1728
rect 750 1723 756 1724
rect 822 1728 828 1729
rect 822 1724 823 1728
rect 827 1724 828 1728
rect 822 1723 828 1724
rect 886 1728 892 1729
rect 886 1724 887 1728
rect 891 1724 892 1728
rect 886 1723 892 1724
rect 958 1728 964 1729
rect 958 1724 959 1728
rect 963 1724 964 1728
rect 958 1723 964 1724
rect 1030 1728 1036 1729
rect 1030 1724 1031 1728
rect 1035 1724 1036 1728
rect 1030 1723 1036 1724
rect 136 1707 138 1723
rect 200 1707 202 1723
rect 296 1707 298 1723
rect 400 1707 402 1723
rect 496 1707 498 1723
rect 592 1707 594 1723
rect 672 1707 674 1723
rect 752 1707 754 1723
rect 824 1707 826 1723
rect 888 1707 890 1723
rect 960 1707 962 1723
rect 1032 1707 1034 1723
rect 1096 1707 1098 1731
rect 1135 1729 1139 1730
rect 1263 1734 1267 1735
rect 1263 1729 1267 1730
rect 1311 1734 1315 1735
rect 1311 1729 1315 1730
rect 1319 1734 1323 1735
rect 1319 1729 1323 1730
rect 1351 1734 1355 1735
rect 1351 1729 1355 1730
rect 1383 1734 1387 1735
rect 1383 1729 1387 1730
rect 1391 1734 1395 1735
rect 1391 1729 1395 1730
rect 1431 1734 1435 1735
rect 1431 1729 1435 1730
rect 1455 1734 1459 1735
rect 1455 1729 1459 1730
rect 1471 1734 1475 1735
rect 1471 1729 1475 1730
rect 1511 1734 1515 1735
rect 1511 1729 1515 1730
rect 1535 1734 1539 1735
rect 1535 1729 1539 1730
rect 1551 1734 1555 1735
rect 1551 1729 1555 1730
rect 1607 1734 1611 1735
rect 1607 1729 1611 1730
rect 1615 1734 1619 1735
rect 1615 1729 1619 1730
rect 1679 1734 1683 1735
rect 1679 1729 1683 1730
rect 1687 1734 1691 1735
rect 1687 1729 1691 1730
rect 1759 1734 1763 1735
rect 1759 1729 1763 1730
rect 1767 1734 1771 1735
rect 1767 1729 1771 1730
rect 1831 1734 1835 1735
rect 1831 1729 1835 1730
rect 1871 1734 1875 1735
rect 1871 1729 1875 1730
rect 1895 1734 1899 1735
rect 1895 1729 1899 1730
rect 1959 1734 1963 1735
rect 1959 1729 1963 1730
rect 1983 1734 1987 1735
rect 1983 1729 1987 1730
rect 2023 1734 2027 1735
rect 2023 1729 2027 1730
rect 2071 1734 2075 1735
rect 2071 1729 2075 1730
rect 2119 1734 2123 1735
rect 2119 1729 2123 1730
rect 1136 1726 1138 1729
rect 1262 1728 1268 1729
rect 1134 1725 1140 1726
rect 1134 1721 1135 1725
rect 1139 1721 1140 1725
rect 1262 1724 1263 1728
rect 1267 1724 1268 1728
rect 1262 1723 1268 1724
rect 1318 1728 1324 1729
rect 1318 1724 1319 1728
rect 1323 1724 1324 1728
rect 1318 1723 1324 1724
rect 1382 1728 1388 1729
rect 1382 1724 1383 1728
rect 1387 1724 1388 1728
rect 1382 1723 1388 1724
rect 1454 1728 1460 1729
rect 1454 1724 1455 1728
rect 1459 1724 1460 1728
rect 1454 1723 1460 1724
rect 1534 1728 1540 1729
rect 1534 1724 1535 1728
rect 1539 1724 1540 1728
rect 1534 1723 1540 1724
rect 1614 1728 1620 1729
rect 1614 1724 1615 1728
rect 1619 1724 1620 1728
rect 1614 1723 1620 1724
rect 1686 1728 1692 1729
rect 1686 1724 1687 1728
rect 1691 1724 1692 1728
rect 1686 1723 1692 1724
rect 1758 1728 1764 1729
rect 1758 1724 1759 1728
rect 1763 1724 1764 1728
rect 1758 1723 1764 1724
rect 1830 1728 1836 1729
rect 1830 1724 1831 1728
rect 1835 1724 1836 1728
rect 1830 1723 1836 1724
rect 1894 1728 1900 1729
rect 1894 1724 1895 1728
rect 1899 1724 1900 1728
rect 1894 1723 1900 1724
rect 1958 1728 1964 1729
rect 1958 1724 1959 1728
rect 1963 1724 1964 1728
rect 1958 1723 1964 1724
rect 2022 1728 2028 1729
rect 2022 1724 2023 1728
rect 2027 1724 2028 1728
rect 2022 1723 2028 1724
rect 2070 1728 2076 1729
rect 2070 1724 2071 1728
rect 2075 1724 2076 1728
rect 2120 1726 2122 1729
rect 2070 1723 2076 1724
rect 2118 1725 2124 1726
rect 1134 1720 1140 1721
rect 2118 1721 2119 1725
rect 2123 1721 2124 1725
rect 2118 1720 2124 1721
rect 1134 1708 1140 1709
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 135 1706 139 1707
rect 135 1701 139 1702
rect 151 1706 155 1707
rect 151 1701 155 1702
rect 199 1706 203 1707
rect 199 1701 203 1702
rect 223 1706 227 1707
rect 223 1701 227 1702
rect 295 1706 299 1707
rect 295 1701 299 1702
rect 303 1706 307 1707
rect 303 1701 307 1702
rect 383 1706 387 1707
rect 383 1701 387 1702
rect 399 1706 403 1707
rect 399 1701 403 1702
rect 463 1706 467 1707
rect 463 1701 467 1702
rect 495 1706 499 1707
rect 495 1701 499 1702
rect 535 1706 539 1707
rect 535 1701 539 1702
rect 591 1706 595 1707
rect 591 1701 595 1702
rect 607 1706 611 1707
rect 607 1701 611 1702
rect 671 1706 675 1707
rect 671 1701 675 1702
rect 735 1706 739 1707
rect 735 1701 739 1702
rect 751 1706 755 1707
rect 751 1701 755 1702
rect 807 1706 811 1707
rect 807 1701 811 1702
rect 823 1706 827 1707
rect 823 1701 827 1702
rect 879 1706 883 1707
rect 879 1701 883 1702
rect 887 1706 891 1707
rect 887 1701 891 1702
rect 959 1706 963 1707
rect 959 1701 963 1702
rect 1031 1706 1035 1707
rect 1031 1701 1035 1702
rect 1095 1706 1099 1707
rect 1134 1704 1135 1708
rect 1139 1704 1140 1708
rect 1134 1703 1140 1704
rect 2118 1708 2124 1709
rect 2118 1704 2119 1708
rect 2123 1704 2124 1708
rect 2118 1703 2124 1704
rect 1095 1701 1099 1702
rect 112 1681 114 1701
rect 152 1689 154 1701
rect 224 1689 226 1701
rect 304 1689 306 1701
rect 384 1689 386 1701
rect 464 1689 466 1701
rect 536 1689 538 1701
rect 608 1689 610 1701
rect 672 1689 674 1701
rect 736 1689 738 1701
rect 808 1689 810 1701
rect 880 1689 882 1701
rect 150 1688 156 1689
rect 150 1684 151 1688
rect 155 1684 156 1688
rect 150 1683 156 1684
rect 222 1688 228 1689
rect 222 1684 223 1688
rect 227 1684 228 1688
rect 222 1683 228 1684
rect 302 1688 308 1689
rect 302 1684 303 1688
rect 307 1684 308 1688
rect 302 1683 308 1684
rect 382 1688 388 1689
rect 382 1684 383 1688
rect 387 1684 388 1688
rect 382 1683 388 1684
rect 462 1688 468 1689
rect 462 1684 463 1688
rect 467 1684 468 1688
rect 462 1683 468 1684
rect 534 1688 540 1689
rect 534 1684 535 1688
rect 539 1684 540 1688
rect 534 1683 540 1684
rect 606 1688 612 1689
rect 606 1684 607 1688
rect 611 1684 612 1688
rect 606 1683 612 1684
rect 670 1688 676 1689
rect 670 1684 671 1688
rect 675 1684 676 1688
rect 670 1683 676 1684
rect 734 1688 740 1689
rect 734 1684 735 1688
rect 739 1684 740 1688
rect 734 1683 740 1684
rect 806 1688 812 1689
rect 806 1684 807 1688
rect 811 1684 812 1688
rect 806 1683 812 1684
rect 878 1688 884 1689
rect 878 1684 879 1688
rect 883 1684 884 1688
rect 878 1683 884 1684
rect 1096 1681 1098 1701
rect 1136 1683 1138 1703
rect 1262 1700 1268 1701
rect 1262 1696 1263 1700
rect 1267 1696 1268 1700
rect 1262 1695 1268 1696
rect 1318 1700 1324 1701
rect 1318 1696 1319 1700
rect 1323 1696 1324 1700
rect 1318 1695 1324 1696
rect 1382 1700 1388 1701
rect 1382 1696 1383 1700
rect 1387 1696 1388 1700
rect 1382 1695 1388 1696
rect 1454 1700 1460 1701
rect 1454 1696 1455 1700
rect 1459 1696 1460 1700
rect 1454 1695 1460 1696
rect 1534 1700 1540 1701
rect 1534 1696 1535 1700
rect 1539 1696 1540 1700
rect 1534 1695 1540 1696
rect 1614 1700 1620 1701
rect 1614 1696 1615 1700
rect 1619 1696 1620 1700
rect 1614 1695 1620 1696
rect 1686 1700 1692 1701
rect 1686 1696 1687 1700
rect 1691 1696 1692 1700
rect 1686 1695 1692 1696
rect 1758 1700 1764 1701
rect 1758 1696 1759 1700
rect 1763 1696 1764 1700
rect 1758 1695 1764 1696
rect 1830 1700 1836 1701
rect 1830 1696 1831 1700
rect 1835 1696 1836 1700
rect 1830 1695 1836 1696
rect 1894 1700 1900 1701
rect 1894 1696 1895 1700
rect 1899 1696 1900 1700
rect 1894 1695 1900 1696
rect 1958 1700 1964 1701
rect 1958 1696 1959 1700
rect 1963 1696 1964 1700
rect 1958 1695 1964 1696
rect 2022 1700 2028 1701
rect 2022 1696 2023 1700
rect 2027 1696 2028 1700
rect 2022 1695 2028 1696
rect 2070 1700 2076 1701
rect 2070 1696 2071 1700
rect 2075 1696 2076 1700
rect 2070 1695 2076 1696
rect 1264 1683 1266 1695
rect 1320 1683 1322 1695
rect 1384 1683 1386 1695
rect 1456 1683 1458 1695
rect 1536 1683 1538 1695
rect 1616 1683 1618 1695
rect 1688 1683 1690 1695
rect 1760 1683 1762 1695
rect 1832 1683 1834 1695
rect 1896 1683 1898 1695
rect 1960 1683 1962 1695
rect 2024 1683 2026 1695
rect 2072 1683 2074 1695
rect 2120 1683 2122 1703
rect 1135 1682 1139 1683
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 1094 1680 1100 1681
rect 1094 1676 1095 1680
rect 1099 1676 1100 1680
rect 1135 1677 1139 1678
rect 1167 1682 1171 1683
rect 1167 1677 1171 1678
rect 1247 1682 1251 1683
rect 1247 1677 1251 1678
rect 1263 1682 1267 1683
rect 1263 1677 1267 1678
rect 1319 1682 1323 1683
rect 1319 1677 1323 1678
rect 1335 1682 1339 1683
rect 1335 1677 1339 1678
rect 1383 1682 1387 1683
rect 1383 1677 1387 1678
rect 1423 1682 1427 1683
rect 1423 1677 1427 1678
rect 1455 1682 1459 1683
rect 1455 1677 1459 1678
rect 1511 1682 1515 1683
rect 1511 1677 1515 1678
rect 1535 1682 1539 1683
rect 1535 1677 1539 1678
rect 1599 1682 1603 1683
rect 1599 1677 1603 1678
rect 1615 1682 1619 1683
rect 1615 1677 1619 1678
rect 1679 1682 1683 1683
rect 1679 1677 1683 1678
rect 1687 1682 1691 1683
rect 1687 1677 1691 1678
rect 1751 1682 1755 1683
rect 1751 1677 1755 1678
rect 1759 1682 1763 1683
rect 1759 1677 1763 1678
rect 1815 1682 1819 1683
rect 1815 1677 1819 1678
rect 1831 1682 1835 1683
rect 1831 1677 1835 1678
rect 1871 1682 1875 1683
rect 1871 1677 1875 1678
rect 1895 1682 1899 1683
rect 1895 1677 1899 1678
rect 1927 1682 1931 1683
rect 1927 1677 1931 1678
rect 1959 1682 1963 1683
rect 1959 1677 1963 1678
rect 1983 1682 1987 1683
rect 1983 1677 1987 1678
rect 2023 1682 2027 1683
rect 2023 1677 2027 1678
rect 2031 1682 2035 1683
rect 2031 1677 2035 1678
rect 2071 1682 2075 1683
rect 2071 1677 2075 1678
rect 2119 1682 2123 1683
rect 2119 1677 2123 1678
rect 1094 1675 1100 1676
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 1094 1663 1100 1664
rect 110 1658 116 1659
rect 150 1660 156 1661
rect 112 1651 114 1658
rect 150 1656 151 1660
rect 155 1656 156 1660
rect 150 1655 156 1656
rect 222 1660 228 1661
rect 222 1656 223 1660
rect 227 1656 228 1660
rect 222 1655 228 1656
rect 302 1660 308 1661
rect 302 1656 303 1660
rect 307 1656 308 1660
rect 302 1655 308 1656
rect 382 1660 388 1661
rect 382 1656 383 1660
rect 387 1656 388 1660
rect 382 1655 388 1656
rect 462 1660 468 1661
rect 462 1656 463 1660
rect 467 1656 468 1660
rect 462 1655 468 1656
rect 534 1660 540 1661
rect 534 1656 535 1660
rect 539 1656 540 1660
rect 534 1655 540 1656
rect 606 1660 612 1661
rect 606 1656 607 1660
rect 611 1656 612 1660
rect 606 1655 612 1656
rect 670 1660 676 1661
rect 670 1656 671 1660
rect 675 1656 676 1660
rect 670 1655 676 1656
rect 734 1660 740 1661
rect 734 1656 735 1660
rect 739 1656 740 1660
rect 734 1655 740 1656
rect 806 1660 812 1661
rect 806 1656 807 1660
rect 811 1656 812 1660
rect 806 1655 812 1656
rect 878 1660 884 1661
rect 878 1656 879 1660
rect 883 1656 884 1660
rect 1094 1659 1095 1663
rect 1099 1659 1100 1663
rect 1094 1658 1100 1659
rect 878 1655 884 1656
rect 152 1651 154 1655
rect 224 1651 226 1655
rect 304 1651 306 1655
rect 384 1651 386 1655
rect 464 1651 466 1655
rect 536 1651 538 1655
rect 608 1651 610 1655
rect 672 1651 674 1655
rect 736 1651 738 1655
rect 808 1651 810 1655
rect 880 1651 882 1655
rect 1096 1651 1098 1658
rect 1136 1657 1138 1677
rect 1168 1665 1170 1677
rect 1248 1665 1250 1677
rect 1336 1665 1338 1677
rect 1424 1665 1426 1677
rect 1512 1665 1514 1677
rect 1600 1665 1602 1677
rect 1680 1665 1682 1677
rect 1752 1665 1754 1677
rect 1816 1665 1818 1677
rect 1872 1665 1874 1677
rect 1928 1665 1930 1677
rect 1984 1665 1986 1677
rect 2032 1665 2034 1677
rect 2072 1665 2074 1677
rect 1166 1664 1172 1665
rect 1166 1660 1167 1664
rect 1171 1660 1172 1664
rect 1166 1659 1172 1660
rect 1246 1664 1252 1665
rect 1246 1660 1247 1664
rect 1251 1660 1252 1664
rect 1246 1659 1252 1660
rect 1334 1664 1340 1665
rect 1334 1660 1335 1664
rect 1339 1660 1340 1664
rect 1334 1659 1340 1660
rect 1422 1664 1428 1665
rect 1422 1660 1423 1664
rect 1427 1660 1428 1664
rect 1422 1659 1428 1660
rect 1510 1664 1516 1665
rect 1510 1660 1511 1664
rect 1515 1660 1516 1664
rect 1510 1659 1516 1660
rect 1598 1664 1604 1665
rect 1598 1660 1599 1664
rect 1603 1660 1604 1664
rect 1598 1659 1604 1660
rect 1678 1664 1684 1665
rect 1678 1660 1679 1664
rect 1683 1660 1684 1664
rect 1678 1659 1684 1660
rect 1750 1664 1756 1665
rect 1750 1660 1751 1664
rect 1755 1660 1756 1664
rect 1750 1659 1756 1660
rect 1814 1664 1820 1665
rect 1814 1660 1815 1664
rect 1819 1660 1820 1664
rect 1814 1659 1820 1660
rect 1870 1664 1876 1665
rect 1870 1660 1871 1664
rect 1875 1660 1876 1664
rect 1870 1659 1876 1660
rect 1926 1664 1932 1665
rect 1926 1660 1927 1664
rect 1931 1660 1932 1664
rect 1926 1659 1932 1660
rect 1982 1664 1988 1665
rect 1982 1660 1983 1664
rect 1987 1660 1988 1664
rect 1982 1659 1988 1660
rect 2030 1664 2036 1665
rect 2030 1660 2031 1664
rect 2035 1660 2036 1664
rect 2030 1659 2036 1660
rect 2070 1664 2076 1665
rect 2070 1660 2071 1664
rect 2075 1660 2076 1664
rect 2070 1659 2076 1660
rect 2120 1657 2122 1677
rect 1134 1656 1140 1657
rect 1134 1652 1135 1656
rect 1139 1652 1140 1656
rect 1134 1651 1140 1652
rect 2118 1656 2124 1657
rect 2118 1652 2119 1656
rect 2123 1652 2124 1656
rect 2118 1651 2124 1652
rect 111 1650 115 1651
rect 111 1645 115 1646
rect 151 1650 155 1651
rect 151 1645 155 1646
rect 175 1650 179 1651
rect 175 1645 179 1646
rect 215 1650 219 1651
rect 215 1645 219 1646
rect 223 1650 227 1651
rect 223 1645 227 1646
rect 255 1650 259 1651
rect 255 1645 259 1646
rect 303 1650 307 1651
rect 303 1645 307 1646
rect 359 1650 363 1651
rect 359 1645 363 1646
rect 383 1650 387 1651
rect 383 1645 387 1646
rect 407 1650 411 1651
rect 407 1645 411 1646
rect 455 1650 459 1651
rect 455 1645 459 1646
rect 463 1650 467 1651
rect 463 1645 467 1646
rect 503 1650 507 1651
rect 503 1645 507 1646
rect 535 1650 539 1651
rect 535 1645 539 1646
rect 551 1650 555 1651
rect 551 1645 555 1646
rect 607 1650 611 1651
rect 607 1645 611 1646
rect 663 1650 667 1651
rect 663 1645 667 1646
rect 671 1650 675 1651
rect 671 1645 675 1646
rect 719 1650 723 1651
rect 719 1645 723 1646
rect 735 1650 739 1651
rect 735 1645 739 1646
rect 807 1650 811 1651
rect 807 1645 811 1646
rect 879 1650 883 1651
rect 879 1645 883 1646
rect 1095 1650 1099 1651
rect 1095 1645 1099 1646
rect 112 1642 114 1645
rect 174 1644 180 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 174 1640 175 1644
rect 179 1640 180 1644
rect 174 1639 180 1640
rect 214 1644 220 1645
rect 214 1640 215 1644
rect 219 1640 220 1644
rect 214 1639 220 1640
rect 254 1644 260 1645
rect 254 1640 255 1644
rect 259 1640 260 1644
rect 254 1639 260 1640
rect 302 1644 308 1645
rect 302 1640 303 1644
rect 307 1640 308 1644
rect 302 1639 308 1640
rect 358 1644 364 1645
rect 358 1640 359 1644
rect 363 1640 364 1644
rect 358 1639 364 1640
rect 406 1644 412 1645
rect 406 1640 407 1644
rect 411 1640 412 1644
rect 406 1639 412 1640
rect 454 1644 460 1645
rect 454 1640 455 1644
rect 459 1640 460 1644
rect 454 1639 460 1640
rect 502 1644 508 1645
rect 502 1640 503 1644
rect 507 1640 508 1644
rect 502 1639 508 1640
rect 550 1644 556 1645
rect 550 1640 551 1644
rect 555 1640 556 1644
rect 550 1639 556 1640
rect 606 1644 612 1645
rect 606 1640 607 1644
rect 611 1640 612 1644
rect 606 1639 612 1640
rect 662 1644 668 1645
rect 662 1640 663 1644
rect 667 1640 668 1644
rect 662 1639 668 1640
rect 718 1644 724 1645
rect 718 1640 719 1644
rect 723 1640 724 1644
rect 1096 1642 1098 1645
rect 718 1639 724 1640
rect 1094 1641 1100 1642
rect 110 1636 116 1637
rect 1094 1637 1095 1641
rect 1099 1637 1100 1641
rect 1094 1636 1100 1637
rect 1134 1639 1140 1640
rect 1134 1635 1135 1639
rect 1139 1635 1140 1639
rect 2118 1639 2124 1640
rect 1134 1634 1140 1635
rect 1166 1636 1172 1637
rect 1136 1627 1138 1634
rect 1166 1632 1167 1636
rect 1171 1632 1172 1636
rect 1166 1631 1172 1632
rect 1246 1636 1252 1637
rect 1246 1632 1247 1636
rect 1251 1632 1252 1636
rect 1246 1631 1252 1632
rect 1334 1636 1340 1637
rect 1334 1632 1335 1636
rect 1339 1632 1340 1636
rect 1334 1631 1340 1632
rect 1422 1636 1428 1637
rect 1422 1632 1423 1636
rect 1427 1632 1428 1636
rect 1422 1631 1428 1632
rect 1510 1636 1516 1637
rect 1510 1632 1511 1636
rect 1515 1632 1516 1636
rect 1510 1631 1516 1632
rect 1598 1636 1604 1637
rect 1598 1632 1599 1636
rect 1603 1632 1604 1636
rect 1598 1631 1604 1632
rect 1678 1636 1684 1637
rect 1678 1632 1679 1636
rect 1683 1632 1684 1636
rect 1678 1631 1684 1632
rect 1750 1636 1756 1637
rect 1750 1632 1751 1636
rect 1755 1632 1756 1636
rect 1750 1631 1756 1632
rect 1814 1636 1820 1637
rect 1814 1632 1815 1636
rect 1819 1632 1820 1636
rect 1814 1631 1820 1632
rect 1870 1636 1876 1637
rect 1870 1632 1871 1636
rect 1875 1632 1876 1636
rect 1870 1631 1876 1632
rect 1926 1636 1932 1637
rect 1926 1632 1927 1636
rect 1931 1632 1932 1636
rect 1926 1631 1932 1632
rect 1982 1636 1988 1637
rect 1982 1632 1983 1636
rect 1987 1632 1988 1636
rect 1982 1631 1988 1632
rect 2030 1636 2036 1637
rect 2030 1632 2031 1636
rect 2035 1632 2036 1636
rect 2030 1631 2036 1632
rect 2070 1636 2076 1637
rect 2070 1632 2071 1636
rect 2075 1632 2076 1636
rect 2118 1635 2119 1639
rect 2123 1635 2124 1639
rect 2118 1634 2124 1635
rect 2070 1631 2076 1632
rect 1168 1627 1170 1631
rect 1248 1627 1250 1631
rect 1336 1627 1338 1631
rect 1424 1627 1426 1631
rect 1512 1627 1514 1631
rect 1600 1627 1602 1631
rect 1680 1627 1682 1631
rect 1752 1627 1754 1631
rect 1816 1627 1818 1631
rect 1872 1627 1874 1631
rect 1928 1627 1930 1631
rect 1984 1627 1986 1631
rect 2032 1627 2034 1631
rect 2072 1627 2074 1631
rect 2120 1627 2122 1634
rect 1135 1626 1139 1627
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 1094 1624 1100 1625
rect 1094 1620 1095 1624
rect 1099 1620 1100 1624
rect 1135 1621 1139 1622
rect 1159 1626 1163 1627
rect 1159 1621 1163 1622
rect 1167 1626 1171 1627
rect 1167 1621 1171 1622
rect 1199 1626 1203 1627
rect 1199 1621 1203 1622
rect 1247 1626 1251 1627
rect 1247 1621 1251 1622
rect 1319 1626 1323 1627
rect 1319 1621 1323 1622
rect 1335 1626 1339 1627
rect 1335 1621 1339 1622
rect 1391 1626 1395 1627
rect 1391 1621 1395 1622
rect 1423 1626 1427 1627
rect 1423 1621 1427 1622
rect 1463 1626 1467 1627
rect 1463 1621 1467 1622
rect 1511 1626 1515 1627
rect 1511 1621 1515 1622
rect 1535 1626 1539 1627
rect 1535 1621 1539 1622
rect 1599 1626 1603 1627
rect 1599 1621 1603 1622
rect 1607 1626 1611 1627
rect 1607 1621 1611 1622
rect 1679 1626 1683 1627
rect 1679 1621 1683 1622
rect 1751 1626 1755 1627
rect 1751 1621 1755 1622
rect 1815 1626 1819 1627
rect 1815 1621 1819 1622
rect 1831 1626 1835 1627
rect 1831 1621 1835 1622
rect 1871 1626 1875 1627
rect 1871 1621 1875 1622
rect 1927 1626 1931 1627
rect 1927 1621 1931 1622
rect 1983 1626 1987 1627
rect 1983 1621 1987 1622
rect 2031 1626 2035 1627
rect 2031 1621 2035 1622
rect 2071 1626 2075 1627
rect 2071 1621 2075 1622
rect 2119 1626 2123 1627
rect 2119 1621 2123 1622
rect 1094 1619 1100 1620
rect 112 1591 114 1619
rect 174 1616 180 1617
rect 174 1612 175 1616
rect 179 1612 180 1616
rect 174 1611 180 1612
rect 214 1616 220 1617
rect 214 1612 215 1616
rect 219 1612 220 1616
rect 214 1611 220 1612
rect 254 1616 260 1617
rect 254 1612 255 1616
rect 259 1612 260 1616
rect 254 1611 260 1612
rect 302 1616 308 1617
rect 302 1612 303 1616
rect 307 1612 308 1616
rect 302 1611 308 1612
rect 358 1616 364 1617
rect 358 1612 359 1616
rect 363 1612 364 1616
rect 358 1611 364 1612
rect 406 1616 412 1617
rect 406 1612 407 1616
rect 411 1612 412 1616
rect 406 1611 412 1612
rect 454 1616 460 1617
rect 454 1612 455 1616
rect 459 1612 460 1616
rect 454 1611 460 1612
rect 502 1616 508 1617
rect 502 1612 503 1616
rect 507 1612 508 1616
rect 502 1611 508 1612
rect 550 1616 556 1617
rect 550 1612 551 1616
rect 555 1612 556 1616
rect 550 1611 556 1612
rect 606 1616 612 1617
rect 606 1612 607 1616
rect 611 1612 612 1616
rect 606 1611 612 1612
rect 662 1616 668 1617
rect 662 1612 663 1616
rect 667 1612 668 1616
rect 662 1611 668 1612
rect 718 1616 724 1617
rect 718 1612 719 1616
rect 723 1612 724 1616
rect 718 1611 724 1612
rect 176 1591 178 1611
rect 216 1591 218 1611
rect 256 1591 258 1611
rect 304 1591 306 1611
rect 360 1591 362 1611
rect 408 1591 410 1611
rect 456 1591 458 1611
rect 504 1591 506 1611
rect 552 1591 554 1611
rect 608 1591 610 1611
rect 664 1591 666 1611
rect 720 1591 722 1611
rect 1096 1591 1098 1619
rect 1136 1618 1138 1621
rect 1158 1620 1164 1621
rect 1134 1617 1140 1618
rect 1134 1613 1135 1617
rect 1139 1613 1140 1617
rect 1158 1616 1159 1620
rect 1163 1616 1164 1620
rect 1158 1615 1164 1616
rect 1198 1620 1204 1621
rect 1198 1616 1199 1620
rect 1203 1616 1204 1620
rect 1198 1615 1204 1616
rect 1246 1620 1252 1621
rect 1246 1616 1247 1620
rect 1251 1616 1252 1620
rect 1246 1615 1252 1616
rect 1318 1620 1324 1621
rect 1318 1616 1319 1620
rect 1323 1616 1324 1620
rect 1318 1615 1324 1616
rect 1390 1620 1396 1621
rect 1390 1616 1391 1620
rect 1395 1616 1396 1620
rect 1390 1615 1396 1616
rect 1462 1620 1468 1621
rect 1462 1616 1463 1620
rect 1467 1616 1468 1620
rect 1462 1615 1468 1616
rect 1534 1620 1540 1621
rect 1534 1616 1535 1620
rect 1539 1616 1540 1620
rect 1534 1615 1540 1616
rect 1606 1620 1612 1621
rect 1606 1616 1607 1620
rect 1611 1616 1612 1620
rect 1606 1615 1612 1616
rect 1678 1620 1684 1621
rect 1678 1616 1679 1620
rect 1683 1616 1684 1620
rect 1678 1615 1684 1616
rect 1750 1620 1756 1621
rect 1750 1616 1751 1620
rect 1755 1616 1756 1620
rect 1750 1615 1756 1616
rect 1830 1620 1836 1621
rect 1830 1616 1831 1620
rect 1835 1616 1836 1620
rect 2120 1618 2122 1621
rect 1830 1615 1836 1616
rect 2118 1617 2124 1618
rect 1134 1612 1140 1613
rect 2118 1613 2119 1617
rect 2123 1613 2124 1617
rect 2118 1612 2124 1613
rect 1134 1600 1140 1601
rect 1134 1596 1135 1600
rect 1139 1596 1140 1600
rect 1134 1595 1140 1596
rect 2118 1600 2124 1601
rect 2118 1596 2119 1600
rect 2123 1596 2124 1600
rect 2118 1595 2124 1596
rect 111 1590 115 1591
rect 111 1585 115 1586
rect 143 1590 147 1591
rect 143 1585 147 1586
rect 175 1590 179 1591
rect 175 1585 179 1586
rect 183 1590 187 1591
rect 183 1585 187 1586
rect 215 1590 219 1591
rect 215 1585 219 1586
rect 231 1590 235 1591
rect 231 1585 235 1586
rect 255 1590 259 1591
rect 255 1585 259 1586
rect 287 1590 291 1591
rect 287 1585 291 1586
rect 303 1590 307 1591
rect 303 1585 307 1586
rect 351 1590 355 1591
rect 351 1585 355 1586
rect 359 1590 363 1591
rect 359 1585 363 1586
rect 407 1590 411 1591
rect 407 1585 411 1586
rect 415 1590 419 1591
rect 415 1585 419 1586
rect 455 1590 459 1591
rect 455 1585 459 1586
rect 479 1590 483 1591
rect 479 1585 483 1586
rect 503 1590 507 1591
rect 503 1585 507 1586
rect 543 1590 547 1591
rect 543 1585 547 1586
rect 551 1590 555 1591
rect 551 1585 555 1586
rect 607 1590 611 1591
rect 607 1585 611 1586
rect 663 1590 667 1591
rect 663 1585 667 1586
rect 719 1590 723 1591
rect 719 1585 723 1586
rect 727 1590 731 1591
rect 727 1585 731 1586
rect 791 1590 795 1591
rect 791 1585 795 1586
rect 855 1590 859 1591
rect 855 1585 859 1586
rect 1095 1590 1099 1591
rect 1095 1585 1099 1586
rect 112 1565 114 1585
rect 144 1573 146 1585
rect 184 1573 186 1585
rect 232 1573 234 1585
rect 288 1573 290 1585
rect 352 1573 354 1585
rect 416 1573 418 1585
rect 480 1573 482 1585
rect 544 1573 546 1585
rect 608 1573 610 1585
rect 664 1573 666 1585
rect 728 1573 730 1585
rect 792 1573 794 1585
rect 856 1573 858 1585
rect 142 1572 148 1573
rect 142 1568 143 1572
rect 147 1568 148 1572
rect 142 1567 148 1568
rect 182 1572 188 1573
rect 182 1568 183 1572
rect 187 1568 188 1572
rect 182 1567 188 1568
rect 230 1572 236 1573
rect 230 1568 231 1572
rect 235 1568 236 1572
rect 230 1567 236 1568
rect 286 1572 292 1573
rect 286 1568 287 1572
rect 291 1568 292 1572
rect 286 1567 292 1568
rect 350 1572 356 1573
rect 350 1568 351 1572
rect 355 1568 356 1572
rect 350 1567 356 1568
rect 414 1572 420 1573
rect 414 1568 415 1572
rect 419 1568 420 1572
rect 414 1567 420 1568
rect 478 1572 484 1573
rect 478 1568 479 1572
rect 483 1568 484 1572
rect 478 1567 484 1568
rect 542 1572 548 1573
rect 542 1568 543 1572
rect 547 1568 548 1572
rect 542 1567 548 1568
rect 606 1572 612 1573
rect 606 1568 607 1572
rect 611 1568 612 1572
rect 606 1567 612 1568
rect 662 1572 668 1573
rect 662 1568 663 1572
rect 667 1568 668 1572
rect 662 1567 668 1568
rect 726 1572 732 1573
rect 726 1568 727 1572
rect 731 1568 732 1572
rect 726 1567 732 1568
rect 790 1572 796 1573
rect 790 1568 791 1572
rect 795 1568 796 1572
rect 790 1567 796 1568
rect 854 1572 860 1573
rect 854 1568 855 1572
rect 859 1568 860 1572
rect 854 1567 860 1568
rect 1096 1565 1098 1585
rect 1136 1575 1138 1595
rect 1158 1592 1164 1593
rect 1158 1588 1159 1592
rect 1163 1588 1164 1592
rect 1158 1587 1164 1588
rect 1198 1592 1204 1593
rect 1198 1588 1199 1592
rect 1203 1588 1204 1592
rect 1198 1587 1204 1588
rect 1246 1592 1252 1593
rect 1246 1588 1247 1592
rect 1251 1588 1252 1592
rect 1246 1587 1252 1588
rect 1318 1592 1324 1593
rect 1318 1588 1319 1592
rect 1323 1588 1324 1592
rect 1318 1587 1324 1588
rect 1390 1592 1396 1593
rect 1390 1588 1391 1592
rect 1395 1588 1396 1592
rect 1390 1587 1396 1588
rect 1462 1592 1468 1593
rect 1462 1588 1463 1592
rect 1467 1588 1468 1592
rect 1462 1587 1468 1588
rect 1534 1592 1540 1593
rect 1534 1588 1535 1592
rect 1539 1588 1540 1592
rect 1534 1587 1540 1588
rect 1606 1592 1612 1593
rect 1606 1588 1607 1592
rect 1611 1588 1612 1592
rect 1606 1587 1612 1588
rect 1678 1592 1684 1593
rect 1678 1588 1679 1592
rect 1683 1588 1684 1592
rect 1678 1587 1684 1588
rect 1750 1592 1756 1593
rect 1750 1588 1751 1592
rect 1755 1588 1756 1592
rect 1750 1587 1756 1588
rect 1830 1592 1836 1593
rect 1830 1588 1831 1592
rect 1835 1588 1836 1592
rect 1830 1587 1836 1588
rect 1160 1575 1162 1587
rect 1200 1575 1202 1587
rect 1248 1575 1250 1587
rect 1320 1575 1322 1587
rect 1392 1575 1394 1587
rect 1464 1575 1466 1587
rect 1536 1575 1538 1587
rect 1608 1575 1610 1587
rect 1680 1575 1682 1587
rect 1752 1575 1754 1587
rect 1832 1575 1834 1587
rect 2120 1575 2122 1595
rect 1135 1574 1139 1575
rect 1135 1569 1139 1570
rect 1159 1574 1163 1575
rect 1159 1569 1163 1570
rect 1199 1574 1203 1575
rect 1199 1569 1203 1570
rect 1239 1574 1243 1575
rect 1239 1569 1243 1570
rect 1247 1574 1251 1575
rect 1247 1569 1251 1570
rect 1279 1574 1283 1575
rect 1279 1569 1283 1570
rect 1319 1574 1323 1575
rect 1319 1569 1323 1570
rect 1327 1574 1331 1575
rect 1327 1569 1331 1570
rect 1375 1574 1379 1575
rect 1375 1569 1379 1570
rect 1391 1574 1395 1575
rect 1391 1569 1395 1570
rect 1423 1574 1427 1575
rect 1423 1569 1427 1570
rect 1463 1574 1467 1575
rect 1463 1569 1467 1570
rect 1471 1574 1475 1575
rect 1471 1569 1475 1570
rect 1519 1574 1523 1575
rect 1519 1569 1523 1570
rect 1535 1574 1539 1575
rect 1535 1569 1539 1570
rect 1567 1574 1571 1575
rect 1567 1569 1571 1570
rect 1607 1574 1611 1575
rect 1607 1569 1611 1570
rect 1623 1574 1627 1575
rect 1623 1569 1627 1570
rect 1679 1574 1683 1575
rect 1679 1569 1683 1570
rect 1735 1574 1739 1575
rect 1735 1569 1739 1570
rect 1751 1574 1755 1575
rect 1751 1569 1755 1570
rect 1831 1574 1835 1575
rect 1831 1569 1835 1570
rect 2119 1574 2123 1575
rect 2119 1569 2123 1570
rect 110 1564 116 1565
rect 110 1560 111 1564
rect 115 1560 116 1564
rect 110 1559 116 1560
rect 1094 1564 1100 1565
rect 1094 1560 1095 1564
rect 1099 1560 1100 1564
rect 1094 1559 1100 1560
rect 1136 1549 1138 1569
rect 1240 1557 1242 1569
rect 1280 1557 1282 1569
rect 1328 1557 1330 1569
rect 1376 1557 1378 1569
rect 1424 1557 1426 1569
rect 1472 1557 1474 1569
rect 1520 1557 1522 1569
rect 1568 1557 1570 1569
rect 1624 1557 1626 1569
rect 1680 1557 1682 1569
rect 1736 1557 1738 1569
rect 1238 1556 1244 1557
rect 1238 1552 1239 1556
rect 1243 1552 1244 1556
rect 1238 1551 1244 1552
rect 1278 1556 1284 1557
rect 1278 1552 1279 1556
rect 1283 1552 1284 1556
rect 1278 1551 1284 1552
rect 1326 1556 1332 1557
rect 1326 1552 1327 1556
rect 1331 1552 1332 1556
rect 1326 1551 1332 1552
rect 1374 1556 1380 1557
rect 1374 1552 1375 1556
rect 1379 1552 1380 1556
rect 1374 1551 1380 1552
rect 1422 1556 1428 1557
rect 1422 1552 1423 1556
rect 1427 1552 1428 1556
rect 1422 1551 1428 1552
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1518 1556 1524 1557
rect 1518 1552 1519 1556
rect 1523 1552 1524 1556
rect 1518 1551 1524 1552
rect 1566 1556 1572 1557
rect 1566 1552 1567 1556
rect 1571 1552 1572 1556
rect 1566 1551 1572 1552
rect 1622 1556 1628 1557
rect 1622 1552 1623 1556
rect 1627 1552 1628 1556
rect 1622 1551 1628 1552
rect 1678 1556 1684 1557
rect 1678 1552 1679 1556
rect 1683 1552 1684 1556
rect 1678 1551 1684 1552
rect 1734 1556 1740 1557
rect 1734 1552 1735 1556
rect 1739 1552 1740 1556
rect 1734 1551 1740 1552
rect 2120 1549 2122 1569
rect 1134 1548 1140 1549
rect 110 1547 116 1548
rect 110 1543 111 1547
rect 115 1543 116 1547
rect 1094 1547 1100 1548
rect 110 1542 116 1543
rect 142 1544 148 1545
rect 112 1531 114 1542
rect 142 1540 143 1544
rect 147 1540 148 1544
rect 142 1539 148 1540
rect 182 1544 188 1545
rect 182 1540 183 1544
rect 187 1540 188 1544
rect 182 1539 188 1540
rect 230 1544 236 1545
rect 230 1540 231 1544
rect 235 1540 236 1544
rect 230 1539 236 1540
rect 286 1544 292 1545
rect 286 1540 287 1544
rect 291 1540 292 1544
rect 286 1539 292 1540
rect 350 1544 356 1545
rect 350 1540 351 1544
rect 355 1540 356 1544
rect 350 1539 356 1540
rect 414 1544 420 1545
rect 414 1540 415 1544
rect 419 1540 420 1544
rect 414 1539 420 1540
rect 478 1544 484 1545
rect 478 1540 479 1544
rect 483 1540 484 1544
rect 478 1539 484 1540
rect 542 1544 548 1545
rect 542 1540 543 1544
rect 547 1540 548 1544
rect 542 1539 548 1540
rect 606 1544 612 1545
rect 606 1540 607 1544
rect 611 1540 612 1544
rect 606 1539 612 1540
rect 662 1544 668 1545
rect 662 1540 663 1544
rect 667 1540 668 1544
rect 662 1539 668 1540
rect 726 1544 732 1545
rect 726 1540 727 1544
rect 731 1540 732 1544
rect 726 1539 732 1540
rect 790 1544 796 1545
rect 790 1540 791 1544
rect 795 1540 796 1544
rect 790 1539 796 1540
rect 854 1544 860 1545
rect 854 1540 855 1544
rect 859 1540 860 1544
rect 1094 1543 1095 1547
rect 1099 1543 1100 1547
rect 1134 1544 1135 1548
rect 1139 1544 1140 1548
rect 1134 1543 1140 1544
rect 2118 1548 2124 1549
rect 2118 1544 2119 1548
rect 2123 1544 2124 1548
rect 2118 1543 2124 1544
rect 1094 1542 1100 1543
rect 854 1539 860 1540
rect 144 1531 146 1539
rect 184 1531 186 1539
rect 232 1531 234 1539
rect 288 1531 290 1539
rect 352 1531 354 1539
rect 416 1531 418 1539
rect 480 1531 482 1539
rect 544 1531 546 1539
rect 608 1531 610 1539
rect 664 1531 666 1539
rect 728 1531 730 1539
rect 792 1531 794 1539
rect 856 1531 858 1539
rect 1096 1531 1098 1542
rect 1134 1531 1140 1532
rect 111 1530 115 1531
rect 111 1525 115 1526
rect 135 1530 139 1531
rect 135 1525 139 1526
rect 143 1530 147 1531
rect 143 1525 147 1526
rect 175 1530 179 1531
rect 175 1525 179 1526
rect 183 1530 187 1531
rect 183 1525 187 1526
rect 215 1530 219 1531
rect 215 1525 219 1526
rect 231 1530 235 1531
rect 231 1525 235 1526
rect 255 1530 259 1531
rect 255 1525 259 1526
rect 287 1530 291 1531
rect 287 1525 291 1526
rect 295 1530 299 1531
rect 295 1525 299 1526
rect 335 1530 339 1531
rect 335 1525 339 1526
rect 351 1530 355 1531
rect 351 1525 355 1526
rect 375 1530 379 1531
rect 375 1525 379 1526
rect 415 1530 419 1531
rect 415 1525 419 1526
rect 455 1530 459 1531
rect 455 1525 459 1526
rect 479 1530 483 1531
rect 479 1525 483 1526
rect 495 1530 499 1531
rect 495 1525 499 1526
rect 535 1530 539 1531
rect 535 1525 539 1526
rect 543 1530 547 1531
rect 543 1525 547 1526
rect 575 1530 579 1531
rect 575 1525 579 1526
rect 607 1530 611 1531
rect 607 1525 611 1526
rect 615 1530 619 1531
rect 615 1525 619 1526
rect 655 1530 659 1531
rect 655 1525 659 1526
rect 663 1530 667 1531
rect 663 1525 667 1526
rect 695 1530 699 1531
rect 695 1525 699 1526
rect 727 1530 731 1531
rect 727 1525 731 1526
rect 735 1530 739 1531
rect 735 1525 739 1526
rect 775 1530 779 1531
rect 775 1525 779 1526
rect 791 1530 795 1531
rect 791 1525 795 1526
rect 831 1530 835 1531
rect 831 1525 835 1526
rect 855 1530 859 1531
rect 855 1525 859 1526
rect 887 1530 891 1531
rect 887 1525 891 1526
rect 1095 1530 1099 1531
rect 1134 1527 1135 1531
rect 1139 1527 1140 1531
rect 2118 1531 2124 1532
rect 1134 1526 1140 1527
rect 1238 1528 1244 1529
rect 1095 1525 1099 1526
rect 112 1522 114 1525
rect 134 1524 140 1525
rect 110 1521 116 1522
rect 110 1517 111 1521
rect 115 1517 116 1521
rect 134 1520 135 1524
rect 139 1520 140 1524
rect 134 1519 140 1520
rect 174 1524 180 1525
rect 174 1520 175 1524
rect 179 1520 180 1524
rect 174 1519 180 1520
rect 214 1524 220 1525
rect 214 1520 215 1524
rect 219 1520 220 1524
rect 214 1519 220 1520
rect 254 1524 260 1525
rect 254 1520 255 1524
rect 259 1520 260 1524
rect 254 1519 260 1520
rect 294 1524 300 1525
rect 294 1520 295 1524
rect 299 1520 300 1524
rect 294 1519 300 1520
rect 334 1524 340 1525
rect 334 1520 335 1524
rect 339 1520 340 1524
rect 334 1519 340 1520
rect 374 1524 380 1525
rect 374 1520 375 1524
rect 379 1520 380 1524
rect 374 1519 380 1520
rect 414 1524 420 1525
rect 414 1520 415 1524
rect 419 1520 420 1524
rect 414 1519 420 1520
rect 454 1524 460 1525
rect 454 1520 455 1524
rect 459 1520 460 1524
rect 454 1519 460 1520
rect 494 1524 500 1525
rect 494 1520 495 1524
rect 499 1520 500 1524
rect 494 1519 500 1520
rect 534 1524 540 1525
rect 534 1520 535 1524
rect 539 1520 540 1524
rect 534 1519 540 1520
rect 574 1524 580 1525
rect 574 1520 575 1524
rect 579 1520 580 1524
rect 574 1519 580 1520
rect 614 1524 620 1525
rect 614 1520 615 1524
rect 619 1520 620 1524
rect 614 1519 620 1520
rect 654 1524 660 1525
rect 654 1520 655 1524
rect 659 1520 660 1524
rect 654 1519 660 1520
rect 694 1524 700 1525
rect 694 1520 695 1524
rect 699 1520 700 1524
rect 694 1519 700 1520
rect 734 1524 740 1525
rect 734 1520 735 1524
rect 739 1520 740 1524
rect 734 1519 740 1520
rect 774 1524 780 1525
rect 774 1520 775 1524
rect 779 1520 780 1524
rect 774 1519 780 1520
rect 830 1524 836 1525
rect 830 1520 831 1524
rect 835 1520 836 1524
rect 830 1519 836 1520
rect 886 1524 892 1525
rect 886 1520 887 1524
rect 891 1520 892 1524
rect 1096 1522 1098 1525
rect 886 1519 892 1520
rect 1094 1521 1100 1522
rect 110 1516 116 1517
rect 1094 1517 1095 1521
rect 1099 1517 1100 1521
rect 1136 1519 1138 1526
rect 1238 1524 1239 1528
rect 1243 1524 1244 1528
rect 1238 1523 1244 1524
rect 1278 1528 1284 1529
rect 1278 1524 1279 1528
rect 1283 1524 1284 1528
rect 1278 1523 1284 1524
rect 1326 1528 1332 1529
rect 1326 1524 1327 1528
rect 1331 1524 1332 1528
rect 1326 1523 1332 1524
rect 1374 1528 1380 1529
rect 1374 1524 1375 1528
rect 1379 1524 1380 1528
rect 1374 1523 1380 1524
rect 1422 1528 1428 1529
rect 1422 1524 1423 1528
rect 1427 1524 1428 1528
rect 1422 1523 1428 1524
rect 1470 1528 1476 1529
rect 1470 1524 1471 1528
rect 1475 1524 1476 1528
rect 1470 1523 1476 1524
rect 1518 1528 1524 1529
rect 1518 1524 1519 1528
rect 1523 1524 1524 1528
rect 1518 1523 1524 1524
rect 1566 1528 1572 1529
rect 1566 1524 1567 1528
rect 1571 1524 1572 1528
rect 1566 1523 1572 1524
rect 1622 1528 1628 1529
rect 1622 1524 1623 1528
rect 1627 1524 1628 1528
rect 1622 1523 1628 1524
rect 1678 1528 1684 1529
rect 1678 1524 1679 1528
rect 1683 1524 1684 1528
rect 1678 1523 1684 1524
rect 1734 1528 1740 1529
rect 1734 1524 1735 1528
rect 1739 1524 1740 1528
rect 2118 1527 2119 1531
rect 2123 1527 2124 1531
rect 2118 1526 2124 1527
rect 1734 1523 1740 1524
rect 1240 1519 1242 1523
rect 1280 1519 1282 1523
rect 1328 1519 1330 1523
rect 1376 1519 1378 1523
rect 1424 1519 1426 1523
rect 1472 1519 1474 1523
rect 1520 1519 1522 1523
rect 1568 1519 1570 1523
rect 1624 1519 1626 1523
rect 1680 1519 1682 1523
rect 1736 1519 1738 1523
rect 2120 1519 2122 1526
rect 1094 1516 1100 1517
rect 1135 1518 1139 1519
rect 1135 1513 1139 1514
rect 1239 1518 1243 1519
rect 1239 1513 1243 1514
rect 1279 1518 1283 1519
rect 1279 1513 1283 1514
rect 1319 1518 1323 1519
rect 1319 1513 1323 1514
rect 1327 1518 1331 1519
rect 1327 1513 1331 1514
rect 1359 1518 1363 1519
rect 1359 1513 1363 1514
rect 1375 1518 1379 1519
rect 1375 1513 1379 1514
rect 1399 1518 1403 1519
rect 1399 1513 1403 1514
rect 1423 1518 1427 1519
rect 1423 1513 1427 1514
rect 1439 1518 1443 1519
rect 1439 1513 1443 1514
rect 1471 1518 1475 1519
rect 1471 1513 1475 1514
rect 1479 1518 1483 1519
rect 1479 1513 1483 1514
rect 1519 1518 1523 1519
rect 1519 1513 1523 1514
rect 1559 1518 1563 1519
rect 1559 1513 1563 1514
rect 1567 1518 1571 1519
rect 1567 1513 1571 1514
rect 1607 1518 1611 1519
rect 1607 1513 1611 1514
rect 1623 1518 1627 1519
rect 1623 1513 1627 1514
rect 1663 1518 1667 1519
rect 1663 1513 1667 1514
rect 1679 1518 1683 1519
rect 1679 1513 1683 1514
rect 1735 1518 1739 1519
rect 1735 1513 1739 1514
rect 1815 1518 1819 1519
rect 1815 1513 1819 1514
rect 1903 1518 1907 1519
rect 1903 1513 1907 1514
rect 1991 1518 1995 1519
rect 1991 1513 1995 1514
rect 2071 1518 2075 1519
rect 2071 1513 2075 1514
rect 2119 1518 2123 1519
rect 2119 1513 2123 1514
rect 1136 1510 1138 1513
rect 1318 1512 1324 1513
rect 1134 1509 1140 1510
rect 1134 1505 1135 1509
rect 1139 1505 1140 1509
rect 1318 1508 1319 1512
rect 1323 1508 1324 1512
rect 1318 1507 1324 1508
rect 1358 1512 1364 1513
rect 1358 1508 1359 1512
rect 1363 1508 1364 1512
rect 1358 1507 1364 1508
rect 1398 1512 1404 1513
rect 1398 1508 1399 1512
rect 1403 1508 1404 1512
rect 1398 1507 1404 1508
rect 1438 1512 1444 1513
rect 1438 1508 1439 1512
rect 1443 1508 1444 1512
rect 1438 1507 1444 1508
rect 1478 1512 1484 1513
rect 1478 1508 1479 1512
rect 1483 1508 1484 1512
rect 1478 1507 1484 1508
rect 1518 1512 1524 1513
rect 1518 1508 1519 1512
rect 1523 1508 1524 1512
rect 1518 1507 1524 1508
rect 1558 1512 1564 1513
rect 1558 1508 1559 1512
rect 1563 1508 1564 1512
rect 1558 1507 1564 1508
rect 1606 1512 1612 1513
rect 1606 1508 1607 1512
rect 1611 1508 1612 1512
rect 1606 1507 1612 1508
rect 1662 1512 1668 1513
rect 1662 1508 1663 1512
rect 1667 1508 1668 1512
rect 1662 1507 1668 1508
rect 1734 1512 1740 1513
rect 1734 1508 1735 1512
rect 1739 1508 1740 1512
rect 1734 1507 1740 1508
rect 1814 1512 1820 1513
rect 1814 1508 1815 1512
rect 1819 1508 1820 1512
rect 1814 1507 1820 1508
rect 1902 1512 1908 1513
rect 1902 1508 1903 1512
rect 1907 1508 1908 1512
rect 1902 1507 1908 1508
rect 1990 1512 1996 1513
rect 1990 1508 1991 1512
rect 1995 1508 1996 1512
rect 1990 1507 1996 1508
rect 2070 1512 2076 1513
rect 2070 1508 2071 1512
rect 2075 1508 2076 1512
rect 2120 1510 2122 1513
rect 2070 1507 2076 1508
rect 2118 1509 2124 1510
rect 110 1504 116 1505
rect 110 1500 111 1504
rect 115 1500 116 1504
rect 110 1499 116 1500
rect 1094 1504 1100 1505
rect 1134 1504 1140 1505
rect 2118 1505 2119 1509
rect 2123 1505 2124 1509
rect 2118 1504 2124 1505
rect 1094 1500 1095 1504
rect 1099 1500 1100 1504
rect 1094 1499 1100 1500
rect 112 1471 114 1499
rect 134 1496 140 1497
rect 134 1492 135 1496
rect 139 1492 140 1496
rect 134 1491 140 1492
rect 174 1496 180 1497
rect 174 1492 175 1496
rect 179 1492 180 1496
rect 174 1491 180 1492
rect 214 1496 220 1497
rect 214 1492 215 1496
rect 219 1492 220 1496
rect 214 1491 220 1492
rect 254 1496 260 1497
rect 254 1492 255 1496
rect 259 1492 260 1496
rect 254 1491 260 1492
rect 294 1496 300 1497
rect 294 1492 295 1496
rect 299 1492 300 1496
rect 294 1491 300 1492
rect 334 1496 340 1497
rect 334 1492 335 1496
rect 339 1492 340 1496
rect 334 1491 340 1492
rect 374 1496 380 1497
rect 374 1492 375 1496
rect 379 1492 380 1496
rect 374 1491 380 1492
rect 414 1496 420 1497
rect 414 1492 415 1496
rect 419 1492 420 1496
rect 414 1491 420 1492
rect 454 1496 460 1497
rect 454 1492 455 1496
rect 459 1492 460 1496
rect 454 1491 460 1492
rect 494 1496 500 1497
rect 494 1492 495 1496
rect 499 1492 500 1496
rect 494 1491 500 1492
rect 534 1496 540 1497
rect 534 1492 535 1496
rect 539 1492 540 1496
rect 534 1491 540 1492
rect 574 1496 580 1497
rect 574 1492 575 1496
rect 579 1492 580 1496
rect 574 1491 580 1492
rect 614 1496 620 1497
rect 614 1492 615 1496
rect 619 1492 620 1496
rect 614 1491 620 1492
rect 654 1496 660 1497
rect 654 1492 655 1496
rect 659 1492 660 1496
rect 654 1491 660 1492
rect 694 1496 700 1497
rect 694 1492 695 1496
rect 699 1492 700 1496
rect 694 1491 700 1492
rect 734 1496 740 1497
rect 734 1492 735 1496
rect 739 1492 740 1496
rect 734 1491 740 1492
rect 774 1496 780 1497
rect 774 1492 775 1496
rect 779 1492 780 1496
rect 774 1491 780 1492
rect 830 1496 836 1497
rect 830 1492 831 1496
rect 835 1492 836 1496
rect 830 1491 836 1492
rect 886 1496 892 1497
rect 886 1492 887 1496
rect 891 1492 892 1496
rect 886 1491 892 1492
rect 136 1471 138 1491
rect 176 1471 178 1491
rect 216 1471 218 1491
rect 256 1471 258 1491
rect 296 1471 298 1491
rect 336 1471 338 1491
rect 376 1471 378 1491
rect 416 1471 418 1491
rect 456 1471 458 1491
rect 496 1471 498 1491
rect 536 1471 538 1491
rect 576 1471 578 1491
rect 616 1471 618 1491
rect 656 1471 658 1491
rect 696 1471 698 1491
rect 736 1471 738 1491
rect 776 1471 778 1491
rect 832 1471 834 1491
rect 888 1471 890 1491
rect 1096 1471 1098 1499
rect 1134 1492 1140 1493
rect 1134 1488 1135 1492
rect 1139 1488 1140 1492
rect 1134 1487 1140 1488
rect 2118 1492 2124 1493
rect 2118 1488 2119 1492
rect 2123 1488 2124 1492
rect 2118 1487 2124 1488
rect 111 1470 115 1471
rect 111 1465 115 1466
rect 135 1470 139 1471
rect 135 1465 139 1466
rect 175 1470 179 1471
rect 175 1465 179 1466
rect 215 1470 219 1471
rect 215 1465 219 1466
rect 255 1470 259 1471
rect 255 1465 259 1466
rect 295 1470 299 1471
rect 295 1465 299 1466
rect 335 1470 339 1471
rect 335 1465 339 1466
rect 375 1470 379 1471
rect 375 1465 379 1466
rect 415 1470 419 1471
rect 415 1465 419 1466
rect 455 1470 459 1471
rect 455 1465 459 1466
rect 495 1470 499 1471
rect 495 1465 499 1466
rect 519 1470 523 1471
rect 519 1465 523 1466
rect 535 1470 539 1471
rect 535 1465 539 1466
rect 559 1470 563 1471
rect 559 1465 563 1466
rect 575 1470 579 1471
rect 575 1465 579 1466
rect 599 1470 603 1471
rect 599 1465 603 1466
rect 615 1470 619 1471
rect 615 1465 619 1466
rect 647 1470 651 1471
rect 647 1465 651 1466
rect 655 1470 659 1471
rect 655 1465 659 1466
rect 695 1470 699 1471
rect 695 1465 699 1466
rect 735 1470 739 1471
rect 735 1465 739 1466
rect 751 1470 755 1471
rect 751 1465 755 1466
rect 775 1470 779 1471
rect 775 1465 779 1466
rect 807 1470 811 1471
rect 807 1465 811 1466
rect 831 1470 835 1471
rect 831 1465 835 1466
rect 871 1470 875 1471
rect 871 1465 875 1466
rect 887 1470 891 1471
rect 887 1465 891 1466
rect 935 1470 939 1471
rect 935 1465 939 1466
rect 1095 1470 1099 1471
rect 1136 1467 1138 1487
rect 1318 1484 1324 1485
rect 1318 1480 1319 1484
rect 1323 1480 1324 1484
rect 1318 1479 1324 1480
rect 1358 1484 1364 1485
rect 1358 1480 1359 1484
rect 1363 1480 1364 1484
rect 1358 1479 1364 1480
rect 1398 1484 1404 1485
rect 1398 1480 1399 1484
rect 1403 1480 1404 1484
rect 1398 1479 1404 1480
rect 1438 1484 1444 1485
rect 1438 1480 1439 1484
rect 1443 1480 1444 1484
rect 1438 1479 1444 1480
rect 1478 1484 1484 1485
rect 1478 1480 1479 1484
rect 1483 1480 1484 1484
rect 1478 1479 1484 1480
rect 1518 1484 1524 1485
rect 1518 1480 1519 1484
rect 1523 1480 1524 1484
rect 1518 1479 1524 1480
rect 1558 1484 1564 1485
rect 1558 1480 1559 1484
rect 1563 1480 1564 1484
rect 1558 1479 1564 1480
rect 1606 1484 1612 1485
rect 1606 1480 1607 1484
rect 1611 1480 1612 1484
rect 1606 1479 1612 1480
rect 1662 1484 1668 1485
rect 1662 1480 1663 1484
rect 1667 1480 1668 1484
rect 1662 1479 1668 1480
rect 1734 1484 1740 1485
rect 1734 1480 1735 1484
rect 1739 1480 1740 1484
rect 1734 1479 1740 1480
rect 1814 1484 1820 1485
rect 1814 1480 1815 1484
rect 1819 1480 1820 1484
rect 1814 1479 1820 1480
rect 1902 1484 1908 1485
rect 1902 1480 1903 1484
rect 1907 1480 1908 1484
rect 1902 1479 1908 1480
rect 1990 1484 1996 1485
rect 1990 1480 1991 1484
rect 1995 1480 1996 1484
rect 1990 1479 1996 1480
rect 2070 1484 2076 1485
rect 2070 1480 2071 1484
rect 2075 1480 2076 1484
rect 2070 1479 2076 1480
rect 1320 1467 1322 1479
rect 1360 1467 1362 1479
rect 1400 1467 1402 1479
rect 1440 1467 1442 1479
rect 1480 1467 1482 1479
rect 1520 1467 1522 1479
rect 1560 1467 1562 1479
rect 1608 1467 1610 1479
rect 1664 1467 1666 1479
rect 1736 1467 1738 1479
rect 1816 1467 1818 1479
rect 1904 1467 1906 1479
rect 1992 1467 1994 1479
rect 2072 1467 2074 1479
rect 2120 1467 2122 1487
rect 1095 1465 1099 1466
rect 1135 1466 1139 1467
rect 112 1445 114 1465
rect 520 1453 522 1465
rect 560 1453 562 1465
rect 600 1453 602 1465
rect 648 1453 650 1465
rect 696 1453 698 1465
rect 752 1453 754 1465
rect 808 1453 810 1465
rect 872 1453 874 1465
rect 936 1453 938 1465
rect 518 1452 524 1453
rect 518 1448 519 1452
rect 523 1448 524 1452
rect 518 1447 524 1448
rect 558 1452 564 1453
rect 558 1448 559 1452
rect 563 1448 564 1452
rect 558 1447 564 1448
rect 598 1452 604 1453
rect 598 1448 599 1452
rect 603 1448 604 1452
rect 598 1447 604 1448
rect 646 1452 652 1453
rect 646 1448 647 1452
rect 651 1448 652 1452
rect 646 1447 652 1448
rect 694 1452 700 1453
rect 694 1448 695 1452
rect 699 1448 700 1452
rect 694 1447 700 1448
rect 750 1452 756 1453
rect 750 1448 751 1452
rect 755 1448 756 1452
rect 750 1447 756 1448
rect 806 1452 812 1453
rect 806 1448 807 1452
rect 811 1448 812 1452
rect 806 1447 812 1448
rect 870 1452 876 1453
rect 870 1448 871 1452
rect 875 1448 876 1452
rect 870 1447 876 1448
rect 934 1452 940 1453
rect 934 1448 935 1452
rect 939 1448 940 1452
rect 934 1447 940 1448
rect 1096 1445 1098 1465
rect 1135 1461 1139 1462
rect 1231 1466 1235 1467
rect 1231 1461 1235 1462
rect 1279 1466 1283 1467
rect 1279 1461 1283 1462
rect 1319 1466 1323 1467
rect 1319 1461 1323 1462
rect 1335 1466 1339 1467
rect 1335 1461 1339 1462
rect 1359 1466 1363 1467
rect 1359 1461 1363 1462
rect 1391 1466 1395 1467
rect 1391 1461 1395 1462
rect 1399 1466 1403 1467
rect 1399 1461 1403 1462
rect 1439 1466 1443 1467
rect 1439 1461 1443 1462
rect 1455 1466 1459 1467
rect 1455 1461 1459 1462
rect 1479 1466 1483 1467
rect 1479 1461 1483 1462
rect 1519 1466 1523 1467
rect 1519 1461 1523 1462
rect 1559 1466 1563 1467
rect 1559 1461 1563 1462
rect 1583 1466 1587 1467
rect 1583 1461 1587 1462
rect 1607 1466 1611 1467
rect 1607 1461 1611 1462
rect 1647 1466 1651 1467
rect 1647 1461 1651 1462
rect 1663 1466 1667 1467
rect 1663 1461 1667 1462
rect 1719 1466 1723 1467
rect 1719 1461 1723 1462
rect 1735 1466 1739 1467
rect 1735 1461 1739 1462
rect 1807 1466 1811 1467
rect 1807 1461 1811 1462
rect 1815 1466 1819 1467
rect 1815 1461 1819 1462
rect 1895 1466 1899 1467
rect 1895 1461 1899 1462
rect 1903 1466 1907 1467
rect 1903 1461 1907 1462
rect 1991 1466 1995 1467
rect 1991 1461 1995 1462
rect 2071 1466 2075 1467
rect 2071 1461 2075 1462
rect 2119 1466 2123 1467
rect 2119 1461 2123 1462
rect 110 1444 116 1445
rect 110 1440 111 1444
rect 115 1440 116 1444
rect 110 1439 116 1440
rect 1094 1444 1100 1445
rect 1094 1440 1095 1444
rect 1099 1440 1100 1444
rect 1136 1441 1138 1461
rect 1232 1449 1234 1461
rect 1280 1449 1282 1461
rect 1336 1449 1338 1461
rect 1392 1449 1394 1461
rect 1456 1449 1458 1461
rect 1520 1449 1522 1461
rect 1584 1449 1586 1461
rect 1648 1449 1650 1461
rect 1720 1449 1722 1461
rect 1808 1449 1810 1461
rect 1896 1449 1898 1461
rect 1992 1449 1994 1461
rect 2072 1449 2074 1461
rect 1230 1448 1236 1449
rect 1230 1444 1231 1448
rect 1235 1444 1236 1448
rect 1230 1443 1236 1444
rect 1278 1448 1284 1449
rect 1278 1444 1279 1448
rect 1283 1444 1284 1448
rect 1278 1443 1284 1444
rect 1334 1448 1340 1449
rect 1334 1444 1335 1448
rect 1339 1444 1340 1448
rect 1334 1443 1340 1444
rect 1390 1448 1396 1449
rect 1390 1444 1391 1448
rect 1395 1444 1396 1448
rect 1390 1443 1396 1444
rect 1454 1448 1460 1449
rect 1454 1444 1455 1448
rect 1459 1444 1460 1448
rect 1454 1443 1460 1444
rect 1518 1448 1524 1449
rect 1518 1444 1519 1448
rect 1523 1444 1524 1448
rect 1518 1443 1524 1444
rect 1582 1448 1588 1449
rect 1582 1444 1583 1448
rect 1587 1444 1588 1448
rect 1582 1443 1588 1444
rect 1646 1448 1652 1449
rect 1646 1444 1647 1448
rect 1651 1444 1652 1448
rect 1646 1443 1652 1444
rect 1718 1448 1724 1449
rect 1718 1444 1719 1448
rect 1723 1444 1724 1448
rect 1718 1443 1724 1444
rect 1806 1448 1812 1449
rect 1806 1444 1807 1448
rect 1811 1444 1812 1448
rect 1806 1443 1812 1444
rect 1894 1448 1900 1449
rect 1894 1444 1895 1448
rect 1899 1444 1900 1448
rect 1894 1443 1900 1444
rect 1990 1448 1996 1449
rect 1990 1444 1991 1448
rect 1995 1444 1996 1448
rect 1990 1443 1996 1444
rect 2070 1448 2076 1449
rect 2070 1444 2071 1448
rect 2075 1444 2076 1448
rect 2070 1443 2076 1444
rect 2120 1441 2122 1461
rect 1094 1439 1100 1440
rect 1134 1440 1140 1441
rect 1134 1436 1135 1440
rect 1139 1436 1140 1440
rect 1134 1435 1140 1436
rect 2118 1440 2124 1441
rect 2118 1436 2119 1440
rect 2123 1436 2124 1440
rect 2118 1435 2124 1436
rect 110 1427 116 1428
rect 110 1423 111 1427
rect 115 1423 116 1427
rect 1094 1427 1100 1428
rect 110 1422 116 1423
rect 518 1424 524 1425
rect 112 1415 114 1422
rect 518 1420 519 1424
rect 523 1420 524 1424
rect 518 1419 524 1420
rect 558 1424 564 1425
rect 558 1420 559 1424
rect 563 1420 564 1424
rect 558 1419 564 1420
rect 598 1424 604 1425
rect 598 1420 599 1424
rect 603 1420 604 1424
rect 598 1419 604 1420
rect 646 1424 652 1425
rect 646 1420 647 1424
rect 651 1420 652 1424
rect 646 1419 652 1420
rect 694 1424 700 1425
rect 694 1420 695 1424
rect 699 1420 700 1424
rect 694 1419 700 1420
rect 750 1424 756 1425
rect 750 1420 751 1424
rect 755 1420 756 1424
rect 750 1419 756 1420
rect 806 1424 812 1425
rect 806 1420 807 1424
rect 811 1420 812 1424
rect 806 1419 812 1420
rect 870 1424 876 1425
rect 870 1420 871 1424
rect 875 1420 876 1424
rect 870 1419 876 1420
rect 934 1424 940 1425
rect 934 1420 935 1424
rect 939 1420 940 1424
rect 1094 1423 1095 1427
rect 1099 1423 1100 1427
rect 1094 1422 1100 1423
rect 1134 1423 1140 1424
rect 934 1419 940 1420
rect 520 1415 522 1419
rect 560 1415 562 1419
rect 600 1415 602 1419
rect 648 1415 650 1419
rect 696 1415 698 1419
rect 752 1415 754 1419
rect 808 1415 810 1419
rect 872 1415 874 1419
rect 936 1415 938 1419
rect 1096 1415 1098 1422
rect 1134 1419 1135 1423
rect 1139 1419 1140 1423
rect 2118 1423 2124 1424
rect 1134 1418 1140 1419
rect 1230 1420 1236 1421
rect 111 1414 115 1415
rect 111 1409 115 1410
rect 431 1414 435 1415
rect 431 1409 435 1410
rect 471 1414 475 1415
rect 471 1409 475 1410
rect 519 1414 523 1415
rect 519 1409 523 1410
rect 559 1414 563 1415
rect 559 1409 563 1410
rect 575 1414 579 1415
rect 575 1409 579 1410
rect 599 1414 603 1415
rect 599 1409 603 1410
rect 631 1414 635 1415
rect 631 1409 635 1410
rect 647 1414 651 1415
rect 647 1409 651 1410
rect 695 1414 699 1415
rect 695 1409 699 1410
rect 751 1414 755 1415
rect 751 1409 755 1410
rect 759 1414 763 1415
rect 759 1409 763 1410
rect 807 1414 811 1415
rect 807 1409 811 1410
rect 823 1414 827 1415
rect 823 1409 827 1410
rect 871 1414 875 1415
rect 871 1409 875 1410
rect 895 1414 899 1415
rect 895 1409 899 1410
rect 935 1414 939 1415
rect 935 1409 939 1410
rect 967 1414 971 1415
rect 967 1409 971 1410
rect 1095 1414 1099 1415
rect 1136 1411 1138 1418
rect 1230 1416 1231 1420
rect 1235 1416 1236 1420
rect 1230 1415 1236 1416
rect 1278 1420 1284 1421
rect 1278 1416 1279 1420
rect 1283 1416 1284 1420
rect 1278 1415 1284 1416
rect 1334 1420 1340 1421
rect 1334 1416 1335 1420
rect 1339 1416 1340 1420
rect 1334 1415 1340 1416
rect 1390 1420 1396 1421
rect 1390 1416 1391 1420
rect 1395 1416 1396 1420
rect 1390 1415 1396 1416
rect 1454 1420 1460 1421
rect 1454 1416 1455 1420
rect 1459 1416 1460 1420
rect 1454 1415 1460 1416
rect 1518 1420 1524 1421
rect 1518 1416 1519 1420
rect 1523 1416 1524 1420
rect 1518 1415 1524 1416
rect 1582 1420 1588 1421
rect 1582 1416 1583 1420
rect 1587 1416 1588 1420
rect 1582 1415 1588 1416
rect 1646 1420 1652 1421
rect 1646 1416 1647 1420
rect 1651 1416 1652 1420
rect 1646 1415 1652 1416
rect 1718 1420 1724 1421
rect 1718 1416 1719 1420
rect 1723 1416 1724 1420
rect 1718 1415 1724 1416
rect 1806 1420 1812 1421
rect 1806 1416 1807 1420
rect 1811 1416 1812 1420
rect 1806 1415 1812 1416
rect 1894 1420 1900 1421
rect 1894 1416 1895 1420
rect 1899 1416 1900 1420
rect 1894 1415 1900 1416
rect 1990 1420 1996 1421
rect 1990 1416 1991 1420
rect 1995 1416 1996 1420
rect 1990 1415 1996 1416
rect 2070 1420 2076 1421
rect 2070 1416 2071 1420
rect 2075 1416 2076 1420
rect 2118 1419 2119 1423
rect 2123 1419 2124 1423
rect 2118 1418 2124 1419
rect 2070 1415 2076 1416
rect 1232 1411 1234 1415
rect 1280 1411 1282 1415
rect 1336 1411 1338 1415
rect 1392 1411 1394 1415
rect 1456 1411 1458 1415
rect 1520 1411 1522 1415
rect 1584 1411 1586 1415
rect 1648 1411 1650 1415
rect 1720 1411 1722 1415
rect 1808 1411 1810 1415
rect 1896 1411 1898 1415
rect 1992 1411 1994 1415
rect 2072 1411 2074 1415
rect 2120 1411 2122 1418
rect 1095 1409 1099 1410
rect 1135 1410 1139 1411
rect 112 1406 114 1409
rect 430 1408 436 1409
rect 110 1405 116 1406
rect 110 1401 111 1405
rect 115 1401 116 1405
rect 430 1404 431 1408
rect 435 1404 436 1408
rect 430 1403 436 1404
rect 470 1408 476 1409
rect 470 1404 471 1408
rect 475 1404 476 1408
rect 470 1403 476 1404
rect 518 1408 524 1409
rect 518 1404 519 1408
rect 523 1404 524 1408
rect 518 1403 524 1404
rect 574 1408 580 1409
rect 574 1404 575 1408
rect 579 1404 580 1408
rect 574 1403 580 1404
rect 630 1408 636 1409
rect 630 1404 631 1408
rect 635 1404 636 1408
rect 630 1403 636 1404
rect 694 1408 700 1409
rect 694 1404 695 1408
rect 699 1404 700 1408
rect 694 1403 700 1404
rect 758 1408 764 1409
rect 758 1404 759 1408
rect 763 1404 764 1408
rect 758 1403 764 1404
rect 822 1408 828 1409
rect 822 1404 823 1408
rect 827 1404 828 1408
rect 822 1403 828 1404
rect 894 1408 900 1409
rect 894 1404 895 1408
rect 899 1404 900 1408
rect 894 1403 900 1404
rect 966 1408 972 1409
rect 966 1404 967 1408
rect 971 1404 972 1408
rect 1096 1406 1098 1409
rect 966 1403 972 1404
rect 1094 1405 1100 1406
rect 1135 1405 1139 1406
rect 1159 1410 1163 1411
rect 1159 1405 1163 1406
rect 1199 1410 1203 1411
rect 1199 1405 1203 1406
rect 1231 1410 1235 1411
rect 1231 1405 1235 1406
rect 1263 1410 1267 1411
rect 1263 1405 1267 1406
rect 1279 1410 1283 1411
rect 1279 1405 1283 1406
rect 1335 1410 1339 1411
rect 1335 1405 1339 1406
rect 1351 1410 1355 1411
rect 1351 1405 1355 1406
rect 1391 1410 1395 1411
rect 1391 1405 1395 1406
rect 1447 1410 1451 1411
rect 1447 1405 1451 1406
rect 1455 1410 1459 1411
rect 1455 1405 1459 1406
rect 1519 1410 1523 1411
rect 1519 1405 1523 1406
rect 1543 1410 1547 1411
rect 1543 1405 1547 1406
rect 1583 1410 1587 1411
rect 1583 1405 1587 1406
rect 1631 1410 1635 1411
rect 1631 1405 1635 1406
rect 1647 1410 1651 1411
rect 1647 1405 1651 1406
rect 1719 1410 1723 1411
rect 1719 1405 1723 1406
rect 1799 1410 1803 1411
rect 1799 1405 1803 1406
rect 1807 1410 1811 1411
rect 1807 1405 1811 1406
rect 1871 1410 1875 1411
rect 1871 1405 1875 1406
rect 1895 1410 1899 1411
rect 1895 1405 1899 1406
rect 1943 1410 1947 1411
rect 1943 1405 1947 1406
rect 1991 1410 1995 1411
rect 1991 1405 1995 1406
rect 2015 1410 2019 1411
rect 2015 1405 2019 1406
rect 2071 1410 2075 1411
rect 2071 1405 2075 1406
rect 2119 1410 2123 1411
rect 2119 1405 2123 1406
rect 110 1400 116 1401
rect 1094 1401 1095 1405
rect 1099 1401 1100 1405
rect 1136 1402 1138 1405
rect 1158 1404 1164 1405
rect 1094 1400 1100 1401
rect 1134 1401 1140 1402
rect 1134 1397 1135 1401
rect 1139 1397 1140 1401
rect 1158 1400 1159 1404
rect 1163 1400 1164 1404
rect 1158 1399 1164 1400
rect 1198 1404 1204 1405
rect 1198 1400 1199 1404
rect 1203 1400 1204 1404
rect 1198 1399 1204 1400
rect 1262 1404 1268 1405
rect 1262 1400 1263 1404
rect 1267 1400 1268 1404
rect 1262 1399 1268 1400
rect 1350 1404 1356 1405
rect 1350 1400 1351 1404
rect 1355 1400 1356 1404
rect 1350 1399 1356 1400
rect 1446 1404 1452 1405
rect 1446 1400 1447 1404
rect 1451 1400 1452 1404
rect 1446 1399 1452 1400
rect 1542 1404 1548 1405
rect 1542 1400 1543 1404
rect 1547 1400 1548 1404
rect 1542 1399 1548 1400
rect 1630 1404 1636 1405
rect 1630 1400 1631 1404
rect 1635 1400 1636 1404
rect 1630 1399 1636 1400
rect 1718 1404 1724 1405
rect 1718 1400 1719 1404
rect 1723 1400 1724 1404
rect 1718 1399 1724 1400
rect 1798 1404 1804 1405
rect 1798 1400 1799 1404
rect 1803 1400 1804 1404
rect 1798 1399 1804 1400
rect 1870 1404 1876 1405
rect 1870 1400 1871 1404
rect 1875 1400 1876 1404
rect 1870 1399 1876 1400
rect 1942 1404 1948 1405
rect 1942 1400 1943 1404
rect 1947 1400 1948 1404
rect 1942 1399 1948 1400
rect 2014 1404 2020 1405
rect 2014 1400 2015 1404
rect 2019 1400 2020 1404
rect 2014 1399 2020 1400
rect 2070 1404 2076 1405
rect 2070 1400 2071 1404
rect 2075 1400 2076 1404
rect 2120 1402 2122 1405
rect 2070 1399 2076 1400
rect 2118 1401 2124 1402
rect 1134 1396 1140 1397
rect 2118 1397 2119 1401
rect 2123 1397 2124 1401
rect 2118 1396 2124 1397
rect 110 1388 116 1389
rect 110 1384 111 1388
rect 115 1384 116 1388
rect 110 1383 116 1384
rect 1094 1388 1100 1389
rect 1094 1384 1095 1388
rect 1099 1384 1100 1388
rect 1094 1383 1100 1384
rect 1134 1384 1140 1385
rect 112 1363 114 1383
rect 430 1380 436 1381
rect 430 1376 431 1380
rect 435 1376 436 1380
rect 430 1375 436 1376
rect 470 1380 476 1381
rect 470 1376 471 1380
rect 475 1376 476 1380
rect 470 1375 476 1376
rect 518 1380 524 1381
rect 518 1376 519 1380
rect 523 1376 524 1380
rect 518 1375 524 1376
rect 574 1380 580 1381
rect 574 1376 575 1380
rect 579 1376 580 1380
rect 574 1375 580 1376
rect 630 1380 636 1381
rect 630 1376 631 1380
rect 635 1376 636 1380
rect 630 1375 636 1376
rect 694 1380 700 1381
rect 694 1376 695 1380
rect 699 1376 700 1380
rect 694 1375 700 1376
rect 758 1380 764 1381
rect 758 1376 759 1380
rect 763 1376 764 1380
rect 758 1375 764 1376
rect 822 1380 828 1381
rect 822 1376 823 1380
rect 827 1376 828 1380
rect 822 1375 828 1376
rect 894 1380 900 1381
rect 894 1376 895 1380
rect 899 1376 900 1380
rect 894 1375 900 1376
rect 966 1380 972 1381
rect 966 1376 967 1380
rect 971 1376 972 1380
rect 966 1375 972 1376
rect 432 1363 434 1375
rect 472 1363 474 1375
rect 520 1363 522 1375
rect 576 1363 578 1375
rect 632 1363 634 1375
rect 696 1363 698 1375
rect 760 1363 762 1375
rect 824 1363 826 1375
rect 896 1363 898 1375
rect 968 1363 970 1375
rect 1096 1363 1098 1383
rect 1134 1380 1135 1384
rect 1139 1380 1140 1384
rect 1134 1379 1140 1380
rect 2118 1384 2124 1385
rect 2118 1380 2119 1384
rect 2123 1380 2124 1384
rect 2118 1379 2124 1380
rect 111 1362 115 1363
rect 111 1357 115 1358
rect 375 1362 379 1363
rect 375 1357 379 1358
rect 423 1362 427 1363
rect 423 1357 427 1358
rect 431 1362 435 1363
rect 431 1357 435 1358
rect 471 1362 475 1363
rect 471 1357 475 1358
rect 479 1362 483 1363
rect 479 1357 483 1358
rect 519 1362 523 1363
rect 519 1357 523 1358
rect 543 1362 547 1363
rect 543 1357 547 1358
rect 575 1362 579 1363
rect 575 1357 579 1358
rect 607 1362 611 1363
rect 607 1357 611 1358
rect 631 1362 635 1363
rect 631 1357 635 1358
rect 671 1362 675 1363
rect 671 1357 675 1358
rect 695 1362 699 1363
rect 695 1357 699 1358
rect 735 1362 739 1363
rect 735 1357 739 1358
rect 759 1362 763 1363
rect 759 1357 763 1358
rect 799 1362 803 1363
rect 799 1357 803 1358
rect 823 1362 827 1363
rect 823 1357 827 1358
rect 863 1362 867 1363
rect 863 1357 867 1358
rect 895 1362 899 1363
rect 895 1357 899 1358
rect 927 1362 931 1363
rect 927 1357 931 1358
rect 967 1362 971 1363
rect 967 1357 971 1358
rect 999 1362 1003 1363
rect 999 1357 1003 1358
rect 1047 1362 1051 1363
rect 1047 1357 1051 1358
rect 1095 1362 1099 1363
rect 1095 1357 1099 1358
rect 112 1337 114 1357
rect 376 1345 378 1357
rect 424 1345 426 1357
rect 480 1345 482 1357
rect 544 1345 546 1357
rect 608 1345 610 1357
rect 672 1345 674 1357
rect 736 1345 738 1357
rect 800 1345 802 1357
rect 864 1345 866 1357
rect 928 1345 930 1357
rect 1000 1345 1002 1357
rect 1048 1345 1050 1357
rect 374 1344 380 1345
rect 374 1340 375 1344
rect 379 1340 380 1344
rect 374 1339 380 1340
rect 422 1344 428 1345
rect 422 1340 423 1344
rect 427 1340 428 1344
rect 422 1339 428 1340
rect 478 1344 484 1345
rect 478 1340 479 1344
rect 483 1340 484 1344
rect 478 1339 484 1340
rect 542 1344 548 1345
rect 542 1340 543 1344
rect 547 1340 548 1344
rect 542 1339 548 1340
rect 606 1344 612 1345
rect 606 1340 607 1344
rect 611 1340 612 1344
rect 606 1339 612 1340
rect 670 1344 676 1345
rect 670 1340 671 1344
rect 675 1340 676 1344
rect 670 1339 676 1340
rect 734 1344 740 1345
rect 734 1340 735 1344
rect 739 1340 740 1344
rect 734 1339 740 1340
rect 798 1344 804 1345
rect 798 1340 799 1344
rect 803 1340 804 1344
rect 798 1339 804 1340
rect 862 1344 868 1345
rect 862 1340 863 1344
rect 867 1340 868 1344
rect 862 1339 868 1340
rect 926 1344 932 1345
rect 926 1340 927 1344
rect 931 1340 932 1344
rect 926 1339 932 1340
rect 998 1344 1004 1345
rect 998 1340 999 1344
rect 1003 1340 1004 1344
rect 998 1339 1004 1340
rect 1046 1344 1052 1345
rect 1046 1340 1047 1344
rect 1051 1340 1052 1344
rect 1046 1339 1052 1340
rect 1096 1337 1098 1357
rect 1136 1355 1138 1379
rect 1158 1376 1164 1377
rect 1158 1372 1159 1376
rect 1163 1372 1164 1376
rect 1158 1371 1164 1372
rect 1198 1376 1204 1377
rect 1198 1372 1199 1376
rect 1203 1372 1204 1376
rect 1198 1371 1204 1372
rect 1262 1376 1268 1377
rect 1262 1372 1263 1376
rect 1267 1372 1268 1376
rect 1262 1371 1268 1372
rect 1350 1376 1356 1377
rect 1350 1372 1351 1376
rect 1355 1372 1356 1376
rect 1350 1371 1356 1372
rect 1446 1376 1452 1377
rect 1446 1372 1447 1376
rect 1451 1372 1452 1376
rect 1446 1371 1452 1372
rect 1542 1376 1548 1377
rect 1542 1372 1543 1376
rect 1547 1372 1548 1376
rect 1542 1371 1548 1372
rect 1630 1376 1636 1377
rect 1630 1372 1631 1376
rect 1635 1372 1636 1376
rect 1630 1371 1636 1372
rect 1718 1376 1724 1377
rect 1718 1372 1719 1376
rect 1723 1372 1724 1376
rect 1718 1371 1724 1372
rect 1798 1376 1804 1377
rect 1798 1372 1799 1376
rect 1803 1372 1804 1376
rect 1798 1371 1804 1372
rect 1870 1376 1876 1377
rect 1870 1372 1871 1376
rect 1875 1372 1876 1376
rect 1870 1371 1876 1372
rect 1942 1376 1948 1377
rect 1942 1372 1943 1376
rect 1947 1372 1948 1376
rect 1942 1371 1948 1372
rect 2014 1376 2020 1377
rect 2014 1372 2015 1376
rect 2019 1372 2020 1376
rect 2014 1371 2020 1372
rect 2070 1376 2076 1377
rect 2070 1372 2071 1376
rect 2075 1372 2076 1376
rect 2070 1371 2076 1372
rect 1160 1355 1162 1371
rect 1200 1355 1202 1371
rect 1264 1355 1266 1371
rect 1352 1355 1354 1371
rect 1448 1355 1450 1371
rect 1544 1355 1546 1371
rect 1632 1355 1634 1371
rect 1720 1355 1722 1371
rect 1800 1355 1802 1371
rect 1872 1355 1874 1371
rect 1944 1355 1946 1371
rect 2016 1355 2018 1371
rect 2072 1355 2074 1371
rect 2120 1355 2122 1379
rect 1135 1354 1139 1355
rect 1135 1349 1139 1350
rect 1159 1354 1163 1355
rect 1159 1349 1163 1350
rect 1199 1354 1203 1355
rect 1199 1349 1203 1350
rect 1255 1354 1259 1355
rect 1255 1349 1259 1350
rect 1263 1354 1267 1355
rect 1263 1349 1267 1350
rect 1351 1354 1355 1355
rect 1351 1349 1355 1350
rect 1375 1354 1379 1355
rect 1375 1349 1379 1350
rect 1447 1354 1451 1355
rect 1447 1349 1451 1350
rect 1487 1354 1491 1355
rect 1487 1349 1491 1350
rect 1543 1354 1547 1355
rect 1543 1349 1547 1350
rect 1591 1354 1595 1355
rect 1591 1349 1595 1350
rect 1631 1354 1635 1355
rect 1631 1349 1635 1350
rect 1679 1354 1683 1355
rect 1679 1349 1683 1350
rect 1719 1354 1723 1355
rect 1719 1349 1723 1350
rect 1759 1354 1763 1355
rect 1759 1349 1763 1350
rect 1799 1354 1803 1355
rect 1799 1349 1803 1350
rect 1831 1354 1835 1355
rect 1831 1349 1835 1350
rect 1871 1354 1875 1355
rect 1871 1349 1875 1350
rect 1903 1354 1907 1355
rect 1903 1349 1907 1350
rect 1943 1354 1947 1355
rect 1943 1349 1947 1350
rect 1967 1354 1971 1355
rect 1967 1349 1971 1350
rect 2015 1354 2019 1355
rect 2015 1349 2019 1350
rect 2031 1354 2035 1355
rect 2031 1349 2035 1350
rect 2071 1354 2075 1355
rect 2071 1349 2075 1350
rect 2119 1354 2123 1355
rect 2119 1349 2123 1350
rect 110 1336 116 1337
rect 110 1332 111 1336
rect 115 1332 116 1336
rect 110 1331 116 1332
rect 1094 1336 1100 1337
rect 1094 1332 1095 1336
rect 1099 1332 1100 1336
rect 1094 1331 1100 1332
rect 1136 1329 1138 1349
rect 1160 1337 1162 1349
rect 1256 1337 1258 1349
rect 1376 1337 1378 1349
rect 1488 1337 1490 1349
rect 1592 1337 1594 1349
rect 1680 1337 1682 1349
rect 1760 1337 1762 1349
rect 1832 1337 1834 1349
rect 1904 1337 1906 1349
rect 1968 1337 1970 1349
rect 2032 1337 2034 1349
rect 2072 1337 2074 1349
rect 1158 1336 1164 1337
rect 1158 1332 1159 1336
rect 1163 1332 1164 1336
rect 1158 1331 1164 1332
rect 1254 1336 1260 1337
rect 1254 1332 1255 1336
rect 1259 1332 1260 1336
rect 1254 1331 1260 1332
rect 1374 1336 1380 1337
rect 1374 1332 1375 1336
rect 1379 1332 1380 1336
rect 1374 1331 1380 1332
rect 1486 1336 1492 1337
rect 1486 1332 1487 1336
rect 1491 1332 1492 1336
rect 1486 1331 1492 1332
rect 1590 1336 1596 1337
rect 1590 1332 1591 1336
rect 1595 1332 1596 1336
rect 1590 1331 1596 1332
rect 1678 1336 1684 1337
rect 1678 1332 1679 1336
rect 1683 1332 1684 1336
rect 1678 1331 1684 1332
rect 1758 1336 1764 1337
rect 1758 1332 1759 1336
rect 1763 1332 1764 1336
rect 1758 1331 1764 1332
rect 1830 1336 1836 1337
rect 1830 1332 1831 1336
rect 1835 1332 1836 1336
rect 1830 1331 1836 1332
rect 1902 1336 1908 1337
rect 1902 1332 1903 1336
rect 1907 1332 1908 1336
rect 1902 1331 1908 1332
rect 1966 1336 1972 1337
rect 1966 1332 1967 1336
rect 1971 1332 1972 1336
rect 1966 1331 1972 1332
rect 2030 1336 2036 1337
rect 2030 1332 2031 1336
rect 2035 1332 2036 1336
rect 2030 1331 2036 1332
rect 2070 1336 2076 1337
rect 2070 1332 2071 1336
rect 2075 1332 2076 1336
rect 2070 1331 2076 1332
rect 2120 1329 2122 1349
rect 1134 1328 1140 1329
rect 1134 1324 1135 1328
rect 1139 1324 1140 1328
rect 1134 1323 1140 1324
rect 2118 1328 2124 1329
rect 2118 1324 2119 1328
rect 2123 1324 2124 1328
rect 2118 1323 2124 1324
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 1094 1319 1100 1320
rect 110 1314 116 1315
rect 374 1316 380 1317
rect 112 1311 114 1314
rect 374 1312 375 1316
rect 379 1312 380 1316
rect 374 1311 380 1312
rect 422 1316 428 1317
rect 422 1312 423 1316
rect 427 1312 428 1316
rect 422 1311 428 1312
rect 478 1316 484 1317
rect 478 1312 479 1316
rect 483 1312 484 1316
rect 478 1311 484 1312
rect 542 1316 548 1317
rect 542 1312 543 1316
rect 547 1312 548 1316
rect 542 1311 548 1312
rect 606 1316 612 1317
rect 606 1312 607 1316
rect 611 1312 612 1316
rect 606 1311 612 1312
rect 670 1316 676 1317
rect 670 1312 671 1316
rect 675 1312 676 1316
rect 670 1311 676 1312
rect 734 1316 740 1317
rect 734 1312 735 1316
rect 739 1312 740 1316
rect 734 1311 740 1312
rect 798 1316 804 1317
rect 798 1312 799 1316
rect 803 1312 804 1316
rect 798 1311 804 1312
rect 862 1316 868 1317
rect 862 1312 863 1316
rect 867 1312 868 1316
rect 862 1311 868 1312
rect 926 1316 932 1317
rect 926 1312 927 1316
rect 931 1312 932 1316
rect 926 1311 932 1312
rect 998 1316 1004 1317
rect 998 1312 999 1316
rect 1003 1312 1004 1316
rect 998 1311 1004 1312
rect 1046 1316 1052 1317
rect 1046 1312 1047 1316
rect 1051 1312 1052 1316
rect 1094 1315 1095 1319
rect 1099 1315 1100 1319
rect 1094 1314 1100 1315
rect 1046 1311 1052 1312
rect 1096 1311 1098 1314
rect 1134 1311 1140 1312
rect 111 1310 115 1311
rect 111 1305 115 1306
rect 335 1310 339 1311
rect 335 1305 339 1306
rect 375 1310 379 1311
rect 375 1305 379 1306
rect 391 1310 395 1311
rect 391 1305 395 1306
rect 423 1310 427 1311
rect 423 1305 427 1306
rect 455 1310 459 1311
rect 455 1305 459 1306
rect 479 1310 483 1311
rect 479 1305 483 1306
rect 527 1310 531 1311
rect 527 1305 531 1306
rect 543 1310 547 1311
rect 543 1305 547 1306
rect 599 1310 603 1311
rect 599 1305 603 1306
rect 607 1310 611 1311
rect 607 1305 611 1306
rect 671 1310 675 1311
rect 671 1305 675 1306
rect 735 1310 739 1311
rect 735 1305 739 1306
rect 743 1310 747 1311
rect 743 1305 747 1306
rect 799 1310 803 1311
rect 799 1305 803 1306
rect 823 1310 827 1311
rect 823 1305 827 1306
rect 863 1310 867 1311
rect 863 1305 867 1306
rect 903 1310 907 1311
rect 903 1305 907 1306
rect 927 1310 931 1311
rect 927 1305 931 1306
rect 983 1310 987 1311
rect 983 1305 987 1306
rect 999 1310 1003 1311
rect 999 1305 1003 1306
rect 1047 1310 1051 1311
rect 1047 1305 1051 1306
rect 1095 1310 1099 1311
rect 1134 1307 1135 1311
rect 1139 1307 1140 1311
rect 2118 1311 2124 1312
rect 1134 1306 1140 1307
rect 1158 1308 1164 1309
rect 1095 1305 1099 1306
rect 112 1302 114 1305
rect 334 1304 340 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 334 1300 335 1304
rect 339 1300 340 1304
rect 334 1299 340 1300
rect 390 1304 396 1305
rect 390 1300 391 1304
rect 395 1300 396 1304
rect 390 1299 396 1300
rect 454 1304 460 1305
rect 454 1300 455 1304
rect 459 1300 460 1304
rect 454 1299 460 1300
rect 526 1304 532 1305
rect 526 1300 527 1304
rect 531 1300 532 1304
rect 526 1299 532 1300
rect 598 1304 604 1305
rect 598 1300 599 1304
rect 603 1300 604 1304
rect 598 1299 604 1300
rect 670 1304 676 1305
rect 670 1300 671 1304
rect 675 1300 676 1304
rect 670 1299 676 1300
rect 742 1304 748 1305
rect 742 1300 743 1304
rect 747 1300 748 1304
rect 742 1299 748 1300
rect 822 1304 828 1305
rect 822 1300 823 1304
rect 827 1300 828 1304
rect 822 1299 828 1300
rect 902 1304 908 1305
rect 902 1300 903 1304
rect 907 1300 908 1304
rect 902 1299 908 1300
rect 982 1304 988 1305
rect 982 1300 983 1304
rect 987 1300 988 1304
rect 982 1299 988 1300
rect 1046 1304 1052 1305
rect 1046 1300 1047 1304
rect 1051 1300 1052 1304
rect 1096 1302 1098 1305
rect 1046 1299 1052 1300
rect 1094 1301 1100 1302
rect 110 1296 116 1297
rect 1094 1297 1095 1301
rect 1099 1297 1100 1301
rect 1136 1299 1138 1306
rect 1158 1304 1159 1308
rect 1163 1304 1164 1308
rect 1158 1303 1164 1304
rect 1254 1308 1260 1309
rect 1254 1304 1255 1308
rect 1259 1304 1260 1308
rect 1254 1303 1260 1304
rect 1374 1308 1380 1309
rect 1374 1304 1375 1308
rect 1379 1304 1380 1308
rect 1374 1303 1380 1304
rect 1486 1308 1492 1309
rect 1486 1304 1487 1308
rect 1491 1304 1492 1308
rect 1486 1303 1492 1304
rect 1590 1308 1596 1309
rect 1590 1304 1591 1308
rect 1595 1304 1596 1308
rect 1590 1303 1596 1304
rect 1678 1308 1684 1309
rect 1678 1304 1679 1308
rect 1683 1304 1684 1308
rect 1678 1303 1684 1304
rect 1758 1308 1764 1309
rect 1758 1304 1759 1308
rect 1763 1304 1764 1308
rect 1758 1303 1764 1304
rect 1830 1308 1836 1309
rect 1830 1304 1831 1308
rect 1835 1304 1836 1308
rect 1830 1303 1836 1304
rect 1902 1308 1908 1309
rect 1902 1304 1903 1308
rect 1907 1304 1908 1308
rect 1902 1303 1908 1304
rect 1966 1308 1972 1309
rect 1966 1304 1967 1308
rect 1971 1304 1972 1308
rect 1966 1303 1972 1304
rect 2030 1308 2036 1309
rect 2030 1304 2031 1308
rect 2035 1304 2036 1308
rect 2030 1303 2036 1304
rect 2070 1308 2076 1309
rect 2070 1304 2071 1308
rect 2075 1304 2076 1308
rect 2118 1307 2119 1311
rect 2123 1307 2124 1311
rect 2118 1306 2124 1307
rect 2070 1303 2076 1304
rect 1160 1299 1162 1303
rect 1256 1299 1258 1303
rect 1376 1299 1378 1303
rect 1488 1299 1490 1303
rect 1592 1299 1594 1303
rect 1680 1299 1682 1303
rect 1760 1299 1762 1303
rect 1832 1299 1834 1303
rect 1904 1299 1906 1303
rect 1968 1299 1970 1303
rect 2032 1299 2034 1303
rect 2072 1299 2074 1303
rect 2120 1299 2122 1306
rect 1094 1296 1100 1297
rect 1135 1298 1139 1299
rect 1135 1293 1139 1294
rect 1159 1298 1163 1299
rect 1159 1293 1163 1294
rect 1199 1298 1203 1299
rect 1199 1293 1203 1294
rect 1247 1298 1251 1299
rect 1247 1293 1251 1294
rect 1255 1298 1259 1299
rect 1255 1293 1259 1294
rect 1319 1298 1323 1299
rect 1319 1293 1323 1294
rect 1375 1298 1379 1299
rect 1375 1293 1379 1294
rect 1399 1298 1403 1299
rect 1399 1293 1403 1294
rect 1479 1298 1483 1299
rect 1479 1293 1483 1294
rect 1487 1298 1491 1299
rect 1487 1293 1491 1294
rect 1559 1298 1563 1299
rect 1559 1293 1563 1294
rect 1591 1298 1595 1299
rect 1591 1293 1595 1294
rect 1639 1298 1643 1299
rect 1639 1293 1643 1294
rect 1679 1298 1683 1299
rect 1679 1293 1683 1294
rect 1719 1298 1723 1299
rect 1719 1293 1723 1294
rect 1759 1298 1763 1299
rect 1759 1293 1763 1294
rect 1799 1298 1803 1299
rect 1799 1293 1803 1294
rect 1831 1298 1835 1299
rect 1831 1293 1835 1294
rect 1879 1298 1883 1299
rect 1879 1293 1883 1294
rect 1903 1298 1907 1299
rect 1903 1293 1907 1294
rect 1967 1298 1971 1299
rect 1967 1293 1971 1294
rect 2031 1298 2035 1299
rect 2031 1293 2035 1294
rect 2055 1298 2059 1299
rect 2055 1293 2059 1294
rect 2071 1298 2075 1299
rect 2071 1293 2075 1294
rect 2119 1298 2123 1299
rect 2119 1293 2123 1294
rect 1136 1290 1138 1293
rect 1158 1292 1164 1293
rect 1134 1289 1140 1290
rect 1134 1285 1135 1289
rect 1139 1285 1140 1289
rect 1158 1288 1159 1292
rect 1163 1288 1164 1292
rect 1158 1287 1164 1288
rect 1198 1292 1204 1293
rect 1198 1288 1199 1292
rect 1203 1288 1204 1292
rect 1198 1287 1204 1288
rect 1246 1292 1252 1293
rect 1246 1288 1247 1292
rect 1251 1288 1252 1292
rect 1246 1287 1252 1288
rect 1318 1292 1324 1293
rect 1318 1288 1319 1292
rect 1323 1288 1324 1292
rect 1318 1287 1324 1288
rect 1398 1292 1404 1293
rect 1398 1288 1399 1292
rect 1403 1288 1404 1292
rect 1398 1287 1404 1288
rect 1478 1292 1484 1293
rect 1478 1288 1479 1292
rect 1483 1288 1484 1292
rect 1478 1287 1484 1288
rect 1558 1292 1564 1293
rect 1558 1288 1559 1292
rect 1563 1288 1564 1292
rect 1558 1287 1564 1288
rect 1638 1292 1644 1293
rect 1638 1288 1639 1292
rect 1643 1288 1644 1292
rect 1638 1287 1644 1288
rect 1718 1292 1724 1293
rect 1718 1288 1719 1292
rect 1723 1288 1724 1292
rect 1718 1287 1724 1288
rect 1798 1292 1804 1293
rect 1798 1288 1799 1292
rect 1803 1288 1804 1292
rect 1798 1287 1804 1288
rect 1878 1292 1884 1293
rect 1878 1288 1879 1292
rect 1883 1288 1884 1292
rect 1878 1287 1884 1288
rect 1966 1292 1972 1293
rect 1966 1288 1967 1292
rect 1971 1288 1972 1292
rect 1966 1287 1972 1288
rect 2054 1292 2060 1293
rect 2054 1288 2055 1292
rect 2059 1288 2060 1292
rect 2120 1290 2122 1293
rect 2054 1287 2060 1288
rect 2118 1289 2124 1290
rect 110 1284 116 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 110 1279 116 1280
rect 1094 1284 1100 1285
rect 1134 1284 1140 1285
rect 2118 1285 2119 1289
rect 2123 1285 2124 1289
rect 2118 1284 2124 1285
rect 1094 1280 1095 1284
rect 1099 1280 1100 1284
rect 1094 1279 1100 1280
rect 112 1255 114 1279
rect 334 1276 340 1277
rect 334 1272 335 1276
rect 339 1272 340 1276
rect 334 1271 340 1272
rect 390 1276 396 1277
rect 390 1272 391 1276
rect 395 1272 396 1276
rect 390 1271 396 1272
rect 454 1276 460 1277
rect 454 1272 455 1276
rect 459 1272 460 1276
rect 454 1271 460 1272
rect 526 1276 532 1277
rect 526 1272 527 1276
rect 531 1272 532 1276
rect 526 1271 532 1272
rect 598 1276 604 1277
rect 598 1272 599 1276
rect 603 1272 604 1276
rect 598 1271 604 1272
rect 670 1276 676 1277
rect 670 1272 671 1276
rect 675 1272 676 1276
rect 670 1271 676 1272
rect 742 1276 748 1277
rect 742 1272 743 1276
rect 747 1272 748 1276
rect 742 1271 748 1272
rect 822 1276 828 1277
rect 822 1272 823 1276
rect 827 1272 828 1276
rect 822 1271 828 1272
rect 902 1276 908 1277
rect 902 1272 903 1276
rect 907 1272 908 1276
rect 902 1271 908 1272
rect 982 1276 988 1277
rect 982 1272 983 1276
rect 987 1272 988 1276
rect 982 1271 988 1272
rect 1046 1276 1052 1277
rect 1046 1272 1047 1276
rect 1051 1272 1052 1276
rect 1046 1271 1052 1272
rect 336 1255 338 1271
rect 392 1255 394 1271
rect 456 1255 458 1271
rect 528 1255 530 1271
rect 600 1255 602 1271
rect 672 1255 674 1271
rect 744 1255 746 1271
rect 824 1255 826 1271
rect 904 1255 906 1271
rect 984 1255 986 1271
rect 1048 1255 1050 1271
rect 1096 1255 1098 1279
rect 1134 1272 1140 1273
rect 1134 1268 1135 1272
rect 1139 1268 1140 1272
rect 1134 1267 1140 1268
rect 2118 1272 2124 1273
rect 2118 1268 2119 1272
rect 2123 1268 2124 1272
rect 2118 1267 2124 1268
rect 111 1254 115 1255
rect 111 1249 115 1250
rect 263 1254 267 1255
rect 263 1249 267 1250
rect 311 1254 315 1255
rect 311 1249 315 1250
rect 335 1254 339 1255
rect 335 1249 339 1250
rect 359 1254 363 1255
rect 359 1249 363 1250
rect 391 1254 395 1255
rect 391 1249 395 1250
rect 415 1254 419 1255
rect 415 1249 419 1250
rect 455 1254 459 1255
rect 455 1249 459 1250
rect 479 1254 483 1255
rect 479 1249 483 1250
rect 527 1254 531 1255
rect 527 1249 531 1250
rect 543 1254 547 1255
rect 543 1249 547 1250
rect 599 1254 603 1255
rect 599 1249 603 1250
rect 607 1254 611 1255
rect 607 1249 611 1250
rect 671 1254 675 1255
rect 671 1249 675 1250
rect 735 1254 739 1255
rect 735 1249 739 1250
rect 743 1254 747 1255
rect 743 1249 747 1250
rect 799 1254 803 1255
rect 799 1249 803 1250
rect 823 1254 827 1255
rect 823 1249 827 1250
rect 863 1254 867 1255
rect 863 1249 867 1250
rect 903 1254 907 1255
rect 903 1249 907 1250
rect 927 1254 931 1255
rect 927 1249 931 1250
rect 983 1254 987 1255
rect 983 1249 987 1250
rect 1047 1254 1051 1255
rect 1047 1249 1051 1250
rect 1095 1254 1099 1255
rect 1095 1249 1099 1250
rect 112 1229 114 1249
rect 264 1237 266 1249
rect 312 1237 314 1249
rect 360 1237 362 1249
rect 416 1237 418 1249
rect 480 1237 482 1249
rect 544 1237 546 1249
rect 608 1237 610 1249
rect 672 1237 674 1249
rect 736 1237 738 1249
rect 800 1237 802 1249
rect 864 1237 866 1249
rect 928 1237 930 1249
rect 262 1236 268 1237
rect 262 1232 263 1236
rect 267 1232 268 1236
rect 262 1231 268 1232
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 358 1236 364 1237
rect 358 1232 359 1236
rect 363 1232 364 1236
rect 358 1231 364 1232
rect 414 1236 420 1237
rect 414 1232 415 1236
rect 419 1232 420 1236
rect 414 1231 420 1232
rect 478 1236 484 1237
rect 478 1232 479 1236
rect 483 1232 484 1236
rect 478 1231 484 1232
rect 542 1236 548 1237
rect 542 1232 543 1236
rect 547 1232 548 1236
rect 542 1231 548 1232
rect 606 1236 612 1237
rect 606 1232 607 1236
rect 611 1232 612 1236
rect 606 1231 612 1232
rect 670 1236 676 1237
rect 670 1232 671 1236
rect 675 1232 676 1236
rect 670 1231 676 1232
rect 734 1236 740 1237
rect 734 1232 735 1236
rect 739 1232 740 1236
rect 734 1231 740 1232
rect 798 1236 804 1237
rect 798 1232 799 1236
rect 803 1232 804 1236
rect 798 1231 804 1232
rect 862 1236 868 1237
rect 862 1232 863 1236
rect 867 1232 868 1236
rect 862 1231 868 1232
rect 926 1236 932 1237
rect 926 1232 927 1236
rect 931 1232 932 1236
rect 926 1231 932 1232
rect 1096 1229 1098 1249
rect 1136 1243 1138 1267
rect 1158 1264 1164 1265
rect 1158 1260 1159 1264
rect 1163 1260 1164 1264
rect 1158 1259 1164 1260
rect 1198 1264 1204 1265
rect 1198 1260 1199 1264
rect 1203 1260 1204 1264
rect 1198 1259 1204 1260
rect 1246 1264 1252 1265
rect 1246 1260 1247 1264
rect 1251 1260 1252 1264
rect 1246 1259 1252 1260
rect 1318 1264 1324 1265
rect 1318 1260 1319 1264
rect 1323 1260 1324 1264
rect 1318 1259 1324 1260
rect 1398 1264 1404 1265
rect 1398 1260 1399 1264
rect 1403 1260 1404 1264
rect 1398 1259 1404 1260
rect 1478 1264 1484 1265
rect 1478 1260 1479 1264
rect 1483 1260 1484 1264
rect 1478 1259 1484 1260
rect 1558 1264 1564 1265
rect 1558 1260 1559 1264
rect 1563 1260 1564 1264
rect 1558 1259 1564 1260
rect 1638 1264 1644 1265
rect 1638 1260 1639 1264
rect 1643 1260 1644 1264
rect 1638 1259 1644 1260
rect 1718 1264 1724 1265
rect 1718 1260 1719 1264
rect 1723 1260 1724 1264
rect 1718 1259 1724 1260
rect 1798 1264 1804 1265
rect 1798 1260 1799 1264
rect 1803 1260 1804 1264
rect 1798 1259 1804 1260
rect 1878 1264 1884 1265
rect 1878 1260 1879 1264
rect 1883 1260 1884 1264
rect 1878 1259 1884 1260
rect 1966 1264 1972 1265
rect 1966 1260 1967 1264
rect 1971 1260 1972 1264
rect 1966 1259 1972 1260
rect 2054 1264 2060 1265
rect 2054 1260 2055 1264
rect 2059 1260 2060 1264
rect 2054 1259 2060 1260
rect 1160 1243 1162 1259
rect 1200 1243 1202 1259
rect 1248 1243 1250 1259
rect 1320 1243 1322 1259
rect 1400 1243 1402 1259
rect 1480 1243 1482 1259
rect 1560 1243 1562 1259
rect 1640 1243 1642 1259
rect 1720 1243 1722 1259
rect 1800 1243 1802 1259
rect 1880 1243 1882 1259
rect 1968 1243 1970 1259
rect 2056 1243 2058 1259
rect 2120 1243 2122 1267
rect 1135 1242 1139 1243
rect 1135 1237 1139 1238
rect 1159 1242 1163 1243
rect 1159 1237 1163 1238
rect 1199 1242 1203 1243
rect 1199 1237 1203 1238
rect 1239 1242 1243 1243
rect 1239 1237 1243 1238
rect 1247 1242 1251 1243
rect 1247 1237 1251 1238
rect 1279 1242 1283 1243
rect 1279 1237 1283 1238
rect 1319 1242 1323 1243
rect 1319 1237 1323 1238
rect 1327 1242 1331 1243
rect 1327 1237 1331 1238
rect 1375 1242 1379 1243
rect 1375 1237 1379 1238
rect 1399 1242 1403 1243
rect 1399 1237 1403 1238
rect 1423 1242 1427 1243
rect 1423 1237 1427 1238
rect 1471 1242 1475 1243
rect 1471 1237 1475 1238
rect 1479 1242 1483 1243
rect 1479 1237 1483 1238
rect 1535 1242 1539 1243
rect 1535 1237 1539 1238
rect 1559 1242 1563 1243
rect 1559 1237 1563 1238
rect 1615 1242 1619 1243
rect 1615 1237 1619 1238
rect 1639 1242 1643 1243
rect 1639 1237 1643 1238
rect 1719 1242 1723 1243
rect 1719 1237 1723 1238
rect 1799 1242 1803 1243
rect 1799 1237 1803 1238
rect 1839 1242 1843 1243
rect 1839 1237 1843 1238
rect 1879 1242 1883 1243
rect 1879 1237 1883 1238
rect 1967 1242 1971 1243
rect 1967 1237 1971 1238
rect 2055 1242 2059 1243
rect 2055 1237 2059 1238
rect 2071 1242 2075 1243
rect 2071 1237 2075 1238
rect 2119 1242 2123 1243
rect 2119 1237 2123 1238
rect 110 1228 116 1229
rect 110 1224 111 1228
rect 115 1224 116 1228
rect 110 1223 116 1224
rect 1094 1228 1100 1229
rect 1094 1224 1095 1228
rect 1099 1224 1100 1228
rect 1094 1223 1100 1224
rect 1136 1217 1138 1237
rect 1160 1225 1162 1237
rect 1200 1225 1202 1237
rect 1240 1225 1242 1237
rect 1280 1225 1282 1237
rect 1328 1225 1330 1237
rect 1376 1225 1378 1237
rect 1424 1225 1426 1237
rect 1472 1225 1474 1237
rect 1536 1225 1538 1237
rect 1616 1225 1618 1237
rect 1720 1225 1722 1237
rect 1840 1225 1842 1237
rect 1968 1225 1970 1237
rect 2072 1225 2074 1237
rect 1158 1224 1164 1225
rect 1158 1220 1159 1224
rect 1163 1220 1164 1224
rect 1158 1219 1164 1220
rect 1198 1224 1204 1225
rect 1198 1220 1199 1224
rect 1203 1220 1204 1224
rect 1198 1219 1204 1220
rect 1238 1224 1244 1225
rect 1238 1220 1239 1224
rect 1243 1220 1244 1224
rect 1238 1219 1244 1220
rect 1278 1224 1284 1225
rect 1278 1220 1279 1224
rect 1283 1220 1284 1224
rect 1278 1219 1284 1220
rect 1326 1224 1332 1225
rect 1326 1220 1327 1224
rect 1331 1220 1332 1224
rect 1326 1219 1332 1220
rect 1374 1224 1380 1225
rect 1374 1220 1375 1224
rect 1379 1220 1380 1224
rect 1374 1219 1380 1220
rect 1422 1224 1428 1225
rect 1422 1220 1423 1224
rect 1427 1220 1428 1224
rect 1422 1219 1428 1220
rect 1470 1224 1476 1225
rect 1470 1220 1471 1224
rect 1475 1220 1476 1224
rect 1470 1219 1476 1220
rect 1534 1224 1540 1225
rect 1534 1220 1535 1224
rect 1539 1220 1540 1224
rect 1534 1219 1540 1220
rect 1614 1224 1620 1225
rect 1614 1220 1615 1224
rect 1619 1220 1620 1224
rect 1614 1219 1620 1220
rect 1718 1224 1724 1225
rect 1718 1220 1719 1224
rect 1723 1220 1724 1224
rect 1718 1219 1724 1220
rect 1838 1224 1844 1225
rect 1838 1220 1839 1224
rect 1843 1220 1844 1224
rect 1838 1219 1844 1220
rect 1966 1224 1972 1225
rect 1966 1220 1967 1224
rect 1971 1220 1972 1224
rect 1966 1219 1972 1220
rect 2070 1224 2076 1225
rect 2070 1220 2071 1224
rect 2075 1220 2076 1224
rect 2070 1219 2076 1220
rect 2120 1217 2122 1237
rect 1134 1216 1140 1217
rect 1134 1212 1135 1216
rect 1139 1212 1140 1216
rect 110 1211 116 1212
rect 110 1207 111 1211
rect 115 1207 116 1211
rect 1094 1211 1100 1212
rect 1134 1211 1140 1212
rect 2118 1216 2124 1217
rect 2118 1212 2119 1216
rect 2123 1212 2124 1216
rect 2118 1211 2124 1212
rect 110 1206 116 1207
rect 262 1208 268 1209
rect 112 1203 114 1206
rect 262 1204 263 1208
rect 267 1204 268 1208
rect 262 1203 268 1204
rect 310 1208 316 1209
rect 310 1204 311 1208
rect 315 1204 316 1208
rect 310 1203 316 1204
rect 358 1208 364 1209
rect 358 1204 359 1208
rect 363 1204 364 1208
rect 358 1203 364 1204
rect 414 1208 420 1209
rect 414 1204 415 1208
rect 419 1204 420 1208
rect 414 1203 420 1204
rect 478 1208 484 1209
rect 478 1204 479 1208
rect 483 1204 484 1208
rect 478 1203 484 1204
rect 542 1208 548 1209
rect 542 1204 543 1208
rect 547 1204 548 1208
rect 542 1203 548 1204
rect 606 1208 612 1209
rect 606 1204 607 1208
rect 611 1204 612 1208
rect 606 1203 612 1204
rect 670 1208 676 1209
rect 670 1204 671 1208
rect 675 1204 676 1208
rect 670 1203 676 1204
rect 734 1208 740 1209
rect 734 1204 735 1208
rect 739 1204 740 1208
rect 734 1203 740 1204
rect 798 1208 804 1209
rect 798 1204 799 1208
rect 803 1204 804 1208
rect 798 1203 804 1204
rect 862 1208 868 1209
rect 862 1204 863 1208
rect 867 1204 868 1208
rect 862 1203 868 1204
rect 926 1208 932 1209
rect 926 1204 927 1208
rect 931 1204 932 1208
rect 1094 1207 1095 1211
rect 1099 1207 1100 1211
rect 1094 1206 1100 1207
rect 926 1203 932 1204
rect 1096 1203 1098 1206
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 223 1202 227 1203
rect 223 1197 227 1198
rect 263 1202 267 1203
rect 263 1197 267 1198
rect 279 1202 283 1203
rect 279 1197 283 1198
rect 311 1202 315 1203
rect 311 1197 315 1198
rect 343 1202 347 1203
rect 343 1197 347 1198
rect 359 1202 363 1203
rect 359 1197 363 1198
rect 407 1202 411 1203
rect 407 1197 411 1198
rect 415 1202 419 1203
rect 415 1197 419 1198
rect 479 1202 483 1203
rect 479 1197 483 1198
rect 543 1202 547 1203
rect 543 1197 547 1198
rect 551 1202 555 1203
rect 551 1197 555 1198
rect 607 1202 611 1203
rect 607 1197 611 1198
rect 631 1202 635 1203
rect 631 1197 635 1198
rect 671 1202 675 1203
rect 671 1197 675 1198
rect 711 1202 715 1203
rect 711 1197 715 1198
rect 735 1202 739 1203
rect 735 1197 739 1198
rect 791 1202 795 1203
rect 791 1197 795 1198
rect 799 1202 803 1203
rect 799 1197 803 1198
rect 863 1202 867 1203
rect 863 1197 867 1198
rect 871 1202 875 1203
rect 871 1197 875 1198
rect 927 1202 931 1203
rect 927 1197 931 1198
rect 959 1202 963 1203
rect 959 1197 963 1198
rect 1095 1202 1099 1203
rect 1095 1197 1099 1198
rect 1134 1199 1140 1200
rect 112 1194 114 1197
rect 222 1196 228 1197
rect 110 1193 116 1194
rect 110 1189 111 1193
rect 115 1189 116 1193
rect 222 1192 223 1196
rect 227 1192 228 1196
rect 222 1191 228 1192
rect 278 1196 284 1197
rect 278 1192 279 1196
rect 283 1192 284 1196
rect 278 1191 284 1192
rect 342 1196 348 1197
rect 342 1192 343 1196
rect 347 1192 348 1196
rect 342 1191 348 1192
rect 406 1196 412 1197
rect 406 1192 407 1196
rect 411 1192 412 1196
rect 406 1191 412 1192
rect 478 1196 484 1197
rect 478 1192 479 1196
rect 483 1192 484 1196
rect 478 1191 484 1192
rect 550 1196 556 1197
rect 550 1192 551 1196
rect 555 1192 556 1196
rect 550 1191 556 1192
rect 630 1196 636 1197
rect 630 1192 631 1196
rect 635 1192 636 1196
rect 630 1191 636 1192
rect 710 1196 716 1197
rect 710 1192 711 1196
rect 715 1192 716 1196
rect 710 1191 716 1192
rect 790 1196 796 1197
rect 790 1192 791 1196
rect 795 1192 796 1196
rect 790 1191 796 1192
rect 870 1196 876 1197
rect 870 1192 871 1196
rect 875 1192 876 1196
rect 870 1191 876 1192
rect 958 1196 964 1197
rect 958 1192 959 1196
rect 963 1192 964 1196
rect 1096 1194 1098 1197
rect 1134 1195 1135 1199
rect 1139 1195 1140 1199
rect 2118 1199 2124 1200
rect 1134 1194 1140 1195
rect 1158 1196 1164 1197
rect 958 1191 964 1192
rect 1094 1193 1100 1194
rect 110 1188 116 1189
rect 1094 1189 1095 1193
rect 1099 1189 1100 1193
rect 1136 1191 1138 1194
rect 1158 1192 1159 1196
rect 1163 1192 1164 1196
rect 1158 1191 1164 1192
rect 1198 1196 1204 1197
rect 1198 1192 1199 1196
rect 1203 1192 1204 1196
rect 1198 1191 1204 1192
rect 1238 1196 1244 1197
rect 1238 1192 1239 1196
rect 1243 1192 1244 1196
rect 1238 1191 1244 1192
rect 1278 1196 1284 1197
rect 1278 1192 1279 1196
rect 1283 1192 1284 1196
rect 1278 1191 1284 1192
rect 1326 1196 1332 1197
rect 1326 1192 1327 1196
rect 1331 1192 1332 1196
rect 1326 1191 1332 1192
rect 1374 1196 1380 1197
rect 1374 1192 1375 1196
rect 1379 1192 1380 1196
rect 1374 1191 1380 1192
rect 1422 1196 1428 1197
rect 1422 1192 1423 1196
rect 1427 1192 1428 1196
rect 1422 1191 1428 1192
rect 1470 1196 1476 1197
rect 1470 1192 1471 1196
rect 1475 1192 1476 1196
rect 1470 1191 1476 1192
rect 1534 1196 1540 1197
rect 1534 1192 1535 1196
rect 1539 1192 1540 1196
rect 1534 1191 1540 1192
rect 1614 1196 1620 1197
rect 1614 1192 1615 1196
rect 1619 1192 1620 1196
rect 1614 1191 1620 1192
rect 1718 1196 1724 1197
rect 1718 1192 1719 1196
rect 1723 1192 1724 1196
rect 1718 1191 1724 1192
rect 1838 1196 1844 1197
rect 1838 1192 1839 1196
rect 1843 1192 1844 1196
rect 1838 1191 1844 1192
rect 1966 1196 1972 1197
rect 1966 1192 1967 1196
rect 1971 1192 1972 1196
rect 1966 1191 1972 1192
rect 2070 1196 2076 1197
rect 2070 1192 2071 1196
rect 2075 1192 2076 1196
rect 2118 1195 2119 1199
rect 2123 1195 2124 1199
rect 2118 1194 2124 1195
rect 2070 1191 2076 1192
rect 2120 1191 2122 1194
rect 1094 1188 1100 1189
rect 1135 1190 1139 1191
rect 1135 1185 1139 1186
rect 1159 1190 1163 1191
rect 1159 1185 1163 1186
rect 1199 1190 1203 1191
rect 1199 1185 1203 1186
rect 1239 1190 1243 1191
rect 1239 1185 1243 1186
rect 1279 1190 1283 1191
rect 1279 1185 1283 1186
rect 1287 1190 1291 1191
rect 1287 1185 1291 1186
rect 1327 1190 1331 1191
rect 1327 1185 1331 1186
rect 1367 1190 1371 1191
rect 1367 1185 1371 1186
rect 1375 1190 1379 1191
rect 1375 1185 1379 1186
rect 1415 1190 1419 1191
rect 1415 1185 1419 1186
rect 1423 1190 1427 1191
rect 1423 1185 1427 1186
rect 1471 1190 1475 1191
rect 1471 1185 1475 1186
rect 1527 1190 1531 1191
rect 1527 1185 1531 1186
rect 1535 1190 1539 1191
rect 1535 1185 1539 1186
rect 1583 1190 1587 1191
rect 1583 1185 1587 1186
rect 1615 1190 1619 1191
rect 1615 1185 1619 1186
rect 1639 1190 1643 1191
rect 1639 1185 1643 1186
rect 1703 1190 1707 1191
rect 1703 1185 1707 1186
rect 1719 1190 1723 1191
rect 1719 1185 1723 1186
rect 1767 1190 1771 1191
rect 1767 1185 1771 1186
rect 1839 1190 1843 1191
rect 1839 1185 1843 1186
rect 1919 1190 1923 1191
rect 1919 1185 1923 1186
rect 1967 1190 1971 1191
rect 1967 1185 1971 1186
rect 2007 1190 2011 1191
rect 2007 1185 2011 1186
rect 2071 1190 2075 1191
rect 2071 1185 2075 1186
rect 2119 1190 2123 1191
rect 2119 1185 2123 1186
rect 1136 1182 1138 1185
rect 1286 1184 1292 1185
rect 1134 1181 1140 1182
rect 1134 1177 1135 1181
rect 1139 1177 1140 1181
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1286 1179 1292 1180
rect 1326 1184 1332 1185
rect 1326 1180 1327 1184
rect 1331 1180 1332 1184
rect 1326 1179 1332 1180
rect 1366 1184 1372 1185
rect 1366 1180 1367 1184
rect 1371 1180 1372 1184
rect 1366 1179 1372 1180
rect 1414 1184 1420 1185
rect 1414 1180 1415 1184
rect 1419 1180 1420 1184
rect 1414 1179 1420 1180
rect 1470 1184 1476 1185
rect 1470 1180 1471 1184
rect 1475 1180 1476 1184
rect 1470 1179 1476 1180
rect 1526 1184 1532 1185
rect 1526 1180 1527 1184
rect 1531 1180 1532 1184
rect 1526 1179 1532 1180
rect 1582 1184 1588 1185
rect 1582 1180 1583 1184
rect 1587 1180 1588 1184
rect 1582 1179 1588 1180
rect 1638 1184 1644 1185
rect 1638 1180 1639 1184
rect 1643 1180 1644 1184
rect 1638 1179 1644 1180
rect 1702 1184 1708 1185
rect 1702 1180 1703 1184
rect 1707 1180 1708 1184
rect 1702 1179 1708 1180
rect 1766 1184 1772 1185
rect 1766 1180 1767 1184
rect 1771 1180 1772 1184
rect 1766 1179 1772 1180
rect 1838 1184 1844 1185
rect 1838 1180 1839 1184
rect 1843 1180 1844 1184
rect 1838 1179 1844 1180
rect 1918 1184 1924 1185
rect 1918 1180 1919 1184
rect 1923 1180 1924 1184
rect 1918 1179 1924 1180
rect 2006 1184 2012 1185
rect 2006 1180 2007 1184
rect 2011 1180 2012 1184
rect 2006 1179 2012 1180
rect 2070 1184 2076 1185
rect 2070 1180 2071 1184
rect 2075 1180 2076 1184
rect 2120 1182 2122 1185
rect 2070 1179 2076 1180
rect 2118 1181 2124 1182
rect 110 1176 116 1177
rect 110 1172 111 1176
rect 115 1172 116 1176
rect 110 1171 116 1172
rect 1094 1176 1100 1177
rect 1134 1176 1140 1177
rect 2118 1177 2119 1181
rect 2123 1177 2124 1181
rect 2118 1176 2124 1177
rect 1094 1172 1095 1176
rect 1099 1172 1100 1176
rect 1094 1171 1100 1172
rect 112 1151 114 1171
rect 222 1168 228 1169
rect 222 1164 223 1168
rect 227 1164 228 1168
rect 222 1163 228 1164
rect 278 1168 284 1169
rect 278 1164 279 1168
rect 283 1164 284 1168
rect 278 1163 284 1164
rect 342 1168 348 1169
rect 342 1164 343 1168
rect 347 1164 348 1168
rect 342 1163 348 1164
rect 406 1168 412 1169
rect 406 1164 407 1168
rect 411 1164 412 1168
rect 406 1163 412 1164
rect 478 1168 484 1169
rect 478 1164 479 1168
rect 483 1164 484 1168
rect 478 1163 484 1164
rect 550 1168 556 1169
rect 550 1164 551 1168
rect 555 1164 556 1168
rect 550 1163 556 1164
rect 630 1168 636 1169
rect 630 1164 631 1168
rect 635 1164 636 1168
rect 630 1163 636 1164
rect 710 1168 716 1169
rect 710 1164 711 1168
rect 715 1164 716 1168
rect 710 1163 716 1164
rect 790 1168 796 1169
rect 790 1164 791 1168
rect 795 1164 796 1168
rect 790 1163 796 1164
rect 870 1168 876 1169
rect 870 1164 871 1168
rect 875 1164 876 1168
rect 870 1163 876 1164
rect 958 1168 964 1169
rect 958 1164 959 1168
rect 963 1164 964 1168
rect 958 1163 964 1164
rect 224 1151 226 1163
rect 280 1151 282 1163
rect 344 1151 346 1163
rect 408 1151 410 1163
rect 480 1151 482 1163
rect 552 1151 554 1163
rect 632 1151 634 1163
rect 712 1151 714 1163
rect 792 1151 794 1163
rect 872 1151 874 1163
rect 960 1151 962 1163
rect 1096 1151 1098 1171
rect 1134 1164 1140 1165
rect 1134 1160 1135 1164
rect 1139 1160 1140 1164
rect 1134 1159 1140 1160
rect 2118 1164 2124 1165
rect 2118 1160 2119 1164
rect 2123 1160 2124 1164
rect 2118 1159 2124 1160
rect 111 1150 115 1151
rect 111 1145 115 1146
rect 159 1150 163 1151
rect 159 1145 163 1146
rect 199 1150 203 1151
rect 199 1145 203 1146
rect 223 1150 227 1151
rect 223 1145 227 1146
rect 247 1150 251 1151
rect 247 1145 251 1146
rect 279 1150 283 1151
rect 279 1145 283 1146
rect 303 1150 307 1151
rect 303 1145 307 1146
rect 343 1150 347 1151
rect 343 1145 347 1146
rect 367 1150 371 1151
rect 367 1145 371 1146
rect 407 1150 411 1151
rect 407 1145 411 1146
rect 439 1150 443 1151
rect 439 1145 443 1146
rect 479 1150 483 1151
rect 479 1145 483 1146
rect 511 1150 515 1151
rect 511 1145 515 1146
rect 551 1150 555 1151
rect 551 1145 555 1146
rect 591 1150 595 1151
rect 591 1145 595 1146
rect 631 1150 635 1151
rect 631 1145 635 1146
rect 679 1150 683 1151
rect 679 1145 683 1146
rect 711 1150 715 1151
rect 711 1145 715 1146
rect 775 1150 779 1151
rect 775 1145 779 1146
rect 791 1150 795 1151
rect 791 1145 795 1146
rect 871 1150 875 1151
rect 871 1145 875 1146
rect 879 1150 883 1151
rect 879 1145 883 1146
rect 959 1150 963 1151
rect 959 1145 963 1146
rect 991 1150 995 1151
rect 991 1145 995 1146
rect 1095 1150 1099 1151
rect 1095 1145 1099 1146
rect 112 1125 114 1145
rect 160 1133 162 1145
rect 200 1133 202 1145
rect 248 1133 250 1145
rect 304 1133 306 1145
rect 368 1133 370 1145
rect 440 1133 442 1145
rect 512 1133 514 1145
rect 592 1133 594 1145
rect 680 1133 682 1145
rect 776 1133 778 1145
rect 880 1133 882 1145
rect 992 1133 994 1145
rect 158 1132 164 1133
rect 158 1128 159 1132
rect 163 1128 164 1132
rect 158 1127 164 1128
rect 198 1132 204 1133
rect 198 1128 199 1132
rect 203 1128 204 1132
rect 198 1127 204 1128
rect 246 1132 252 1133
rect 246 1128 247 1132
rect 251 1128 252 1132
rect 246 1127 252 1128
rect 302 1132 308 1133
rect 302 1128 303 1132
rect 307 1128 308 1132
rect 302 1127 308 1128
rect 366 1132 372 1133
rect 366 1128 367 1132
rect 371 1128 372 1132
rect 366 1127 372 1128
rect 438 1132 444 1133
rect 438 1128 439 1132
rect 443 1128 444 1132
rect 438 1127 444 1128
rect 510 1132 516 1133
rect 510 1128 511 1132
rect 515 1128 516 1132
rect 510 1127 516 1128
rect 590 1132 596 1133
rect 590 1128 591 1132
rect 595 1128 596 1132
rect 590 1127 596 1128
rect 678 1132 684 1133
rect 678 1128 679 1132
rect 683 1128 684 1132
rect 678 1127 684 1128
rect 774 1132 780 1133
rect 774 1128 775 1132
rect 779 1128 780 1132
rect 774 1127 780 1128
rect 878 1132 884 1133
rect 878 1128 879 1132
rect 883 1128 884 1132
rect 878 1127 884 1128
rect 990 1132 996 1133
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 1096 1125 1098 1145
rect 1136 1131 1138 1159
rect 1286 1156 1292 1157
rect 1286 1152 1287 1156
rect 1291 1152 1292 1156
rect 1286 1151 1292 1152
rect 1326 1156 1332 1157
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1326 1151 1332 1152
rect 1366 1156 1372 1157
rect 1366 1152 1367 1156
rect 1371 1152 1372 1156
rect 1366 1151 1372 1152
rect 1414 1156 1420 1157
rect 1414 1152 1415 1156
rect 1419 1152 1420 1156
rect 1414 1151 1420 1152
rect 1470 1156 1476 1157
rect 1470 1152 1471 1156
rect 1475 1152 1476 1156
rect 1470 1151 1476 1152
rect 1526 1156 1532 1157
rect 1526 1152 1527 1156
rect 1531 1152 1532 1156
rect 1526 1151 1532 1152
rect 1582 1156 1588 1157
rect 1582 1152 1583 1156
rect 1587 1152 1588 1156
rect 1582 1151 1588 1152
rect 1638 1156 1644 1157
rect 1638 1152 1639 1156
rect 1643 1152 1644 1156
rect 1638 1151 1644 1152
rect 1702 1156 1708 1157
rect 1702 1152 1703 1156
rect 1707 1152 1708 1156
rect 1702 1151 1708 1152
rect 1766 1156 1772 1157
rect 1766 1152 1767 1156
rect 1771 1152 1772 1156
rect 1766 1151 1772 1152
rect 1838 1156 1844 1157
rect 1838 1152 1839 1156
rect 1843 1152 1844 1156
rect 1838 1151 1844 1152
rect 1918 1156 1924 1157
rect 1918 1152 1919 1156
rect 1923 1152 1924 1156
rect 1918 1151 1924 1152
rect 2006 1156 2012 1157
rect 2006 1152 2007 1156
rect 2011 1152 2012 1156
rect 2006 1151 2012 1152
rect 2070 1156 2076 1157
rect 2070 1152 2071 1156
rect 2075 1152 2076 1156
rect 2070 1151 2076 1152
rect 1288 1131 1290 1151
rect 1328 1131 1330 1151
rect 1368 1131 1370 1151
rect 1416 1131 1418 1151
rect 1472 1131 1474 1151
rect 1528 1131 1530 1151
rect 1584 1131 1586 1151
rect 1640 1131 1642 1151
rect 1704 1131 1706 1151
rect 1768 1131 1770 1151
rect 1840 1131 1842 1151
rect 1920 1131 1922 1151
rect 2008 1131 2010 1151
rect 2072 1131 2074 1151
rect 2120 1131 2122 1159
rect 1135 1130 1139 1131
rect 1135 1125 1139 1126
rect 1287 1130 1291 1131
rect 1287 1125 1291 1126
rect 1327 1130 1331 1131
rect 1327 1125 1331 1126
rect 1367 1130 1371 1131
rect 1367 1125 1371 1126
rect 1383 1130 1387 1131
rect 1383 1125 1387 1126
rect 1415 1130 1419 1131
rect 1415 1125 1419 1126
rect 1423 1130 1427 1131
rect 1423 1125 1427 1126
rect 1471 1130 1475 1131
rect 1471 1125 1475 1126
rect 1527 1130 1531 1131
rect 1527 1125 1531 1126
rect 1583 1130 1587 1131
rect 1583 1125 1587 1126
rect 1591 1130 1595 1131
rect 1591 1125 1595 1126
rect 1639 1130 1643 1131
rect 1639 1125 1643 1126
rect 1655 1130 1659 1131
rect 1655 1125 1659 1126
rect 1703 1130 1707 1131
rect 1703 1125 1707 1126
rect 1711 1130 1715 1131
rect 1711 1125 1715 1126
rect 1767 1130 1771 1131
rect 1767 1125 1771 1126
rect 1823 1130 1827 1131
rect 1823 1125 1827 1126
rect 1839 1130 1843 1131
rect 1839 1125 1843 1126
rect 1871 1130 1875 1131
rect 1871 1125 1875 1126
rect 1919 1130 1923 1131
rect 1919 1125 1923 1126
rect 1927 1130 1931 1131
rect 1927 1125 1931 1126
rect 1983 1130 1987 1131
rect 1983 1125 1987 1126
rect 2007 1130 2011 1131
rect 2007 1125 2011 1126
rect 2031 1130 2035 1131
rect 2031 1125 2035 1126
rect 2071 1130 2075 1131
rect 2071 1125 2075 1126
rect 2119 1130 2123 1131
rect 2119 1125 2123 1126
rect 110 1124 116 1125
rect 110 1120 111 1124
rect 115 1120 116 1124
rect 110 1119 116 1120
rect 1094 1124 1100 1125
rect 1094 1120 1095 1124
rect 1099 1120 1100 1124
rect 1094 1119 1100 1120
rect 110 1107 116 1108
rect 110 1103 111 1107
rect 115 1103 116 1107
rect 1094 1107 1100 1108
rect 110 1102 116 1103
rect 158 1104 164 1105
rect 112 1091 114 1102
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 198 1104 204 1105
rect 198 1100 199 1104
rect 203 1100 204 1104
rect 198 1099 204 1100
rect 246 1104 252 1105
rect 246 1100 247 1104
rect 251 1100 252 1104
rect 246 1099 252 1100
rect 302 1104 308 1105
rect 302 1100 303 1104
rect 307 1100 308 1104
rect 302 1099 308 1100
rect 366 1104 372 1105
rect 366 1100 367 1104
rect 371 1100 372 1104
rect 366 1099 372 1100
rect 438 1104 444 1105
rect 438 1100 439 1104
rect 443 1100 444 1104
rect 438 1099 444 1100
rect 510 1104 516 1105
rect 510 1100 511 1104
rect 515 1100 516 1104
rect 510 1099 516 1100
rect 590 1104 596 1105
rect 590 1100 591 1104
rect 595 1100 596 1104
rect 590 1099 596 1100
rect 678 1104 684 1105
rect 678 1100 679 1104
rect 683 1100 684 1104
rect 678 1099 684 1100
rect 774 1104 780 1105
rect 774 1100 775 1104
rect 779 1100 780 1104
rect 774 1099 780 1100
rect 878 1104 884 1105
rect 878 1100 879 1104
rect 883 1100 884 1104
rect 878 1099 884 1100
rect 990 1104 996 1105
rect 990 1100 991 1104
rect 995 1100 996 1104
rect 1094 1103 1095 1107
rect 1099 1103 1100 1107
rect 1136 1105 1138 1125
rect 1384 1113 1386 1125
rect 1424 1113 1426 1125
rect 1472 1113 1474 1125
rect 1528 1113 1530 1125
rect 1592 1113 1594 1125
rect 1656 1113 1658 1125
rect 1712 1113 1714 1125
rect 1768 1113 1770 1125
rect 1824 1113 1826 1125
rect 1872 1113 1874 1125
rect 1928 1113 1930 1125
rect 1984 1113 1986 1125
rect 2032 1113 2034 1125
rect 2072 1113 2074 1125
rect 1382 1112 1388 1113
rect 1382 1108 1383 1112
rect 1387 1108 1388 1112
rect 1382 1107 1388 1108
rect 1422 1112 1428 1113
rect 1422 1108 1423 1112
rect 1427 1108 1428 1112
rect 1422 1107 1428 1108
rect 1470 1112 1476 1113
rect 1470 1108 1471 1112
rect 1475 1108 1476 1112
rect 1470 1107 1476 1108
rect 1526 1112 1532 1113
rect 1526 1108 1527 1112
rect 1531 1108 1532 1112
rect 1526 1107 1532 1108
rect 1590 1112 1596 1113
rect 1590 1108 1591 1112
rect 1595 1108 1596 1112
rect 1590 1107 1596 1108
rect 1654 1112 1660 1113
rect 1654 1108 1655 1112
rect 1659 1108 1660 1112
rect 1654 1107 1660 1108
rect 1710 1112 1716 1113
rect 1710 1108 1711 1112
rect 1715 1108 1716 1112
rect 1710 1107 1716 1108
rect 1766 1112 1772 1113
rect 1766 1108 1767 1112
rect 1771 1108 1772 1112
rect 1766 1107 1772 1108
rect 1822 1112 1828 1113
rect 1822 1108 1823 1112
rect 1827 1108 1828 1112
rect 1822 1107 1828 1108
rect 1870 1112 1876 1113
rect 1870 1108 1871 1112
rect 1875 1108 1876 1112
rect 1870 1107 1876 1108
rect 1926 1112 1932 1113
rect 1926 1108 1927 1112
rect 1931 1108 1932 1112
rect 1926 1107 1932 1108
rect 1982 1112 1988 1113
rect 1982 1108 1983 1112
rect 1987 1108 1988 1112
rect 1982 1107 1988 1108
rect 2030 1112 2036 1113
rect 2030 1108 2031 1112
rect 2035 1108 2036 1112
rect 2030 1107 2036 1108
rect 2070 1112 2076 1113
rect 2070 1108 2071 1112
rect 2075 1108 2076 1112
rect 2070 1107 2076 1108
rect 2120 1105 2122 1125
rect 1094 1102 1100 1103
rect 1134 1104 1140 1105
rect 990 1099 996 1100
rect 160 1091 162 1099
rect 200 1091 202 1099
rect 248 1091 250 1099
rect 304 1091 306 1099
rect 368 1091 370 1099
rect 440 1091 442 1099
rect 512 1091 514 1099
rect 592 1091 594 1099
rect 680 1091 682 1099
rect 776 1091 778 1099
rect 880 1091 882 1099
rect 992 1091 994 1099
rect 1096 1091 1098 1102
rect 1134 1100 1135 1104
rect 1139 1100 1140 1104
rect 1134 1099 1140 1100
rect 2118 1104 2124 1105
rect 2118 1100 2119 1104
rect 2123 1100 2124 1104
rect 2118 1099 2124 1100
rect 111 1090 115 1091
rect 111 1085 115 1086
rect 159 1090 163 1091
rect 159 1085 163 1086
rect 199 1090 203 1091
rect 199 1085 203 1086
rect 247 1090 251 1091
rect 247 1085 251 1086
rect 303 1090 307 1091
rect 303 1085 307 1086
rect 367 1090 371 1091
rect 367 1085 371 1086
rect 431 1090 435 1091
rect 431 1085 435 1086
rect 439 1090 443 1091
rect 439 1085 443 1086
rect 503 1090 507 1091
rect 503 1085 507 1086
rect 511 1090 515 1091
rect 511 1085 515 1086
rect 575 1090 579 1091
rect 575 1085 579 1086
rect 591 1090 595 1091
rect 591 1085 595 1086
rect 647 1090 651 1091
rect 647 1085 651 1086
rect 679 1090 683 1091
rect 679 1085 683 1086
rect 719 1090 723 1091
rect 719 1085 723 1086
rect 775 1090 779 1091
rect 775 1085 779 1086
rect 783 1090 787 1091
rect 783 1085 787 1086
rect 839 1090 843 1091
rect 839 1085 843 1086
rect 879 1090 883 1091
rect 879 1085 883 1086
rect 895 1090 899 1091
rect 895 1085 899 1086
rect 951 1090 955 1091
rect 951 1085 955 1086
rect 991 1090 995 1091
rect 991 1085 995 1086
rect 1007 1090 1011 1091
rect 1007 1085 1011 1086
rect 1047 1090 1051 1091
rect 1047 1085 1051 1086
rect 1095 1090 1099 1091
rect 1095 1085 1099 1086
rect 1134 1087 1140 1088
rect 112 1082 114 1085
rect 198 1084 204 1085
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 198 1080 199 1084
rect 203 1080 204 1084
rect 198 1079 204 1080
rect 246 1084 252 1085
rect 246 1080 247 1084
rect 251 1080 252 1084
rect 246 1079 252 1080
rect 302 1084 308 1085
rect 302 1080 303 1084
rect 307 1080 308 1084
rect 302 1079 308 1080
rect 366 1084 372 1085
rect 366 1080 367 1084
rect 371 1080 372 1084
rect 366 1079 372 1080
rect 430 1084 436 1085
rect 430 1080 431 1084
rect 435 1080 436 1084
rect 430 1079 436 1080
rect 502 1084 508 1085
rect 502 1080 503 1084
rect 507 1080 508 1084
rect 502 1079 508 1080
rect 574 1084 580 1085
rect 574 1080 575 1084
rect 579 1080 580 1084
rect 574 1079 580 1080
rect 646 1084 652 1085
rect 646 1080 647 1084
rect 651 1080 652 1084
rect 646 1079 652 1080
rect 718 1084 724 1085
rect 718 1080 719 1084
rect 723 1080 724 1084
rect 718 1079 724 1080
rect 782 1084 788 1085
rect 782 1080 783 1084
rect 787 1080 788 1084
rect 782 1079 788 1080
rect 838 1084 844 1085
rect 838 1080 839 1084
rect 843 1080 844 1084
rect 838 1079 844 1080
rect 894 1084 900 1085
rect 894 1080 895 1084
rect 899 1080 900 1084
rect 894 1079 900 1080
rect 950 1084 956 1085
rect 950 1080 951 1084
rect 955 1080 956 1084
rect 950 1079 956 1080
rect 1006 1084 1012 1085
rect 1006 1080 1007 1084
rect 1011 1080 1012 1084
rect 1006 1079 1012 1080
rect 1046 1084 1052 1085
rect 1046 1080 1047 1084
rect 1051 1080 1052 1084
rect 1096 1082 1098 1085
rect 1134 1083 1135 1087
rect 1139 1083 1140 1087
rect 2118 1087 2124 1088
rect 1134 1082 1140 1083
rect 1382 1084 1388 1085
rect 1046 1079 1052 1080
rect 1094 1081 1100 1082
rect 110 1076 116 1077
rect 1094 1077 1095 1081
rect 1099 1077 1100 1081
rect 1136 1079 1138 1082
rect 1382 1080 1383 1084
rect 1387 1080 1388 1084
rect 1382 1079 1388 1080
rect 1422 1084 1428 1085
rect 1422 1080 1423 1084
rect 1427 1080 1428 1084
rect 1422 1079 1428 1080
rect 1470 1084 1476 1085
rect 1470 1080 1471 1084
rect 1475 1080 1476 1084
rect 1470 1079 1476 1080
rect 1526 1084 1532 1085
rect 1526 1080 1527 1084
rect 1531 1080 1532 1084
rect 1526 1079 1532 1080
rect 1590 1084 1596 1085
rect 1590 1080 1591 1084
rect 1595 1080 1596 1084
rect 1590 1079 1596 1080
rect 1654 1084 1660 1085
rect 1654 1080 1655 1084
rect 1659 1080 1660 1084
rect 1654 1079 1660 1080
rect 1710 1084 1716 1085
rect 1710 1080 1711 1084
rect 1715 1080 1716 1084
rect 1710 1079 1716 1080
rect 1766 1084 1772 1085
rect 1766 1080 1767 1084
rect 1771 1080 1772 1084
rect 1766 1079 1772 1080
rect 1822 1084 1828 1085
rect 1822 1080 1823 1084
rect 1827 1080 1828 1084
rect 1822 1079 1828 1080
rect 1870 1084 1876 1085
rect 1870 1080 1871 1084
rect 1875 1080 1876 1084
rect 1870 1079 1876 1080
rect 1926 1084 1932 1085
rect 1926 1080 1927 1084
rect 1931 1080 1932 1084
rect 1926 1079 1932 1080
rect 1982 1084 1988 1085
rect 1982 1080 1983 1084
rect 1987 1080 1988 1084
rect 1982 1079 1988 1080
rect 2030 1084 2036 1085
rect 2030 1080 2031 1084
rect 2035 1080 2036 1084
rect 2030 1079 2036 1080
rect 2070 1084 2076 1085
rect 2070 1080 2071 1084
rect 2075 1080 2076 1084
rect 2118 1083 2119 1087
rect 2123 1083 2124 1087
rect 2118 1082 2124 1083
rect 2070 1079 2076 1080
rect 2120 1079 2122 1082
rect 1094 1076 1100 1077
rect 1135 1078 1139 1079
rect 1135 1073 1139 1074
rect 1159 1078 1163 1079
rect 1159 1073 1163 1074
rect 1247 1078 1251 1079
rect 1247 1073 1251 1074
rect 1359 1078 1363 1079
rect 1359 1073 1363 1074
rect 1383 1078 1387 1079
rect 1383 1073 1387 1074
rect 1423 1078 1427 1079
rect 1423 1073 1427 1074
rect 1471 1078 1475 1079
rect 1471 1073 1475 1074
rect 1527 1078 1531 1079
rect 1527 1073 1531 1074
rect 1575 1078 1579 1079
rect 1575 1073 1579 1074
rect 1591 1078 1595 1079
rect 1591 1073 1595 1074
rect 1655 1078 1659 1079
rect 1655 1073 1659 1074
rect 1671 1078 1675 1079
rect 1671 1073 1675 1074
rect 1711 1078 1715 1079
rect 1711 1073 1715 1074
rect 1759 1078 1763 1079
rect 1759 1073 1763 1074
rect 1767 1078 1771 1079
rect 1767 1073 1771 1074
rect 1823 1078 1827 1079
rect 1823 1073 1827 1074
rect 1847 1078 1851 1079
rect 1847 1073 1851 1074
rect 1871 1078 1875 1079
rect 1871 1073 1875 1074
rect 1927 1078 1931 1079
rect 1927 1073 1931 1074
rect 1983 1078 1987 1079
rect 1983 1073 1987 1074
rect 2007 1078 2011 1079
rect 2007 1073 2011 1074
rect 2031 1078 2035 1079
rect 2031 1073 2035 1074
rect 2071 1078 2075 1079
rect 2071 1073 2075 1074
rect 2119 1078 2123 1079
rect 2119 1073 2123 1074
rect 1136 1070 1138 1073
rect 1158 1072 1164 1073
rect 1134 1069 1140 1070
rect 1134 1065 1135 1069
rect 1139 1065 1140 1069
rect 1158 1068 1159 1072
rect 1163 1068 1164 1072
rect 1158 1067 1164 1068
rect 1246 1072 1252 1073
rect 1246 1068 1247 1072
rect 1251 1068 1252 1072
rect 1246 1067 1252 1068
rect 1358 1072 1364 1073
rect 1358 1068 1359 1072
rect 1363 1068 1364 1072
rect 1358 1067 1364 1068
rect 1470 1072 1476 1073
rect 1470 1068 1471 1072
rect 1475 1068 1476 1072
rect 1470 1067 1476 1068
rect 1574 1072 1580 1073
rect 1574 1068 1575 1072
rect 1579 1068 1580 1072
rect 1574 1067 1580 1068
rect 1670 1072 1676 1073
rect 1670 1068 1671 1072
rect 1675 1068 1676 1072
rect 1670 1067 1676 1068
rect 1758 1072 1764 1073
rect 1758 1068 1759 1072
rect 1763 1068 1764 1072
rect 1758 1067 1764 1068
rect 1846 1072 1852 1073
rect 1846 1068 1847 1072
rect 1851 1068 1852 1072
rect 1846 1067 1852 1068
rect 1926 1072 1932 1073
rect 1926 1068 1927 1072
rect 1931 1068 1932 1072
rect 1926 1067 1932 1068
rect 2006 1072 2012 1073
rect 2006 1068 2007 1072
rect 2011 1068 2012 1072
rect 2006 1067 2012 1068
rect 2070 1072 2076 1073
rect 2070 1068 2071 1072
rect 2075 1068 2076 1072
rect 2120 1070 2122 1073
rect 2070 1067 2076 1068
rect 2118 1069 2124 1070
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 110 1059 116 1060
rect 1094 1064 1100 1065
rect 1134 1064 1140 1065
rect 2118 1065 2119 1069
rect 2123 1065 2124 1069
rect 2118 1064 2124 1065
rect 1094 1060 1095 1064
rect 1099 1060 1100 1064
rect 1094 1059 1100 1060
rect 112 1035 114 1059
rect 198 1056 204 1057
rect 198 1052 199 1056
rect 203 1052 204 1056
rect 198 1051 204 1052
rect 246 1056 252 1057
rect 246 1052 247 1056
rect 251 1052 252 1056
rect 246 1051 252 1052
rect 302 1056 308 1057
rect 302 1052 303 1056
rect 307 1052 308 1056
rect 302 1051 308 1052
rect 366 1056 372 1057
rect 366 1052 367 1056
rect 371 1052 372 1056
rect 366 1051 372 1052
rect 430 1056 436 1057
rect 430 1052 431 1056
rect 435 1052 436 1056
rect 430 1051 436 1052
rect 502 1056 508 1057
rect 502 1052 503 1056
rect 507 1052 508 1056
rect 502 1051 508 1052
rect 574 1056 580 1057
rect 574 1052 575 1056
rect 579 1052 580 1056
rect 574 1051 580 1052
rect 646 1056 652 1057
rect 646 1052 647 1056
rect 651 1052 652 1056
rect 646 1051 652 1052
rect 718 1056 724 1057
rect 718 1052 719 1056
rect 723 1052 724 1056
rect 718 1051 724 1052
rect 782 1056 788 1057
rect 782 1052 783 1056
rect 787 1052 788 1056
rect 782 1051 788 1052
rect 838 1056 844 1057
rect 838 1052 839 1056
rect 843 1052 844 1056
rect 838 1051 844 1052
rect 894 1056 900 1057
rect 894 1052 895 1056
rect 899 1052 900 1056
rect 894 1051 900 1052
rect 950 1056 956 1057
rect 950 1052 951 1056
rect 955 1052 956 1056
rect 950 1051 956 1052
rect 1006 1056 1012 1057
rect 1006 1052 1007 1056
rect 1011 1052 1012 1056
rect 1006 1051 1012 1052
rect 1046 1056 1052 1057
rect 1046 1052 1047 1056
rect 1051 1052 1052 1056
rect 1046 1051 1052 1052
rect 200 1035 202 1051
rect 248 1035 250 1051
rect 304 1035 306 1051
rect 368 1035 370 1051
rect 432 1035 434 1051
rect 504 1035 506 1051
rect 576 1035 578 1051
rect 648 1035 650 1051
rect 720 1035 722 1051
rect 784 1035 786 1051
rect 840 1035 842 1051
rect 896 1035 898 1051
rect 952 1035 954 1051
rect 1008 1035 1010 1051
rect 1048 1035 1050 1051
rect 1096 1035 1098 1059
rect 1134 1052 1140 1053
rect 1134 1048 1135 1052
rect 1139 1048 1140 1052
rect 1134 1047 1140 1048
rect 2118 1052 2124 1053
rect 2118 1048 2119 1052
rect 2123 1048 2124 1052
rect 2118 1047 2124 1048
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 199 1034 203 1035
rect 199 1029 203 1030
rect 223 1034 227 1035
rect 223 1029 227 1030
rect 247 1034 251 1035
rect 247 1029 251 1030
rect 271 1034 275 1035
rect 271 1029 275 1030
rect 303 1034 307 1035
rect 303 1029 307 1030
rect 335 1034 339 1035
rect 335 1029 339 1030
rect 367 1034 371 1035
rect 367 1029 371 1030
rect 407 1034 411 1035
rect 407 1029 411 1030
rect 431 1034 435 1035
rect 431 1029 435 1030
rect 479 1034 483 1035
rect 479 1029 483 1030
rect 503 1034 507 1035
rect 503 1029 507 1030
rect 559 1034 563 1035
rect 559 1029 563 1030
rect 575 1034 579 1035
rect 575 1029 579 1030
rect 631 1034 635 1035
rect 631 1029 635 1030
rect 647 1034 651 1035
rect 647 1029 651 1030
rect 703 1034 707 1035
rect 703 1029 707 1030
rect 719 1034 723 1035
rect 719 1029 723 1030
rect 775 1034 779 1035
rect 775 1029 779 1030
rect 783 1034 787 1035
rect 783 1029 787 1030
rect 839 1034 843 1035
rect 839 1029 843 1030
rect 895 1034 899 1035
rect 895 1029 899 1030
rect 903 1034 907 1035
rect 903 1029 907 1030
rect 951 1034 955 1035
rect 951 1029 955 1030
rect 967 1034 971 1035
rect 967 1029 971 1030
rect 1007 1034 1011 1035
rect 1007 1029 1011 1030
rect 1039 1034 1043 1035
rect 1039 1029 1043 1030
rect 1047 1034 1051 1035
rect 1047 1029 1051 1030
rect 1095 1034 1099 1035
rect 1095 1029 1099 1030
rect 112 1009 114 1029
rect 224 1017 226 1029
rect 272 1017 274 1029
rect 336 1017 338 1029
rect 408 1017 410 1029
rect 480 1017 482 1029
rect 560 1017 562 1029
rect 632 1017 634 1029
rect 704 1017 706 1029
rect 776 1017 778 1029
rect 840 1017 842 1029
rect 904 1017 906 1029
rect 968 1017 970 1029
rect 1040 1017 1042 1029
rect 222 1016 228 1017
rect 222 1012 223 1016
rect 227 1012 228 1016
rect 222 1011 228 1012
rect 270 1016 276 1017
rect 270 1012 271 1016
rect 275 1012 276 1016
rect 270 1011 276 1012
rect 334 1016 340 1017
rect 334 1012 335 1016
rect 339 1012 340 1016
rect 334 1011 340 1012
rect 406 1016 412 1017
rect 406 1012 407 1016
rect 411 1012 412 1016
rect 406 1011 412 1012
rect 478 1016 484 1017
rect 478 1012 479 1016
rect 483 1012 484 1016
rect 478 1011 484 1012
rect 558 1016 564 1017
rect 558 1012 559 1016
rect 563 1012 564 1016
rect 558 1011 564 1012
rect 630 1016 636 1017
rect 630 1012 631 1016
rect 635 1012 636 1016
rect 630 1011 636 1012
rect 702 1016 708 1017
rect 702 1012 703 1016
rect 707 1012 708 1016
rect 702 1011 708 1012
rect 774 1016 780 1017
rect 774 1012 775 1016
rect 779 1012 780 1016
rect 774 1011 780 1012
rect 838 1016 844 1017
rect 838 1012 839 1016
rect 843 1012 844 1016
rect 838 1011 844 1012
rect 902 1016 908 1017
rect 902 1012 903 1016
rect 907 1012 908 1016
rect 902 1011 908 1012
rect 966 1016 972 1017
rect 966 1012 967 1016
rect 971 1012 972 1016
rect 966 1011 972 1012
rect 1038 1016 1044 1017
rect 1038 1012 1039 1016
rect 1043 1012 1044 1016
rect 1038 1011 1044 1012
rect 1096 1009 1098 1029
rect 1136 1027 1138 1047
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1246 1044 1252 1045
rect 1246 1040 1247 1044
rect 1251 1040 1252 1044
rect 1246 1039 1252 1040
rect 1358 1044 1364 1045
rect 1358 1040 1359 1044
rect 1363 1040 1364 1044
rect 1358 1039 1364 1040
rect 1470 1044 1476 1045
rect 1470 1040 1471 1044
rect 1475 1040 1476 1044
rect 1470 1039 1476 1040
rect 1574 1044 1580 1045
rect 1574 1040 1575 1044
rect 1579 1040 1580 1044
rect 1574 1039 1580 1040
rect 1670 1044 1676 1045
rect 1670 1040 1671 1044
rect 1675 1040 1676 1044
rect 1670 1039 1676 1040
rect 1758 1044 1764 1045
rect 1758 1040 1759 1044
rect 1763 1040 1764 1044
rect 1758 1039 1764 1040
rect 1846 1044 1852 1045
rect 1846 1040 1847 1044
rect 1851 1040 1852 1044
rect 1846 1039 1852 1040
rect 1926 1044 1932 1045
rect 1926 1040 1927 1044
rect 1931 1040 1932 1044
rect 1926 1039 1932 1040
rect 2006 1044 2012 1045
rect 2006 1040 2007 1044
rect 2011 1040 2012 1044
rect 2006 1039 2012 1040
rect 2070 1044 2076 1045
rect 2070 1040 2071 1044
rect 2075 1040 2076 1044
rect 2070 1039 2076 1040
rect 1160 1027 1162 1039
rect 1248 1027 1250 1039
rect 1360 1027 1362 1039
rect 1472 1027 1474 1039
rect 1576 1027 1578 1039
rect 1672 1027 1674 1039
rect 1760 1027 1762 1039
rect 1848 1027 1850 1039
rect 1928 1027 1930 1039
rect 2008 1027 2010 1039
rect 2072 1027 2074 1039
rect 2120 1027 2122 1047
rect 1135 1026 1139 1027
rect 1135 1021 1139 1022
rect 1159 1026 1163 1027
rect 1159 1021 1163 1022
rect 1231 1026 1235 1027
rect 1231 1021 1235 1022
rect 1247 1026 1251 1027
rect 1247 1021 1251 1022
rect 1303 1026 1307 1027
rect 1303 1021 1307 1022
rect 1359 1026 1363 1027
rect 1359 1021 1363 1022
rect 1383 1026 1387 1027
rect 1383 1021 1387 1022
rect 1463 1026 1467 1027
rect 1463 1021 1467 1022
rect 1471 1026 1475 1027
rect 1471 1021 1475 1022
rect 1543 1026 1547 1027
rect 1543 1021 1547 1022
rect 1575 1026 1579 1027
rect 1575 1021 1579 1022
rect 1623 1026 1627 1027
rect 1623 1021 1627 1022
rect 1671 1026 1675 1027
rect 1671 1021 1675 1022
rect 1695 1026 1699 1027
rect 1695 1021 1699 1022
rect 1759 1026 1763 1027
rect 1759 1021 1763 1022
rect 1823 1026 1827 1027
rect 1823 1021 1827 1022
rect 1847 1026 1851 1027
rect 1847 1021 1851 1022
rect 1887 1026 1891 1027
rect 1887 1021 1891 1022
rect 1927 1026 1931 1027
rect 1927 1021 1931 1022
rect 1951 1026 1955 1027
rect 1951 1021 1955 1022
rect 2007 1026 2011 1027
rect 2007 1021 2011 1022
rect 2071 1026 2075 1027
rect 2071 1021 2075 1022
rect 2119 1026 2123 1027
rect 2119 1021 2123 1022
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 1094 1008 1100 1009
rect 1094 1004 1095 1008
rect 1099 1004 1100 1008
rect 1094 1003 1100 1004
rect 1136 1001 1138 1021
rect 1160 1009 1162 1021
rect 1232 1009 1234 1021
rect 1304 1009 1306 1021
rect 1384 1009 1386 1021
rect 1464 1009 1466 1021
rect 1544 1009 1546 1021
rect 1624 1009 1626 1021
rect 1696 1009 1698 1021
rect 1760 1009 1762 1021
rect 1824 1009 1826 1021
rect 1888 1009 1890 1021
rect 1952 1009 1954 1021
rect 1158 1008 1164 1009
rect 1158 1004 1159 1008
rect 1163 1004 1164 1008
rect 1158 1003 1164 1004
rect 1230 1008 1236 1009
rect 1230 1004 1231 1008
rect 1235 1004 1236 1008
rect 1230 1003 1236 1004
rect 1302 1008 1308 1009
rect 1302 1004 1303 1008
rect 1307 1004 1308 1008
rect 1302 1003 1308 1004
rect 1382 1008 1388 1009
rect 1382 1004 1383 1008
rect 1387 1004 1388 1008
rect 1382 1003 1388 1004
rect 1462 1008 1468 1009
rect 1462 1004 1463 1008
rect 1467 1004 1468 1008
rect 1462 1003 1468 1004
rect 1542 1008 1548 1009
rect 1542 1004 1543 1008
rect 1547 1004 1548 1008
rect 1542 1003 1548 1004
rect 1622 1008 1628 1009
rect 1622 1004 1623 1008
rect 1627 1004 1628 1008
rect 1622 1003 1628 1004
rect 1694 1008 1700 1009
rect 1694 1004 1695 1008
rect 1699 1004 1700 1008
rect 1694 1003 1700 1004
rect 1758 1008 1764 1009
rect 1758 1004 1759 1008
rect 1763 1004 1764 1008
rect 1758 1003 1764 1004
rect 1822 1008 1828 1009
rect 1822 1004 1823 1008
rect 1827 1004 1828 1008
rect 1822 1003 1828 1004
rect 1886 1008 1892 1009
rect 1886 1004 1887 1008
rect 1891 1004 1892 1008
rect 1886 1003 1892 1004
rect 1950 1008 1956 1009
rect 1950 1004 1951 1008
rect 1955 1004 1956 1008
rect 1950 1003 1956 1004
rect 2120 1001 2122 1021
rect 1134 1000 1140 1001
rect 1134 996 1135 1000
rect 1139 996 1140 1000
rect 1134 995 1140 996
rect 2118 1000 2124 1001
rect 2118 996 2119 1000
rect 2123 996 2124 1000
rect 2118 995 2124 996
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1094 991 1100 992
rect 110 986 116 987
rect 222 988 228 989
rect 112 979 114 986
rect 222 984 223 988
rect 227 984 228 988
rect 222 983 228 984
rect 270 988 276 989
rect 270 984 271 988
rect 275 984 276 988
rect 270 983 276 984
rect 334 988 340 989
rect 334 984 335 988
rect 339 984 340 988
rect 334 983 340 984
rect 406 988 412 989
rect 406 984 407 988
rect 411 984 412 988
rect 406 983 412 984
rect 478 988 484 989
rect 478 984 479 988
rect 483 984 484 988
rect 478 983 484 984
rect 558 988 564 989
rect 558 984 559 988
rect 563 984 564 988
rect 558 983 564 984
rect 630 988 636 989
rect 630 984 631 988
rect 635 984 636 988
rect 630 983 636 984
rect 702 988 708 989
rect 702 984 703 988
rect 707 984 708 988
rect 702 983 708 984
rect 774 988 780 989
rect 774 984 775 988
rect 779 984 780 988
rect 774 983 780 984
rect 838 988 844 989
rect 838 984 839 988
rect 843 984 844 988
rect 838 983 844 984
rect 902 988 908 989
rect 902 984 903 988
rect 907 984 908 988
rect 902 983 908 984
rect 966 988 972 989
rect 966 984 967 988
rect 971 984 972 988
rect 966 983 972 984
rect 1038 988 1044 989
rect 1038 984 1039 988
rect 1043 984 1044 988
rect 1094 987 1095 991
rect 1099 987 1100 991
rect 1094 986 1100 987
rect 1038 983 1044 984
rect 224 979 226 983
rect 272 979 274 983
rect 336 979 338 983
rect 408 979 410 983
rect 480 979 482 983
rect 560 979 562 983
rect 632 979 634 983
rect 704 979 706 983
rect 776 979 778 983
rect 840 979 842 983
rect 904 979 906 983
rect 968 979 970 983
rect 1040 979 1042 983
rect 1096 979 1098 986
rect 1134 983 1140 984
rect 1134 979 1135 983
rect 1139 979 1140 983
rect 2118 983 2124 984
rect 111 978 115 979
rect 111 973 115 974
rect 151 978 155 979
rect 151 973 155 974
rect 215 978 219 979
rect 215 973 219 974
rect 223 978 227 979
rect 223 973 227 974
rect 271 978 275 979
rect 271 973 275 974
rect 287 978 291 979
rect 287 973 291 974
rect 335 978 339 979
rect 335 973 339 974
rect 367 978 371 979
rect 367 973 371 974
rect 407 978 411 979
rect 407 973 411 974
rect 447 978 451 979
rect 447 973 451 974
rect 479 978 483 979
rect 479 973 483 974
rect 527 978 531 979
rect 527 973 531 974
rect 559 978 563 979
rect 559 973 563 974
rect 599 978 603 979
rect 599 973 603 974
rect 631 978 635 979
rect 631 973 635 974
rect 671 978 675 979
rect 671 973 675 974
rect 703 978 707 979
rect 703 973 707 974
rect 735 978 739 979
rect 735 973 739 974
rect 775 978 779 979
rect 775 973 779 974
rect 799 978 803 979
rect 799 973 803 974
rect 839 978 843 979
rect 839 973 843 974
rect 863 978 867 979
rect 863 973 867 974
rect 903 978 907 979
rect 903 973 907 974
rect 927 978 931 979
rect 927 973 931 974
rect 967 978 971 979
rect 967 973 971 974
rect 991 978 995 979
rect 991 973 995 974
rect 1039 978 1043 979
rect 1039 973 1043 974
rect 1047 978 1051 979
rect 1047 973 1051 974
rect 1095 978 1099 979
rect 1134 978 1140 979
rect 1158 980 1164 981
rect 1136 975 1138 978
rect 1158 976 1159 980
rect 1163 976 1164 980
rect 1158 975 1164 976
rect 1230 980 1236 981
rect 1230 976 1231 980
rect 1235 976 1236 980
rect 1230 975 1236 976
rect 1302 980 1308 981
rect 1302 976 1303 980
rect 1307 976 1308 980
rect 1302 975 1308 976
rect 1382 980 1388 981
rect 1382 976 1383 980
rect 1387 976 1388 980
rect 1382 975 1388 976
rect 1462 980 1468 981
rect 1462 976 1463 980
rect 1467 976 1468 980
rect 1462 975 1468 976
rect 1542 980 1548 981
rect 1542 976 1543 980
rect 1547 976 1548 980
rect 1542 975 1548 976
rect 1622 980 1628 981
rect 1622 976 1623 980
rect 1627 976 1628 980
rect 1622 975 1628 976
rect 1694 980 1700 981
rect 1694 976 1695 980
rect 1699 976 1700 980
rect 1694 975 1700 976
rect 1758 980 1764 981
rect 1758 976 1759 980
rect 1763 976 1764 980
rect 1758 975 1764 976
rect 1822 980 1828 981
rect 1822 976 1823 980
rect 1827 976 1828 980
rect 1822 975 1828 976
rect 1886 980 1892 981
rect 1886 976 1887 980
rect 1891 976 1892 980
rect 1886 975 1892 976
rect 1950 980 1956 981
rect 1950 976 1951 980
rect 1955 976 1956 980
rect 2118 979 2119 983
rect 2123 979 2124 983
rect 2118 978 2124 979
rect 1950 975 1956 976
rect 2120 975 2122 978
rect 1095 973 1099 974
rect 1135 974 1139 975
rect 112 970 114 973
rect 150 972 156 973
rect 110 969 116 970
rect 110 965 111 969
rect 115 965 116 969
rect 150 968 151 972
rect 155 968 156 972
rect 150 967 156 968
rect 214 972 220 973
rect 214 968 215 972
rect 219 968 220 972
rect 214 967 220 968
rect 286 972 292 973
rect 286 968 287 972
rect 291 968 292 972
rect 286 967 292 968
rect 366 972 372 973
rect 366 968 367 972
rect 371 968 372 972
rect 366 967 372 968
rect 446 972 452 973
rect 446 968 447 972
rect 451 968 452 972
rect 446 967 452 968
rect 526 972 532 973
rect 526 968 527 972
rect 531 968 532 972
rect 526 967 532 968
rect 598 972 604 973
rect 598 968 599 972
rect 603 968 604 972
rect 598 967 604 968
rect 670 972 676 973
rect 670 968 671 972
rect 675 968 676 972
rect 670 967 676 968
rect 734 972 740 973
rect 734 968 735 972
rect 739 968 740 972
rect 734 967 740 968
rect 798 972 804 973
rect 798 968 799 972
rect 803 968 804 972
rect 798 967 804 968
rect 862 972 868 973
rect 862 968 863 972
rect 867 968 868 972
rect 862 967 868 968
rect 926 972 932 973
rect 926 968 927 972
rect 931 968 932 972
rect 926 967 932 968
rect 990 972 996 973
rect 990 968 991 972
rect 995 968 996 972
rect 990 967 996 968
rect 1046 972 1052 973
rect 1046 968 1047 972
rect 1051 968 1052 972
rect 1096 970 1098 973
rect 1046 967 1052 968
rect 1094 969 1100 970
rect 1135 969 1139 970
rect 1159 974 1163 975
rect 1159 969 1163 970
rect 1231 974 1235 975
rect 1231 969 1235 970
rect 1239 974 1243 975
rect 1239 969 1243 970
rect 1303 974 1307 975
rect 1303 969 1307 970
rect 1375 974 1379 975
rect 1375 969 1379 970
rect 1383 974 1387 975
rect 1383 969 1387 970
rect 1439 974 1443 975
rect 1439 969 1443 970
rect 1463 974 1467 975
rect 1463 969 1467 970
rect 1511 974 1515 975
rect 1511 969 1515 970
rect 1543 974 1547 975
rect 1543 969 1547 970
rect 1583 974 1587 975
rect 1583 969 1587 970
rect 1623 974 1627 975
rect 1623 969 1627 970
rect 1655 974 1659 975
rect 1655 969 1659 970
rect 1695 974 1699 975
rect 1695 969 1699 970
rect 1727 974 1731 975
rect 1727 969 1731 970
rect 1759 974 1763 975
rect 1759 969 1763 970
rect 1799 974 1803 975
rect 1799 969 1803 970
rect 1823 974 1827 975
rect 1823 969 1827 970
rect 1871 974 1875 975
rect 1871 969 1875 970
rect 1887 974 1891 975
rect 1887 969 1891 970
rect 1943 974 1947 975
rect 1943 969 1947 970
rect 1951 974 1955 975
rect 1951 969 1955 970
rect 2015 974 2019 975
rect 2015 969 2019 970
rect 2071 974 2075 975
rect 2071 969 2075 970
rect 2119 974 2123 975
rect 2119 969 2123 970
rect 110 964 116 965
rect 1094 965 1095 969
rect 1099 965 1100 969
rect 1136 966 1138 969
rect 1238 968 1244 969
rect 1094 964 1100 965
rect 1134 965 1140 966
rect 1134 961 1135 965
rect 1139 961 1140 965
rect 1238 964 1239 968
rect 1243 964 1244 968
rect 1238 963 1244 964
rect 1302 968 1308 969
rect 1302 964 1303 968
rect 1307 964 1308 968
rect 1302 963 1308 964
rect 1374 968 1380 969
rect 1374 964 1375 968
rect 1379 964 1380 968
rect 1374 963 1380 964
rect 1438 968 1444 969
rect 1438 964 1439 968
rect 1443 964 1444 968
rect 1438 963 1444 964
rect 1510 968 1516 969
rect 1510 964 1511 968
rect 1515 964 1516 968
rect 1510 963 1516 964
rect 1582 968 1588 969
rect 1582 964 1583 968
rect 1587 964 1588 968
rect 1582 963 1588 964
rect 1654 968 1660 969
rect 1654 964 1655 968
rect 1659 964 1660 968
rect 1654 963 1660 964
rect 1726 968 1732 969
rect 1726 964 1727 968
rect 1731 964 1732 968
rect 1726 963 1732 964
rect 1798 968 1804 969
rect 1798 964 1799 968
rect 1803 964 1804 968
rect 1798 963 1804 964
rect 1870 968 1876 969
rect 1870 964 1871 968
rect 1875 964 1876 968
rect 1870 963 1876 964
rect 1942 968 1948 969
rect 1942 964 1943 968
rect 1947 964 1948 968
rect 1942 963 1948 964
rect 2014 968 2020 969
rect 2014 964 2015 968
rect 2019 964 2020 968
rect 2014 963 2020 964
rect 2070 968 2076 969
rect 2070 964 2071 968
rect 2075 964 2076 968
rect 2120 966 2122 969
rect 2070 963 2076 964
rect 2118 965 2124 966
rect 1134 960 1140 961
rect 2118 961 2119 965
rect 2123 961 2124 965
rect 2118 960 2124 961
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 110 947 116 948
rect 1094 952 1100 953
rect 1094 948 1095 952
rect 1099 948 1100 952
rect 1094 947 1100 948
rect 1134 948 1140 949
rect 112 927 114 947
rect 150 944 156 945
rect 150 940 151 944
rect 155 940 156 944
rect 150 939 156 940
rect 214 944 220 945
rect 214 940 215 944
rect 219 940 220 944
rect 214 939 220 940
rect 286 944 292 945
rect 286 940 287 944
rect 291 940 292 944
rect 286 939 292 940
rect 366 944 372 945
rect 366 940 367 944
rect 371 940 372 944
rect 366 939 372 940
rect 446 944 452 945
rect 446 940 447 944
rect 451 940 452 944
rect 446 939 452 940
rect 526 944 532 945
rect 526 940 527 944
rect 531 940 532 944
rect 526 939 532 940
rect 598 944 604 945
rect 598 940 599 944
rect 603 940 604 944
rect 598 939 604 940
rect 670 944 676 945
rect 670 940 671 944
rect 675 940 676 944
rect 670 939 676 940
rect 734 944 740 945
rect 734 940 735 944
rect 739 940 740 944
rect 734 939 740 940
rect 798 944 804 945
rect 798 940 799 944
rect 803 940 804 944
rect 798 939 804 940
rect 862 944 868 945
rect 862 940 863 944
rect 867 940 868 944
rect 862 939 868 940
rect 926 944 932 945
rect 926 940 927 944
rect 931 940 932 944
rect 926 939 932 940
rect 990 944 996 945
rect 990 940 991 944
rect 995 940 996 944
rect 990 939 996 940
rect 1046 944 1052 945
rect 1046 940 1047 944
rect 1051 940 1052 944
rect 1046 939 1052 940
rect 152 927 154 939
rect 216 927 218 939
rect 288 927 290 939
rect 368 927 370 939
rect 448 927 450 939
rect 528 927 530 939
rect 600 927 602 939
rect 672 927 674 939
rect 736 927 738 939
rect 800 927 802 939
rect 864 927 866 939
rect 928 927 930 939
rect 992 927 994 939
rect 1048 927 1050 939
rect 1096 927 1098 947
rect 1134 944 1135 948
rect 1139 944 1140 948
rect 1134 943 1140 944
rect 2118 948 2124 949
rect 2118 944 2119 948
rect 2123 944 2124 948
rect 2118 943 2124 944
rect 111 926 115 927
rect 111 921 115 922
rect 135 926 139 927
rect 135 921 139 922
rect 151 926 155 927
rect 151 921 155 922
rect 183 926 187 927
rect 183 921 187 922
rect 215 926 219 927
rect 215 921 219 922
rect 255 926 259 927
rect 255 921 259 922
rect 287 926 291 927
rect 287 921 291 922
rect 327 926 331 927
rect 327 921 331 922
rect 367 926 371 927
rect 367 921 371 922
rect 399 926 403 927
rect 399 921 403 922
rect 447 926 451 927
rect 447 921 451 922
rect 463 926 467 927
rect 463 921 467 922
rect 527 926 531 927
rect 527 921 531 922
rect 599 926 603 927
rect 599 921 603 922
rect 671 926 675 927
rect 671 921 675 922
rect 735 926 739 927
rect 735 921 739 922
rect 743 926 747 927
rect 743 921 747 922
rect 799 926 803 927
rect 799 921 803 922
rect 815 926 819 927
rect 815 921 819 922
rect 863 926 867 927
rect 863 921 867 922
rect 895 926 899 927
rect 895 921 899 922
rect 927 926 931 927
rect 927 921 931 922
rect 983 926 987 927
rect 983 921 987 922
rect 991 926 995 927
rect 991 921 995 922
rect 1047 926 1051 927
rect 1047 921 1051 922
rect 1095 926 1099 927
rect 1095 921 1099 922
rect 112 901 114 921
rect 136 909 138 921
rect 184 909 186 921
rect 256 909 258 921
rect 328 909 330 921
rect 400 909 402 921
rect 464 909 466 921
rect 528 909 530 921
rect 600 909 602 921
rect 672 909 674 921
rect 744 909 746 921
rect 816 909 818 921
rect 896 909 898 921
rect 984 909 986 921
rect 1048 909 1050 921
rect 134 908 140 909
rect 134 904 135 908
rect 139 904 140 908
rect 134 903 140 904
rect 182 908 188 909
rect 182 904 183 908
rect 187 904 188 908
rect 182 903 188 904
rect 254 908 260 909
rect 254 904 255 908
rect 259 904 260 908
rect 254 903 260 904
rect 326 908 332 909
rect 326 904 327 908
rect 331 904 332 908
rect 326 903 332 904
rect 398 908 404 909
rect 398 904 399 908
rect 403 904 404 908
rect 398 903 404 904
rect 462 908 468 909
rect 462 904 463 908
rect 467 904 468 908
rect 462 903 468 904
rect 526 908 532 909
rect 526 904 527 908
rect 531 904 532 908
rect 526 903 532 904
rect 598 908 604 909
rect 598 904 599 908
rect 603 904 604 908
rect 598 903 604 904
rect 670 908 676 909
rect 670 904 671 908
rect 675 904 676 908
rect 670 903 676 904
rect 742 908 748 909
rect 742 904 743 908
rect 747 904 748 908
rect 742 903 748 904
rect 814 908 820 909
rect 814 904 815 908
rect 819 904 820 908
rect 814 903 820 904
rect 894 908 900 909
rect 894 904 895 908
rect 899 904 900 908
rect 894 903 900 904
rect 982 908 988 909
rect 982 904 983 908
rect 987 904 988 908
rect 982 903 988 904
rect 1046 908 1052 909
rect 1046 904 1047 908
rect 1051 904 1052 908
rect 1046 903 1052 904
rect 1096 901 1098 921
rect 1136 919 1138 943
rect 1238 940 1244 941
rect 1238 936 1239 940
rect 1243 936 1244 940
rect 1238 935 1244 936
rect 1302 940 1308 941
rect 1302 936 1303 940
rect 1307 936 1308 940
rect 1302 935 1308 936
rect 1374 940 1380 941
rect 1374 936 1375 940
rect 1379 936 1380 940
rect 1374 935 1380 936
rect 1438 940 1444 941
rect 1438 936 1439 940
rect 1443 936 1444 940
rect 1438 935 1444 936
rect 1510 940 1516 941
rect 1510 936 1511 940
rect 1515 936 1516 940
rect 1510 935 1516 936
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1654 940 1660 941
rect 1654 936 1655 940
rect 1659 936 1660 940
rect 1654 935 1660 936
rect 1726 940 1732 941
rect 1726 936 1727 940
rect 1731 936 1732 940
rect 1726 935 1732 936
rect 1798 940 1804 941
rect 1798 936 1799 940
rect 1803 936 1804 940
rect 1798 935 1804 936
rect 1870 940 1876 941
rect 1870 936 1871 940
rect 1875 936 1876 940
rect 1870 935 1876 936
rect 1942 940 1948 941
rect 1942 936 1943 940
rect 1947 936 1948 940
rect 1942 935 1948 936
rect 2014 940 2020 941
rect 2014 936 2015 940
rect 2019 936 2020 940
rect 2014 935 2020 936
rect 2070 940 2076 941
rect 2070 936 2071 940
rect 2075 936 2076 940
rect 2070 935 2076 936
rect 1240 919 1242 935
rect 1304 919 1306 935
rect 1376 919 1378 935
rect 1440 919 1442 935
rect 1512 919 1514 935
rect 1584 919 1586 935
rect 1656 919 1658 935
rect 1728 919 1730 935
rect 1800 919 1802 935
rect 1872 919 1874 935
rect 1944 919 1946 935
rect 2016 919 2018 935
rect 2072 919 2074 935
rect 2120 919 2122 943
rect 1135 918 1139 919
rect 1135 913 1139 914
rect 1239 918 1243 919
rect 1239 913 1243 914
rect 1287 918 1291 919
rect 1287 913 1291 914
rect 1303 918 1307 919
rect 1303 913 1307 914
rect 1327 918 1331 919
rect 1327 913 1331 914
rect 1375 918 1379 919
rect 1375 913 1379 914
rect 1423 918 1427 919
rect 1423 913 1427 914
rect 1439 918 1443 919
rect 1439 913 1443 914
rect 1479 918 1483 919
rect 1479 913 1483 914
rect 1511 918 1515 919
rect 1511 913 1515 914
rect 1551 918 1555 919
rect 1551 913 1555 914
rect 1583 918 1587 919
rect 1583 913 1587 914
rect 1623 918 1627 919
rect 1623 913 1627 914
rect 1655 918 1659 919
rect 1655 913 1659 914
rect 1703 918 1707 919
rect 1703 913 1707 914
rect 1727 918 1731 919
rect 1727 913 1731 914
rect 1791 918 1795 919
rect 1791 913 1795 914
rect 1799 918 1803 919
rect 1799 913 1803 914
rect 1871 918 1875 919
rect 1871 913 1875 914
rect 1879 918 1883 919
rect 1879 913 1883 914
rect 1943 918 1947 919
rect 1943 913 1947 914
rect 1967 918 1971 919
rect 1967 913 1971 914
rect 2015 918 2019 919
rect 2015 913 2019 914
rect 2063 918 2067 919
rect 2063 913 2067 914
rect 2071 918 2075 919
rect 2071 913 2075 914
rect 2119 918 2123 919
rect 2119 913 2123 914
rect 110 900 116 901
rect 110 896 111 900
rect 115 896 116 900
rect 110 895 116 896
rect 1094 900 1100 901
rect 1094 896 1095 900
rect 1099 896 1100 900
rect 1094 895 1100 896
rect 1136 893 1138 913
rect 1288 901 1290 913
rect 1328 901 1330 913
rect 1376 901 1378 913
rect 1424 901 1426 913
rect 1480 901 1482 913
rect 1552 901 1554 913
rect 1624 901 1626 913
rect 1704 901 1706 913
rect 1792 901 1794 913
rect 1880 901 1882 913
rect 1968 901 1970 913
rect 2064 901 2066 913
rect 1286 900 1292 901
rect 1286 896 1287 900
rect 1291 896 1292 900
rect 1286 895 1292 896
rect 1326 900 1332 901
rect 1326 896 1327 900
rect 1331 896 1332 900
rect 1326 895 1332 896
rect 1374 900 1380 901
rect 1374 896 1375 900
rect 1379 896 1380 900
rect 1374 895 1380 896
rect 1422 900 1428 901
rect 1422 896 1423 900
rect 1427 896 1428 900
rect 1422 895 1428 896
rect 1478 900 1484 901
rect 1478 896 1479 900
rect 1483 896 1484 900
rect 1478 895 1484 896
rect 1550 900 1556 901
rect 1550 896 1551 900
rect 1555 896 1556 900
rect 1550 895 1556 896
rect 1622 900 1628 901
rect 1622 896 1623 900
rect 1627 896 1628 900
rect 1622 895 1628 896
rect 1702 900 1708 901
rect 1702 896 1703 900
rect 1707 896 1708 900
rect 1702 895 1708 896
rect 1790 900 1796 901
rect 1790 896 1791 900
rect 1795 896 1796 900
rect 1790 895 1796 896
rect 1878 900 1884 901
rect 1878 896 1879 900
rect 1883 896 1884 900
rect 1878 895 1884 896
rect 1966 900 1972 901
rect 1966 896 1967 900
rect 1971 896 1972 900
rect 1966 895 1972 896
rect 2062 900 2068 901
rect 2062 896 2063 900
rect 2067 896 2068 900
rect 2062 895 2068 896
rect 2120 893 2122 913
rect 1134 892 1140 893
rect 1134 888 1135 892
rect 1139 888 1140 892
rect 1134 887 1140 888
rect 2118 892 2124 893
rect 2118 888 2119 892
rect 2123 888 2124 892
rect 2118 887 2124 888
rect 110 883 116 884
rect 110 879 111 883
rect 115 879 116 883
rect 1094 883 1100 884
rect 110 878 116 879
rect 134 880 140 881
rect 112 871 114 878
rect 134 876 135 880
rect 139 876 140 880
rect 134 875 140 876
rect 182 880 188 881
rect 182 876 183 880
rect 187 876 188 880
rect 182 875 188 876
rect 254 880 260 881
rect 254 876 255 880
rect 259 876 260 880
rect 254 875 260 876
rect 326 880 332 881
rect 326 876 327 880
rect 331 876 332 880
rect 326 875 332 876
rect 398 880 404 881
rect 398 876 399 880
rect 403 876 404 880
rect 398 875 404 876
rect 462 880 468 881
rect 462 876 463 880
rect 467 876 468 880
rect 462 875 468 876
rect 526 880 532 881
rect 526 876 527 880
rect 531 876 532 880
rect 526 875 532 876
rect 598 880 604 881
rect 598 876 599 880
rect 603 876 604 880
rect 598 875 604 876
rect 670 880 676 881
rect 670 876 671 880
rect 675 876 676 880
rect 670 875 676 876
rect 742 880 748 881
rect 742 876 743 880
rect 747 876 748 880
rect 742 875 748 876
rect 814 880 820 881
rect 814 876 815 880
rect 819 876 820 880
rect 814 875 820 876
rect 894 880 900 881
rect 894 876 895 880
rect 899 876 900 880
rect 894 875 900 876
rect 982 880 988 881
rect 982 876 983 880
rect 987 876 988 880
rect 982 875 988 876
rect 1046 880 1052 881
rect 1046 876 1047 880
rect 1051 876 1052 880
rect 1094 879 1095 883
rect 1099 879 1100 883
rect 1094 878 1100 879
rect 1046 875 1052 876
rect 136 871 138 875
rect 184 871 186 875
rect 256 871 258 875
rect 328 871 330 875
rect 400 871 402 875
rect 464 871 466 875
rect 528 871 530 875
rect 600 871 602 875
rect 672 871 674 875
rect 744 871 746 875
rect 816 871 818 875
rect 896 871 898 875
rect 984 871 986 875
rect 1048 871 1050 875
rect 1096 871 1098 878
rect 1134 875 1140 876
rect 1134 871 1135 875
rect 1139 871 1140 875
rect 2118 875 2124 876
rect 111 870 115 871
rect 111 865 115 866
rect 135 870 139 871
rect 135 865 139 866
rect 175 870 179 871
rect 175 865 179 866
rect 183 870 187 871
rect 183 865 187 866
rect 215 870 219 871
rect 215 865 219 866
rect 255 870 259 871
rect 255 865 259 866
rect 279 870 283 871
rect 279 865 283 866
rect 327 870 331 871
rect 327 865 331 866
rect 343 870 347 871
rect 343 865 347 866
rect 399 870 403 871
rect 399 865 403 866
rect 463 870 467 871
rect 463 865 467 866
rect 527 870 531 871
rect 527 865 531 866
rect 535 870 539 871
rect 535 865 539 866
rect 599 870 603 871
rect 599 865 603 866
rect 615 870 619 871
rect 615 865 619 866
rect 671 870 675 871
rect 671 865 675 866
rect 711 870 715 871
rect 711 865 715 866
rect 743 870 747 871
rect 743 865 747 866
rect 815 870 819 871
rect 815 865 819 866
rect 823 870 827 871
rect 823 865 827 866
rect 895 870 899 871
rect 895 865 899 866
rect 943 870 947 871
rect 943 865 947 866
rect 983 870 987 871
rect 983 865 987 866
rect 1047 870 1051 871
rect 1047 865 1051 866
rect 1095 870 1099 871
rect 1134 870 1140 871
rect 1286 872 1292 873
rect 1136 867 1138 870
rect 1286 868 1287 872
rect 1291 868 1292 872
rect 1286 867 1292 868
rect 1326 872 1332 873
rect 1326 868 1327 872
rect 1331 868 1332 872
rect 1326 867 1332 868
rect 1374 872 1380 873
rect 1374 868 1375 872
rect 1379 868 1380 872
rect 1374 867 1380 868
rect 1422 872 1428 873
rect 1422 868 1423 872
rect 1427 868 1428 872
rect 1422 867 1428 868
rect 1478 872 1484 873
rect 1478 868 1479 872
rect 1483 868 1484 872
rect 1478 867 1484 868
rect 1550 872 1556 873
rect 1550 868 1551 872
rect 1555 868 1556 872
rect 1550 867 1556 868
rect 1622 872 1628 873
rect 1622 868 1623 872
rect 1627 868 1628 872
rect 1622 867 1628 868
rect 1702 872 1708 873
rect 1702 868 1703 872
rect 1707 868 1708 872
rect 1702 867 1708 868
rect 1790 872 1796 873
rect 1790 868 1791 872
rect 1795 868 1796 872
rect 1790 867 1796 868
rect 1878 872 1884 873
rect 1878 868 1879 872
rect 1883 868 1884 872
rect 1878 867 1884 868
rect 1966 872 1972 873
rect 1966 868 1967 872
rect 1971 868 1972 872
rect 1966 867 1972 868
rect 2062 872 2068 873
rect 2062 868 2063 872
rect 2067 868 2068 872
rect 2118 871 2119 875
rect 2123 871 2124 875
rect 2118 870 2124 871
rect 2062 867 2068 868
rect 2120 867 2122 870
rect 1095 865 1099 866
rect 1135 866 1139 867
rect 112 862 114 865
rect 134 864 140 865
rect 110 861 116 862
rect 110 857 111 861
rect 115 857 116 861
rect 134 860 135 864
rect 139 860 140 864
rect 134 859 140 860
rect 174 864 180 865
rect 174 860 175 864
rect 179 860 180 864
rect 174 859 180 860
rect 214 864 220 865
rect 214 860 215 864
rect 219 860 220 864
rect 214 859 220 860
rect 278 864 284 865
rect 278 860 279 864
rect 283 860 284 864
rect 278 859 284 860
rect 342 864 348 865
rect 342 860 343 864
rect 347 860 348 864
rect 342 859 348 860
rect 398 864 404 865
rect 398 860 399 864
rect 403 860 404 864
rect 398 859 404 860
rect 462 864 468 865
rect 462 860 463 864
rect 467 860 468 864
rect 462 859 468 860
rect 534 864 540 865
rect 534 860 535 864
rect 539 860 540 864
rect 534 859 540 860
rect 614 864 620 865
rect 614 860 615 864
rect 619 860 620 864
rect 614 859 620 860
rect 710 864 716 865
rect 710 860 711 864
rect 715 860 716 864
rect 710 859 716 860
rect 822 864 828 865
rect 822 860 823 864
rect 827 860 828 864
rect 822 859 828 860
rect 942 864 948 865
rect 942 860 943 864
rect 947 860 948 864
rect 942 859 948 860
rect 1046 864 1052 865
rect 1046 860 1047 864
rect 1051 860 1052 864
rect 1096 862 1098 865
rect 1046 859 1052 860
rect 1094 861 1100 862
rect 1135 861 1139 862
rect 1159 866 1163 867
rect 1159 861 1163 862
rect 1199 866 1203 867
rect 1199 861 1203 862
rect 1263 866 1267 867
rect 1263 861 1267 862
rect 1287 866 1291 867
rect 1287 861 1291 862
rect 1327 866 1331 867
rect 1327 861 1331 862
rect 1375 866 1379 867
rect 1375 861 1379 862
rect 1399 866 1403 867
rect 1399 861 1403 862
rect 1423 866 1427 867
rect 1423 861 1427 862
rect 1471 866 1475 867
rect 1471 861 1475 862
rect 1479 866 1483 867
rect 1479 861 1483 862
rect 1543 866 1547 867
rect 1543 861 1547 862
rect 1551 866 1555 867
rect 1551 861 1555 862
rect 1623 866 1627 867
rect 1623 861 1627 862
rect 1703 866 1707 867
rect 1703 861 1707 862
rect 1775 866 1779 867
rect 1775 861 1779 862
rect 1791 866 1795 867
rect 1791 861 1795 862
rect 1855 866 1859 867
rect 1855 861 1859 862
rect 1879 866 1883 867
rect 1879 861 1883 862
rect 1935 866 1939 867
rect 1935 861 1939 862
rect 1967 866 1971 867
rect 1967 861 1971 862
rect 2015 866 2019 867
rect 2015 861 2019 862
rect 2063 866 2067 867
rect 2063 861 2067 862
rect 2071 866 2075 867
rect 2071 861 2075 862
rect 2119 866 2123 867
rect 2119 861 2123 862
rect 110 856 116 857
rect 1094 857 1095 861
rect 1099 857 1100 861
rect 1136 858 1138 861
rect 1158 860 1164 861
rect 1094 856 1100 857
rect 1134 857 1140 858
rect 1134 853 1135 857
rect 1139 853 1140 857
rect 1158 856 1159 860
rect 1163 856 1164 860
rect 1158 855 1164 856
rect 1198 860 1204 861
rect 1198 856 1199 860
rect 1203 856 1204 860
rect 1198 855 1204 856
rect 1262 860 1268 861
rect 1262 856 1263 860
rect 1267 856 1268 860
rect 1262 855 1268 856
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1398 860 1404 861
rect 1398 856 1399 860
rect 1403 856 1404 860
rect 1398 855 1404 856
rect 1470 860 1476 861
rect 1470 856 1471 860
rect 1475 856 1476 860
rect 1470 855 1476 856
rect 1542 860 1548 861
rect 1542 856 1543 860
rect 1547 856 1548 860
rect 1542 855 1548 856
rect 1622 860 1628 861
rect 1622 856 1623 860
rect 1627 856 1628 860
rect 1622 855 1628 856
rect 1702 860 1708 861
rect 1702 856 1703 860
rect 1707 856 1708 860
rect 1702 855 1708 856
rect 1774 860 1780 861
rect 1774 856 1775 860
rect 1779 856 1780 860
rect 1774 855 1780 856
rect 1854 860 1860 861
rect 1854 856 1855 860
rect 1859 856 1860 860
rect 1854 855 1860 856
rect 1934 860 1940 861
rect 1934 856 1935 860
rect 1939 856 1940 860
rect 1934 855 1940 856
rect 2014 860 2020 861
rect 2014 856 2015 860
rect 2019 856 2020 860
rect 2014 855 2020 856
rect 2070 860 2076 861
rect 2070 856 2071 860
rect 2075 856 2076 860
rect 2120 858 2122 861
rect 2070 855 2076 856
rect 2118 857 2124 858
rect 1134 852 1140 853
rect 2118 853 2119 857
rect 2123 853 2124 857
rect 2118 852 2124 853
rect 110 844 116 845
rect 110 840 111 844
rect 115 840 116 844
rect 110 839 116 840
rect 1094 844 1100 845
rect 1094 840 1095 844
rect 1099 840 1100 844
rect 1094 839 1100 840
rect 1134 840 1140 841
rect 112 819 114 839
rect 134 836 140 837
rect 134 832 135 836
rect 139 832 140 836
rect 134 831 140 832
rect 174 836 180 837
rect 174 832 175 836
rect 179 832 180 836
rect 174 831 180 832
rect 214 836 220 837
rect 214 832 215 836
rect 219 832 220 836
rect 214 831 220 832
rect 278 836 284 837
rect 278 832 279 836
rect 283 832 284 836
rect 278 831 284 832
rect 342 836 348 837
rect 342 832 343 836
rect 347 832 348 836
rect 342 831 348 832
rect 398 836 404 837
rect 398 832 399 836
rect 403 832 404 836
rect 398 831 404 832
rect 462 836 468 837
rect 462 832 463 836
rect 467 832 468 836
rect 462 831 468 832
rect 534 836 540 837
rect 534 832 535 836
rect 539 832 540 836
rect 534 831 540 832
rect 614 836 620 837
rect 614 832 615 836
rect 619 832 620 836
rect 614 831 620 832
rect 710 836 716 837
rect 710 832 711 836
rect 715 832 716 836
rect 710 831 716 832
rect 822 836 828 837
rect 822 832 823 836
rect 827 832 828 836
rect 822 831 828 832
rect 942 836 948 837
rect 942 832 943 836
rect 947 832 948 836
rect 942 831 948 832
rect 1046 836 1052 837
rect 1046 832 1047 836
rect 1051 832 1052 836
rect 1046 831 1052 832
rect 136 819 138 831
rect 176 819 178 831
rect 216 819 218 831
rect 280 819 282 831
rect 344 819 346 831
rect 400 819 402 831
rect 464 819 466 831
rect 536 819 538 831
rect 616 819 618 831
rect 712 819 714 831
rect 824 819 826 831
rect 944 819 946 831
rect 1048 819 1050 831
rect 1096 819 1098 839
rect 1134 836 1135 840
rect 1139 836 1140 840
rect 1134 835 1140 836
rect 2118 840 2124 841
rect 2118 836 2119 840
rect 2123 836 2124 840
rect 2118 835 2124 836
rect 111 818 115 819
rect 111 813 115 814
rect 135 818 139 819
rect 135 813 139 814
rect 175 818 179 819
rect 175 813 179 814
rect 215 818 219 819
rect 215 813 219 814
rect 279 818 283 819
rect 279 813 283 814
rect 335 818 339 819
rect 335 813 339 814
rect 343 818 347 819
rect 343 813 347 814
rect 391 818 395 819
rect 391 813 395 814
rect 399 818 403 819
rect 399 813 403 814
rect 455 818 459 819
rect 455 813 459 814
rect 463 818 467 819
rect 463 813 467 814
rect 519 818 523 819
rect 519 813 523 814
rect 535 818 539 819
rect 535 813 539 814
rect 583 818 587 819
rect 583 813 587 814
rect 615 818 619 819
rect 615 813 619 814
rect 655 818 659 819
rect 655 813 659 814
rect 711 818 715 819
rect 711 813 715 814
rect 735 818 739 819
rect 735 813 739 814
rect 815 818 819 819
rect 815 813 819 814
rect 823 818 827 819
rect 823 813 827 814
rect 895 818 899 819
rect 895 813 899 814
rect 943 818 947 819
rect 943 813 947 814
rect 983 818 987 819
rect 983 813 987 814
rect 1047 818 1051 819
rect 1047 813 1051 814
rect 1095 818 1099 819
rect 1095 813 1099 814
rect 112 793 114 813
rect 136 801 138 813
rect 176 801 178 813
rect 216 801 218 813
rect 280 801 282 813
rect 336 801 338 813
rect 392 801 394 813
rect 456 801 458 813
rect 520 801 522 813
rect 584 801 586 813
rect 656 801 658 813
rect 736 801 738 813
rect 816 801 818 813
rect 896 801 898 813
rect 984 801 986 813
rect 1048 801 1050 813
rect 134 800 140 801
rect 134 796 135 800
rect 139 796 140 800
rect 134 795 140 796
rect 174 800 180 801
rect 174 796 175 800
rect 179 796 180 800
rect 174 795 180 796
rect 214 800 220 801
rect 214 796 215 800
rect 219 796 220 800
rect 214 795 220 796
rect 278 800 284 801
rect 278 796 279 800
rect 283 796 284 800
rect 278 795 284 796
rect 334 800 340 801
rect 334 796 335 800
rect 339 796 340 800
rect 334 795 340 796
rect 390 800 396 801
rect 390 796 391 800
rect 395 796 396 800
rect 390 795 396 796
rect 454 800 460 801
rect 454 796 455 800
rect 459 796 460 800
rect 454 795 460 796
rect 518 800 524 801
rect 518 796 519 800
rect 523 796 524 800
rect 518 795 524 796
rect 582 800 588 801
rect 582 796 583 800
rect 587 796 588 800
rect 582 795 588 796
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 654 795 660 796
rect 734 800 740 801
rect 734 796 735 800
rect 739 796 740 800
rect 734 795 740 796
rect 814 800 820 801
rect 814 796 815 800
rect 819 796 820 800
rect 814 795 820 796
rect 894 800 900 801
rect 894 796 895 800
rect 899 796 900 800
rect 894 795 900 796
rect 982 800 988 801
rect 982 796 983 800
rect 987 796 988 800
rect 982 795 988 796
rect 1046 800 1052 801
rect 1046 796 1047 800
rect 1051 796 1052 800
rect 1046 795 1052 796
rect 1096 793 1098 813
rect 1136 807 1138 835
rect 1158 832 1164 833
rect 1158 828 1159 832
rect 1163 828 1164 832
rect 1158 827 1164 828
rect 1198 832 1204 833
rect 1198 828 1199 832
rect 1203 828 1204 832
rect 1198 827 1204 828
rect 1262 832 1268 833
rect 1262 828 1263 832
rect 1267 828 1268 832
rect 1262 827 1268 828
rect 1326 832 1332 833
rect 1326 828 1327 832
rect 1331 828 1332 832
rect 1326 827 1332 828
rect 1398 832 1404 833
rect 1398 828 1399 832
rect 1403 828 1404 832
rect 1398 827 1404 828
rect 1470 832 1476 833
rect 1470 828 1471 832
rect 1475 828 1476 832
rect 1470 827 1476 828
rect 1542 832 1548 833
rect 1542 828 1543 832
rect 1547 828 1548 832
rect 1542 827 1548 828
rect 1622 832 1628 833
rect 1622 828 1623 832
rect 1627 828 1628 832
rect 1622 827 1628 828
rect 1702 832 1708 833
rect 1702 828 1703 832
rect 1707 828 1708 832
rect 1702 827 1708 828
rect 1774 832 1780 833
rect 1774 828 1775 832
rect 1779 828 1780 832
rect 1774 827 1780 828
rect 1854 832 1860 833
rect 1854 828 1855 832
rect 1859 828 1860 832
rect 1854 827 1860 828
rect 1934 832 1940 833
rect 1934 828 1935 832
rect 1939 828 1940 832
rect 1934 827 1940 828
rect 2014 832 2020 833
rect 2014 828 2015 832
rect 2019 828 2020 832
rect 2014 827 2020 828
rect 2070 832 2076 833
rect 2070 828 2071 832
rect 2075 828 2076 832
rect 2070 827 2076 828
rect 1160 807 1162 827
rect 1200 807 1202 827
rect 1264 807 1266 827
rect 1328 807 1330 827
rect 1400 807 1402 827
rect 1472 807 1474 827
rect 1544 807 1546 827
rect 1624 807 1626 827
rect 1704 807 1706 827
rect 1776 807 1778 827
rect 1856 807 1858 827
rect 1936 807 1938 827
rect 2016 807 2018 827
rect 2072 807 2074 827
rect 2120 807 2122 835
rect 1135 806 1139 807
rect 1135 801 1139 802
rect 1159 806 1163 807
rect 1159 801 1163 802
rect 1199 806 1203 807
rect 1199 801 1203 802
rect 1239 806 1243 807
rect 1239 801 1243 802
rect 1263 806 1267 807
rect 1263 801 1267 802
rect 1327 806 1331 807
rect 1327 801 1331 802
rect 1343 806 1347 807
rect 1343 801 1347 802
rect 1399 806 1403 807
rect 1399 801 1403 802
rect 1447 806 1451 807
rect 1447 801 1451 802
rect 1471 806 1475 807
rect 1471 801 1475 802
rect 1543 806 1547 807
rect 1543 801 1547 802
rect 1551 806 1555 807
rect 1551 801 1555 802
rect 1623 806 1627 807
rect 1623 801 1627 802
rect 1655 806 1659 807
rect 1655 801 1659 802
rect 1703 806 1707 807
rect 1703 801 1707 802
rect 1751 806 1755 807
rect 1751 801 1755 802
rect 1775 806 1779 807
rect 1775 801 1779 802
rect 1839 806 1843 807
rect 1839 801 1843 802
rect 1855 806 1859 807
rect 1855 801 1859 802
rect 1919 806 1923 807
rect 1919 801 1923 802
rect 1935 806 1939 807
rect 1935 801 1939 802
rect 2007 806 2011 807
rect 2007 801 2011 802
rect 2015 806 2019 807
rect 2015 801 2019 802
rect 2071 806 2075 807
rect 2071 801 2075 802
rect 2119 806 2123 807
rect 2119 801 2123 802
rect 110 792 116 793
rect 110 788 111 792
rect 115 788 116 792
rect 110 787 116 788
rect 1094 792 1100 793
rect 1094 788 1095 792
rect 1099 788 1100 792
rect 1094 787 1100 788
rect 1136 781 1138 801
rect 1160 789 1162 801
rect 1240 789 1242 801
rect 1344 789 1346 801
rect 1448 789 1450 801
rect 1552 789 1554 801
rect 1656 789 1658 801
rect 1752 789 1754 801
rect 1840 789 1842 801
rect 1920 789 1922 801
rect 2008 789 2010 801
rect 2072 789 2074 801
rect 1158 788 1164 789
rect 1158 784 1159 788
rect 1163 784 1164 788
rect 1158 783 1164 784
rect 1238 788 1244 789
rect 1238 784 1239 788
rect 1243 784 1244 788
rect 1238 783 1244 784
rect 1342 788 1348 789
rect 1342 784 1343 788
rect 1347 784 1348 788
rect 1342 783 1348 784
rect 1446 788 1452 789
rect 1446 784 1447 788
rect 1451 784 1452 788
rect 1446 783 1452 784
rect 1550 788 1556 789
rect 1550 784 1551 788
rect 1555 784 1556 788
rect 1550 783 1556 784
rect 1654 788 1660 789
rect 1654 784 1655 788
rect 1659 784 1660 788
rect 1654 783 1660 784
rect 1750 788 1756 789
rect 1750 784 1751 788
rect 1755 784 1756 788
rect 1750 783 1756 784
rect 1838 788 1844 789
rect 1838 784 1839 788
rect 1843 784 1844 788
rect 1838 783 1844 784
rect 1918 788 1924 789
rect 1918 784 1919 788
rect 1923 784 1924 788
rect 1918 783 1924 784
rect 2006 788 2012 789
rect 2006 784 2007 788
rect 2011 784 2012 788
rect 2006 783 2012 784
rect 2070 788 2076 789
rect 2070 784 2071 788
rect 2075 784 2076 788
rect 2070 783 2076 784
rect 2120 781 2122 801
rect 1134 780 1140 781
rect 1134 776 1135 780
rect 1139 776 1140 780
rect 110 775 116 776
rect 110 771 111 775
rect 115 771 116 775
rect 1094 775 1100 776
rect 1134 775 1140 776
rect 2118 780 2124 781
rect 2118 776 2119 780
rect 2123 776 2124 780
rect 2118 775 2124 776
rect 110 770 116 771
rect 134 772 140 773
rect 112 767 114 770
rect 134 768 135 772
rect 139 768 140 772
rect 134 767 140 768
rect 174 772 180 773
rect 174 768 175 772
rect 179 768 180 772
rect 174 767 180 768
rect 214 772 220 773
rect 214 768 215 772
rect 219 768 220 772
rect 214 767 220 768
rect 278 772 284 773
rect 278 768 279 772
rect 283 768 284 772
rect 278 767 284 768
rect 334 772 340 773
rect 334 768 335 772
rect 339 768 340 772
rect 334 767 340 768
rect 390 772 396 773
rect 390 768 391 772
rect 395 768 396 772
rect 390 767 396 768
rect 454 772 460 773
rect 454 768 455 772
rect 459 768 460 772
rect 454 767 460 768
rect 518 772 524 773
rect 518 768 519 772
rect 523 768 524 772
rect 518 767 524 768
rect 582 772 588 773
rect 582 768 583 772
rect 587 768 588 772
rect 582 767 588 768
rect 654 772 660 773
rect 654 768 655 772
rect 659 768 660 772
rect 654 767 660 768
rect 734 772 740 773
rect 734 768 735 772
rect 739 768 740 772
rect 734 767 740 768
rect 814 772 820 773
rect 814 768 815 772
rect 819 768 820 772
rect 814 767 820 768
rect 894 772 900 773
rect 894 768 895 772
rect 899 768 900 772
rect 894 767 900 768
rect 982 772 988 773
rect 982 768 983 772
rect 987 768 988 772
rect 982 767 988 768
rect 1046 772 1052 773
rect 1046 768 1047 772
rect 1051 768 1052 772
rect 1094 771 1095 775
rect 1099 771 1100 775
rect 1094 770 1100 771
rect 1046 767 1052 768
rect 1096 767 1098 770
rect 111 766 115 767
rect 111 761 115 762
rect 135 766 139 767
rect 135 761 139 762
rect 175 766 179 767
rect 175 761 179 762
rect 207 766 211 767
rect 207 761 211 762
rect 215 766 219 767
rect 215 761 219 762
rect 279 766 283 767
rect 279 761 283 762
rect 295 766 299 767
rect 295 761 299 762
rect 335 766 339 767
rect 335 761 339 762
rect 375 766 379 767
rect 375 761 379 762
rect 391 766 395 767
rect 391 761 395 762
rect 447 766 451 767
rect 447 761 451 762
rect 455 766 459 767
rect 455 761 459 762
rect 519 766 523 767
rect 519 761 523 762
rect 583 766 587 767
rect 583 761 587 762
rect 639 766 643 767
rect 639 761 643 762
rect 655 766 659 767
rect 655 761 659 762
rect 687 766 691 767
rect 687 761 691 762
rect 735 766 739 767
rect 735 761 739 762
rect 743 766 747 767
rect 743 761 747 762
rect 799 766 803 767
rect 799 761 803 762
rect 815 766 819 767
rect 815 761 819 762
rect 855 766 859 767
rect 855 761 859 762
rect 895 766 899 767
rect 895 761 899 762
rect 983 766 987 767
rect 983 761 987 762
rect 1047 766 1051 767
rect 1047 761 1051 762
rect 1095 766 1099 767
rect 1095 761 1099 762
rect 1134 763 1140 764
rect 112 758 114 761
rect 134 760 140 761
rect 110 757 116 758
rect 110 753 111 757
rect 115 753 116 757
rect 134 756 135 760
rect 139 756 140 760
rect 134 755 140 756
rect 206 760 212 761
rect 206 756 207 760
rect 211 756 212 760
rect 206 755 212 756
rect 294 760 300 761
rect 294 756 295 760
rect 299 756 300 760
rect 294 755 300 756
rect 374 760 380 761
rect 374 756 375 760
rect 379 756 380 760
rect 374 755 380 756
rect 446 760 452 761
rect 446 756 447 760
rect 451 756 452 760
rect 446 755 452 756
rect 518 760 524 761
rect 518 756 519 760
rect 523 756 524 760
rect 518 755 524 756
rect 582 760 588 761
rect 582 756 583 760
rect 587 756 588 760
rect 582 755 588 756
rect 638 760 644 761
rect 638 756 639 760
rect 643 756 644 760
rect 638 755 644 756
rect 686 760 692 761
rect 686 756 687 760
rect 691 756 692 760
rect 686 755 692 756
rect 742 760 748 761
rect 742 756 743 760
rect 747 756 748 760
rect 742 755 748 756
rect 798 760 804 761
rect 798 756 799 760
rect 803 756 804 760
rect 798 755 804 756
rect 854 760 860 761
rect 854 756 855 760
rect 859 756 860 760
rect 1096 758 1098 761
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 2118 763 2124 764
rect 1134 758 1140 759
rect 1158 760 1164 761
rect 854 755 860 756
rect 1094 757 1100 758
rect 110 752 116 753
rect 1094 753 1095 757
rect 1099 753 1100 757
rect 1136 755 1138 758
rect 1158 756 1159 760
rect 1163 756 1164 760
rect 1158 755 1164 756
rect 1238 760 1244 761
rect 1238 756 1239 760
rect 1243 756 1244 760
rect 1238 755 1244 756
rect 1342 760 1348 761
rect 1342 756 1343 760
rect 1347 756 1348 760
rect 1342 755 1348 756
rect 1446 760 1452 761
rect 1446 756 1447 760
rect 1451 756 1452 760
rect 1446 755 1452 756
rect 1550 760 1556 761
rect 1550 756 1551 760
rect 1555 756 1556 760
rect 1550 755 1556 756
rect 1654 760 1660 761
rect 1654 756 1655 760
rect 1659 756 1660 760
rect 1654 755 1660 756
rect 1750 760 1756 761
rect 1750 756 1751 760
rect 1755 756 1756 760
rect 1750 755 1756 756
rect 1838 760 1844 761
rect 1838 756 1839 760
rect 1843 756 1844 760
rect 1838 755 1844 756
rect 1918 760 1924 761
rect 1918 756 1919 760
rect 1923 756 1924 760
rect 1918 755 1924 756
rect 2006 760 2012 761
rect 2006 756 2007 760
rect 2011 756 2012 760
rect 2006 755 2012 756
rect 2070 760 2076 761
rect 2070 756 2071 760
rect 2075 756 2076 760
rect 2118 759 2119 763
rect 2123 759 2124 763
rect 2118 758 2124 759
rect 2070 755 2076 756
rect 2120 755 2122 758
rect 1094 752 1100 753
rect 1135 754 1139 755
rect 1135 749 1139 750
rect 1159 754 1163 755
rect 1159 749 1163 750
rect 1199 754 1203 755
rect 1199 749 1203 750
rect 1239 754 1243 755
rect 1239 749 1243 750
rect 1287 754 1291 755
rect 1287 749 1291 750
rect 1343 754 1347 755
rect 1343 749 1347 750
rect 1359 754 1363 755
rect 1359 749 1363 750
rect 1439 754 1443 755
rect 1439 749 1443 750
rect 1447 754 1451 755
rect 1447 749 1451 750
rect 1527 754 1531 755
rect 1527 749 1531 750
rect 1551 754 1555 755
rect 1551 749 1555 750
rect 1615 754 1619 755
rect 1615 749 1619 750
rect 1655 754 1659 755
rect 1655 749 1659 750
rect 1711 754 1715 755
rect 1711 749 1715 750
rect 1751 754 1755 755
rect 1751 749 1755 750
rect 1807 754 1811 755
rect 1807 749 1811 750
rect 1839 754 1843 755
rect 1839 749 1843 750
rect 1903 754 1907 755
rect 1903 749 1907 750
rect 1919 754 1923 755
rect 1919 749 1923 750
rect 1999 754 2003 755
rect 1999 749 2003 750
rect 2007 754 2011 755
rect 2007 749 2011 750
rect 2071 754 2075 755
rect 2071 749 2075 750
rect 2119 754 2123 755
rect 2119 749 2123 750
rect 1136 746 1138 749
rect 1158 748 1164 749
rect 1134 745 1140 746
rect 1134 741 1135 745
rect 1139 741 1140 745
rect 1158 744 1159 748
rect 1163 744 1164 748
rect 1158 743 1164 744
rect 1198 748 1204 749
rect 1198 744 1199 748
rect 1203 744 1204 748
rect 1198 743 1204 744
rect 1238 748 1244 749
rect 1238 744 1239 748
rect 1243 744 1244 748
rect 1238 743 1244 744
rect 1286 748 1292 749
rect 1286 744 1287 748
rect 1291 744 1292 748
rect 1286 743 1292 744
rect 1358 748 1364 749
rect 1358 744 1359 748
rect 1363 744 1364 748
rect 1358 743 1364 744
rect 1438 748 1444 749
rect 1438 744 1439 748
rect 1443 744 1444 748
rect 1438 743 1444 744
rect 1526 748 1532 749
rect 1526 744 1527 748
rect 1531 744 1532 748
rect 1526 743 1532 744
rect 1614 748 1620 749
rect 1614 744 1615 748
rect 1619 744 1620 748
rect 1614 743 1620 744
rect 1710 748 1716 749
rect 1710 744 1711 748
rect 1715 744 1716 748
rect 1710 743 1716 744
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 1806 743 1812 744
rect 1902 748 1908 749
rect 1902 744 1903 748
rect 1907 744 1908 748
rect 1902 743 1908 744
rect 1998 748 2004 749
rect 1998 744 1999 748
rect 2003 744 2004 748
rect 1998 743 2004 744
rect 2070 748 2076 749
rect 2070 744 2071 748
rect 2075 744 2076 748
rect 2120 746 2122 749
rect 2070 743 2076 744
rect 2118 745 2124 746
rect 110 740 116 741
rect 110 736 111 740
rect 115 736 116 740
rect 110 735 116 736
rect 1094 740 1100 741
rect 1134 740 1140 741
rect 2118 741 2119 745
rect 2123 741 2124 745
rect 2118 740 2124 741
rect 1094 736 1095 740
rect 1099 736 1100 740
rect 1094 735 1100 736
rect 112 711 114 735
rect 134 732 140 733
rect 134 728 135 732
rect 139 728 140 732
rect 134 727 140 728
rect 206 732 212 733
rect 206 728 207 732
rect 211 728 212 732
rect 206 727 212 728
rect 294 732 300 733
rect 294 728 295 732
rect 299 728 300 732
rect 294 727 300 728
rect 374 732 380 733
rect 374 728 375 732
rect 379 728 380 732
rect 374 727 380 728
rect 446 732 452 733
rect 446 728 447 732
rect 451 728 452 732
rect 446 727 452 728
rect 518 732 524 733
rect 518 728 519 732
rect 523 728 524 732
rect 518 727 524 728
rect 582 732 588 733
rect 582 728 583 732
rect 587 728 588 732
rect 582 727 588 728
rect 638 732 644 733
rect 638 728 639 732
rect 643 728 644 732
rect 638 727 644 728
rect 686 732 692 733
rect 686 728 687 732
rect 691 728 692 732
rect 686 727 692 728
rect 742 732 748 733
rect 742 728 743 732
rect 747 728 748 732
rect 742 727 748 728
rect 798 732 804 733
rect 798 728 799 732
rect 803 728 804 732
rect 798 727 804 728
rect 854 732 860 733
rect 854 728 855 732
rect 859 728 860 732
rect 854 727 860 728
rect 136 711 138 727
rect 208 711 210 727
rect 296 711 298 727
rect 376 711 378 727
rect 448 711 450 727
rect 520 711 522 727
rect 584 711 586 727
rect 640 711 642 727
rect 688 711 690 727
rect 744 711 746 727
rect 800 711 802 727
rect 856 711 858 727
rect 1096 711 1098 735
rect 1134 728 1140 729
rect 1134 724 1135 728
rect 1139 724 1140 728
rect 1134 723 1140 724
rect 2118 728 2124 729
rect 2118 724 2119 728
rect 2123 724 2124 728
rect 2118 723 2124 724
rect 111 710 115 711
rect 111 705 115 706
rect 135 710 139 711
rect 135 705 139 706
rect 183 710 187 711
rect 183 705 187 706
rect 207 710 211 711
rect 207 705 211 706
rect 247 710 251 711
rect 247 705 251 706
rect 295 710 299 711
rect 295 705 299 706
rect 311 710 315 711
rect 311 705 315 706
rect 375 710 379 711
rect 375 705 379 706
rect 383 710 387 711
rect 383 705 387 706
rect 447 710 451 711
rect 447 705 451 706
rect 455 710 459 711
rect 455 705 459 706
rect 519 710 523 711
rect 519 705 523 706
rect 583 710 587 711
rect 583 705 587 706
rect 639 710 643 711
rect 639 705 643 706
rect 647 710 651 711
rect 647 705 651 706
rect 687 710 691 711
rect 687 705 691 706
rect 711 710 715 711
rect 711 705 715 706
rect 743 710 747 711
rect 743 705 747 706
rect 767 710 771 711
rect 767 705 771 706
rect 799 710 803 711
rect 799 705 803 706
rect 823 710 827 711
rect 823 705 827 706
rect 855 710 859 711
rect 855 705 859 706
rect 879 710 883 711
rect 879 705 883 706
rect 943 710 947 711
rect 943 705 947 706
rect 1095 710 1099 711
rect 1095 705 1099 706
rect 112 685 114 705
rect 136 693 138 705
rect 184 693 186 705
rect 248 693 250 705
rect 312 693 314 705
rect 384 693 386 705
rect 456 693 458 705
rect 520 693 522 705
rect 584 693 586 705
rect 648 693 650 705
rect 712 693 714 705
rect 768 693 770 705
rect 824 693 826 705
rect 880 693 882 705
rect 944 693 946 705
rect 134 692 140 693
rect 134 688 135 692
rect 139 688 140 692
rect 134 687 140 688
rect 182 692 188 693
rect 182 688 183 692
rect 187 688 188 692
rect 182 687 188 688
rect 246 692 252 693
rect 246 688 247 692
rect 251 688 252 692
rect 246 687 252 688
rect 310 692 316 693
rect 310 688 311 692
rect 315 688 316 692
rect 310 687 316 688
rect 382 692 388 693
rect 382 688 383 692
rect 387 688 388 692
rect 382 687 388 688
rect 454 692 460 693
rect 454 688 455 692
rect 459 688 460 692
rect 454 687 460 688
rect 518 692 524 693
rect 518 688 519 692
rect 523 688 524 692
rect 518 687 524 688
rect 582 692 588 693
rect 582 688 583 692
rect 587 688 588 692
rect 582 687 588 688
rect 646 692 652 693
rect 646 688 647 692
rect 651 688 652 692
rect 646 687 652 688
rect 710 692 716 693
rect 710 688 711 692
rect 715 688 716 692
rect 710 687 716 688
rect 766 692 772 693
rect 766 688 767 692
rect 771 688 772 692
rect 766 687 772 688
rect 822 692 828 693
rect 822 688 823 692
rect 827 688 828 692
rect 822 687 828 688
rect 878 692 884 693
rect 878 688 879 692
rect 883 688 884 692
rect 878 687 884 688
rect 942 692 948 693
rect 942 688 943 692
rect 947 688 948 692
rect 942 687 948 688
rect 1096 685 1098 705
rect 1136 699 1138 723
rect 1158 720 1164 721
rect 1158 716 1159 720
rect 1163 716 1164 720
rect 1158 715 1164 716
rect 1198 720 1204 721
rect 1198 716 1199 720
rect 1203 716 1204 720
rect 1198 715 1204 716
rect 1238 720 1244 721
rect 1238 716 1239 720
rect 1243 716 1244 720
rect 1238 715 1244 716
rect 1286 720 1292 721
rect 1286 716 1287 720
rect 1291 716 1292 720
rect 1286 715 1292 716
rect 1358 720 1364 721
rect 1358 716 1359 720
rect 1363 716 1364 720
rect 1358 715 1364 716
rect 1438 720 1444 721
rect 1438 716 1439 720
rect 1443 716 1444 720
rect 1438 715 1444 716
rect 1526 720 1532 721
rect 1526 716 1527 720
rect 1531 716 1532 720
rect 1526 715 1532 716
rect 1614 720 1620 721
rect 1614 716 1615 720
rect 1619 716 1620 720
rect 1614 715 1620 716
rect 1710 720 1716 721
rect 1710 716 1711 720
rect 1715 716 1716 720
rect 1710 715 1716 716
rect 1806 720 1812 721
rect 1806 716 1807 720
rect 1811 716 1812 720
rect 1806 715 1812 716
rect 1902 720 1908 721
rect 1902 716 1903 720
rect 1907 716 1908 720
rect 1902 715 1908 716
rect 1998 720 2004 721
rect 1998 716 1999 720
rect 2003 716 2004 720
rect 1998 715 2004 716
rect 2070 720 2076 721
rect 2070 716 2071 720
rect 2075 716 2076 720
rect 2070 715 2076 716
rect 1160 699 1162 715
rect 1200 699 1202 715
rect 1240 699 1242 715
rect 1288 699 1290 715
rect 1360 699 1362 715
rect 1440 699 1442 715
rect 1528 699 1530 715
rect 1616 699 1618 715
rect 1712 699 1714 715
rect 1808 699 1810 715
rect 1904 699 1906 715
rect 2000 699 2002 715
rect 2072 699 2074 715
rect 2120 699 2122 723
rect 1135 698 1139 699
rect 1135 693 1139 694
rect 1159 698 1163 699
rect 1159 693 1163 694
rect 1199 698 1203 699
rect 1199 693 1203 694
rect 1239 698 1243 699
rect 1239 693 1243 694
rect 1287 698 1291 699
rect 1287 693 1291 694
rect 1335 698 1339 699
rect 1335 693 1339 694
rect 1359 698 1363 699
rect 1359 693 1363 694
rect 1391 698 1395 699
rect 1391 693 1395 694
rect 1439 698 1443 699
rect 1439 693 1443 694
rect 1447 698 1451 699
rect 1447 693 1451 694
rect 1511 698 1515 699
rect 1511 693 1515 694
rect 1527 698 1531 699
rect 1527 693 1531 694
rect 1575 698 1579 699
rect 1575 693 1579 694
rect 1615 698 1619 699
rect 1615 693 1619 694
rect 1639 698 1643 699
rect 1639 693 1643 694
rect 1703 698 1707 699
rect 1703 693 1707 694
rect 1711 698 1715 699
rect 1711 693 1715 694
rect 1767 698 1771 699
rect 1767 693 1771 694
rect 1807 698 1811 699
rect 1807 693 1811 694
rect 1831 698 1835 699
rect 1831 693 1835 694
rect 1895 698 1899 699
rect 1895 693 1899 694
rect 1903 698 1907 699
rect 1903 693 1907 694
rect 1959 698 1963 699
rect 1959 693 1963 694
rect 1999 698 2003 699
rect 1999 693 2003 694
rect 2023 698 2027 699
rect 2023 693 2027 694
rect 2071 698 2075 699
rect 2071 693 2075 694
rect 2119 698 2123 699
rect 2119 693 2123 694
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 110 679 116 680
rect 1094 684 1100 685
rect 1094 680 1095 684
rect 1099 680 1100 684
rect 1094 679 1100 680
rect 1136 673 1138 693
rect 1240 681 1242 693
rect 1288 681 1290 693
rect 1336 681 1338 693
rect 1392 681 1394 693
rect 1448 681 1450 693
rect 1512 681 1514 693
rect 1576 681 1578 693
rect 1640 681 1642 693
rect 1704 681 1706 693
rect 1768 681 1770 693
rect 1832 681 1834 693
rect 1896 681 1898 693
rect 1960 681 1962 693
rect 2024 681 2026 693
rect 2072 681 2074 693
rect 1238 680 1244 681
rect 1238 676 1239 680
rect 1243 676 1244 680
rect 1238 675 1244 676
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 1334 680 1340 681
rect 1334 676 1335 680
rect 1339 676 1340 680
rect 1334 675 1340 676
rect 1390 680 1396 681
rect 1390 676 1391 680
rect 1395 676 1396 680
rect 1390 675 1396 676
rect 1446 680 1452 681
rect 1446 676 1447 680
rect 1451 676 1452 680
rect 1446 675 1452 676
rect 1510 680 1516 681
rect 1510 676 1511 680
rect 1515 676 1516 680
rect 1510 675 1516 676
rect 1574 680 1580 681
rect 1574 676 1575 680
rect 1579 676 1580 680
rect 1574 675 1580 676
rect 1638 680 1644 681
rect 1638 676 1639 680
rect 1643 676 1644 680
rect 1638 675 1644 676
rect 1702 680 1708 681
rect 1702 676 1703 680
rect 1707 676 1708 680
rect 1702 675 1708 676
rect 1766 680 1772 681
rect 1766 676 1767 680
rect 1771 676 1772 680
rect 1766 675 1772 676
rect 1830 680 1836 681
rect 1830 676 1831 680
rect 1835 676 1836 680
rect 1830 675 1836 676
rect 1894 680 1900 681
rect 1894 676 1895 680
rect 1899 676 1900 680
rect 1894 675 1900 676
rect 1958 680 1964 681
rect 1958 676 1959 680
rect 1963 676 1964 680
rect 1958 675 1964 676
rect 2022 680 2028 681
rect 2022 676 2023 680
rect 2027 676 2028 680
rect 2022 675 2028 676
rect 2070 680 2076 681
rect 2070 676 2071 680
rect 2075 676 2076 680
rect 2070 675 2076 676
rect 2120 673 2122 693
rect 1134 672 1140 673
rect 1134 668 1135 672
rect 1139 668 1140 672
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 1094 667 1100 668
rect 1134 667 1140 668
rect 2118 672 2124 673
rect 2118 668 2119 672
rect 2123 668 2124 672
rect 2118 667 2124 668
rect 110 662 116 663
rect 134 664 140 665
rect 112 651 114 662
rect 134 660 135 664
rect 139 660 140 664
rect 134 659 140 660
rect 182 664 188 665
rect 182 660 183 664
rect 187 660 188 664
rect 182 659 188 660
rect 246 664 252 665
rect 246 660 247 664
rect 251 660 252 664
rect 246 659 252 660
rect 310 664 316 665
rect 310 660 311 664
rect 315 660 316 664
rect 310 659 316 660
rect 382 664 388 665
rect 382 660 383 664
rect 387 660 388 664
rect 382 659 388 660
rect 454 664 460 665
rect 454 660 455 664
rect 459 660 460 664
rect 454 659 460 660
rect 518 664 524 665
rect 518 660 519 664
rect 523 660 524 664
rect 518 659 524 660
rect 582 664 588 665
rect 582 660 583 664
rect 587 660 588 664
rect 582 659 588 660
rect 646 664 652 665
rect 646 660 647 664
rect 651 660 652 664
rect 646 659 652 660
rect 710 664 716 665
rect 710 660 711 664
rect 715 660 716 664
rect 710 659 716 660
rect 766 664 772 665
rect 766 660 767 664
rect 771 660 772 664
rect 766 659 772 660
rect 822 664 828 665
rect 822 660 823 664
rect 827 660 828 664
rect 822 659 828 660
rect 878 664 884 665
rect 878 660 879 664
rect 883 660 884 664
rect 878 659 884 660
rect 942 664 948 665
rect 942 660 943 664
rect 947 660 948 664
rect 1094 663 1095 667
rect 1099 663 1100 667
rect 1094 662 1100 663
rect 942 659 948 660
rect 136 651 138 659
rect 184 651 186 659
rect 248 651 250 659
rect 312 651 314 659
rect 384 651 386 659
rect 456 651 458 659
rect 520 651 522 659
rect 584 651 586 659
rect 648 651 650 659
rect 712 651 714 659
rect 768 651 770 659
rect 824 651 826 659
rect 880 651 882 659
rect 944 651 946 659
rect 1096 651 1098 662
rect 1134 655 1140 656
rect 1134 651 1135 655
rect 1139 651 1140 655
rect 2118 655 2124 656
rect 111 650 115 651
rect 111 645 115 646
rect 135 650 139 651
rect 135 645 139 646
rect 159 650 163 651
rect 159 645 163 646
rect 183 650 187 651
rect 183 645 187 646
rect 215 650 219 651
rect 215 645 219 646
rect 247 650 251 651
rect 247 645 251 646
rect 287 650 291 651
rect 287 645 291 646
rect 311 650 315 651
rect 311 645 315 646
rect 367 650 371 651
rect 367 645 371 646
rect 383 650 387 651
rect 383 645 387 646
rect 455 650 459 651
rect 455 645 459 646
rect 519 650 523 651
rect 519 645 523 646
rect 543 650 547 651
rect 543 645 547 646
rect 583 650 587 651
rect 583 645 587 646
rect 631 650 635 651
rect 631 645 635 646
rect 647 650 651 651
rect 647 645 651 646
rect 711 650 715 651
rect 711 645 715 646
rect 719 650 723 651
rect 719 645 723 646
rect 767 650 771 651
rect 767 645 771 646
rect 799 650 803 651
rect 799 645 803 646
rect 823 650 827 651
rect 823 645 827 646
rect 871 650 875 651
rect 871 645 875 646
rect 879 650 883 651
rect 879 645 883 646
rect 943 650 947 651
rect 943 645 947 646
rect 951 650 955 651
rect 951 645 955 646
rect 1031 650 1035 651
rect 1031 645 1035 646
rect 1095 650 1099 651
rect 1134 650 1140 651
rect 1238 652 1244 653
rect 1136 647 1138 650
rect 1238 648 1239 652
rect 1243 648 1244 652
rect 1238 647 1244 648
rect 1286 652 1292 653
rect 1286 648 1287 652
rect 1291 648 1292 652
rect 1286 647 1292 648
rect 1334 652 1340 653
rect 1334 648 1335 652
rect 1339 648 1340 652
rect 1334 647 1340 648
rect 1390 652 1396 653
rect 1390 648 1391 652
rect 1395 648 1396 652
rect 1390 647 1396 648
rect 1446 652 1452 653
rect 1446 648 1447 652
rect 1451 648 1452 652
rect 1446 647 1452 648
rect 1510 652 1516 653
rect 1510 648 1511 652
rect 1515 648 1516 652
rect 1510 647 1516 648
rect 1574 652 1580 653
rect 1574 648 1575 652
rect 1579 648 1580 652
rect 1574 647 1580 648
rect 1638 652 1644 653
rect 1638 648 1639 652
rect 1643 648 1644 652
rect 1638 647 1644 648
rect 1702 652 1708 653
rect 1702 648 1703 652
rect 1707 648 1708 652
rect 1702 647 1708 648
rect 1766 652 1772 653
rect 1766 648 1767 652
rect 1771 648 1772 652
rect 1766 647 1772 648
rect 1830 652 1836 653
rect 1830 648 1831 652
rect 1835 648 1836 652
rect 1830 647 1836 648
rect 1894 652 1900 653
rect 1894 648 1895 652
rect 1899 648 1900 652
rect 1894 647 1900 648
rect 1958 652 1964 653
rect 1958 648 1959 652
rect 1963 648 1964 652
rect 1958 647 1964 648
rect 2022 652 2028 653
rect 2022 648 2023 652
rect 2027 648 2028 652
rect 2022 647 2028 648
rect 2070 652 2076 653
rect 2070 648 2071 652
rect 2075 648 2076 652
rect 2118 651 2119 655
rect 2123 651 2124 655
rect 2118 650 2124 651
rect 2070 647 2076 648
rect 2120 647 2122 650
rect 1095 645 1099 646
rect 1135 646 1139 647
rect 112 642 114 645
rect 158 644 164 645
rect 110 641 116 642
rect 110 637 111 641
rect 115 637 116 641
rect 158 640 159 644
rect 163 640 164 644
rect 158 639 164 640
rect 214 644 220 645
rect 214 640 215 644
rect 219 640 220 644
rect 214 639 220 640
rect 286 644 292 645
rect 286 640 287 644
rect 291 640 292 644
rect 286 639 292 640
rect 366 644 372 645
rect 366 640 367 644
rect 371 640 372 644
rect 366 639 372 640
rect 454 644 460 645
rect 454 640 455 644
rect 459 640 460 644
rect 454 639 460 640
rect 542 644 548 645
rect 542 640 543 644
rect 547 640 548 644
rect 542 639 548 640
rect 630 644 636 645
rect 630 640 631 644
rect 635 640 636 644
rect 630 639 636 640
rect 718 644 724 645
rect 718 640 719 644
rect 723 640 724 644
rect 718 639 724 640
rect 798 644 804 645
rect 798 640 799 644
rect 803 640 804 644
rect 798 639 804 640
rect 870 644 876 645
rect 870 640 871 644
rect 875 640 876 644
rect 870 639 876 640
rect 950 644 956 645
rect 950 640 951 644
rect 955 640 956 644
rect 950 639 956 640
rect 1030 644 1036 645
rect 1030 640 1031 644
rect 1035 640 1036 644
rect 1096 642 1098 645
rect 1030 639 1036 640
rect 1094 641 1100 642
rect 1135 641 1139 642
rect 1239 646 1243 647
rect 1239 641 1243 642
rect 1279 646 1283 647
rect 1279 641 1283 642
rect 1287 646 1291 647
rect 1287 641 1291 642
rect 1319 646 1323 647
rect 1319 641 1323 642
rect 1335 646 1339 647
rect 1335 641 1339 642
rect 1367 646 1371 647
rect 1367 641 1371 642
rect 1391 646 1395 647
rect 1391 641 1395 642
rect 1423 646 1427 647
rect 1423 641 1427 642
rect 1447 646 1451 647
rect 1447 641 1451 642
rect 1479 646 1483 647
rect 1479 641 1483 642
rect 1511 646 1515 647
rect 1511 641 1515 642
rect 1535 646 1539 647
rect 1535 641 1539 642
rect 1575 646 1579 647
rect 1575 641 1579 642
rect 1591 646 1595 647
rect 1591 641 1595 642
rect 1639 646 1643 647
rect 1639 641 1643 642
rect 1647 646 1651 647
rect 1647 641 1651 642
rect 1703 646 1707 647
rect 1703 641 1707 642
rect 1719 646 1723 647
rect 1719 641 1723 642
rect 1767 646 1771 647
rect 1767 641 1771 642
rect 1799 646 1803 647
rect 1799 641 1803 642
rect 1831 646 1835 647
rect 1831 641 1835 642
rect 1879 646 1883 647
rect 1879 641 1883 642
rect 1895 646 1899 647
rect 1895 641 1899 642
rect 1959 646 1963 647
rect 1959 641 1963 642
rect 1967 646 1971 647
rect 1967 641 1971 642
rect 2023 646 2027 647
rect 2023 641 2027 642
rect 2063 646 2067 647
rect 2063 641 2067 642
rect 2071 646 2075 647
rect 2071 641 2075 642
rect 2119 646 2123 647
rect 2119 641 2123 642
rect 110 636 116 637
rect 1094 637 1095 641
rect 1099 637 1100 641
rect 1136 638 1138 641
rect 1278 640 1284 641
rect 1094 636 1100 637
rect 1134 637 1140 638
rect 1134 633 1135 637
rect 1139 633 1140 637
rect 1278 636 1279 640
rect 1283 636 1284 640
rect 1278 635 1284 636
rect 1318 640 1324 641
rect 1318 636 1319 640
rect 1323 636 1324 640
rect 1318 635 1324 636
rect 1366 640 1372 641
rect 1366 636 1367 640
rect 1371 636 1372 640
rect 1366 635 1372 636
rect 1422 640 1428 641
rect 1422 636 1423 640
rect 1427 636 1428 640
rect 1422 635 1428 636
rect 1478 640 1484 641
rect 1478 636 1479 640
rect 1483 636 1484 640
rect 1478 635 1484 636
rect 1534 640 1540 641
rect 1534 636 1535 640
rect 1539 636 1540 640
rect 1534 635 1540 636
rect 1590 640 1596 641
rect 1590 636 1591 640
rect 1595 636 1596 640
rect 1590 635 1596 636
rect 1646 640 1652 641
rect 1646 636 1647 640
rect 1651 636 1652 640
rect 1646 635 1652 636
rect 1718 640 1724 641
rect 1718 636 1719 640
rect 1723 636 1724 640
rect 1718 635 1724 636
rect 1798 640 1804 641
rect 1798 636 1799 640
rect 1803 636 1804 640
rect 1798 635 1804 636
rect 1878 640 1884 641
rect 1878 636 1879 640
rect 1883 636 1884 640
rect 1878 635 1884 636
rect 1966 640 1972 641
rect 1966 636 1967 640
rect 1971 636 1972 640
rect 1966 635 1972 636
rect 2062 640 2068 641
rect 2062 636 2063 640
rect 2067 636 2068 640
rect 2120 638 2122 641
rect 2062 635 2068 636
rect 2118 637 2124 638
rect 1134 632 1140 633
rect 2118 633 2119 637
rect 2123 633 2124 637
rect 2118 632 2124 633
rect 110 624 116 625
rect 110 620 111 624
rect 115 620 116 624
rect 110 619 116 620
rect 1094 624 1100 625
rect 1094 620 1095 624
rect 1099 620 1100 624
rect 1094 619 1100 620
rect 1134 620 1140 621
rect 112 595 114 619
rect 158 616 164 617
rect 158 612 159 616
rect 163 612 164 616
rect 158 611 164 612
rect 214 616 220 617
rect 214 612 215 616
rect 219 612 220 616
rect 214 611 220 612
rect 286 616 292 617
rect 286 612 287 616
rect 291 612 292 616
rect 286 611 292 612
rect 366 616 372 617
rect 366 612 367 616
rect 371 612 372 616
rect 366 611 372 612
rect 454 616 460 617
rect 454 612 455 616
rect 459 612 460 616
rect 454 611 460 612
rect 542 616 548 617
rect 542 612 543 616
rect 547 612 548 616
rect 542 611 548 612
rect 630 616 636 617
rect 630 612 631 616
rect 635 612 636 616
rect 630 611 636 612
rect 718 616 724 617
rect 718 612 719 616
rect 723 612 724 616
rect 718 611 724 612
rect 798 616 804 617
rect 798 612 799 616
rect 803 612 804 616
rect 798 611 804 612
rect 870 616 876 617
rect 870 612 871 616
rect 875 612 876 616
rect 870 611 876 612
rect 950 616 956 617
rect 950 612 951 616
rect 955 612 956 616
rect 950 611 956 612
rect 1030 616 1036 617
rect 1030 612 1031 616
rect 1035 612 1036 616
rect 1030 611 1036 612
rect 160 595 162 611
rect 216 595 218 611
rect 288 595 290 611
rect 368 595 370 611
rect 456 595 458 611
rect 544 595 546 611
rect 632 595 634 611
rect 720 595 722 611
rect 800 595 802 611
rect 872 595 874 611
rect 952 595 954 611
rect 1032 595 1034 611
rect 1096 595 1098 619
rect 1134 616 1135 620
rect 1139 616 1140 620
rect 1134 615 1140 616
rect 2118 620 2124 621
rect 2118 616 2119 620
rect 2123 616 2124 620
rect 2118 615 2124 616
rect 1136 595 1138 615
rect 1278 612 1284 613
rect 1278 608 1279 612
rect 1283 608 1284 612
rect 1278 607 1284 608
rect 1318 612 1324 613
rect 1318 608 1319 612
rect 1323 608 1324 612
rect 1318 607 1324 608
rect 1366 612 1372 613
rect 1366 608 1367 612
rect 1371 608 1372 612
rect 1366 607 1372 608
rect 1422 612 1428 613
rect 1422 608 1423 612
rect 1427 608 1428 612
rect 1422 607 1428 608
rect 1478 612 1484 613
rect 1478 608 1479 612
rect 1483 608 1484 612
rect 1478 607 1484 608
rect 1534 612 1540 613
rect 1534 608 1535 612
rect 1539 608 1540 612
rect 1534 607 1540 608
rect 1590 612 1596 613
rect 1590 608 1591 612
rect 1595 608 1596 612
rect 1590 607 1596 608
rect 1646 612 1652 613
rect 1646 608 1647 612
rect 1651 608 1652 612
rect 1646 607 1652 608
rect 1718 612 1724 613
rect 1718 608 1719 612
rect 1723 608 1724 612
rect 1718 607 1724 608
rect 1798 612 1804 613
rect 1798 608 1799 612
rect 1803 608 1804 612
rect 1798 607 1804 608
rect 1878 612 1884 613
rect 1878 608 1879 612
rect 1883 608 1884 612
rect 1878 607 1884 608
rect 1966 612 1972 613
rect 1966 608 1967 612
rect 1971 608 1972 612
rect 1966 607 1972 608
rect 2062 612 2068 613
rect 2062 608 2063 612
rect 2067 608 2068 612
rect 2062 607 2068 608
rect 1280 595 1282 607
rect 1320 595 1322 607
rect 1368 595 1370 607
rect 1424 595 1426 607
rect 1480 595 1482 607
rect 1536 595 1538 607
rect 1592 595 1594 607
rect 1648 595 1650 607
rect 1720 595 1722 607
rect 1800 595 1802 607
rect 1880 595 1882 607
rect 1968 595 1970 607
rect 2064 595 2066 607
rect 2120 595 2122 615
rect 111 594 115 595
rect 111 589 115 590
rect 159 594 163 595
rect 159 589 163 590
rect 207 594 211 595
rect 207 589 211 590
rect 215 594 219 595
rect 215 589 219 590
rect 255 594 259 595
rect 255 589 259 590
rect 287 594 291 595
rect 287 589 291 590
rect 311 594 315 595
rect 311 589 315 590
rect 367 594 371 595
rect 367 589 371 590
rect 383 594 387 595
rect 383 589 387 590
rect 455 594 459 595
rect 455 589 459 590
rect 463 594 467 595
rect 463 589 467 590
rect 543 594 547 595
rect 543 589 547 590
rect 623 594 627 595
rect 623 589 627 590
rect 631 594 635 595
rect 631 589 635 590
rect 703 594 707 595
rect 703 589 707 590
rect 719 594 723 595
rect 719 589 723 590
rect 783 594 787 595
rect 783 589 787 590
rect 799 594 803 595
rect 799 589 803 590
rect 855 594 859 595
rect 855 589 859 590
rect 871 594 875 595
rect 871 589 875 590
rect 927 594 931 595
rect 927 589 931 590
rect 951 594 955 595
rect 951 589 955 590
rect 999 594 1003 595
rect 999 589 1003 590
rect 1031 594 1035 595
rect 1031 589 1035 590
rect 1047 594 1051 595
rect 1047 589 1051 590
rect 1095 594 1099 595
rect 1095 589 1099 590
rect 1135 594 1139 595
rect 1135 589 1139 590
rect 1279 594 1283 595
rect 1279 589 1283 590
rect 1319 594 1323 595
rect 1319 589 1323 590
rect 1335 594 1339 595
rect 1335 589 1339 590
rect 1367 594 1371 595
rect 1367 589 1371 590
rect 1375 594 1379 595
rect 1375 589 1379 590
rect 1415 594 1419 595
rect 1415 589 1419 590
rect 1423 594 1427 595
rect 1423 589 1427 590
rect 1463 594 1467 595
rect 1463 589 1467 590
rect 1479 594 1483 595
rect 1479 589 1483 590
rect 1519 594 1523 595
rect 1519 589 1523 590
rect 1535 594 1539 595
rect 1535 589 1539 590
rect 1583 594 1587 595
rect 1583 589 1587 590
rect 1591 594 1595 595
rect 1591 589 1595 590
rect 1647 594 1651 595
rect 1647 589 1651 590
rect 1655 594 1659 595
rect 1655 589 1659 590
rect 1719 594 1723 595
rect 1719 589 1723 590
rect 1727 594 1731 595
rect 1727 589 1731 590
rect 1799 594 1803 595
rect 1799 589 1803 590
rect 1807 594 1811 595
rect 1807 589 1811 590
rect 1879 594 1883 595
rect 1879 589 1883 590
rect 1887 594 1891 595
rect 1887 589 1891 590
rect 1967 594 1971 595
rect 1967 589 1971 590
rect 1975 594 1979 595
rect 1975 589 1979 590
rect 2063 594 2067 595
rect 2063 589 2067 590
rect 2119 594 2123 595
rect 2119 589 2123 590
rect 112 569 114 589
rect 160 577 162 589
rect 208 577 210 589
rect 256 577 258 589
rect 312 577 314 589
rect 384 577 386 589
rect 464 577 466 589
rect 544 577 546 589
rect 624 577 626 589
rect 704 577 706 589
rect 784 577 786 589
rect 856 577 858 589
rect 928 577 930 589
rect 1000 577 1002 589
rect 1048 577 1050 589
rect 158 576 164 577
rect 158 572 159 576
rect 163 572 164 576
rect 158 571 164 572
rect 206 576 212 577
rect 206 572 207 576
rect 211 572 212 576
rect 206 571 212 572
rect 254 576 260 577
rect 254 572 255 576
rect 259 572 260 576
rect 254 571 260 572
rect 310 576 316 577
rect 310 572 311 576
rect 315 572 316 576
rect 310 571 316 572
rect 382 576 388 577
rect 382 572 383 576
rect 387 572 388 576
rect 382 571 388 572
rect 462 576 468 577
rect 462 572 463 576
rect 467 572 468 576
rect 462 571 468 572
rect 542 576 548 577
rect 542 572 543 576
rect 547 572 548 576
rect 542 571 548 572
rect 622 576 628 577
rect 622 572 623 576
rect 627 572 628 576
rect 622 571 628 572
rect 702 576 708 577
rect 702 572 703 576
rect 707 572 708 576
rect 702 571 708 572
rect 782 576 788 577
rect 782 572 783 576
rect 787 572 788 576
rect 782 571 788 572
rect 854 576 860 577
rect 854 572 855 576
rect 859 572 860 576
rect 854 571 860 572
rect 926 576 932 577
rect 926 572 927 576
rect 931 572 932 576
rect 926 571 932 572
rect 998 576 1004 577
rect 998 572 999 576
rect 1003 572 1004 576
rect 998 571 1004 572
rect 1046 576 1052 577
rect 1046 572 1047 576
rect 1051 572 1052 576
rect 1046 571 1052 572
rect 1096 569 1098 589
rect 1136 569 1138 589
rect 1336 577 1338 589
rect 1376 577 1378 589
rect 1416 577 1418 589
rect 1464 577 1466 589
rect 1520 577 1522 589
rect 1584 577 1586 589
rect 1656 577 1658 589
rect 1728 577 1730 589
rect 1808 577 1810 589
rect 1888 577 1890 589
rect 1976 577 1978 589
rect 2064 577 2066 589
rect 1334 576 1340 577
rect 1334 572 1335 576
rect 1339 572 1340 576
rect 1334 571 1340 572
rect 1374 576 1380 577
rect 1374 572 1375 576
rect 1379 572 1380 576
rect 1374 571 1380 572
rect 1414 576 1420 577
rect 1414 572 1415 576
rect 1419 572 1420 576
rect 1414 571 1420 572
rect 1462 576 1468 577
rect 1462 572 1463 576
rect 1467 572 1468 576
rect 1462 571 1468 572
rect 1518 576 1524 577
rect 1518 572 1519 576
rect 1523 572 1524 576
rect 1518 571 1524 572
rect 1582 576 1588 577
rect 1582 572 1583 576
rect 1587 572 1588 576
rect 1582 571 1588 572
rect 1654 576 1660 577
rect 1654 572 1655 576
rect 1659 572 1660 576
rect 1654 571 1660 572
rect 1726 576 1732 577
rect 1726 572 1727 576
rect 1731 572 1732 576
rect 1726 571 1732 572
rect 1806 576 1812 577
rect 1806 572 1807 576
rect 1811 572 1812 576
rect 1806 571 1812 572
rect 1886 576 1892 577
rect 1886 572 1887 576
rect 1891 572 1892 576
rect 1886 571 1892 572
rect 1974 576 1980 577
rect 1974 572 1975 576
rect 1979 572 1980 576
rect 1974 571 1980 572
rect 2062 576 2068 577
rect 2062 572 2063 576
rect 2067 572 2068 576
rect 2062 571 2068 572
rect 2120 569 2122 589
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 110 563 116 564
rect 1094 568 1100 569
rect 1094 564 1095 568
rect 1099 564 1100 568
rect 1094 563 1100 564
rect 1134 568 1140 569
rect 1134 564 1135 568
rect 1139 564 1140 568
rect 1134 563 1140 564
rect 2118 568 2124 569
rect 2118 564 2119 568
rect 2123 564 2124 568
rect 2118 563 2124 564
rect 110 551 116 552
rect 110 547 111 551
rect 115 547 116 551
rect 1094 551 1100 552
rect 110 546 116 547
rect 158 548 164 549
rect 112 535 114 546
rect 158 544 159 548
rect 163 544 164 548
rect 158 543 164 544
rect 206 548 212 549
rect 206 544 207 548
rect 211 544 212 548
rect 206 543 212 544
rect 254 548 260 549
rect 254 544 255 548
rect 259 544 260 548
rect 254 543 260 544
rect 310 548 316 549
rect 310 544 311 548
rect 315 544 316 548
rect 310 543 316 544
rect 382 548 388 549
rect 382 544 383 548
rect 387 544 388 548
rect 382 543 388 544
rect 462 548 468 549
rect 462 544 463 548
rect 467 544 468 548
rect 462 543 468 544
rect 542 548 548 549
rect 542 544 543 548
rect 547 544 548 548
rect 542 543 548 544
rect 622 548 628 549
rect 622 544 623 548
rect 627 544 628 548
rect 622 543 628 544
rect 702 548 708 549
rect 702 544 703 548
rect 707 544 708 548
rect 702 543 708 544
rect 782 548 788 549
rect 782 544 783 548
rect 787 544 788 548
rect 782 543 788 544
rect 854 548 860 549
rect 854 544 855 548
rect 859 544 860 548
rect 854 543 860 544
rect 926 548 932 549
rect 926 544 927 548
rect 931 544 932 548
rect 926 543 932 544
rect 998 548 1004 549
rect 998 544 999 548
rect 1003 544 1004 548
rect 998 543 1004 544
rect 1046 548 1052 549
rect 1046 544 1047 548
rect 1051 544 1052 548
rect 1094 547 1095 551
rect 1099 547 1100 551
rect 1094 546 1100 547
rect 1134 551 1140 552
rect 1134 547 1135 551
rect 1139 547 1140 551
rect 2118 551 2124 552
rect 1134 546 1140 547
rect 1334 548 1340 549
rect 1046 543 1052 544
rect 160 535 162 543
rect 208 535 210 543
rect 256 535 258 543
rect 312 535 314 543
rect 384 535 386 543
rect 464 535 466 543
rect 544 535 546 543
rect 624 535 626 543
rect 704 535 706 543
rect 784 535 786 543
rect 856 535 858 543
rect 928 535 930 543
rect 1000 535 1002 543
rect 1048 535 1050 543
rect 1096 535 1098 546
rect 1136 539 1138 546
rect 1334 544 1335 548
rect 1339 544 1340 548
rect 1334 543 1340 544
rect 1374 548 1380 549
rect 1374 544 1375 548
rect 1379 544 1380 548
rect 1374 543 1380 544
rect 1414 548 1420 549
rect 1414 544 1415 548
rect 1419 544 1420 548
rect 1414 543 1420 544
rect 1462 548 1468 549
rect 1462 544 1463 548
rect 1467 544 1468 548
rect 1462 543 1468 544
rect 1518 548 1524 549
rect 1518 544 1519 548
rect 1523 544 1524 548
rect 1518 543 1524 544
rect 1582 548 1588 549
rect 1582 544 1583 548
rect 1587 544 1588 548
rect 1582 543 1588 544
rect 1654 548 1660 549
rect 1654 544 1655 548
rect 1659 544 1660 548
rect 1654 543 1660 544
rect 1726 548 1732 549
rect 1726 544 1727 548
rect 1731 544 1732 548
rect 1726 543 1732 544
rect 1806 548 1812 549
rect 1806 544 1807 548
rect 1811 544 1812 548
rect 1806 543 1812 544
rect 1886 548 1892 549
rect 1886 544 1887 548
rect 1891 544 1892 548
rect 1886 543 1892 544
rect 1974 548 1980 549
rect 1974 544 1975 548
rect 1979 544 1980 548
rect 1974 543 1980 544
rect 2062 548 2068 549
rect 2062 544 2063 548
rect 2067 544 2068 548
rect 2118 547 2119 551
rect 2123 547 2124 551
rect 2118 546 2124 547
rect 2062 543 2068 544
rect 1336 539 1338 543
rect 1376 539 1378 543
rect 1416 539 1418 543
rect 1464 539 1466 543
rect 1520 539 1522 543
rect 1584 539 1586 543
rect 1656 539 1658 543
rect 1728 539 1730 543
rect 1808 539 1810 543
rect 1888 539 1890 543
rect 1976 539 1978 543
rect 2064 539 2066 543
rect 2120 539 2122 546
rect 1135 538 1139 539
rect 111 534 115 535
rect 111 529 115 530
rect 159 534 163 535
rect 159 529 163 530
rect 167 534 171 535
rect 167 529 171 530
rect 207 534 211 535
rect 207 529 211 530
rect 223 534 227 535
rect 223 529 227 530
rect 255 534 259 535
rect 255 529 259 530
rect 287 534 291 535
rect 287 529 291 530
rect 311 534 315 535
rect 311 529 315 530
rect 359 534 363 535
rect 359 529 363 530
rect 383 534 387 535
rect 383 529 387 530
rect 431 534 435 535
rect 431 529 435 530
rect 463 534 467 535
rect 463 529 467 530
rect 511 534 515 535
rect 511 529 515 530
rect 543 534 547 535
rect 543 529 547 530
rect 591 534 595 535
rect 591 529 595 530
rect 623 534 627 535
rect 623 529 627 530
rect 663 534 667 535
rect 663 529 667 530
rect 703 534 707 535
rect 703 529 707 530
rect 735 534 739 535
rect 735 529 739 530
rect 783 534 787 535
rect 783 529 787 530
rect 807 534 811 535
rect 807 529 811 530
rect 855 534 859 535
rect 855 529 859 530
rect 871 534 875 535
rect 871 529 875 530
rect 927 534 931 535
rect 927 529 931 530
rect 935 534 939 535
rect 935 529 939 530
rect 999 534 1003 535
rect 999 529 1003 530
rect 1047 534 1051 535
rect 1047 529 1051 530
rect 1095 534 1099 535
rect 1135 533 1139 534
rect 1191 538 1195 539
rect 1191 533 1195 534
rect 1239 538 1243 539
rect 1239 533 1243 534
rect 1287 538 1291 539
rect 1287 533 1291 534
rect 1335 538 1339 539
rect 1335 533 1339 534
rect 1343 538 1347 539
rect 1343 533 1347 534
rect 1375 538 1379 539
rect 1375 533 1379 534
rect 1407 538 1411 539
rect 1407 533 1411 534
rect 1415 538 1419 539
rect 1415 533 1419 534
rect 1463 538 1467 539
rect 1463 533 1467 534
rect 1479 538 1483 539
rect 1479 533 1483 534
rect 1519 538 1523 539
rect 1519 533 1523 534
rect 1543 538 1547 539
rect 1543 533 1547 534
rect 1583 538 1587 539
rect 1583 533 1587 534
rect 1607 538 1611 539
rect 1607 533 1611 534
rect 1655 538 1659 539
rect 1655 533 1659 534
rect 1671 538 1675 539
rect 1671 533 1675 534
rect 1727 538 1731 539
rect 1727 533 1731 534
rect 1735 538 1739 539
rect 1735 533 1739 534
rect 1799 538 1803 539
rect 1799 533 1803 534
rect 1807 538 1811 539
rect 1807 533 1811 534
rect 1863 538 1867 539
rect 1863 533 1867 534
rect 1887 538 1891 539
rect 1887 533 1891 534
rect 1935 538 1939 539
rect 1935 533 1939 534
rect 1975 538 1979 539
rect 1975 533 1979 534
rect 2007 538 2011 539
rect 2007 533 2011 534
rect 2063 538 2067 539
rect 2063 533 2067 534
rect 2071 538 2075 539
rect 2071 533 2075 534
rect 2119 538 2123 539
rect 2119 533 2123 534
rect 1136 530 1138 533
rect 1190 532 1196 533
rect 1095 529 1099 530
rect 1134 529 1140 530
rect 112 526 114 529
rect 166 528 172 529
rect 110 525 116 526
rect 110 521 111 525
rect 115 521 116 525
rect 166 524 167 528
rect 171 524 172 528
rect 166 523 172 524
rect 222 528 228 529
rect 222 524 223 528
rect 227 524 228 528
rect 222 523 228 524
rect 286 528 292 529
rect 286 524 287 528
rect 291 524 292 528
rect 286 523 292 524
rect 358 528 364 529
rect 358 524 359 528
rect 363 524 364 528
rect 358 523 364 524
rect 430 528 436 529
rect 430 524 431 528
rect 435 524 436 528
rect 430 523 436 524
rect 510 528 516 529
rect 510 524 511 528
rect 515 524 516 528
rect 510 523 516 524
rect 590 528 596 529
rect 590 524 591 528
rect 595 524 596 528
rect 590 523 596 524
rect 662 528 668 529
rect 662 524 663 528
rect 667 524 668 528
rect 662 523 668 524
rect 734 528 740 529
rect 734 524 735 528
rect 739 524 740 528
rect 734 523 740 524
rect 806 528 812 529
rect 806 524 807 528
rect 811 524 812 528
rect 806 523 812 524
rect 870 528 876 529
rect 870 524 871 528
rect 875 524 876 528
rect 870 523 876 524
rect 934 528 940 529
rect 934 524 935 528
rect 939 524 940 528
rect 934 523 940 524
rect 998 528 1004 529
rect 998 524 999 528
rect 1003 524 1004 528
rect 998 523 1004 524
rect 1046 528 1052 529
rect 1046 524 1047 528
rect 1051 524 1052 528
rect 1096 526 1098 529
rect 1046 523 1052 524
rect 1094 525 1100 526
rect 110 520 116 521
rect 1094 521 1095 525
rect 1099 521 1100 525
rect 1134 525 1135 529
rect 1139 525 1140 529
rect 1190 528 1191 532
rect 1195 528 1196 532
rect 1190 527 1196 528
rect 1238 532 1244 533
rect 1238 528 1239 532
rect 1243 528 1244 532
rect 1238 527 1244 528
rect 1286 532 1292 533
rect 1286 528 1287 532
rect 1291 528 1292 532
rect 1286 527 1292 528
rect 1342 532 1348 533
rect 1342 528 1343 532
rect 1347 528 1348 532
rect 1342 527 1348 528
rect 1406 532 1412 533
rect 1406 528 1407 532
rect 1411 528 1412 532
rect 1406 527 1412 528
rect 1478 532 1484 533
rect 1478 528 1479 532
rect 1483 528 1484 532
rect 1478 527 1484 528
rect 1542 532 1548 533
rect 1542 528 1543 532
rect 1547 528 1548 532
rect 1542 527 1548 528
rect 1606 532 1612 533
rect 1606 528 1607 532
rect 1611 528 1612 532
rect 1606 527 1612 528
rect 1670 532 1676 533
rect 1670 528 1671 532
rect 1675 528 1676 532
rect 1670 527 1676 528
rect 1734 532 1740 533
rect 1734 528 1735 532
rect 1739 528 1740 532
rect 1734 527 1740 528
rect 1798 532 1804 533
rect 1798 528 1799 532
rect 1803 528 1804 532
rect 1798 527 1804 528
rect 1862 532 1868 533
rect 1862 528 1863 532
rect 1867 528 1868 532
rect 1862 527 1868 528
rect 1934 532 1940 533
rect 1934 528 1935 532
rect 1939 528 1940 532
rect 1934 527 1940 528
rect 2006 532 2012 533
rect 2006 528 2007 532
rect 2011 528 2012 532
rect 2006 527 2012 528
rect 2070 532 2076 533
rect 2070 528 2071 532
rect 2075 528 2076 532
rect 2120 530 2122 533
rect 2070 527 2076 528
rect 2118 529 2124 530
rect 1134 524 1140 525
rect 2118 525 2119 529
rect 2123 525 2124 529
rect 2118 524 2124 525
rect 1094 520 1100 521
rect 1134 512 1140 513
rect 110 508 116 509
rect 110 504 111 508
rect 115 504 116 508
rect 110 503 116 504
rect 1094 508 1100 509
rect 1094 504 1095 508
rect 1099 504 1100 508
rect 1134 508 1135 512
rect 1139 508 1140 512
rect 1134 507 1140 508
rect 2118 512 2124 513
rect 2118 508 2119 512
rect 2123 508 2124 512
rect 2118 507 2124 508
rect 1094 503 1100 504
rect 112 483 114 503
rect 166 500 172 501
rect 166 496 167 500
rect 171 496 172 500
rect 166 495 172 496
rect 222 500 228 501
rect 222 496 223 500
rect 227 496 228 500
rect 222 495 228 496
rect 286 500 292 501
rect 286 496 287 500
rect 291 496 292 500
rect 286 495 292 496
rect 358 500 364 501
rect 358 496 359 500
rect 363 496 364 500
rect 358 495 364 496
rect 430 500 436 501
rect 430 496 431 500
rect 435 496 436 500
rect 430 495 436 496
rect 510 500 516 501
rect 510 496 511 500
rect 515 496 516 500
rect 510 495 516 496
rect 590 500 596 501
rect 590 496 591 500
rect 595 496 596 500
rect 590 495 596 496
rect 662 500 668 501
rect 662 496 663 500
rect 667 496 668 500
rect 662 495 668 496
rect 734 500 740 501
rect 734 496 735 500
rect 739 496 740 500
rect 734 495 740 496
rect 806 500 812 501
rect 806 496 807 500
rect 811 496 812 500
rect 806 495 812 496
rect 870 500 876 501
rect 870 496 871 500
rect 875 496 876 500
rect 870 495 876 496
rect 934 500 940 501
rect 934 496 935 500
rect 939 496 940 500
rect 934 495 940 496
rect 998 500 1004 501
rect 998 496 999 500
rect 1003 496 1004 500
rect 998 495 1004 496
rect 1046 500 1052 501
rect 1046 496 1047 500
rect 1051 496 1052 500
rect 1046 495 1052 496
rect 168 483 170 495
rect 224 483 226 495
rect 288 483 290 495
rect 360 483 362 495
rect 432 483 434 495
rect 512 483 514 495
rect 592 483 594 495
rect 664 483 666 495
rect 736 483 738 495
rect 808 483 810 495
rect 872 483 874 495
rect 936 483 938 495
rect 1000 483 1002 495
rect 1048 483 1050 495
rect 1096 483 1098 503
rect 1136 487 1138 507
rect 1190 504 1196 505
rect 1190 500 1191 504
rect 1195 500 1196 504
rect 1190 499 1196 500
rect 1238 504 1244 505
rect 1238 500 1239 504
rect 1243 500 1244 504
rect 1238 499 1244 500
rect 1286 504 1292 505
rect 1286 500 1287 504
rect 1291 500 1292 504
rect 1286 499 1292 500
rect 1342 504 1348 505
rect 1342 500 1343 504
rect 1347 500 1348 504
rect 1342 499 1348 500
rect 1406 504 1412 505
rect 1406 500 1407 504
rect 1411 500 1412 504
rect 1406 499 1412 500
rect 1478 504 1484 505
rect 1478 500 1479 504
rect 1483 500 1484 504
rect 1478 499 1484 500
rect 1542 504 1548 505
rect 1542 500 1543 504
rect 1547 500 1548 504
rect 1542 499 1548 500
rect 1606 504 1612 505
rect 1606 500 1607 504
rect 1611 500 1612 504
rect 1606 499 1612 500
rect 1670 504 1676 505
rect 1670 500 1671 504
rect 1675 500 1676 504
rect 1670 499 1676 500
rect 1734 504 1740 505
rect 1734 500 1735 504
rect 1739 500 1740 504
rect 1734 499 1740 500
rect 1798 504 1804 505
rect 1798 500 1799 504
rect 1803 500 1804 504
rect 1798 499 1804 500
rect 1862 504 1868 505
rect 1862 500 1863 504
rect 1867 500 1868 504
rect 1862 499 1868 500
rect 1934 504 1940 505
rect 1934 500 1935 504
rect 1939 500 1940 504
rect 1934 499 1940 500
rect 2006 504 2012 505
rect 2006 500 2007 504
rect 2011 500 2012 504
rect 2006 499 2012 500
rect 2070 504 2076 505
rect 2070 500 2071 504
rect 2075 500 2076 504
rect 2070 499 2076 500
rect 1192 487 1194 499
rect 1240 487 1242 499
rect 1288 487 1290 499
rect 1344 487 1346 499
rect 1408 487 1410 499
rect 1480 487 1482 499
rect 1544 487 1546 499
rect 1608 487 1610 499
rect 1672 487 1674 499
rect 1736 487 1738 499
rect 1800 487 1802 499
rect 1864 487 1866 499
rect 1936 487 1938 499
rect 2008 487 2010 499
rect 2072 487 2074 499
rect 2120 487 2122 507
rect 1135 486 1139 487
rect 111 482 115 483
rect 111 477 115 478
rect 167 482 171 483
rect 167 477 171 478
rect 223 482 227 483
rect 223 477 227 478
rect 231 482 235 483
rect 231 477 235 478
rect 287 482 291 483
rect 287 477 291 478
rect 303 482 307 483
rect 303 477 307 478
rect 359 482 363 483
rect 359 477 363 478
rect 375 482 379 483
rect 375 477 379 478
rect 431 482 435 483
rect 431 477 435 478
rect 455 482 459 483
rect 455 477 459 478
rect 511 482 515 483
rect 511 477 515 478
rect 535 482 539 483
rect 535 477 539 478
rect 591 482 595 483
rect 591 477 595 478
rect 607 482 611 483
rect 607 477 611 478
rect 663 482 667 483
rect 663 477 667 478
rect 679 482 683 483
rect 679 477 683 478
rect 735 482 739 483
rect 735 477 739 478
rect 743 482 747 483
rect 743 477 747 478
rect 799 482 803 483
rect 799 477 803 478
rect 807 482 811 483
rect 807 477 811 478
rect 855 482 859 483
rect 855 477 859 478
rect 871 482 875 483
rect 871 477 875 478
rect 903 482 907 483
rect 903 477 907 478
rect 935 482 939 483
rect 935 477 939 478
rect 959 482 963 483
rect 959 477 963 478
rect 999 482 1003 483
rect 999 477 1003 478
rect 1007 482 1011 483
rect 1007 477 1011 478
rect 1047 482 1051 483
rect 1047 477 1051 478
rect 1095 482 1099 483
rect 1135 481 1139 482
rect 1159 486 1163 487
rect 1159 481 1163 482
rect 1191 486 1195 487
rect 1191 481 1195 482
rect 1239 486 1243 487
rect 1239 481 1243 482
rect 1263 486 1267 487
rect 1263 481 1267 482
rect 1287 486 1291 487
rect 1287 481 1291 482
rect 1343 486 1347 487
rect 1343 481 1347 482
rect 1383 486 1387 487
rect 1383 481 1387 482
rect 1407 486 1411 487
rect 1407 481 1411 482
rect 1479 486 1483 487
rect 1479 481 1483 482
rect 1495 486 1499 487
rect 1495 481 1499 482
rect 1543 486 1547 487
rect 1543 481 1547 482
rect 1599 486 1603 487
rect 1599 481 1603 482
rect 1607 486 1611 487
rect 1607 481 1611 482
rect 1671 486 1675 487
rect 1671 481 1675 482
rect 1703 486 1707 487
rect 1703 481 1707 482
rect 1735 486 1739 487
rect 1735 481 1739 482
rect 1799 486 1803 487
rect 1799 481 1803 482
rect 1863 486 1867 487
rect 1863 481 1867 482
rect 1887 486 1891 487
rect 1887 481 1891 482
rect 1935 486 1939 487
rect 1935 481 1939 482
rect 1983 486 1987 487
rect 1983 481 1987 482
rect 2007 486 2011 487
rect 2007 481 2011 482
rect 2071 486 2075 487
rect 2071 481 2075 482
rect 2119 486 2123 487
rect 2119 481 2123 482
rect 1095 477 1099 478
rect 112 457 114 477
rect 168 465 170 477
rect 232 465 234 477
rect 304 465 306 477
rect 376 465 378 477
rect 456 465 458 477
rect 536 465 538 477
rect 608 465 610 477
rect 680 465 682 477
rect 744 465 746 477
rect 800 465 802 477
rect 856 465 858 477
rect 904 465 906 477
rect 960 465 962 477
rect 1008 465 1010 477
rect 1048 465 1050 477
rect 166 464 172 465
rect 166 460 167 464
rect 171 460 172 464
rect 166 459 172 460
rect 230 464 236 465
rect 230 460 231 464
rect 235 460 236 464
rect 230 459 236 460
rect 302 464 308 465
rect 302 460 303 464
rect 307 460 308 464
rect 302 459 308 460
rect 374 464 380 465
rect 374 460 375 464
rect 379 460 380 464
rect 374 459 380 460
rect 454 464 460 465
rect 454 460 455 464
rect 459 460 460 464
rect 454 459 460 460
rect 534 464 540 465
rect 534 460 535 464
rect 539 460 540 464
rect 534 459 540 460
rect 606 464 612 465
rect 606 460 607 464
rect 611 460 612 464
rect 606 459 612 460
rect 678 464 684 465
rect 678 460 679 464
rect 683 460 684 464
rect 678 459 684 460
rect 742 464 748 465
rect 742 460 743 464
rect 747 460 748 464
rect 742 459 748 460
rect 798 464 804 465
rect 798 460 799 464
rect 803 460 804 464
rect 798 459 804 460
rect 854 464 860 465
rect 854 460 855 464
rect 859 460 860 464
rect 854 459 860 460
rect 902 464 908 465
rect 902 460 903 464
rect 907 460 908 464
rect 902 459 908 460
rect 958 464 964 465
rect 958 460 959 464
rect 963 460 964 464
rect 958 459 964 460
rect 1006 464 1012 465
rect 1006 460 1007 464
rect 1011 460 1012 464
rect 1006 459 1012 460
rect 1046 464 1052 465
rect 1046 460 1047 464
rect 1051 460 1052 464
rect 1046 459 1052 460
rect 1096 457 1098 477
rect 1136 461 1138 481
rect 1160 469 1162 481
rect 1264 469 1266 481
rect 1384 469 1386 481
rect 1496 469 1498 481
rect 1600 469 1602 481
rect 1704 469 1706 481
rect 1800 469 1802 481
rect 1888 469 1890 481
rect 1984 469 1986 481
rect 2072 469 2074 481
rect 1158 468 1164 469
rect 1158 464 1159 468
rect 1163 464 1164 468
rect 1158 463 1164 464
rect 1262 468 1268 469
rect 1262 464 1263 468
rect 1267 464 1268 468
rect 1262 463 1268 464
rect 1382 468 1388 469
rect 1382 464 1383 468
rect 1387 464 1388 468
rect 1382 463 1388 464
rect 1494 468 1500 469
rect 1494 464 1495 468
rect 1499 464 1500 468
rect 1494 463 1500 464
rect 1598 468 1604 469
rect 1598 464 1599 468
rect 1603 464 1604 468
rect 1598 463 1604 464
rect 1702 468 1708 469
rect 1702 464 1703 468
rect 1707 464 1708 468
rect 1702 463 1708 464
rect 1798 468 1804 469
rect 1798 464 1799 468
rect 1803 464 1804 468
rect 1798 463 1804 464
rect 1886 468 1892 469
rect 1886 464 1887 468
rect 1891 464 1892 468
rect 1886 463 1892 464
rect 1982 468 1988 469
rect 1982 464 1983 468
rect 1987 464 1988 468
rect 1982 463 1988 464
rect 2070 468 2076 469
rect 2070 464 2071 468
rect 2075 464 2076 468
rect 2070 463 2076 464
rect 2120 461 2122 481
rect 1134 460 1140 461
rect 110 456 116 457
rect 110 452 111 456
rect 115 452 116 456
rect 110 451 116 452
rect 1094 456 1100 457
rect 1094 452 1095 456
rect 1099 452 1100 456
rect 1134 456 1135 460
rect 1139 456 1140 460
rect 1134 455 1140 456
rect 2118 460 2124 461
rect 2118 456 2119 460
rect 2123 456 2124 460
rect 2118 455 2124 456
rect 1094 451 1100 452
rect 1134 443 1140 444
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 1094 439 1100 440
rect 110 434 116 435
rect 166 436 172 437
rect 112 431 114 434
rect 166 432 167 436
rect 171 432 172 436
rect 166 431 172 432
rect 230 436 236 437
rect 230 432 231 436
rect 235 432 236 436
rect 230 431 236 432
rect 302 436 308 437
rect 302 432 303 436
rect 307 432 308 436
rect 302 431 308 432
rect 374 436 380 437
rect 374 432 375 436
rect 379 432 380 436
rect 374 431 380 432
rect 454 436 460 437
rect 454 432 455 436
rect 459 432 460 436
rect 454 431 460 432
rect 534 436 540 437
rect 534 432 535 436
rect 539 432 540 436
rect 534 431 540 432
rect 606 436 612 437
rect 606 432 607 436
rect 611 432 612 436
rect 606 431 612 432
rect 678 436 684 437
rect 678 432 679 436
rect 683 432 684 436
rect 678 431 684 432
rect 742 436 748 437
rect 742 432 743 436
rect 747 432 748 436
rect 742 431 748 432
rect 798 436 804 437
rect 798 432 799 436
rect 803 432 804 436
rect 798 431 804 432
rect 854 436 860 437
rect 854 432 855 436
rect 859 432 860 436
rect 854 431 860 432
rect 902 436 908 437
rect 902 432 903 436
rect 907 432 908 436
rect 902 431 908 432
rect 958 436 964 437
rect 958 432 959 436
rect 963 432 964 436
rect 958 431 964 432
rect 1006 436 1012 437
rect 1006 432 1007 436
rect 1011 432 1012 436
rect 1006 431 1012 432
rect 1046 436 1052 437
rect 1046 432 1047 436
rect 1051 432 1052 436
rect 1094 435 1095 439
rect 1099 435 1100 439
rect 1134 439 1135 443
rect 1139 439 1140 443
rect 2118 443 2124 444
rect 1134 438 1140 439
rect 1158 440 1164 441
rect 1136 435 1138 438
rect 1158 436 1159 440
rect 1163 436 1164 440
rect 1158 435 1164 436
rect 1262 440 1268 441
rect 1262 436 1263 440
rect 1267 436 1268 440
rect 1262 435 1268 436
rect 1382 440 1388 441
rect 1382 436 1383 440
rect 1387 436 1388 440
rect 1382 435 1388 436
rect 1494 440 1500 441
rect 1494 436 1495 440
rect 1499 436 1500 440
rect 1494 435 1500 436
rect 1598 440 1604 441
rect 1598 436 1599 440
rect 1603 436 1604 440
rect 1598 435 1604 436
rect 1702 440 1708 441
rect 1702 436 1703 440
rect 1707 436 1708 440
rect 1702 435 1708 436
rect 1798 440 1804 441
rect 1798 436 1799 440
rect 1803 436 1804 440
rect 1798 435 1804 436
rect 1886 440 1892 441
rect 1886 436 1887 440
rect 1891 436 1892 440
rect 1886 435 1892 436
rect 1982 440 1988 441
rect 1982 436 1983 440
rect 1987 436 1988 440
rect 1982 435 1988 436
rect 2070 440 2076 441
rect 2070 436 2071 440
rect 2075 436 2076 440
rect 2118 439 2119 443
rect 2123 439 2124 443
rect 2118 438 2124 439
rect 2070 435 2076 436
rect 2120 435 2122 438
rect 1094 434 1100 435
rect 1135 434 1139 435
rect 1046 431 1052 432
rect 1096 431 1098 434
rect 111 430 115 431
rect 111 425 115 426
rect 151 430 155 431
rect 151 425 155 426
rect 167 430 171 431
rect 167 425 171 426
rect 215 430 219 431
rect 215 425 219 426
rect 231 430 235 431
rect 231 425 235 426
rect 279 430 283 431
rect 279 425 283 426
rect 303 430 307 431
rect 303 425 307 426
rect 351 430 355 431
rect 351 425 355 426
rect 375 430 379 431
rect 375 425 379 426
rect 423 430 427 431
rect 423 425 427 426
rect 455 430 459 431
rect 455 425 459 426
rect 487 430 491 431
rect 487 425 491 426
rect 535 430 539 431
rect 535 425 539 426
rect 551 430 555 431
rect 551 425 555 426
rect 607 430 611 431
rect 607 425 611 426
rect 615 430 619 431
rect 615 425 619 426
rect 671 430 675 431
rect 671 425 675 426
rect 679 430 683 431
rect 679 425 683 426
rect 727 430 731 431
rect 727 425 731 426
rect 743 430 747 431
rect 743 425 747 426
rect 791 430 795 431
rect 791 425 795 426
rect 799 430 803 431
rect 799 425 803 426
rect 855 430 859 431
rect 855 425 859 426
rect 903 430 907 431
rect 903 425 907 426
rect 959 430 963 431
rect 959 425 963 426
rect 1007 430 1011 431
rect 1007 425 1011 426
rect 1047 430 1051 431
rect 1047 425 1051 426
rect 1095 430 1099 431
rect 1135 429 1139 430
rect 1159 434 1163 435
rect 1159 429 1163 430
rect 1199 434 1203 435
rect 1199 429 1203 430
rect 1255 434 1259 435
rect 1255 429 1259 430
rect 1263 434 1267 435
rect 1263 429 1267 430
rect 1335 434 1339 435
rect 1335 429 1339 430
rect 1383 434 1387 435
rect 1383 429 1387 430
rect 1415 434 1419 435
rect 1415 429 1419 430
rect 1495 434 1499 435
rect 1495 429 1499 430
rect 1503 434 1507 435
rect 1503 429 1507 430
rect 1591 434 1595 435
rect 1591 429 1595 430
rect 1599 434 1603 435
rect 1599 429 1603 430
rect 1671 434 1675 435
rect 1671 429 1675 430
rect 1703 434 1707 435
rect 1703 429 1707 430
rect 1751 434 1755 435
rect 1751 429 1755 430
rect 1799 434 1803 435
rect 1799 429 1803 430
rect 1823 434 1827 435
rect 1823 429 1827 430
rect 1887 434 1891 435
rect 1887 429 1891 430
rect 1951 434 1955 435
rect 1951 429 1955 430
rect 1983 434 1987 435
rect 1983 429 1987 430
rect 2023 434 2027 435
rect 2023 429 2027 430
rect 2071 434 2075 435
rect 2071 429 2075 430
rect 2119 434 2123 435
rect 2119 429 2123 430
rect 1136 426 1138 429
rect 1158 428 1164 429
rect 1095 425 1099 426
rect 1134 425 1140 426
rect 112 422 114 425
rect 150 424 156 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 150 420 151 424
rect 155 420 156 424
rect 150 419 156 420
rect 214 424 220 425
rect 214 420 215 424
rect 219 420 220 424
rect 214 419 220 420
rect 278 424 284 425
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 350 424 356 425
rect 350 420 351 424
rect 355 420 356 424
rect 350 419 356 420
rect 422 424 428 425
rect 422 420 423 424
rect 427 420 428 424
rect 422 419 428 420
rect 486 424 492 425
rect 486 420 487 424
rect 491 420 492 424
rect 486 419 492 420
rect 550 424 556 425
rect 550 420 551 424
rect 555 420 556 424
rect 550 419 556 420
rect 614 424 620 425
rect 614 420 615 424
rect 619 420 620 424
rect 614 419 620 420
rect 670 424 676 425
rect 670 420 671 424
rect 675 420 676 424
rect 670 419 676 420
rect 726 424 732 425
rect 726 420 727 424
rect 731 420 732 424
rect 726 419 732 420
rect 790 424 796 425
rect 790 420 791 424
rect 795 420 796 424
rect 790 419 796 420
rect 854 424 860 425
rect 854 420 855 424
rect 859 420 860 424
rect 1096 422 1098 425
rect 854 419 860 420
rect 1094 421 1100 422
rect 110 416 116 417
rect 1094 417 1095 421
rect 1099 417 1100 421
rect 1134 421 1135 425
rect 1139 421 1140 425
rect 1158 424 1159 428
rect 1163 424 1164 428
rect 1158 423 1164 424
rect 1198 428 1204 429
rect 1198 424 1199 428
rect 1203 424 1204 428
rect 1198 423 1204 424
rect 1254 428 1260 429
rect 1254 424 1255 428
rect 1259 424 1260 428
rect 1254 423 1260 424
rect 1334 428 1340 429
rect 1334 424 1335 428
rect 1339 424 1340 428
rect 1334 423 1340 424
rect 1414 428 1420 429
rect 1414 424 1415 428
rect 1419 424 1420 428
rect 1414 423 1420 424
rect 1502 428 1508 429
rect 1502 424 1503 428
rect 1507 424 1508 428
rect 1502 423 1508 424
rect 1590 428 1596 429
rect 1590 424 1591 428
rect 1595 424 1596 428
rect 1590 423 1596 424
rect 1670 428 1676 429
rect 1670 424 1671 428
rect 1675 424 1676 428
rect 1670 423 1676 424
rect 1750 428 1756 429
rect 1750 424 1751 428
rect 1755 424 1756 428
rect 1750 423 1756 424
rect 1822 428 1828 429
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1822 423 1828 424
rect 1886 428 1892 429
rect 1886 424 1887 428
rect 1891 424 1892 428
rect 1886 423 1892 424
rect 1950 428 1956 429
rect 1950 424 1951 428
rect 1955 424 1956 428
rect 1950 423 1956 424
rect 2022 428 2028 429
rect 2022 424 2023 428
rect 2027 424 2028 428
rect 2022 423 2028 424
rect 2070 428 2076 429
rect 2070 424 2071 428
rect 2075 424 2076 428
rect 2120 426 2122 429
rect 2070 423 2076 424
rect 2118 425 2124 426
rect 1134 420 1140 421
rect 2118 421 2119 425
rect 2123 421 2124 425
rect 2118 420 2124 421
rect 1094 416 1100 417
rect 1134 408 1140 409
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 1094 404 1100 405
rect 1094 400 1095 404
rect 1099 400 1100 404
rect 1134 404 1135 408
rect 1139 404 1140 408
rect 1134 403 1140 404
rect 2118 408 2124 409
rect 2118 404 2119 408
rect 2123 404 2124 408
rect 2118 403 2124 404
rect 1094 399 1100 400
rect 112 379 114 399
rect 150 396 156 397
rect 150 392 151 396
rect 155 392 156 396
rect 150 391 156 392
rect 214 396 220 397
rect 214 392 215 396
rect 219 392 220 396
rect 214 391 220 392
rect 278 396 284 397
rect 278 392 279 396
rect 283 392 284 396
rect 278 391 284 392
rect 350 396 356 397
rect 350 392 351 396
rect 355 392 356 396
rect 350 391 356 392
rect 422 396 428 397
rect 422 392 423 396
rect 427 392 428 396
rect 422 391 428 392
rect 486 396 492 397
rect 486 392 487 396
rect 491 392 492 396
rect 486 391 492 392
rect 550 396 556 397
rect 550 392 551 396
rect 555 392 556 396
rect 550 391 556 392
rect 614 396 620 397
rect 614 392 615 396
rect 619 392 620 396
rect 614 391 620 392
rect 670 396 676 397
rect 670 392 671 396
rect 675 392 676 396
rect 670 391 676 392
rect 726 396 732 397
rect 726 392 727 396
rect 731 392 732 396
rect 726 391 732 392
rect 790 396 796 397
rect 790 392 791 396
rect 795 392 796 396
rect 790 391 796 392
rect 854 396 860 397
rect 854 392 855 396
rect 859 392 860 396
rect 854 391 860 392
rect 152 379 154 391
rect 216 379 218 391
rect 280 379 282 391
rect 352 379 354 391
rect 424 379 426 391
rect 488 379 490 391
rect 552 379 554 391
rect 616 379 618 391
rect 672 379 674 391
rect 728 379 730 391
rect 792 379 794 391
rect 856 379 858 391
rect 1096 379 1098 399
rect 1136 379 1138 403
rect 1158 400 1164 401
rect 1158 396 1159 400
rect 1163 396 1164 400
rect 1158 395 1164 396
rect 1198 400 1204 401
rect 1198 396 1199 400
rect 1203 396 1204 400
rect 1198 395 1204 396
rect 1254 400 1260 401
rect 1254 396 1255 400
rect 1259 396 1260 400
rect 1254 395 1260 396
rect 1334 400 1340 401
rect 1334 396 1335 400
rect 1339 396 1340 400
rect 1334 395 1340 396
rect 1414 400 1420 401
rect 1414 396 1415 400
rect 1419 396 1420 400
rect 1414 395 1420 396
rect 1502 400 1508 401
rect 1502 396 1503 400
rect 1507 396 1508 400
rect 1502 395 1508 396
rect 1590 400 1596 401
rect 1590 396 1591 400
rect 1595 396 1596 400
rect 1590 395 1596 396
rect 1670 400 1676 401
rect 1670 396 1671 400
rect 1675 396 1676 400
rect 1670 395 1676 396
rect 1750 400 1756 401
rect 1750 396 1751 400
rect 1755 396 1756 400
rect 1750 395 1756 396
rect 1822 400 1828 401
rect 1822 396 1823 400
rect 1827 396 1828 400
rect 1822 395 1828 396
rect 1886 400 1892 401
rect 1886 396 1887 400
rect 1891 396 1892 400
rect 1886 395 1892 396
rect 1950 400 1956 401
rect 1950 396 1951 400
rect 1955 396 1956 400
rect 1950 395 1956 396
rect 2022 400 2028 401
rect 2022 396 2023 400
rect 2027 396 2028 400
rect 2022 395 2028 396
rect 2070 400 2076 401
rect 2070 396 2071 400
rect 2075 396 2076 400
rect 2070 395 2076 396
rect 1160 379 1162 395
rect 1200 379 1202 395
rect 1256 379 1258 395
rect 1336 379 1338 395
rect 1416 379 1418 395
rect 1504 379 1506 395
rect 1592 379 1594 395
rect 1672 379 1674 395
rect 1752 379 1754 395
rect 1824 379 1826 395
rect 1888 379 1890 395
rect 1952 379 1954 395
rect 2024 379 2026 395
rect 2072 379 2074 395
rect 2120 379 2122 403
rect 111 378 115 379
rect 111 373 115 374
rect 135 378 139 379
rect 135 373 139 374
rect 151 378 155 379
rect 151 373 155 374
rect 175 378 179 379
rect 175 373 179 374
rect 215 378 219 379
rect 215 373 219 374
rect 271 378 275 379
rect 271 373 275 374
rect 279 378 283 379
rect 279 373 283 374
rect 335 378 339 379
rect 335 373 339 374
rect 351 378 355 379
rect 351 373 355 374
rect 399 378 403 379
rect 399 373 403 374
rect 423 378 427 379
rect 423 373 427 374
rect 463 378 467 379
rect 463 373 467 374
rect 487 378 491 379
rect 487 373 491 374
rect 519 378 523 379
rect 519 373 523 374
rect 551 378 555 379
rect 551 373 555 374
rect 575 378 579 379
rect 575 373 579 374
rect 615 378 619 379
rect 615 373 619 374
rect 631 378 635 379
rect 631 373 635 374
rect 671 378 675 379
rect 671 373 675 374
rect 687 378 691 379
rect 687 373 691 374
rect 727 378 731 379
rect 727 373 731 374
rect 751 378 755 379
rect 751 373 755 374
rect 791 378 795 379
rect 791 373 795 374
rect 855 378 859 379
rect 855 373 859 374
rect 1095 378 1099 379
rect 1095 373 1099 374
rect 1135 378 1139 379
rect 1135 373 1139 374
rect 1159 378 1163 379
rect 1159 373 1163 374
rect 1199 378 1203 379
rect 1199 373 1203 374
rect 1255 378 1259 379
rect 1255 373 1259 374
rect 1303 378 1307 379
rect 1303 373 1307 374
rect 1335 378 1339 379
rect 1335 373 1339 374
rect 1343 378 1347 379
rect 1343 373 1347 374
rect 1383 378 1387 379
rect 1383 373 1387 374
rect 1415 378 1419 379
rect 1415 373 1419 374
rect 1423 378 1427 379
rect 1423 373 1427 374
rect 1463 378 1467 379
rect 1463 373 1467 374
rect 1503 378 1507 379
rect 1503 373 1507 374
rect 1551 378 1555 379
rect 1551 373 1555 374
rect 1591 378 1595 379
rect 1591 373 1595 374
rect 1615 378 1619 379
rect 1615 373 1619 374
rect 1671 378 1675 379
rect 1671 373 1675 374
rect 1679 378 1683 379
rect 1679 373 1683 374
rect 1751 378 1755 379
rect 1751 373 1755 374
rect 1823 378 1827 379
rect 1823 373 1827 374
rect 1831 378 1835 379
rect 1831 373 1835 374
rect 1887 378 1891 379
rect 1887 373 1891 374
rect 1919 378 1923 379
rect 1919 373 1923 374
rect 1951 378 1955 379
rect 1951 373 1955 374
rect 2007 378 2011 379
rect 2007 373 2011 374
rect 2023 378 2027 379
rect 2023 373 2027 374
rect 2071 378 2075 379
rect 2071 373 2075 374
rect 2119 378 2123 379
rect 2119 373 2123 374
rect 112 353 114 373
rect 136 361 138 373
rect 176 361 178 373
rect 216 361 218 373
rect 272 361 274 373
rect 336 361 338 373
rect 400 361 402 373
rect 464 361 466 373
rect 520 361 522 373
rect 576 361 578 373
rect 632 361 634 373
rect 688 361 690 373
rect 752 361 754 373
rect 134 360 140 361
rect 134 356 135 360
rect 139 356 140 360
rect 134 355 140 356
rect 174 360 180 361
rect 174 356 175 360
rect 179 356 180 360
rect 174 355 180 356
rect 214 360 220 361
rect 214 356 215 360
rect 219 356 220 360
rect 214 355 220 356
rect 270 360 276 361
rect 270 356 271 360
rect 275 356 276 360
rect 270 355 276 356
rect 334 360 340 361
rect 334 356 335 360
rect 339 356 340 360
rect 334 355 340 356
rect 398 360 404 361
rect 398 356 399 360
rect 403 356 404 360
rect 398 355 404 356
rect 462 360 468 361
rect 462 356 463 360
rect 467 356 468 360
rect 462 355 468 356
rect 518 360 524 361
rect 518 356 519 360
rect 523 356 524 360
rect 518 355 524 356
rect 574 360 580 361
rect 574 356 575 360
rect 579 356 580 360
rect 574 355 580 356
rect 630 360 636 361
rect 630 356 631 360
rect 635 356 636 360
rect 630 355 636 356
rect 686 360 692 361
rect 686 356 687 360
rect 691 356 692 360
rect 686 355 692 356
rect 750 360 756 361
rect 750 356 751 360
rect 755 356 756 360
rect 750 355 756 356
rect 1096 353 1098 373
rect 1136 353 1138 373
rect 1304 361 1306 373
rect 1344 361 1346 373
rect 1384 361 1386 373
rect 1424 361 1426 373
rect 1464 361 1466 373
rect 1504 361 1506 373
rect 1552 361 1554 373
rect 1616 361 1618 373
rect 1680 361 1682 373
rect 1752 361 1754 373
rect 1832 361 1834 373
rect 1920 361 1922 373
rect 2008 361 2010 373
rect 2072 361 2074 373
rect 1302 360 1308 361
rect 1302 356 1303 360
rect 1307 356 1308 360
rect 1302 355 1308 356
rect 1342 360 1348 361
rect 1342 356 1343 360
rect 1347 356 1348 360
rect 1342 355 1348 356
rect 1382 360 1388 361
rect 1382 356 1383 360
rect 1387 356 1388 360
rect 1382 355 1388 356
rect 1422 360 1428 361
rect 1422 356 1423 360
rect 1427 356 1428 360
rect 1422 355 1428 356
rect 1462 360 1468 361
rect 1462 356 1463 360
rect 1467 356 1468 360
rect 1462 355 1468 356
rect 1502 360 1508 361
rect 1502 356 1503 360
rect 1507 356 1508 360
rect 1502 355 1508 356
rect 1550 360 1556 361
rect 1550 356 1551 360
rect 1555 356 1556 360
rect 1550 355 1556 356
rect 1614 360 1620 361
rect 1614 356 1615 360
rect 1619 356 1620 360
rect 1614 355 1620 356
rect 1678 360 1684 361
rect 1678 356 1679 360
rect 1683 356 1684 360
rect 1678 355 1684 356
rect 1750 360 1756 361
rect 1750 356 1751 360
rect 1755 356 1756 360
rect 1750 355 1756 356
rect 1830 360 1836 361
rect 1830 356 1831 360
rect 1835 356 1836 360
rect 1830 355 1836 356
rect 1918 360 1924 361
rect 1918 356 1919 360
rect 1923 356 1924 360
rect 1918 355 1924 356
rect 2006 360 2012 361
rect 2006 356 2007 360
rect 2011 356 2012 360
rect 2006 355 2012 356
rect 2070 360 2076 361
rect 2070 356 2071 360
rect 2075 356 2076 360
rect 2070 355 2076 356
rect 2120 353 2122 373
rect 110 352 116 353
rect 110 348 111 352
rect 115 348 116 352
rect 110 347 116 348
rect 1094 352 1100 353
rect 1094 348 1095 352
rect 1099 348 1100 352
rect 1094 347 1100 348
rect 1134 352 1140 353
rect 1134 348 1135 352
rect 1139 348 1140 352
rect 1134 347 1140 348
rect 2118 352 2124 353
rect 2118 348 2119 352
rect 2123 348 2124 352
rect 2118 347 2124 348
rect 110 335 116 336
rect 110 331 111 335
rect 115 331 116 335
rect 1094 335 1100 336
rect 110 330 116 331
rect 134 332 140 333
rect 112 323 114 330
rect 134 328 135 332
rect 139 328 140 332
rect 134 327 140 328
rect 174 332 180 333
rect 174 328 175 332
rect 179 328 180 332
rect 174 327 180 328
rect 214 332 220 333
rect 214 328 215 332
rect 219 328 220 332
rect 214 327 220 328
rect 270 332 276 333
rect 270 328 271 332
rect 275 328 276 332
rect 270 327 276 328
rect 334 332 340 333
rect 334 328 335 332
rect 339 328 340 332
rect 334 327 340 328
rect 398 332 404 333
rect 398 328 399 332
rect 403 328 404 332
rect 398 327 404 328
rect 462 332 468 333
rect 462 328 463 332
rect 467 328 468 332
rect 462 327 468 328
rect 518 332 524 333
rect 518 328 519 332
rect 523 328 524 332
rect 518 327 524 328
rect 574 332 580 333
rect 574 328 575 332
rect 579 328 580 332
rect 574 327 580 328
rect 630 332 636 333
rect 630 328 631 332
rect 635 328 636 332
rect 630 327 636 328
rect 686 332 692 333
rect 686 328 687 332
rect 691 328 692 332
rect 686 327 692 328
rect 750 332 756 333
rect 750 328 751 332
rect 755 328 756 332
rect 1094 331 1095 335
rect 1099 331 1100 335
rect 1094 330 1100 331
rect 1134 335 1140 336
rect 1134 331 1135 335
rect 1139 331 1140 335
rect 2118 335 2124 336
rect 1134 330 1140 331
rect 1302 332 1308 333
rect 750 327 756 328
rect 136 323 138 327
rect 176 323 178 327
rect 216 323 218 327
rect 272 323 274 327
rect 336 323 338 327
rect 400 323 402 327
rect 464 323 466 327
rect 520 323 522 327
rect 576 323 578 327
rect 632 323 634 327
rect 688 323 690 327
rect 752 323 754 327
rect 1096 323 1098 330
rect 1136 323 1138 330
rect 1302 328 1303 332
rect 1307 328 1308 332
rect 1302 327 1308 328
rect 1342 332 1348 333
rect 1342 328 1343 332
rect 1347 328 1348 332
rect 1342 327 1348 328
rect 1382 332 1388 333
rect 1382 328 1383 332
rect 1387 328 1388 332
rect 1382 327 1388 328
rect 1422 332 1428 333
rect 1422 328 1423 332
rect 1427 328 1428 332
rect 1422 327 1428 328
rect 1462 332 1468 333
rect 1462 328 1463 332
rect 1467 328 1468 332
rect 1462 327 1468 328
rect 1502 332 1508 333
rect 1502 328 1503 332
rect 1507 328 1508 332
rect 1502 327 1508 328
rect 1550 332 1556 333
rect 1550 328 1551 332
rect 1555 328 1556 332
rect 1550 327 1556 328
rect 1614 332 1620 333
rect 1614 328 1615 332
rect 1619 328 1620 332
rect 1614 327 1620 328
rect 1678 332 1684 333
rect 1678 328 1679 332
rect 1683 328 1684 332
rect 1678 327 1684 328
rect 1750 332 1756 333
rect 1750 328 1751 332
rect 1755 328 1756 332
rect 1750 327 1756 328
rect 1830 332 1836 333
rect 1830 328 1831 332
rect 1835 328 1836 332
rect 1830 327 1836 328
rect 1918 332 1924 333
rect 1918 328 1919 332
rect 1923 328 1924 332
rect 1918 327 1924 328
rect 2006 332 2012 333
rect 2006 328 2007 332
rect 2011 328 2012 332
rect 2006 327 2012 328
rect 2070 332 2076 333
rect 2070 328 2071 332
rect 2075 328 2076 332
rect 2118 331 2119 335
rect 2123 331 2124 335
rect 2118 330 2124 331
rect 2070 327 2076 328
rect 1304 323 1306 327
rect 1344 323 1346 327
rect 1384 323 1386 327
rect 1424 323 1426 327
rect 1464 323 1466 327
rect 1504 323 1506 327
rect 1552 323 1554 327
rect 1616 323 1618 327
rect 1680 323 1682 327
rect 1752 323 1754 327
rect 1832 323 1834 327
rect 1920 323 1922 327
rect 2008 323 2010 327
rect 2072 323 2074 327
rect 2120 323 2122 330
rect 111 322 115 323
rect 111 317 115 318
rect 135 322 139 323
rect 135 317 139 318
rect 175 322 179 323
rect 175 317 179 318
rect 207 322 211 323
rect 207 317 211 318
rect 215 322 219 323
rect 215 317 219 318
rect 271 322 275 323
rect 271 317 275 318
rect 295 322 299 323
rect 295 317 299 318
rect 335 322 339 323
rect 335 317 339 318
rect 383 322 387 323
rect 383 317 387 318
rect 399 322 403 323
rect 399 317 403 318
rect 463 322 467 323
rect 463 317 467 318
rect 471 322 475 323
rect 471 317 475 318
rect 519 322 523 323
rect 519 317 523 318
rect 551 322 555 323
rect 551 317 555 318
rect 575 322 579 323
rect 575 317 579 318
rect 623 322 627 323
rect 623 317 627 318
rect 631 322 635 323
rect 631 317 635 318
rect 687 322 691 323
rect 687 317 691 318
rect 751 322 755 323
rect 751 317 755 318
rect 807 322 811 323
rect 807 317 811 318
rect 871 322 875 323
rect 871 317 875 318
rect 935 322 939 323
rect 935 317 939 318
rect 1095 322 1099 323
rect 1095 317 1099 318
rect 1135 322 1139 323
rect 1135 317 1139 318
rect 1167 322 1171 323
rect 1167 317 1171 318
rect 1207 322 1211 323
rect 1207 317 1211 318
rect 1247 322 1251 323
rect 1247 317 1251 318
rect 1295 322 1299 323
rect 1295 317 1299 318
rect 1303 322 1307 323
rect 1303 317 1307 318
rect 1343 322 1347 323
rect 1343 317 1347 318
rect 1383 322 1387 323
rect 1383 317 1387 318
rect 1391 322 1395 323
rect 1391 317 1395 318
rect 1423 322 1427 323
rect 1423 317 1427 318
rect 1439 322 1443 323
rect 1439 317 1443 318
rect 1463 322 1467 323
rect 1463 317 1467 318
rect 1495 322 1499 323
rect 1495 317 1499 318
rect 1503 322 1507 323
rect 1503 317 1507 318
rect 1551 322 1555 323
rect 1551 317 1555 318
rect 1559 322 1563 323
rect 1559 317 1563 318
rect 1615 322 1619 323
rect 1615 317 1619 318
rect 1623 322 1627 323
rect 1623 317 1627 318
rect 1679 322 1683 323
rect 1679 317 1683 318
rect 1695 322 1699 323
rect 1695 317 1699 318
rect 1751 322 1755 323
rect 1751 317 1755 318
rect 1775 322 1779 323
rect 1775 317 1779 318
rect 1831 322 1835 323
rect 1831 317 1835 318
rect 1855 322 1859 323
rect 1855 317 1859 318
rect 1919 322 1923 323
rect 1919 317 1923 318
rect 1935 322 1939 323
rect 1935 317 1939 318
rect 2007 322 2011 323
rect 2007 317 2011 318
rect 2015 322 2019 323
rect 2015 317 2019 318
rect 2071 322 2075 323
rect 2071 317 2075 318
rect 2119 322 2123 323
rect 2119 317 2123 318
rect 112 314 114 317
rect 134 316 140 317
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 134 312 135 316
rect 139 312 140 316
rect 134 311 140 312
rect 206 316 212 317
rect 206 312 207 316
rect 211 312 212 316
rect 206 311 212 312
rect 294 316 300 317
rect 294 312 295 316
rect 299 312 300 316
rect 294 311 300 312
rect 382 316 388 317
rect 382 312 383 316
rect 387 312 388 316
rect 382 311 388 312
rect 470 316 476 317
rect 470 312 471 316
rect 475 312 476 316
rect 470 311 476 312
rect 550 316 556 317
rect 550 312 551 316
rect 555 312 556 316
rect 550 311 556 312
rect 622 316 628 317
rect 622 312 623 316
rect 627 312 628 316
rect 622 311 628 312
rect 686 316 692 317
rect 686 312 687 316
rect 691 312 692 316
rect 686 311 692 312
rect 750 316 756 317
rect 750 312 751 316
rect 755 312 756 316
rect 750 311 756 312
rect 806 316 812 317
rect 806 312 807 316
rect 811 312 812 316
rect 806 311 812 312
rect 870 316 876 317
rect 870 312 871 316
rect 875 312 876 316
rect 870 311 876 312
rect 934 316 940 317
rect 934 312 935 316
rect 939 312 940 316
rect 1096 314 1098 317
rect 1136 314 1138 317
rect 1166 316 1172 317
rect 934 311 940 312
rect 1094 313 1100 314
rect 110 308 116 309
rect 1094 309 1095 313
rect 1099 309 1100 313
rect 1094 308 1100 309
rect 1134 313 1140 314
rect 1134 309 1135 313
rect 1139 309 1140 313
rect 1166 312 1167 316
rect 1171 312 1172 316
rect 1166 311 1172 312
rect 1206 316 1212 317
rect 1206 312 1207 316
rect 1211 312 1212 316
rect 1206 311 1212 312
rect 1246 316 1252 317
rect 1246 312 1247 316
rect 1251 312 1252 316
rect 1246 311 1252 312
rect 1294 316 1300 317
rect 1294 312 1295 316
rect 1299 312 1300 316
rect 1294 311 1300 312
rect 1342 316 1348 317
rect 1342 312 1343 316
rect 1347 312 1348 316
rect 1342 311 1348 312
rect 1390 316 1396 317
rect 1390 312 1391 316
rect 1395 312 1396 316
rect 1390 311 1396 312
rect 1438 316 1444 317
rect 1438 312 1439 316
rect 1443 312 1444 316
rect 1438 311 1444 312
rect 1494 316 1500 317
rect 1494 312 1495 316
rect 1499 312 1500 316
rect 1494 311 1500 312
rect 1558 316 1564 317
rect 1558 312 1559 316
rect 1563 312 1564 316
rect 1558 311 1564 312
rect 1622 316 1628 317
rect 1622 312 1623 316
rect 1627 312 1628 316
rect 1622 311 1628 312
rect 1694 316 1700 317
rect 1694 312 1695 316
rect 1699 312 1700 316
rect 1694 311 1700 312
rect 1774 316 1780 317
rect 1774 312 1775 316
rect 1779 312 1780 316
rect 1774 311 1780 312
rect 1854 316 1860 317
rect 1854 312 1855 316
rect 1859 312 1860 316
rect 1854 311 1860 312
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 1934 311 1940 312
rect 2014 316 2020 317
rect 2014 312 2015 316
rect 2019 312 2020 316
rect 2014 311 2020 312
rect 2070 316 2076 317
rect 2070 312 2071 316
rect 2075 312 2076 316
rect 2120 314 2122 317
rect 2070 311 2076 312
rect 2118 313 2124 314
rect 1134 308 1140 309
rect 2118 309 2119 313
rect 2123 309 2124 313
rect 2118 308 2124 309
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 1094 296 1100 297
rect 1094 292 1095 296
rect 1099 292 1100 296
rect 1094 291 1100 292
rect 1134 296 1140 297
rect 1134 292 1135 296
rect 1139 292 1140 296
rect 1134 291 1140 292
rect 2118 296 2124 297
rect 2118 292 2119 296
rect 2123 292 2124 296
rect 2118 291 2124 292
rect 112 271 114 291
rect 134 288 140 289
rect 134 284 135 288
rect 139 284 140 288
rect 134 283 140 284
rect 206 288 212 289
rect 206 284 207 288
rect 211 284 212 288
rect 206 283 212 284
rect 294 288 300 289
rect 294 284 295 288
rect 299 284 300 288
rect 294 283 300 284
rect 382 288 388 289
rect 382 284 383 288
rect 387 284 388 288
rect 382 283 388 284
rect 470 288 476 289
rect 470 284 471 288
rect 475 284 476 288
rect 470 283 476 284
rect 550 288 556 289
rect 550 284 551 288
rect 555 284 556 288
rect 550 283 556 284
rect 622 288 628 289
rect 622 284 623 288
rect 627 284 628 288
rect 622 283 628 284
rect 686 288 692 289
rect 686 284 687 288
rect 691 284 692 288
rect 686 283 692 284
rect 750 288 756 289
rect 750 284 751 288
rect 755 284 756 288
rect 750 283 756 284
rect 806 288 812 289
rect 806 284 807 288
rect 811 284 812 288
rect 806 283 812 284
rect 870 288 876 289
rect 870 284 871 288
rect 875 284 876 288
rect 870 283 876 284
rect 934 288 940 289
rect 934 284 935 288
rect 939 284 940 288
rect 934 283 940 284
rect 136 271 138 283
rect 208 271 210 283
rect 296 271 298 283
rect 384 271 386 283
rect 472 271 474 283
rect 552 271 554 283
rect 624 271 626 283
rect 688 271 690 283
rect 752 271 754 283
rect 808 271 810 283
rect 872 271 874 283
rect 936 271 938 283
rect 1096 271 1098 291
rect 111 270 115 271
rect 111 265 115 266
rect 135 270 139 271
rect 135 265 139 266
rect 199 270 203 271
rect 199 265 203 266
rect 207 270 211 271
rect 207 265 211 266
rect 279 270 283 271
rect 279 265 283 266
rect 295 270 299 271
rect 295 265 299 266
rect 359 270 363 271
rect 359 265 363 266
rect 383 270 387 271
rect 383 265 387 266
rect 439 270 443 271
rect 439 265 443 266
rect 471 270 475 271
rect 471 265 475 266
rect 511 270 515 271
rect 511 265 515 266
rect 551 270 555 271
rect 551 265 555 266
rect 583 270 587 271
rect 583 265 587 266
rect 623 270 627 271
rect 623 265 627 266
rect 647 270 651 271
rect 647 265 651 266
rect 687 270 691 271
rect 687 265 691 266
rect 703 270 707 271
rect 703 265 707 266
rect 751 270 755 271
rect 751 265 755 266
rect 759 270 763 271
rect 759 265 763 266
rect 807 270 811 271
rect 807 265 811 266
rect 815 270 819 271
rect 815 265 819 266
rect 871 270 875 271
rect 871 265 875 266
rect 879 270 883 271
rect 879 265 883 266
rect 935 270 939 271
rect 935 265 939 266
rect 1095 270 1099 271
rect 1095 265 1099 266
rect 112 245 114 265
rect 136 253 138 265
rect 200 253 202 265
rect 280 253 282 265
rect 360 253 362 265
rect 440 253 442 265
rect 512 253 514 265
rect 584 253 586 265
rect 648 253 650 265
rect 704 253 706 265
rect 760 253 762 265
rect 816 253 818 265
rect 880 253 882 265
rect 134 252 140 253
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 198 252 204 253
rect 198 248 199 252
rect 203 248 204 252
rect 198 247 204 248
rect 278 252 284 253
rect 278 248 279 252
rect 283 248 284 252
rect 278 247 284 248
rect 358 252 364 253
rect 358 248 359 252
rect 363 248 364 252
rect 358 247 364 248
rect 438 252 444 253
rect 438 248 439 252
rect 443 248 444 252
rect 438 247 444 248
rect 510 252 516 253
rect 510 248 511 252
rect 515 248 516 252
rect 510 247 516 248
rect 582 252 588 253
rect 582 248 583 252
rect 587 248 588 252
rect 582 247 588 248
rect 646 252 652 253
rect 646 248 647 252
rect 651 248 652 252
rect 646 247 652 248
rect 702 252 708 253
rect 702 248 703 252
rect 707 248 708 252
rect 702 247 708 248
rect 758 252 764 253
rect 758 248 759 252
rect 763 248 764 252
rect 758 247 764 248
rect 814 252 820 253
rect 814 248 815 252
rect 819 248 820 252
rect 814 247 820 248
rect 878 252 884 253
rect 878 248 879 252
rect 883 248 884 252
rect 878 247 884 248
rect 1096 245 1098 265
rect 1136 263 1138 291
rect 1166 288 1172 289
rect 1166 284 1167 288
rect 1171 284 1172 288
rect 1166 283 1172 284
rect 1206 288 1212 289
rect 1206 284 1207 288
rect 1211 284 1212 288
rect 1206 283 1212 284
rect 1246 288 1252 289
rect 1246 284 1247 288
rect 1251 284 1252 288
rect 1246 283 1252 284
rect 1294 288 1300 289
rect 1294 284 1295 288
rect 1299 284 1300 288
rect 1294 283 1300 284
rect 1342 288 1348 289
rect 1342 284 1343 288
rect 1347 284 1348 288
rect 1342 283 1348 284
rect 1390 288 1396 289
rect 1390 284 1391 288
rect 1395 284 1396 288
rect 1390 283 1396 284
rect 1438 288 1444 289
rect 1438 284 1439 288
rect 1443 284 1444 288
rect 1438 283 1444 284
rect 1494 288 1500 289
rect 1494 284 1495 288
rect 1499 284 1500 288
rect 1494 283 1500 284
rect 1558 288 1564 289
rect 1558 284 1559 288
rect 1563 284 1564 288
rect 1558 283 1564 284
rect 1622 288 1628 289
rect 1622 284 1623 288
rect 1627 284 1628 288
rect 1622 283 1628 284
rect 1694 288 1700 289
rect 1694 284 1695 288
rect 1699 284 1700 288
rect 1694 283 1700 284
rect 1774 288 1780 289
rect 1774 284 1775 288
rect 1779 284 1780 288
rect 1774 283 1780 284
rect 1854 288 1860 289
rect 1854 284 1855 288
rect 1859 284 1860 288
rect 1854 283 1860 284
rect 1934 288 1940 289
rect 1934 284 1935 288
rect 1939 284 1940 288
rect 1934 283 1940 284
rect 2014 288 2020 289
rect 2014 284 2015 288
rect 2019 284 2020 288
rect 2014 283 2020 284
rect 2070 288 2076 289
rect 2070 284 2071 288
rect 2075 284 2076 288
rect 2070 283 2076 284
rect 1168 263 1170 283
rect 1208 263 1210 283
rect 1248 263 1250 283
rect 1296 263 1298 283
rect 1344 263 1346 283
rect 1392 263 1394 283
rect 1440 263 1442 283
rect 1496 263 1498 283
rect 1560 263 1562 283
rect 1624 263 1626 283
rect 1696 263 1698 283
rect 1776 263 1778 283
rect 1856 263 1858 283
rect 1936 263 1938 283
rect 2016 263 2018 283
rect 2072 263 2074 283
rect 2120 263 2122 291
rect 1135 262 1139 263
rect 1135 257 1139 258
rect 1159 262 1163 263
rect 1159 257 1163 258
rect 1167 262 1171 263
rect 1167 257 1171 258
rect 1207 262 1211 263
rect 1207 257 1211 258
rect 1247 262 1251 263
rect 1247 257 1251 258
rect 1271 262 1275 263
rect 1271 257 1275 258
rect 1295 262 1299 263
rect 1295 257 1299 258
rect 1327 262 1331 263
rect 1327 257 1331 258
rect 1343 262 1347 263
rect 1343 257 1347 258
rect 1391 262 1395 263
rect 1391 257 1395 258
rect 1439 262 1443 263
rect 1439 257 1443 258
rect 1455 262 1459 263
rect 1455 257 1459 258
rect 1495 262 1499 263
rect 1495 257 1499 258
rect 1527 262 1531 263
rect 1527 257 1531 258
rect 1559 262 1563 263
rect 1559 257 1563 258
rect 1607 262 1611 263
rect 1607 257 1611 258
rect 1623 262 1627 263
rect 1623 257 1627 258
rect 1687 262 1691 263
rect 1687 257 1691 258
rect 1695 262 1699 263
rect 1695 257 1699 258
rect 1767 262 1771 263
rect 1767 257 1771 258
rect 1775 262 1779 263
rect 1775 257 1779 258
rect 1839 262 1843 263
rect 1839 257 1843 258
rect 1855 262 1859 263
rect 1855 257 1859 258
rect 1919 262 1923 263
rect 1919 257 1923 258
rect 1935 262 1939 263
rect 1935 257 1939 258
rect 1999 262 2003 263
rect 1999 257 2003 258
rect 2015 262 2019 263
rect 2015 257 2019 258
rect 2071 262 2075 263
rect 2071 257 2075 258
rect 2119 262 2123 263
rect 2119 257 2123 258
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 110 239 116 240
rect 1094 244 1100 245
rect 1094 240 1095 244
rect 1099 240 1100 244
rect 1094 239 1100 240
rect 1136 237 1138 257
rect 1160 245 1162 257
rect 1208 245 1210 257
rect 1272 245 1274 257
rect 1328 245 1330 257
rect 1392 245 1394 257
rect 1456 245 1458 257
rect 1528 245 1530 257
rect 1608 245 1610 257
rect 1688 245 1690 257
rect 1768 245 1770 257
rect 1840 245 1842 257
rect 1920 245 1922 257
rect 2000 245 2002 257
rect 2072 245 2074 257
rect 1158 244 1164 245
rect 1158 240 1159 244
rect 1163 240 1164 244
rect 1158 239 1164 240
rect 1206 244 1212 245
rect 1206 240 1207 244
rect 1211 240 1212 244
rect 1206 239 1212 240
rect 1270 244 1276 245
rect 1270 240 1271 244
rect 1275 240 1276 244
rect 1270 239 1276 240
rect 1326 244 1332 245
rect 1326 240 1327 244
rect 1331 240 1332 244
rect 1326 239 1332 240
rect 1390 244 1396 245
rect 1390 240 1391 244
rect 1395 240 1396 244
rect 1390 239 1396 240
rect 1454 244 1460 245
rect 1454 240 1455 244
rect 1459 240 1460 244
rect 1454 239 1460 240
rect 1526 244 1532 245
rect 1526 240 1527 244
rect 1531 240 1532 244
rect 1526 239 1532 240
rect 1606 244 1612 245
rect 1606 240 1607 244
rect 1611 240 1612 244
rect 1606 239 1612 240
rect 1686 244 1692 245
rect 1686 240 1687 244
rect 1691 240 1692 244
rect 1686 239 1692 240
rect 1766 244 1772 245
rect 1766 240 1767 244
rect 1771 240 1772 244
rect 1766 239 1772 240
rect 1838 244 1844 245
rect 1838 240 1839 244
rect 1843 240 1844 244
rect 1838 239 1844 240
rect 1918 244 1924 245
rect 1918 240 1919 244
rect 1923 240 1924 244
rect 1918 239 1924 240
rect 1998 244 2004 245
rect 1998 240 1999 244
rect 2003 240 2004 244
rect 1998 239 2004 240
rect 2070 244 2076 245
rect 2070 240 2071 244
rect 2075 240 2076 244
rect 2070 239 2076 240
rect 2120 237 2122 257
rect 1134 236 1140 237
rect 1134 232 1135 236
rect 1139 232 1140 236
rect 1134 231 1140 232
rect 2118 236 2124 237
rect 2118 232 2119 236
rect 2123 232 2124 236
rect 2118 231 2124 232
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1094 227 1100 228
rect 110 222 116 223
rect 134 224 140 225
rect 112 215 114 222
rect 134 220 135 224
rect 139 220 140 224
rect 134 219 140 220
rect 198 224 204 225
rect 198 220 199 224
rect 203 220 204 224
rect 198 219 204 220
rect 278 224 284 225
rect 278 220 279 224
rect 283 220 284 224
rect 278 219 284 220
rect 358 224 364 225
rect 358 220 359 224
rect 363 220 364 224
rect 358 219 364 220
rect 438 224 444 225
rect 438 220 439 224
rect 443 220 444 224
rect 438 219 444 220
rect 510 224 516 225
rect 510 220 511 224
rect 515 220 516 224
rect 510 219 516 220
rect 582 224 588 225
rect 582 220 583 224
rect 587 220 588 224
rect 582 219 588 220
rect 646 224 652 225
rect 646 220 647 224
rect 651 220 652 224
rect 646 219 652 220
rect 702 224 708 225
rect 702 220 703 224
rect 707 220 708 224
rect 702 219 708 220
rect 758 224 764 225
rect 758 220 759 224
rect 763 220 764 224
rect 758 219 764 220
rect 814 224 820 225
rect 814 220 815 224
rect 819 220 820 224
rect 814 219 820 220
rect 878 224 884 225
rect 878 220 879 224
rect 883 220 884 224
rect 1094 223 1095 227
rect 1099 223 1100 227
rect 1094 222 1100 223
rect 878 219 884 220
rect 136 215 138 219
rect 200 215 202 219
rect 280 215 282 219
rect 360 215 362 219
rect 440 215 442 219
rect 512 215 514 219
rect 584 215 586 219
rect 648 215 650 219
rect 704 215 706 219
rect 760 215 762 219
rect 816 215 818 219
rect 880 215 882 219
rect 1096 215 1098 222
rect 1134 219 1140 220
rect 1134 215 1135 219
rect 1139 215 1140 219
rect 2118 219 2124 220
rect 111 214 115 215
rect 111 209 115 210
rect 135 214 139 215
rect 135 209 139 210
rect 183 214 187 215
rect 183 209 187 210
rect 199 214 203 215
rect 199 209 203 210
rect 231 214 235 215
rect 231 209 235 210
rect 279 214 283 215
rect 279 209 283 210
rect 327 214 331 215
rect 327 209 331 210
rect 359 214 363 215
rect 359 209 363 210
rect 375 214 379 215
rect 375 209 379 210
rect 415 214 419 215
rect 415 209 419 210
rect 439 214 443 215
rect 439 209 443 210
rect 455 214 459 215
rect 455 209 459 210
rect 503 214 507 215
rect 503 209 507 210
rect 511 214 515 215
rect 511 209 515 210
rect 551 214 555 215
rect 551 209 555 210
rect 583 214 587 215
rect 583 209 587 210
rect 599 214 603 215
rect 599 209 603 210
rect 647 214 651 215
rect 647 209 651 210
rect 695 214 699 215
rect 695 209 699 210
rect 703 214 707 215
rect 703 209 707 210
rect 743 214 747 215
rect 743 209 747 210
rect 759 214 763 215
rect 759 209 763 210
rect 815 214 819 215
rect 815 209 819 210
rect 879 214 883 215
rect 879 209 883 210
rect 1095 214 1099 215
rect 1134 214 1140 215
rect 1158 216 1164 217
rect 1136 211 1138 214
rect 1158 212 1159 216
rect 1163 212 1164 216
rect 1158 211 1164 212
rect 1206 216 1212 217
rect 1206 212 1207 216
rect 1211 212 1212 216
rect 1206 211 1212 212
rect 1270 216 1276 217
rect 1270 212 1271 216
rect 1275 212 1276 216
rect 1270 211 1276 212
rect 1326 216 1332 217
rect 1326 212 1327 216
rect 1331 212 1332 216
rect 1326 211 1332 212
rect 1390 216 1396 217
rect 1390 212 1391 216
rect 1395 212 1396 216
rect 1390 211 1396 212
rect 1454 216 1460 217
rect 1454 212 1455 216
rect 1459 212 1460 216
rect 1454 211 1460 212
rect 1526 216 1532 217
rect 1526 212 1527 216
rect 1531 212 1532 216
rect 1526 211 1532 212
rect 1606 216 1612 217
rect 1606 212 1607 216
rect 1611 212 1612 216
rect 1606 211 1612 212
rect 1686 216 1692 217
rect 1686 212 1687 216
rect 1691 212 1692 216
rect 1686 211 1692 212
rect 1766 216 1772 217
rect 1766 212 1767 216
rect 1771 212 1772 216
rect 1766 211 1772 212
rect 1838 216 1844 217
rect 1838 212 1839 216
rect 1843 212 1844 216
rect 1838 211 1844 212
rect 1918 216 1924 217
rect 1918 212 1919 216
rect 1923 212 1924 216
rect 1918 211 1924 212
rect 1998 216 2004 217
rect 1998 212 1999 216
rect 2003 212 2004 216
rect 1998 211 2004 212
rect 2070 216 2076 217
rect 2070 212 2071 216
rect 2075 212 2076 216
rect 2118 215 2119 219
rect 2123 215 2124 219
rect 2118 214 2124 215
rect 2070 211 2076 212
rect 2120 211 2122 214
rect 1095 209 1099 210
rect 1135 210 1139 211
rect 112 206 114 209
rect 134 208 140 209
rect 110 205 116 206
rect 110 201 111 205
rect 115 201 116 205
rect 134 204 135 208
rect 139 204 140 208
rect 134 203 140 204
rect 182 208 188 209
rect 182 204 183 208
rect 187 204 188 208
rect 182 203 188 204
rect 230 208 236 209
rect 230 204 231 208
rect 235 204 236 208
rect 230 203 236 204
rect 278 208 284 209
rect 278 204 279 208
rect 283 204 284 208
rect 278 203 284 204
rect 326 208 332 209
rect 326 204 327 208
rect 331 204 332 208
rect 326 203 332 204
rect 374 208 380 209
rect 374 204 375 208
rect 379 204 380 208
rect 374 203 380 204
rect 414 208 420 209
rect 414 204 415 208
rect 419 204 420 208
rect 414 203 420 204
rect 454 208 460 209
rect 454 204 455 208
rect 459 204 460 208
rect 454 203 460 204
rect 502 208 508 209
rect 502 204 503 208
rect 507 204 508 208
rect 502 203 508 204
rect 550 208 556 209
rect 550 204 551 208
rect 555 204 556 208
rect 550 203 556 204
rect 598 208 604 209
rect 598 204 599 208
rect 603 204 604 208
rect 598 203 604 204
rect 646 208 652 209
rect 646 204 647 208
rect 651 204 652 208
rect 646 203 652 204
rect 694 208 700 209
rect 694 204 695 208
rect 699 204 700 208
rect 694 203 700 204
rect 742 208 748 209
rect 742 204 743 208
rect 747 204 748 208
rect 1096 206 1098 209
rect 742 203 748 204
rect 1094 205 1100 206
rect 1135 205 1139 206
rect 1159 210 1163 211
rect 1159 205 1163 206
rect 1199 210 1203 211
rect 1199 205 1203 206
rect 1207 210 1211 211
rect 1207 205 1211 206
rect 1263 210 1267 211
rect 1263 205 1267 206
rect 1271 210 1275 211
rect 1271 205 1275 206
rect 1327 210 1331 211
rect 1327 205 1331 206
rect 1391 210 1395 211
rect 1391 205 1395 206
rect 1399 210 1403 211
rect 1399 205 1403 206
rect 1455 210 1459 211
rect 1455 205 1459 206
rect 1471 210 1475 211
rect 1471 205 1475 206
rect 1527 210 1531 211
rect 1527 205 1531 206
rect 1543 210 1547 211
rect 1543 205 1547 206
rect 1607 210 1611 211
rect 1607 205 1611 206
rect 1671 210 1675 211
rect 1671 205 1675 206
rect 1687 210 1691 211
rect 1687 205 1691 206
rect 1735 210 1739 211
rect 1735 205 1739 206
rect 1767 210 1771 211
rect 1767 205 1771 206
rect 1807 210 1811 211
rect 1807 205 1811 206
rect 1839 210 1843 211
rect 1839 205 1843 206
rect 1879 210 1883 211
rect 1879 205 1883 206
rect 1919 210 1923 211
rect 1919 205 1923 206
rect 1951 210 1955 211
rect 1951 205 1955 206
rect 1999 210 2003 211
rect 1999 205 2003 206
rect 2023 210 2027 211
rect 2023 205 2027 206
rect 2071 210 2075 211
rect 2071 205 2075 206
rect 2119 210 2123 211
rect 2119 205 2123 206
rect 110 200 116 201
rect 1094 201 1095 205
rect 1099 201 1100 205
rect 1136 202 1138 205
rect 1158 204 1164 205
rect 1094 200 1100 201
rect 1134 201 1140 202
rect 1134 197 1135 201
rect 1139 197 1140 201
rect 1158 200 1159 204
rect 1163 200 1164 204
rect 1158 199 1164 200
rect 1198 204 1204 205
rect 1198 200 1199 204
rect 1203 200 1204 204
rect 1198 199 1204 200
rect 1262 204 1268 205
rect 1262 200 1263 204
rect 1267 200 1268 204
rect 1262 199 1268 200
rect 1326 204 1332 205
rect 1326 200 1327 204
rect 1331 200 1332 204
rect 1326 199 1332 200
rect 1398 204 1404 205
rect 1398 200 1399 204
rect 1403 200 1404 204
rect 1398 199 1404 200
rect 1470 204 1476 205
rect 1470 200 1471 204
rect 1475 200 1476 204
rect 1470 199 1476 200
rect 1542 204 1548 205
rect 1542 200 1543 204
rect 1547 200 1548 204
rect 1542 199 1548 200
rect 1606 204 1612 205
rect 1606 200 1607 204
rect 1611 200 1612 204
rect 1606 199 1612 200
rect 1670 204 1676 205
rect 1670 200 1671 204
rect 1675 200 1676 204
rect 1670 199 1676 200
rect 1734 204 1740 205
rect 1734 200 1735 204
rect 1739 200 1740 204
rect 1734 199 1740 200
rect 1806 204 1812 205
rect 1806 200 1807 204
rect 1811 200 1812 204
rect 1806 199 1812 200
rect 1878 204 1884 205
rect 1878 200 1879 204
rect 1883 200 1884 204
rect 1878 199 1884 200
rect 1950 204 1956 205
rect 1950 200 1951 204
rect 1955 200 1956 204
rect 1950 199 1956 200
rect 2022 204 2028 205
rect 2022 200 2023 204
rect 2027 200 2028 204
rect 2022 199 2028 200
rect 2070 204 2076 205
rect 2070 200 2071 204
rect 2075 200 2076 204
rect 2120 202 2122 205
rect 2070 199 2076 200
rect 2118 201 2124 202
rect 1134 196 1140 197
rect 2118 197 2119 201
rect 2123 197 2124 201
rect 2118 196 2124 197
rect 110 188 116 189
rect 110 184 111 188
rect 115 184 116 188
rect 110 183 116 184
rect 1094 188 1100 189
rect 1094 184 1095 188
rect 1099 184 1100 188
rect 1094 183 1100 184
rect 1134 184 1140 185
rect 112 139 114 183
rect 134 180 140 181
rect 134 176 135 180
rect 139 176 140 180
rect 134 175 140 176
rect 182 180 188 181
rect 182 176 183 180
rect 187 176 188 180
rect 182 175 188 176
rect 230 180 236 181
rect 230 176 231 180
rect 235 176 236 180
rect 230 175 236 176
rect 278 180 284 181
rect 278 176 279 180
rect 283 176 284 180
rect 278 175 284 176
rect 326 180 332 181
rect 326 176 327 180
rect 331 176 332 180
rect 326 175 332 176
rect 374 180 380 181
rect 374 176 375 180
rect 379 176 380 180
rect 374 175 380 176
rect 414 180 420 181
rect 414 176 415 180
rect 419 176 420 180
rect 414 175 420 176
rect 454 180 460 181
rect 454 176 455 180
rect 459 176 460 180
rect 454 175 460 176
rect 502 180 508 181
rect 502 176 503 180
rect 507 176 508 180
rect 502 175 508 176
rect 550 180 556 181
rect 550 176 551 180
rect 555 176 556 180
rect 550 175 556 176
rect 598 180 604 181
rect 598 176 599 180
rect 603 176 604 180
rect 598 175 604 176
rect 646 180 652 181
rect 646 176 647 180
rect 651 176 652 180
rect 646 175 652 176
rect 694 180 700 181
rect 694 176 695 180
rect 699 176 700 180
rect 694 175 700 176
rect 742 180 748 181
rect 742 176 743 180
rect 747 176 748 180
rect 742 175 748 176
rect 136 139 138 175
rect 184 139 186 175
rect 232 139 234 175
rect 280 139 282 175
rect 328 139 330 175
rect 376 139 378 175
rect 416 139 418 175
rect 456 139 458 175
rect 504 139 506 175
rect 552 139 554 175
rect 600 139 602 175
rect 648 139 650 175
rect 696 139 698 175
rect 744 139 746 175
rect 1096 139 1098 183
rect 1134 180 1135 184
rect 1139 180 1140 184
rect 1134 179 1140 180
rect 2118 184 2124 185
rect 2118 180 2119 184
rect 2123 180 2124 184
rect 2118 179 2124 180
rect 1136 139 1138 179
rect 1158 176 1164 177
rect 1158 172 1159 176
rect 1163 172 1164 176
rect 1158 171 1164 172
rect 1198 176 1204 177
rect 1198 172 1199 176
rect 1203 172 1204 176
rect 1198 171 1204 172
rect 1262 176 1268 177
rect 1262 172 1263 176
rect 1267 172 1268 176
rect 1262 171 1268 172
rect 1326 176 1332 177
rect 1326 172 1327 176
rect 1331 172 1332 176
rect 1326 171 1332 172
rect 1398 176 1404 177
rect 1398 172 1399 176
rect 1403 172 1404 176
rect 1398 171 1404 172
rect 1470 176 1476 177
rect 1470 172 1471 176
rect 1475 172 1476 176
rect 1470 171 1476 172
rect 1542 176 1548 177
rect 1542 172 1543 176
rect 1547 172 1548 176
rect 1542 171 1548 172
rect 1606 176 1612 177
rect 1606 172 1607 176
rect 1611 172 1612 176
rect 1606 171 1612 172
rect 1670 176 1676 177
rect 1670 172 1671 176
rect 1675 172 1676 176
rect 1670 171 1676 172
rect 1734 176 1740 177
rect 1734 172 1735 176
rect 1739 172 1740 176
rect 1734 171 1740 172
rect 1806 176 1812 177
rect 1806 172 1807 176
rect 1811 172 1812 176
rect 1806 171 1812 172
rect 1878 176 1884 177
rect 1878 172 1879 176
rect 1883 172 1884 176
rect 1878 171 1884 172
rect 1950 176 1956 177
rect 1950 172 1951 176
rect 1955 172 1956 176
rect 1950 171 1956 172
rect 2022 176 2028 177
rect 2022 172 2023 176
rect 2027 172 2028 176
rect 2022 171 2028 172
rect 2070 176 2076 177
rect 2070 172 2071 176
rect 2075 172 2076 176
rect 2070 171 2076 172
rect 1160 139 1162 171
rect 1200 139 1202 171
rect 1264 139 1266 171
rect 1328 139 1330 171
rect 1400 139 1402 171
rect 1472 139 1474 171
rect 1544 139 1546 171
rect 1608 139 1610 171
rect 1672 139 1674 171
rect 1736 139 1738 171
rect 1808 139 1810 171
rect 1880 139 1882 171
rect 1952 139 1954 171
rect 2024 139 2026 171
rect 2072 139 2074 171
rect 2120 139 2122 179
rect 111 138 115 139
rect 111 133 115 134
rect 135 138 139 139
rect 135 133 139 134
rect 143 138 147 139
rect 143 133 147 134
rect 183 138 187 139
rect 183 133 187 134
rect 223 138 227 139
rect 223 133 227 134
rect 231 138 235 139
rect 231 133 235 134
rect 263 138 267 139
rect 263 133 267 134
rect 279 138 283 139
rect 279 133 283 134
rect 303 138 307 139
rect 303 133 307 134
rect 327 138 331 139
rect 327 133 331 134
rect 343 138 347 139
rect 343 133 347 134
rect 375 138 379 139
rect 375 133 379 134
rect 383 138 387 139
rect 383 133 387 134
rect 415 138 419 139
rect 415 133 419 134
rect 423 138 427 139
rect 423 133 427 134
rect 455 138 459 139
rect 455 133 459 134
rect 463 138 467 139
rect 463 133 467 134
rect 503 138 507 139
rect 503 133 507 134
rect 543 138 547 139
rect 543 133 547 134
rect 551 138 555 139
rect 551 133 555 134
rect 583 138 587 139
rect 583 133 587 134
rect 599 138 603 139
rect 599 133 603 134
rect 623 138 627 139
rect 623 133 627 134
rect 647 138 651 139
rect 647 133 651 134
rect 663 138 667 139
rect 663 133 667 134
rect 695 138 699 139
rect 695 133 699 134
rect 703 138 707 139
rect 703 133 707 134
rect 743 138 747 139
rect 743 133 747 134
rect 783 138 787 139
rect 783 133 787 134
rect 831 138 835 139
rect 831 133 835 134
rect 879 138 883 139
rect 879 133 883 134
rect 927 138 931 139
rect 927 133 931 134
rect 967 138 971 139
rect 967 133 971 134
rect 1007 138 1011 139
rect 1007 133 1011 134
rect 1047 138 1051 139
rect 1047 133 1051 134
rect 1095 138 1099 139
rect 1095 133 1099 134
rect 1135 138 1139 139
rect 1135 133 1139 134
rect 1159 138 1163 139
rect 1159 133 1163 134
rect 1199 138 1203 139
rect 1199 133 1203 134
rect 1207 138 1211 139
rect 1207 133 1211 134
rect 1263 138 1267 139
rect 1263 133 1267 134
rect 1271 138 1275 139
rect 1271 133 1275 134
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 1335 138 1339 139
rect 1335 133 1339 134
rect 1399 138 1403 139
rect 1399 133 1403 134
rect 1455 138 1459 139
rect 1455 133 1459 134
rect 1471 138 1475 139
rect 1471 133 1475 134
rect 1511 138 1515 139
rect 1511 133 1515 134
rect 1543 138 1547 139
rect 1543 133 1547 134
rect 1559 138 1563 139
rect 1559 133 1563 134
rect 1607 138 1611 139
rect 1607 133 1611 134
rect 1647 138 1651 139
rect 1647 133 1651 134
rect 1671 138 1675 139
rect 1671 133 1675 134
rect 1687 138 1691 139
rect 1687 133 1691 134
rect 1727 138 1731 139
rect 1727 133 1731 134
rect 1735 138 1739 139
rect 1735 133 1739 134
rect 1767 138 1771 139
rect 1767 133 1771 134
rect 1807 138 1811 139
rect 1807 133 1811 134
rect 1855 138 1859 139
rect 1855 133 1859 134
rect 1879 138 1883 139
rect 1879 133 1883 134
rect 1903 138 1907 139
rect 1903 133 1907 134
rect 1951 138 1955 139
rect 1951 133 1955 134
rect 1991 138 1995 139
rect 1991 133 1995 134
rect 2023 138 2027 139
rect 2023 133 2027 134
rect 2031 138 2035 139
rect 2031 133 2035 134
rect 2071 138 2075 139
rect 2071 133 2075 134
rect 2119 138 2123 139
rect 2119 133 2123 134
rect 112 113 114 133
rect 144 121 146 133
rect 184 121 186 133
rect 224 121 226 133
rect 264 121 266 133
rect 304 121 306 133
rect 344 121 346 133
rect 384 121 386 133
rect 424 121 426 133
rect 464 121 466 133
rect 504 121 506 133
rect 544 121 546 133
rect 584 121 586 133
rect 624 121 626 133
rect 664 121 666 133
rect 704 121 706 133
rect 744 121 746 133
rect 784 121 786 133
rect 832 121 834 133
rect 880 121 882 133
rect 928 121 930 133
rect 968 121 970 133
rect 1008 121 1010 133
rect 1048 121 1050 133
rect 142 120 148 121
rect 142 116 143 120
rect 147 116 148 120
rect 142 115 148 116
rect 182 120 188 121
rect 182 116 183 120
rect 187 116 188 120
rect 182 115 188 116
rect 222 120 228 121
rect 222 116 223 120
rect 227 116 228 120
rect 222 115 228 116
rect 262 120 268 121
rect 262 116 263 120
rect 267 116 268 120
rect 262 115 268 116
rect 302 120 308 121
rect 302 116 303 120
rect 307 116 308 120
rect 302 115 308 116
rect 342 120 348 121
rect 342 116 343 120
rect 347 116 348 120
rect 342 115 348 116
rect 382 120 388 121
rect 382 116 383 120
rect 387 116 388 120
rect 382 115 388 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 462 120 468 121
rect 462 116 463 120
rect 467 116 468 120
rect 462 115 468 116
rect 502 120 508 121
rect 502 116 503 120
rect 507 116 508 120
rect 502 115 508 116
rect 542 120 548 121
rect 542 116 543 120
rect 547 116 548 120
rect 542 115 548 116
rect 582 120 588 121
rect 582 116 583 120
rect 587 116 588 120
rect 582 115 588 116
rect 622 120 628 121
rect 622 116 623 120
rect 627 116 628 120
rect 622 115 628 116
rect 662 120 668 121
rect 662 116 663 120
rect 667 116 668 120
rect 662 115 668 116
rect 702 120 708 121
rect 702 116 703 120
rect 707 116 708 120
rect 702 115 708 116
rect 742 120 748 121
rect 742 116 743 120
rect 747 116 748 120
rect 742 115 748 116
rect 782 120 788 121
rect 782 116 783 120
rect 787 116 788 120
rect 782 115 788 116
rect 830 120 836 121
rect 830 116 831 120
rect 835 116 836 120
rect 830 115 836 116
rect 878 120 884 121
rect 878 116 879 120
rect 883 116 884 120
rect 878 115 884 116
rect 926 120 932 121
rect 926 116 927 120
rect 931 116 932 120
rect 926 115 932 116
rect 966 120 972 121
rect 966 116 967 120
rect 971 116 972 120
rect 966 115 972 116
rect 1006 120 1012 121
rect 1006 116 1007 120
rect 1011 116 1012 120
rect 1006 115 1012 116
rect 1046 120 1052 121
rect 1046 116 1047 120
rect 1051 116 1052 120
rect 1046 115 1052 116
rect 1096 113 1098 133
rect 1136 113 1138 133
rect 1160 121 1162 133
rect 1208 121 1210 133
rect 1272 121 1274 133
rect 1336 121 1338 133
rect 1400 121 1402 133
rect 1456 121 1458 133
rect 1512 121 1514 133
rect 1560 121 1562 133
rect 1608 121 1610 133
rect 1648 121 1650 133
rect 1688 121 1690 133
rect 1728 121 1730 133
rect 1768 121 1770 133
rect 1808 121 1810 133
rect 1856 121 1858 133
rect 1904 121 1906 133
rect 1952 121 1954 133
rect 1992 121 1994 133
rect 2032 121 2034 133
rect 2072 121 2074 133
rect 1158 120 1164 121
rect 1158 116 1159 120
rect 1163 116 1164 120
rect 1158 115 1164 116
rect 1206 120 1212 121
rect 1206 116 1207 120
rect 1211 116 1212 120
rect 1206 115 1212 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1334 120 1340 121
rect 1334 116 1335 120
rect 1339 116 1340 120
rect 1334 115 1340 116
rect 1398 120 1404 121
rect 1398 116 1399 120
rect 1403 116 1404 120
rect 1398 115 1404 116
rect 1454 120 1460 121
rect 1454 116 1455 120
rect 1459 116 1460 120
rect 1454 115 1460 116
rect 1510 120 1516 121
rect 1510 116 1511 120
rect 1515 116 1516 120
rect 1510 115 1516 116
rect 1558 120 1564 121
rect 1558 116 1559 120
rect 1563 116 1564 120
rect 1558 115 1564 116
rect 1606 120 1612 121
rect 1606 116 1607 120
rect 1611 116 1612 120
rect 1606 115 1612 116
rect 1646 120 1652 121
rect 1646 116 1647 120
rect 1651 116 1652 120
rect 1646 115 1652 116
rect 1686 120 1692 121
rect 1686 116 1687 120
rect 1691 116 1692 120
rect 1686 115 1692 116
rect 1726 120 1732 121
rect 1726 116 1727 120
rect 1731 116 1732 120
rect 1726 115 1732 116
rect 1766 120 1772 121
rect 1766 116 1767 120
rect 1771 116 1772 120
rect 1766 115 1772 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1854 120 1860 121
rect 1854 116 1855 120
rect 1859 116 1860 120
rect 1854 115 1860 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 1902 115 1908 116
rect 1950 120 1956 121
rect 1950 116 1951 120
rect 1955 116 1956 120
rect 1950 115 1956 116
rect 1990 120 1996 121
rect 1990 116 1991 120
rect 1995 116 1996 120
rect 1990 115 1996 116
rect 2030 120 2036 121
rect 2030 116 2031 120
rect 2035 116 2036 120
rect 2030 115 2036 116
rect 2070 120 2076 121
rect 2070 116 2071 120
rect 2075 116 2076 120
rect 2070 115 2076 116
rect 2120 113 2122 133
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 110 107 116 108
rect 1094 112 1100 113
rect 1094 108 1095 112
rect 1099 108 1100 112
rect 1094 107 1100 108
rect 1134 112 1140 113
rect 1134 108 1135 112
rect 1139 108 1140 112
rect 1134 107 1140 108
rect 2118 112 2124 113
rect 2118 108 2119 112
rect 2123 108 2124 112
rect 2118 107 2124 108
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1094 95 1100 96
rect 110 90 116 91
rect 142 92 148 93
rect 112 87 114 90
rect 142 88 143 92
rect 147 88 148 92
rect 142 87 148 88
rect 182 92 188 93
rect 182 88 183 92
rect 187 88 188 92
rect 182 87 188 88
rect 222 92 228 93
rect 222 88 223 92
rect 227 88 228 92
rect 222 87 228 88
rect 262 92 268 93
rect 262 88 263 92
rect 267 88 268 92
rect 262 87 268 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 342 92 348 93
rect 342 88 343 92
rect 347 88 348 92
rect 342 87 348 88
rect 382 92 388 93
rect 382 88 383 92
rect 387 88 388 92
rect 382 87 388 88
rect 422 92 428 93
rect 422 88 423 92
rect 427 88 428 92
rect 422 87 428 88
rect 462 92 468 93
rect 462 88 463 92
rect 467 88 468 92
rect 462 87 468 88
rect 502 92 508 93
rect 502 88 503 92
rect 507 88 508 92
rect 502 87 508 88
rect 542 92 548 93
rect 542 88 543 92
rect 547 88 548 92
rect 542 87 548 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 622 92 628 93
rect 622 88 623 92
rect 627 88 628 92
rect 622 87 628 88
rect 662 92 668 93
rect 662 88 663 92
rect 667 88 668 92
rect 662 87 668 88
rect 702 92 708 93
rect 702 88 703 92
rect 707 88 708 92
rect 702 87 708 88
rect 742 92 748 93
rect 742 88 743 92
rect 747 88 748 92
rect 742 87 748 88
rect 782 92 788 93
rect 782 88 783 92
rect 787 88 788 92
rect 782 87 788 88
rect 830 92 836 93
rect 830 88 831 92
rect 835 88 836 92
rect 830 87 836 88
rect 878 92 884 93
rect 878 88 879 92
rect 883 88 884 92
rect 878 87 884 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 966 92 972 93
rect 966 88 967 92
rect 971 88 972 92
rect 966 87 972 88
rect 1006 92 1012 93
rect 1006 88 1007 92
rect 1011 88 1012 92
rect 1006 87 1012 88
rect 1046 92 1052 93
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1094 91 1095 95
rect 1099 91 1100 95
rect 1094 90 1100 91
rect 1134 95 1140 96
rect 1134 91 1135 95
rect 1139 91 1140 95
rect 2118 95 2124 96
rect 1134 90 1140 91
rect 1158 92 1164 93
rect 1046 87 1052 88
rect 1096 87 1098 90
rect 1136 87 1138 90
rect 1158 88 1159 92
rect 1163 88 1164 92
rect 1158 87 1164 88
rect 1206 92 1212 93
rect 1206 88 1207 92
rect 1211 88 1212 92
rect 1206 87 1212 88
rect 1270 92 1276 93
rect 1270 88 1271 92
rect 1275 88 1276 92
rect 1270 87 1276 88
rect 1334 92 1340 93
rect 1334 88 1335 92
rect 1339 88 1340 92
rect 1334 87 1340 88
rect 1398 92 1404 93
rect 1398 88 1399 92
rect 1403 88 1404 92
rect 1398 87 1404 88
rect 1454 92 1460 93
rect 1454 88 1455 92
rect 1459 88 1460 92
rect 1454 87 1460 88
rect 1510 92 1516 93
rect 1510 88 1511 92
rect 1515 88 1516 92
rect 1510 87 1516 88
rect 1558 92 1564 93
rect 1558 88 1559 92
rect 1563 88 1564 92
rect 1558 87 1564 88
rect 1606 92 1612 93
rect 1606 88 1607 92
rect 1611 88 1612 92
rect 1606 87 1612 88
rect 1646 92 1652 93
rect 1646 88 1647 92
rect 1651 88 1652 92
rect 1646 87 1652 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1726 92 1732 93
rect 1726 88 1727 92
rect 1731 88 1732 92
rect 1726 87 1732 88
rect 1766 92 1772 93
rect 1766 88 1767 92
rect 1771 88 1772 92
rect 1766 87 1772 88
rect 1806 92 1812 93
rect 1806 88 1807 92
rect 1811 88 1812 92
rect 1806 87 1812 88
rect 1854 92 1860 93
rect 1854 88 1855 92
rect 1859 88 1860 92
rect 1854 87 1860 88
rect 1902 92 1908 93
rect 1902 88 1903 92
rect 1907 88 1908 92
rect 1902 87 1908 88
rect 1950 92 1956 93
rect 1950 88 1951 92
rect 1955 88 1956 92
rect 1950 87 1956 88
rect 1990 92 1996 93
rect 1990 88 1991 92
rect 1995 88 1996 92
rect 1990 87 1996 88
rect 2030 92 2036 93
rect 2030 88 2031 92
rect 2035 88 2036 92
rect 2030 87 2036 88
rect 2070 92 2076 93
rect 2070 88 2071 92
rect 2075 88 2076 92
rect 2118 91 2119 95
rect 2123 91 2124 95
rect 2118 90 2124 91
rect 2070 87 2076 88
rect 2120 87 2122 90
rect 111 86 115 87
rect 111 81 115 82
rect 143 86 147 87
rect 143 81 147 82
rect 183 86 187 87
rect 183 81 187 82
rect 223 86 227 87
rect 223 81 227 82
rect 263 86 267 87
rect 263 81 267 82
rect 303 86 307 87
rect 303 81 307 82
rect 343 86 347 87
rect 343 81 347 82
rect 383 86 387 87
rect 383 81 387 82
rect 423 86 427 87
rect 423 81 427 82
rect 463 86 467 87
rect 463 81 467 82
rect 503 86 507 87
rect 503 81 507 82
rect 543 86 547 87
rect 543 81 547 82
rect 583 86 587 87
rect 583 81 587 82
rect 623 86 627 87
rect 623 81 627 82
rect 663 86 667 87
rect 663 81 667 82
rect 703 86 707 87
rect 703 81 707 82
rect 743 86 747 87
rect 743 81 747 82
rect 783 86 787 87
rect 783 81 787 82
rect 831 86 835 87
rect 831 81 835 82
rect 879 86 883 87
rect 879 81 883 82
rect 927 86 931 87
rect 927 81 931 82
rect 967 86 971 87
rect 967 81 971 82
rect 1007 86 1011 87
rect 1007 81 1011 82
rect 1047 86 1051 87
rect 1047 81 1051 82
rect 1095 86 1099 87
rect 1095 81 1099 82
rect 1135 86 1139 87
rect 1135 81 1139 82
rect 1159 86 1163 87
rect 1159 81 1163 82
rect 1207 86 1211 87
rect 1207 81 1211 82
rect 1271 86 1275 87
rect 1271 81 1275 82
rect 1335 86 1339 87
rect 1335 81 1339 82
rect 1399 86 1403 87
rect 1399 81 1403 82
rect 1455 86 1459 87
rect 1455 81 1459 82
rect 1511 86 1515 87
rect 1511 81 1515 82
rect 1559 86 1563 87
rect 1559 81 1563 82
rect 1607 86 1611 87
rect 1607 81 1611 82
rect 1647 86 1651 87
rect 1647 81 1651 82
rect 1687 86 1691 87
rect 1687 81 1691 82
rect 1727 86 1731 87
rect 1727 81 1731 82
rect 1767 86 1771 87
rect 1767 81 1771 82
rect 1807 86 1811 87
rect 1807 81 1811 82
rect 1855 86 1859 87
rect 1855 81 1859 82
rect 1903 86 1907 87
rect 1903 81 1907 82
rect 1951 86 1955 87
rect 1951 81 1955 82
rect 1991 86 1995 87
rect 1991 81 1995 82
rect 2031 86 2035 87
rect 2031 81 2035 82
rect 2071 86 2075 87
rect 2071 81 2075 82
rect 2119 86 2123 87
rect 2119 81 2123 82
<< m4c >>
rect 1135 2226 1139 2230
rect 1687 2226 1691 2230
rect 1727 2226 1731 2230
rect 1767 2226 1771 2230
rect 1807 2226 1811 2230
rect 2119 2226 2123 2230
rect 111 2210 115 2214
rect 135 2210 139 2214
rect 175 2210 179 2214
rect 215 2210 219 2214
rect 255 2210 259 2214
rect 319 2210 323 2214
rect 383 2210 387 2214
rect 447 2210 451 2214
rect 511 2210 515 2214
rect 575 2210 579 2214
rect 631 2210 635 2214
rect 687 2210 691 2214
rect 735 2210 739 2214
rect 791 2210 795 2214
rect 847 2210 851 2214
rect 903 2210 907 2214
rect 1095 2210 1099 2214
rect 1135 2174 1139 2178
rect 1159 2174 1163 2178
rect 1199 2174 1203 2178
rect 1239 2174 1243 2178
rect 1279 2174 1283 2178
rect 1335 2174 1339 2178
rect 1391 2174 1395 2178
rect 1455 2174 1459 2178
rect 1527 2174 1531 2178
rect 1591 2174 1595 2178
rect 1663 2174 1667 2178
rect 1687 2174 1691 2178
rect 1727 2174 1731 2178
rect 1735 2174 1739 2178
rect 1767 2174 1771 2178
rect 1807 2174 1811 2178
rect 1879 2174 1883 2178
rect 2119 2174 2123 2178
rect 111 2150 115 2154
rect 135 2150 139 2154
rect 175 2150 179 2154
rect 215 2150 219 2154
rect 231 2150 235 2154
rect 255 2150 259 2154
rect 271 2150 275 2154
rect 311 2150 315 2154
rect 319 2150 323 2154
rect 359 2150 363 2154
rect 383 2150 387 2154
rect 423 2150 427 2154
rect 447 2150 451 2154
rect 487 2150 491 2154
rect 511 2150 515 2154
rect 559 2150 563 2154
rect 575 2150 579 2154
rect 631 2150 635 2154
rect 639 2150 643 2154
rect 687 2150 691 2154
rect 719 2150 723 2154
rect 735 2150 739 2154
rect 791 2150 795 2154
rect 799 2150 803 2154
rect 847 2150 851 2154
rect 879 2150 883 2154
rect 903 2150 907 2154
rect 967 2150 971 2154
rect 1095 2150 1099 2154
rect 1135 2122 1139 2126
rect 1159 2122 1163 2126
rect 1199 2122 1203 2126
rect 1239 2122 1243 2126
rect 1279 2122 1283 2126
rect 1295 2122 1299 2126
rect 1335 2122 1339 2126
rect 1367 2122 1371 2126
rect 1391 2122 1395 2126
rect 1439 2122 1443 2126
rect 1455 2122 1459 2126
rect 1519 2122 1523 2126
rect 1527 2122 1531 2126
rect 1591 2122 1595 2126
rect 1599 2122 1603 2126
rect 1663 2122 1667 2126
rect 1679 2122 1683 2126
rect 1735 2122 1739 2126
rect 1751 2122 1755 2126
rect 1807 2122 1811 2126
rect 1823 2122 1827 2126
rect 1879 2122 1883 2126
rect 1887 2122 1891 2126
rect 1951 2122 1955 2126
rect 2023 2122 2027 2126
rect 2071 2122 2075 2126
rect 2119 2122 2123 2126
rect 111 2094 115 2098
rect 231 2094 235 2098
rect 271 2094 275 2098
rect 303 2094 307 2098
rect 311 2094 315 2098
rect 351 2094 355 2098
rect 359 2094 363 2098
rect 407 2094 411 2098
rect 423 2094 427 2098
rect 471 2094 475 2098
rect 487 2094 491 2098
rect 543 2094 547 2098
rect 559 2094 563 2098
rect 623 2094 627 2098
rect 639 2094 643 2098
rect 703 2094 707 2098
rect 719 2094 723 2098
rect 783 2094 787 2098
rect 799 2094 803 2098
rect 863 2094 867 2098
rect 879 2094 883 2098
rect 951 2094 955 2098
rect 967 2094 971 2098
rect 1039 2094 1043 2098
rect 1095 2094 1099 2098
rect 1135 2070 1139 2074
rect 1159 2070 1163 2074
rect 1199 2070 1203 2074
rect 1215 2070 1219 2074
rect 1239 2070 1243 2074
rect 1295 2070 1299 2074
rect 1303 2070 1307 2074
rect 1367 2070 1371 2074
rect 1399 2070 1403 2074
rect 1439 2070 1443 2074
rect 1495 2070 1499 2074
rect 1519 2070 1523 2074
rect 1591 2070 1595 2074
rect 1599 2070 1603 2074
rect 1679 2070 1683 2074
rect 1751 2070 1755 2074
rect 1759 2070 1763 2074
rect 1823 2070 1827 2074
rect 1831 2070 1835 2074
rect 1887 2070 1891 2074
rect 1895 2070 1899 2074
rect 1951 2070 1955 2074
rect 1959 2070 1963 2074
rect 2023 2070 2027 2074
rect 2071 2070 2075 2074
rect 2119 2070 2123 2074
rect 111 2038 115 2042
rect 183 2038 187 2042
rect 279 2038 283 2042
rect 303 2038 307 2042
rect 351 2038 355 2042
rect 375 2038 379 2042
rect 407 2038 411 2042
rect 463 2038 467 2042
rect 471 2038 475 2042
rect 543 2038 547 2042
rect 623 2038 627 2042
rect 695 2038 699 2042
rect 703 2038 707 2042
rect 759 2038 763 2042
rect 783 2038 787 2042
rect 815 2038 819 2042
rect 863 2038 867 2042
rect 911 2038 915 2042
rect 951 2038 955 2042
rect 959 2038 963 2042
rect 1007 2038 1011 2042
rect 1039 2038 1043 2042
rect 1047 2038 1051 2042
rect 1095 2038 1099 2042
rect 1135 2018 1139 2022
rect 1159 2018 1163 2022
rect 1215 2018 1219 2022
rect 1239 2018 1243 2022
rect 1303 2018 1307 2022
rect 1351 2018 1355 2022
rect 1399 2018 1403 2022
rect 1455 2018 1459 2022
rect 1495 2018 1499 2022
rect 1559 2018 1563 2022
rect 1591 2018 1595 2022
rect 1655 2018 1659 2022
rect 1679 2018 1683 2022
rect 1743 2018 1747 2022
rect 1759 2018 1763 2022
rect 1823 2018 1827 2022
rect 1831 2018 1835 2022
rect 1895 2018 1899 2022
rect 1959 2018 1963 2022
rect 2023 2018 2027 2022
rect 2071 2018 2075 2022
rect 2119 2018 2123 2022
rect 111 1986 115 1990
rect 159 1986 163 1990
rect 183 1986 187 1990
rect 231 1986 235 1990
rect 279 1986 283 1990
rect 303 1986 307 1990
rect 375 1986 379 1990
rect 447 1986 451 1990
rect 463 1986 467 1990
rect 527 1986 531 1990
rect 543 1986 547 1990
rect 607 1986 611 1990
rect 623 1986 627 1990
rect 687 1986 691 1990
rect 695 1986 699 1990
rect 759 1986 763 1990
rect 815 1986 819 1990
rect 831 1986 835 1990
rect 863 1986 867 1990
rect 911 1986 915 1990
rect 959 1986 963 1990
rect 991 1986 995 1990
rect 1007 1986 1011 1990
rect 1047 1986 1051 1990
rect 1095 1986 1099 1990
rect 1135 1954 1139 1958
rect 1159 1954 1163 1958
rect 1239 1954 1243 1958
rect 1351 1954 1355 1958
rect 1359 1954 1363 1958
rect 1423 1954 1427 1958
rect 1455 1954 1459 1958
rect 1487 1954 1491 1958
rect 1559 1954 1563 1958
rect 1631 1954 1635 1958
rect 1655 1954 1659 1958
rect 1703 1954 1707 1958
rect 1743 1954 1747 1958
rect 1775 1954 1779 1958
rect 1823 1954 1827 1958
rect 1847 1954 1851 1958
rect 1895 1954 1899 1958
rect 1927 1954 1931 1958
rect 1959 1954 1963 1958
rect 2007 1954 2011 1958
rect 2023 1954 2027 1958
rect 2071 1954 2075 1958
rect 2119 1954 2123 1958
rect 111 1930 115 1934
rect 135 1930 139 1934
rect 159 1930 163 1934
rect 175 1930 179 1934
rect 231 1930 235 1934
rect 295 1930 299 1934
rect 303 1930 307 1934
rect 367 1930 371 1934
rect 375 1930 379 1934
rect 447 1930 451 1934
rect 527 1930 531 1934
rect 607 1930 611 1934
rect 615 1930 619 1934
rect 687 1930 691 1934
rect 703 1930 707 1934
rect 759 1930 763 1934
rect 791 1930 795 1934
rect 831 1930 835 1934
rect 879 1930 883 1934
rect 911 1930 915 1934
rect 991 1930 995 1934
rect 1095 1930 1099 1934
rect 1135 1902 1139 1906
rect 1231 1902 1235 1906
rect 1271 1902 1275 1906
rect 1319 1902 1323 1906
rect 1359 1902 1363 1906
rect 1375 1902 1379 1906
rect 1423 1902 1427 1906
rect 1439 1902 1443 1906
rect 1487 1902 1491 1906
rect 1503 1902 1507 1906
rect 1559 1902 1563 1906
rect 1575 1902 1579 1906
rect 1631 1902 1635 1906
rect 1655 1902 1659 1906
rect 1703 1902 1707 1906
rect 1751 1902 1755 1906
rect 1775 1902 1779 1906
rect 1847 1902 1851 1906
rect 1863 1902 1867 1906
rect 1927 1902 1931 1906
rect 1975 1902 1979 1906
rect 2007 1902 2011 1906
rect 2071 1902 2075 1906
rect 2119 1902 2123 1906
rect 111 1874 115 1878
rect 135 1874 139 1878
rect 175 1874 179 1878
rect 223 1874 227 1878
rect 231 1874 235 1878
rect 287 1874 291 1878
rect 295 1874 299 1878
rect 359 1874 363 1878
rect 367 1874 371 1878
rect 431 1874 435 1878
rect 447 1874 451 1878
rect 503 1874 507 1878
rect 527 1874 531 1878
rect 567 1874 571 1878
rect 615 1874 619 1878
rect 631 1874 635 1878
rect 695 1874 699 1878
rect 703 1874 707 1878
rect 759 1874 763 1878
rect 791 1874 795 1878
rect 831 1874 835 1878
rect 879 1874 883 1878
rect 1095 1874 1099 1878
rect 1135 1846 1139 1850
rect 1159 1846 1163 1850
rect 1199 1846 1203 1850
rect 1231 1846 1235 1850
rect 1239 1846 1243 1850
rect 1271 1846 1275 1850
rect 1303 1846 1307 1850
rect 1319 1846 1323 1850
rect 1367 1846 1371 1850
rect 1375 1846 1379 1850
rect 1431 1846 1435 1850
rect 1439 1846 1443 1850
rect 1503 1846 1507 1850
rect 1575 1846 1579 1850
rect 1583 1846 1587 1850
rect 1655 1846 1659 1850
rect 1671 1846 1675 1850
rect 1751 1846 1755 1850
rect 1767 1846 1771 1850
rect 1863 1846 1867 1850
rect 1871 1846 1875 1850
rect 1975 1846 1979 1850
rect 1983 1846 1987 1850
rect 2071 1846 2075 1850
rect 2119 1846 2123 1850
rect 111 1818 115 1822
rect 135 1818 139 1822
rect 175 1818 179 1822
rect 183 1818 187 1822
rect 223 1818 227 1822
rect 263 1818 267 1822
rect 287 1818 291 1822
rect 351 1818 355 1822
rect 359 1818 363 1822
rect 431 1818 435 1822
rect 439 1818 443 1822
rect 503 1818 507 1822
rect 527 1818 531 1822
rect 567 1818 571 1822
rect 607 1818 611 1822
rect 631 1818 635 1822
rect 687 1818 691 1822
rect 695 1818 699 1822
rect 759 1818 763 1822
rect 767 1818 771 1822
rect 831 1818 835 1822
rect 839 1818 843 1822
rect 911 1818 915 1822
rect 991 1818 995 1822
rect 1047 1818 1051 1822
rect 1095 1818 1099 1822
rect 1135 1786 1139 1790
rect 1159 1786 1163 1790
rect 1199 1786 1203 1790
rect 1239 1786 1243 1790
rect 1303 1786 1307 1790
rect 1311 1786 1315 1790
rect 1351 1786 1355 1790
rect 1367 1786 1371 1790
rect 1391 1786 1395 1790
rect 1431 1786 1435 1790
rect 1471 1786 1475 1790
rect 1503 1786 1507 1790
rect 1511 1786 1515 1790
rect 1551 1786 1555 1790
rect 1583 1786 1587 1790
rect 1607 1786 1611 1790
rect 1671 1786 1675 1790
rect 1679 1786 1683 1790
rect 1767 1786 1771 1790
rect 1871 1786 1875 1790
rect 1983 1786 1987 1790
rect 2071 1786 2075 1790
rect 2119 1786 2123 1790
rect 111 1758 115 1762
rect 135 1758 139 1762
rect 183 1758 187 1762
rect 199 1758 203 1762
rect 263 1758 267 1762
rect 295 1758 299 1762
rect 351 1758 355 1762
rect 399 1758 403 1762
rect 439 1758 443 1762
rect 495 1758 499 1762
rect 527 1758 531 1762
rect 591 1758 595 1762
rect 607 1758 611 1762
rect 671 1758 675 1762
rect 687 1758 691 1762
rect 751 1758 755 1762
rect 767 1758 771 1762
rect 823 1758 827 1762
rect 839 1758 843 1762
rect 887 1758 891 1762
rect 911 1758 915 1762
rect 959 1758 963 1762
rect 991 1758 995 1762
rect 1031 1758 1035 1762
rect 1047 1758 1051 1762
rect 1095 1758 1099 1762
rect 1135 1730 1139 1734
rect 1263 1730 1267 1734
rect 1311 1730 1315 1734
rect 1319 1730 1323 1734
rect 1351 1730 1355 1734
rect 1383 1730 1387 1734
rect 1391 1730 1395 1734
rect 1431 1730 1435 1734
rect 1455 1730 1459 1734
rect 1471 1730 1475 1734
rect 1511 1730 1515 1734
rect 1535 1730 1539 1734
rect 1551 1730 1555 1734
rect 1607 1730 1611 1734
rect 1615 1730 1619 1734
rect 1679 1730 1683 1734
rect 1687 1730 1691 1734
rect 1759 1730 1763 1734
rect 1767 1730 1771 1734
rect 1831 1730 1835 1734
rect 1871 1730 1875 1734
rect 1895 1730 1899 1734
rect 1959 1730 1963 1734
rect 1983 1730 1987 1734
rect 2023 1730 2027 1734
rect 2071 1730 2075 1734
rect 2119 1730 2123 1734
rect 111 1702 115 1706
rect 135 1702 139 1706
rect 151 1702 155 1706
rect 199 1702 203 1706
rect 223 1702 227 1706
rect 295 1702 299 1706
rect 303 1702 307 1706
rect 383 1702 387 1706
rect 399 1702 403 1706
rect 463 1702 467 1706
rect 495 1702 499 1706
rect 535 1702 539 1706
rect 591 1702 595 1706
rect 607 1702 611 1706
rect 671 1702 675 1706
rect 735 1702 739 1706
rect 751 1702 755 1706
rect 807 1702 811 1706
rect 823 1702 827 1706
rect 879 1702 883 1706
rect 887 1702 891 1706
rect 959 1702 963 1706
rect 1031 1702 1035 1706
rect 1095 1702 1099 1706
rect 1135 1678 1139 1682
rect 1167 1678 1171 1682
rect 1247 1678 1251 1682
rect 1263 1678 1267 1682
rect 1319 1678 1323 1682
rect 1335 1678 1339 1682
rect 1383 1678 1387 1682
rect 1423 1678 1427 1682
rect 1455 1678 1459 1682
rect 1511 1678 1515 1682
rect 1535 1678 1539 1682
rect 1599 1678 1603 1682
rect 1615 1678 1619 1682
rect 1679 1678 1683 1682
rect 1687 1678 1691 1682
rect 1751 1678 1755 1682
rect 1759 1678 1763 1682
rect 1815 1678 1819 1682
rect 1831 1678 1835 1682
rect 1871 1678 1875 1682
rect 1895 1678 1899 1682
rect 1927 1678 1931 1682
rect 1959 1678 1963 1682
rect 1983 1678 1987 1682
rect 2023 1678 2027 1682
rect 2031 1678 2035 1682
rect 2071 1678 2075 1682
rect 2119 1678 2123 1682
rect 111 1646 115 1650
rect 151 1646 155 1650
rect 175 1646 179 1650
rect 215 1646 219 1650
rect 223 1646 227 1650
rect 255 1646 259 1650
rect 303 1646 307 1650
rect 359 1646 363 1650
rect 383 1646 387 1650
rect 407 1646 411 1650
rect 455 1646 459 1650
rect 463 1646 467 1650
rect 503 1646 507 1650
rect 535 1646 539 1650
rect 551 1646 555 1650
rect 607 1646 611 1650
rect 663 1646 667 1650
rect 671 1646 675 1650
rect 719 1646 723 1650
rect 735 1646 739 1650
rect 807 1646 811 1650
rect 879 1646 883 1650
rect 1095 1646 1099 1650
rect 1135 1622 1139 1626
rect 1159 1622 1163 1626
rect 1167 1622 1171 1626
rect 1199 1622 1203 1626
rect 1247 1622 1251 1626
rect 1319 1622 1323 1626
rect 1335 1622 1339 1626
rect 1391 1622 1395 1626
rect 1423 1622 1427 1626
rect 1463 1622 1467 1626
rect 1511 1622 1515 1626
rect 1535 1622 1539 1626
rect 1599 1622 1603 1626
rect 1607 1622 1611 1626
rect 1679 1622 1683 1626
rect 1751 1622 1755 1626
rect 1815 1622 1819 1626
rect 1831 1622 1835 1626
rect 1871 1622 1875 1626
rect 1927 1622 1931 1626
rect 1983 1622 1987 1626
rect 2031 1622 2035 1626
rect 2071 1622 2075 1626
rect 2119 1622 2123 1626
rect 111 1586 115 1590
rect 143 1586 147 1590
rect 175 1586 179 1590
rect 183 1586 187 1590
rect 215 1586 219 1590
rect 231 1586 235 1590
rect 255 1586 259 1590
rect 287 1586 291 1590
rect 303 1586 307 1590
rect 351 1586 355 1590
rect 359 1586 363 1590
rect 407 1586 411 1590
rect 415 1586 419 1590
rect 455 1586 459 1590
rect 479 1586 483 1590
rect 503 1586 507 1590
rect 543 1586 547 1590
rect 551 1586 555 1590
rect 607 1586 611 1590
rect 663 1586 667 1590
rect 719 1586 723 1590
rect 727 1586 731 1590
rect 791 1586 795 1590
rect 855 1586 859 1590
rect 1095 1586 1099 1590
rect 1135 1570 1139 1574
rect 1159 1570 1163 1574
rect 1199 1570 1203 1574
rect 1239 1570 1243 1574
rect 1247 1570 1251 1574
rect 1279 1570 1283 1574
rect 1319 1570 1323 1574
rect 1327 1570 1331 1574
rect 1375 1570 1379 1574
rect 1391 1570 1395 1574
rect 1423 1570 1427 1574
rect 1463 1570 1467 1574
rect 1471 1570 1475 1574
rect 1519 1570 1523 1574
rect 1535 1570 1539 1574
rect 1567 1570 1571 1574
rect 1607 1570 1611 1574
rect 1623 1570 1627 1574
rect 1679 1570 1683 1574
rect 1735 1570 1739 1574
rect 1751 1570 1755 1574
rect 1831 1570 1835 1574
rect 2119 1570 2123 1574
rect 111 1526 115 1530
rect 135 1526 139 1530
rect 143 1526 147 1530
rect 175 1526 179 1530
rect 183 1526 187 1530
rect 215 1526 219 1530
rect 231 1526 235 1530
rect 255 1526 259 1530
rect 287 1526 291 1530
rect 295 1526 299 1530
rect 335 1526 339 1530
rect 351 1526 355 1530
rect 375 1526 379 1530
rect 415 1526 419 1530
rect 455 1526 459 1530
rect 479 1526 483 1530
rect 495 1526 499 1530
rect 535 1526 539 1530
rect 543 1526 547 1530
rect 575 1526 579 1530
rect 607 1526 611 1530
rect 615 1526 619 1530
rect 655 1526 659 1530
rect 663 1526 667 1530
rect 695 1526 699 1530
rect 727 1526 731 1530
rect 735 1526 739 1530
rect 775 1526 779 1530
rect 791 1526 795 1530
rect 831 1526 835 1530
rect 855 1526 859 1530
rect 887 1526 891 1530
rect 1095 1526 1099 1530
rect 1135 1514 1139 1518
rect 1239 1514 1243 1518
rect 1279 1514 1283 1518
rect 1319 1514 1323 1518
rect 1327 1514 1331 1518
rect 1359 1514 1363 1518
rect 1375 1514 1379 1518
rect 1399 1514 1403 1518
rect 1423 1514 1427 1518
rect 1439 1514 1443 1518
rect 1471 1514 1475 1518
rect 1479 1514 1483 1518
rect 1519 1514 1523 1518
rect 1559 1514 1563 1518
rect 1567 1514 1571 1518
rect 1607 1514 1611 1518
rect 1623 1514 1627 1518
rect 1663 1514 1667 1518
rect 1679 1514 1683 1518
rect 1735 1514 1739 1518
rect 1815 1514 1819 1518
rect 1903 1514 1907 1518
rect 1991 1514 1995 1518
rect 2071 1514 2075 1518
rect 2119 1514 2123 1518
rect 111 1466 115 1470
rect 135 1466 139 1470
rect 175 1466 179 1470
rect 215 1466 219 1470
rect 255 1466 259 1470
rect 295 1466 299 1470
rect 335 1466 339 1470
rect 375 1466 379 1470
rect 415 1466 419 1470
rect 455 1466 459 1470
rect 495 1466 499 1470
rect 519 1466 523 1470
rect 535 1466 539 1470
rect 559 1466 563 1470
rect 575 1466 579 1470
rect 599 1466 603 1470
rect 615 1466 619 1470
rect 647 1466 651 1470
rect 655 1466 659 1470
rect 695 1466 699 1470
rect 735 1466 739 1470
rect 751 1466 755 1470
rect 775 1466 779 1470
rect 807 1466 811 1470
rect 831 1466 835 1470
rect 871 1466 875 1470
rect 887 1466 891 1470
rect 935 1466 939 1470
rect 1095 1466 1099 1470
rect 1135 1462 1139 1466
rect 1231 1462 1235 1466
rect 1279 1462 1283 1466
rect 1319 1462 1323 1466
rect 1335 1462 1339 1466
rect 1359 1462 1363 1466
rect 1391 1462 1395 1466
rect 1399 1462 1403 1466
rect 1439 1462 1443 1466
rect 1455 1462 1459 1466
rect 1479 1462 1483 1466
rect 1519 1462 1523 1466
rect 1559 1462 1563 1466
rect 1583 1462 1587 1466
rect 1607 1462 1611 1466
rect 1647 1462 1651 1466
rect 1663 1462 1667 1466
rect 1719 1462 1723 1466
rect 1735 1462 1739 1466
rect 1807 1462 1811 1466
rect 1815 1462 1819 1466
rect 1895 1462 1899 1466
rect 1903 1462 1907 1466
rect 1991 1462 1995 1466
rect 2071 1462 2075 1466
rect 2119 1462 2123 1466
rect 111 1410 115 1414
rect 431 1410 435 1414
rect 471 1410 475 1414
rect 519 1410 523 1414
rect 559 1410 563 1414
rect 575 1410 579 1414
rect 599 1410 603 1414
rect 631 1410 635 1414
rect 647 1410 651 1414
rect 695 1410 699 1414
rect 751 1410 755 1414
rect 759 1410 763 1414
rect 807 1410 811 1414
rect 823 1410 827 1414
rect 871 1410 875 1414
rect 895 1410 899 1414
rect 935 1410 939 1414
rect 967 1410 971 1414
rect 1095 1410 1099 1414
rect 1135 1406 1139 1410
rect 1159 1406 1163 1410
rect 1199 1406 1203 1410
rect 1231 1406 1235 1410
rect 1263 1406 1267 1410
rect 1279 1406 1283 1410
rect 1335 1406 1339 1410
rect 1351 1406 1355 1410
rect 1391 1406 1395 1410
rect 1447 1406 1451 1410
rect 1455 1406 1459 1410
rect 1519 1406 1523 1410
rect 1543 1406 1547 1410
rect 1583 1406 1587 1410
rect 1631 1406 1635 1410
rect 1647 1406 1651 1410
rect 1719 1406 1723 1410
rect 1799 1406 1803 1410
rect 1807 1406 1811 1410
rect 1871 1406 1875 1410
rect 1895 1406 1899 1410
rect 1943 1406 1947 1410
rect 1991 1406 1995 1410
rect 2015 1406 2019 1410
rect 2071 1406 2075 1410
rect 2119 1406 2123 1410
rect 111 1358 115 1362
rect 375 1358 379 1362
rect 423 1358 427 1362
rect 431 1358 435 1362
rect 471 1358 475 1362
rect 479 1358 483 1362
rect 519 1358 523 1362
rect 543 1358 547 1362
rect 575 1358 579 1362
rect 607 1358 611 1362
rect 631 1358 635 1362
rect 671 1358 675 1362
rect 695 1358 699 1362
rect 735 1358 739 1362
rect 759 1358 763 1362
rect 799 1358 803 1362
rect 823 1358 827 1362
rect 863 1358 867 1362
rect 895 1358 899 1362
rect 927 1358 931 1362
rect 967 1358 971 1362
rect 999 1358 1003 1362
rect 1047 1358 1051 1362
rect 1095 1358 1099 1362
rect 1135 1350 1139 1354
rect 1159 1350 1163 1354
rect 1199 1350 1203 1354
rect 1255 1350 1259 1354
rect 1263 1350 1267 1354
rect 1351 1350 1355 1354
rect 1375 1350 1379 1354
rect 1447 1350 1451 1354
rect 1487 1350 1491 1354
rect 1543 1350 1547 1354
rect 1591 1350 1595 1354
rect 1631 1350 1635 1354
rect 1679 1350 1683 1354
rect 1719 1350 1723 1354
rect 1759 1350 1763 1354
rect 1799 1350 1803 1354
rect 1831 1350 1835 1354
rect 1871 1350 1875 1354
rect 1903 1350 1907 1354
rect 1943 1350 1947 1354
rect 1967 1350 1971 1354
rect 2015 1350 2019 1354
rect 2031 1350 2035 1354
rect 2071 1350 2075 1354
rect 2119 1350 2123 1354
rect 111 1306 115 1310
rect 335 1306 339 1310
rect 375 1306 379 1310
rect 391 1306 395 1310
rect 423 1306 427 1310
rect 455 1306 459 1310
rect 479 1306 483 1310
rect 527 1306 531 1310
rect 543 1306 547 1310
rect 599 1306 603 1310
rect 607 1306 611 1310
rect 671 1306 675 1310
rect 735 1306 739 1310
rect 743 1306 747 1310
rect 799 1306 803 1310
rect 823 1306 827 1310
rect 863 1306 867 1310
rect 903 1306 907 1310
rect 927 1306 931 1310
rect 983 1306 987 1310
rect 999 1306 1003 1310
rect 1047 1306 1051 1310
rect 1095 1306 1099 1310
rect 1135 1294 1139 1298
rect 1159 1294 1163 1298
rect 1199 1294 1203 1298
rect 1247 1294 1251 1298
rect 1255 1294 1259 1298
rect 1319 1294 1323 1298
rect 1375 1294 1379 1298
rect 1399 1294 1403 1298
rect 1479 1294 1483 1298
rect 1487 1294 1491 1298
rect 1559 1294 1563 1298
rect 1591 1294 1595 1298
rect 1639 1294 1643 1298
rect 1679 1294 1683 1298
rect 1719 1294 1723 1298
rect 1759 1294 1763 1298
rect 1799 1294 1803 1298
rect 1831 1294 1835 1298
rect 1879 1294 1883 1298
rect 1903 1294 1907 1298
rect 1967 1294 1971 1298
rect 2031 1294 2035 1298
rect 2055 1294 2059 1298
rect 2071 1294 2075 1298
rect 2119 1294 2123 1298
rect 111 1250 115 1254
rect 263 1250 267 1254
rect 311 1250 315 1254
rect 335 1250 339 1254
rect 359 1250 363 1254
rect 391 1250 395 1254
rect 415 1250 419 1254
rect 455 1250 459 1254
rect 479 1250 483 1254
rect 527 1250 531 1254
rect 543 1250 547 1254
rect 599 1250 603 1254
rect 607 1250 611 1254
rect 671 1250 675 1254
rect 735 1250 739 1254
rect 743 1250 747 1254
rect 799 1250 803 1254
rect 823 1250 827 1254
rect 863 1250 867 1254
rect 903 1250 907 1254
rect 927 1250 931 1254
rect 983 1250 987 1254
rect 1047 1250 1051 1254
rect 1095 1250 1099 1254
rect 1135 1238 1139 1242
rect 1159 1238 1163 1242
rect 1199 1238 1203 1242
rect 1239 1238 1243 1242
rect 1247 1238 1251 1242
rect 1279 1238 1283 1242
rect 1319 1238 1323 1242
rect 1327 1238 1331 1242
rect 1375 1238 1379 1242
rect 1399 1238 1403 1242
rect 1423 1238 1427 1242
rect 1471 1238 1475 1242
rect 1479 1238 1483 1242
rect 1535 1238 1539 1242
rect 1559 1238 1563 1242
rect 1615 1238 1619 1242
rect 1639 1238 1643 1242
rect 1719 1238 1723 1242
rect 1799 1238 1803 1242
rect 1839 1238 1843 1242
rect 1879 1238 1883 1242
rect 1967 1238 1971 1242
rect 2055 1238 2059 1242
rect 2071 1238 2075 1242
rect 2119 1238 2123 1242
rect 111 1198 115 1202
rect 223 1198 227 1202
rect 263 1198 267 1202
rect 279 1198 283 1202
rect 311 1198 315 1202
rect 343 1198 347 1202
rect 359 1198 363 1202
rect 407 1198 411 1202
rect 415 1198 419 1202
rect 479 1198 483 1202
rect 543 1198 547 1202
rect 551 1198 555 1202
rect 607 1198 611 1202
rect 631 1198 635 1202
rect 671 1198 675 1202
rect 711 1198 715 1202
rect 735 1198 739 1202
rect 791 1198 795 1202
rect 799 1198 803 1202
rect 863 1198 867 1202
rect 871 1198 875 1202
rect 927 1198 931 1202
rect 959 1198 963 1202
rect 1095 1198 1099 1202
rect 1135 1186 1139 1190
rect 1159 1186 1163 1190
rect 1199 1186 1203 1190
rect 1239 1186 1243 1190
rect 1279 1186 1283 1190
rect 1287 1186 1291 1190
rect 1327 1186 1331 1190
rect 1367 1186 1371 1190
rect 1375 1186 1379 1190
rect 1415 1186 1419 1190
rect 1423 1186 1427 1190
rect 1471 1186 1475 1190
rect 1527 1186 1531 1190
rect 1535 1186 1539 1190
rect 1583 1186 1587 1190
rect 1615 1186 1619 1190
rect 1639 1186 1643 1190
rect 1703 1186 1707 1190
rect 1719 1186 1723 1190
rect 1767 1186 1771 1190
rect 1839 1186 1843 1190
rect 1919 1186 1923 1190
rect 1967 1186 1971 1190
rect 2007 1186 2011 1190
rect 2071 1186 2075 1190
rect 2119 1186 2123 1190
rect 111 1146 115 1150
rect 159 1146 163 1150
rect 199 1146 203 1150
rect 223 1146 227 1150
rect 247 1146 251 1150
rect 279 1146 283 1150
rect 303 1146 307 1150
rect 343 1146 347 1150
rect 367 1146 371 1150
rect 407 1146 411 1150
rect 439 1146 443 1150
rect 479 1146 483 1150
rect 511 1146 515 1150
rect 551 1146 555 1150
rect 591 1146 595 1150
rect 631 1146 635 1150
rect 679 1146 683 1150
rect 711 1146 715 1150
rect 775 1146 779 1150
rect 791 1146 795 1150
rect 871 1146 875 1150
rect 879 1146 883 1150
rect 959 1146 963 1150
rect 991 1146 995 1150
rect 1095 1146 1099 1150
rect 1135 1126 1139 1130
rect 1287 1126 1291 1130
rect 1327 1126 1331 1130
rect 1367 1126 1371 1130
rect 1383 1126 1387 1130
rect 1415 1126 1419 1130
rect 1423 1126 1427 1130
rect 1471 1126 1475 1130
rect 1527 1126 1531 1130
rect 1583 1126 1587 1130
rect 1591 1126 1595 1130
rect 1639 1126 1643 1130
rect 1655 1126 1659 1130
rect 1703 1126 1707 1130
rect 1711 1126 1715 1130
rect 1767 1126 1771 1130
rect 1823 1126 1827 1130
rect 1839 1126 1843 1130
rect 1871 1126 1875 1130
rect 1919 1126 1923 1130
rect 1927 1126 1931 1130
rect 1983 1126 1987 1130
rect 2007 1126 2011 1130
rect 2031 1126 2035 1130
rect 2071 1126 2075 1130
rect 2119 1126 2123 1130
rect 111 1086 115 1090
rect 159 1086 163 1090
rect 199 1086 203 1090
rect 247 1086 251 1090
rect 303 1086 307 1090
rect 367 1086 371 1090
rect 431 1086 435 1090
rect 439 1086 443 1090
rect 503 1086 507 1090
rect 511 1086 515 1090
rect 575 1086 579 1090
rect 591 1086 595 1090
rect 647 1086 651 1090
rect 679 1086 683 1090
rect 719 1086 723 1090
rect 775 1086 779 1090
rect 783 1086 787 1090
rect 839 1086 843 1090
rect 879 1086 883 1090
rect 895 1086 899 1090
rect 951 1086 955 1090
rect 991 1086 995 1090
rect 1007 1086 1011 1090
rect 1047 1086 1051 1090
rect 1095 1086 1099 1090
rect 1135 1074 1139 1078
rect 1159 1074 1163 1078
rect 1247 1074 1251 1078
rect 1359 1074 1363 1078
rect 1383 1074 1387 1078
rect 1423 1074 1427 1078
rect 1471 1074 1475 1078
rect 1527 1074 1531 1078
rect 1575 1074 1579 1078
rect 1591 1074 1595 1078
rect 1655 1074 1659 1078
rect 1671 1074 1675 1078
rect 1711 1074 1715 1078
rect 1759 1074 1763 1078
rect 1767 1074 1771 1078
rect 1823 1074 1827 1078
rect 1847 1074 1851 1078
rect 1871 1074 1875 1078
rect 1927 1074 1931 1078
rect 1983 1074 1987 1078
rect 2007 1074 2011 1078
rect 2031 1074 2035 1078
rect 2071 1074 2075 1078
rect 2119 1074 2123 1078
rect 111 1030 115 1034
rect 199 1030 203 1034
rect 223 1030 227 1034
rect 247 1030 251 1034
rect 271 1030 275 1034
rect 303 1030 307 1034
rect 335 1030 339 1034
rect 367 1030 371 1034
rect 407 1030 411 1034
rect 431 1030 435 1034
rect 479 1030 483 1034
rect 503 1030 507 1034
rect 559 1030 563 1034
rect 575 1030 579 1034
rect 631 1030 635 1034
rect 647 1030 651 1034
rect 703 1030 707 1034
rect 719 1030 723 1034
rect 775 1030 779 1034
rect 783 1030 787 1034
rect 839 1030 843 1034
rect 895 1030 899 1034
rect 903 1030 907 1034
rect 951 1030 955 1034
rect 967 1030 971 1034
rect 1007 1030 1011 1034
rect 1039 1030 1043 1034
rect 1047 1030 1051 1034
rect 1095 1030 1099 1034
rect 1135 1022 1139 1026
rect 1159 1022 1163 1026
rect 1231 1022 1235 1026
rect 1247 1022 1251 1026
rect 1303 1022 1307 1026
rect 1359 1022 1363 1026
rect 1383 1022 1387 1026
rect 1463 1022 1467 1026
rect 1471 1022 1475 1026
rect 1543 1022 1547 1026
rect 1575 1022 1579 1026
rect 1623 1022 1627 1026
rect 1671 1022 1675 1026
rect 1695 1022 1699 1026
rect 1759 1022 1763 1026
rect 1823 1022 1827 1026
rect 1847 1022 1851 1026
rect 1887 1022 1891 1026
rect 1927 1022 1931 1026
rect 1951 1022 1955 1026
rect 2007 1022 2011 1026
rect 2071 1022 2075 1026
rect 2119 1022 2123 1026
rect 111 974 115 978
rect 151 974 155 978
rect 215 974 219 978
rect 223 974 227 978
rect 271 974 275 978
rect 287 974 291 978
rect 335 974 339 978
rect 367 974 371 978
rect 407 974 411 978
rect 447 974 451 978
rect 479 974 483 978
rect 527 974 531 978
rect 559 974 563 978
rect 599 974 603 978
rect 631 974 635 978
rect 671 974 675 978
rect 703 974 707 978
rect 735 974 739 978
rect 775 974 779 978
rect 799 974 803 978
rect 839 974 843 978
rect 863 974 867 978
rect 903 974 907 978
rect 927 974 931 978
rect 967 974 971 978
rect 991 974 995 978
rect 1039 974 1043 978
rect 1047 974 1051 978
rect 1095 974 1099 978
rect 1135 970 1139 974
rect 1159 970 1163 974
rect 1231 970 1235 974
rect 1239 970 1243 974
rect 1303 970 1307 974
rect 1375 970 1379 974
rect 1383 970 1387 974
rect 1439 970 1443 974
rect 1463 970 1467 974
rect 1511 970 1515 974
rect 1543 970 1547 974
rect 1583 970 1587 974
rect 1623 970 1627 974
rect 1655 970 1659 974
rect 1695 970 1699 974
rect 1727 970 1731 974
rect 1759 970 1763 974
rect 1799 970 1803 974
rect 1823 970 1827 974
rect 1871 970 1875 974
rect 1887 970 1891 974
rect 1943 970 1947 974
rect 1951 970 1955 974
rect 2015 970 2019 974
rect 2071 970 2075 974
rect 2119 970 2123 974
rect 111 922 115 926
rect 135 922 139 926
rect 151 922 155 926
rect 183 922 187 926
rect 215 922 219 926
rect 255 922 259 926
rect 287 922 291 926
rect 327 922 331 926
rect 367 922 371 926
rect 399 922 403 926
rect 447 922 451 926
rect 463 922 467 926
rect 527 922 531 926
rect 599 922 603 926
rect 671 922 675 926
rect 735 922 739 926
rect 743 922 747 926
rect 799 922 803 926
rect 815 922 819 926
rect 863 922 867 926
rect 895 922 899 926
rect 927 922 931 926
rect 983 922 987 926
rect 991 922 995 926
rect 1047 922 1051 926
rect 1095 922 1099 926
rect 1135 914 1139 918
rect 1239 914 1243 918
rect 1287 914 1291 918
rect 1303 914 1307 918
rect 1327 914 1331 918
rect 1375 914 1379 918
rect 1423 914 1427 918
rect 1439 914 1443 918
rect 1479 914 1483 918
rect 1511 914 1515 918
rect 1551 914 1555 918
rect 1583 914 1587 918
rect 1623 914 1627 918
rect 1655 914 1659 918
rect 1703 914 1707 918
rect 1727 914 1731 918
rect 1791 914 1795 918
rect 1799 914 1803 918
rect 1871 914 1875 918
rect 1879 914 1883 918
rect 1943 914 1947 918
rect 1967 914 1971 918
rect 2015 914 2019 918
rect 2063 914 2067 918
rect 2071 914 2075 918
rect 2119 914 2123 918
rect 111 866 115 870
rect 135 866 139 870
rect 175 866 179 870
rect 183 866 187 870
rect 215 866 219 870
rect 255 866 259 870
rect 279 866 283 870
rect 327 866 331 870
rect 343 866 347 870
rect 399 866 403 870
rect 463 866 467 870
rect 527 866 531 870
rect 535 866 539 870
rect 599 866 603 870
rect 615 866 619 870
rect 671 866 675 870
rect 711 866 715 870
rect 743 866 747 870
rect 815 866 819 870
rect 823 866 827 870
rect 895 866 899 870
rect 943 866 947 870
rect 983 866 987 870
rect 1047 866 1051 870
rect 1095 866 1099 870
rect 1135 862 1139 866
rect 1159 862 1163 866
rect 1199 862 1203 866
rect 1263 862 1267 866
rect 1287 862 1291 866
rect 1327 862 1331 866
rect 1375 862 1379 866
rect 1399 862 1403 866
rect 1423 862 1427 866
rect 1471 862 1475 866
rect 1479 862 1483 866
rect 1543 862 1547 866
rect 1551 862 1555 866
rect 1623 862 1627 866
rect 1703 862 1707 866
rect 1775 862 1779 866
rect 1791 862 1795 866
rect 1855 862 1859 866
rect 1879 862 1883 866
rect 1935 862 1939 866
rect 1967 862 1971 866
rect 2015 862 2019 866
rect 2063 862 2067 866
rect 2071 862 2075 866
rect 2119 862 2123 866
rect 111 814 115 818
rect 135 814 139 818
rect 175 814 179 818
rect 215 814 219 818
rect 279 814 283 818
rect 335 814 339 818
rect 343 814 347 818
rect 391 814 395 818
rect 399 814 403 818
rect 455 814 459 818
rect 463 814 467 818
rect 519 814 523 818
rect 535 814 539 818
rect 583 814 587 818
rect 615 814 619 818
rect 655 814 659 818
rect 711 814 715 818
rect 735 814 739 818
rect 815 814 819 818
rect 823 814 827 818
rect 895 814 899 818
rect 943 814 947 818
rect 983 814 987 818
rect 1047 814 1051 818
rect 1095 814 1099 818
rect 1135 802 1139 806
rect 1159 802 1163 806
rect 1199 802 1203 806
rect 1239 802 1243 806
rect 1263 802 1267 806
rect 1327 802 1331 806
rect 1343 802 1347 806
rect 1399 802 1403 806
rect 1447 802 1451 806
rect 1471 802 1475 806
rect 1543 802 1547 806
rect 1551 802 1555 806
rect 1623 802 1627 806
rect 1655 802 1659 806
rect 1703 802 1707 806
rect 1751 802 1755 806
rect 1775 802 1779 806
rect 1839 802 1843 806
rect 1855 802 1859 806
rect 1919 802 1923 806
rect 1935 802 1939 806
rect 2007 802 2011 806
rect 2015 802 2019 806
rect 2071 802 2075 806
rect 2119 802 2123 806
rect 111 762 115 766
rect 135 762 139 766
rect 175 762 179 766
rect 207 762 211 766
rect 215 762 219 766
rect 279 762 283 766
rect 295 762 299 766
rect 335 762 339 766
rect 375 762 379 766
rect 391 762 395 766
rect 447 762 451 766
rect 455 762 459 766
rect 519 762 523 766
rect 583 762 587 766
rect 639 762 643 766
rect 655 762 659 766
rect 687 762 691 766
rect 735 762 739 766
rect 743 762 747 766
rect 799 762 803 766
rect 815 762 819 766
rect 855 762 859 766
rect 895 762 899 766
rect 983 762 987 766
rect 1047 762 1051 766
rect 1095 762 1099 766
rect 1135 750 1139 754
rect 1159 750 1163 754
rect 1199 750 1203 754
rect 1239 750 1243 754
rect 1287 750 1291 754
rect 1343 750 1347 754
rect 1359 750 1363 754
rect 1439 750 1443 754
rect 1447 750 1451 754
rect 1527 750 1531 754
rect 1551 750 1555 754
rect 1615 750 1619 754
rect 1655 750 1659 754
rect 1711 750 1715 754
rect 1751 750 1755 754
rect 1807 750 1811 754
rect 1839 750 1843 754
rect 1903 750 1907 754
rect 1919 750 1923 754
rect 1999 750 2003 754
rect 2007 750 2011 754
rect 2071 750 2075 754
rect 2119 750 2123 754
rect 111 706 115 710
rect 135 706 139 710
rect 183 706 187 710
rect 207 706 211 710
rect 247 706 251 710
rect 295 706 299 710
rect 311 706 315 710
rect 375 706 379 710
rect 383 706 387 710
rect 447 706 451 710
rect 455 706 459 710
rect 519 706 523 710
rect 583 706 587 710
rect 639 706 643 710
rect 647 706 651 710
rect 687 706 691 710
rect 711 706 715 710
rect 743 706 747 710
rect 767 706 771 710
rect 799 706 803 710
rect 823 706 827 710
rect 855 706 859 710
rect 879 706 883 710
rect 943 706 947 710
rect 1095 706 1099 710
rect 1135 694 1139 698
rect 1159 694 1163 698
rect 1199 694 1203 698
rect 1239 694 1243 698
rect 1287 694 1291 698
rect 1335 694 1339 698
rect 1359 694 1363 698
rect 1391 694 1395 698
rect 1439 694 1443 698
rect 1447 694 1451 698
rect 1511 694 1515 698
rect 1527 694 1531 698
rect 1575 694 1579 698
rect 1615 694 1619 698
rect 1639 694 1643 698
rect 1703 694 1707 698
rect 1711 694 1715 698
rect 1767 694 1771 698
rect 1807 694 1811 698
rect 1831 694 1835 698
rect 1895 694 1899 698
rect 1903 694 1907 698
rect 1959 694 1963 698
rect 1999 694 2003 698
rect 2023 694 2027 698
rect 2071 694 2075 698
rect 2119 694 2123 698
rect 111 646 115 650
rect 135 646 139 650
rect 159 646 163 650
rect 183 646 187 650
rect 215 646 219 650
rect 247 646 251 650
rect 287 646 291 650
rect 311 646 315 650
rect 367 646 371 650
rect 383 646 387 650
rect 455 646 459 650
rect 519 646 523 650
rect 543 646 547 650
rect 583 646 587 650
rect 631 646 635 650
rect 647 646 651 650
rect 711 646 715 650
rect 719 646 723 650
rect 767 646 771 650
rect 799 646 803 650
rect 823 646 827 650
rect 871 646 875 650
rect 879 646 883 650
rect 943 646 947 650
rect 951 646 955 650
rect 1031 646 1035 650
rect 1095 646 1099 650
rect 1135 642 1139 646
rect 1239 642 1243 646
rect 1279 642 1283 646
rect 1287 642 1291 646
rect 1319 642 1323 646
rect 1335 642 1339 646
rect 1367 642 1371 646
rect 1391 642 1395 646
rect 1423 642 1427 646
rect 1447 642 1451 646
rect 1479 642 1483 646
rect 1511 642 1515 646
rect 1535 642 1539 646
rect 1575 642 1579 646
rect 1591 642 1595 646
rect 1639 642 1643 646
rect 1647 642 1651 646
rect 1703 642 1707 646
rect 1719 642 1723 646
rect 1767 642 1771 646
rect 1799 642 1803 646
rect 1831 642 1835 646
rect 1879 642 1883 646
rect 1895 642 1899 646
rect 1959 642 1963 646
rect 1967 642 1971 646
rect 2023 642 2027 646
rect 2063 642 2067 646
rect 2071 642 2075 646
rect 2119 642 2123 646
rect 111 590 115 594
rect 159 590 163 594
rect 207 590 211 594
rect 215 590 219 594
rect 255 590 259 594
rect 287 590 291 594
rect 311 590 315 594
rect 367 590 371 594
rect 383 590 387 594
rect 455 590 459 594
rect 463 590 467 594
rect 543 590 547 594
rect 623 590 627 594
rect 631 590 635 594
rect 703 590 707 594
rect 719 590 723 594
rect 783 590 787 594
rect 799 590 803 594
rect 855 590 859 594
rect 871 590 875 594
rect 927 590 931 594
rect 951 590 955 594
rect 999 590 1003 594
rect 1031 590 1035 594
rect 1047 590 1051 594
rect 1095 590 1099 594
rect 1135 590 1139 594
rect 1279 590 1283 594
rect 1319 590 1323 594
rect 1335 590 1339 594
rect 1367 590 1371 594
rect 1375 590 1379 594
rect 1415 590 1419 594
rect 1423 590 1427 594
rect 1463 590 1467 594
rect 1479 590 1483 594
rect 1519 590 1523 594
rect 1535 590 1539 594
rect 1583 590 1587 594
rect 1591 590 1595 594
rect 1647 590 1651 594
rect 1655 590 1659 594
rect 1719 590 1723 594
rect 1727 590 1731 594
rect 1799 590 1803 594
rect 1807 590 1811 594
rect 1879 590 1883 594
rect 1887 590 1891 594
rect 1967 590 1971 594
rect 1975 590 1979 594
rect 2063 590 2067 594
rect 2119 590 2123 594
rect 111 530 115 534
rect 159 530 163 534
rect 167 530 171 534
rect 207 530 211 534
rect 223 530 227 534
rect 255 530 259 534
rect 287 530 291 534
rect 311 530 315 534
rect 359 530 363 534
rect 383 530 387 534
rect 431 530 435 534
rect 463 530 467 534
rect 511 530 515 534
rect 543 530 547 534
rect 591 530 595 534
rect 623 530 627 534
rect 663 530 667 534
rect 703 530 707 534
rect 735 530 739 534
rect 783 530 787 534
rect 807 530 811 534
rect 855 530 859 534
rect 871 530 875 534
rect 927 530 931 534
rect 935 530 939 534
rect 999 530 1003 534
rect 1047 530 1051 534
rect 1095 530 1099 534
rect 1135 534 1139 538
rect 1191 534 1195 538
rect 1239 534 1243 538
rect 1287 534 1291 538
rect 1335 534 1339 538
rect 1343 534 1347 538
rect 1375 534 1379 538
rect 1407 534 1411 538
rect 1415 534 1419 538
rect 1463 534 1467 538
rect 1479 534 1483 538
rect 1519 534 1523 538
rect 1543 534 1547 538
rect 1583 534 1587 538
rect 1607 534 1611 538
rect 1655 534 1659 538
rect 1671 534 1675 538
rect 1727 534 1731 538
rect 1735 534 1739 538
rect 1799 534 1803 538
rect 1807 534 1811 538
rect 1863 534 1867 538
rect 1887 534 1891 538
rect 1935 534 1939 538
rect 1975 534 1979 538
rect 2007 534 2011 538
rect 2063 534 2067 538
rect 2071 534 2075 538
rect 2119 534 2123 538
rect 111 478 115 482
rect 167 478 171 482
rect 223 478 227 482
rect 231 478 235 482
rect 287 478 291 482
rect 303 478 307 482
rect 359 478 363 482
rect 375 478 379 482
rect 431 478 435 482
rect 455 478 459 482
rect 511 478 515 482
rect 535 478 539 482
rect 591 478 595 482
rect 607 478 611 482
rect 663 478 667 482
rect 679 478 683 482
rect 735 478 739 482
rect 743 478 747 482
rect 799 478 803 482
rect 807 478 811 482
rect 855 478 859 482
rect 871 478 875 482
rect 903 478 907 482
rect 935 478 939 482
rect 959 478 963 482
rect 999 478 1003 482
rect 1007 478 1011 482
rect 1047 478 1051 482
rect 1095 478 1099 482
rect 1135 482 1139 486
rect 1159 482 1163 486
rect 1191 482 1195 486
rect 1239 482 1243 486
rect 1263 482 1267 486
rect 1287 482 1291 486
rect 1343 482 1347 486
rect 1383 482 1387 486
rect 1407 482 1411 486
rect 1479 482 1483 486
rect 1495 482 1499 486
rect 1543 482 1547 486
rect 1599 482 1603 486
rect 1607 482 1611 486
rect 1671 482 1675 486
rect 1703 482 1707 486
rect 1735 482 1739 486
rect 1799 482 1803 486
rect 1863 482 1867 486
rect 1887 482 1891 486
rect 1935 482 1939 486
rect 1983 482 1987 486
rect 2007 482 2011 486
rect 2071 482 2075 486
rect 2119 482 2123 486
rect 111 426 115 430
rect 151 426 155 430
rect 167 426 171 430
rect 215 426 219 430
rect 231 426 235 430
rect 279 426 283 430
rect 303 426 307 430
rect 351 426 355 430
rect 375 426 379 430
rect 423 426 427 430
rect 455 426 459 430
rect 487 426 491 430
rect 535 426 539 430
rect 551 426 555 430
rect 607 426 611 430
rect 615 426 619 430
rect 671 426 675 430
rect 679 426 683 430
rect 727 426 731 430
rect 743 426 747 430
rect 791 426 795 430
rect 799 426 803 430
rect 855 426 859 430
rect 903 426 907 430
rect 959 426 963 430
rect 1007 426 1011 430
rect 1047 426 1051 430
rect 1095 426 1099 430
rect 1135 430 1139 434
rect 1159 430 1163 434
rect 1199 430 1203 434
rect 1255 430 1259 434
rect 1263 430 1267 434
rect 1335 430 1339 434
rect 1383 430 1387 434
rect 1415 430 1419 434
rect 1495 430 1499 434
rect 1503 430 1507 434
rect 1591 430 1595 434
rect 1599 430 1603 434
rect 1671 430 1675 434
rect 1703 430 1707 434
rect 1751 430 1755 434
rect 1799 430 1803 434
rect 1823 430 1827 434
rect 1887 430 1891 434
rect 1951 430 1955 434
rect 1983 430 1987 434
rect 2023 430 2027 434
rect 2071 430 2075 434
rect 2119 430 2123 434
rect 111 374 115 378
rect 135 374 139 378
rect 151 374 155 378
rect 175 374 179 378
rect 215 374 219 378
rect 271 374 275 378
rect 279 374 283 378
rect 335 374 339 378
rect 351 374 355 378
rect 399 374 403 378
rect 423 374 427 378
rect 463 374 467 378
rect 487 374 491 378
rect 519 374 523 378
rect 551 374 555 378
rect 575 374 579 378
rect 615 374 619 378
rect 631 374 635 378
rect 671 374 675 378
rect 687 374 691 378
rect 727 374 731 378
rect 751 374 755 378
rect 791 374 795 378
rect 855 374 859 378
rect 1095 374 1099 378
rect 1135 374 1139 378
rect 1159 374 1163 378
rect 1199 374 1203 378
rect 1255 374 1259 378
rect 1303 374 1307 378
rect 1335 374 1339 378
rect 1343 374 1347 378
rect 1383 374 1387 378
rect 1415 374 1419 378
rect 1423 374 1427 378
rect 1463 374 1467 378
rect 1503 374 1507 378
rect 1551 374 1555 378
rect 1591 374 1595 378
rect 1615 374 1619 378
rect 1671 374 1675 378
rect 1679 374 1683 378
rect 1751 374 1755 378
rect 1823 374 1827 378
rect 1831 374 1835 378
rect 1887 374 1891 378
rect 1919 374 1923 378
rect 1951 374 1955 378
rect 2007 374 2011 378
rect 2023 374 2027 378
rect 2071 374 2075 378
rect 2119 374 2123 378
rect 111 318 115 322
rect 135 318 139 322
rect 175 318 179 322
rect 207 318 211 322
rect 215 318 219 322
rect 271 318 275 322
rect 295 318 299 322
rect 335 318 339 322
rect 383 318 387 322
rect 399 318 403 322
rect 463 318 467 322
rect 471 318 475 322
rect 519 318 523 322
rect 551 318 555 322
rect 575 318 579 322
rect 623 318 627 322
rect 631 318 635 322
rect 687 318 691 322
rect 751 318 755 322
rect 807 318 811 322
rect 871 318 875 322
rect 935 318 939 322
rect 1095 318 1099 322
rect 1135 318 1139 322
rect 1167 318 1171 322
rect 1207 318 1211 322
rect 1247 318 1251 322
rect 1295 318 1299 322
rect 1303 318 1307 322
rect 1343 318 1347 322
rect 1383 318 1387 322
rect 1391 318 1395 322
rect 1423 318 1427 322
rect 1439 318 1443 322
rect 1463 318 1467 322
rect 1495 318 1499 322
rect 1503 318 1507 322
rect 1551 318 1555 322
rect 1559 318 1563 322
rect 1615 318 1619 322
rect 1623 318 1627 322
rect 1679 318 1683 322
rect 1695 318 1699 322
rect 1751 318 1755 322
rect 1775 318 1779 322
rect 1831 318 1835 322
rect 1855 318 1859 322
rect 1919 318 1923 322
rect 1935 318 1939 322
rect 2007 318 2011 322
rect 2015 318 2019 322
rect 2071 318 2075 322
rect 2119 318 2123 322
rect 111 266 115 270
rect 135 266 139 270
rect 199 266 203 270
rect 207 266 211 270
rect 279 266 283 270
rect 295 266 299 270
rect 359 266 363 270
rect 383 266 387 270
rect 439 266 443 270
rect 471 266 475 270
rect 511 266 515 270
rect 551 266 555 270
rect 583 266 587 270
rect 623 266 627 270
rect 647 266 651 270
rect 687 266 691 270
rect 703 266 707 270
rect 751 266 755 270
rect 759 266 763 270
rect 807 266 811 270
rect 815 266 819 270
rect 871 266 875 270
rect 879 266 883 270
rect 935 266 939 270
rect 1095 266 1099 270
rect 1135 258 1139 262
rect 1159 258 1163 262
rect 1167 258 1171 262
rect 1207 258 1211 262
rect 1247 258 1251 262
rect 1271 258 1275 262
rect 1295 258 1299 262
rect 1327 258 1331 262
rect 1343 258 1347 262
rect 1391 258 1395 262
rect 1439 258 1443 262
rect 1455 258 1459 262
rect 1495 258 1499 262
rect 1527 258 1531 262
rect 1559 258 1563 262
rect 1607 258 1611 262
rect 1623 258 1627 262
rect 1687 258 1691 262
rect 1695 258 1699 262
rect 1767 258 1771 262
rect 1775 258 1779 262
rect 1839 258 1843 262
rect 1855 258 1859 262
rect 1919 258 1923 262
rect 1935 258 1939 262
rect 1999 258 2003 262
rect 2015 258 2019 262
rect 2071 258 2075 262
rect 2119 258 2123 262
rect 111 210 115 214
rect 135 210 139 214
rect 183 210 187 214
rect 199 210 203 214
rect 231 210 235 214
rect 279 210 283 214
rect 327 210 331 214
rect 359 210 363 214
rect 375 210 379 214
rect 415 210 419 214
rect 439 210 443 214
rect 455 210 459 214
rect 503 210 507 214
rect 511 210 515 214
rect 551 210 555 214
rect 583 210 587 214
rect 599 210 603 214
rect 647 210 651 214
rect 695 210 699 214
rect 703 210 707 214
rect 743 210 747 214
rect 759 210 763 214
rect 815 210 819 214
rect 879 210 883 214
rect 1095 210 1099 214
rect 1135 206 1139 210
rect 1159 206 1163 210
rect 1199 206 1203 210
rect 1207 206 1211 210
rect 1263 206 1267 210
rect 1271 206 1275 210
rect 1327 206 1331 210
rect 1391 206 1395 210
rect 1399 206 1403 210
rect 1455 206 1459 210
rect 1471 206 1475 210
rect 1527 206 1531 210
rect 1543 206 1547 210
rect 1607 206 1611 210
rect 1671 206 1675 210
rect 1687 206 1691 210
rect 1735 206 1739 210
rect 1767 206 1771 210
rect 1807 206 1811 210
rect 1839 206 1843 210
rect 1879 206 1883 210
rect 1919 206 1923 210
rect 1951 206 1955 210
rect 1999 206 2003 210
rect 2023 206 2027 210
rect 2071 206 2075 210
rect 2119 206 2123 210
rect 111 134 115 138
rect 135 134 139 138
rect 143 134 147 138
rect 183 134 187 138
rect 223 134 227 138
rect 231 134 235 138
rect 263 134 267 138
rect 279 134 283 138
rect 303 134 307 138
rect 327 134 331 138
rect 343 134 347 138
rect 375 134 379 138
rect 383 134 387 138
rect 415 134 419 138
rect 423 134 427 138
rect 455 134 459 138
rect 463 134 467 138
rect 503 134 507 138
rect 543 134 547 138
rect 551 134 555 138
rect 583 134 587 138
rect 599 134 603 138
rect 623 134 627 138
rect 647 134 651 138
rect 663 134 667 138
rect 695 134 699 138
rect 703 134 707 138
rect 743 134 747 138
rect 783 134 787 138
rect 831 134 835 138
rect 879 134 883 138
rect 927 134 931 138
rect 967 134 971 138
rect 1007 134 1011 138
rect 1047 134 1051 138
rect 1095 134 1099 138
rect 1135 134 1139 138
rect 1159 134 1163 138
rect 1199 134 1203 138
rect 1207 134 1211 138
rect 1263 134 1267 138
rect 1271 134 1275 138
rect 1327 134 1331 138
rect 1335 134 1339 138
rect 1399 134 1403 138
rect 1455 134 1459 138
rect 1471 134 1475 138
rect 1511 134 1515 138
rect 1543 134 1547 138
rect 1559 134 1563 138
rect 1607 134 1611 138
rect 1647 134 1651 138
rect 1671 134 1675 138
rect 1687 134 1691 138
rect 1727 134 1731 138
rect 1735 134 1739 138
rect 1767 134 1771 138
rect 1807 134 1811 138
rect 1855 134 1859 138
rect 1879 134 1883 138
rect 1903 134 1907 138
rect 1951 134 1955 138
rect 1991 134 1995 138
rect 2023 134 2027 138
rect 2031 134 2035 138
rect 2071 134 2075 138
rect 2119 134 2123 138
rect 111 82 115 86
rect 143 82 147 86
rect 183 82 187 86
rect 223 82 227 86
rect 263 82 267 86
rect 303 82 307 86
rect 343 82 347 86
rect 383 82 387 86
rect 423 82 427 86
rect 463 82 467 86
rect 503 82 507 86
rect 543 82 547 86
rect 583 82 587 86
rect 623 82 627 86
rect 663 82 667 86
rect 703 82 707 86
rect 743 82 747 86
rect 783 82 787 86
rect 831 82 835 86
rect 879 82 883 86
rect 927 82 931 86
rect 967 82 971 86
rect 1007 82 1011 86
rect 1047 82 1051 86
rect 1095 82 1099 86
rect 1135 82 1139 86
rect 1159 82 1163 86
rect 1207 82 1211 86
rect 1271 82 1275 86
rect 1335 82 1339 86
rect 1399 82 1403 86
rect 1455 82 1459 86
rect 1511 82 1515 86
rect 1559 82 1563 86
rect 1607 82 1611 86
rect 1647 82 1651 86
rect 1687 82 1691 86
rect 1727 82 1731 86
rect 1767 82 1771 86
rect 1807 82 1811 86
rect 1855 82 1859 86
rect 1903 82 1907 86
rect 1951 82 1955 86
rect 1991 82 1995 86
rect 2031 82 2035 86
rect 2071 82 2075 86
rect 2119 82 2123 86
<< m4 >>
rect 1118 2225 1119 2231
rect 1125 2230 2155 2231
rect 1125 2226 1135 2230
rect 1139 2226 1687 2230
rect 1691 2226 1727 2230
rect 1731 2226 1767 2230
rect 1771 2226 1807 2230
rect 1811 2226 2119 2230
rect 2123 2226 2155 2230
rect 1125 2225 2155 2226
rect 2161 2225 2162 2231
rect 84 2209 85 2215
rect 91 2214 1107 2215
rect 91 2210 111 2214
rect 115 2210 135 2214
rect 139 2210 175 2214
rect 179 2210 215 2214
rect 219 2210 255 2214
rect 259 2210 319 2214
rect 323 2210 383 2214
rect 387 2210 447 2214
rect 451 2210 511 2214
rect 515 2210 575 2214
rect 579 2210 631 2214
rect 635 2210 687 2214
rect 691 2210 735 2214
rect 739 2210 791 2214
rect 795 2210 847 2214
rect 851 2210 903 2214
rect 907 2210 1095 2214
rect 1099 2210 1107 2214
rect 91 2209 1107 2210
rect 1113 2209 1114 2215
rect 1106 2173 1107 2179
rect 1113 2178 2143 2179
rect 1113 2174 1135 2178
rect 1139 2174 1159 2178
rect 1163 2174 1199 2178
rect 1203 2174 1239 2178
rect 1243 2174 1279 2178
rect 1283 2174 1335 2178
rect 1339 2174 1391 2178
rect 1395 2174 1455 2178
rect 1459 2174 1527 2178
rect 1531 2174 1591 2178
rect 1595 2174 1663 2178
rect 1667 2174 1687 2178
rect 1691 2174 1727 2178
rect 1731 2174 1735 2178
rect 1739 2174 1767 2178
rect 1771 2174 1807 2178
rect 1811 2174 1879 2178
rect 1883 2174 2119 2178
rect 2123 2174 2143 2178
rect 1113 2173 2143 2174
rect 2149 2173 2150 2179
rect 96 2149 97 2155
rect 103 2154 1119 2155
rect 103 2150 111 2154
rect 115 2150 135 2154
rect 139 2150 175 2154
rect 179 2150 215 2154
rect 219 2150 231 2154
rect 235 2150 255 2154
rect 259 2150 271 2154
rect 275 2150 311 2154
rect 315 2150 319 2154
rect 323 2150 359 2154
rect 363 2150 383 2154
rect 387 2150 423 2154
rect 427 2150 447 2154
rect 451 2150 487 2154
rect 491 2150 511 2154
rect 515 2150 559 2154
rect 563 2150 575 2154
rect 579 2150 631 2154
rect 635 2150 639 2154
rect 643 2150 687 2154
rect 691 2150 719 2154
rect 723 2150 735 2154
rect 739 2150 791 2154
rect 795 2150 799 2154
rect 803 2150 847 2154
rect 851 2150 879 2154
rect 883 2150 903 2154
rect 907 2150 967 2154
rect 971 2150 1095 2154
rect 1099 2150 1119 2154
rect 103 2149 1119 2150
rect 1125 2149 1126 2155
rect 1118 2121 1119 2127
rect 1125 2126 2155 2127
rect 1125 2122 1135 2126
rect 1139 2122 1159 2126
rect 1163 2122 1199 2126
rect 1203 2122 1239 2126
rect 1243 2122 1279 2126
rect 1283 2122 1295 2126
rect 1299 2122 1335 2126
rect 1339 2122 1367 2126
rect 1371 2122 1391 2126
rect 1395 2122 1439 2126
rect 1443 2122 1455 2126
rect 1459 2122 1519 2126
rect 1523 2122 1527 2126
rect 1531 2122 1591 2126
rect 1595 2122 1599 2126
rect 1603 2122 1663 2126
rect 1667 2122 1679 2126
rect 1683 2122 1735 2126
rect 1739 2122 1751 2126
rect 1755 2122 1807 2126
rect 1811 2122 1823 2126
rect 1827 2122 1879 2126
rect 1883 2122 1887 2126
rect 1891 2122 1951 2126
rect 1955 2122 2023 2126
rect 2027 2122 2071 2126
rect 2075 2122 2119 2126
rect 2123 2122 2155 2126
rect 1125 2121 2155 2122
rect 2161 2121 2162 2127
rect 84 2093 85 2099
rect 91 2098 1107 2099
rect 91 2094 111 2098
rect 115 2094 231 2098
rect 235 2094 271 2098
rect 275 2094 303 2098
rect 307 2094 311 2098
rect 315 2094 351 2098
rect 355 2094 359 2098
rect 363 2094 407 2098
rect 411 2094 423 2098
rect 427 2094 471 2098
rect 475 2094 487 2098
rect 491 2094 543 2098
rect 547 2094 559 2098
rect 563 2094 623 2098
rect 627 2094 639 2098
rect 643 2094 703 2098
rect 707 2094 719 2098
rect 723 2094 783 2098
rect 787 2094 799 2098
rect 803 2094 863 2098
rect 867 2094 879 2098
rect 883 2094 951 2098
rect 955 2094 967 2098
rect 971 2094 1039 2098
rect 1043 2094 1095 2098
rect 1099 2094 1107 2098
rect 91 2093 1107 2094
rect 1113 2093 1114 2099
rect 1106 2069 1107 2075
rect 1113 2074 2143 2075
rect 1113 2070 1135 2074
rect 1139 2070 1159 2074
rect 1163 2070 1199 2074
rect 1203 2070 1215 2074
rect 1219 2070 1239 2074
rect 1243 2070 1295 2074
rect 1299 2070 1303 2074
rect 1307 2070 1367 2074
rect 1371 2070 1399 2074
rect 1403 2070 1439 2074
rect 1443 2070 1495 2074
rect 1499 2070 1519 2074
rect 1523 2070 1591 2074
rect 1595 2070 1599 2074
rect 1603 2070 1679 2074
rect 1683 2070 1751 2074
rect 1755 2070 1759 2074
rect 1763 2070 1823 2074
rect 1827 2070 1831 2074
rect 1835 2070 1887 2074
rect 1891 2070 1895 2074
rect 1899 2070 1951 2074
rect 1955 2070 1959 2074
rect 1963 2070 2023 2074
rect 2027 2070 2071 2074
rect 2075 2070 2119 2074
rect 2123 2070 2143 2074
rect 1113 2069 2143 2070
rect 2149 2069 2150 2075
rect 96 2037 97 2043
rect 103 2042 1119 2043
rect 103 2038 111 2042
rect 115 2038 183 2042
rect 187 2038 279 2042
rect 283 2038 303 2042
rect 307 2038 351 2042
rect 355 2038 375 2042
rect 379 2038 407 2042
rect 411 2038 463 2042
rect 467 2038 471 2042
rect 475 2038 543 2042
rect 547 2038 623 2042
rect 627 2038 695 2042
rect 699 2038 703 2042
rect 707 2038 759 2042
rect 763 2038 783 2042
rect 787 2038 815 2042
rect 819 2038 863 2042
rect 867 2038 911 2042
rect 915 2038 951 2042
rect 955 2038 959 2042
rect 963 2038 1007 2042
rect 1011 2038 1039 2042
rect 1043 2038 1047 2042
rect 1051 2038 1095 2042
rect 1099 2038 1119 2042
rect 103 2037 1119 2038
rect 1125 2037 1126 2043
rect 1118 2017 1119 2023
rect 1125 2022 2155 2023
rect 1125 2018 1135 2022
rect 1139 2018 1159 2022
rect 1163 2018 1215 2022
rect 1219 2018 1239 2022
rect 1243 2018 1303 2022
rect 1307 2018 1351 2022
rect 1355 2018 1399 2022
rect 1403 2018 1455 2022
rect 1459 2018 1495 2022
rect 1499 2018 1559 2022
rect 1563 2018 1591 2022
rect 1595 2018 1655 2022
rect 1659 2018 1679 2022
rect 1683 2018 1743 2022
rect 1747 2018 1759 2022
rect 1763 2018 1823 2022
rect 1827 2018 1831 2022
rect 1835 2018 1895 2022
rect 1899 2018 1959 2022
rect 1963 2018 2023 2022
rect 2027 2018 2071 2022
rect 2075 2018 2119 2022
rect 2123 2018 2155 2022
rect 1125 2017 2155 2018
rect 2161 2017 2162 2023
rect 84 1985 85 1991
rect 91 1990 1107 1991
rect 91 1986 111 1990
rect 115 1986 159 1990
rect 163 1986 183 1990
rect 187 1986 231 1990
rect 235 1986 279 1990
rect 283 1986 303 1990
rect 307 1986 375 1990
rect 379 1986 447 1990
rect 451 1986 463 1990
rect 467 1986 527 1990
rect 531 1986 543 1990
rect 547 1986 607 1990
rect 611 1986 623 1990
rect 627 1986 687 1990
rect 691 1986 695 1990
rect 699 1986 759 1990
rect 763 1986 815 1990
rect 819 1986 831 1990
rect 835 1986 863 1990
rect 867 1986 911 1990
rect 915 1986 959 1990
rect 963 1986 991 1990
rect 995 1986 1007 1990
rect 1011 1986 1047 1990
rect 1051 1986 1095 1990
rect 1099 1986 1107 1990
rect 91 1985 1107 1986
rect 1113 1985 1114 1991
rect 1106 1953 1107 1959
rect 1113 1958 2143 1959
rect 1113 1954 1135 1958
rect 1139 1954 1159 1958
rect 1163 1954 1239 1958
rect 1243 1954 1351 1958
rect 1355 1954 1359 1958
rect 1363 1954 1423 1958
rect 1427 1954 1455 1958
rect 1459 1954 1487 1958
rect 1491 1954 1559 1958
rect 1563 1954 1631 1958
rect 1635 1954 1655 1958
rect 1659 1954 1703 1958
rect 1707 1954 1743 1958
rect 1747 1954 1775 1958
rect 1779 1954 1823 1958
rect 1827 1954 1847 1958
rect 1851 1954 1895 1958
rect 1899 1954 1927 1958
rect 1931 1954 1959 1958
rect 1963 1954 2007 1958
rect 2011 1954 2023 1958
rect 2027 1954 2071 1958
rect 2075 1954 2119 1958
rect 2123 1954 2143 1958
rect 1113 1953 2143 1954
rect 2149 1953 2150 1959
rect 96 1929 97 1935
rect 103 1934 1119 1935
rect 103 1930 111 1934
rect 115 1930 135 1934
rect 139 1930 159 1934
rect 163 1930 175 1934
rect 179 1930 231 1934
rect 235 1930 295 1934
rect 299 1930 303 1934
rect 307 1930 367 1934
rect 371 1930 375 1934
rect 379 1930 447 1934
rect 451 1930 527 1934
rect 531 1930 607 1934
rect 611 1930 615 1934
rect 619 1930 687 1934
rect 691 1930 703 1934
rect 707 1930 759 1934
rect 763 1930 791 1934
rect 795 1930 831 1934
rect 835 1930 879 1934
rect 883 1930 911 1934
rect 915 1930 991 1934
rect 995 1930 1095 1934
rect 1099 1930 1119 1934
rect 103 1929 1119 1930
rect 1125 1929 1126 1935
rect 1118 1901 1119 1907
rect 1125 1906 2155 1907
rect 1125 1902 1135 1906
rect 1139 1902 1231 1906
rect 1235 1902 1271 1906
rect 1275 1902 1319 1906
rect 1323 1902 1359 1906
rect 1363 1902 1375 1906
rect 1379 1902 1423 1906
rect 1427 1902 1439 1906
rect 1443 1902 1487 1906
rect 1491 1902 1503 1906
rect 1507 1902 1559 1906
rect 1563 1902 1575 1906
rect 1579 1902 1631 1906
rect 1635 1902 1655 1906
rect 1659 1902 1703 1906
rect 1707 1902 1751 1906
rect 1755 1902 1775 1906
rect 1779 1902 1847 1906
rect 1851 1902 1863 1906
rect 1867 1902 1927 1906
rect 1931 1902 1975 1906
rect 1979 1902 2007 1906
rect 2011 1902 2071 1906
rect 2075 1902 2119 1906
rect 2123 1902 2155 1906
rect 1125 1901 2155 1902
rect 2161 1901 2162 1907
rect 84 1873 85 1879
rect 91 1878 1107 1879
rect 91 1874 111 1878
rect 115 1874 135 1878
rect 139 1874 175 1878
rect 179 1874 223 1878
rect 227 1874 231 1878
rect 235 1874 287 1878
rect 291 1874 295 1878
rect 299 1874 359 1878
rect 363 1874 367 1878
rect 371 1874 431 1878
rect 435 1874 447 1878
rect 451 1874 503 1878
rect 507 1874 527 1878
rect 531 1874 567 1878
rect 571 1874 615 1878
rect 619 1874 631 1878
rect 635 1874 695 1878
rect 699 1874 703 1878
rect 707 1874 759 1878
rect 763 1874 791 1878
rect 795 1874 831 1878
rect 835 1874 879 1878
rect 883 1874 1095 1878
rect 1099 1874 1107 1878
rect 91 1873 1107 1874
rect 1113 1873 1114 1879
rect 1106 1845 1107 1851
rect 1113 1850 2143 1851
rect 1113 1846 1135 1850
rect 1139 1846 1159 1850
rect 1163 1846 1199 1850
rect 1203 1846 1231 1850
rect 1235 1846 1239 1850
rect 1243 1846 1271 1850
rect 1275 1846 1303 1850
rect 1307 1846 1319 1850
rect 1323 1846 1367 1850
rect 1371 1846 1375 1850
rect 1379 1846 1431 1850
rect 1435 1846 1439 1850
rect 1443 1846 1503 1850
rect 1507 1846 1575 1850
rect 1579 1846 1583 1850
rect 1587 1846 1655 1850
rect 1659 1846 1671 1850
rect 1675 1846 1751 1850
rect 1755 1846 1767 1850
rect 1771 1846 1863 1850
rect 1867 1846 1871 1850
rect 1875 1846 1975 1850
rect 1979 1846 1983 1850
rect 1987 1846 2071 1850
rect 2075 1846 2119 1850
rect 2123 1846 2143 1850
rect 1113 1845 2143 1846
rect 2149 1845 2150 1851
rect 96 1817 97 1823
rect 103 1822 1119 1823
rect 103 1818 111 1822
rect 115 1818 135 1822
rect 139 1818 175 1822
rect 179 1818 183 1822
rect 187 1818 223 1822
rect 227 1818 263 1822
rect 267 1818 287 1822
rect 291 1818 351 1822
rect 355 1818 359 1822
rect 363 1818 431 1822
rect 435 1818 439 1822
rect 443 1818 503 1822
rect 507 1818 527 1822
rect 531 1818 567 1822
rect 571 1818 607 1822
rect 611 1818 631 1822
rect 635 1818 687 1822
rect 691 1818 695 1822
rect 699 1818 759 1822
rect 763 1818 767 1822
rect 771 1818 831 1822
rect 835 1818 839 1822
rect 843 1818 911 1822
rect 915 1818 991 1822
rect 995 1818 1047 1822
rect 1051 1818 1095 1822
rect 1099 1818 1119 1822
rect 103 1817 1119 1818
rect 1125 1817 1126 1823
rect 1118 1785 1119 1791
rect 1125 1790 2155 1791
rect 1125 1786 1135 1790
rect 1139 1786 1159 1790
rect 1163 1786 1199 1790
rect 1203 1786 1239 1790
rect 1243 1786 1303 1790
rect 1307 1786 1311 1790
rect 1315 1786 1351 1790
rect 1355 1786 1367 1790
rect 1371 1786 1391 1790
rect 1395 1786 1431 1790
rect 1435 1786 1471 1790
rect 1475 1786 1503 1790
rect 1507 1786 1511 1790
rect 1515 1786 1551 1790
rect 1555 1786 1583 1790
rect 1587 1786 1607 1790
rect 1611 1786 1671 1790
rect 1675 1786 1679 1790
rect 1683 1786 1767 1790
rect 1771 1786 1871 1790
rect 1875 1786 1983 1790
rect 1987 1786 2071 1790
rect 2075 1786 2119 1790
rect 2123 1786 2155 1790
rect 1125 1785 2155 1786
rect 2161 1785 2162 1791
rect 84 1757 85 1763
rect 91 1762 1107 1763
rect 91 1758 111 1762
rect 115 1758 135 1762
rect 139 1758 183 1762
rect 187 1758 199 1762
rect 203 1758 263 1762
rect 267 1758 295 1762
rect 299 1758 351 1762
rect 355 1758 399 1762
rect 403 1758 439 1762
rect 443 1758 495 1762
rect 499 1758 527 1762
rect 531 1758 591 1762
rect 595 1758 607 1762
rect 611 1758 671 1762
rect 675 1758 687 1762
rect 691 1758 751 1762
rect 755 1758 767 1762
rect 771 1758 823 1762
rect 827 1758 839 1762
rect 843 1758 887 1762
rect 891 1758 911 1762
rect 915 1758 959 1762
rect 963 1758 991 1762
rect 995 1758 1031 1762
rect 1035 1758 1047 1762
rect 1051 1758 1095 1762
rect 1099 1758 1107 1762
rect 91 1757 1107 1758
rect 1113 1757 1114 1763
rect 1106 1729 1107 1735
rect 1113 1734 2143 1735
rect 1113 1730 1135 1734
rect 1139 1730 1263 1734
rect 1267 1730 1311 1734
rect 1315 1730 1319 1734
rect 1323 1730 1351 1734
rect 1355 1730 1383 1734
rect 1387 1730 1391 1734
rect 1395 1730 1431 1734
rect 1435 1730 1455 1734
rect 1459 1730 1471 1734
rect 1475 1730 1511 1734
rect 1515 1730 1535 1734
rect 1539 1730 1551 1734
rect 1555 1730 1607 1734
rect 1611 1730 1615 1734
rect 1619 1730 1679 1734
rect 1683 1730 1687 1734
rect 1691 1730 1759 1734
rect 1763 1730 1767 1734
rect 1771 1730 1831 1734
rect 1835 1730 1871 1734
rect 1875 1730 1895 1734
rect 1899 1730 1959 1734
rect 1963 1730 1983 1734
rect 1987 1730 2023 1734
rect 2027 1730 2071 1734
rect 2075 1730 2119 1734
rect 2123 1730 2143 1734
rect 1113 1729 2143 1730
rect 2149 1729 2150 1735
rect 96 1701 97 1707
rect 103 1706 1119 1707
rect 103 1702 111 1706
rect 115 1702 135 1706
rect 139 1702 151 1706
rect 155 1702 199 1706
rect 203 1702 223 1706
rect 227 1702 295 1706
rect 299 1702 303 1706
rect 307 1702 383 1706
rect 387 1702 399 1706
rect 403 1702 463 1706
rect 467 1702 495 1706
rect 499 1702 535 1706
rect 539 1702 591 1706
rect 595 1702 607 1706
rect 611 1702 671 1706
rect 675 1702 735 1706
rect 739 1702 751 1706
rect 755 1702 807 1706
rect 811 1702 823 1706
rect 827 1702 879 1706
rect 883 1702 887 1706
rect 891 1702 959 1706
rect 963 1702 1031 1706
rect 1035 1702 1095 1706
rect 1099 1702 1119 1706
rect 103 1701 1119 1702
rect 1125 1701 1126 1707
rect 1118 1677 1119 1683
rect 1125 1682 2155 1683
rect 1125 1678 1135 1682
rect 1139 1678 1167 1682
rect 1171 1678 1247 1682
rect 1251 1678 1263 1682
rect 1267 1678 1319 1682
rect 1323 1678 1335 1682
rect 1339 1678 1383 1682
rect 1387 1678 1423 1682
rect 1427 1678 1455 1682
rect 1459 1678 1511 1682
rect 1515 1678 1535 1682
rect 1539 1678 1599 1682
rect 1603 1678 1615 1682
rect 1619 1678 1679 1682
rect 1683 1678 1687 1682
rect 1691 1678 1751 1682
rect 1755 1678 1759 1682
rect 1763 1678 1815 1682
rect 1819 1678 1831 1682
rect 1835 1678 1871 1682
rect 1875 1678 1895 1682
rect 1899 1678 1927 1682
rect 1931 1678 1959 1682
rect 1963 1678 1983 1682
rect 1987 1678 2023 1682
rect 2027 1678 2031 1682
rect 2035 1678 2071 1682
rect 2075 1678 2119 1682
rect 2123 1678 2155 1682
rect 1125 1677 2155 1678
rect 2161 1677 2162 1683
rect 84 1645 85 1651
rect 91 1650 1107 1651
rect 91 1646 111 1650
rect 115 1646 151 1650
rect 155 1646 175 1650
rect 179 1646 215 1650
rect 219 1646 223 1650
rect 227 1646 255 1650
rect 259 1646 303 1650
rect 307 1646 359 1650
rect 363 1646 383 1650
rect 387 1646 407 1650
rect 411 1646 455 1650
rect 459 1646 463 1650
rect 467 1646 503 1650
rect 507 1646 535 1650
rect 539 1646 551 1650
rect 555 1646 607 1650
rect 611 1646 663 1650
rect 667 1646 671 1650
rect 675 1646 719 1650
rect 723 1646 735 1650
rect 739 1646 807 1650
rect 811 1646 879 1650
rect 883 1646 1095 1650
rect 1099 1646 1107 1650
rect 91 1645 1107 1646
rect 1113 1645 1114 1651
rect 1106 1621 1107 1627
rect 1113 1626 2143 1627
rect 1113 1622 1135 1626
rect 1139 1622 1159 1626
rect 1163 1622 1167 1626
rect 1171 1622 1199 1626
rect 1203 1622 1247 1626
rect 1251 1622 1319 1626
rect 1323 1622 1335 1626
rect 1339 1622 1391 1626
rect 1395 1622 1423 1626
rect 1427 1622 1463 1626
rect 1467 1622 1511 1626
rect 1515 1622 1535 1626
rect 1539 1622 1599 1626
rect 1603 1622 1607 1626
rect 1611 1622 1679 1626
rect 1683 1622 1751 1626
rect 1755 1622 1815 1626
rect 1819 1622 1831 1626
rect 1835 1622 1871 1626
rect 1875 1622 1927 1626
rect 1931 1622 1983 1626
rect 1987 1622 2031 1626
rect 2035 1622 2071 1626
rect 2075 1622 2119 1626
rect 2123 1622 2143 1626
rect 1113 1621 2143 1622
rect 2149 1621 2150 1627
rect 96 1585 97 1591
rect 103 1590 1119 1591
rect 103 1586 111 1590
rect 115 1586 143 1590
rect 147 1586 175 1590
rect 179 1586 183 1590
rect 187 1586 215 1590
rect 219 1586 231 1590
rect 235 1586 255 1590
rect 259 1586 287 1590
rect 291 1586 303 1590
rect 307 1586 351 1590
rect 355 1586 359 1590
rect 363 1586 407 1590
rect 411 1586 415 1590
rect 419 1586 455 1590
rect 459 1586 479 1590
rect 483 1586 503 1590
rect 507 1586 543 1590
rect 547 1586 551 1590
rect 555 1586 607 1590
rect 611 1586 663 1590
rect 667 1586 719 1590
rect 723 1586 727 1590
rect 731 1586 791 1590
rect 795 1586 855 1590
rect 859 1586 1095 1590
rect 1099 1586 1119 1590
rect 103 1585 1119 1586
rect 1125 1585 1126 1591
rect 1118 1569 1119 1575
rect 1125 1574 2155 1575
rect 1125 1570 1135 1574
rect 1139 1570 1159 1574
rect 1163 1570 1199 1574
rect 1203 1570 1239 1574
rect 1243 1570 1247 1574
rect 1251 1570 1279 1574
rect 1283 1570 1319 1574
rect 1323 1570 1327 1574
rect 1331 1570 1375 1574
rect 1379 1570 1391 1574
rect 1395 1570 1423 1574
rect 1427 1570 1463 1574
rect 1467 1570 1471 1574
rect 1475 1570 1519 1574
rect 1523 1570 1535 1574
rect 1539 1570 1567 1574
rect 1571 1570 1607 1574
rect 1611 1570 1623 1574
rect 1627 1570 1679 1574
rect 1683 1570 1735 1574
rect 1739 1570 1751 1574
rect 1755 1570 1831 1574
rect 1835 1570 2119 1574
rect 2123 1570 2155 1574
rect 1125 1569 2155 1570
rect 2161 1569 2162 1575
rect 84 1525 85 1531
rect 91 1530 1107 1531
rect 91 1526 111 1530
rect 115 1526 135 1530
rect 139 1526 143 1530
rect 147 1526 175 1530
rect 179 1526 183 1530
rect 187 1526 215 1530
rect 219 1526 231 1530
rect 235 1526 255 1530
rect 259 1526 287 1530
rect 291 1526 295 1530
rect 299 1526 335 1530
rect 339 1526 351 1530
rect 355 1526 375 1530
rect 379 1526 415 1530
rect 419 1526 455 1530
rect 459 1526 479 1530
rect 483 1526 495 1530
rect 499 1526 535 1530
rect 539 1526 543 1530
rect 547 1526 575 1530
rect 579 1526 607 1530
rect 611 1526 615 1530
rect 619 1526 655 1530
rect 659 1526 663 1530
rect 667 1526 695 1530
rect 699 1526 727 1530
rect 731 1526 735 1530
rect 739 1526 775 1530
rect 779 1526 791 1530
rect 795 1526 831 1530
rect 835 1526 855 1530
rect 859 1526 887 1530
rect 891 1526 1095 1530
rect 1099 1526 1107 1530
rect 91 1525 1107 1526
rect 1113 1525 1114 1531
rect 1106 1513 1107 1519
rect 1113 1518 2143 1519
rect 1113 1514 1135 1518
rect 1139 1514 1239 1518
rect 1243 1514 1279 1518
rect 1283 1514 1319 1518
rect 1323 1514 1327 1518
rect 1331 1514 1359 1518
rect 1363 1514 1375 1518
rect 1379 1514 1399 1518
rect 1403 1514 1423 1518
rect 1427 1514 1439 1518
rect 1443 1514 1471 1518
rect 1475 1514 1479 1518
rect 1483 1514 1519 1518
rect 1523 1514 1559 1518
rect 1563 1514 1567 1518
rect 1571 1514 1607 1518
rect 1611 1514 1623 1518
rect 1627 1514 1663 1518
rect 1667 1514 1679 1518
rect 1683 1514 1735 1518
rect 1739 1514 1815 1518
rect 1819 1514 1903 1518
rect 1907 1514 1991 1518
rect 1995 1514 2071 1518
rect 2075 1514 2119 1518
rect 2123 1514 2143 1518
rect 1113 1513 2143 1514
rect 2149 1513 2150 1519
rect 96 1465 97 1471
rect 103 1470 1119 1471
rect 103 1466 111 1470
rect 115 1466 135 1470
rect 139 1466 175 1470
rect 179 1466 215 1470
rect 219 1466 255 1470
rect 259 1466 295 1470
rect 299 1466 335 1470
rect 339 1466 375 1470
rect 379 1466 415 1470
rect 419 1466 455 1470
rect 459 1466 495 1470
rect 499 1466 519 1470
rect 523 1466 535 1470
rect 539 1466 559 1470
rect 563 1466 575 1470
rect 579 1466 599 1470
rect 603 1466 615 1470
rect 619 1466 647 1470
rect 651 1466 655 1470
rect 659 1466 695 1470
rect 699 1466 735 1470
rect 739 1466 751 1470
rect 755 1466 775 1470
rect 779 1466 807 1470
rect 811 1466 831 1470
rect 835 1466 871 1470
rect 875 1466 887 1470
rect 891 1466 935 1470
rect 939 1466 1095 1470
rect 1099 1466 1119 1470
rect 103 1465 1119 1466
rect 1125 1467 1126 1471
rect 1125 1466 2162 1467
rect 1125 1465 1135 1466
rect 1118 1462 1135 1465
rect 1139 1462 1231 1466
rect 1235 1462 1279 1466
rect 1283 1462 1319 1466
rect 1323 1462 1335 1466
rect 1339 1462 1359 1466
rect 1363 1462 1391 1466
rect 1395 1462 1399 1466
rect 1403 1462 1439 1466
rect 1443 1462 1455 1466
rect 1459 1462 1479 1466
rect 1483 1462 1519 1466
rect 1523 1462 1559 1466
rect 1563 1462 1583 1466
rect 1587 1462 1607 1466
rect 1611 1462 1647 1466
rect 1651 1462 1663 1466
rect 1667 1462 1719 1466
rect 1723 1462 1735 1466
rect 1739 1462 1807 1466
rect 1811 1462 1815 1466
rect 1819 1462 1895 1466
rect 1899 1462 1903 1466
rect 1907 1462 1991 1466
rect 1995 1462 2071 1466
rect 2075 1462 2119 1466
rect 2123 1462 2162 1466
rect 1118 1461 2162 1462
rect 84 1409 85 1415
rect 91 1414 1107 1415
rect 91 1410 111 1414
rect 115 1410 431 1414
rect 435 1410 471 1414
rect 475 1410 519 1414
rect 523 1410 559 1414
rect 563 1410 575 1414
rect 579 1410 599 1414
rect 603 1410 631 1414
rect 635 1410 647 1414
rect 651 1410 695 1414
rect 699 1410 751 1414
rect 755 1410 759 1414
rect 763 1410 807 1414
rect 811 1410 823 1414
rect 827 1410 871 1414
rect 875 1410 895 1414
rect 899 1410 935 1414
rect 939 1410 967 1414
rect 971 1410 1095 1414
rect 1099 1410 1107 1414
rect 91 1409 1107 1410
rect 1113 1411 1114 1415
rect 1113 1410 2150 1411
rect 1113 1409 1135 1410
rect 1106 1406 1135 1409
rect 1139 1406 1159 1410
rect 1163 1406 1199 1410
rect 1203 1406 1231 1410
rect 1235 1406 1263 1410
rect 1267 1406 1279 1410
rect 1283 1406 1335 1410
rect 1339 1406 1351 1410
rect 1355 1406 1391 1410
rect 1395 1406 1447 1410
rect 1451 1406 1455 1410
rect 1459 1406 1519 1410
rect 1523 1406 1543 1410
rect 1547 1406 1583 1410
rect 1587 1406 1631 1410
rect 1635 1406 1647 1410
rect 1651 1406 1719 1410
rect 1723 1406 1799 1410
rect 1803 1406 1807 1410
rect 1811 1406 1871 1410
rect 1875 1406 1895 1410
rect 1899 1406 1943 1410
rect 1947 1406 1991 1410
rect 1995 1406 2015 1410
rect 2019 1406 2071 1410
rect 2075 1406 2119 1410
rect 2123 1406 2150 1410
rect 1106 1405 2150 1406
rect 96 1357 97 1363
rect 103 1362 1119 1363
rect 103 1358 111 1362
rect 115 1358 375 1362
rect 379 1358 423 1362
rect 427 1358 431 1362
rect 435 1358 471 1362
rect 475 1358 479 1362
rect 483 1358 519 1362
rect 523 1358 543 1362
rect 547 1358 575 1362
rect 579 1358 607 1362
rect 611 1358 631 1362
rect 635 1358 671 1362
rect 675 1358 695 1362
rect 699 1358 735 1362
rect 739 1358 759 1362
rect 763 1358 799 1362
rect 803 1358 823 1362
rect 827 1358 863 1362
rect 867 1358 895 1362
rect 899 1358 927 1362
rect 931 1358 967 1362
rect 971 1358 999 1362
rect 1003 1358 1047 1362
rect 1051 1358 1095 1362
rect 1099 1358 1119 1362
rect 103 1357 1119 1358
rect 1125 1357 1126 1363
rect 1118 1355 1126 1357
rect 1118 1349 1119 1355
rect 1125 1354 2155 1355
rect 1125 1350 1135 1354
rect 1139 1350 1159 1354
rect 1163 1350 1199 1354
rect 1203 1350 1255 1354
rect 1259 1350 1263 1354
rect 1267 1350 1351 1354
rect 1355 1350 1375 1354
rect 1379 1350 1447 1354
rect 1451 1350 1487 1354
rect 1491 1350 1543 1354
rect 1547 1350 1591 1354
rect 1595 1350 1631 1354
rect 1635 1350 1679 1354
rect 1683 1350 1719 1354
rect 1723 1350 1759 1354
rect 1763 1350 1799 1354
rect 1803 1350 1831 1354
rect 1835 1350 1871 1354
rect 1875 1350 1903 1354
rect 1907 1350 1943 1354
rect 1947 1350 1967 1354
rect 1971 1350 2015 1354
rect 2019 1350 2031 1354
rect 2035 1350 2071 1354
rect 2075 1350 2119 1354
rect 2123 1350 2155 1354
rect 1125 1349 2155 1350
rect 2161 1349 2162 1355
rect 84 1305 85 1311
rect 91 1310 1107 1311
rect 91 1306 111 1310
rect 115 1306 335 1310
rect 339 1306 375 1310
rect 379 1306 391 1310
rect 395 1306 423 1310
rect 427 1306 455 1310
rect 459 1306 479 1310
rect 483 1306 527 1310
rect 531 1306 543 1310
rect 547 1306 599 1310
rect 603 1306 607 1310
rect 611 1306 671 1310
rect 675 1306 735 1310
rect 739 1306 743 1310
rect 747 1306 799 1310
rect 803 1306 823 1310
rect 827 1306 863 1310
rect 867 1306 903 1310
rect 907 1306 927 1310
rect 931 1306 983 1310
rect 987 1306 999 1310
rect 1003 1306 1047 1310
rect 1051 1306 1095 1310
rect 1099 1306 1107 1310
rect 91 1305 1107 1306
rect 1113 1305 1114 1311
rect 1106 1293 1107 1299
rect 1113 1298 2143 1299
rect 1113 1294 1135 1298
rect 1139 1294 1159 1298
rect 1163 1294 1199 1298
rect 1203 1294 1247 1298
rect 1251 1294 1255 1298
rect 1259 1294 1319 1298
rect 1323 1294 1375 1298
rect 1379 1294 1399 1298
rect 1403 1294 1479 1298
rect 1483 1294 1487 1298
rect 1491 1294 1559 1298
rect 1563 1294 1591 1298
rect 1595 1294 1639 1298
rect 1643 1294 1679 1298
rect 1683 1294 1719 1298
rect 1723 1294 1759 1298
rect 1763 1294 1799 1298
rect 1803 1294 1831 1298
rect 1835 1294 1879 1298
rect 1883 1294 1903 1298
rect 1907 1294 1967 1298
rect 1971 1294 2031 1298
rect 2035 1294 2055 1298
rect 2059 1294 2071 1298
rect 2075 1294 2119 1298
rect 2123 1294 2143 1298
rect 1113 1293 2143 1294
rect 2149 1293 2150 1299
rect 96 1249 97 1255
rect 103 1254 1119 1255
rect 103 1250 111 1254
rect 115 1250 263 1254
rect 267 1250 311 1254
rect 315 1250 335 1254
rect 339 1250 359 1254
rect 363 1250 391 1254
rect 395 1250 415 1254
rect 419 1250 455 1254
rect 459 1250 479 1254
rect 483 1250 527 1254
rect 531 1250 543 1254
rect 547 1250 599 1254
rect 603 1250 607 1254
rect 611 1250 671 1254
rect 675 1250 735 1254
rect 739 1250 743 1254
rect 747 1250 799 1254
rect 803 1250 823 1254
rect 827 1250 863 1254
rect 867 1250 903 1254
rect 907 1250 927 1254
rect 931 1250 983 1254
rect 987 1250 1047 1254
rect 1051 1250 1095 1254
rect 1099 1250 1119 1254
rect 103 1249 1119 1250
rect 1125 1249 1126 1255
rect 1118 1237 1119 1243
rect 1125 1242 2155 1243
rect 1125 1238 1135 1242
rect 1139 1238 1159 1242
rect 1163 1238 1199 1242
rect 1203 1238 1239 1242
rect 1243 1238 1247 1242
rect 1251 1238 1279 1242
rect 1283 1238 1319 1242
rect 1323 1238 1327 1242
rect 1331 1238 1375 1242
rect 1379 1238 1399 1242
rect 1403 1238 1423 1242
rect 1427 1238 1471 1242
rect 1475 1238 1479 1242
rect 1483 1238 1535 1242
rect 1539 1238 1559 1242
rect 1563 1238 1615 1242
rect 1619 1238 1639 1242
rect 1643 1238 1719 1242
rect 1723 1238 1799 1242
rect 1803 1238 1839 1242
rect 1843 1238 1879 1242
rect 1883 1238 1967 1242
rect 1971 1238 2055 1242
rect 2059 1238 2071 1242
rect 2075 1238 2119 1242
rect 2123 1238 2155 1242
rect 1125 1237 2155 1238
rect 2161 1237 2162 1243
rect 84 1197 85 1203
rect 91 1202 1107 1203
rect 91 1198 111 1202
rect 115 1198 223 1202
rect 227 1198 263 1202
rect 267 1198 279 1202
rect 283 1198 311 1202
rect 315 1198 343 1202
rect 347 1198 359 1202
rect 363 1198 407 1202
rect 411 1198 415 1202
rect 419 1198 479 1202
rect 483 1198 543 1202
rect 547 1198 551 1202
rect 555 1198 607 1202
rect 611 1198 631 1202
rect 635 1198 671 1202
rect 675 1198 711 1202
rect 715 1198 735 1202
rect 739 1198 791 1202
rect 795 1198 799 1202
rect 803 1198 863 1202
rect 867 1198 871 1202
rect 875 1198 927 1202
rect 931 1198 959 1202
rect 963 1198 1095 1202
rect 1099 1198 1107 1202
rect 91 1197 1107 1198
rect 1113 1197 1114 1203
rect 1106 1185 1107 1191
rect 1113 1190 2143 1191
rect 1113 1186 1135 1190
rect 1139 1186 1159 1190
rect 1163 1186 1199 1190
rect 1203 1186 1239 1190
rect 1243 1186 1279 1190
rect 1283 1186 1287 1190
rect 1291 1186 1327 1190
rect 1331 1186 1367 1190
rect 1371 1186 1375 1190
rect 1379 1186 1415 1190
rect 1419 1186 1423 1190
rect 1427 1186 1471 1190
rect 1475 1186 1527 1190
rect 1531 1186 1535 1190
rect 1539 1186 1583 1190
rect 1587 1186 1615 1190
rect 1619 1186 1639 1190
rect 1643 1186 1703 1190
rect 1707 1186 1719 1190
rect 1723 1186 1767 1190
rect 1771 1186 1839 1190
rect 1843 1186 1919 1190
rect 1923 1186 1967 1190
rect 1971 1186 2007 1190
rect 2011 1186 2071 1190
rect 2075 1186 2119 1190
rect 2123 1186 2143 1190
rect 1113 1185 2143 1186
rect 2149 1185 2150 1191
rect 96 1145 97 1151
rect 103 1150 1119 1151
rect 103 1146 111 1150
rect 115 1146 159 1150
rect 163 1146 199 1150
rect 203 1146 223 1150
rect 227 1146 247 1150
rect 251 1146 279 1150
rect 283 1146 303 1150
rect 307 1146 343 1150
rect 347 1146 367 1150
rect 371 1146 407 1150
rect 411 1146 439 1150
rect 443 1146 479 1150
rect 483 1146 511 1150
rect 515 1146 551 1150
rect 555 1146 591 1150
rect 595 1146 631 1150
rect 635 1146 679 1150
rect 683 1146 711 1150
rect 715 1146 775 1150
rect 779 1146 791 1150
rect 795 1146 871 1150
rect 875 1146 879 1150
rect 883 1146 959 1150
rect 963 1146 991 1150
rect 995 1146 1095 1150
rect 1099 1146 1119 1150
rect 103 1145 1119 1146
rect 1125 1145 1126 1151
rect 1118 1125 1119 1131
rect 1125 1130 2155 1131
rect 1125 1126 1135 1130
rect 1139 1126 1287 1130
rect 1291 1126 1327 1130
rect 1331 1126 1367 1130
rect 1371 1126 1383 1130
rect 1387 1126 1415 1130
rect 1419 1126 1423 1130
rect 1427 1126 1471 1130
rect 1475 1126 1527 1130
rect 1531 1126 1583 1130
rect 1587 1126 1591 1130
rect 1595 1126 1639 1130
rect 1643 1126 1655 1130
rect 1659 1126 1703 1130
rect 1707 1126 1711 1130
rect 1715 1126 1767 1130
rect 1771 1126 1823 1130
rect 1827 1126 1839 1130
rect 1843 1126 1871 1130
rect 1875 1126 1919 1130
rect 1923 1126 1927 1130
rect 1931 1126 1983 1130
rect 1987 1126 2007 1130
rect 2011 1126 2031 1130
rect 2035 1126 2071 1130
rect 2075 1126 2119 1130
rect 2123 1126 2155 1130
rect 1125 1125 2155 1126
rect 2161 1125 2162 1131
rect 84 1085 85 1091
rect 91 1090 1107 1091
rect 91 1086 111 1090
rect 115 1086 159 1090
rect 163 1086 199 1090
rect 203 1086 247 1090
rect 251 1086 303 1090
rect 307 1086 367 1090
rect 371 1086 431 1090
rect 435 1086 439 1090
rect 443 1086 503 1090
rect 507 1086 511 1090
rect 515 1086 575 1090
rect 579 1086 591 1090
rect 595 1086 647 1090
rect 651 1086 679 1090
rect 683 1086 719 1090
rect 723 1086 775 1090
rect 779 1086 783 1090
rect 787 1086 839 1090
rect 843 1086 879 1090
rect 883 1086 895 1090
rect 899 1086 951 1090
rect 955 1086 991 1090
rect 995 1086 1007 1090
rect 1011 1086 1047 1090
rect 1051 1086 1095 1090
rect 1099 1086 1107 1090
rect 91 1085 1107 1086
rect 1113 1085 1114 1091
rect 1106 1073 1107 1079
rect 1113 1078 2143 1079
rect 1113 1074 1135 1078
rect 1139 1074 1159 1078
rect 1163 1074 1247 1078
rect 1251 1074 1359 1078
rect 1363 1074 1383 1078
rect 1387 1074 1423 1078
rect 1427 1074 1471 1078
rect 1475 1074 1527 1078
rect 1531 1074 1575 1078
rect 1579 1074 1591 1078
rect 1595 1074 1655 1078
rect 1659 1074 1671 1078
rect 1675 1074 1711 1078
rect 1715 1074 1759 1078
rect 1763 1074 1767 1078
rect 1771 1074 1823 1078
rect 1827 1074 1847 1078
rect 1851 1074 1871 1078
rect 1875 1074 1927 1078
rect 1931 1074 1983 1078
rect 1987 1074 2007 1078
rect 2011 1074 2031 1078
rect 2035 1074 2071 1078
rect 2075 1074 2119 1078
rect 2123 1074 2143 1078
rect 1113 1073 2143 1074
rect 2149 1073 2150 1079
rect 96 1029 97 1035
rect 103 1034 1119 1035
rect 103 1030 111 1034
rect 115 1030 199 1034
rect 203 1030 223 1034
rect 227 1030 247 1034
rect 251 1030 271 1034
rect 275 1030 303 1034
rect 307 1030 335 1034
rect 339 1030 367 1034
rect 371 1030 407 1034
rect 411 1030 431 1034
rect 435 1030 479 1034
rect 483 1030 503 1034
rect 507 1030 559 1034
rect 563 1030 575 1034
rect 579 1030 631 1034
rect 635 1030 647 1034
rect 651 1030 703 1034
rect 707 1030 719 1034
rect 723 1030 775 1034
rect 779 1030 783 1034
rect 787 1030 839 1034
rect 843 1030 895 1034
rect 899 1030 903 1034
rect 907 1030 951 1034
rect 955 1030 967 1034
rect 971 1030 1007 1034
rect 1011 1030 1039 1034
rect 1043 1030 1047 1034
rect 1051 1030 1095 1034
rect 1099 1030 1119 1034
rect 103 1029 1119 1030
rect 1125 1029 1126 1035
rect 1118 1027 1126 1029
rect 1118 1021 1119 1027
rect 1125 1026 2155 1027
rect 1125 1022 1135 1026
rect 1139 1022 1159 1026
rect 1163 1022 1231 1026
rect 1235 1022 1247 1026
rect 1251 1022 1303 1026
rect 1307 1022 1359 1026
rect 1363 1022 1383 1026
rect 1387 1022 1463 1026
rect 1467 1022 1471 1026
rect 1475 1022 1543 1026
rect 1547 1022 1575 1026
rect 1579 1022 1623 1026
rect 1627 1022 1671 1026
rect 1675 1022 1695 1026
rect 1699 1022 1759 1026
rect 1763 1022 1823 1026
rect 1827 1022 1847 1026
rect 1851 1022 1887 1026
rect 1891 1022 1927 1026
rect 1931 1022 1951 1026
rect 1955 1022 2007 1026
rect 2011 1022 2071 1026
rect 2075 1022 2119 1026
rect 2123 1022 2155 1026
rect 1125 1021 2155 1022
rect 2161 1021 2162 1027
rect 84 973 85 979
rect 91 978 1107 979
rect 91 974 111 978
rect 115 974 151 978
rect 155 974 215 978
rect 219 974 223 978
rect 227 974 271 978
rect 275 974 287 978
rect 291 974 335 978
rect 339 974 367 978
rect 371 974 407 978
rect 411 974 447 978
rect 451 974 479 978
rect 483 974 527 978
rect 531 974 559 978
rect 563 974 599 978
rect 603 974 631 978
rect 635 974 671 978
rect 675 974 703 978
rect 707 974 735 978
rect 739 974 775 978
rect 779 974 799 978
rect 803 974 839 978
rect 843 974 863 978
rect 867 974 903 978
rect 907 974 927 978
rect 931 974 967 978
rect 971 974 991 978
rect 995 974 1039 978
rect 1043 974 1047 978
rect 1051 974 1095 978
rect 1099 974 1107 978
rect 91 973 1107 974
rect 1113 975 1114 979
rect 1113 974 2150 975
rect 1113 973 1135 974
rect 1106 970 1135 973
rect 1139 970 1159 974
rect 1163 970 1231 974
rect 1235 970 1239 974
rect 1243 970 1303 974
rect 1307 970 1375 974
rect 1379 970 1383 974
rect 1387 970 1439 974
rect 1443 970 1463 974
rect 1467 970 1511 974
rect 1515 970 1543 974
rect 1547 970 1583 974
rect 1587 970 1623 974
rect 1627 970 1655 974
rect 1659 970 1695 974
rect 1699 970 1727 974
rect 1731 970 1759 974
rect 1763 970 1799 974
rect 1803 970 1823 974
rect 1827 970 1871 974
rect 1875 970 1887 974
rect 1891 970 1943 974
rect 1947 970 1951 974
rect 1955 970 2015 974
rect 2019 970 2071 974
rect 2075 970 2119 974
rect 2123 970 2150 974
rect 1106 969 2150 970
rect 96 921 97 927
rect 103 926 1119 927
rect 103 922 111 926
rect 115 922 135 926
rect 139 922 151 926
rect 155 922 183 926
rect 187 922 215 926
rect 219 922 255 926
rect 259 922 287 926
rect 291 922 327 926
rect 331 922 367 926
rect 371 922 399 926
rect 403 922 447 926
rect 451 922 463 926
rect 467 922 527 926
rect 531 922 599 926
rect 603 922 671 926
rect 675 922 735 926
rect 739 922 743 926
rect 747 922 799 926
rect 803 922 815 926
rect 819 922 863 926
rect 867 922 895 926
rect 899 922 927 926
rect 931 922 983 926
rect 987 922 991 926
rect 995 922 1047 926
rect 1051 922 1095 926
rect 1099 922 1119 926
rect 103 921 1119 922
rect 1125 921 1126 927
rect 1118 919 1126 921
rect 1118 913 1119 919
rect 1125 918 2155 919
rect 1125 914 1135 918
rect 1139 914 1239 918
rect 1243 914 1287 918
rect 1291 914 1303 918
rect 1307 914 1327 918
rect 1331 914 1375 918
rect 1379 914 1423 918
rect 1427 914 1439 918
rect 1443 914 1479 918
rect 1483 914 1511 918
rect 1515 914 1551 918
rect 1555 914 1583 918
rect 1587 914 1623 918
rect 1627 914 1655 918
rect 1659 914 1703 918
rect 1707 914 1727 918
rect 1731 914 1791 918
rect 1795 914 1799 918
rect 1803 914 1871 918
rect 1875 914 1879 918
rect 1883 914 1943 918
rect 1947 914 1967 918
rect 1971 914 2015 918
rect 2019 914 2063 918
rect 2067 914 2071 918
rect 2075 914 2119 918
rect 2123 914 2155 918
rect 1125 913 2155 914
rect 2161 913 2162 919
rect 84 865 85 871
rect 91 870 1107 871
rect 91 866 111 870
rect 115 866 135 870
rect 139 866 175 870
rect 179 866 183 870
rect 187 866 215 870
rect 219 866 255 870
rect 259 866 279 870
rect 283 866 327 870
rect 331 866 343 870
rect 347 866 399 870
rect 403 866 463 870
rect 467 866 527 870
rect 531 866 535 870
rect 539 866 599 870
rect 603 866 615 870
rect 619 866 671 870
rect 675 866 711 870
rect 715 866 743 870
rect 747 866 815 870
rect 819 866 823 870
rect 827 866 895 870
rect 899 866 943 870
rect 947 866 983 870
rect 987 866 1047 870
rect 1051 866 1095 870
rect 1099 866 1107 870
rect 91 865 1107 866
rect 1113 867 1114 871
rect 1113 866 2150 867
rect 1113 865 1135 866
rect 1106 862 1135 865
rect 1139 862 1159 866
rect 1163 862 1199 866
rect 1203 862 1263 866
rect 1267 862 1287 866
rect 1291 862 1327 866
rect 1331 862 1375 866
rect 1379 862 1399 866
rect 1403 862 1423 866
rect 1427 862 1471 866
rect 1475 862 1479 866
rect 1483 862 1543 866
rect 1547 862 1551 866
rect 1555 862 1623 866
rect 1627 862 1703 866
rect 1707 862 1775 866
rect 1779 862 1791 866
rect 1795 862 1855 866
rect 1859 862 1879 866
rect 1883 862 1935 866
rect 1939 862 1967 866
rect 1971 862 2015 866
rect 2019 862 2063 866
rect 2067 862 2071 866
rect 2075 862 2119 866
rect 2123 862 2150 866
rect 1106 861 2150 862
rect 96 813 97 819
rect 103 818 1119 819
rect 103 814 111 818
rect 115 814 135 818
rect 139 814 175 818
rect 179 814 215 818
rect 219 814 279 818
rect 283 814 335 818
rect 339 814 343 818
rect 347 814 391 818
rect 395 814 399 818
rect 403 814 455 818
rect 459 814 463 818
rect 467 814 519 818
rect 523 814 535 818
rect 539 814 583 818
rect 587 814 615 818
rect 619 814 655 818
rect 659 814 711 818
rect 715 814 735 818
rect 739 814 815 818
rect 819 814 823 818
rect 827 814 895 818
rect 899 814 943 818
rect 947 814 983 818
rect 987 814 1047 818
rect 1051 814 1095 818
rect 1099 814 1119 818
rect 103 813 1119 814
rect 1125 813 1126 819
rect 1118 801 1119 807
rect 1125 806 2155 807
rect 1125 802 1135 806
rect 1139 802 1159 806
rect 1163 802 1199 806
rect 1203 802 1239 806
rect 1243 802 1263 806
rect 1267 802 1327 806
rect 1331 802 1343 806
rect 1347 802 1399 806
rect 1403 802 1447 806
rect 1451 802 1471 806
rect 1475 802 1543 806
rect 1547 802 1551 806
rect 1555 802 1623 806
rect 1627 802 1655 806
rect 1659 802 1703 806
rect 1707 802 1751 806
rect 1755 802 1775 806
rect 1779 802 1839 806
rect 1843 802 1855 806
rect 1859 802 1919 806
rect 1923 802 1935 806
rect 1939 802 2007 806
rect 2011 802 2015 806
rect 2019 802 2071 806
rect 2075 802 2119 806
rect 2123 802 2155 806
rect 1125 801 2155 802
rect 2161 801 2162 807
rect 84 761 85 767
rect 91 766 1107 767
rect 91 762 111 766
rect 115 762 135 766
rect 139 762 175 766
rect 179 762 207 766
rect 211 762 215 766
rect 219 762 279 766
rect 283 762 295 766
rect 299 762 335 766
rect 339 762 375 766
rect 379 762 391 766
rect 395 762 447 766
rect 451 762 455 766
rect 459 762 519 766
rect 523 762 583 766
rect 587 762 639 766
rect 643 762 655 766
rect 659 762 687 766
rect 691 762 735 766
rect 739 762 743 766
rect 747 762 799 766
rect 803 762 815 766
rect 819 762 855 766
rect 859 762 895 766
rect 899 762 983 766
rect 987 762 1047 766
rect 1051 762 1095 766
rect 1099 762 1107 766
rect 91 761 1107 762
rect 1113 761 1114 767
rect 1106 749 1107 755
rect 1113 754 2143 755
rect 1113 750 1135 754
rect 1139 750 1159 754
rect 1163 750 1199 754
rect 1203 750 1239 754
rect 1243 750 1287 754
rect 1291 750 1343 754
rect 1347 750 1359 754
rect 1363 750 1439 754
rect 1443 750 1447 754
rect 1451 750 1527 754
rect 1531 750 1551 754
rect 1555 750 1615 754
rect 1619 750 1655 754
rect 1659 750 1711 754
rect 1715 750 1751 754
rect 1755 750 1807 754
rect 1811 750 1839 754
rect 1843 750 1903 754
rect 1907 750 1919 754
rect 1923 750 1999 754
rect 2003 750 2007 754
rect 2011 750 2071 754
rect 2075 750 2119 754
rect 2123 750 2143 754
rect 1113 749 2143 750
rect 2149 749 2150 755
rect 96 705 97 711
rect 103 710 1119 711
rect 103 706 111 710
rect 115 706 135 710
rect 139 706 183 710
rect 187 706 207 710
rect 211 706 247 710
rect 251 706 295 710
rect 299 706 311 710
rect 315 706 375 710
rect 379 706 383 710
rect 387 706 447 710
rect 451 706 455 710
rect 459 706 519 710
rect 523 706 583 710
rect 587 706 639 710
rect 643 706 647 710
rect 651 706 687 710
rect 691 706 711 710
rect 715 706 743 710
rect 747 706 767 710
rect 771 706 799 710
rect 803 706 823 710
rect 827 706 855 710
rect 859 706 879 710
rect 883 706 943 710
rect 947 706 1095 710
rect 1099 706 1119 710
rect 103 705 1119 706
rect 1125 705 1126 711
rect 1118 693 1119 699
rect 1125 698 2155 699
rect 1125 694 1135 698
rect 1139 694 1159 698
rect 1163 694 1199 698
rect 1203 694 1239 698
rect 1243 694 1287 698
rect 1291 694 1335 698
rect 1339 694 1359 698
rect 1363 694 1391 698
rect 1395 694 1439 698
rect 1443 694 1447 698
rect 1451 694 1511 698
rect 1515 694 1527 698
rect 1531 694 1575 698
rect 1579 694 1615 698
rect 1619 694 1639 698
rect 1643 694 1703 698
rect 1707 694 1711 698
rect 1715 694 1767 698
rect 1771 694 1807 698
rect 1811 694 1831 698
rect 1835 694 1895 698
rect 1899 694 1903 698
rect 1907 694 1959 698
rect 1963 694 1999 698
rect 2003 694 2023 698
rect 2027 694 2071 698
rect 2075 694 2119 698
rect 2123 694 2155 698
rect 1125 693 2155 694
rect 2161 693 2162 699
rect 84 645 85 651
rect 91 650 1107 651
rect 91 646 111 650
rect 115 646 135 650
rect 139 646 159 650
rect 163 646 183 650
rect 187 646 215 650
rect 219 646 247 650
rect 251 646 287 650
rect 291 646 311 650
rect 315 646 367 650
rect 371 646 383 650
rect 387 646 455 650
rect 459 646 519 650
rect 523 646 543 650
rect 547 646 583 650
rect 587 646 631 650
rect 635 646 647 650
rect 651 646 711 650
rect 715 646 719 650
rect 723 646 767 650
rect 771 646 799 650
rect 803 646 823 650
rect 827 646 871 650
rect 875 646 879 650
rect 883 646 943 650
rect 947 646 951 650
rect 955 646 1031 650
rect 1035 646 1095 650
rect 1099 646 1107 650
rect 91 645 1107 646
rect 1113 647 1114 651
rect 1113 646 2150 647
rect 1113 645 1135 646
rect 1106 642 1135 645
rect 1139 642 1239 646
rect 1243 642 1279 646
rect 1283 642 1287 646
rect 1291 642 1319 646
rect 1323 642 1335 646
rect 1339 642 1367 646
rect 1371 642 1391 646
rect 1395 642 1423 646
rect 1427 642 1447 646
rect 1451 642 1479 646
rect 1483 642 1511 646
rect 1515 642 1535 646
rect 1539 642 1575 646
rect 1579 642 1591 646
rect 1595 642 1639 646
rect 1643 642 1647 646
rect 1651 642 1703 646
rect 1707 642 1719 646
rect 1723 642 1767 646
rect 1771 642 1799 646
rect 1803 642 1831 646
rect 1835 642 1879 646
rect 1883 642 1895 646
rect 1899 642 1959 646
rect 1963 642 1967 646
rect 1971 642 2023 646
rect 2027 642 2063 646
rect 2067 642 2071 646
rect 2075 642 2119 646
rect 2123 642 2150 646
rect 1106 641 2150 642
rect 96 589 97 595
rect 103 594 1119 595
rect 103 590 111 594
rect 115 590 159 594
rect 163 590 207 594
rect 211 590 215 594
rect 219 590 255 594
rect 259 590 287 594
rect 291 590 311 594
rect 315 590 367 594
rect 371 590 383 594
rect 387 590 455 594
rect 459 590 463 594
rect 467 590 543 594
rect 547 590 623 594
rect 627 590 631 594
rect 635 590 703 594
rect 707 590 719 594
rect 723 590 783 594
rect 787 590 799 594
rect 803 590 855 594
rect 859 590 871 594
rect 875 590 927 594
rect 931 590 951 594
rect 955 590 999 594
rect 1003 590 1031 594
rect 1035 590 1047 594
rect 1051 590 1095 594
rect 1099 590 1119 594
rect 103 589 1119 590
rect 1125 594 2162 595
rect 1125 590 1135 594
rect 1139 590 1279 594
rect 1283 590 1319 594
rect 1323 590 1335 594
rect 1339 590 1367 594
rect 1371 590 1375 594
rect 1379 590 1415 594
rect 1419 590 1423 594
rect 1427 590 1463 594
rect 1467 590 1479 594
rect 1483 590 1519 594
rect 1523 590 1535 594
rect 1539 590 1583 594
rect 1587 590 1591 594
rect 1595 590 1647 594
rect 1651 590 1655 594
rect 1659 590 1719 594
rect 1723 590 1727 594
rect 1731 590 1799 594
rect 1803 590 1807 594
rect 1811 590 1879 594
rect 1883 590 1887 594
rect 1891 590 1967 594
rect 1971 590 1975 594
rect 1979 590 2063 594
rect 2067 590 2119 594
rect 2123 590 2162 594
rect 1125 589 2162 590
rect 1106 538 2150 539
rect 1106 535 1135 538
rect 84 529 85 535
rect 91 534 1107 535
rect 91 530 111 534
rect 115 530 159 534
rect 163 530 167 534
rect 171 530 207 534
rect 211 530 223 534
rect 227 530 255 534
rect 259 530 287 534
rect 291 530 311 534
rect 315 530 359 534
rect 363 530 383 534
rect 387 530 431 534
rect 435 530 463 534
rect 467 530 511 534
rect 515 530 543 534
rect 547 530 591 534
rect 595 530 623 534
rect 627 530 663 534
rect 667 530 703 534
rect 707 530 735 534
rect 739 530 783 534
rect 787 530 807 534
rect 811 530 855 534
rect 859 530 871 534
rect 875 530 927 534
rect 931 530 935 534
rect 939 530 999 534
rect 1003 530 1047 534
rect 1051 530 1095 534
rect 1099 530 1107 534
rect 91 529 1107 530
rect 1113 534 1135 535
rect 1139 534 1191 538
rect 1195 534 1239 538
rect 1243 534 1287 538
rect 1291 534 1335 538
rect 1339 534 1343 538
rect 1347 534 1375 538
rect 1379 534 1407 538
rect 1411 534 1415 538
rect 1419 534 1463 538
rect 1467 534 1479 538
rect 1483 534 1519 538
rect 1523 534 1543 538
rect 1547 534 1583 538
rect 1587 534 1607 538
rect 1611 534 1655 538
rect 1659 534 1671 538
rect 1675 534 1727 538
rect 1731 534 1735 538
rect 1739 534 1799 538
rect 1803 534 1807 538
rect 1811 534 1863 538
rect 1867 534 1887 538
rect 1891 534 1935 538
rect 1939 534 1975 538
rect 1979 534 2007 538
rect 2011 534 2063 538
rect 2067 534 2071 538
rect 2075 534 2119 538
rect 2123 534 2150 538
rect 1113 533 2150 534
rect 1113 529 1114 533
rect 1118 486 2162 487
rect 1118 483 1135 486
rect 96 477 97 483
rect 103 482 1119 483
rect 103 478 111 482
rect 115 478 167 482
rect 171 478 223 482
rect 227 478 231 482
rect 235 478 287 482
rect 291 478 303 482
rect 307 478 359 482
rect 363 478 375 482
rect 379 478 431 482
rect 435 478 455 482
rect 459 478 511 482
rect 515 478 535 482
rect 539 478 591 482
rect 595 478 607 482
rect 611 478 663 482
rect 667 478 679 482
rect 683 478 735 482
rect 739 478 743 482
rect 747 478 799 482
rect 803 478 807 482
rect 811 478 855 482
rect 859 478 871 482
rect 875 478 903 482
rect 907 478 935 482
rect 939 478 959 482
rect 963 478 999 482
rect 1003 478 1007 482
rect 1011 478 1047 482
rect 1051 478 1095 482
rect 1099 478 1119 482
rect 103 477 1119 478
rect 1125 482 1135 483
rect 1139 482 1159 486
rect 1163 482 1191 486
rect 1195 482 1239 486
rect 1243 482 1263 486
rect 1267 482 1287 486
rect 1291 482 1343 486
rect 1347 482 1383 486
rect 1387 482 1407 486
rect 1411 482 1479 486
rect 1483 482 1495 486
rect 1499 482 1543 486
rect 1547 482 1599 486
rect 1603 482 1607 486
rect 1611 482 1671 486
rect 1675 482 1703 486
rect 1707 482 1735 486
rect 1739 482 1799 486
rect 1803 482 1863 486
rect 1867 482 1887 486
rect 1891 482 1935 486
rect 1939 482 1983 486
rect 1987 482 2007 486
rect 2011 482 2071 486
rect 2075 482 2119 486
rect 2123 482 2162 486
rect 1125 481 2162 482
rect 1125 477 1126 481
rect 1106 434 2150 435
rect 1106 431 1135 434
rect 84 425 85 431
rect 91 430 1107 431
rect 91 426 111 430
rect 115 426 151 430
rect 155 426 167 430
rect 171 426 215 430
rect 219 426 231 430
rect 235 426 279 430
rect 283 426 303 430
rect 307 426 351 430
rect 355 426 375 430
rect 379 426 423 430
rect 427 426 455 430
rect 459 426 487 430
rect 491 426 535 430
rect 539 426 551 430
rect 555 426 607 430
rect 611 426 615 430
rect 619 426 671 430
rect 675 426 679 430
rect 683 426 727 430
rect 731 426 743 430
rect 747 426 791 430
rect 795 426 799 430
rect 803 426 855 430
rect 859 426 903 430
rect 907 426 959 430
rect 963 426 1007 430
rect 1011 426 1047 430
rect 1051 426 1095 430
rect 1099 426 1107 430
rect 91 425 1107 426
rect 1113 430 1135 431
rect 1139 430 1159 434
rect 1163 430 1199 434
rect 1203 430 1255 434
rect 1259 430 1263 434
rect 1267 430 1335 434
rect 1339 430 1383 434
rect 1387 430 1415 434
rect 1419 430 1495 434
rect 1499 430 1503 434
rect 1507 430 1591 434
rect 1595 430 1599 434
rect 1603 430 1671 434
rect 1675 430 1703 434
rect 1707 430 1751 434
rect 1755 430 1799 434
rect 1803 430 1823 434
rect 1827 430 1887 434
rect 1891 430 1951 434
rect 1955 430 1983 434
rect 1987 430 2023 434
rect 2027 430 2071 434
rect 2075 430 2119 434
rect 2123 430 2150 434
rect 1113 429 2150 430
rect 1113 425 1114 429
rect 96 373 97 379
rect 103 378 1119 379
rect 103 374 111 378
rect 115 374 135 378
rect 139 374 151 378
rect 155 374 175 378
rect 179 374 215 378
rect 219 374 271 378
rect 275 374 279 378
rect 283 374 335 378
rect 339 374 351 378
rect 355 374 399 378
rect 403 374 423 378
rect 427 374 463 378
rect 467 374 487 378
rect 491 374 519 378
rect 523 374 551 378
rect 555 374 575 378
rect 579 374 615 378
rect 619 374 631 378
rect 635 374 671 378
rect 675 374 687 378
rect 691 374 727 378
rect 731 374 751 378
rect 755 374 791 378
rect 795 374 855 378
rect 859 374 1095 378
rect 1099 374 1119 378
rect 103 373 1119 374
rect 1125 378 2162 379
rect 1125 374 1135 378
rect 1139 374 1159 378
rect 1163 374 1199 378
rect 1203 374 1255 378
rect 1259 374 1303 378
rect 1307 374 1335 378
rect 1339 374 1343 378
rect 1347 374 1383 378
rect 1387 374 1415 378
rect 1419 374 1423 378
rect 1427 374 1463 378
rect 1467 374 1503 378
rect 1507 374 1551 378
rect 1555 374 1591 378
rect 1595 374 1615 378
rect 1619 374 1671 378
rect 1675 374 1679 378
rect 1683 374 1751 378
rect 1755 374 1823 378
rect 1827 374 1831 378
rect 1835 374 1887 378
rect 1891 374 1919 378
rect 1923 374 1951 378
rect 1955 374 2007 378
rect 2011 374 2023 378
rect 2027 374 2071 378
rect 2075 374 2119 378
rect 2123 374 2162 378
rect 1125 373 2162 374
rect 84 317 85 323
rect 91 322 1107 323
rect 91 318 111 322
rect 115 318 135 322
rect 139 318 175 322
rect 179 318 207 322
rect 211 318 215 322
rect 219 318 271 322
rect 275 318 295 322
rect 299 318 335 322
rect 339 318 383 322
rect 387 318 399 322
rect 403 318 463 322
rect 467 318 471 322
rect 475 318 519 322
rect 523 318 551 322
rect 555 318 575 322
rect 579 318 623 322
rect 627 318 631 322
rect 635 318 687 322
rect 691 318 751 322
rect 755 318 807 322
rect 811 318 871 322
rect 875 318 935 322
rect 939 318 1095 322
rect 1099 318 1107 322
rect 91 317 1107 318
rect 1113 322 2150 323
rect 1113 318 1135 322
rect 1139 318 1167 322
rect 1171 318 1207 322
rect 1211 318 1247 322
rect 1251 318 1295 322
rect 1299 318 1303 322
rect 1307 318 1343 322
rect 1347 318 1383 322
rect 1387 318 1391 322
rect 1395 318 1423 322
rect 1427 318 1439 322
rect 1443 318 1463 322
rect 1467 318 1495 322
rect 1499 318 1503 322
rect 1507 318 1551 322
rect 1555 318 1559 322
rect 1563 318 1615 322
rect 1619 318 1623 322
rect 1627 318 1679 322
rect 1683 318 1695 322
rect 1699 318 1751 322
rect 1755 318 1775 322
rect 1779 318 1831 322
rect 1835 318 1855 322
rect 1859 318 1919 322
rect 1923 318 1935 322
rect 1939 318 2007 322
rect 2011 318 2015 322
rect 2019 318 2071 322
rect 2075 318 2119 322
rect 2123 318 2150 322
rect 1113 317 2150 318
rect 96 265 97 271
rect 103 270 1119 271
rect 103 266 111 270
rect 115 266 135 270
rect 139 266 199 270
rect 203 266 207 270
rect 211 266 279 270
rect 283 266 295 270
rect 299 266 359 270
rect 363 266 383 270
rect 387 266 439 270
rect 443 266 471 270
rect 475 266 511 270
rect 515 266 551 270
rect 555 266 583 270
rect 587 266 623 270
rect 627 266 647 270
rect 651 266 687 270
rect 691 266 703 270
rect 707 266 751 270
rect 755 266 759 270
rect 763 266 807 270
rect 811 266 815 270
rect 819 266 871 270
rect 875 266 879 270
rect 883 266 935 270
rect 939 266 1095 270
rect 1099 266 1119 270
rect 103 265 1119 266
rect 1125 265 1126 271
rect 1118 263 1126 265
rect 1118 257 1119 263
rect 1125 262 2155 263
rect 1125 258 1135 262
rect 1139 258 1159 262
rect 1163 258 1167 262
rect 1171 258 1207 262
rect 1211 258 1247 262
rect 1251 258 1271 262
rect 1275 258 1295 262
rect 1299 258 1327 262
rect 1331 258 1343 262
rect 1347 258 1391 262
rect 1395 258 1439 262
rect 1443 258 1455 262
rect 1459 258 1495 262
rect 1499 258 1527 262
rect 1531 258 1559 262
rect 1563 258 1607 262
rect 1611 258 1623 262
rect 1627 258 1687 262
rect 1691 258 1695 262
rect 1699 258 1767 262
rect 1771 258 1775 262
rect 1779 258 1839 262
rect 1843 258 1855 262
rect 1859 258 1919 262
rect 1923 258 1935 262
rect 1939 258 1999 262
rect 2003 258 2015 262
rect 2019 258 2071 262
rect 2075 258 2119 262
rect 2123 258 2155 262
rect 1125 257 2155 258
rect 2161 257 2162 263
rect 84 209 85 215
rect 91 214 1107 215
rect 91 210 111 214
rect 115 210 135 214
rect 139 210 183 214
rect 187 210 199 214
rect 203 210 231 214
rect 235 210 279 214
rect 283 210 327 214
rect 331 210 359 214
rect 363 210 375 214
rect 379 210 415 214
rect 419 210 439 214
rect 443 210 455 214
rect 459 210 503 214
rect 507 210 511 214
rect 515 210 551 214
rect 555 210 583 214
rect 587 210 599 214
rect 603 210 647 214
rect 651 210 695 214
rect 699 210 703 214
rect 707 210 743 214
rect 747 210 759 214
rect 763 210 815 214
rect 819 210 879 214
rect 883 210 1095 214
rect 1099 210 1107 214
rect 91 209 1107 210
rect 1113 211 1114 215
rect 1113 210 2150 211
rect 1113 209 1135 210
rect 1106 206 1135 209
rect 1139 206 1159 210
rect 1163 206 1199 210
rect 1203 206 1207 210
rect 1211 206 1263 210
rect 1267 206 1271 210
rect 1275 206 1327 210
rect 1331 206 1391 210
rect 1395 206 1399 210
rect 1403 206 1455 210
rect 1459 206 1471 210
rect 1475 206 1527 210
rect 1531 206 1543 210
rect 1547 206 1607 210
rect 1611 206 1671 210
rect 1675 206 1687 210
rect 1691 206 1735 210
rect 1739 206 1767 210
rect 1771 206 1807 210
rect 1811 206 1839 210
rect 1843 206 1879 210
rect 1883 206 1919 210
rect 1923 206 1951 210
rect 1955 206 1999 210
rect 2003 206 2023 210
rect 2027 206 2071 210
rect 2075 206 2119 210
rect 2123 206 2150 210
rect 1106 205 2150 206
rect 96 133 97 139
rect 103 138 1119 139
rect 103 134 111 138
rect 115 134 135 138
rect 139 134 143 138
rect 147 134 183 138
rect 187 134 223 138
rect 227 134 231 138
rect 235 134 263 138
rect 267 134 279 138
rect 283 134 303 138
rect 307 134 327 138
rect 331 134 343 138
rect 347 134 375 138
rect 379 134 383 138
rect 387 134 415 138
rect 419 134 423 138
rect 427 134 455 138
rect 459 134 463 138
rect 467 134 503 138
rect 507 134 543 138
rect 547 134 551 138
rect 555 134 583 138
rect 587 134 599 138
rect 603 134 623 138
rect 627 134 647 138
rect 651 134 663 138
rect 667 134 695 138
rect 699 134 703 138
rect 707 134 743 138
rect 747 134 783 138
rect 787 134 831 138
rect 835 134 879 138
rect 883 134 927 138
rect 931 134 967 138
rect 971 134 1007 138
rect 1011 134 1047 138
rect 1051 134 1095 138
rect 1099 134 1119 138
rect 103 133 1119 134
rect 1125 138 2162 139
rect 1125 134 1135 138
rect 1139 134 1159 138
rect 1163 134 1199 138
rect 1203 134 1207 138
rect 1211 134 1263 138
rect 1267 134 1271 138
rect 1275 134 1327 138
rect 1331 134 1335 138
rect 1339 134 1399 138
rect 1403 134 1455 138
rect 1459 134 1471 138
rect 1475 134 1511 138
rect 1515 134 1543 138
rect 1547 134 1559 138
rect 1563 134 1607 138
rect 1611 134 1647 138
rect 1651 134 1671 138
rect 1675 134 1687 138
rect 1691 134 1727 138
rect 1731 134 1735 138
rect 1739 134 1767 138
rect 1771 134 1807 138
rect 1811 134 1855 138
rect 1859 134 1879 138
rect 1883 134 1903 138
rect 1907 134 1951 138
rect 1955 134 1991 138
rect 1995 134 2023 138
rect 2027 134 2031 138
rect 2035 134 2071 138
rect 2075 134 2119 138
rect 2123 134 2162 138
rect 1125 133 2162 134
rect 84 81 85 87
rect 91 86 1107 87
rect 91 82 111 86
rect 115 82 143 86
rect 147 82 183 86
rect 187 82 223 86
rect 227 82 263 86
rect 267 82 303 86
rect 307 82 343 86
rect 347 82 383 86
rect 387 82 423 86
rect 427 82 463 86
rect 467 82 503 86
rect 507 82 543 86
rect 547 82 583 86
rect 587 82 623 86
rect 627 82 663 86
rect 667 82 703 86
rect 707 82 743 86
rect 747 82 783 86
rect 787 82 831 86
rect 835 82 879 86
rect 883 82 927 86
rect 931 82 967 86
rect 971 82 1007 86
rect 1011 82 1047 86
rect 1051 82 1095 86
rect 1099 82 1107 86
rect 91 81 1107 82
rect 1113 86 2150 87
rect 1113 82 1135 86
rect 1139 82 1159 86
rect 1163 82 1207 86
rect 1211 82 1271 86
rect 1275 82 1335 86
rect 1339 82 1399 86
rect 1403 82 1455 86
rect 1459 82 1511 86
rect 1515 82 1559 86
rect 1563 82 1607 86
rect 1611 82 1647 86
rect 1651 82 1687 86
rect 1691 82 1727 86
rect 1731 82 1767 86
rect 1771 82 1807 86
rect 1811 82 1855 86
rect 1859 82 1903 86
rect 1907 82 1951 86
rect 1955 82 1991 86
rect 1995 82 2031 86
rect 2035 82 2071 86
rect 2075 82 2119 86
rect 2123 82 2150 86
rect 1113 81 2150 82
<< m5c >>
rect 1119 2225 1125 2231
rect 2155 2225 2161 2231
rect 85 2209 91 2215
rect 1107 2209 1113 2215
rect 1107 2173 1113 2179
rect 2143 2173 2149 2179
rect 97 2149 103 2155
rect 1119 2149 1125 2155
rect 1119 2121 1125 2127
rect 2155 2121 2161 2127
rect 85 2093 91 2099
rect 1107 2093 1113 2099
rect 1107 2069 1113 2075
rect 2143 2069 2149 2075
rect 97 2037 103 2043
rect 1119 2037 1125 2043
rect 1119 2017 1125 2023
rect 2155 2017 2161 2023
rect 85 1985 91 1991
rect 1107 1985 1113 1991
rect 1107 1953 1113 1959
rect 2143 1953 2149 1959
rect 97 1929 103 1935
rect 1119 1929 1125 1935
rect 1119 1901 1125 1907
rect 2155 1901 2161 1907
rect 85 1873 91 1879
rect 1107 1873 1113 1879
rect 1107 1845 1113 1851
rect 2143 1845 2149 1851
rect 97 1817 103 1823
rect 1119 1817 1125 1823
rect 1119 1785 1125 1791
rect 2155 1785 2161 1791
rect 85 1757 91 1763
rect 1107 1757 1113 1763
rect 1107 1729 1113 1735
rect 2143 1729 2149 1735
rect 97 1701 103 1707
rect 1119 1701 1125 1707
rect 1119 1677 1125 1683
rect 2155 1677 2161 1683
rect 85 1645 91 1651
rect 1107 1645 1113 1651
rect 1107 1621 1113 1627
rect 2143 1621 2149 1627
rect 97 1585 103 1591
rect 1119 1585 1125 1591
rect 1119 1569 1125 1575
rect 2155 1569 2161 1575
rect 85 1525 91 1531
rect 1107 1525 1113 1531
rect 1107 1513 1113 1519
rect 2143 1513 2149 1519
rect 97 1465 103 1471
rect 1119 1465 1125 1471
rect 85 1409 91 1415
rect 1107 1409 1113 1415
rect 97 1357 103 1363
rect 1119 1357 1125 1363
rect 1119 1349 1125 1355
rect 2155 1349 2161 1355
rect 85 1305 91 1311
rect 1107 1305 1113 1311
rect 1107 1293 1113 1299
rect 2143 1293 2149 1299
rect 97 1249 103 1255
rect 1119 1249 1125 1255
rect 1119 1237 1125 1243
rect 2155 1237 2161 1243
rect 85 1197 91 1203
rect 1107 1197 1113 1203
rect 1107 1185 1113 1191
rect 2143 1185 2149 1191
rect 97 1145 103 1151
rect 1119 1145 1125 1151
rect 1119 1125 1125 1131
rect 2155 1125 2161 1131
rect 85 1085 91 1091
rect 1107 1085 1113 1091
rect 1107 1073 1113 1079
rect 2143 1073 2149 1079
rect 97 1029 103 1035
rect 1119 1029 1125 1035
rect 1119 1021 1125 1027
rect 2155 1021 2161 1027
rect 85 973 91 979
rect 1107 973 1113 979
rect 97 921 103 927
rect 1119 921 1125 927
rect 1119 913 1125 919
rect 2155 913 2161 919
rect 85 865 91 871
rect 1107 865 1113 871
rect 97 813 103 819
rect 1119 813 1125 819
rect 1119 801 1125 807
rect 2155 801 2161 807
rect 85 761 91 767
rect 1107 761 1113 767
rect 1107 749 1113 755
rect 2143 749 2149 755
rect 97 705 103 711
rect 1119 705 1125 711
rect 1119 693 1125 699
rect 2155 693 2161 699
rect 85 645 91 651
rect 1107 645 1113 651
rect 97 589 103 595
rect 1119 589 1125 595
rect 85 529 91 535
rect 1107 529 1113 535
rect 97 477 103 483
rect 1119 477 1125 483
rect 85 425 91 431
rect 1107 425 1113 431
rect 97 373 103 379
rect 1119 373 1125 379
rect 85 317 91 323
rect 1107 317 1113 323
rect 97 265 103 271
rect 1119 265 1125 271
rect 1119 257 1125 263
rect 2155 257 2161 263
rect 85 209 91 215
rect 1107 209 1113 215
rect 97 133 103 139
rect 1119 133 1125 139
rect 85 81 91 87
rect 1107 81 1113 87
<< m5 >>
rect 84 2215 92 2232
rect 84 2209 85 2215
rect 91 2209 92 2215
rect 84 2099 92 2209
rect 84 2093 85 2099
rect 91 2093 92 2099
rect 84 1991 92 2093
rect 84 1985 85 1991
rect 91 1985 92 1991
rect 84 1879 92 1985
rect 84 1873 85 1879
rect 91 1873 92 1879
rect 84 1763 92 1873
rect 84 1757 85 1763
rect 91 1757 92 1763
rect 84 1651 92 1757
rect 84 1645 85 1651
rect 91 1645 92 1651
rect 84 1531 92 1645
rect 84 1525 85 1531
rect 91 1525 92 1531
rect 84 1415 92 1525
rect 84 1409 85 1415
rect 91 1409 92 1415
rect 84 1311 92 1409
rect 84 1305 85 1311
rect 91 1305 92 1311
rect 84 1203 92 1305
rect 84 1197 85 1203
rect 91 1197 92 1203
rect 84 1091 92 1197
rect 84 1085 85 1091
rect 91 1085 92 1091
rect 84 979 92 1085
rect 84 973 85 979
rect 91 973 92 979
rect 84 871 92 973
rect 84 865 85 871
rect 91 865 92 871
rect 84 767 92 865
rect 84 761 85 767
rect 91 761 92 767
rect 84 651 92 761
rect 84 645 85 651
rect 91 645 92 651
rect 84 535 92 645
rect 84 529 85 535
rect 91 529 92 535
rect 84 431 92 529
rect 84 425 85 431
rect 91 425 92 431
rect 84 323 92 425
rect 84 317 85 323
rect 91 317 92 323
rect 84 215 92 317
rect 84 209 85 215
rect 91 209 92 215
rect 84 87 92 209
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2155 104 2232
rect 96 2149 97 2155
rect 103 2149 104 2155
rect 96 2043 104 2149
rect 96 2037 97 2043
rect 103 2037 104 2043
rect 96 1935 104 2037
rect 96 1929 97 1935
rect 103 1929 104 1935
rect 96 1823 104 1929
rect 96 1817 97 1823
rect 103 1817 104 1823
rect 96 1707 104 1817
rect 96 1701 97 1707
rect 103 1701 104 1707
rect 96 1591 104 1701
rect 96 1585 97 1591
rect 103 1585 104 1591
rect 96 1471 104 1585
rect 96 1465 97 1471
rect 103 1465 104 1471
rect 96 1363 104 1465
rect 96 1357 97 1363
rect 103 1357 104 1363
rect 96 1255 104 1357
rect 96 1249 97 1255
rect 103 1249 104 1255
rect 96 1151 104 1249
rect 96 1145 97 1151
rect 103 1145 104 1151
rect 96 1035 104 1145
rect 96 1029 97 1035
rect 103 1029 104 1035
rect 96 927 104 1029
rect 96 921 97 927
rect 103 921 104 927
rect 96 819 104 921
rect 96 813 97 819
rect 103 813 104 819
rect 96 711 104 813
rect 96 705 97 711
rect 103 705 104 711
rect 96 595 104 705
rect 96 589 97 595
rect 103 589 104 595
rect 96 483 104 589
rect 96 477 97 483
rect 103 477 104 483
rect 96 379 104 477
rect 96 373 97 379
rect 103 373 104 379
rect 96 271 104 373
rect 96 265 97 271
rect 103 265 104 271
rect 96 139 104 265
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1106 2215 1114 2232
rect 1106 2209 1107 2215
rect 1113 2209 1114 2215
rect 1106 2179 1114 2209
rect 1106 2173 1107 2179
rect 1113 2173 1114 2179
rect 1106 2099 1114 2173
rect 1106 2093 1107 2099
rect 1113 2093 1114 2099
rect 1106 2075 1114 2093
rect 1106 2069 1107 2075
rect 1113 2069 1114 2075
rect 1106 1991 1114 2069
rect 1106 1985 1107 1991
rect 1113 1985 1114 1991
rect 1106 1959 1114 1985
rect 1106 1953 1107 1959
rect 1113 1953 1114 1959
rect 1106 1879 1114 1953
rect 1106 1873 1107 1879
rect 1113 1873 1114 1879
rect 1106 1851 1114 1873
rect 1106 1845 1107 1851
rect 1113 1845 1114 1851
rect 1106 1763 1114 1845
rect 1106 1757 1107 1763
rect 1113 1757 1114 1763
rect 1106 1735 1114 1757
rect 1106 1729 1107 1735
rect 1113 1729 1114 1735
rect 1106 1651 1114 1729
rect 1106 1645 1107 1651
rect 1113 1645 1114 1651
rect 1106 1627 1114 1645
rect 1106 1621 1107 1627
rect 1113 1621 1114 1627
rect 1106 1531 1114 1621
rect 1106 1525 1107 1531
rect 1113 1525 1114 1531
rect 1106 1519 1114 1525
rect 1106 1513 1107 1519
rect 1113 1513 1114 1519
rect 1106 1415 1114 1513
rect 1106 1409 1107 1415
rect 1113 1409 1114 1415
rect 1106 1311 1114 1409
rect 1106 1305 1107 1311
rect 1113 1305 1114 1311
rect 1106 1299 1114 1305
rect 1106 1293 1107 1299
rect 1113 1293 1114 1299
rect 1106 1203 1114 1293
rect 1106 1197 1107 1203
rect 1113 1197 1114 1203
rect 1106 1191 1114 1197
rect 1106 1185 1107 1191
rect 1113 1185 1114 1191
rect 1106 1091 1114 1185
rect 1106 1085 1107 1091
rect 1113 1085 1114 1091
rect 1106 1079 1114 1085
rect 1106 1073 1107 1079
rect 1113 1073 1114 1079
rect 1106 979 1114 1073
rect 1106 973 1107 979
rect 1113 973 1114 979
rect 1106 871 1114 973
rect 1106 865 1107 871
rect 1113 865 1114 871
rect 1106 767 1114 865
rect 1106 761 1107 767
rect 1113 761 1114 767
rect 1106 755 1114 761
rect 1106 749 1107 755
rect 1113 749 1114 755
rect 1106 651 1114 749
rect 1106 645 1107 651
rect 1113 645 1114 651
rect 1106 535 1114 645
rect 1106 529 1107 535
rect 1113 529 1114 535
rect 1106 431 1114 529
rect 1106 425 1107 431
rect 1113 425 1114 431
rect 1106 323 1114 425
rect 1106 317 1107 323
rect 1113 317 1114 323
rect 1106 215 1114 317
rect 1106 209 1107 215
rect 1113 209 1114 215
rect 1106 87 1114 209
rect 1106 81 1107 87
rect 1113 81 1114 87
rect 1106 72 1114 81
rect 1118 2231 1126 2232
rect 1118 2225 1119 2231
rect 1125 2225 1126 2231
rect 1118 2155 1126 2225
rect 1118 2149 1119 2155
rect 1125 2149 1126 2155
rect 1118 2127 1126 2149
rect 1118 2121 1119 2127
rect 1125 2121 1126 2127
rect 1118 2043 1126 2121
rect 1118 2037 1119 2043
rect 1125 2037 1126 2043
rect 1118 2023 1126 2037
rect 1118 2017 1119 2023
rect 1125 2017 1126 2023
rect 1118 1935 1126 2017
rect 1118 1929 1119 1935
rect 1125 1929 1126 1935
rect 1118 1907 1126 1929
rect 1118 1901 1119 1907
rect 1125 1901 1126 1907
rect 1118 1823 1126 1901
rect 1118 1817 1119 1823
rect 1125 1817 1126 1823
rect 1118 1791 1126 1817
rect 1118 1785 1119 1791
rect 1125 1785 1126 1791
rect 1118 1707 1126 1785
rect 1118 1701 1119 1707
rect 1125 1701 1126 1707
rect 1118 1683 1126 1701
rect 1118 1677 1119 1683
rect 1125 1677 1126 1683
rect 1118 1591 1126 1677
rect 1118 1585 1119 1591
rect 1125 1585 1126 1591
rect 1118 1575 1126 1585
rect 1118 1569 1119 1575
rect 1125 1569 1126 1575
rect 1118 1471 1126 1569
rect 1118 1465 1119 1471
rect 1125 1465 1126 1471
rect 1118 1363 1126 1465
rect 1118 1357 1119 1363
rect 1125 1357 1126 1363
rect 1118 1355 1126 1357
rect 1118 1349 1119 1355
rect 1125 1349 1126 1355
rect 1118 1255 1126 1349
rect 1118 1249 1119 1255
rect 1125 1249 1126 1255
rect 1118 1243 1126 1249
rect 1118 1237 1119 1243
rect 1125 1237 1126 1243
rect 1118 1151 1126 1237
rect 1118 1145 1119 1151
rect 1125 1145 1126 1151
rect 1118 1131 1126 1145
rect 1118 1125 1119 1131
rect 1125 1125 1126 1131
rect 1118 1035 1126 1125
rect 1118 1029 1119 1035
rect 1125 1029 1126 1035
rect 1118 1027 1126 1029
rect 1118 1021 1119 1027
rect 1125 1021 1126 1027
rect 1118 927 1126 1021
rect 1118 921 1119 927
rect 1125 921 1126 927
rect 1118 919 1126 921
rect 1118 913 1119 919
rect 1125 913 1126 919
rect 1118 819 1126 913
rect 1118 813 1119 819
rect 1125 813 1126 819
rect 1118 807 1126 813
rect 1118 801 1119 807
rect 1125 801 1126 807
rect 1118 711 1126 801
rect 1118 705 1119 711
rect 1125 705 1126 711
rect 1118 699 1126 705
rect 1118 693 1119 699
rect 1125 693 1126 699
rect 1118 595 1126 693
rect 1118 589 1119 595
rect 1125 589 1126 595
rect 1118 483 1126 589
rect 1118 477 1119 483
rect 1125 477 1126 483
rect 1118 379 1126 477
rect 1118 373 1119 379
rect 1125 373 1126 379
rect 1118 271 1126 373
rect 1118 265 1119 271
rect 1125 265 1126 271
rect 1118 263 1126 265
rect 1118 257 1119 263
rect 1125 257 1126 263
rect 1118 139 1126 257
rect 1118 133 1119 139
rect 1125 133 1126 139
rect 1118 72 1126 133
rect 2142 2179 2150 2232
rect 2142 2173 2143 2179
rect 2149 2173 2150 2179
rect 2142 2075 2150 2173
rect 2142 2069 2143 2075
rect 2149 2069 2150 2075
rect 2142 1959 2150 2069
rect 2142 1953 2143 1959
rect 2149 1953 2150 1959
rect 2142 1851 2150 1953
rect 2142 1845 2143 1851
rect 2149 1845 2150 1851
rect 2142 1735 2150 1845
rect 2142 1729 2143 1735
rect 2149 1729 2150 1735
rect 2142 1627 2150 1729
rect 2142 1621 2143 1627
rect 2149 1621 2150 1627
rect 2142 1519 2150 1621
rect 2142 1513 2143 1519
rect 2149 1513 2150 1519
rect 2142 1299 2150 1513
rect 2142 1293 2143 1299
rect 2149 1293 2150 1299
rect 2142 1191 2150 1293
rect 2142 1185 2143 1191
rect 2149 1185 2150 1191
rect 2142 1079 2150 1185
rect 2142 1073 2143 1079
rect 2149 1073 2150 1079
rect 2142 755 2150 1073
rect 2142 749 2143 755
rect 2149 749 2150 755
rect 2142 72 2150 749
rect 2154 2231 2162 2232
rect 2154 2225 2155 2231
rect 2161 2225 2162 2231
rect 2154 2127 2162 2225
rect 2154 2121 2155 2127
rect 2161 2121 2162 2127
rect 2154 2023 2162 2121
rect 2154 2017 2155 2023
rect 2161 2017 2162 2023
rect 2154 1907 2162 2017
rect 2154 1901 2155 1907
rect 2161 1901 2162 1907
rect 2154 1791 2162 1901
rect 2154 1785 2155 1791
rect 2161 1785 2162 1791
rect 2154 1683 2162 1785
rect 2154 1677 2155 1683
rect 2161 1677 2162 1683
rect 2154 1575 2162 1677
rect 2154 1569 2155 1575
rect 2161 1569 2162 1575
rect 2154 1355 2162 1569
rect 2154 1349 2155 1355
rect 2161 1349 2162 1355
rect 2154 1243 2162 1349
rect 2154 1237 2155 1243
rect 2161 1237 2162 1243
rect 2154 1131 2162 1237
rect 2154 1125 2155 1131
rect 2161 1125 2162 1131
rect 2154 1027 2162 1125
rect 2154 1021 2155 1027
rect 2161 1021 2162 1027
rect 2154 919 2162 1021
rect 2154 913 2155 919
rect 2161 913 2162 919
rect 2154 807 2162 913
rect 2154 801 2155 807
rect 2161 801 2162 807
rect 2154 699 2162 801
rect 2154 693 2155 699
rect 2161 693 2162 699
rect 2154 263 2162 693
rect 2154 257 2155 263
rect 2161 257 2162 263
rect 2154 72 2162 257
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__153
timestamp 1731220618
transform 1 0 2112 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220618
transform 1 0 1128 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220618
transform 1 0 2112 0 -1 2172
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220618
transform 1 0 1128 0 -1 2172
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220618
transform 1 0 2112 0 1 2076
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220618
transform 1 0 1128 0 1 2076
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220618
transform 1 0 2112 0 -1 2068
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220618
transform 1 0 1128 0 -1 2068
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220618
transform 1 0 2112 0 1 1972
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220618
transform 1 0 1128 0 1 1972
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220618
transform 1 0 2112 0 -1 1952
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220618
transform 1 0 1128 0 -1 1952
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220618
transform 1 0 2112 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220618
transform 1 0 1128 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220618
transform 1 0 2112 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220618
transform 1 0 1128 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220618
transform 1 0 2112 0 1 1740
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220618
transform 1 0 1128 0 1 1740
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220618
transform 1 0 2112 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220618
transform 1 0 1128 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220618
transform 1 0 2112 0 1 1632
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220618
transform 1 0 1128 0 1 1632
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220618
transform 1 0 2112 0 -1 1620
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220618
transform 1 0 1128 0 -1 1620
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220618
transform 1 0 2112 0 1 1524
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220618
transform 1 0 1128 0 1 1524
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220618
transform 1 0 2112 0 -1 1512
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220618
transform 1 0 1128 0 -1 1512
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220618
transform 1 0 2112 0 1 1416
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220618
transform 1 0 1128 0 1 1416
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220618
transform 1 0 2112 0 -1 1404
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220618
transform 1 0 1128 0 -1 1404
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220618
transform 1 0 2112 0 1 1304
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220618
transform 1 0 1128 0 1 1304
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220618
transform 1 0 2112 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220618
transform 1 0 1128 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220618
transform 1 0 2112 0 1 1192
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220618
transform 1 0 1128 0 1 1192
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220618
transform 1 0 2112 0 -1 1184
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220618
transform 1 0 1128 0 -1 1184
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220618
transform 1 0 2112 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220618
transform 1 0 1128 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220618
transform 1 0 2112 0 -1 1072
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220618
transform 1 0 1128 0 -1 1072
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220618
transform 1 0 2112 0 1 976
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220618
transform 1 0 1128 0 1 976
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220618
transform 1 0 2112 0 -1 968
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220618
transform 1 0 1128 0 -1 968
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220618
transform 1 0 2112 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220618
transform 1 0 1128 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220618
transform 1 0 2112 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220618
transform 1 0 1128 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220618
transform 1 0 2112 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220618
transform 1 0 1128 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220618
transform 1 0 2112 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220618
transform 1 0 1128 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220618
transform 1 0 2112 0 1 648
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220618
transform 1 0 1128 0 1 648
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220618
transform 1 0 2112 0 -1 640
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220618
transform 1 0 1128 0 -1 640
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220618
transform 1 0 2112 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220618
transform 1 0 1128 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220618
transform 1 0 2112 0 -1 532
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220618
transform 1 0 1128 0 -1 532
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220618
transform 1 0 2112 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220618
transform 1 0 1128 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220618
transform 1 0 2112 0 -1 428
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220618
transform 1 0 1128 0 -1 428
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220618
transform 1 0 2112 0 1 328
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220618
transform 1 0 1128 0 1 328
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220618
transform 1 0 2112 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220618
transform 1 0 1128 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220618
transform 1 0 2112 0 1 212
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220618
transform 1 0 1128 0 1 212
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220618
transform 1 0 2112 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220618
transform 1 0 1128 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220618
transform 1 0 2112 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220618
transform 1 0 1128 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220618
transform 1 0 1088 0 -1 2208
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220618
transform 1 0 104 0 -1 2208
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220618
transform 1 0 1088 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220618
transform 1 0 104 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220618
transform 1 0 1088 0 -1 2092
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220618
transform 1 0 104 0 -1 2092
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220618
transform 1 0 1088 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220618
transform 1 0 104 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220618
transform 1 0 1088 0 -1 1984
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220618
transform 1 0 104 0 -1 1984
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220618
transform 1 0 1088 0 1 1884
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220618
transform 1 0 104 0 1 1884
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220618
transform 1 0 1088 0 -1 1872
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220618
transform 1 0 104 0 -1 1872
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220618
transform 1 0 1088 0 1 1772
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220618
transform 1 0 104 0 1 1772
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220618
transform 1 0 1088 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220618
transform 1 0 104 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220618
transform 1 0 1088 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220618
transform 1 0 104 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220618
transform 1 0 1088 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220618
transform 1 0 104 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220618
transform 1 0 1088 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220618
transform 1 0 104 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220618
transform 1 0 1088 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220618
transform 1 0 104 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220618
transform 1 0 1088 0 1 1420
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220618
transform 1 0 104 0 1 1420
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220618
transform 1 0 1088 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220618
transform 1 0 104 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220618
transform 1 0 1088 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220618
transform 1 0 104 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220618
transform 1 0 1088 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220618
transform 1 0 104 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220618
transform 1 0 1088 0 1 1204
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220618
transform 1 0 104 0 1 1204
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220618
transform 1 0 1088 0 -1 1196
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220618
transform 1 0 104 0 -1 1196
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220618
transform 1 0 1088 0 1 1100
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220618
transform 1 0 104 0 1 1100
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220618
transform 1 0 1088 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220618
transform 1 0 104 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220618
transform 1 0 1088 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220618
transform 1 0 104 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220618
transform 1 0 1088 0 -1 972
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220618
transform 1 0 104 0 -1 972
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220618
transform 1 0 1088 0 1 876
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220618
transform 1 0 104 0 1 876
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220618
transform 1 0 1088 0 -1 864
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220618
transform 1 0 104 0 -1 864
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220618
transform 1 0 1088 0 1 768
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220618
transform 1 0 104 0 1 768
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220618
transform 1 0 1088 0 -1 760
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220618
transform 1 0 104 0 -1 760
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220618
transform 1 0 1088 0 1 660
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220618
transform 1 0 104 0 1 660
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220618
transform 1 0 1088 0 -1 644
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220618
transform 1 0 104 0 -1 644
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220618
transform 1 0 1088 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220618
transform 1 0 104 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220618
transform 1 0 1088 0 -1 528
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220618
transform 1 0 104 0 -1 528
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220618
transform 1 0 1088 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220618
transform 1 0 104 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220618
transform 1 0 1088 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220618
transform 1 0 104 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220618
transform 1 0 1088 0 1 328
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220618
transform 1 0 104 0 1 328
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220618
transform 1 0 1088 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220618
transform 1 0 104 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220618
transform 1 0 1088 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220618
transform 1 0 104 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220618
transform 1 0 1088 0 -1 208
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220618
transform 1 0 104 0 -1 208
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220618
transform 1 0 1088 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220618
transform 1 0 104 0 1 88
box 7 3 12 24
use _0_0std_0_0cells_0_0NOR2X1  tst_5999_6
timestamp 1731220618
transform 1 0 1984 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5998_6
timestamp 1731220618
transform 1 0 2024 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5997_6
timestamp 1731220618
transform 1 0 2064 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5996_6
timestamp 1731220618
transform 1 0 2064 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5995_6
timestamp 1731220618
transform 1 0 2064 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5994_6
timestamp 1731220618
transform 1 0 1992 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5993_6
timestamp 1731220618
transform 1 0 2008 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5992_6
timestamp 1731220618
transform 1 0 2064 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5991_6
timestamp 1731220618
transform 1 0 2064 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5990_6
timestamp 1731220618
transform 1 0 2064 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5989_6
timestamp 1731220618
transform 1 0 2016 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5988_6
timestamp 1731220618
transform 1 0 2064 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5987_6
timestamp 1731220618
transform 1 0 2064 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5986_6
timestamp 1731220618
transform 1 0 2000 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5985_6
timestamp 1731220618
transform 1 0 1968 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5984_6
timestamp 1731220618
transform 1 0 2056 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5983_6
timestamp 1731220618
transform 1 0 2056 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5982_6
timestamp 1731220618
transform 1 0 2016 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5981_6
timestamp 1731220618
transform 1 0 2064 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5980_6
timestamp 1731220618
transform 1 0 2064 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5979_6
timestamp 1731220618
transform 1 0 2064 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5978_6
timestamp 1731220618
transform 1 0 2064 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5977_6
timestamp 1731220618
transform 1 0 2008 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5976_6
timestamp 1731220618
transform 1 0 1936 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5975_6
timestamp 1731220618
transform 1 0 2008 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5974_6
timestamp 1731220618
transform 1 0 2064 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5973_6
timestamp 1731220618
transform 1 0 2056 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5972_6
timestamp 1731220618
transform 1 0 1960 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5971_6
timestamp 1731220618
transform 1 0 1872 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5970_6
timestamp 1731220618
transform 1 0 1848 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5969_6
timestamp 1731220618
transform 1 0 1928 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5968_6
timestamp 1731220618
transform 1 0 2000 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5967_6
timestamp 1731220618
transform 1 0 1912 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5966_6
timestamp 1731220618
transform 1 0 1832 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5965_6
timestamp 1731220618
transform 1 0 1800 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5964_6
timestamp 1731220618
transform 1 0 1896 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5963_6
timestamp 1731220618
transform 1 0 1992 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5962_6
timestamp 1731220618
transform 1 0 1952 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5961_6
timestamp 1731220618
transform 1 0 1888 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5960_6
timestamp 1731220618
transform 1 0 1824 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5959_6
timestamp 1731220618
transform 1 0 1760 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5958_6
timestamp 1731220618
transform 1 0 1696 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5957_6
timestamp 1731220618
transform 1 0 1960 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5956_6
timestamp 1731220618
transform 1 0 1872 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5955_6
timestamp 1731220618
transform 1 0 1792 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5954_6
timestamp 1731220618
transform 1 0 1712 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5953_6
timestamp 1731220618
transform 1 0 1640 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5952_6
timestamp 1731220618
transform 1 0 1584 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5951_6
timestamp 1731220618
transform 1 0 1720 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5950_6
timestamp 1731220618
transform 1 0 1800 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5949_6
timestamp 1731220618
transform 1 0 1880 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5948_6
timestamp 1731220618
transform 1 0 1856 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5947_6
timestamp 1731220618
transform 1 0 1792 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5946_6
timestamp 1731220618
transform 1 0 1728 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5945_6
timestamp 1731220618
transform 1 0 1928 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5944_6
timestamp 1731220618
transform 1 0 1976 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5943_6
timestamp 1731220618
transform 1 0 1880 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5942_6
timestamp 1731220618
transform 1 0 1792 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5941_6
timestamp 1731220618
transform 1 0 1816 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5940_6
timestamp 1731220618
transform 1 0 1880 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5939_6
timestamp 1731220618
transform 1 0 1944 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5938_6
timestamp 1731220618
transform 1 0 2000 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5937_6
timestamp 1731220618
transform 1 0 1912 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5936_6
timestamp 1731220618
transform 1 0 1928 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5935_6
timestamp 1731220618
transform 1 0 1848 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5934_6
timestamp 1731220618
transform 1 0 1832 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5933_6
timestamp 1731220618
transform 1 0 1912 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5932_6
timestamp 1731220618
transform 1 0 2016 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5931_6
timestamp 1731220618
transform 1 0 1944 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5930_6
timestamp 1731220618
transform 1 0 1872 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5929_6
timestamp 1731220618
transform 1 0 1800 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5928_6
timestamp 1731220618
transform 1 0 1944 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5927_6
timestamp 1731220618
transform 1 0 1896 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5926_6
timestamp 1731220618
transform 1 0 1848 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5925_6
timestamp 1731220618
transform 1 0 1800 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5924_6
timestamp 1731220618
transform 1 0 1760 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5923_6
timestamp 1731220618
transform 1 0 1720 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5922_6
timestamp 1731220618
transform 1 0 1680 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5921_6
timestamp 1731220618
transform 1 0 1640 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5920_6
timestamp 1731220618
transform 1 0 1600 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5919_6
timestamp 1731220618
transform 1 0 1552 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5918_6
timestamp 1731220618
transform 1 0 1600 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5917_6
timestamp 1731220618
transform 1 0 1664 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5916_6
timestamp 1731220618
transform 1 0 1728 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5915_6
timestamp 1731220618
transform 1 0 1760 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5914_6
timestamp 1731220618
transform 1 0 1680 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5913_6
timestamp 1731220618
transform 1 0 1600 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5912_6
timestamp 1731220618
transform 1 0 1688 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5911_6
timestamp 1731220618
transform 1 0 1768 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5910_6
timestamp 1731220618
transform 1 0 1824 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5909_6
timestamp 1731220618
transform 1 0 1744 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5908_6
timestamp 1731220618
transform 1 0 1664 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5907_6
timestamp 1731220618
transform 1 0 1584 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5906_6
timestamp 1731220618
transform 1 0 1488 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5905_6
timestamp 1731220618
transform 1 0 1592 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5904_6
timestamp 1731220618
transform 1 0 1696 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5903_6
timestamp 1731220618
transform 1 0 1664 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5902_6
timestamp 1731220618
transform 1 0 1600 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5901_6
timestamp 1731220618
transform 1 0 1536 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5900_6
timestamp 1731220618
transform 1 0 1648 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5899_6
timestamp 1731220618
transform 1 0 1576 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5898_6
timestamp 1731220618
transform 1 0 1528 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5897_6
timestamp 1731220618
transform 1 0 1472 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5896_6
timestamp 1731220618
transform 1 0 1440 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5895_6
timestamp 1731220618
transform 1 0 1384 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5894_6
timestamp 1731220618
transform 1 0 1504 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5893_6
timestamp 1731220618
transform 1 0 1568 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5892_6
timestamp 1731220618
transform 1 0 1632 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5891_6
timestamp 1731220618
transform 1 0 1704 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5890_6
timestamp 1731220618
transform 1 0 1608 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5889_6
timestamp 1731220618
transform 1 0 1520 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5888_6
timestamp 1731220618
transform 1 0 1440 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5887_6
timestamp 1731220618
transform 1 0 1544 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5886_6
timestamp 1731220618
transform 1 0 1648 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5885_6
timestamp 1731220618
transform 1 0 1744 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5884_6
timestamp 1731220618
transform 1 0 1768 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5883_6
timestamp 1731220618
transform 1 0 1696 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5882_6
timestamp 1731220618
transform 1 0 1616 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5881_6
timestamp 1731220618
transform 1 0 1536 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5880_6
timestamp 1731220618
transform 1 0 1544 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5879_6
timestamp 1731220618
transform 1 0 1616 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5878_6
timestamp 1731220618
transform 1 0 1696 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5877_6
timestamp 1731220618
transform 1 0 1784 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5876_6
timestamp 1731220618
transform 1 0 1720 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5875_6
timestamp 1731220618
transform 1 0 1648 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5874_6
timestamp 1731220618
transform 1 0 1576 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5873_6
timestamp 1731220618
transform 1 0 1864 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5872_6
timestamp 1731220618
transform 1 0 1792 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5871_6
timestamp 1731220618
transform 1 0 1752 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5870_6
timestamp 1731220618
transform 1 0 1688 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5869_6
timestamp 1731220618
transform 1 0 1616 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5868_6
timestamp 1731220618
transform 1 0 1944 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5867_6
timestamp 1731220618
transform 1 0 1880 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5866_6
timestamp 1731220618
transform 1 0 1816 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5865_6
timestamp 1731220618
transform 1 0 1752 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5864_6
timestamp 1731220618
transform 1 0 1664 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5863_6
timestamp 1731220618
transform 1 0 1840 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5862_6
timestamp 1731220618
transform 1 0 1920 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5861_6
timestamp 1731220618
transform 1 0 2000 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5860_6
timestamp 1731220618
transform 1 0 1976 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5859_6
timestamp 1731220618
transform 1 0 1920 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5858_6
timestamp 1731220618
transform 1 0 1864 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5857_6
timestamp 1731220618
transform 1 0 1816 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5856_6
timestamp 1731220618
transform 1 0 1760 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5855_6
timestamp 1731220618
transform 1 0 1704 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5854_6
timestamp 1731220618
transform 1 0 1912 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5853_6
timestamp 1731220618
transform 1 0 1832 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5852_6
timestamp 1731220618
transform 1 0 1760 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5851_6
timestamp 1731220618
transform 1 0 1696 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5850_6
timestamp 1731220618
transform 1 0 1632 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5849_6
timestamp 1731220618
transform 1 0 1576 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5848_6
timestamp 1731220618
transform 1 0 1712 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5847_6
timestamp 1731220618
transform 1 0 1608 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5846_6
timestamp 1731220618
transform 1 0 1528 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5845_6
timestamp 1731220618
transform 1 0 1464 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5844_6
timestamp 1731220618
transform 1 0 1960 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5843_6
timestamp 1731220618
transform 1 0 1832 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5842_6
timestamp 1731220618
transform 1 0 1712 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5841_6
timestamp 1731220618
transform 1 0 1632 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5840_6
timestamp 1731220618
transform 1 0 1552 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5839_6
timestamp 1731220618
transform 1 0 1792 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5838_6
timestamp 1731220618
transform 1 0 1872 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5837_6
timestamp 1731220618
transform 1 0 1960 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5836_6
timestamp 1731220618
transform 1 0 1896 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5835_6
timestamp 1731220618
transform 1 0 1960 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5834_6
timestamp 1731220618
transform 1 0 2024 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5833_6
timestamp 1731220618
transform 1 0 2048 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5832_6
timestamp 1731220618
transform 1 0 2000 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5831_6
timestamp 1731220618
transform 1 0 2024 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5830_6
timestamp 1731220618
transform 1 0 2064 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5829_6
timestamp 1731220618
transform 1 0 2064 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5828_6
timestamp 1731220618
transform 1 0 2064 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5827_6
timestamp 1731220618
transform 1 0 2064 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5826_6
timestamp 1731220618
transform 1 0 2064 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5825_6
timestamp 1731220618
transform 1 0 2064 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5824_6
timestamp 1731220618
transform 1 0 2064 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5823_6
timestamp 1731220618
transform 1 0 2064 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5822_6
timestamp 1731220618
transform 1 0 1984 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5821_6
timestamp 1731220618
transform 1 0 2008 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5820_6
timestamp 1731220618
transform 1 0 1936 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5819_6
timestamp 1731220618
transform 1 0 1824 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5818_6
timestamp 1731220618
transform 1 0 1752 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5817_6
timestamp 1731220618
transform 1 0 1672 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5816_6
timestamp 1731220618
transform 1 0 1584 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5815_6
timestamp 1731220618
transform 1 0 1864 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5814_6
timestamp 1731220618
transform 1 0 1792 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5813_6
timestamp 1731220618
transform 1 0 1712 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5812_6
timestamp 1731220618
transform 1 0 1624 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5811_6
timestamp 1731220618
transform 1 0 1984 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5810_6
timestamp 1731220618
transform 1 0 1888 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5809_6
timestamp 1731220618
transform 1 0 1800 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5808_6
timestamp 1731220618
transform 1 0 1712 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5807_6
timestamp 1731220618
transform 1 0 1640 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5806_6
timestamp 1731220618
transform 1 0 1576 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5805_6
timestamp 1731220618
transform 1 0 1896 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5804_6
timestamp 1731220618
transform 1 0 1808 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5803_6
timestamp 1731220618
transform 1 0 1728 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5802_6
timestamp 1731220618
transform 1 0 1656 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5801_6
timestamp 1731220618
transform 1 0 1600 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5800_6
timestamp 1731220618
transform 1 0 1552 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5799_6
timestamp 1731220618
transform 1 0 1512 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5798_6
timestamp 1731220618
transform 1 0 1464 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5797_6
timestamp 1731220618
transform 1 0 1560 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5796_6
timestamp 1731220618
transform 1 0 1728 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5795_6
timestamp 1731220618
transform 1 0 1672 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5794_6
timestamp 1731220618
transform 1 0 1616 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5793_6
timestamp 1731220618
transform 1 0 1600 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5792_6
timestamp 1731220618
transform 1 0 1528 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5791_6
timestamp 1731220618
transform 1 0 1672 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5790_6
timestamp 1731220618
transform 1 0 1824 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5789_6
timestamp 1731220618
transform 1 0 1744 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5788_6
timestamp 1731220618
transform 1 0 1672 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5787_6
timestamp 1731220618
transform 1 0 1592 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5786_6
timestamp 1731220618
transform 1 0 1744 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5785_6
timestamp 1731220618
transform 1 0 1808 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5784_6
timestamp 1731220618
transform 1 0 1752 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5783_6
timestamp 1731220618
transform 1 0 1680 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5782_6
timestamp 1731220618
transform 1 0 1824 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5781_6
timestamp 1731220618
transform 1 0 1888 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5780_6
timestamp 1731220618
transform 1 0 1952 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5779_6
timestamp 1731220618
transform 1 0 2016 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5778_6
timestamp 1731220618
transform 1 0 1976 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5777_6
timestamp 1731220618
transform 1 0 1920 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5776_6
timestamp 1731220618
transform 1 0 1864 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5775_6
timestamp 1731220618
transform 1 0 2024 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5774_6
timestamp 1731220618
transform 1 0 2064 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5773_6
timestamp 1731220618
transform 1 0 2064 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5772_6
timestamp 1731220618
transform 1 0 2064 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5771_6
timestamp 1731220618
transform 1 0 2064 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5770_6
timestamp 1731220618
transform 1 0 1976 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5769_6
timestamp 1731220618
transform 1 0 2064 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5768_6
timestamp 1731220618
transform 1 0 2064 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5767_6
timestamp 1731220618
transform 1 0 2000 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5766_6
timestamp 1731220618
transform 1 0 2064 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5765_6
timestamp 1731220618
transform 1 0 2064 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5764_6
timestamp 1731220618
transform 1 0 2016 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5763_6
timestamp 1731220618
transform 1 0 2064 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5762_6
timestamp 1731220618
transform 1 0 2016 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5761_6
timestamp 1731220618
transform 1 0 1944 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5760_6
timestamp 1731220618
transform 1 0 1952 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5759_6
timestamp 1731220618
transform 1 0 2016 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5758_6
timestamp 1731220618
transform 1 0 1952 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5757_6
timestamp 1731220618
transform 1 0 1888 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5756_6
timestamp 1731220618
transform 1 0 1816 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5755_6
timestamp 1731220618
transform 1 0 1736 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5754_6
timestamp 1731220618
transform 1 0 1752 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5753_6
timestamp 1731220618
transform 1 0 1824 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5752_6
timestamp 1731220618
transform 1 0 1888 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5751_6
timestamp 1731220618
transform 1 0 1880 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5750_6
timestamp 1731220618
transform 1 0 1816 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5749_6
timestamp 1731220618
transform 1 0 1744 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5748_6
timestamp 1731220618
transform 1 0 1728 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5747_6
timestamp 1731220618
transform 1 0 1872 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5746_6
timestamp 1731220618
transform 1 0 1800 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5745_6
timestamp 1731220618
transform 1 0 1800 0 1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5744_6
timestamp 1731220618
transform 1 0 1760 0 1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5743_6
timestamp 1731220618
transform 1 0 1720 0 1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5742_6
timestamp 1731220618
transform 1 0 1680 0 1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5741_6
timestamp 1731220618
transform 1 0 1656 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5740_6
timestamp 1731220618
transform 1 0 1584 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5739_6
timestamp 1731220618
transform 1 0 1672 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5738_6
timestamp 1731220618
transform 1 0 1592 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5737_6
timestamp 1731220618
transform 1 0 1584 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5736_6
timestamp 1731220618
transform 1 0 1672 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5735_6
timestamp 1731220618
transform 1 0 1648 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5734_6
timestamp 1731220618
transform 1 0 1624 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5733_6
timestamp 1731220618
transform 1 0 1696 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5732_6
timestamp 1731220618
transform 1 0 1768 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5731_6
timestamp 1731220618
transform 1 0 1840 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5730_6
timestamp 1731220618
transform 1 0 1920 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5729_6
timestamp 1731220618
transform 1 0 1968 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5728_6
timestamp 1731220618
transform 1 0 1856 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5727_6
timestamp 1731220618
transform 1 0 1744 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5726_6
timestamp 1731220618
transform 1 0 1648 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5725_6
timestamp 1731220618
transform 1 0 1568 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5724_6
timestamp 1731220618
transform 1 0 1864 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5723_6
timestamp 1731220618
transform 1 0 1760 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5722_6
timestamp 1731220618
transform 1 0 1664 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5721_6
timestamp 1731220618
transform 1 0 1576 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5720_6
timestamp 1731220618
transform 1 0 1496 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5719_6
timestamp 1731220618
transform 1 0 1424 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5718_6
timestamp 1731220618
transform 1 0 1976 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5717_6
timestamp 1731220618
transform 1 0 1864 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5716_6
timestamp 1731220618
transform 1 0 1760 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5715_6
timestamp 1731220618
transform 1 0 1672 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5714_6
timestamp 1731220618
transform 1 0 1600 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5713_6
timestamp 1731220618
transform 1 0 1544 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5712_6
timestamp 1731220618
transform 1 0 1504 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5711_6
timestamp 1731220618
transform 1 0 1464 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5710_6
timestamp 1731220618
transform 1 0 1424 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5709_6
timestamp 1731220618
transform 1 0 1384 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5708_6
timestamp 1731220618
transform 1 0 1344 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5707_6
timestamp 1731220618
transform 1 0 1304 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5706_6
timestamp 1731220618
transform 1 0 1608 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5705_6
timestamp 1731220618
transform 1 0 1528 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5704_6
timestamp 1731220618
transform 1 0 1448 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5703_6
timestamp 1731220618
transform 1 0 1376 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5702_6
timestamp 1731220618
transform 1 0 1312 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5701_6
timestamp 1731220618
transform 1 0 1256 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5700_6
timestamp 1731220618
transform 1 0 1504 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5699_6
timestamp 1731220618
transform 1 0 1416 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5698_6
timestamp 1731220618
transform 1 0 1328 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5697_6
timestamp 1731220618
transform 1 0 1240 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5696_6
timestamp 1731220618
transform 1 0 1160 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5695_6
timestamp 1731220618
transform 1 0 1312 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5694_6
timestamp 1731220618
transform 1 0 1240 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5693_6
timestamp 1731220618
transform 1 0 1192 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5692_6
timestamp 1731220618
transform 1 0 1152 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5691_6
timestamp 1731220618
transform 1 0 1456 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5690_6
timestamp 1731220618
transform 1 0 1384 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5689_6
timestamp 1731220618
transform 1 0 1320 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5688_6
timestamp 1731220618
transform 1 0 1272 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5687_6
timestamp 1731220618
transform 1 0 1232 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5686_6
timestamp 1731220618
transform 1 0 1368 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5685_6
timestamp 1731220618
transform 1 0 1416 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5684_6
timestamp 1731220618
transform 1 0 1512 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5683_6
timestamp 1731220618
transform 1 0 1472 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5682_6
timestamp 1731220618
transform 1 0 1432 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5681_6
timestamp 1731220618
transform 1 0 1392 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5680_6
timestamp 1731220618
transform 1 0 1352 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5679_6
timestamp 1731220618
transform 1 0 1312 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5678_6
timestamp 1731220618
transform 1 0 1512 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5677_6
timestamp 1731220618
transform 1 0 1448 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5676_6
timestamp 1731220618
transform 1 0 1384 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5675_6
timestamp 1731220618
transform 1 0 1328 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5674_6
timestamp 1731220618
transform 1 0 1272 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5673_6
timestamp 1731220618
transform 1 0 1224 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5672_6
timestamp 1731220618
transform 1 0 1536 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5671_6
timestamp 1731220618
transform 1 0 1440 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5670_6
timestamp 1731220618
transform 1 0 1344 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5669_6
timestamp 1731220618
transform 1 0 1256 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5668_6
timestamp 1731220618
transform 1 0 1192 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5667_6
timestamp 1731220618
transform 1 0 1152 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5666_6
timestamp 1731220618
transform 1 0 1480 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5665_6
timestamp 1731220618
transform 1 0 1368 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5664_6
timestamp 1731220618
transform 1 0 1248 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5663_6
timestamp 1731220618
transform 1 0 1152 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5662_6
timestamp 1731220618
transform 1 0 1040 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5661_6
timestamp 1731220618
transform 1 0 1040 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5660_6
timestamp 1731220618
transform 1 0 1152 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5659_6
timestamp 1731220618
transform 1 0 1192 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5658_6
timestamp 1731220618
transform 1 0 1240 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5657_6
timestamp 1731220618
transform 1 0 1472 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5656_6
timestamp 1731220618
transform 1 0 1392 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5655_6
timestamp 1731220618
transform 1 0 1312 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5654_6
timestamp 1731220618
transform 1 0 1232 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5653_6
timestamp 1731220618
transform 1 0 1192 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5652_6
timestamp 1731220618
transform 1 0 1152 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5651_6
timestamp 1731220618
transform 1 0 1272 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5650_6
timestamp 1731220618
transform 1 0 1320 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5649_6
timestamp 1731220618
transform 1 0 1416 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5648_6
timestamp 1731220618
transform 1 0 1368 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5647_6
timestamp 1731220618
transform 1 0 1360 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5646_6
timestamp 1731220618
transform 1 0 1320 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5645_6
timestamp 1731220618
transform 1 0 1280 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5644_6
timestamp 1731220618
transform 1 0 1408 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5643_6
timestamp 1731220618
transform 1 0 1520 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5642_6
timestamp 1731220618
transform 1 0 1464 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5641_6
timestamp 1731220618
transform 1 0 1464 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5640_6
timestamp 1731220618
transform 1 0 1416 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5639_6
timestamp 1731220618
transform 1 0 1376 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5638_6
timestamp 1731220618
transform 1 0 1520 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5637_6
timestamp 1731220618
transform 1 0 1648 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5636_6
timestamp 1731220618
transform 1 0 1584 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5635_6
timestamp 1731220618
transform 1 0 1568 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5634_6
timestamp 1731220618
transform 1 0 1464 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5633_6
timestamp 1731220618
transform 1 0 1456 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5632_6
timestamp 1731220618
transform 1 0 1536 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5631_6
timestamp 1731220618
transform 1 0 1504 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5630_6
timestamp 1731220618
transform 1 0 1432 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5629_6
timestamp 1731220618
transform 1 0 1416 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5628_6
timestamp 1731220618
transform 1 0 1472 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5627_6
timestamp 1731220618
transform 1 0 1464 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5626_6
timestamp 1731220618
transform 1 0 1392 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5625_6
timestamp 1731220618
transform 1 0 1320 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5624_6
timestamp 1731220618
transform 1 0 1256 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5623_6
timestamp 1731220618
transform 1 0 1192 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5622_6
timestamp 1731220618
transform 1 0 1280 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5621_6
timestamp 1731220618
transform 1 0 1320 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5620_6
timestamp 1731220618
transform 1 0 1368 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5619_6
timestamp 1731220618
transform 1 0 1368 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5618_6
timestamp 1731220618
transform 1 0 1296 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5617_6
timestamp 1731220618
transform 1 0 1232 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5616_6
timestamp 1731220618
transform 1 0 1376 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5615_6
timestamp 1731220618
transform 1 0 1296 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5614_6
timestamp 1731220618
transform 1 0 1224 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5613_6
timestamp 1731220618
transform 1 0 1152 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5612_6
timestamp 1731220618
transform 1 0 1352 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5611_6
timestamp 1731220618
transform 1 0 1240 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5610_6
timestamp 1731220618
transform 1 0 1152 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5609_6
timestamp 1731220618
transform 1 0 1040 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5608_6
timestamp 1731220618
transform 1 0 1000 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5607_6
timestamp 1731220618
transform 1 0 944 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5606_6
timestamp 1731220618
transform 1 0 888 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5605_6
timestamp 1731220618
transform 1 0 896 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5604_6
timestamp 1731220618
transform 1 0 832 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5603_6
timestamp 1731220618
transform 1 0 768 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5602_6
timestamp 1731220618
transform 1 0 696 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5601_6
timestamp 1731220618
transform 1 0 920 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5600_6
timestamp 1731220618
transform 1 0 856 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5599_6
timestamp 1731220618
transform 1 0 792 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5598_6
timestamp 1731220618
transform 1 0 728 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5597_6
timestamp 1731220618
transform 1 0 664 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5596_6
timestamp 1731220618
transform 1 0 592 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5595_6
timestamp 1731220618
transform 1 0 888 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5594_6
timestamp 1731220618
transform 1 0 808 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5593_6
timestamp 1731220618
transform 1 0 736 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5592_6
timestamp 1731220618
transform 1 0 664 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5591_6
timestamp 1731220618
transform 1 0 592 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5590_6
timestamp 1731220618
transform 1 0 520 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5589_6
timestamp 1731220618
transform 1 0 816 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5588_6
timestamp 1731220618
transform 1 0 704 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5587_6
timestamp 1731220618
transform 1 0 608 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5586_6
timestamp 1731220618
transform 1 0 528 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5585_6
timestamp 1731220618
transform 1 0 648 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5584_6
timestamp 1731220618
transform 1 0 576 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5583_6
timestamp 1731220618
transform 1 0 576 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5582_6
timestamp 1731220618
transform 1 0 640 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5581_6
timestamp 1731220618
transform 1 0 624 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5580_6
timestamp 1731220618
transform 1 0 616 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5579_6
timestamp 1731220618
transform 1 0 696 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5578_6
timestamp 1731220618
transform 1 0 656 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5577_6
timestamp 1731220618
transform 1 0 600 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5576_6
timestamp 1731220618
transform 1 0 544 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5575_6
timestamp 1731220618
transform 1 0 512 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5574_6
timestamp 1731220618
transform 1 0 456 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5573_6
timestamp 1731220618
transform 1 0 376 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5572_6
timestamp 1731220618
transform 1 0 464 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5571_6
timestamp 1731220618
transform 1 0 544 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5570_6
timestamp 1731220618
transform 1 0 504 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5569_6
timestamp 1731220618
transform 1 0 432 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5568_6
timestamp 1731220618
transform 1 0 352 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5567_6
timestamp 1731220618
transform 1 0 320 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5566_6
timestamp 1731220618
transform 1 0 368 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5565_6
timestamp 1731220618
transform 1 0 408 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5564_6
timestamp 1731220618
transform 1 0 496 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5563_6
timestamp 1731220618
transform 1 0 456 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5562_6
timestamp 1731220618
transform 1 0 416 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5561_6
timestamp 1731220618
transform 1 0 376 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5560_6
timestamp 1731220618
transform 1 0 336 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5559_6
timestamp 1731220618
transform 1 0 296 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5558_6
timestamp 1731220618
transform 1 0 256 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5557_6
timestamp 1731220618
transform 1 0 216 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5556_6
timestamp 1731220618
transform 1 0 176 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5555_6
timestamp 1731220618
transform 1 0 136 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5554_6
timestamp 1731220618
transform 1 0 272 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5553_6
timestamp 1731220618
transform 1 0 224 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5552_6
timestamp 1731220618
transform 1 0 176 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5551_6
timestamp 1731220618
transform 1 0 128 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5550_6
timestamp 1731220618
transform 1 0 128 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5549_6
timestamp 1731220618
transform 1 0 192 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5548_6
timestamp 1731220618
transform 1 0 272 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5547_6
timestamp 1731220618
transform 1 0 288 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5546_6
timestamp 1731220618
transform 1 0 200 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5545_6
timestamp 1731220618
transform 1 0 128 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5544_6
timestamp 1731220618
transform 1 0 128 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5543_6
timestamp 1731220618
transform 1 0 168 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5542_6
timestamp 1731220618
transform 1 0 328 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5541_6
timestamp 1731220618
transform 1 0 264 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5540_6
timestamp 1731220618
transform 1 0 208 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5539_6
timestamp 1731220618
transform 1 0 144 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5538_6
timestamp 1731220618
transform 1 0 160 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5537_6
timestamp 1731220618
transform 1 0 160 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5536_6
timestamp 1731220618
transform 1 0 216 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5535_6
timestamp 1731220618
transform 1 0 200 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5534_6
timestamp 1731220618
transform 1 0 248 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5533_6
timestamp 1731220618
transform 1 0 280 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5532_6
timestamp 1731220618
transform 1 0 240 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5531_6
timestamp 1731220618
transform 1 0 304 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5530_6
timestamp 1731220618
transform 1 0 288 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5529_6
timestamp 1731220618
transform 1 0 200 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5528_6
timestamp 1731220618
transform 1 0 272 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5527_6
timestamp 1731220618
transform 1 0 328 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5526_6
timestamp 1731220618
transform 1 0 384 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5525_6
timestamp 1731220618
transform 1 0 392 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5524_6
timestamp 1731220618
transform 1 0 336 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5523_6
timestamp 1731220618
transform 1 0 320 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5522_6
timestamp 1731220618
transform 1 0 392 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5521_6
timestamp 1731220618
transform 1 0 456 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5520_6
timestamp 1731220618
transform 1 0 440 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5519_6
timestamp 1731220618
transform 1 0 520 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5518_6
timestamp 1731220618
transform 1 0 472 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5517_6
timestamp 1731220618
transform 1 0 552 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5516_6
timestamp 1731220618
transform 1 0 624 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5515_6
timestamp 1731220618
transform 1 0 640 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5514_6
timestamp 1731220618
transform 1 0 568 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5513_6
timestamp 1731220618
transform 1 0 496 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5512_6
timestamp 1731220618
transform 1 0 504 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5511_6
timestamp 1731220618
transform 1 0 584 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5510_6
timestamp 1731220618
transform 1 0 672 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5509_6
timestamp 1731220618
transform 1 0 768 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5508_6
timestamp 1731220618
transform 1 0 784 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5507_6
timestamp 1731220618
transform 1 0 704 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5506_6
timestamp 1731220618
transform 1 0 624 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5505_6
timestamp 1731220618
transform 1 0 544 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5504_6
timestamp 1731220618
transform 1 0 600 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5503_6
timestamp 1731220618
transform 1 0 664 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5502_6
timestamp 1731220618
transform 1 0 728 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5501_6
timestamp 1731220618
transform 1 0 792 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5500_6
timestamp 1731220618
transform 1 0 736 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5499_6
timestamp 1731220618
transform 1 0 664 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5498_6
timestamp 1731220618
transform 1 0 816 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5497_6
timestamp 1731220618
transform 1 0 856 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5496_6
timestamp 1731220618
transform 1 0 792 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5495_6
timestamp 1731220618
transform 1 0 728 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5494_6
timestamp 1731220618
transform 1 0 664 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5493_6
timestamp 1731220618
transform 1 0 688 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5492_6
timestamp 1731220618
transform 1 0 752 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5491_6
timestamp 1731220618
transform 1 0 816 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5490_6
timestamp 1731220618
transform 1 0 800 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5489_6
timestamp 1731220618
transform 1 0 744 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5488_6
timestamp 1731220618
transform 1 0 688 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5487_6
timestamp 1731220618
transform 1 0 640 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5486_6
timestamp 1731220618
transform 1 0 768 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5485_6
timestamp 1731220618
transform 1 0 728 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5484_6
timestamp 1731220618
transform 1 0 688 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5483_6
timestamp 1731220618
transform 1 0 648 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5482_6
timestamp 1731220618
transform 1 0 608 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5481_6
timestamp 1731220618
transform 1 0 568 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5480_6
timestamp 1731220618
transform 1 0 512 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5479_6
timestamp 1731220618
transform 1 0 552 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5478_6
timestamp 1731220618
transform 1 0 592 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5477_6
timestamp 1731220618
transform 1 0 624 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5476_6
timestamp 1731220618
transform 1 0 568 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5475_6
timestamp 1731220618
transform 1 0 512 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5474_6
timestamp 1731220618
transform 1 0 464 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5473_6
timestamp 1731220618
transform 1 0 424 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5472_6
timestamp 1731220618
transform 1 0 600 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5471_6
timestamp 1731220618
transform 1 0 536 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5470_6
timestamp 1731220618
transform 1 0 472 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5469_6
timestamp 1731220618
transform 1 0 416 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5468_6
timestamp 1731220618
transform 1 0 368 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5467_6
timestamp 1731220618
transform 1 0 592 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5466_6
timestamp 1731220618
transform 1 0 520 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5465_6
timestamp 1731220618
transform 1 0 448 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5464_6
timestamp 1731220618
transform 1 0 384 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5463_6
timestamp 1731220618
transform 1 0 328 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5462_6
timestamp 1731220618
transform 1 0 536 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5461_6
timestamp 1731220618
transform 1 0 472 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5460_6
timestamp 1731220618
transform 1 0 408 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5459_6
timestamp 1731220618
transform 1 0 352 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5458_6
timestamp 1731220618
transform 1 0 304 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5457_6
timestamp 1731220618
transform 1 0 256 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5456_6
timestamp 1731220618
transform 1 0 472 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5455_6
timestamp 1731220618
transform 1 0 400 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5454_6
timestamp 1731220618
transform 1 0 336 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5453_6
timestamp 1731220618
transform 1 0 272 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5452_6
timestamp 1731220618
transform 1 0 216 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5451_6
timestamp 1731220618
transform 1 0 432 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5450_6
timestamp 1731220618
transform 1 0 360 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5449_6
timestamp 1731220618
transform 1 0 296 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5448_6
timestamp 1731220618
transform 1 0 240 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5447_6
timestamp 1731220618
transform 1 0 192 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5446_6
timestamp 1731220618
transform 1 0 152 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5445_6
timestamp 1731220618
transform 1 0 192 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5444_6
timestamp 1731220618
transform 1 0 240 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5443_6
timestamp 1731220618
transform 1 0 296 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5442_6
timestamp 1731220618
transform 1 0 360 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5441_6
timestamp 1731220618
transform 1 0 424 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5440_6
timestamp 1731220618
transform 1 0 400 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5439_6
timestamp 1731220618
transform 1 0 328 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5438_6
timestamp 1731220618
transform 1 0 264 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5437_6
timestamp 1731220618
transform 1 0 216 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5436_6
timestamp 1731220618
transform 1 0 360 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5435_6
timestamp 1731220618
transform 1 0 280 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5434_6
timestamp 1731220618
transform 1 0 208 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5433_6
timestamp 1731220618
transform 1 0 144 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5432_6
timestamp 1731220618
transform 1 0 128 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5431_6
timestamp 1731220618
transform 1 0 176 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5430_6
timestamp 1731220618
transform 1 0 248 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5429_6
timestamp 1731220618
transform 1 0 272 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5428_6
timestamp 1731220618
transform 1 0 208 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5427_6
timestamp 1731220618
transform 1 0 168 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5426_6
timestamp 1731220618
transform 1 0 128 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5425_6
timestamp 1731220618
transform 1 0 128 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5424_6
timestamp 1731220618
transform 1 0 208 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5423_6
timestamp 1731220618
transform 1 0 168 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5422_6
timestamp 1731220618
transform 1 0 128 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5421_6
timestamp 1731220618
transform 1 0 128 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5420_6
timestamp 1731220618
transform 1 0 176 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5419_6
timestamp 1731220618
transform 1 0 208 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5418_6
timestamp 1731220618
transform 1 0 152 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5417_6
timestamp 1731220618
transform 1 0 152 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5416_6
timestamp 1731220618
transform 1 0 304 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5415_6
timestamp 1731220618
transform 1 0 352 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5414_6
timestamp 1731220618
transform 1 0 280 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5413_6
timestamp 1731220618
transform 1 0 224 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5412_6
timestamp 1731220618
transform 1 0 296 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5411_6
timestamp 1731220618
transform 1 0 272 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5410_6
timestamp 1731220618
transform 1 0 208 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5409_6
timestamp 1731220618
transform 1 0 392 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5408_6
timestamp 1731220618
transform 1 0 344 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5407_6
timestamp 1731220618
transform 1 0 416 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5406_6
timestamp 1731220618
transform 1 0 480 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5405_6
timestamp 1731220618
transform 1 0 528 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5404_6
timestamp 1731220618
transform 1 0 448 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5403_6
timestamp 1731220618
transform 1 0 368 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5402_6
timestamp 1731220618
transform 1 0 424 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5401_6
timestamp 1731220618
transform 1 0 504 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5400_6
timestamp 1731220618
transform 1 0 584 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5399_6
timestamp 1731220618
transform 1 0 536 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5398_6
timestamp 1731220618
transform 1 0 456 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5397_6
timestamp 1731220618
transform 1 0 376 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5396_6
timestamp 1731220618
transform 1 0 360 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5395_6
timestamp 1731220618
transform 1 0 448 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5394_6
timestamp 1731220618
transform 1 0 536 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5393_6
timestamp 1731220618
transform 1 0 512 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5392_6
timestamp 1731220618
transform 1 0 448 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5391_6
timestamp 1731220618
transform 1 0 376 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5390_6
timestamp 1731220618
transform 1 0 368 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5389_6
timestamp 1731220618
transform 1 0 440 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5388_6
timestamp 1731220618
transform 1 0 512 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5387_6
timestamp 1731220618
transform 1 0 576 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5386_6
timestamp 1731220618
transform 1 0 512 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5385_6
timestamp 1731220618
transform 1 0 448 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5384_6
timestamp 1731220618
transform 1 0 456 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5383_6
timestamp 1731220618
transform 1 0 936 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5382_6
timestamp 1731220618
transform 1 0 808 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5381_6
timestamp 1731220618
transform 1 0 728 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5380_6
timestamp 1731220618
transform 1 0 680 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5379_6
timestamp 1731220618
transform 1 0 632 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5378_6
timestamp 1731220618
transform 1 0 736 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5377_6
timestamp 1731220618
transform 1 0 848 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5376_6
timestamp 1731220618
transform 1 0 792 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5375_6
timestamp 1731220618
transform 1 0 760 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5374_6
timestamp 1731220618
transform 1 0 704 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5373_6
timestamp 1731220618
transform 1 0 936 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5372_6
timestamp 1731220618
transform 1 0 872 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5371_6
timestamp 1731220618
transform 1 0 816 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5370_6
timestamp 1731220618
transform 1 0 792 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5369_6
timestamp 1731220618
transform 1 0 712 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5368_6
timestamp 1731220618
transform 1 0 1024 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5367_6
timestamp 1731220618
transform 1 0 944 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5366_6
timestamp 1731220618
transform 1 0 864 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5365_6
timestamp 1731220618
transform 1 0 848 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5364_6
timestamp 1731220618
transform 1 0 776 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5363_6
timestamp 1731220618
transform 1 0 920 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5362_6
timestamp 1731220618
transform 1 0 992 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5361_6
timestamp 1731220618
transform 1 0 1040 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5360_6
timestamp 1731220618
transform 1 0 1040 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5359_6
timestamp 1731220618
transform 1 0 992 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5358_6
timestamp 1731220618
transform 1 0 928 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5357_6
timestamp 1731220618
transform 1 0 864 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5356_6
timestamp 1731220618
transform 1 0 800 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5355_6
timestamp 1731220618
transform 1 0 728 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5354_6
timestamp 1731220618
transform 1 0 896 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5353_6
timestamp 1731220618
transform 1 0 848 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5352_6
timestamp 1731220618
transform 1 0 792 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5351_6
timestamp 1731220618
transform 1 0 736 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5350_6
timestamp 1731220618
transform 1 0 672 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5349_6
timestamp 1731220618
transform 1 0 848 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5348_6
timestamp 1731220618
transform 1 0 784 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5347_6
timestamp 1731220618
transform 1 0 720 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5346_6
timestamp 1731220618
transform 1 0 664 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5345_6
timestamp 1731220618
transform 1 0 608 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5344_6
timestamp 1731220618
transform 1 0 568 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5343_6
timestamp 1731220618
transform 1 0 744 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5342_6
timestamp 1731220618
transform 1 0 680 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5341_6
timestamp 1731220618
transform 1 0 624 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5340_6
timestamp 1731220618
transform 1 0 616 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5339_6
timestamp 1731220618
transform 1 0 680 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5338_6
timestamp 1731220618
transform 1 0 744 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5337_6
timestamp 1731220618
transform 1 0 800 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5336_6
timestamp 1731220618
transform 1 0 864 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5335_6
timestamp 1731220618
transform 1 0 928 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5334_6
timestamp 1731220618
transform 1 0 872 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5333_6
timestamp 1731220618
transform 1 0 808 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5332_6
timestamp 1731220618
transform 1 0 752 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5331_6
timestamp 1731220618
transform 1 0 696 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5330_6
timestamp 1731220618
transform 1 0 640 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5329_6
timestamp 1731220618
transform 1 0 576 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5328_6
timestamp 1731220618
transform 1 0 736 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5327_6
timestamp 1731220618
transform 1 0 688 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5326_6
timestamp 1731220618
transform 1 0 640 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5325_6
timestamp 1731220618
transform 1 0 592 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5324_6
timestamp 1731220618
transform 1 0 544 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5323_6
timestamp 1731220618
transform 1 0 496 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5322_6
timestamp 1731220618
transform 1 0 448 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5321_6
timestamp 1731220618
transform 1 0 536 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5320_6
timestamp 1731220618
transform 1 0 576 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5319_6
timestamp 1731220618
transform 1 0 616 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5318_6
timestamp 1731220618
transform 1 0 656 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5317_6
timestamp 1731220618
transform 1 0 696 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5316_6
timestamp 1731220618
transform 1 0 736 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5315_6
timestamp 1731220618
transform 1 0 776 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5314_6
timestamp 1731220618
transform 1 0 824 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5313_6
timestamp 1731220618
transform 1 0 872 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5312_6
timestamp 1731220618
transform 1 0 920 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5311_6
timestamp 1731220618
transform 1 0 960 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5310_6
timestamp 1731220618
transform 1 0 1000 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5309_6
timestamp 1731220618
transform 1 0 1040 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5308_6
timestamp 1731220618
transform 1 0 1152 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5307_6
timestamp 1731220618
transform 1 0 1152 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5306_6
timestamp 1731220618
transform 1 0 1192 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5305_6
timestamp 1731220618
transform 1 0 1256 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5304_6
timestamp 1731220618
transform 1 0 1264 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5303_6
timestamp 1731220618
transform 1 0 1200 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5302_6
timestamp 1731220618
transform 1 0 1152 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5301_6
timestamp 1731220618
transform 1 0 1160 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5300_6
timestamp 1731220618
transform 1 0 1200 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5299_6
timestamp 1731220618
transform 1 0 1240 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5298_6
timestamp 1731220618
transform 1 0 1288 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5297_6
timestamp 1731220618
transform 1 0 1384 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5296_6
timestamp 1731220618
transform 1 0 1336 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5295_6
timestamp 1731220618
transform 1 0 1320 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5294_6
timestamp 1731220618
transform 1 0 1384 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5293_6
timestamp 1731220618
transform 1 0 1392 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5292_6
timestamp 1731220618
transform 1 0 1320 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5291_6
timestamp 1731220618
transform 1 0 1264 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5290_6
timestamp 1731220618
transform 1 0 1200 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5289_6
timestamp 1731220618
transform 1 0 1328 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5288_6
timestamp 1731220618
transform 1 0 1392 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5287_6
timestamp 1731220618
transform 1 0 1448 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5286_6
timestamp 1731220618
transform 1 0 1504 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5285_6
timestamp 1731220618
transform 1 0 1536 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5284_6
timestamp 1731220618
transform 1 0 1464 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5283_6
timestamp 1731220618
transform 1 0 1448 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5282_6
timestamp 1731220618
transform 1 0 1520 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5281_6
timestamp 1731220618
transform 1 0 1488 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5280_6
timestamp 1731220618
transform 1 0 1432 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5279_6
timestamp 1731220618
transform 1 0 1616 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5278_6
timestamp 1731220618
transform 1 0 1744 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5277_6
timestamp 1731220618
transform 1 0 1672 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5276_6
timestamp 1731220618
transform 1 0 1608 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5275_6
timestamp 1731220618
transform 1 0 1544 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5274_6
timestamp 1731220618
transform 1 0 1552 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5273_6
timestamp 1731220618
transform 1 0 1496 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5272_6
timestamp 1731220618
transform 1 0 1456 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5271_6
timestamp 1731220618
transform 1 0 1416 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5270_6
timestamp 1731220618
transform 1 0 1376 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5269_6
timestamp 1731220618
transform 1 0 1336 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5268_6
timestamp 1731220618
transform 1 0 1296 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5267_6
timestamp 1731220618
transform 1 0 1496 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5266_6
timestamp 1731220618
transform 1 0 1408 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5265_6
timestamp 1731220618
transform 1 0 1328 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5264_6
timestamp 1731220618
transform 1 0 1248 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5263_6
timestamp 1731220618
transform 1 0 1192 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5262_6
timestamp 1731220618
transform 1 0 1152 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5261_6
timestamp 1731220618
transform 1 0 1152 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5260_6
timestamp 1731220618
transform 1 0 1040 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5259_6
timestamp 1731220618
transform 1 0 1000 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5258_6
timestamp 1731220618
transform 1 0 952 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5257_6
timestamp 1731220618
transform 1 0 1256 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5256_6
timestamp 1731220618
transform 1 0 1376 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5255_6
timestamp 1731220618
transform 1 0 1280 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5254_6
timestamp 1731220618
transform 1 0 1232 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5253_6
timestamp 1731220618
transform 1 0 1184 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5252_6
timestamp 1731220618
transform 1 0 1336 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5251_6
timestamp 1731220618
transform 1 0 1400 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5250_6
timestamp 1731220618
transform 1 0 1472 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5249_6
timestamp 1731220618
transform 1 0 1512 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5248_6
timestamp 1731220618
transform 1 0 1456 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5247_6
timestamp 1731220618
transform 1 0 1408 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5246_6
timestamp 1731220618
transform 1 0 1368 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5245_6
timestamp 1731220618
transform 1 0 1328 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5244_6
timestamp 1731220618
transform 1 0 1416 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5243_6
timestamp 1731220618
transform 1 0 1360 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5242_6
timestamp 1731220618
transform 1 0 1312 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5241_6
timestamp 1731220618
transform 1 0 1272 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5240_6
timestamp 1731220618
transform 1 0 1232 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5239_6
timestamp 1731220618
transform 1 0 1280 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5238_6
timestamp 1731220618
transform 1 0 1328 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5237_6
timestamp 1731220618
transform 1 0 1432 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5236_6
timestamp 1731220618
transform 1 0 1352 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5235_6
timestamp 1731220618
transform 1 0 1280 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5234_6
timestamp 1731220618
transform 1 0 1232 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5233_6
timestamp 1731220618
transform 1 0 1192 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5232_6
timestamp 1731220618
transform 1 0 1152 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5231_6
timestamp 1731220618
transform 1 0 1336 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5230_6
timestamp 1731220618
transform 1 0 1232 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5229_6
timestamp 1731220618
transform 1 0 1152 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5228_6
timestamp 1731220618
transform 1 0 1040 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5227_6
timestamp 1731220618
transform 1 0 976 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5226_6
timestamp 1731220618
transform 1 0 888 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5225_6
timestamp 1731220618
transform 1 0 1040 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5224_6
timestamp 1731220618
transform 1 0 1152 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5223_6
timestamp 1731220618
transform 1 0 1040 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5222_6
timestamp 1731220618
transform 1 0 976 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5221_6
timestamp 1731220618
transform 1 0 984 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5220_6
timestamp 1731220618
transform 1 0 1040 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5219_6
timestamp 1731220618
transform 1 0 1032 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5218_6
timestamp 1731220618
transform 1 0 960 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5217_6
timestamp 1731220618
transform 1 0 832 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5216_6
timestamp 1731220618
transform 1 0 776 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5215_6
timestamp 1731220618
transform 1 0 712 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5214_6
timestamp 1731220618
transform 1 0 872 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5213_6
timestamp 1731220618
transform 1 0 984 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5212_6
timestamp 1731220618
transform 1 0 952 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5211_6
timestamp 1731220618
transform 1 0 864 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5210_6
timestamp 1731220618
transform 1 0 856 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5209_6
timestamp 1731220618
transform 1 0 920 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5208_6
timestamp 1731220618
transform 1 0 896 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5207_6
timestamp 1731220618
transform 1 0 976 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5206_6
timestamp 1731220618
transform 1 0 920 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5205_6
timestamp 1731220618
transform 1 0 992 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5204_6
timestamp 1731220618
transform 1 0 960 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5203_6
timestamp 1731220618
transform 1 0 888 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5202_6
timestamp 1731220618
transform 1 0 864 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5201_6
timestamp 1731220618
transform 1 0 928 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5200_6
timestamp 1731220618
transform 1 0 880 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5199_6
timestamp 1731220618
transform 1 0 824 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5198_6
timestamp 1731220618
transform 1 0 848 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5197_6
timestamp 1731220618
transform 1 0 784 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5196_6
timestamp 1731220618
transform 1 0 720 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5195_6
timestamp 1731220618
transform 1 0 656 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5194_6
timestamp 1731220618
transform 1 0 600 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5193_6
timestamp 1731220618
transform 1 0 536 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5192_6
timestamp 1731220618
transform 1 0 600 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5191_6
timestamp 1731220618
transform 1 0 544 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5190_6
timestamp 1731220618
transform 1 0 496 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5189_6
timestamp 1731220618
transform 1 0 448 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5188_6
timestamp 1731220618
transform 1 0 712 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5187_6
timestamp 1731220618
transform 1 0 656 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5186_6
timestamp 1731220618
transform 1 0 600 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5185_6
timestamp 1731220618
transform 1 0 664 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5184_6
timestamp 1731220618
transform 1 0 728 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5183_6
timestamp 1731220618
transform 1 0 872 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5182_6
timestamp 1731220618
transform 1 0 800 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5181_6
timestamp 1731220618
transform 1 0 744 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5180_6
timestamp 1731220618
transform 1 0 664 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5179_6
timestamp 1731220618
transform 1 0 816 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5178_6
timestamp 1731220618
transform 1 0 880 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5177_6
timestamp 1731220618
transform 1 0 1024 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5176_6
timestamp 1731220618
transform 1 0 952 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5175_6
timestamp 1731220618
transform 1 0 904 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5174_6
timestamp 1731220618
transform 1 0 832 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5173_6
timestamp 1731220618
transform 1 0 984 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5172_6
timestamp 1731220618
transform 1 0 1040 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5171_6
timestamp 1731220618
transform 1 0 1152 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5170_6
timestamp 1731220618
transform 1 0 1192 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5169_6
timestamp 1731220618
transform 1 0 1232 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5168_6
timestamp 1731220618
transform 1 0 1360 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5167_6
timestamp 1731220618
transform 1 0 1296 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5166_6
timestamp 1731220618
transform 1 0 1264 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5165_6
timestamp 1731220618
transform 1 0 1224 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5164_6
timestamp 1731220618
transform 1 0 1312 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5163_6
timestamp 1731220618
transform 1 0 1368 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5162_6
timestamp 1731220618
transform 1 0 1496 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5161_6
timestamp 1731220618
transform 1 0 1432 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5160_6
timestamp 1731220618
transform 1 0 1416 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5159_6
timestamp 1731220618
transform 1 0 1352 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5158_6
timestamp 1731220618
transform 1 0 1480 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5157_6
timestamp 1731220618
transform 1 0 1552 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5156_6
timestamp 1731220618
transform 1 0 1552 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5155_6
timestamp 1731220618
transform 1 0 1448 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5154_6
timestamp 1731220618
transform 1 0 1344 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5153_6
timestamp 1731220618
transform 1 0 1392 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5152_6
timestamp 1731220618
transform 1 0 1488 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5151_6
timestamp 1731220618
transform 1 0 1432 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5150_6
timestamp 1731220618
transform 1 0 1360 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5149_6
timestamp 1731220618
transform 1 0 1512 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5148_6
timestamp 1731220618
transform 1 0 1520 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5147_6
timestamp 1731220618
transform 1 0 1448 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5146_6
timestamp 1731220618
transform 1 0 1384 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5145_6
timestamp 1731220618
transform 1 0 1328 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5144_6
timestamp 1731220618
transform 1 0 1272 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5143_6
timestamp 1731220618
transform 1 0 1232 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5142_6
timestamp 1731220618
transform 1 0 1192 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5141_6
timestamp 1731220618
transform 1 0 1152 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5140_6
timestamp 1731220618
transform 1 0 1288 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5139_6
timestamp 1731220618
transform 1 0 1232 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5138_6
timestamp 1731220618
transform 1 0 1192 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5137_6
timestamp 1731220618
transform 1 0 1152 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5136_6
timestamp 1731220618
transform 1 0 1152 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5135_6
timestamp 1731220618
transform 1 0 1208 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5134_6
timestamp 1731220618
transform 1 0 1296 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5133_6
timestamp 1731220618
transform 1 0 1232 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5132_6
timestamp 1731220618
transform 1 0 1152 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5131_6
timestamp 1731220618
transform 1 0 1040 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5130_6
timestamp 1731220618
transform 1 0 1000 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5129_6
timestamp 1731220618
transform 1 0 952 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5128_6
timestamp 1731220618
transform 1 0 904 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5127_6
timestamp 1731220618
transform 1 0 856 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5126_6
timestamp 1731220618
transform 1 0 808 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5125_6
timestamp 1731220618
transform 1 0 856 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5124_6
timestamp 1731220618
transform 1 0 944 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5123_6
timestamp 1731220618
transform 1 0 1032 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5122_6
timestamp 1731220618
transform 1 0 960 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5121_6
timestamp 1731220618
transform 1 0 872 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5120_6
timestamp 1731220618
transform 1 0 792 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5119_6
timestamp 1731220618
transform 1 0 896 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5118_6
timestamp 1731220618
transform 1 0 840 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5117_6
timestamp 1731220618
transform 1 0 784 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5116_6
timestamp 1731220618
transform 1 0 728 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5115_6
timestamp 1731220618
transform 1 0 680 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5114_6
timestamp 1731220618
transform 1 0 624 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5113_6
timestamp 1731220618
transform 1 0 568 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5112_6
timestamp 1731220618
transform 1 0 504 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5111_6
timestamp 1731220618
transform 1 0 552 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5110_6
timestamp 1731220618
transform 1 0 632 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5109_6
timestamp 1731220618
transform 1 0 712 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5108_6
timestamp 1731220618
transform 1 0 696 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5107_6
timestamp 1731220618
transform 1 0 776 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5106_6
timestamp 1731220618
transform 1 0 752 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5105_6
timestamp 1731220618
transform 1 0 688 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5104_6
timestamp 1731220618
transform 1 0 616 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5103_6
timestamp 1731220618
transform 1 0 752 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5102_6
timestamp 1731220618
transform 1 0 824 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5101_6
timestamp 1731220618
transform 1 0 984 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5100_6
timestamp 1731220618
transform 1 0 904 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_599_6
timestamp 1731220618
transform 1 0 872 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_598_6
timestamp 1731220618
transform 1 0 784 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_597_6
timestamp 1731220618
transform 1 0 824 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_596_6
timestamp 1731220618
transform 1 0 752 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_595_6
timestamp 1731220618
transform 1 0 688 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_594_6
timestamp 1731220618
transform 1 0 760 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_593_6
timestamp 1731220618
transform 1 0 680 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_592_6
timestamp 1731220618
transform 1 0 600 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_591_6
timestamp 1731220618
transform 1 0 560 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_590_6
timestamp 1731220618
transform 1 0 496 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_589_6
timestamp 1731220618
transform 1 0 624 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_588_6
timestamp 1731220618
transform 1 0 608 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_587_6
timestamp 1731220618
transform 1 0 520 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_586_6
timestamp 1731220618
transform 1 0 696 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_585_6
timestamp 1731220618
transform 1 0 680 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_584_6
timestamp 1731220618
transform 1 0 600 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_583_6
timestamp 1731220618
transform 1 0 520 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_582_6
timestamp 1731220618
transform 1 0 440 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_581_6
timestamp 1731220618
transform 1 0 456 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_580_6
timestamp 1731220618
transform 1 0 536 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_579_6
timestamp 1731220618
transform 1 0 616 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_578_6
timestamp 1731220618
transform 1 0 536 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_577_6
timestamp 1731220618
transform 1 0 464 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_576_6
timestamp 1731220618
transform 1 0 400 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_575_6
timestamp 1731220618
transform 1 0 344 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_574_6
timestamp 1731220618
transform 1 0 368 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_573_6
timestamp 1731220618
transform 1 0 368 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_572_6
timestamp 1731220618
transform 1 0 296 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_571_6
timestamp 1731220618
transform 1 0 224 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_570_6
timestamp 1731220618
transform 1 0 440 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_569_6
timestamp 1731220618
transform 1 0 360 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_568_6
timestamp 1731220618
transform 1 0 288 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_567_6
timestamp 1731220618
transform 1 0 224 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_566_6
timestamp 1731220618
transform 1 0 280 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_565_6
timestamp 1731220618
transform 1 0 424 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_564_6
timestamp 1731220618
transform 1 0 352 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_563_6
timestamp 1731220618
transform 1 0 344 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_562_6
timestamp 1731220618
transform 1 0 256 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_561_6
timestamp 1731220618
transform 1 0 432 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_560_6
timestamp 1731220618
transform 1 0 520 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_559_6
timestamp 1731220618
transform 1 0 488 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_558_6
timestamp 1731220618
transform 1 0 392 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_557_6
timestamp 1731220618
transform 1 0 584 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_556_6
timestamp 1731220618
transform 1 0 528 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_555_6
timestamp 1731220618
transform 1 0 456 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_554_6
timestamp 1731220618
transform 1 0 376 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_553_6
timestamp 1731220618
transform 1 0 296 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_552_6
timestamp 1731220618
transform 1 0 296 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_551_6
timestamp 1731220618
transform 1 0 400 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_550_6
timestamp 1731220618
transform 1 0 352 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_549_6
timestamp 1731220618
transform 1 0 344 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_548_6
timestamp 1731220618
transform 1 0 408 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_547_6
timestamp 1731220618
transform 1 0 472 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_546_6
timestamp 1731220618
transform 1 0 528 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_545_6
timestamp 1731220618
transform 1 0 488 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_544_6
timestamp 1731220618
transform 1 0 448 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_543_6
timestamp 1731220618
transform 1 0 408 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_542_6
timestamp 1731220618
transform 1 0 368 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_541_6
timestamp 1731220618
transform 1 0 328 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_540_6
timestamp 1731220618
transform 1 0 288 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_539_6
timestamp 1731220618
transform 1 0 248 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_538_6
timestamp 1731220618
transform 1 0 208 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_537_6
timestamp 1731220618
transform 1 0 168 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_536_6
timestamp 1731220618
transform 1 0 128 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_535_6
timestamp 1731220618
transform 1 0 136 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_534_6
timestamp 1731220618
transform 1 0 176 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_533_6
timestamp 1731220618
transform 1 0 224 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_532_6
timestamp 1731220618
transform 1 0 280 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_531_6
timestamp 1731220618
transform 1 0 248 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_530_6
timestamp 1731220618
transform 1 0 208 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_529_6
timestamp 1731220618
transform 1 0 168 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_528_6
timestamp 1731220618
transform 1 0 144 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_527_6
timestamp 1731220618
transform 1 0 216 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_526_6
timestamp 1731220618
transform 1 0 288 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_525_6
timestamp 1731220618
transform 1 0 192 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_524_6
timestamp 1731220618
transform 1 0 128 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_523_6
timestamp 1731220618
transform 1 0 176 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_522_6
timestamp 1731220618
transform 1 0 128 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_521_6
timestamp 1731220618
transform 1 0 128 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_520_6
timestamp 1731220618
transform 1 0 216 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_519_6
timestamp 1731220618
transform 1 0 168 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_518_6
timestamp 1731220618
transform 1 0 128 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_517_6
timestamp 1731220618
transform 1 0 168 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_516_6
timestamp 1731220618
transform 1 0 152 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_515_6
timestamp 1731220618
transform 1 0 176 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_514_6
timestamp 1731220618
transform 1 0 272 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_513_6
timestamp 1731220618
transform 1 0 296 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_512_6
timestamp 1731220618
transform 1 0 480 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_511_6
timestamp 1731220618
transform 1 0 416 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_510_6
timestamp 1731220618
transform 1 0 352 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_59_6
timestamp 1731220618
transform 1 0 304 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_58_6
timestamp 1731220618
transform 1 0 264 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_57_6
timestamp 1731220618
transform 1 0 224 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_56_6
timestamp 1731220618
transform 1 0 440 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_55_6
timestamp 1731220618
transform 1 0 376 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_54_6
timestamp 1731220618
transform 1 0 312 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_53_6
timestamp 1731220618
transform 1 0 248 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_52_6
timestamp 1731220618
transform 1 0 208 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_51_6
timestamp 1731220618
transform 1 0 168 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_50_6
timestamp 1731220618
transform 1 0 128 0 -1 2212
box 4 6 36 48
<< end >>
