magic
tech sky130l
timestamp 1731001050
<< m1 >>
rect 352 1035 356 1055
rect 128 767 132 847
rect 768 807 772 895
rect 1008 891 1012 919
rect 400 767 404 787
rect 1008 767 1012 847
rect 856 719 860 763
rect 1008 615 1012 703
rect 560 455 564 491
rect 664 431 668 451
rect 128 323 132 351
rect 968 331 972 411
rect 192 175 196 215
rect 472 195 476 279
<< m2c >>
rect 111 1197 115 1201
rect 1111 1197 1115 1201
rect 111 1179 115 1183
rect 1111 1179 1115 1183
rect 111 1129 115 1133
rect 1111 1129 1115 1133
rect 111 1111 115 1115
rect 1111 1111 1115 1115
rect 111 1069 115 1073
rect 1111 1069 1115 1073
rect 352 1055 356 1059
rect 111 1051 115 1055
rect 1111 1051 1115 1055
rect 352 1031 356 1035
rect 111 993 115 997
rect 1111 993 1115 997
rect 111 975 115 979
rect 1111 975 1115 979
rect 111 933 115 937
rect 1111 933 1115 937
rect 1008 919 1012 923
rect 111 915 115 919
rect 768 895 772 899
rect 111 865 115 869
rect 111 847 115 851
rect 128 847 132 851
rect 111 801 115 805
rect 111 783 115 787
rect 1111 915 1115 919
rect 1008 887 1012 891
rect 1111 865 1115 869
rect 768 803 772 807
rect 1008 847 1012 851
rect 1111 847 1115 851
rect 128 763 132 767
rect 400 787 404 791
rect 1111 801 1115 805
rect 1111 783 1115 787
rect 400 763 404 767
rect 856 763 860 767
rect 1008 763 1012 767
rect 111 721 115 725
rect 1111 721 1115 725
rect 856 715 860 719
rect 111 703 115 707
rect 1008 703 1012 707
rect 1111 703 1115 707
rect 111 649 115 653
rect 111 631 115 635
rect 1111 649 1115 653
rect 1111 631 1115 635
rect 1008 611 1012 615
rect 111 573 115 577
rect 1111 573 1115 577
rect 111 555 115 559
rect 1111 555 1115 559
rect 111 505 115 509
rect 1111 505 1115 509
rect 560 491 564 495
rect 111 487 115 491
rect 1111 487 1115 491
rect 560 451 564 455
rect 664 451 668 455
rect 111 429 115 433
rect 664 427 668 431
rect 1111 429 1115 433
rect 111 411 115 415
rect 968 411 972 415
rect 1111 411 1115 415
rect 111 365 115 369
rect 128 351 132 355
rect 111 347 115 351
rect 1111 365 1115 369
rect 1111 347 1115 351
rect 968 327 972 331
rect 128 319 132 323
rect 111 297 115 301
rect 1111 297 1115 301
rect 111 279 115 283
rect 472 279 476 283
rect 1111 279 1115 283
rect 111 229 115 233
rect 192 215 196 219
rect 111 211 115 215
rect 1111 229 1115 233
rect 1111 211 1115 215
rect 472 191 476 195
rect 192 171 196 175
rect 111 149 115 153
rect 1111 149 1115 153
rect 111 131 115 135
rect 1111 131 1115 135
<< m2 >>
rect 134 1216 140 1217
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 222 1216 228 1217
rect 222 1212 223 1216
rect 227 1212 228 1216
rect 222 1211 228 1212
rect 310 1216 316 1217
rect 310 1212 311 1216
rect 315 1212 316 1216
rect 310 1211 316 1212
rect 398 1216 404 1217
rect 398 1212 399 1216
rect 403 1212 404 1216
rect 398 1211 404 1212
rect 110 1201 116 1202
rect 110 1197 111 1201
rect 115 1197 116 1201
rect 110 1196 116 1197
rect 1110 1201 1116 1202
rect 1110 1197 1111 1201
rect 1115 1197 1116 1201
rect 1110 1196 1116 1197
rect 202 1187 208 1188
rect 202 1186 203 1187
rect 197 1184 203 1186
rect 110 1183 116 1184
rect 110 1179 111 1183
rect 115 1179 116 1183
rect 202 1183 203 1184
rect 207 1183 208 1187
rect 290 1187 296 1188
rect 290 1186 291 1187
rect 285 1184 291 1186
rect 202 1182 208 1183
rect 290 1183 291 1184
rect 295 1183 296 1187
rect 378 1187 384 1188
rect 378 1186 379 1187
rect 373 1184 379 1186
rect 290 1182 296 1183
rect 378 1183 379 1184
rect 383 1183 384 1187
rect 378 1182 384 1183
rect 386 1187 392 1188
rect 386 1183 387 1187
rect 391 1186 392 1187
rect 391 1184 425 1186
rect 391 1183 392 1184
rect 386 1182 392 1183
rect 1110 1183 1116 1184
rect 110 1178 116 1179
rect 1110 1179 1111 1183
rect 1115 1179 1116 1183
rect 1110 1178 1116 1179
rect 142 1171 148 1172
rect 142 1167 143 1171
rect 147 1167 148 1171
rect 142 1166 148 1167
rect 230 1171 236 1172
rect 230 1167 231 1171
rect 235 1167 236 1171
rect 230 1166 236 1167
rect 318 1171 324 1172
rect 318 1167 319 1171
rect 323 1167 324 1171
rect 318 1166 324 1167
rect 406 1171 412 1172
rect 406 1167 407 1171
rect 411 1167 412 1171
rect 406 1166 412 1167
rect 202 1163 208 1164
rect 202 1159 203 1163
rect 207 1162 208 1163
rect 290 1163 296 1164
rect 207 1160 225 1162
rect 207 1159 208 1160
rect 202 1158 208 1159
rect 290 1159 291 1163
rect 295 1162 296 1163
rect 378 1163 384 1164
rect 295 1160 313 1162
rect 295 1159 296 1160
rect 290 1158 296 1159
rect 378 1159 379 1163
rect 383 1162 384 1163
rect 383 1160 401 1162
rect 383 1159 384 1160
rect 378 1158 384 1159
rect 150 1155 156 1156
rect 150 1154 151 1155
rect 141 1152 151 1154
rect 150 1151 151 1152
rect 155 1151 156 1155
rect 150 1150 156 1151
rect 202 1155 208 1156
rect 202 1151 203 1155
rect 207 1154 208 1155
rect 290 1155 296 1156
rect 207 1152 225 1154
rect 207 1151 208 1152
rect 202 1150 208 1151
rect 290 1151 291 1155
rect 295 1154 296 1155
rect 378 1155 384 1156
rect 295 1152 313 1154
rect 295 1151 296 1152
rect 290 1150 296 1151
rect 378 1151 379 1155
rect 383 1154 384 1155
rect 383 1152 401 1154
rect 383 1151 384 1152
rect 378 1150 384 1151
rect 142 1145 148 1146
rect 142 1141 143 1145
rect 147 1141 148 1145
rect 142 1140 148 1141
rect 230 1145 236 1146
rect 230 1141 231 1145
rect 235 1141 236 1145
rect 230 1140 236 1141
rect 318 1145 324 1146
rect 318 1141 319 1145
rect 323 1141 324 1145
rect 318 1140 324 1141
rect 406 1145 412 1146
rect 406 1141 407 1145
rect 411 1141 412 1145
rect 406 1140 412 1141
rect 110 1133 116 1134
rect 110 1129 111 1133
rect 115 1129 116 1133
rect 1110 1133 1116 1134
rect 202 1131 208 1132
rect 202 1130 203 1131
rect 110 1128 116 1129
rect 197 1128 203 1130
rect 202 1127 203 1128
rect 207 1127 208 1131
rect 290 1131 296 1132
rect 290 1130 291 1131
rect 285 1128 291 1130
rect 202 1126 208 1127
rect 290 1127 291 1128
rect 295 1127 296 1131
rect 378 1131 384 1132
rect 378 1130 379 1131
rect 373 1128 379 1130
rect 290 1126 296 1127
rect 378 1127 379 1128
rect 383 1127 384 1131
rect 1110 1129 1111 1133
rect 1115 1129 1116 1133
rect 1110 1128 1116 1129
rect 378 1126 384 1127
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 1110 1115 1116 1116
rect 384 1112 417 1114
rect 110 1110 116 1111
rect 382 1111 388 1112
rect 382 1107 383 1111
rect 387 1107 388 1111
rect 1110 1111 1111 1115
rect 1115 1111 1116 1115
rect 1110 1110 1116 1111
rect 382 1106 388 1107
rect 134 1100 140 1101
rect 134 1096 135 1100
rect 139 1096 140 1100
rect 134 1095 140 1096
rect 222 1100 228 1101
rect 222 1096 223 1100
rect 227 1096 228 1100
rect 222 1095 228 1096
rect 310 1100 316 1101
rect 310 1096 311 1100
rect 315 1096 316 1100
rect 310 1095 316 1096
rect 398 1100 404 1101
rect 398 1096 399 1100
rect 403 1096 404 1100
rect 398 1095 404 1096
rect 278 1088 284 1089
rect 278 1084 279 1088
rect 283 1084 284 1088
rect 278 1083 284 1084
rect 366 1088 372 1089
rect 366 1084 367 1088
rect 371 1084 372 1088
rect 366 1083 372 1084
rect 454 1088 460 1089
rect 454 1084 455 1088
rect 459 1084 460 1088
rect 454 1083 460 1084
rect 542 1088 548 1089
rect 542 1084 543 1088
rect 547 1084 548 1088
rect 542 1083 548 1084
rect 630 1088 636 1089
rect 630 1084 631 1088
rect 635 1084 636 1088
rect 630 1083 636 1084
rect 110 1073 116 1074
rect 110 1069 111 1073
rect 115 1069 116 1073
rect 110 1068 116 1069
rect 1110 1073 1116 1074
rect 1110 1069 1111 1073
rect 1115 1069 1116 1073
rect 1110 1068 1116 1069
rect 351 1059 357 1060
rect 351 1058 352 1059
rect 341 1056 352 1058
rect 110 1055 116 1056
rect 110 1051 111 1055
rect 115 1051 116 1055
rect 351 1055 352 1056
rect 356 1055 357 1059
rect 434 1059 440 1060
rect 434 1058 435 1059
rect 429 1056 435 1058
rect 351 1054 357 1055
rect 434 1055 435 1056
rect 439 1055 440 1059
rect 522 1059 528 1060
rect 522 1058 523 1059
rect 517 1056 523 1058
rect 434 1054 440 1055
rect 522 1055 523 1056
rect 527 1055 528 1059
rect 610 1059 616 1060
rect 610 1058 611 1059
rect 605 1056 611 1058
rect 522 1054 528 1055
rect 610 1055 611 1056
rect 615 1055 616 1059
rect 610 1054 616 1055
rect 618 1059 624 1060
rect 618 1055 619 1059
rect 623 1058 624 1059
rect 623 1056 657 1058
rect 623 1055 624 1056
rect 618 1054 624 1055
rect 1110 1055 1116 1056
rect 110 1050 116 1051
rect 1110 1051 1111 1055
rect 1115 1051 1116 1055
rect 1110 1050 1116 1051
rect 286 1043 292 1044
rect 286 1039 287 1043
rect 291 1039 292 1043
rect 286 1038 292 1039
rect 374 1043 380 1044
rect 374 1039 375 1043
rect 379 1039 380 1043
rect 374 1038 380 1039
rect 462 1043 468 1044
rect 462 1039 463 1043
rect 467 1039 468 1043
rect 462 1038 468 1039
rect 550 1043 556 1044
rect 550 1039 551 1043
rect 555 1039 556 1043
rect 550 1038 556 1039
rect 638 1043 644 1044
rect 638 1039 639 1043
rect 643 1039 644 1043
rect 638 1038 644 1039
rect 351 1035 357 1036
rect 351 1031 352 1035
rect 356 1034 357 1035
rect 434 1035 440 1036
rect 356 1032 369 1034
rect 356 1031 357 1032
rect 351 1030 357 1031
rect 434 1031 435 1035
rect 439 1034 440 1035
rect 522 1035 528 1036
rect 439 1032 457 1034
rect 439 1031 440 1032
rect 434 1030 440 1031
rect 522 1031 523 1035
rect 527 1034 528 1035
rect 610 1035 616 1036
rect 527 1032 545 1034
rect 527 1031 528 1032
rect 522 1030 528 1031
rect 610 1031 611 1035
rect 615 1034 616 1035
rect 615 1032 633 1034
rect 615 1031 616 1032
rect 610 1030 616 1031
rect 280 1026 282 1029
rect 382 1027 388 1028
rect 382 1026 383 1027
rect 280 1024 383 1026
rect 382 1023 383 1024
rect 387 1023 388 1027
rect 618 1027 624 1028
rect 618 1026 619 1027
rect 382 1022 388 1023
rect 532 1024 619 1026
rect 532 1018 534 1024
rect 618 1023 619 1024
rect 623 1023 624 1027
rect 618 1022 624 1023
rect 517 1016 534 1018
rect 578 1019 584 1020
rect 578 1015 579 1019
rect 583 1018 584 1019
rect 666 1019 672 1020
rect 583 1016 601 1018
rect 583 1015 584 1016
rect 578 1014 584 1015
rect 666 1015 667 1019
rect 671 1018 672 1019
rect 762 1019 768 1020
rect 671 1016 697 1018
rect 671 1015 672 1016
rect 666 1014 672 1015
rect 762 1015 763 1019
rect 767 1018 768 1019
rect 918 1019 924 1020
rect 918 1018 919 1019
rect 767 1016 801 1018
rect 909 1016 919 1018
rect 767 1015 768 1016
rect 762 1014 768 1015
rect 918 1015 919 1016
rect 923 1015 924 1019
rect 918 1014 924 1015
rect 970 1019 976 1020
rect 970 1015 971 1019
rect 975 1018 976 1019
rect 975 1016 1009 1018
rect 975 1015 976 1016
rect 970 1014 976 1015
rect 518 1009 524 1010
rect 518 1005 519 1009
rect 523 1005 524 1009
rect 518 1004 524 1005
rect 606 1009 612 1010
rect 606 1005 607 1009
rect 611 1005 612 1009
rect 606 1004 612 1005
rect 702 1009 708 1010
rect 702 1005 703 1009
rect 707 1005 708 1009
rect 702 1004 708 1005
rect 806 1009 812 1010
rect 806 1005 807 1009
rect 811 1005 812 1009
rect 806 1004 812 1005
rect 910 1009 916 1010
rect 910 1005 911 1009
rect 915 1005 916 1009
rect 910 1004 916 1005
rect 1014 1009 1020 1010
rect 1014 1005 1015 1009
rect 1019 1005 1020 1009
rect 1014 1004 1020 1005
rect 110 997 116 998
rect 110 993 111 997
rect 115 993 116 997
rect 1110 997 1116 998
rect 578 995 584 996
rect 578 994 579 995
rect 110 992 116 993
rect 573 992 579 994
rect 578 991 579 992
rect 583 991 584 995
rect 666 995 672 996
rect 666 994 667 995
rect 661 992 667 994
rect 578 990 584 991
rect 666 991 667 992
rect 671 991 672 995
rect 762 995 768 996
rect 762 994 763 995
rect 757 992 763 994
rect 666 990 672 991
rect 762 991 763 992
rect 767 991 768 995
rect 970 995 976 996
rect 970 994 971 995
rect 965 992 971 994
rect 762 990 768 991
rect 970 991 971 992
rect 975 991 976 995
rect 1110 993 1111 997
rect 1115 993 1116 997
rect 1110 992 1116 993
rect 970 990 976 991
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 806 979 812 980
rect 806 975 807 979
rect 811 978 812 979
rect 978 979 984 980
rect 811 976 817 978
rect 811 975 812 976
rect 806 974 812 975
rect 978 975 979 979
rect 983 978 984 979
rect 1110 979 1116 980
rect 983 976 1025 978
rect 983 975 984 976
rect 978 974 984 975
rect 1110 975 1111 979
rect 1115 975 1116 979
rect 1110 974 1116 975
rect 510 964 516 965
rect 510 960 511 964
rect 515 960 516 964
rect 510 959 516 960
rect 598 964 604 965
rect 598 960 599 964
rect 603 960 604 964
rect 598 959 604 960
rect 694 964 700 965
rect 694 960 695 964
rect 699 960 700 964
rect 694 959 700 960
rect 798 964 804 965
rect 798 960 799 964
rect 803 960 804 964
rect 798 959 804 960
rect 902 964 908 965
rect 902 960 903 964
rect 907 960 908 964
rect 902 959 908 960
rect 1006 964 1012 965
rect 1006 960 1007 964
rect 1011 960 1012 964
rect 1006 959 1012 960
rect 398 952 404 953
rect 398 948 399 952
rect 403 948 404 952
rect 398 947 404 948
rect 486 952 492 953
rect 486 948 487 952
rect 491 948 492 952
rect 486 947 492 948
rect 574 952 580 953
rect 574 948 575 952
rect 579 948 580 952
rect 574 947 580 948
rect 662 952 668 953
rect 662 948 663 952
rect 667 948 668 952
rect 662 947 668 948
rect 750 952 756 953
rect 750 948 751 952
rect 755 948 756 952
rect 750 947 756 948
rect 838 952 844 953
rect 838 948 839 952
rect 843 948 844 952
rect 838 947 844 948
rect 926 952 932 953
rect 926 948 927 952
rect 931 948 932 952
rect 926 947 932 948
rect 1014 952 1020 953
rect 1014 948 1015 952
rect 1019 948 1020 952
rect 1014 947 1020 948
rect 918 939 924 940
rect 918 938 919 939
rect 110 937 116 938
rect 110 933 111 937
rect 115 933 116 937
rect 897 936 919 938
rect 918 935 919 936
rect 923 935 924 939
rect 918 934 924 935
rect 1110 937 1116 938
rect 110 932 116 933
rect 1110 933 1111 937
rect 1115 933 1116 937
rect 1110 932 1116 933
rect 466 923 472 924
rect 466 922 467 923
rect 461 920 467 922
rect 110 919 116 920
rect 110 915 111 919
rect 115 915 116 919
rect 466 919 467 920
rect 471 919 472 923
rect 554 923 560 924
rect 554 922 555 923
rect 549 920 555 922
rect 466 918 472 919
rect 554 919 555 920
rect 559 919 560 923
rect 642 923 648 924
rect 554 918 560 919
rect 110 914 116 915
rect 636 916 638 921
rect 642 919 643 923
rect 647 922 648 923
rect 818 923 824 924
rect 818 922 819 923
rect 647 920 689 922
rect 813 920 819 922
rect 647 919 648 920
rect 642 918 648 919
rect 818 919 819 920
rect 823 919 824 923
rect 994 923 1000 924
rect 994 922 995 923
rect 989 920 995 922
rect 818 918 824 919
rect 994 919 995 920
rect 999 919 1000 923
rect 994 918 1000 919
rect 1007 923 1013 924
rect 1007 919 1008 923
rect 1012 922 1013 923
rect 1012 920 1041 922
rect 1012 919 1013 920
rect 1007 918 1013 919
rect 1110 919 1116 920
rect 636 915 644 916
rect 636 912 639 915
rect 638 911 639 912
rect 643 911 644 915
rect 1110 915 1111 919
rect 1115 915 1116 919
rect 1110 914 1116 915
rect 638 910 644 911
rect 406 907 412 908
rect 406 903 407 907
rect 411 903 412 907
rect 406 902 412 903
rect 494 907 500 908
rect 494 903 495 907
rect 499 903 500 907
rect 494 902 500 903
rect 582 907 588 908
rect 582 903 583 907
rect 587 903 588 907
rect 582 902 588 903
rect 670 907 676 908
rect 670 903 671 907
rect 675 903 676 907
rect 670 902 676 903
rect 758 907 764 908
rect 758 903 759 907
rect 763 903 764 907
rect 758 902 764 903
rect 846 907 852 908
rect 846 903 847 907
rect 851 903 852 907
rect 846 902 852 903
rect 934 907 940 908
rect 934 903 935 907
rect 939 903 940 907
rect 934 902 940 903
rect 1022 907 1028 908
rect 1022 903 1023 907
rect 1027 903 1028 907
rect 1022 902 1028 903
rect 210 899 216 900
rect 210 898 211 899
rect 140 896 211 898
rect 140 889 142 896
rect 210 895 211 896
rect 215 895 216 899
rect 350 899 356 900
rect 350 898 351 899
rect 210 894 216 895
rect 268 896 351 898
rect 268 889 270 896
rect 350 895 351 896
rect 355 895 356 899
rect 414 899 420 900
rect 414 898 415 899
rect 405 896 415 898
rect 350 894 356 895
rect 414 895 415 896
rect 419 895 420 899
rect 414 894 420 895
rect 466 899 472 900
rect 466 895 467 899
rect 471 898 472 899
rect 554 899 560 900
rect 471 896 489 898
rect 471 895 472 896
rect 466 894 472 895
rect 554 895 555 899
rect 559 898 560 899
rect 767 899 773 900
rect 767 898 768 899
rect 559 896 577 898
rect 669 896 686 898
rect 757 896 768 898
rect 559 895 560 896
rect 554 894 560 895
rect 446 891 452 892
rect 446 890 447 891
rect 437 888 447 890
rect 446 887 447 888
rect 451 887 452 891
rect 638 891 644 892
rect 638 890 639 891
rect 629 888 639 890
rect 446 886 452 887
rect 638 887 639 888
rect 643 887 644 891
rect 684 890 686 896
rect 767 895 768 896
rect 772 895 773 899
rect 767 894 773 895
rect 818 899 824 900
rect 818 895 819 899
rect 823 898 824 899
rect 994 899 1000 900
rect 823 896 841 898
rect 823 895 824 896
rect 818 894 824 895
rect 994 895 995 899
rect 999 898 1000 899
rect 999 896 1017 898
rect 999 895 1000 896
rect 994 894 1000 895
rect 806 891 812 892
rect 806 890 807 891
rect 684 888 807 890
rect 638 886 644 887
rect 806 887 807 888
rect 811 887 812 891
rect 806 886 812 887
rect 814 891 820 892
rect 814 887 815 891
rect 819 890 820 891
rect 928 890 930 893
rect 978 891 984 892
rect 978 890 979 891
rect 819 888 833 890
rect 928 888 979 890
rect 819 887 820 888
rect 814 886 820 887
rect 978 887 979 888
rect 983 887 984 891
rect 978 886 984 887
rect 1007 891 1013 892
rect 1007 887 1008 891
rect 1012 890 1013 891
rect 1012 888 1017 890
rect 1012 887 1013 888
rect 1007 886 1013 887
rect 142 881 148 882
rect 142 877 143 881
rect 147 877 148 881
rect 142 876 148 877
rect 270 881 276 882
rect 270 877 271 881
rect 275 877 276 881
rect 270 876 276 877
rect 438 881 444 882
rect 438 877 439 881
rect 443 877 444 881
rect 438 876 444 877
rect 630 881 636 882
rect 630 877 631 881
rect 635 877 636 881
rect 630 876 636 877
rect 838 881 844 882
rect 838 877 839 881
rect 843 877 844 881
rect 838 876 844 877
rect 1022 881 1028 882
rect 1022 877 1023 881
rect 1027 877 1028 881
rect 1022 876 1028 877
rect 814 871 820 872
rect 814 870 815 871
rect 110 869 116 870
rect 110 865 111 869
rect 115 865 116 869
rect 684 868 815 870
rect 684 865 686 868
rect 814 867 815 868
rect 819 867 820 871
rect 814 866 820 867
rect 1110 869 1116 870
rect 1110 865 1111 869
rect 1115 865 1116 869
rect 110 864 116 865
rect 1110 864 1116 865
rect 210 863 216 864
rect 210 859 211 863
rect 215 862 216 863
rect 350 863 356 864
rect 215 860 289 862
rect 215 859 216 860
rect 210 858 216 859
rect 350 859 351 863
rect 355 862 356 863
rect 738 863 744 864
rect 355 860 457 862
rect 355 859 356 860
rect 350 858 356 859
rect 738 859 739 863
rect 743 862 744 863
rect 743 860 857 862
rect 743 859 744 860
rect 738 858 744 859
rect 110 851 116 852
rect 110 847 111 851
rect 115 847 116 851
rect 110 846 116 847
rect 127 851 133 852
rect 127 847 128 851
rect 132 850 133 851
rect 1007 851 1013 852
rect 132 848 153 850
rect 132 847 133 848
rect 127 846 133 847
rect 1007 847 1008 851
rect 1012 850 1013 851
rect 1110 851 1116 852
rect 1012 848 1033 850
rect 1012 847 1013 848
rect 1007 846 1013 847
rect 1110 847 1111 851
rect 1115 847 1116 851
rect 1110 846 1116 847
rect 134 836 140 837
rect 134 832 135 836
rect 139 832 140 836
rect 134 831 140 832
rect 262 836 268 837
rect 262 832 263 836
rect 267 832 268 836
rect 262 831 268 832
rect 430 836 436 837
rect 430 832 431 836
rect 435 832 436 836
rect 430 831 436 832
rect 622 836 628 837
rect 622 832 623 836
rect 627 832 628 836
rect 622 831 628 832
rect 830 836 836 837
rect 830 832 831 836
rect 835 832 836 836
rect 830 831 836 832
rect 1014 836 1020 837
rect 1014 832 1015 836
rect 1019 832 1020 836
rect 1014 831 1020 832
rect 134 820 140 821
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 278 820 284 821
rect 278 816 279 820
rect 283 816 284 820
rect 278 815 284 816
rect 462 820 468 821
rect 462 816 463 820
rect 467 816 468 820
rect 462 815 468 816
rect 646 820 652 821
rect 646 816 647 820
rect 651 816 652 820
rect 646 815 652 816
rect 838 820 844 821
rect 838 816 839 820
rect 843 816 844 820
rect 838 815 844 816
rect 1014 820 1020 821
rect 1014 816 1015 820
rect 1019 816 1020 820
rect 1014 815 1020 816
rect 767 807 773 808
rect 110 805 116 806
rect 110 801 111 805
rect 115 801 116 805
rect 767 803 768 807
rect 772 806 773 807
rect 772 804 857 806
rect 1110 805 1116 806
rect 772 803 773 804
rect 767 802 773 803
rect 110 800 116 801
rect 1110 801 1111 805
rect 1115 801 1116 805
rect 1110 800 1116 801
rect 1014 795 1020 796
rect 218 791 224 792
rect 218 790 219 791
rect 197 788 219 790
rect 110 787 116 788
rect 110 783 111 787
rect 115 783 116 787
rect 218 787 219 788
rect 223 787 224 791
rect 399 791 405 792
rect 399 790 400 791
rect 341 788 400 790
rect 218 786 224 787
rect 399 787 400 788
rect 404 787 405 791
rect 566 791 572 792
rect 566 790 567 791
rect 525 788 567 790
rect 399 786 405 787
rect 566 787 567 788
rect 571 787 572 791
rect 566 786 572 787
rect 574 791 580 792
rect 574 787 575 791
rect 579 790 580 791
rect 1014 791 1015 795
rect 1019 791 1020 795
rect 1014 790 1020 791
rect 579 788 673 790
rect 1016 788 1041 790
rect 579 787 580 788
rect 574 786 580 787
rect 1110 787 1116 788
rect 110 782 116 783
rect 1110 783 1111 787
rect 1115 783 1116 787
rect 1110 782 1116 783
rect 142 775 148 776
rect 142 771 143 775
rect 147 771 148 775
rect 142 770 148 771
rect 286 775 292 776
rect 286 771 287 775
rect 291 771 292 775
rect 286 770 292 771
rect 470 775 476 776
rect 470 771 471 775
rect 475 771 476 775
rect 470 770 476 771
rect 654 775 660 776
rect 654 771 655 775
rect 659 771 660 775
rect 654 770 660 771
rect 846 775 852 776
rect 846 771 847 775
rect 851 771 852 775
rect 846 770 852 771
rect 1022 775 1028 776
rect 1022 771 1023 775
rect 1027 771 1028 775
rect 1022 770 1028 771
rect 127 767 133 768
rect 127 763 128 767
rect 132 766 133 767
rect 218 767 224 768
rect 132 764 137 766
rect 132 763 133 764
rect 127 762 133 763
rect 218 763 219 767
rect 223 766 224 767
rect 399 767 405 768
rect 223 764 281 766
rect 223 763 224 764
rect 218 762 224 763
rect 399 763 400 767
rect 404 766 405 767
rect 566 767 572 768
rect 404 764 465 766
rect 404 763 405 764
rect 399 762 405 763
rect 566 763 567 767
rect 571 766 572 767
rect 855 767 861 768
rect 855 766 856 767
rect 571 764 649 766
rect 845 764 856 766
rect 571 763 572 764
rect 566 762 572 763
rect 855 763 856 764
rect 860 763 861 767
rect 855 762 861 763
rect 1007 767 1013 768
rect 1007 763 1008 767
rect 1012 766 1013 767
rect 1012 764 1017 766
rect 1012 763 1013 764
rect 1007 762 1013 763
rect 190 747 196 748
rect 190 746 191 747
rect 181 744 191 746
rect 190 743 191 744
rect 195 743 196 747
rect 190 742 196 743
rect 242 747 248 748
rect 242 743 243 747
rect 247 746 248 747
rect 394 747 400 748
rect 247 744 297 746
rect 247 743 248 744
rect 242 742 248 743
rect 394 743 395 747
rect 399 746 400 747
rect 498 747 504 748
rect 399 744 425 746
rect 399 743 400 744
rect 394 742 400 743
rect 498 743 499 747
rect 503 746 504 747
rect 642 747 648 748
rect 503 744 561 746
rect 503 743 504 744
rect 498 742 504 743
rect 642 743 643 747
rect 647 746 648 747
rect 886 747 892 748
rect 886 746 887 747
rect 647 744 713 746
rect 877 744 887 746
rect 647 743 648 744
rect 642 742 648 743
rect 886 743 887 744
rect 891 743 892 747
rect 886 742 892 743
rect 1014 747 1020 748
rect 1014 743 1015 747
rect 1019 743 1020 747
rect 1014 742 1020 743
rect 182 737 188 738
rect 182 733 183 737
rect 187 733 188 737
rect 182 732 188 733
rect 302 737 308 738
rect 302 733 303 737
rect 307 733 308 737
rect 302 732 308 733
rect 430 737 436 738
rect 430 733 431 737
rect 435 733 436 737
rect 430 732 436 733
rect 566 737 572 738
rect 566 733 567 737
rect 571 733 572 737
rect 566 732 572 733
rect 718 737 724 738
rect 718 733 719 737
rect 723 733 724 737
rect 718 732 724 733
rect 878 737 884 738
rect 878 733 879 737
rect 883 733 884 737
rect 878 732 884 733
rect 1022 737 1028 738
rect 1022 733 1023 737
rect 1027 733 1028 737
rect 1022 732 1028 733
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 1110 725 1116 726
rect 242 723 248 724
rect 242 722 243 723
rect 110 720 116 721
rect 237 720 243 722
rect 242 719 243 720
rect 247 719 248 723
rect 394 723 400 724
rect 394 722 395 723
rect 357 720 395 722
rect 242 718 248 719
rect 394 719 395 720
rect 399 719 400 723
rect 498 723 504 724
rect 498 722 499 723
rect 485 720 499 722
rect 394 718 400 719
rect 498 719 499 720
rect 503 719 504 723
rect 642 723 648 724
rect 642 722 643 723
rect 621 720 643 722
rect 498 718 504 719
rect 642 719 643 720
rect 647 719 648 723
rect 1110 721 1111 725
rect 1115 721 1116 725
rect 1110 720 1116 721
rect 642 718 648 719
rect 855 719 861 720
rect 855 715 856 719
rect 860 718 861 719
rect 860 716 897 718
rect 860 715 861 716
rect 855 714 861 715
rect 110 707 116 708
rect 110 703 111 707
rect 115 703 116 707
rect 110 702 116 703
rect 634 707 640 708
rect 634 703 635 707
rect 639 706 640 707
rect 1007 707 1013 708
rect 639 704 729 706
rect 639 703 640 704
rect 634 702 640 703
rect 1007 703 1008 707
rect 1012 706 1013 707
rect 1110 707 1116 708
rect 1012 704 1033 706
rect 1012 703 1013 704
rect 1007 702 1013 703
rect 1110 703 1111 707
rect 1115 703 1116 707
rect 1110 702 1116 703
rect 174 692 180 693
rect 174 688 175 692
rect 179 688 180 692
rect 174 687 180 688
rect 294 692 300 693
rect 294 688 295 692
rect 299 688 300 692
rect 294 687 300 688
rect 422 692 428 693
rect 422 688 423 692
rect 427 688 428 692
rect 422 687 428 688
rect 558 692 564 693
rect 558 688 559 692
rect 563 688 564 692
rect 558 687 564 688
rect 710 692 716 693
rect 710 688 711 692
rect 715 688 716 692
rect 710 687 716 688
rect 870 692 876 693
rect 870 688 871 692
rect 875 688 876 692
rect 870 687 876 688
rect 1014 692 1020 693
rect 1014 688 1015 692
rect 1019 688 1020 692
rect 1014 687 1020 688
rect 342 668 348 669
rect 342 664 343 668
rect 347 664 348 668
rect 342 663 348 664
rect 454 668 460 669
rect 454 664 455 668
rect 459 664 460 668
rect 454 663 460 664
rect 582 668 588 669
rect 582 664 583 668
rect 587 664 588 668
rect 582 663 588 664
rect 718 668 724 669
rect 718 664 719 668
rect 723 664 724 668
rect 718 663 724 664
rect 862 668 868 669
rect 862 664 863 668
rect 867 664 868 668
rect 862 663 868 664
rect 1014 668 1020 669
rect 1014 664 1015 668
rect 1019 664 1020 668
rect 1014 663 1020 664
rect 110 653 116 654
rect 110 649 111 653
rect 115 649 116 653
rect 110 648 116 649
rect 1110 653 1116 654
rect 1110 649 1111 653
rect 1115 649 1116 653
rect 1110 648 1116 649
rect 410 639 416 640
rect 410 638 411 639
rect 405 636 411 638
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 410 635 411 636
rect 415 635 416 639
rect 530 639 536 640
rect 530 638 531 639
rect 517 636 531 638
rect 410 634 416 635
rect 530 635 531 636
rect 535 635 536 639
rect 662 639 668 640
rect 662 638 663 639
rect 645 636 663 638
rect 530 634 536 635
rect 662 635 663 636
rect 667 635 668 639
rect 802 639 808 640
rect 802 638 803 639
rect 781 636 803 638
rect 662 634 668 635
rect 802 635 803 636
rect 807 635 808 639
rect 802 634 808 635
rect 810 639 816 640
rect 810 635 811 639
rect 815 638 816 639
rect 998 639 1004 640
rect 815 636 889 638
rect 815 635 816 636
rect 810 634 816 635
rect 998 635 999 639
rect 1003 638 1004 639
rect 1003 636 1041 638
rect 1003 635 1004 636
rect 998 634 1004 635
rect 1110 635 1116 636
rect 110 630 116 631
rect 1110 631 1111 635
rect 1115 631 1116 635
rect 1110 630 1116 631
rect 350 623 356 624
rect 350 619 351 623
rect 355 619 356 623
rect 350 618 356 619
rect 462 623 468 624
rect 462 619 463 623
rect 467 619 468 623
rect 462 618 468 619
rect 590 623 596 624
rect 590 619 591 623
rect 595 619 596 623
rect 590 618 596 619
rect 726 623 732 624
rect 726 619 727 623
rect 731 619 732 623
rect 726 618 732 619
rect 870 623 876 624
rect 870 619 871 623
rect 875 619 876 623
rect 870 618 876 619
rect 1022 623 1028 624
rect 1022 619 1023 623
rect 1027 619 1028 623
rect 1022 618 1028 619
rect 358 615 364 616
rect 358 614 359 615
rect 349 612 359 614
rect 358 611 359 612
rect 363 611 364 615
rect 358 610 364 611
rect 410 615 416 616
rect 410 611 411 615
rect 415 614 416 615
rect 530 615 536 616
rect 415 612 457 614
rect 415 611 416 612
rect 410 610 416 611
rect 530 611 531 615
rect 535 614 536 615
rect 662 615 668 616
rect 535 612 585 614
rect 535 611 536 612
rect 530 610 536 611
rect 662 611 663 615
rect 667 614 668 615
rect 802 615 808 616
rect 667 612 721 614
rect 667 611 668 612
rect 662 610 668 611
rect 802 611 803 615
rect 807 614 808 615
rect 1007 615 1013 616
rect 807 612 865 614
rect 807 611 808 612
rect 802 610 808 611
rect 1007 611 1008 615
rect 1012 614 1013 615
rect 1012 612 1017 614
rect 1012 611 1013 612
rect 1007 610 1013 611
rect 550 599 556 600
rect 550 598 551 599
rect 541 596 551 598
rect 550 595 551 596
rect 555 595 556 599
rect 550 594 556 595
rect 602 599 608 600
rect 602 595 603 599
rect 607 598 608 599
rect 690 599 696 600
rect 607 596 625 598
rect 607 595 608 596
rect 602 594 608 595
rect 690 595 691 599
rect 695 598 696 599
rect 778 599 784 600
rect 695 596 713 598
rect 695 595 696 596
rect 690 594 696 595
rect 778 595 779 599
rect 783 598 784 599
rect 910 599 916 600
rect 910 598 911 599
rect 783 596 801 598
rect 901 596 911 598
rect 783 595 784 596
rect 778 594 784 595
rect 910 595 911 596
rect 915 595 916 599
rect 910 594 916 595
rect 998 599 1004 600
rect 998 595 999 599
rect 1003 595 1004 599
rect 998 594 1004 595
rect 542 589 548 590
rect 542 585 543 589
rect 547 585 548 589
rect 542 584 548 585
rect 630 589 636 590
rect 630 585 631 589
rect 635 585 636 589
rect 630 584 636 585
rect 718 589 724 590
rect 718 585 719 589
rect 723 585 724 589
rect 718 584 724 585
rect 806 589 812 590
rect 806 585 807 589
rect 811 585 812 589
rect 806 584 812 585
rect 902 589 908 590
rect 902 585 903 589
rect 907 585 908 589
rect 902 584 908 585
rect 1006 589 1012 590
rect 1006 585 1007 589
rect 1011 585 1012 589
rect 1006 584 1012 585
rect 110 577 116 578
rect 110 573 111 577
rect 115 573 116 577
rect 1110 577 1116 578
rect 602 575 608 576
rect 602 574 603 575
rect 110 572 116 573
rect 597 572 603 574
rect 602 571 603 572
rect 607 571 608 575
rect 690 575 696 576
rect 690 574 691 575
rect 685 572 691 574
rect 602 570 608 571
rect 690 571 691 572
rect 695 571 696 575
rect 778 575 784 576
rect 778 574 779 575
rect 773 572 779 574
rect 690 570 696 571
rect 778 571 779 572
rect 783 571 784 575
rect 1110 573 1111 577
rect 1115 573 1116 577
rect 1110 572 1116 573
rect 778 570 784 571
rect 886 571 892 572
rect 886 567 887 571
rect 891 570 892 571
rect 891 568 921 570
rect 891 567 892 568
rect 886 566 892 567
rect 110 559 116 560
rect 110 555 111 559
rect 115 555 116 559
rect 110 554 116 555
rect 806 559 812 560
rect 806 555 807 559
rect 811 558 812 559
rect 990 559 996 560
rect 811 556 817 558
rect 811 555 812 556
rect 806 554 812 555
rect 990 555 991 559
rect 995 558 996 559
rect 1110 559 1116 560
rect 995 556 1017 558
rect 995 555 996 556
rect 990 554 996 555
rect 1110 555 1111 559
rect 1115 555 1116 559
rect 1110 554 1116 555
rect 534 544 540 545
rect 534 540 535 544
rect 539 540 540 544
rect 534 539 540 540
rect 622 544 628 545
rect 622 540 623 544
rect 627 540 628 544
rect 622 539 628 540
rect 710 544 716 545
rect 710 540 711 544
rect 715 540 716 544
rect 710 539 716 540
rect 798 544 804 545
rect 798 540 799 544
rect 803 540 804 544
rect 798 539 804 540
rect 894 544 900 545
rect 894 540 895 544
rect 899 540 900 544
rect 894 539 900 540
rect 998 544 1004 545
rect 998 540 999 544
rect 1003 540 1004 544
rect 998 539 1004 540
rect 478 524 484 525
rect 478 520 479 524
rect 483 520 484 524
rect 478 519 484 520
rect 566 524 572 525
rect 566 520 567 524
rect 571 520 572 524
rect 566 519 572 520
rect 654 524 660 525
rect 654 520 655 524
rect 659 520 660 524
rect 654 519 660 520
rect 742 524 748 525
rect 742 520 743 524
rect 747 520 748 524
rect 742 519 748 520
rect 830 524 836 525
rect 830 520 831 524
rect 835 520 836 524
rect 830 519 836 520
rect 918 524 924 525
rect 918 520 919 524
rect 923 520 924 524
rect 918 519 924 520
rect 910 511 916 512
rect 110 509 116 510
rect 110 505 111 509
rect 115 505 116 509
rect 910 507 911 511
rect 915 510 916 511
rect 915 508 937 510
rect 1110 509 1116 510
rect 915 507 916 508
rect 910 506 916 507
rect 110 504 116 505
rect 1110 505 1111 509
rect 1115 505 1116 509
rect 1110 504 1116 505
rect 546 495 552 496
rect 546 494 547 495
rect 541 492 547 494
rect 110 491 116 492
rect 110 487 111 491
rect 115 487 116 491
rect 546 491 547 492
rect 551 491 552 495
rect 546 490 552 491
rect 559 495 565 496
rect 559 491 560 495
rect 564 494 565 495
rect 634 495 640 496
rect 564 492 593 494
rect 564 491 565 492
rect 559 490 565 491
rect 634 491 635 495
rect 639 494 640 495
rect 726 495 732 496
rect 639 492 681 494
rect 639 491 640 492
rect 634 490 640 491
rect 726 491 727 495
rect 731 494 732 495
rect 814 495 820 496
rect 731 492 769 494
rect 731 491 732 492
rect 726 490 732 491
rect 814 491 815 495
rect 819 494 820 495
rect 819 492 857 494
rect 819 491 820 492
rect 814 490 820 491
rect 1110 491 1116 492
rect 110 486 116 487
rect 1110 487 1111 491
rect 1115 487 1116 491
rect 1110 486 1116 487
rect 486 479 492 480
rect 486 475 487 479
rect 491 475 492 479
rect 486 474 492 475
rect 574 479 580 480
rect 574 475 575 479
rect 579 475 580 479
rect 574 474 580 475
rect 662 479 668 480
rect 662 475 663 479
rect 667 475 668 479
rect 662 474 668 475
rect 750 479 756 480
rect 750 475 751 479
rect 755 475 756 479
rect 750 474 756 475
rect 838 479 844 480
rect 838 475 839 479
rect 843 475 844 479
rect 838 474 844 475
rect 926 479 932 480
rect 926 475 927 479
rect 931 475 932 479
rect 926 474 932 475
rect 546 471 552 472
rect 546 467 547 471
rect 551 470 552 471
rect 806 471 812 472
rect 551 468 569 470
rect 551 467 552 468
rect 546 466 552 467
rect 806 467 807 471
rect 811 470 812 471
rect 918 471 924 472
rect 811 468 833 470
rect 811 467 812 468
rect 806 466 812 467
rect 918 467 919 471
rect 923 467 924 471
rect 918 466 924 467
rect 442 463 448 464
rect 442 462 443 463
rect 268 460 443 462
rect 268 453 270 460
rect 442 459 443 460
rect 447 459 448 463
rect 480 462 482 465
rect 634 463 640 464
rect 634 462 635 463
rect 480 460 635 462
rect 442 458 448 459
rect 634 459 635 460
rect 639 459 640 463
rect 656 462 658 465
rect 726 463 732 464
rect 726 462 727 463
rect 656 460 727 462
rect 634 458 640 459
rect 726 459 727 460
rect 731 459 732 463
rect 744 462 746 465
rect 814 463 820 464
rect 814 462 815 463
rect 744 460 815 462
rect 726 458 732 459
rect 814 459 815 460
rect 819 459 820 463
rect 814 458 820 459
rect 342 455 348 456
rect 342 451 343 455
rect 347 454 348 455
rect 494 455 500 456
rect 494 454 495 455
rect 347 452 369 454
rect 485 452 495 454
rect 347 451 348 452
rect 342 450 348 451
rect 494 451 495 452
rect 499 451 500 455
rect 494 450 500 451
rect 559 455 565 456
rect 559 451 560 455
rect 564 454 565 455
rect 663 455 669 456
rect 564 452 593 454
rect 564 451 565 452
rect 559 450 565 451
rect 663 451 664 455
rect 668 454 669 455
rect 854 455 860 456
rect 854 454 855 455
rect 668 452 713 454
rect 845 452 855 454
rect 668 451 669 452
rect 663 450 669 451
rect 854 451 855 452
rect 859 451 860 455
rect 990 455 996 456
rect 990 454 991 455
rect 981 452 991 454
rect 854 450 860 451
rect 990 451 991 452
rect 995 451 996 455
rect 990 450 996 451
rect 270 445 276 446
rect 270 441 271 445
rect 275 441 276 445
rect 270 440 276 441
rect 374 445 380 446
rect 374 441 375 445
rect 379 441 380 445
rect 374 440 380 441
rect 486 445 492 446
rect 486 441 487 445
rect 491 441 492 445
rect 486 440 492 441
rect 598 445 604 446
rect 598 441 599 445
rect 603 441 604 445
rect 598 440 604 441
rect 718 445 724 446
rect 718 441 719 445
rect 723 441 724 445
rect 718 440 724 441
rect 846 445 852 446
rect 846 441 847 445
rect 851 441 852 445
rect 846 440 852 441
rect 982 445 988 446
rect 982 441 983 445
rect 987 441 988 445
rect 982 440 988 441
rect 110 433 116 434
rect 110 429 111 433
rect 115 429 116 433
rect 1110 433 1116 434
rect 342 431 348 432
rect 342 430 343 431
rect 110 428 116 429
rect 325 428 343 430
rect 342 427 343 428
rect 347 427 348 431
rect 663 431 669 432
rect 663 430 664 431
rect 653 428 664 430
rect 342 426 348 427
rect 442 427 448 428
rect 442 423 443 427
rect 447 426 448 427
rect 663 427 664 428
rect 668 427 669 431
rect 918 431 924 432
rect 918 430 919 431
rect 901 428 919 430
rect 663 426 669 427
rect 918 427 919 428
rect 923 427 924 431
rect 1110 429 1111 433
rect 1115 429 1116 433
rect 1110 428 1116 429
rect 918 426 924 427
rect 447 424 505 426
rect 447 423 448 424
rect 442 422 448 423
rect 110 415 116 416
rect 110 411 111 415
rect 115 411 116 415
rect 446 415 452 416
rect 446 414 447 415
rect 425 412 447 414
rect 110 410 116 411
rect 446 411 447 412
rect 451 411 452 415
rect 446 410 452 411
rect 666 415 672 416
rect 666 411 667 415
rect 671 414 672 415
rect 967 415 973 416
rect 671 412 729 414
rect 671 411 672 412
rect 666 410 672 411
rect 967 411 968 415
rect 972 414 973 415
rect 1110 415 1116 416
rect 972 412 993 414
rect 972 411 973 412
rect 967 410 973 411
rect 1110 411 1111 415
rect 1115 411 1116 415
rect 1110 410 1116 411
rect 262 400 268 401
rect 262 396 263 400
rect 267 396 268 400
rect 262 395 268 396
rect 366 400 372 401
rect 366 396 367 400
rect 371 396 372 400
rect 366 395 372 396
rect 478 400 484 401
rect 478 396 479 400
rect 483 396 484 400
rect 478 395 484 396
rect 590 400 596 401
rect 590 396 591 400
rect 595 396 596 400
rect 590 395 596 396
rect 710 400 716 401
rect 710 396 711 400
rect 715 396 716 400
rect 710 395 716 396
rect 838 400 844 401
rect 838 396 839 400
rect 843 396 844 400
rect 838 395 844 396
rect 974 400 980 401
rect 974 396 975 400
rect 979 396 980 400
rect 974 395 980 396
rect 494 391 500 392
rect 494 387 495 391
rect 499 390 500 391
rect 666 391 672 392
rect 666 390 667 391
rect 499 388 667 390
rect 499 387 500 388
rect 494 386 500 387
rect 666 387 667 388
rect 671 387 672 391
rect 666 386 672 387
rect 134 384 140 385
rect 134 380 135 384
rect 139 380 140 384
rect 134 379 140 380
rect 262 384 268 385
rect 262 380 263 384
rect 267 380 268 384
rect 262 379 268 380
rect 430 384 436 385
rect 430 380 431 384
rect 435 380 436 384
rect 430 379 436 380
rect 606 384 612 385
rect 606 380 607 384
rect 611 380 612 384
rect 606 379 612 380
rect 790 384 796 385
rect 790 380 791 384
rect 795 380 796 384
rect 790 379 796 380
rect 974 384 980 385
rect 974 380 975 384
rect 979 380 980 384
rect 974 379 980 380
rect 858 371 864 372
rect 858 370 859 371
rect 110 369 116 370
rect 110 365 111 369
rect 115 365 116 369
rect 849 368 859 370
rect 858 367 859 368
rect 863 367 864 371
rect 858 366 864 367
rect 1110 369 1116 370
rect 110 364 116 365
rect 1110 365 1111 369
rect 1115 365 1116 369
rect 1110 364 1116 365
rect 127 355 133 356
rect 110 351 116 352
rect 110 347 111 351
rect 115 347 116 351
rect 127 351 128 355
rect 132 354 133 355
rect 202 355 208 356
rect 132 352 161 354
rect 132 351 133 352
rect 127 350 133 351
rect 202 351 203 355
rect 207 354 208 355
rect 530 355 536 356
rect 530 354 531 355
rect 207 352 289 354
rect 493 352 531 354
rect 207 351 208 352
rect 202 350 208 351
rect 530 351 531 352
rect 535 351 536 355
rect 530 350 536 351
rect 538 355 544 356
rect 538 351 539 355
rect 543 354 544 355
rect 543 352 633 354
rect 543 351 544 352
rect 538 350 544 351
rect 110 346 116 347
rect 142 339 148 340
rect 142 335 143 339
rect 147 335 148 339
rect 142 334 148 335
rect 270 339 276 340
rect 270 335 271 339
rect 275 335 276 339
rect 270 334 276 335
rect 438 339 444 340
rect 438 335 439 339
rect 443 335 444 339
rect 438 334 444 335
rect 614 339 620 340
rect 614 335 615 339
rect 619 335 620 339
rect 614 334 620 335
rect 798 339 804 340
rect 798 335 799 339
rect 803 335 804 339
rect 798 334 804 335
rect 982 339 988 340
rect 982 335 983 339
rect 987 335 988 339
rect 982 334 988 335
rect 150 331 156 332
rect 150 330 151 331
rect 141 328 151 330
rect 150 327 151 328
rect 155 327 156 331
rect 278 331 284 332
rect 278 330 279 331
rect 269 328 279 330
rect 150 326 156 327
rect 278 327 279 328
rect 283 327 284 331
rect 446 331 452 332
rect 446 330 447 331
rect 437 328 447 330
rect 278 326 284 327
rect 446 327 447 328
rect 451 327 452 331
rect 446 326 452 327
rect 530 331 536 332
rect 530 327 531 331
rect 535 330 536 331
rect 790 331 796 332
rect 535 328 609 330
rect 535 327 536 328
rect 530 326 536 327
rect 790 327 791 331
rect 795 327 796 331
rect 938 331 944 332
rect 938 330 939 331
rect 790 326 796 327
rect 852 328 939 330
rect 127 323 133 324
rect 127 319 128 323
rect 132 322 133 323
rect 222 323 228 324
rect 132 320 137 322
rect 132 319 133 320
rect 127 318 133 319
rect 222 319 223 323
rect 227 322 228 323
rect 394 323 400 324
rect 227 320 297 322
rect 227 319 228 320
rect 222 318 228 319
rect 394 319 395 323
rect 399 322 400 323
rect 678 323 684 324
rect 678 322 679 323
rect 399 320 481 322
rect 669 320 679 322
rect 399 319 400 320
rect 394 318 400 319
rect 678 319 679 320
rect 683 319 684 323
rect 852 321 854 328
rect 938 327 939 328
rect 943 327 944 331
rect 938 326 944 327
rect 967 331 973 332
rect 967 327 968 331
rect 972 330 973 331
rect 972 328 977 330
rect 972 327 973 328
rect 967 326 973 327
rect 1036 322 1038 353
rect 1110 351 1116 352
rect 1110 347 1111 351
rect 1115 347 1116 351
rect 1110 346 1116 347
rect 1021 320 1038 322
rect 678 318 684 319
rect 142 313 148 314
rect 142 309 143 313
rect 147 309 148 313
rect 142 308 148 309
rect 302 313 308 314
rect 302 309 303 313
rect 307 309 308 313
rect 302 308 308 309
rect 486 313 492 314
rect 486 309 487 313
rect 491 309 492 313
rect 486 308 492 309
rect 670 313 676 314
rect 670 309 671 313
rect 675 309 676 313
rect 670 308 676 309
rect 854 313 860 314
rect 854 309 855 313
rect 859 309 860 313
rect 854 308 860 309
rect 1022 313 1028 314
rect 1022 309 1023 313
rect 1027 309 1028 313
rect 1022 308 1028 309
rect 110 301 116 302
rect 110 297 111 301
rect 115 297 116 301
rect 1110 301 1116 302
rect 222 299 228 300
rect 222 298 223 299
rect 110 296 116 297
rect 197 296 223 298
rect 222 295 223 296
rect 227 295 228 299
rect 394 299 400 300
rect 394 298 395 299
rect 357 296 395 298
rect 222 294 228 295
rect 394 295 395 296
rect 399 295 400 299
rect 790 299 796 300
rect 790 298 791 299
rect 725 296 791 298
rect 394 294 400 295
rect 790 295 791 296
rect 795 295 796 299
rect 1110 297 1111 301
rect 1115 297 1116 301
rect 1110 296 1116 297
rect 790 294 796 295
rect 938 295 944 296
rect 938 291 939 295
rect 943 294 944 295
rect 943 292 1041 294
rect 943 291 944 292
rect 938 290 944 291
rect 110 283 116 284
rect 110 279 111 283
rect 115 279 116 283
rect 110 278 116 279
rect 471 283 477 284
rect 471 279 472 283
rect 476 282 477 283
rect 1110 283 1116 284
rect 476 280 497 282
rect 905 280 918 282
rect 476 279 477 280
rect 471 278 477 279
rect 914 279 920 280
rect 914 275 915 279
rect 919 275 920 279
rect 1110 279 1111 283
rect 1115 279 1116 283
rect 1110 278 1116 279
rect 914 274 920 275
rect 134 268 140 269
rect 134 264 135 268
rect 139 264 140 268
rect 134 263 140 264
rect 294 268 300 269
rect 294 264 295 268
rect 299 264 300 268
rect 294 263 300 264
rect 478 268 484 269
rect 478 264 479 268
rect 483 264 484 268
rect 478 263 484 264
rect 662 268 668 269
rect 662 264 663 268
rect 667 264 668 268
rect 662 263 668 264
rect 846 268 852 269
rect 846 264 847 268
rect 851 264 852 268
rect 846 263 852 264
rect 1014 268 1020 269
rect 1014 264 1015 268
rect 1019 264 1020 268
rect 1014 263 1020 264
rect 198 248 204 249
rect 198 244 199 248
rect 203 244 204 248
rect 198 243 204 244
rect 342 248 348 249
rect 342 244 343 248
rect 347 244 348 248
rect 342 243 348 244
rect 478 248 484 249
rect 478 244 479 248
rect 483 244 484 248
rect 478 243 484 244
rect 614 248 620 249
rect 614 244 615 248
rect 619 244 620 248
rect 614 243 620 244
rect 750 248 756 249
rect 750 244 751 248
rect 755 244 756 248
rect 750 243 756 244
rect 894 248 900 249
rect 894 244 895 248
rect 899 244 900 248
rect 894 243 900 244
rect 1014 248 1020 249
rect 1014 244 1015 248
rect 1019 244 1020 248
rect 1014 243 1020 244
rect 682 235 688 236
rect 682 234 683 235
rect 110 233 116 234
rect 110 229 111 233
rect 115 229 116 233
rect 673 232 683 234
rect 682 231 683 232
rect 687 231 688 235
rect 682 230 688 231
rect 1110 233 1116 234
rect 110 228 116 229
rect 1110 229 1111 233
rect 1115 229 1116 233
rect 1110 228 1116 229
rect 1014 223 1020 224
rect 191 219 197 220
rect 110 215 116 216
rect 110 211 111 215
rect 115 211 116 215
rect 191 215 192 219
rect 196 218 197 219
rect 266 219 272 220
rect 196 216 225 218
rect 196 215 197 216
rect 191 214 197 215
rect 266 215 267 219
rect 271 218 272 219
rect 422 219 428 220
rect 271 216 369 218
rect 271 215 272 216
rect 266 214 272 215
rect 422 215 423 219
rect 427 218 428 219
rect 694 219 700 220
rect 427 216 505 218
rect 427 215 428 216
rect 422 214 428 215
rect 694 215 695 219
rect 699 218 700 219
rect 1002 219 1008 220
rect 1002 218 1003 219
rect 699 216 777 218
rect 957 216 1003 218
rect 699 215 700 216
rect 694 214 700 215
rect 1002 215 1003 216
rect 1007 215 1008 219
rect 1014 219 1015 223
rect 1019 219 1020 223
rect 1014 218 1020 219
rect 1016 216 1041 218
rect 1002 214 1008 215
rect 1110 215 1116 216
rect 110 210 116 211
rect 1110 211 1111 215
rect 1115 211 1116 215
rect 1110 210 1116 211
rect 206 203 212 204
rect 206 199 207 203
rect 211 199 212 203
rect 206 198 212 199
rect 350 203 356 204
rect 350 199 351 203
rect 355 199 356 203
rect 350 198 356 199
rect 486 203 492 204
rect 486 199 487 203
rect 491 199 492 203
rect 486 198 492 199
rect 622 203 628 204
rect 622 199 623 203
rect 627 199 628 203
rect 622 198 628 199
rect 758 203 764 204
rect 758 199 759 203
rect 763 199 764 203
rect 758 198 764 199
rect 902 203 908 204
rect 902 199 903 203
rect 907 199 908 203
rect 902 198 908 199
rect 1022 203 1028 204
rect 1022 199 1023 203
rect 1027 199 1028 203
rect 1022 198 1028 199
rect 471 195 477 196
rect 471 191 472 195
rect 476 194 477 195
rect 910 195 916 196
rect 910 194 911 195
rect 476 192 481 194
rect 901 192 911 194
rect 476 191 477 192
rect 471 190 477 191
rect 910 191 911 192
rect 915 191 916 195
rect 910 190 916 191
rect 1002 195 1008 196
rect 1002 191 1003 195
rect 1007 194 1008 195
rect 1007 192 1017 194
rect 1007 191 1008 192
rect 1002 190 1008 191
rect 200 186 202 189
rect 266 187 272 188
rect 266 186 267 187
rect 200 184 267 186
rect 266 183 267 184
rect 271 183 272 187
rect 344 186 346 189
rect 422 187 428 188
rect 422 186 423 187
rect 344 184 423 186
rect 266 182 272 183
rect 422 183 423 184
rect 427 183 428 187
rect 616 186 618 189
rect 694 187 700 188
rect 694 186 695 187
rect 616 184 695 186
rect 422 182 428 183
rect 694 183 695 184
rect 699 183 700 187
rect 752 186 754 189
rect 826 187 832 188
rect 826 186 827 187
rect 752 184 827 186
rect 694 182 700 183
rect 826 183 827 184
rect 831 183 832 187
rect 826 182 832 183
rect 1002 183 1008 184
rect 1002 182 1003 183
rect 932 180 1003 182
rect 191 175 197 176
rect 191 171 192 175
rect 196 174 197 175
rect 290 175 296 176
rect 196 172 225 174
rect 196 171 197 172
rect 191 170 197 171
rect 290 171 291 175
rect 295 174 296 175
rect 378 175 384 176
rect 295 172 313 174
rect 295 171 296 172
rect 290 170 296 171
rect 378 171 379 175
rect 383 174 384 175
rect 466 175 472 176
rect 383 172 401 174
rect 383 171 384 172
rect 378 170 384 171
rect 466 171 467 175
rect 471 174 472 175
rect 554 175 560 176
rect 471 172 489 174
rect 471 171 472 172
rect 466 170 472 171
rect 554 171 555 175
rect 559 174 560 175
rect 642 175 648 176
rect 559 172 577 174
rect 559 171 560 172
rect 554 170 560 171
rect 642 171 643 175
rect 647 174 648 175
rect 730 175 736 176
rect 647 172 665 174
rect 647 171 648 172
rect 642 170 648 171
rect 730 171 731 175
rect 735 174 736 175
rect 818 175 824 176
rect 735 172 753 174
rect 735 171 736 172
rect 730 170 736 171
rect 818 171 819 175
rect 823 174 824 175
rect 823 172 841 174
rect 932 173 934 180
rect 1002 179 1003 180
rect 1007 179 1008 183
rect 1002 178 1008 179
rect 1014 175 1020 176
rect 823 171 824 172
rect 818 170 824 171
rect 1014 171 1015 175
rect 1019 171 1020 175
rect 1014 170 1020 171
rect 230 165 236 166
rect 230 161 231 165
rect 235 161 236 165
rect 230 160 236 161
rect 318 165 324 166
rect 318 161 319 165
rect 323 161 324 165
rect 318 160 324 161
rect 406 165 412 166
rect 406 161 407 165
rect 411 161 412 165
rect 406 160 412 161
rect 494 165 500 166
rect 494 161 495 165
rect 499 161 500 165
rect 494 160 500 161
rect 582 165 588 166
rect 582 161 583 165
rect 587 161 588 165
rect 582 160 588 161
rect 670 165 676 166
rect 670 161 671 165
rect 675 161 676 165
rect 670 160 676 161
rect 758 165 764 166
rect 758 161 759 165
rect 763 161 764 165
rect 758 160 764 161
rect 846 165 852 166
rect 846 161 847 165
rect 851 161 852 165
rect 846 160 852 161
rect 934 165 940 166
rect 934 161 935 165
rect 939 161 940 165
rect 934 160 940 161
rect 1022 165 1028 166
rect 1022 161 1023 165
rect 1027 161 1028 165
rect 1022 160 1028 161
rect 110 153 116 154
rect 110 149 111 153
rect 115 149 116 153
rect 1110 153 1116 154
rect 290 151 296 152
rect 290 150 291 151
rect 110 148 116 149
rect 285 148 291 150
rect 290 147 291 148
rect 295 147 296 151
rect 378 151 384 152
rect 378 150 379 151
rect 373 148 379 150
rect 290 146 296 147
rect 378 147 379 148
rect 383 147 384 151
rect 466 151 472 152
rect 466 150 467 151
rect 461 148 467 150
rect 378 146 384 147
rect 466 147 467 148
rect 471 147 472 151
rect 554 151 560 152
rect 554 150 555 151
rect 549 148 555 150
rect 466 146 472 147
rect 554 147 555 148
rect 559 147 560 151
rect 642 151 648 152
rect 642 150 643 151
rect 637 148 643 150
rect 554 146 560 147
rect 642 147 643 148
rect 647 147 648 151
rect 730 151 736 152
rect 730 150 731 151
rect 725 148 731 150
rect 642 146 648 147
rect 730 147 731 148
rect 735 147 736 151
rect 818 151 824 152
rect 818 150 819 151
rect 813 148 819 150
rect 730 146 736 147
rect 818 147 819 148
rect 823 147 824 151
rect 1110 149 1111 153
rect 1115 149 1116 153
rect 1110 148 1116 149
rect 818 146 824 147
rect 826 147 832 148
rect 826 143 827 147
rect 831 146 832 147
rect 1002 147 1008 148
rect 831 144 865 146
rect 831 143 832 144
rect 826 142 832 143
rect 1002 143 1003 147
rect 1007 146 1008 147
rect 1007 144 1041 146
rect 1007 143 1008 144
rect 1002 142 1008 143
rect 110 135 116 136
rect 110 131 111 135
rect 115 131 116 135
rect 110 130 116 131
rect 1110 135 1116 136
rect 1110 131 1111 135
rect 1115 131 1116 135
rect 1110 130 1116 131
rect 222 120 228 121
rect 222 116 223 120
rect 227 116 228 120
rect 222 115 228 116
rect 310 120 316 121
rect 310 116 311 120
rect 315 116 316 120
rect 310 115 316 116
rect 398 120 404 121
rect 398 116 399 120
rect 403 116 404 120
rect 398 115 404 116
rect 486 120 492 121
rect 486 116 487 120
rect 491 116 492 120
rect 486 115 492 116
rect 574 120 580 121
rect 574 116 575 120
rect 579 116 580 120
rect 574 115 580 116
rect 662 120 668 121
rect 662 116 663 120
rect 667 116 668 120
rect 662 115 668 116
rect 750 120 756 121
rect 750 116 751 120
rect 755 116 756 120
rect 750 115 756 116
rect 838 120 844 121
rect 838 116 839 120
rect 843 116 844 120
rect 838 115 844 116
rect 926 120 932 121
rect 926 116 927 120
rect 931 116 932 120
rect 926 115 932 116
rect 1014 120 1020 121
rect 1014 116 1015 120
rect 1019 116 1020 120
rect 1014 115 1020 116
<< m3c >>
rect 135 1212 139 1216
rect 223 1212 227 1216
rect 311 1212 315 1216
rect 399 1212 403 1216
rect 111 1197 115 1201
rect 1111 1197 1115 1201
rect 111 1179 115 1183
rect 203 1183 207 1187
rect 291 1183 295 1187
rect 379 1183 383 1187
rect 387 1183 391 1187
rect 1111 1179 1115 1183
rect 143 1167 147 1171
rect 231 1167 235 1171
rect 319 1167 323 1171
rect 407 1167 411 1171
rect 203 1159 207 1163
rect 291 1159 295 1163
rect 379 1159 383 1163
rect 151 1151 155 1155
rect 203 1151 207 1155
rect 291 1151 295 1155
rect 379 1151 383 1155
rect 143 1141 147 1145
rect 231 1141 235 1145
rect 319 1141 323 1145
rect 407 1141 411 1145
rect 111 1129 115 1133
rect 203 1127 207 1131
rect 291 1127 295 1131
rect 379 1127 383 1131
rect 1111 1129 1115 1133
rect 111 1111 115 1115
rect 383 1107 387 1111
rect 1111 1111 1115 1115
rect 135 1096 139 1100
rect 223 1096 227 1100
rect 311 1096 315 1100
rect 399 1096 403 1100
rect 279 1084 283 1088
rect 367 1084 371 1088
rect 455 1084 459 1088
rect 543 1084 547 1088
rect 631 1084 635 1088
rect 111 1069 115 1073
rect 1111 1069 1115 1073
rect 111 1051 115 1055
rect 435 1055 439 1059
rect 523 1055 527 1059
rect 611 1055 615 1059
rect 619 1055 623 1059
rect 1111 1051 1115 1055
rect 287 1039 291 1043
rect 375 1039 379 1043
rect 463 1039 467 1043
rect 551 1039 555 1043
rect 639 1039 643 1043
rect 435 1031 439 1035
rect 523 1031 527 1035
rect 611 1031 615 1035
rect 383 1023 387 1027
rect 619 1023 623 1027
rect 579 1015 583 1019
rect 667 1015 671 1019
rect 763 1015 767 1019
rect 919 1015 923 1019
rect 971 1015 975 1019
rect 519 1005 523 1009
rect 607 1005 611 1009
rect 703 1005 707 1009
rect 807 1005 811 1009
rect 911 1005 915 1009
rect 1015 1005 1019 1009
rect 111 993 115 997
rect 579 991 583 995
rect 667 991 671 995
rect 763 991 767 995
rect 971 991 975 995
rect 1111 993 1115 997
rect 111 975 115 979
rect 807 975 811 979
rect 979 975 983 979
rect 1111 975 1115 979
rect 511 960 515 964
rect 599 960 603 964
rect 695 960 699 964
rect 799 960 803 964
rect 903 960 907 964
rect 1007 960 1011 964
rect 399 948 403 952
rect 487 948 491 952
rect 575 948 579 952
rect 663 948 667 952
rect 751 948 755 952
rect 839 948 843 952
rect 927 948 931 952
rect 1015 948 1019 952
rect 111 933 115 937
rect 919 935 923 939
rect 1111 933 1115 937
rect 111 915 115 919
rect 467 919 471 923
rect 555 919 559 923
rect 643 919 647 923
rect 819 919 823 923
rect 995 919 999 923
rect 639 911 643 915
rect 1111 915 1115 919
rect 407 903 411 907
rect 495 903 499 907
rect 583 903 587 907
rect 671 903 675 907
rect 759 903 763 907
rect 847 903 851 907
rect 935 903 939 907
rect 1023 903 1027 907
rect 211 895 215 899
rect 351 895 355 899
rect 415 895 419 899
rect 467 895 471 899
rect 555 895 559 899
rect 447 887 451 891
rect 639 887 643 891
rect 819 895 823 899
rect 995 895 999 899
rect 807 887 811 891
rect 815 887 819 891
rect 979 887 983 891
rect 143 877 147 881
rect 271 877 275 881
rect 439 877 443 881
rect 631 877 635 881
rect 839 877 843 881
rect 1023 877 1027 881
rect 111 865 115 869
rect 815 867 819 871
rect 1111 865 1115 869
rect 211 859 215 863
rect 351 859 355 863
rect 739 859 743 863
rect 111 847 115 851
rect 1111 847 1115 851
rect 135 832 139 836
rect 263 832 267 836
rect 431 832 435 836
rect 623 832 627 836
rect 831 832 835 836
rect 1015 832 1019 836
rect 135 816 139 820
rect 279 816 283 820
rect 463 816 467 820
rect 647 816 651 820
rect 839 816 843 820
rect 1015 816 1019 820
rect 111 801 115 805
rect 1111 801 1115 805
rect 111 783 115 787
rect 219 787 223 791
rect 567 787 571 791
rect 575 787 579 791
rect 1015 791 1019 795
rect 1111 783 1115 787
rect 143 771 147 775
rect 287 771 291 775
rect 471 771 475 775
rect 655 771 659 775
rect 847 771 851 775
rect 1023 771 1027 775
rect 219 763 223 767
rect 567 763 571 767
rect 191 743 195 747
rect 243 743 247 747
rect 395 743 399 747
rect 499 743 503 747
rect 643 743 647 747
rect 887 743 891 747
rect 1015 743 1019 747
rect 183 733 187 737
rect 303 733 307 737
rect 431 733 435 737
rect 567 733 571 737
rect 719 733 723 737
rect 879 733 883 737
rect 1023 733 1027 737
rect 111 721 115 725
rect 243 719 247 723
rect 395 719 399 723
rect 499 719 503 723
rect 643 719 647 723
rect 1111 721 1115 725
rect 111 703 115 707
rect 635 703 639 707
rect 1111 703 1115 707
rect 175 688 179 692
rect 295 688 299 692
rect 423 688 427 692
rect 559 688 563 692
rect 711 688 715 692
rect 871 688 875 692
rect 1015 688 1019 692
rect 343 664 347 668
rect 455 664 459 668
rect 583 664 587 668
rect 719 664 723 668
rect 863 664 867 668
rect 1015 664 1019 668
rect 111 649 115 653
rect 1111 649 1115 653
rect 111 631 115 635
rect 411 635 415 639
rect 531 635 535 639
rect 663 635 667 639
rect 803 635 807 639
rect 811 635 815 639
rect 999 635 1003 639
rect 1111 631 1115 635
rect 351 619 355 623
rect 463 619 467 623
rect 591 619 595 623
rect 727 619 731 623
rect 871 619 875 623
rect 1023 619 1027 623
rect 359 611 363 615
rect 411 611 415 615
rect 531 611 535 615
rect 663 611 667 615
rect 803 611 807 615
rect 551 595 555 599
rect 603 595 607 599
rect 691 595 695 599
rect 779 595 783 599
rect 911 595 915 599
rect 999 595 1003 599
rect 543 585 547 589
rect 631 585 635 589
rect 719 585 723 589
rect 807 585 811 589
rect 903 585 907 589
rect 1007 585 1011 589
rect 111 573 115 577
rect 603 571 607 575
rect 691 571 695 575
rect 779 571 783 575
rect 1111 573 1115 577
rect 887 567 891 571
rect 111 555 115 559
rect 807 555 811 559
rect 991 555 995 559
rect 1111 555 1115 559
rect 535 540 539 544
rect 623 540 627 544
rect 711 540 715 544
rect 799 540 803 544
rect 895 540 899 544
rect 999 540 1003 544
rect 479 520 483 524
rect 567 520 571 524
rect 655 520 659 524
rect 743 520 747 524
rect 831 520 835 524
rect 919 520 923 524
rect 111 505 115 509
rect 911 507 915 511
rect 1111 505 1115 509
rect 111 487 115 491
rect 547 491 551 495
rect 635 491 639 495
rect 727 491 731 495
rect 815 491 819 495
rect 1111 487 1115 491
rect 487 475 491 479
rect 575 475 579 479
rect 663 475 667 479
rect 751 475 755 479
rect 839 475 843 479
rect 927 475 931 479
rect 547 467 551 471
rect 807 467 811 471
rect 919 467 923 471
rect 443 459 447 463
rect 635 459 639 463
rect 727 459 731 463
rect 815 459 819 463
rect 343 451 347 455
rect 495 451 499 455
rect 855 451 859 455
rect 991 451 995 455
rect 271 441 275 445
rect 375 441 379 445
rect 487 441 491 445
rect 599 441 603 445
rect 719 441 723 445
rect 847 441 851 445
rect 983 441 987 445
rect 111 429 115 433
rect 343 427 347 431
rect 443 423 447 427
rect 919 427 923 431
rect 1111 429 1115 433
rect 111 411 115 415
rect 447 411 451 415
rect 667 411 671 415
rect 1111 411 1115 415
rect 263 396 267 400
rect 367 396 371 400
rect 479 396 483 400
rect 591 396 595 400
rect 711 396 715 400
rect 839 396 843 400
rect 975 396 979 400
rect 495 387 499 391
rect 667 387 671 391
rect 135 380 139 384
rect 263 380 267 384
rect 431 380 435 384
rect 607 380 611 384
rect 791 380 795 384
rect 975 380 979 384
rect 111 365 115 369
rect 859 367 863 371
rect 1111 365 1115 369
rect 111 347 115 351
rect 203 351 207 355
rect 531 351 535 355
rect 539 351 543 355
rect 143 335 147 339
rect 271 335 275 339
rect 439 335 443 339
rect 615 335 619 339
rect 799 335 803 339
rect 983 335 987 339
rect 151 327 155 331
rect 279 327 283 331
rect 447 327 451 331
rect 531 327 535 331
rect 791 327 795 331
rect 223 319 227 323
rect 395 319 399 323
rect 679 319 683 323
rect 939 327 943 331
rect 1111 347 1115 351
rect 143 309 147 313
rect 303 309 307 313
rect 487 309 491 313
rect 671 309 675 313
rect 855 309 859 313
rect 1023 309 1027 313
rect 111 297 115 301
rect 223 295 227 299
rect 395 295 399 299
rect 791 295 795 299
rect 1111 297 1115 301
rect 939 291 943 295
rect 111 279 115 283
rect 915 275 919 279
rect 1111 279 1115 283
rect 135 264 139 268
rect 295 264 299 268
rect 479 264 483 268
rect 663 264 667 268
rect 847 264 851 268
rect 1015 264 1019 268
rect 199 244 203 248
rect 343 244 347 248
rect 479 244 483 248
rect 615 244 619 248
rect 751 244 755 248
rect 895 244 899 248
rect 1015 244 1019 248
rect 111 229 115 233
rect 683 231 687 235
rect 1111 229 1115 233
rect 111 211 115 215
rect 267 215 271 219
rect 423 215 427 219
rect 695 215 699 219
rect 1003 215 1007 219
rect 1015 219 1019 223
rect 1111 211 1115 215
rect 207 199 211 203
rect 351 199 355 203
rect 487 199 491 203
rect 623 199 627 203
rect 759 199 763 203
rect 903 199 907 203
rect 1023 199 1027 203
rect 911 191 915 195
rect 1003 191 1007 195
rect 267 183 271 187
rect 423 183 427 187
rect 695 183 699 187
rect 827 183 831 187
rect 291 171 295 175
rect 379 171 383 175
rect 467 171 471 175
rect 555 171 559 175
rect 643 171 647 175
rect 731 171 735 175
rect 819 171 823 175
rect 1003 179 1007 183
rect 1015 171 1019 175
rect 231 161 235 165
rect 319 161 323 165
rect 407 161 411 165
rect 495 161 499 165
rect 583 161 587 165
rect 671 161 675 165
rect 759 161 763 165
rect 847 161 851 165
rect 935 161 939 165
rect 1023 161 1027 165
rect 111 149 115 153
rect 291 147 295 151
rect 379 147 383 151
rect 467 147 471 151
rect 555 147 559 151
rect 643 147 647 151
rect 731 147 735 151
rect 819 147 823 151
rect 1111 149 1115 153
rect 827 143 831 147
rect 1003 143 1007 147
rect 111 131 115 135
rect 1111 131 1115 135
rect 223 116 227 120
rect 311 116 315 120
rect 399 116 403 120
rect 487 116 491 120
rect 575 116 579 120
rect 663 116 667 120
rect 751 116 755 120
rect 839 116 843 120
rect 927 116 931 120
rect 1015 116 1019 120
<< m3 >>
rect 111 1222 115 1223
rect 111 1217 115 1218
rect 135 1222 139 1223
rect 135 1217 139 1218
rect 223 1222 227 1223
rect 223 1217 227 1218
rect 311 1222 315 1223
rect 311 1217 315 1218
rect 399 1222 403 1223
rect 399 1217 403 1218
rect 1111 1222 1115 1223
rect 1111 1217 1115 1218
rect 112 1202 114 1217
rect 134 1216 140 1217
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 222 1216 228 1217
rect 222 1212 223 1216
rect 227 1212 228 1216
rect 222 1211 228 1212
rect 310 1216 316 1217
rect 310 1212 311 1216
rect 315 1212 316 1216
rect 310 1211 316 1212
rect 398 1216 404 1217
rect 398 1212 399 1216
rect 403 1212 404 1216
rect 398 1211 404 1212
rect 1112 1202 1114 1217
rect 110 1201 116 1202
rect 110 1197 111 1201
rect 115 1197 116 1201
rect 110 1196 116 1197
rect 1110 1201 1116 1202
rect 1110 1197 1111 1201
rect 1115 1197 1116 1201
rect 1110 1196 1116 1197
rect 202 1187 208 1188
rect 110 1183 116 1184
rect 110 1179 111 1183
rect 115 1179 116 1183
rect 202 1183 203 1187
rect 207 1183 208 1187
rect 202 1182 208 1183
rect 290 1187 296 1188
rect 290 1183 291 1187
rect 295 1183 296 1187
rect 290 1182 296 1183
rect 378 1187 384 1188
rect 378 1183 379 1187
rect 383 1183 384 1187
rect 378 1182 384 1183
rect 386 1187 392 1188
rect 386 1183 387 1187
rect 391 1183 392 1187
rect 386 1182 392 1183
rect 1110 1183 1116 1184
rect 110 1178 116 1179
rect 112 1159 114 1178
rect 151 1172 155 1173
rect 142 1171 148 1172
rect 142 1167 143 1171
rect 147 1167 148 1171
rect 151 1167 155 1168
rect 142 1166 148 1167
rect 144 1159 146 1166
rect 111 1158 115 1159
rect 111 1153 115 1154
rect 143 1158 147 1159
rect 152 1156 154 1167
rect 204 1164 206 1182
rect 230 1171 236 1172
rect 230 1167 231 1171
rect 235 1167 236 1171
rect 230 1166 236 1167
rect 202 1163 208 1164
rect 202 1159 203 1163
rect 207 1159 208 1163
rect 232 1159 234 1166
rect 292 1164 294 1182
rect 318 1171 324 1172
rect 318 1167 319 1171
rect 323 1167 324 1171
rect 318 1166 324 1167
rect 290 1163 296 1164
rect 290 1159 291 1163
rect 295 1159 296 1163
rect 320 1159 322 1166
rect 380 1164 382 1182
rect 388 1173 390 1182
rect 1110 1179 1111 1183
rect 1115 1179 1116 1183
rect 1110 1178 1116 1179
rect 387 1172 391 1173
rect 387 1167 391 1168
rect 406 1171 412 1172
rect 406 1167 407 1171
rect 411 1167 412 1171
rect 406 1166 412 1167
rect 378 1163 384 1164
rect 378 1159 379 1163
rect 383 1159 384 1163
rect 408 1159 410 1166
rect 1112 1159 1114 1178
rect 202 1158 208 1159
rect 231 1158 235 1159
rect 290 1158 296 1159
rect 319 1158 323 1159
rect 378 1158 384 1159
rect 407 1158 411 1159
rect 143 1153 147 1154
rect 150 1155 156 1156
rect 112 1134 114 1153
rect 144 1146 146 1153
rect 150 1151 151 1155
rect 155 1151 156 1155
rect 150 1150 156 1151
rect 202 1155 208 1156
rect 202 1151 203 1155
rect 207 1151 208 1155
rect 231 1153 235 1154
rect 290 1155 296 1156
rect 202 1150 208 1151
rect 142 1145 148 1146
rect 142 1141 143 1145
rect 147 1141 148 1145
rect 142 1140 148 1141
rect 110 1133 116 1134
rect 110 1129 111 1133
rect 115 1129 116 1133
rect 204 1132 206 1150
rect 232 1146 234 1153
rect 290 1151 291 1155
rect 295 1151 296 1155
rect 319 1153 323 1154
rect 378 1155 384 1156
rect 290 1150 296 1151
rect 230 1145 236 1146
rect 230 1141 231 1145
rect 235 1141 236 1145
rect 230 1140 236 1141
rect 292 1132 294 1150
rect 320 1146 322 1153
rect 378 1151 379 1155
rect 383 1151 384 1155
rect 407 1153 411 1154
rect 1111 1158 1115 1159
rect 1111 1153 1115 1154
rect 378 1150 384 1151
rect 318 1145 324 1146
rect 318 1141 319 1145
rect 323 1141 324 1145
rect 318 1140 324 1141
rect 380 1132 382 1150
rect 408 1146 410 1153
rect 406 1145 412 1146
rect 406 1141 407 1145
rect 411 1141 412 1145
rect 406 1140 412 1141
rect 1112 1134 1114 1153
rect 1110 1133 1116 1134
rect 110 1128 116 1129
rect 202 1131 208 1132
rect 202 1127 203 1131
rect 207 1127 208 1131
rect 202 1126 208 1127
rect 290 1131 296 1132
rect 290 1127 291 1131
rect 295 1127 296 1131
rect 290 1126 296 1127
rect 378 1131 384 1132
rect 378 1127 379 1131
rect 383 1127 384 1131
rect 1110 1129 1111 1133
rect 1115 1129 1116 1133
rect 1110 1128 1116 1129
rect 378 1126 384 1127
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 1110 1115 1116 1116
rect 110 1110 116 1111
rect 382 1111 388 1112
rect 112 1095 114 1110
rect 382 1107 383 1111
rect 387 1107 388 1111
rect 1110 1111 1111 1115
rect 1115 1111 1116 1115
rect 1110 1110 1116 1111
rect 382 1106 388 1107
rect 134 1100 140 1101
rect 134 1096 135 1100
rect 139 1096 140 1100
rect 134 1095 140 1096
rect 222 1100 228 1101
rect 222 1096 223 1100
rect 227 1096 228 1100
rect 222 1095 228 1096
rect 310 1100 316 1101
rect 310 1096 311 1100
rect 315 1096 316 1100
rect 310 1095 316 1096
rect 111 1094 115 1095
rect 111 1089 115 1090
rect 135 1094 139 1095
rect 135 1089 139 1090
rect 223 1094 227 1095
rect 223 1089 227 1090
rect 279 1094 283 1095
rect 279 1089 283 1090
rect 311 1094 315 1095
rect 311 1089 315 1090
rect 367 1094 371 1095
rect 367 1089 371 1090
rect 112 1074 114 1089
rect 278 1088 284 1089
rect 278 1084 279 1088
rect 283 1084 284 1088
rect 278 1083 284 1084
rect 366 1088 372 1089
rect 366 1084 367 1088
rect 371 1084 372 1088
rect 366 1083 372 1084
rect 110 1073 116 1074
rect 110 1069 111 1073
rect 115 1069 116 1073
rect 110 1068 116 1069
rect 110 1055 116 1056
rect 110 1051 111 1055
rect 115 1051 116 1055
rect 110 1050 116 1051
rect 112 1023 114 1050
rect 286 1043 292 1044
rect 286 1039 287 1043
rect 291 1039 292 1043
rect 286 1038 292 1039
rect 374 1043 380 1044
rect 374 1039 375 1043
rect 379 1039 380 1043
rect 374 1038 380 1039
rect 288 1023 290 1038
rect 376 1023 378 1038
rect 384 1028 386 1106
rect 398 1100 404 1101
rect 398 1096 399 1100
rect 403 1096 404 1100
rect 398 1095 404 1096
rect 1112 1095 1114 1110
rect 399 1094 403 1095
rect 399 1089 403 1090
rect 455 1094 459 1095
rect 455 1089 459 1090
rect 543 1094 547 1095
rect 543 1089 547 1090
rect 631 1094 635 1095
rect 631 1089 635 1090
rect 1111 1094 1115 1095
rect 1111 1089 1115 1090
rect 454 1088 460 1089
rect 454 1084 455 1088
rect 459 1084 460 1088
rect 454 1083 460 1084
rect 542 1088 548 1089
rect 542 1084 543 1088
rect 547 1084 548 1088
rect 542 1083 548 1084
rect 630 1088 636 1089
rect 630 1084 631 1088
rect 635 1084 636 1088
rect 630 1083 636 1084
rect 1112 1074 1114 1089
rect 1110 1073 1116 1074
rect 1110 1069 1111 1073
rect 1115 1069 1116 1073
rect 1110 1068 1116 1069
rect 434 1059 440 1060
rect 434 1055 435 1059
rect 439 1055 440 1059
rect 434 1054 440 1055
rect 522 1059 528 1060
rect 522 1055 523 1059
rect 527 1055 528 1059
rect 522 1054 528 1055
rect 610 1059 616 1060
rect 610 1055 611 1059
rect 615 1055 616 1059
rect 610 1054 616 1055
rect 618 1059 624 1060
rect 618 1055 619 1059
rect 623 1055 624 1059
rect 618 1054 624 1055
rect 1110 1055 1116 1056
rect 436 1036 438 1054
rect 462 1043 468 1044
rect 462 1039 463 1043
rect 467 1039 468 1043
rect 462 1038 468 1039
rect 434 1035 440 1036
rect 434 1031 435 1035
rect 439 1031 440 1035
rect 434 1030 440 1031
rect 382 1027 388 1028
rect 382 1023 383 1027
rect 387 1023 388 1027
rect 464 1023 466 1038
rect 524 1036 526 1054
rect 550 1043 556 1044
rect 550 1039 551 1043
rect 555 1039 556 1043
rect 550 1038 556 1039
rect 522 1035 528 1036
rect 522 1031 523 1035
rect 527 1031 528 1035
rect 522 1030 528 1031
rect 552 1023 554 1038
rect 612 1036 614 1054
rect 610 1035 616 1036
rect 610 1031 611 1035
rect 615 1031 616 1035
rect 610 1030 616 1031
rect 620 1028 622 1054
rect 1110 1051 1111 1055
rect 1115 1051 1116 1055
rect 1110 1050 1116 1051
rect 638 1043 644 1044
rect 638 1039 639 1043
rect 643 1039 644 1043
rect 638 1038 644 1039
rect 618 1027 624 1028
rect 618 1023 619 1027
rect 623 1023 624 1027
rect 640 1023 642 1038
rect 1112 1023 1114 1050
rect 111 1022 115 1023
rect 111 1017 115 1018
rect 287 1022 291 1023
rect 287 1017 291 1018
rect 375 1022 379 1023
rect 382 1022 388 1023
rect 463 1022 467 1023
rect 375 1017 379 1018
rect 463 1017 467 1018
rect 519 1022 523 1023
rect 519 1017 523 1018
rect 551 1022 555 1023
rect 607 1022 611 1023
rect 618 1022 624 1023
rect 639 1022 643 1023
rect 551 1017 555 1018
rect 578 1019 584 1020
rect 112 998 114 1017
rect 520 1010 522 1017
rect 578 1015 579 1019
rect 583 1015 584 1019
rect 607 1017 611 1018
rect 703 1022 707 1023
rect 639 1017 643 1018
rect 666 1019 672 1020
rect 578 1014 584 1015
rect 518 1009 524 1010
rect 518 1005 519 1009
rect 523 1005 524 1009
rect 518 1004 524 1005
rect 110 997 116 998
rect 110 993 111 997
rect 115 993 116 997
rect 580 996 582 1014
rect 608 1010 610 1017
rect 666 1015 667 1019
rect 671 1015 672 1019
rect 807 1022 811 1023
rect 703 1017 707 1018
rect 762 1019 768 1020
rect 666 1014 672 1015
rect 606 1009 612 1010
rect 606 1005 607 1009
rect 611 1005 612 1009
rect 606 1004 612 1005
rect 668 996 670 1014
rect 704 1010 706 1017
rect 762 1015 763 1019
rect 767 1015 768 1019
rect 807 1017 811 1018
rect 911 1022 915 1023
rect 1015 1022 1019 1023
rect 911 1017 915 1018
rect 918 1019 924 1020
rect 762 1014 768 1015
rect 702 1009 708 1010
rect 702 1005 703 1009
rect 707 1005 708 1009
rect 702 1004 708 1005
rect 764 996 766 1014
rect 808 1010 810 1017
rect 912 1010 914 1017
rect 918 1015 919 1019
rect 923 1015 924 1019
rect 918 1014 924 1015
rect 970 1019 976 1020
rect 970 1015 971 1019
rect 975 1015 976 1019
rect 1015 1017 1019 1018
rect 1111 1022 1115 1023
rect 1111 1017 1115 1018
rect 970 1014 976 1015
rect 806 1009 812 1010
rect 806 1005 807 1009
rect 811 1005 812 1009
rect 806 1004 812 1005
rect 910 1009 916 1010
rect 910 1005 911 1009
rect 915 1005 916 1009
rect 910 1004 916 1005
rect 110 992 116 993
rect 578 995 584 996
rect 578 991 579 995
rect 583 991 584 995
rect 578 990 584 991
rect 666 995 672 996
rect 666 991 667 995
rect 671 991 672 995
rect 666 990 672 991
rect 762 995 768 996
rect 762 991 763 995
rect 767 991 768 995
rect 762 990 768 991
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 806 979 812 980
rect 806 975 807 979
rect 811 975 812 979
rect 806 974 812 975
rect 112 959 114 974
rect 510 964 516 965
rect 510 960 511 964
rect 515 960 516 964
rect 510 959 516 960
rect 598 964 604 965
rect 598 960 599 964
rect 603 960 604 964
rect 598 959 604 960
rect 694 964 700 965
rect 694 960 695 964
rect 699 960 700 964
rect 694 959 700 960
rect 798 964 804 965
rect 798 960 799 964
rect 803 960 804 964
rect 798 959 804 960
rect 111 958 115 959
rect 111 953 115 954
rect 399 958 403 959
rect 399 953 403 954
rect 487 958 491 959
rect 487 953 491 954
rect 511 958 515 959
rect 511 953 515 954
rect 575 958 579 959
rect 575 953 579 954
rect 599 958 603 959
rect 599 953 603 954
rect 663 958 667 959
rect 663 953 667 954
rect 695 958 699 959
rect 695 953 699 954
rect 751 958 755 959
rect 751 953 755 954
rect 799 958 803 959
rect 799 953 803 954
rect 112 938 114 953
rect 398 952 404 953
rect 398 948 399 952
rect 403 948 404 952
rect 398 947 404 948
rect 486 952 492 953
rect 486 948 487 952
rect 491 948 492 952
rect 486 947 492 948
rect 574 952 580 953
rect 574 948 575 952
rect 579 948 580 952
rect 574 947 580 948
rect 662 952 668 953
rect 662 948 663 952
rect 667 948 668 952
rect 662 947 668 948
rect 750 952 756 953
rect 750 948 751 952
rect 755 948 756 952
rect 750 947 756 948
rect 110 937 116 938
rect 110 933 111 937
rect 115 933 116 937
rect 110 932 116 933
rect 415 924 419 925
rect 643 924 647 925
rect 110 919 116 920
rect 415 919 419 920
rect 466 923 472 924
rect 466 919 467 923
rect 471 919 472 923
rect 110 915 111 919
rect 115 915 116 919
rect 110 914 116 915
rect 112 895 114 914
rect 406 907 412 908
rect 406 903 407 907
rect 411 903 412 907
rect 406 902 412 903
rect 210 899 216 900
rect 210 895 211 899
rect 215 895 216 899
rect 350 899 356 900
rect 350 895 351 899
rect 355 895 356 899
rect 408 895 410 902
rect 416 900 418 919
rect 466 918 472 919
rect 554 923 560 924
rect 554 919 555 923
rect 559 919 560 923
rect 554 918 560 919
rect 642 919 643 924
rect 647 919 648 924
rect 642 918 648 919
rect 468 900 470 918
rect 494 907 500 908
rect 494 903 495 907
rect 499 903 500 907
rect 494 902 500 903
rect 414 899 420 900
rect 414 895 415 899
rect 419 895 420 899
rect 466 899 472 900
rect 466 895 467 899
rect 471 895 472 899
rect 496 895 498 902
rect 556 900 558 918
rect 638 915 644 916
rect 638 911 639 915
rect 643 911 644 915
rect 638 910 644 911
rect 582 907 588 908
rect 582 903 583 907
rect 587 903 588 907
rect 582 902 588 903
rect 554 899 560 900
rect 554 895 555 899
rect 559 895 560 899
rect 584 895 586 902
rect 111 894 115 895
rect 111 889 115 890
rect 143 894 147 895
rect 210 894 216 895
rect 271 894 275 895
rect 350 894 356 895
rect 407 894 411 895
rect 414 894 420 895
rect 439 894 443 895
rect 466 894 472 895
rect 495 894 499 895
rect 554 894 560 895
rect 583 894 587 895
rect 143 889 147 890
rect 112 870 114 889
rect 144 882 146 889
rect 142 881 148 882
rect 142 877 143 881
rect 147 877 148 881
rect 142 876 148 877
rect 110 869 116 870
rect 110 865 111 869
rect 115 865 116 869
rect 110 864 116 865
rect 212 864 214 894
rect 271 889 275 890
rect 272 882 274 889
rect 270 881 276 882
rect 270 877 271 881
rect 275 877 276 881
rect 270 876 276 877
rect 352 864 354 894
rect 407 889 411 890
rect 439 889 443 890
rect 446 891 452 892
rect 440 882 442 889
rect 446 887 447 891
rect 451 887 452 891
rect 495 889 499 890
rect 583 889 587 890
rect 631 894 635 895
rect 640 892 642 910
rect 670 907 676 908
rect 670 903 671 907
rect 675 903 676 907
rect 670 902 676 903
rect 758 907 764 908
rect 758 903 759 907
rect 763 903 764 907
rect 758 902 764 903
rect 672 895 674 902
rect 760 895 762 902
rect 671 894 675 895
rect 631 889 635 890
rect 638 891 644 892
rect 446 886 452 887
rect 438 881 444 882
rect 438 877 439 881
rect 443 877 444 881
rect 448 877 450 886
rect 632 882 634 889
rect 638 887 639 891
rect 643 887 644 891
rect 671 889 675 890
rect 759 894 763 895
rect 808 892 810 974
rect 902 964 908 965
rect 902 960 903 964
rect 907 960 908 964
rect 902 959 908 960
rect 839 958 843 959
rect 839 953 843 954
rect 903 958 907 959
rect 903 953 907 954
rect 838 952 844 953
rect 838 948 839 952
rect 843 948 844 952
rect 838 947 844 948
rect 920 940 922 1014
rect 972 996 974 1014
rect 1016 1010 1018 1017
rect 1014 1009 1020 1010
rect 1014 1005 1015 1009
rect 1019 1005 1020 1009
rect 1014 1004 1020 1005
rect 1112 998 1114 1017
rect 1110 997 1116 998
rect 970 995 976 996
rect 970 991 971 995
rect 975 991 976 995
rect 1110 993 1111 997
rect 1115 993 1116 997
rect 1110 992 1116 993
rect 970 990 976 991
rect 978 979 984 980
rect 978 975 979 979
rect 983 975 984 979
rect 978 974 984 975
rect 1110 979 1116 980
rect 1110 975 1111 979
rect 1115 975 1116 979
rect 1110 974 1116 975
rect 927 958 931 959
rect 927 953 931 954
rect 926 952 932 953
rect 926 948 927 952
rect 931 948 932 952
rect 926 947 932 948
rect 918 939 924 940
rect 918 935 919 939
rect 923 935 924 939
rect 918 934 924 935
rect 818 923 824 924
rect 818 919 819 923
rect 823 919 824 923
rect 818 918 824 919
rect 820 900 822 918
rect 846 907 852 908
rect 846 903 847 907
rect 851 903 852 907
rect 846 902 852 903
rect 934 907 940 908
rect 934 903 935 907
rect 939 903 940 907
rect 934 902 940 903
rect 818 899 824 900
rect 818 895 819 899
rect 823 895 824 899
rect 848 895 850 902
rect 936 895 938 902
rect 818 894 824 895
rect 839 894 843 895
rect 759 889 763 890
rect 806 891 812 892
rect 638 886 644 887
rect 806 887 807 891
rect 811 887 812 891
rect 806 886 812 887
rect 814 891 820 892
rect 814 887 815 891
rect 819 887 820 891
rect 839 889 843 890
rect 847 894 851 895
rect 847 889 851 890
rect 935 894 939 895
rect 980 892 982 974
rect 1006 964 1012 965
rect 1006 960 1007 964
rect 1011 960 1012 964
rect 1006 959 1012 960
rect 1112 959 1114 974
rect 1007 958 1011 959
rect 1007 953 1011 954
rect 1015 958 1019 959
rect 1015 953 1019 954
rect 1111 958 1115 959
rect 1111 953 1115 954
rect 1014 952 1020 953
rect 1014 948 1015 952
rect 1019 948 1020 952
rect 1014 947 1020 948
rect 1112 938 1114 953
rect 1110 937 1116 938
rect 1110 933 1111 937
rect 1115 933 1116 937
rect 1110 932 1116 933
rect 994 923 1000 924
rect 994 919 995 923
rect 999 919 1000 923
rect 994 918 1000 919
rect 1110 919 1116 920
rect 996 900 998 918
rect 1110 915 1111 919
rect 1115 915 1116 919
rect 1110 914 1116 915
rect 1022 907 1028 908
rect 1022 903 1023 907
rect 1027 903 1028 907
rect 1022 902 1028 903
rect 994 899 1000 900
rect 994 895 995 899
rect 999 895 1000 899
rect 1024 895 1026 902
rect 1112 895 1114 914
rect 994 894 1000 895
rect 1023 894 1027 895
rect 935 889 939 890
rect 978 891 984 892
rect 814 886 820 887
rect 630 881 636 882
rect 630 877 631 881
rect 635 877 636 881
rect 438 876 444 877
rect 447 876 451 877
rect 630 876 636 877
rect 739 876 743 877
rect 447 871 451 872
rect 816 872 818 886
rect 840 882 842 889
rect 978 887 979 891
rect 983 887 984 891
rect 1023 889 1027 890
rect 1111 894 1115 895
rect 1111 889 1115 890
rect 978 886 984 887
rect 1024 882 1026 889
rect 838 881 844 882
rect 838 877 839 881
rect 843 877 844 881
rect 838 876 844 877
rect 1022 881 1028 882
rect 1022 877 1023 881
rect 1027 877 1028 881
rect 1022 876 1028 877
rect 739 871 743 872
rect 814 871 820 872
rect 740 864 742 871
rect 814 867 815 871
rect 819 867 820 871
rect 1112 870 1114 889
rect 814 866 820 867
rect 1110 869 1116 870
rect 1110 865 1111 869
rect 1115 865 1116 869
rect 1110 864 1116 865
rect 210 863 216 864
rect 210 859 211 863
rect 215 859 216 863
rect 210 858 216 859
rect 350 863 356 864
rect 350 859 351 863
rect 355 859 356 863
rect 350 858 356 859
rect 738 863 744 864
rect 738 859 739 863
rect 743 859 744 863
rect 738 858 744 859
rect 110 851 116 852
rect 110 847 111 851
rect 115 847 116 851
rect 110 846 116 847
rect 1110 851 1116 852
rect 1110 847 1111 851
rect 1115 847 1116 851
rect 1110 846 1116 847
rect 112 827 114 846
rect 134 836 140 837
rect 134 832 135 836
rect 139 832 140 836
rect 134 831 140 832
rect 262 836 268 837
rect 262 832 263 836
rect 267 832 268 836
rect 262 831 268 832
rect 430 836 436 837
rect 430 832 431 836
rect 435 832 436 836
rect 430 831 436 832
rect 622 836 628 837
rect 622 832 623 836
rect 627 832 628 836
rect 622 831 628 832
rect 830 836 836 837
rect 830 832 831 836
rect 835 832 836 836
rect 830 831 836 832
rect 1014 836 1020 837
rect 1014 832 1015 836
rect 1019 832 1020 836
rect 1014 831 1020 832
rect 136 827 138 831
rect 264 827 266 831
rect 432 827 434 831
rect 624 827 626 831
rect 832 827 834 831
rect 1016 827 1018 831
rect 1112 827 1114 846
rect 111 826 115 827
rect 111 821 115 822
rect 135 826 139 827
rect 135 821 139 822
rect 263 826 267 827
rect 263 821 267 822
rect 279 826 283 827
rect 279 821 283 822
rect 431 826 435 827
rect 431 821 435 822
rect 463 826 467 827
rect 463 821 467 822
rect 623 826 627 827
rect 623 821 627 822
rect 647 826 651 827
rect 647 821 651 822
rect 831 826 835 827
rect 831 821 835 822
rect 839 826 843 827
rect 839 821 843 822
rect 1015 826 1019 827
rect 1015 821 1019 822
rect 1111 826 1115 827
rect 1111 821 1115 822
rect 112 806 114 821
rect 134 820 140 821
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 278 820 284 821
rect 278 816 279 820
rect 283 816 284 820
rect 278 815 284 816
rect 462 820 468 821
rect 462 816 463 820
rect 467 816 468 820
rect 462 815 468 816
rect 646 820 652 821
rect 646 816 647 820
rect 651 816 652 820
rect 646 815 652 816
rect 838 820 844 821
rect 838 816 839 820
rect 843 816 844 820
rect 838 815 844 816
rect 1014 820 1020 821
rect 1014 816 1015 820
rect 1019 816 1020 820
rect 1014 815 1020 816
rect 1112 806 1114 821
rect 110 805 116 806
rect 110 801 111 805
rect 115 801 116 805
rect 110 800 116 801
rect 1110 805 1116 806
rect 1110 801 1111 805
rect 1115 801 1116 805
rect 1110 800 1116 801
rect 1014 795 1020 796
rect 218 791 224 792
rect 191 788 195 789
rect 110 787 116 788
rect 110 783 111 787
rect 115 783 116 787
rect 218 787 219 791
rect 223 787 224 791
rect 218 786 224 787
rect 566 791 572 792
rect 566 787 567 791
rect 571 787 572 791
rect 566 786 572 787
rect 574 791 580 792
rect 574 786 575 791
rect 191 783 195 784
rect 110 782 116 783
rect 112 751 114 782
rect 142 775 148 776
rect 142 771 143 775
rect 147 771 148 775
rect 142 770 148 771
rect 144 751 146 770
rect 111 750 115 751
rect 111 745 115 746
rect 143 750 147 751
rect 143 745 147 746
rect 183 750 187 751
rect 192 748 194 783
rect 220 768 222 786
rect 286 775 292 776
rect 286 771 287 775
rect 291 771 292 775
rect 286 770 292 771
rect 470 775 476 776
rect 470 771 471 775
rect 475 771 476 775
rect 470 770 476 771
rect 218 767 224 768
rect 218 763 219 767
rect 223 763 224 767
rect 218 762 224 763
rect 288 751 290 770
rect 472 751 474 770
rect 568 768 570 786
rect 579 786 580 791
rect 1014 791 1015 795
rect 1019 791 1020 795
rect 1014 790 1020 791
rect 575 783 579 784
rect 654 775 660 776
rect 654 771 655 775
rect 659 771 660 775
rect 654 770 660 771
rect 846 775 852 776
rect 846 771 847 775
rect 851 771 852 775
rect 846 770 852 771
rect 566 767 572 768
rect 566 763 567 767
rect 571 763 572 767
rect 566 762 572 763
rect 656 751 658 770
rect 848 751 850 770
rect 287 750 291 751
rect 183 745 187 746
rect 190 747 196 748
rect 112 726 114 745
rect 184 738 186 745
rect 190 743 191 747
rect 195 743 196 747
rect 190 742 196 743
rect 242 747 248 748
rect 242 743 243 747
rect 247 743 248 747
rect 287 745 291 746
rect 303 750 307 751
rect 431 750 435 751
rect 303 745 307 746
rect 394 747 400 748
rect 242 742 248 743
rect 182 737 188 738
rect 182 733 183 737
rect 187 733 188 737
rect 182 732 188 733
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 244 724 246 742
rect 304 738 306 745
rect 394 743 395 747
rect 399 743 400 747
rect 431 745 435 746
rect 471 750 475 751
rect 567 750 571 751
rect 471 745 475 746
rect 498 747 504 748
rect 394 742 400 743
rect 302 737 308 738
rect 302 733 303 737
rect 307 733 308 737
rect 302 732 308 733
rect 396 724 398 742
rect 432 738 434 745
rect 498 743 499 747
rect 503 743 504 747
rect 655 750 659 751
rect 567 745 571 746
rect 642 747 648 748
rect 498 742 504 743
rect 430 737 436 738
rect 430 733 431 737
rect 435 733 436 737
rect 430 732 436 733
rect 500 724 502 742
rect 568 738 570 745
rect 642 743 643 747
rect 647 743 648 747
rect 655 745 659 746
rect 719 750 723 751
rect 719 745 723 746
rect 847 750 851 751
rect 847 745 851 746
rect 879 750 883 751
rect 1016 748 1018 790
rect 1110 787 1116 788
rect 1110 783 1111 787
rect 1115 783 1116 787
rect 1110 782 1116 783
rect 1022 775 1028 776
rect 1022 771 1023 775
rect 1027 771 1028 775
rect 1022 770 1028 771
rect 1024 751 1026 770
rect 1112 751 1114 782
rect 1023 750 1027 751
rect 879 745 883 746
rect 886 747 892 748
rect 642 742 648 743
rect 566 737 572 738
rect 566 733 567 737
rect 571 733 572 737
rect 566 732 572 733
rect 644 724 646 742
rect 720 738 722 745
rect 880 738 882 745
rect 886 743 887 747
rect 891 743 892 747
rect 886 742 892 743
rect 1014 747 1020 748
rect 1014 743 1015 747
rect 1019 743 1020 747
rect 1023 745 1027 746
rect 1111 750 1115 751
rect 1111 745 1115 746
rect 1014 742 1020 743
rect 718 737 724 738
rect 718 733 719 737
rect 723 733 724 737
rect 718 732 724 733
rect 878 737 884 738
rect 878 733 879 737
rect 883 733 884 737
rect 878 732 884 733
rect 110 720 116 721
rect 242 723 248 724
rect 242 719 243 723
rect 247 719 248 723
rect 242 718 248 719
rect 394 723 400 724
rect 394 719 395 723
rect 399 719 400 723
rect 394 718 400 719
rect 498 723 504 724
rect 498 719 499 723
rect 503 719 504 723
rect 498 718 504 719
rect 642 723 648 724
rect 642 719 643 723
rect 647 719 648 723
rect 642 718 648 719
rect 110 707 116 708
rect 110 703 111 707
rect 115 703 116 707
rect 110 702 116 703
rect 634 707 640 708
rect 634 703 635 707
rect 639 703 640 707
rect 634 702 640 703
rect 112 675 114 702
rect 174 692 180 693
rect 174 688 175 692
rect 179 688 180 692
rect 174 687 180 688
rect 294 692 300 693
rect 294 688 295 692
rect 299 688 300 692
rect 294 687 300 688
rect 422 692 428 693
rect 422 688 423 692
rect 427 688 428 692
rect 422 687 428 688
rect 558 692 564 693
rect 558 688 559 692
rect 563 688 564 692
rect 558 687 564 688
rect 176 675 178 687
rect 296 675 298 687
rect 424 675 426 687
rect 560 675 562 687
rect 111 674 115 675
rect 111 669 115 670
rect 175 674 179 675
rect 175 669 179 670
rect 295 674 299 675
rect 295 669 299 670
rect 343 674 347 675
rect 343 669 347 670
rect 423 674 427 675
rect 423 669 427 670
rect 455 674 459 675
rect 455 669 459 670
rect 559 674 563 675
rect 559 669 563 670
rect 583 674 587 675
rect 583 669 587 670
rect 112 654 114 669
rect 342 668 348 669
rect 342 664 343 668
rect 347 664 348 668
rect 342 663 348 664
rect 454 668 460 669
rect 454 664 455 668
rect 459 664 460 668
rect 454 663 460 664
rect 582 668 588 669
rect 582 664 583 668
rect 587 664 588 668
rect 582 663 588 664
rect 636 661 638 702
rect 710 692 716 693
rect 710 688 711 692
rect 715 688 716 692
rect 710 687 716 688
rect 870 692 876 693
rect 870 688 871 692
rect 875 688 876 692
rect 870 687 876 688
rect 712 675 714 687
rect 872 675 874 687
rect 711 674 715 675
rect 711 669 715 670
rect 719 674 723 675
rect 719 669 723 670
rect 863 674 867 675
rect 863 669 867 670
rect 871 674 875 675
rect 871 669 875 670
rect 718 668 724 669
rect 718 664 719 668
rect 723 664 724 668
rect 718 663 724 664
rect 862 668 868 669
rect 862 664 863 668
rect 867 664 868 668
rect 862 663 868 664
rect 359 660 363 661
rect 359 655 363 656
rect 635 660 639 661
rect 635 655 639 656
rect 110 653 116 654
rect 110 649 111 653
rect 115 649 116 653
rect 110 648 116 649
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 110 630 116 631
rect 112 603 114 630
rect 350 623 356 624
rect 350 619 351 623
rect 355 619 356 623
rect 350 618 356 619
rect 352 603 354 618
rect 360 616 362 655
rect 410 639 416 640
rect 410 635 411 639
rect 415 635 416 639
rect 410 634 416 635
rect 530 639 536 640
rect 530 635 531 639
rect 535 635 536 639
rect 530 634 536 635
rect 662 639 668 640
rect 662 635 663 639
rect 667 635 668 639
rect 662 634 668 635
rect 802 639 808 640
rect 802 635 803 639
rect 807 635 808 639
rect 802 634 808 635
rect 810 639 816 640
rect 810 635 811 639
rect 815 635 816 639
rect 810 634 816 635
rect 412 616 414 634
rect 462 623 468 624
rect 462 619 463 623
rect 467 619 468 623
rect 462 618 468 619
rect 358 615 364 616
rect 358 611 359 615
rect 363 611 364 615
rect 358 610 364 611
rect 410 615 416 616
rect 410 611 411 615
rect 415 611 416 615
rect 410 610 416 611
rect 464 603 466 618
rect 532 616 534 634
rect 590 623 596 624
rect 551 620 555 621
rect 590 619 591 623
rect 595 619 596 623
rect 590 618 596 619
rect 530 615 536 616
rect 551 615 555 616
rect 530 611 531 615
rect 535 611 536 615
rect 530 610 536 611
rect 111 602 115 603
rect 111 597 115 598
rect 351 602 355 603
rect 351 597 355 598
rect 463 602 467 603
rect 463 597 467 598
rect 543 602 547 603
rect 552 600 554 615
rect 592 603 594 618
rect 664 616 666 634
rect 726 623 732 624
rect 726 619 727 623
rect 731 619 732 623
rect 726 618 732 619
rect 662 615 668 616
rect 662 611 663 615
rect 667 611 668 615
rect 662 610 668 611
rect 728 603 730 618
rect 804 616 806 634
rect 812 621 814 634
rect 870 623 876 624
rect 811 620 815 621
rect 870 619 871 623
rect 875 619 876 623
rect 870 618 876 619
rect 802 615 808 616
rect 811 615 815 616
rect 802 611 803 615
rect 807 611 808 615
rect 802 610 808 611
rect 872 603 874 618
rect 591 602 595 603
rect 543 597 547 598
rect 550 599 556 600
rect 112 578 114 597
rect 544 590 546 597
rect 550 595 551 599
rect 555 595 556 599
rect 631 602 635 603
rect 591 597 595 598
rect 602 599 608 600
rect 550 594 556 595
rect 602 595 603 599
rect 607 595 608 599
rect 719 602 723 603
rect 631 597 635 598
rect 690 599 696 600
rect 602 594 608 595
rect 542 589 548 590
rect 542 585 543 589
rect 547 585 548 589
rect 542 584 548 585
rect 110 577 116 578
rect 110 573 111 577
rect 115 573 116 577
rect 604 576 606 594
rect 632 590 634 597
rect 690 595 691 599
rect 695 595 696 599
rect 719 597 723 598
rect 727 602 731 603
rect 807 602 811 603
rect 727 597 731 598
rect 778 599 784 600
rect 690 594 696 595
rect 630 589 636 590
rect 630 585 631 589
rect 635 585 636 589
rect 630 584 636 585
rect 692 576 694 594
rect 720 590 722 597
rect 778 595 779 599
rect 783 595 784 599
rect 807 597 811 598
rect 871 602 875 603
rect 871 597 875 598
rect 778 594 784 595
rect 718 589 724 590
rect 718 585 719 589
rect 723 585 724 589
rect 718 584 724 585
rect 780 576 782 594
rect 808 590 810 597
rect 806 589 812 590
rect 806 585 807 589
rect 811 585 812 589
rect 806 584 812 585
rect 110 572 116 573
rect 602 575 608 576
rect 602 571 603 575
rect 607 571 608 575
rect 602 570 608 571
rect 690 575 696 576
rect 690 571 691 575
rect 695 571 696 575
rect 690 570 696 571
rect 778 575 784 576
rect 778 571 779 575
rect 783 571 784 575
rect 888 572 890 742
rect 1024 738 1026 745
rect 1022 737 1028 738
rect 1022 733 1023 737
rect 1027 733 1028 737
rect 1022 732 1028 733
rect 1112 726 1114 745
rect 1110 725 1116 726
rect 1110 721 1111 725
rect 1115 721 1116 725
rect 1110 720 1116 721
rect 1110 707 1116 708
rect 1110 703 1111 707
rect 1115 703 1116 707
rect 1110 702 1116 703
rect 1014 692 1020 693
rect 1014 688 1015 692
rect 1019 688 1020 692
rect 1014 687 1020 688
rect 1016 675 1018 687
rect 1112 675 1114 702
rect 1015 674 1019 675
rect 1015 669 1019 670
rect 1111 674 1115 675
rect 1111 669 1115 670
rect 1014 668 1020 669
rect 1014 664 1015 668
rect 1019 664 1020 668
rect 1014 663 1020 664
rect 1112 654 1114 669
rect 1110 653 1116 654
rect 1110 649 1111 653
rect 1115 649 1116 653
rect 1110 648 1116 649
rect 998 639 1004 640
rect 998 635 999 639
rect 1003 635 1004 639
rect 998 634 1004 635
rect 1110 635 1116 636
rect 903 602 907 603
rect 1000 600 1002 634
rect 1110 631 1111 635
rect 1115 631 1116 635
rect 1110 630 1116 631
rect 1022 623 1028 624
rect 1022 619 1023 623
rect 1027 619 1028 623
rect 1022 618 1028 619
rect 1024 603 1026 618
rect 1112 603 1114 630
rect 1007 602 1011 603
rect 903 597 907 598
rect 910 599 916 600
rect 904 590 906 597
rect 910 595 911 599
rect 915 595 916 599
rect 910 594 916 595
rect 998 599 1004 600
rect 998 595 999 599
rect 1003 595 1004 599
rect 1007 597 1011 598
rect 1023 602 1027 603
rect 1023 597 1027 598
rect 1111 602 1115 603
rect 1111 597 1115 598
rect 998 594 1004 595
rect 902 589 908 590
rect 902 585 903 589
rect 907 585 908 589
rect 902 584 908 585
rect 778 570 784 571
rect 886 571 892 572
rect 886 567 887 571
rect 891 567 892 571
rect 886 566 892 567
rect 110 559 116 560
rect 110 555 111 559
rect 115 555 116 559
rect 110 554 116 555
rect 806 559 812 560
rect 806 555 807 559
rect 811 555 812 559
rect 806 554 812 555
rect 112 531 114 554
rect 534 544 540 545
rect 534 540 535 544
rect 539 540 540 544
rect 534 539 540 540
rect 622 544 628 545
rect 622 540 623 544
rect 627 540 628 544
rect 622 539 628 540
rect 710 544 716 545
rect 710 540 711 544
rect 715 540 716 544
rect 710 539 716 540
rect 798 544 804 545
rect 798 540 799 544
rect 803 540 804 544
rect 798 539 804 540
rect 536 531 538 539
rect 624 531 626 539
rect 712 531 714 539
rect 800 531 802 539
rect 111 530 115 531
rect 111 525 115 526
rect 479 530 483 531
rect 479 525 483 526
rect 535 530 539 531
rect 535 525 539 526
rect 567 530 571 531
rect 567 525 571 526
rect 623 530 627 531
rect 623 525 627 526
rect 655 530 659 531
rect 655 525 659 526
rect 711 530 715 531
rect 711 525 715 526
rect 743 530 747 531
rect 743 525 747 526
rect 799 530 803 531
rect 799 525 803 526
rect 112 510 114 525
rect 478 524 484 525
rect 478 520 479 524
rect 483 520 484 524
rect 478 519 484 520
rect 566 524 572 525
rect 566 520 567 524
rect 571 520 572 524
rect 566 519 572 520
rect 654 524 660 525
rect 654 520 655 524
rect 659 520 660 524
rect 654 519 660 520
rect 742 524 748 525
rect 742 520 743 524
rect 747 520 748 524
rect 742 519 748 520
rect 110 509 116 510
rect 110 505 111 509
rect 115 505 116 509
rect 110 504 116 505
rect 546 495 552 496
rect 110 491 116 492
rect 110 487 111 491
rect 115 487 116 491
rect 546 491 547 495
rect 551 491 552 495
rect 546 490 552 491
rect 634 495 640 496
rect 634 491 635 495
rect 639 491 640 495
rect 634 490 640 491
rect 726 495 732 496
rect 726 491 727 495
rect 731 491 732 495
rect 726 490 732 491
rect 110 486 116 487
rect 112 459 114 486
rect 486 479 492 480
rect 486 475 487 479
rect 491 475 492 479
rect 486 474 492 475
rect 442 463 448 464
rect 442 459 443 463
rect 447 459 448 463
rect 488 459 490 474
rect 548 472 550 490
rect 574 479 580 480
rect 574 475 575 479
rect 579 475 580 479
rect 574 474 580 475
rect 546 471 552 472
rect 546 467 547 471
rect 551 467 552 471
rect 546 466 552 467
rect 576 459 578 474
rect 636 464 638 490
rect 662 479 668 480
rect 662 475 663 479
rect 667 475 668 479
rect 662 474 668 475
rect 634 463 640 464
rect 634 459 635 463
rect 639 459 640 463
rect 664 459 666 474
rect 728 464 730 490
rect 750 479 756 480
rect 750 475 751 479
rect 755 475 756 479
rect 750 474 756 475
rect 726 463 732 464
rect 726 459 727 463
rect 731 459 732 463
rect 752 459 754 474
rect 808 472 810 554
rect 894 544 900 545
rect 894 540 895 544
rect 899 540 900 544
rect 894 539 900 540
rect 896 531 898 539
rect 831 530 835 531
rect 831 525 835 526
rect 895 530 899 531
rect 895 525 899 526
rect 830 524 836 525
rect 830 520 831 524
rect 835 520 836 524
rect 830 519 836 520
rect 912 512 914 594
rect 1008 590 1010 597
rect 1006 589 1012 590
rect 1006 585 1007 589
rect 1011 585 1012 589
rect 1006 584 1012 585
rect 1112 578 1114 597
rect 1110 577 1116 578
rect 1110 573 1111 577
rect 1115 573 1116 577
rect 1110 572 1116 573
rect 990 559 996 560
rect 990 555 991 559
rect 995 555 996 559
rect 990 554 996 555
rect 1110 559 1116 560
rect 1110 555 1111 559
rect 1115 555 1116 559
rect 1110 554 1116 555
rect 919 530 923 531
rect 919 525 923 526
rect 918 524 924 525
rect 918 520 919 524
rect 923 520 924 524
rect 918 519 924 520
rect 910 511 916 512
rect 910 507 911 511
rect 915 507 916 511
rect 910 506 916 507
rect 814 495 820 496
rect 814 491 815 495
rect 819 491 820 495
rect 814 490 820 491
rect 806 471 812 472
rect 806 467 807 471
rect 811 467 812 471
rect 806 466 812 467
rect 816 464 818 490
rect 838 479 844 480
rect 838 475 839 479
rect 843 475 844 479
rect 838 474 844 475
rect 926 479 932 480
rect 926 475 927 479
rect 931 475 932 479
rect 926 474 932 475
rect 814 463 820 464
rect 814 459 815 463
rect 819 459 820 463
rect 840 459 842 474
rect 918 471 924 472
rect 918 467 919 471
rect 923 467 924 471
rect 918 466 924 467
rect 111 458 115 459
rect 111 453 115 454
rect 271 458 275 459
rect 375 458 379 459
rect 442 458 448 459
rect 487 458 491 459
rect 271 453 275 454
rect 342 455 348 456
rect 112 434 114 453
rect 272 446 274 453
rect 342 451 343 455
rect 347 451 348 455
rect 375 453 379 454
rect 342 450 348 451
rect 270 445 276 446
rect 270 441 271 445
rect 275 441 276 445
rect 270 440 276 441
rect 110 433 116 434
rect 110 429 111 433
rect 115 429 116 433
rect 344 432 346 450
rect 376 446 378 453
rect 374 445 380 446
rect 374 441 375 445
rect 379 441 380 445
rect 374 440 380 441
rect 110 428 116 429
rect 342 431 348 432
rect 342 427 343 431
rect 347 427 348 431
rect 444 428 446 458
rect 575 458 579 459
rect 487 453 491 454
rect 494 455 500 456
rect 488 446 490 453
rect 494 451 495 455
rect 499 451 500 455
rect 575 453 579 454
rect 599 458 603 459
rect 634 458 640 459
rect 663 458 667 459
rect 599 453 603 454
rect 663 453 667 454
rect 719 458 723 459
rect 726 458 732 459
rect 751 458 755 459
rect 814 458 820 459
rect 839 458 843 459
rect 719 453 723 454
rect 751 453 755 454
rect 839 453 843 454
rect 847 458 851 459
rect 847 453 851 454
rect 854 455 860 456
rect 494 450 500 451
rect 486 445 492 446
rect 486 441 487 445
rect 491 441 492 445
rect 486 440 492 441
rect 342 426 348 427
rect 442 427 448 428
rect 442 423 443 427
rect 447 423 448 427
rect 442 422 448 423
rect 110 415 116 416
rect 110 411 111 415
rect 115 411 116 415
rect 110 410 116 411
rect 446 415 452 416
rect 446 411 447 415
rect 451 411 452 415
rect 446 410 452 411
rect 112 391 114 410
rect 262 400 268 401
rect 262 396 263 400
rect 267 396 268 400
rect 262 395 268 396
rect 366 400 372 401
rect 366 396 367 400
rect 371 396 372 400
rect 366 395 372 396
rect 264 391 266 395
rect 368 391 370 395
rect 111 390 115 391
rect 111 385 115 386
rect 135 390 139 391
rect 135 385 139 386
rect 263 390 267 391
rect 263 385 267 386
rect 367 390 371 391
rect 367 385 371 386
rect 431 390 435 391
rect 431 385 435 386
rect 112 370 114 385
rect 134 384 140 385
rect 134 380 135 384
rect 139 380 140 384
rect 134 379 140 380
rect 262 384 268 385
rect 262 380 263 384
rect 267 380 268 384
rect 262 379 268 380
rect 430 384 436 385
rect 430 380 431 384
rect 435 380 436 384
rect 430 379 436 380
rect 110 369 116 370
rect 110 365 111 369
rect 115 365 116 369
rect 110 364 116 365
rect 202 355 208 356
rect 110 351 116 352
rect 110 347 111 351
rect 115 347 116 351
rect 202 351 203 355
rect 207 351 208 355
rect 202 350 208 351
rect 110 346 116 347
rect 112 327 114 346
rect 204 341 206 350
rect 151 340 155 341
rect 142 339 148 340
rect 142 335 143 339
rect 147 335 148 339
rect 151 335 155 336
rect 203 340 207 341
rect 279 340 283 341
rect 203 335 207 336
rect 270 339 276 340
rect 270 335 271 339
rect 275 335 276 339
rect 279 335 283 336
rect 438 339 444 340
rect 438 335 439 339
rect 443 335 444 339
rect 142 334 148 335
rect 144 327 146 334
rect 152 332 154 335
rect 270 334 276 335
rect 150 331 156 332
rect 150 327 151 331
rect 155 327 156 331
rect 272 327 274 334
rect 280 332 282 335
rect 438 334 444 335
rect 278 331 284 332
rect 278 327 279 331
rect 283 327 284 331
rect 440 327 442 334
rect 448 332 450 410
rect 478 400 484 401
rect 478 396 479 400
rect 483 396 484 400
rect 478 395 484 396
rect 480 391 482 395
rect 496 392 498 450
rect 600 446 602 453
rect 720 446 722 453
rect 848 446 850 453
rect 854 451 855 455
rect 859 451 860 455
rect 854 450 862 451
rect 856 449 862 450
rect 598 445 604 446
rect 598 441 599 445
rect 603 441 604 445
rect 598 440 604 441
rect 718 445 724 446
rect 718 441 719 445
rect 723 441 724 445
rect 718 440 724 441
rect 846 445 852 446
rect 846 441 847 445
rect 851 441 852 445
rect 846 440 852 441
rect 666 415 672 416
rect 666 411 667 415
rect 671 411 672 415
rect 666 410 672 411
rect 590 400 596 401
rect 590 396 591 400
rect 595 396 596 400
rect 590 395 596 396
rect 494 391 500 392
rect 592 391 594 395
rect 668 392 670 410
rect 710 400 716 401
rect 710 396 711 400
rect 715 396 716 400
rect 710 395 716 396
rect 838 400 844 401
rect 838 396 839 400
rect 843 396 844 400
rect 838 395 844 396
rect 666 391 672 392
rect 712 391 714 395
rect 840 391 842 395
rect 479 390 483 391
rect 494 387 495 391
rect 499 387 500 391
rect 494 386 500 387
rect 591 390 595 391
rect 479 385 483 386
rect 591 385 595 386
rect 607 390 611 391
rect 666 387 667 391
rect 671 387 672 391
rect 666 386 672 387
rect 711 390 715 391
rect 607 385 611 386
rect 711 385 715 386
rect 791 390 795 391
rect 791 385 795 386
rect 839 390 843 391
rect 839 385 843 386
rect 606 384 612 385
rect 606 380 607 384
rect 611 380 612 384
rect 606 379 612 380
rect 790 384 796 385
rect 790 380 791 384
rect 795 380 796 384
rect 790 379 796 380
rect 860 372 862 449
rect 920 432 922 466
rect 928 459 930 474
rect 927 458 931 459
rect 927 453 931 454
rect 983 458 987 459
rect 992 456 994 554
rect 998 544 1004 545
rect 998 540 999 544
rect 1003 540 1004 544
rect 998 539 1004 540
rect 1000 531 1002 539
rect 1112 531 1114 554
rect 999 530 1003 531
rect 999 525 1003 526
rect 1111 530 1115 531
rect 1111 525 1115 526
rect 1112 510 1114 525
rect 1110 509 1116 510
rect 1110 505 1111 509
rect 1115 505 1116 509
rect 1110 504 1116 505
rect 1110 491 1116 492
rect 1110 487 1111 491
rect 1115 487 1116 491
rect 1110 486 1116 487
rect 1112 459 1114 486
rect 1111 458 1115 459
rect 983 453 987 454
rect 990 455 996 456
rect 984 446 986 453
rect 990 451 991 455
rect 995 451 996 455
rect 1111 453 1115 454
rect 990 450 996 451
rect 982 445 988 446
rect 982 441 983 445
rect 987 441 988 445
rect 982 440 988 441
rect 1112 434 1114 453
rect 1110 433 1116 434
rect 918 431 924 432
rect 918 427 919 431
rect 923 427 924 431
rect 1110 429 1111 433
rect 1115 429 1116 433
rect 1110 428 1116 429
rect 918 426 924 427
rect 1110 415 1116 416
rect 1110 411 1111 415
rect 1115 411 1116 415
rect 1110 410 1116 411
rect 974 400 980 401
rect 974 396 975 400
rect 979 396 980 400
rect 974 395 980 396
rect 976 391 978 395
rect 1112 391 1114 410
rect 975 390 979 391
rect 975 385 979 386
rect 1111 390 1115 391
rect 1111 385 1115 386
rect 974 384 980 385
rect 974 380 975 384
rect 979 380 980 384
rect 974 379 980 380
rect 858 371 864 372
rect 858 367 859 371
rect 863 367 864 371
rect 1112 370 1114 385
rect 858 366 864 367
rect 1110 369 1116 370
rect 1110 365 1111 369
rect 1115 365 1116 369
rect 1110 364 1116 365
rect 530 355 536 356
rect 530 351 531 355
rect 535 351 536 355
rect 530 350 536 351
rect 538 355 544 356
rect 538 351 539 355
rect 543 351 544 355
rect 538 350 544 351
rect 1110 351 1116 352
rect 532 332 534 350
rect 540 341 542 350
rect 1110 347 1111 351
rect 1115 347 1116 351
rect 1110 346 1116 347
rect 539 340 543 341
rect 539 335 543 336
rect 614 339 620 340
rect 614 335 615 339
rect 619 335 620 339
rect 614 334 620 335
rect 798 339 804 340
rect 798 335 799 339
rect 803 335 804 339
rect 798 334 804 335
rect 982 339 988 340
rect 982 335 983 339
rect 987 335 988 339
rect 982 334 988 335
rect 446 331 452 332
rect 446 327 447 331
rect 451 327 452 331
rect 530 331 536 332
rect 530 327 531 331
rect 535 327 536 331
rect 616 327 618 334
rect 790 331 796 332
rect 790 327 791 331
rect 795 327 796 331
rect 800 327 802 334
rect 938 331 944 332
rect 938 327 939 331
rect 943 327 944 331
rect 984 327 986 334
rect 1112 327 1114 346
rect 111 326 115 327
rect 111 321 115 322
rect 143 326 147 327
rect 150 326 156 327
rect 271 326 275 327
rect 278 326 284 327
rect 303 326 307 327
rect 143 321 147 322
rect 222 323 228 324
rect 112 302 114 321
rect 144 314 146 321
rect 222 319 223 323
rect 227 319 228 323
rect 271 321 275 322
rect 439 326 443 327
rect 446 326 452 327
rect 487 326 491 327
rect 530 326 536 327
rect 615 326 619 327
rect 303 321 307 322
rect 394 323 400 324
rect 222 318 228 319
rect 142 313 148 314
rect 142 309 143 313
rect 147 309 148 313
rect 142 308 148 309
rect 110 301 116 302
rect 110 297 111 301
rect 115 297 116 301
rect 224 300 226 318
rect 304 314 306 321
rect 394 319 395 323
rect 399 319 400 323
rect 439 321 443 322
rect 487 321 491 322
rect 615 321 619 322
rect 671 326 675 327
rect 790 326 796 327
rect 799 326 803 327
rect 671 321 675 322
rect 678 323 684 324
rect 394 318 400 319
rect 302 313 308 314
rect 302 309 303 313
rect 307 309 308 313
rect 302 308 308 309
rect 396 300 398 318
rect 488 314 490 321
rect 672 314 674 321
rect 678 319 679 323
rect 683 319 684 323
rect 678 318 684 319
rect 486 313 492 314
rect 486 309 487 313
rect 491 309 492 313
rect 486 308 492 309
rect 670 313 676 314
rect 670 309 671 313
rect 675 309 676 313
rect 680 313 682 318
rect 680 311 686 313
rect 670 308 676 309
rect 110 296 116 297
rect 222 299 228 300
rect 222 295 223 299
rect 227 295 228 299
rect 222 294 228 295
rect 394 299 400 300
rect 394 295 395 299
rect 399 295 400 299
rect 394 294 400 295
rect 110 283 116 284
rect 110 279 111 283
rect 115 279 116 283
rect 110 278 116 279
rect 112 255 114 278
rect 134 268 140 269
rect 134 264 135 268
rect 139 264 140 268
rect 134 263 140 264
rect 294 268 300 269
rect 294 264 295 268
rect 299 264 300 268
rect 294 263 300 264
rect 478 268 484 269
rect 478 264 479 268
rect 483 264 484 268
rect 478 263 484 264
rect 662 268 668 269
rect 662 264 663 268
rect 667 264 668 268
rect 662 263 668 264
rect 136 255 138 263
rect 296 255 298 263
rect 480 255 482 263
rect 664 255 666 263
rect 111 254 115 255
rect 111 249 115 250
rect 135 254 139 255
rect 135 249 139 250
rect 199 254 203 255
rect 199 249 203 250
rect 295 254 299 255
rect 295 249 299 250
rect 343 254 347 255
rect 343 249 347 250
rect 479 254 483 255
rect 479 249 483 250
rect 615 254 619 255
rect 615 249 619 250
rect 663 254 667 255
rect 663 249 667 250
rect 112 234 114 249
rect 198 248 204 249
rect 198 244 199 248
rect 203 244 204 248
rect 198 243 204 244
rect 342 248 348 249
rect 342 244 343 248
rect 347 244 348 248
rect 342 243 348 244
rect 478 248 484 249
rect 478 244 479 248
rect 483 244 484 248
rect 478 243 484 244
rect 614 248 620 249
rect 614 244 615 248
rect 619 244 620 248
rect 614 243 620 244
rect 684 236 686 311
rect 792 300 794 326
rect 799 321 803 322
rect 855 326 859 327
rect 938 326 944 327
rect 983 326 987 327
rect 855 321 859 322
rect 856 314 858 321
rect 854 313 860 314
rect 854 309 855 313
rect 859 309 860 313
rect 854 308 860 309
rect 790 299 796 300
rect 790 295 791 299
rect 795 295 796 299
rect 940 296 942 326
rect 983 321 987 322
rect 1023 326 1027 327
rect 1023 321 1027 322
rect 1111 326 1115 327
rect 1111 321 1115 322
rect 1024 314 1026 321
rect 1022 313 1028 314
rect 1022 309 1023 313
rect 1027 309 1028 313
rect 1022 308 1028 309
rect 1112 302 1114 321
rect 1110 301 1116 302
rect 1110 297 1111 301
rect 1115 297 1116 301
rect 1110 296 1116 297
rect 790 294 796 295
rect 938 295 944 296
rect 938 291 939 295
rect 943 291 944 295
rect 938 290 944 291
rect 1110 283 1116 284
rect 914 279 920 280
rect 914 275 915 279
rect 919 275 920 279
rect 1110 279 1111 283
rect 1115 279 1116 283
rect 1110 278 1116 279
rect 914 274 920 275
rect 846 268 852 269
rect 846 264 847 268
rect 851 264 852 268
rect 846 263 852 264
rect 848 255 850 263
rect 751 254 755 255
rect 751 249 755 250
rect 847 254 851 255
rect 847 249 851 250
rect 895 254 899 255
rect 895 249 899 250
rect 750 248 756 249
rect 750 244 751 248
rect 755 244 756 248
rect 750 243 756 244
rect 894 248 900 249
rect 894 244 895 248
rect 899 244 900 248
rect 894 243 900 244
rect 682 235 688 236
rect 110 233 116 234
rect 110 229 111 233
rect 115 229 116 233
rect 682 231 683 235
rect 687 231 688 235
rect 682 230 688 231
rect 110 228 116 229
rect 266 219 272 220
rect 110 215 116 216
rect 110 211 111 215
rect 115 211 116 215
rect 266 215 267 219
rect 271 215 272 219
rect 266 214 272 215
rect 422 219 428 220
rect 422 215 423 219
rect 427 215 428 219
rect 422 214 428 215
rect 694 219 700 220
rect 694 215 695 219
rect 699 215 700 219
rect 694 214 700 215
rect 110 210 116 211
rect 112 179 114 210
rect 206 203 212 204
rect 206 199 207 203
rect 211 199 212 203
rect 206 198 212 199
rect 208 179 210 198
rect 268 188 270 214
rect 350 203 356 204
rect 350 199 351 203
rect 355 199 356 203
rect 350 198 356 199
rect 266 187 272 188
rect 266 183 267 187
rect 271 183 272 187
rect 266 182 272 183
rect 352 179 354 198
rect 424 188 426 214
rect 486 203 492 204
rect 486 199 487 203
rect 491 199 492 203
rect 486 198 492 199
rect 622 203 628 204
rect 622 199 623 203
rect 627 199 628 203
rect 622 198 628 199
rect 422 187 428 188
rect 422 183 423 187
rect 427 183 428 187
rect 422 182 428 183
rect 488 179 490 198
rect 624 179 626 198
rect 696 188 698 214
rect 758 203 764 204
rect 758 199 759 203
rect 763 199 764 203
rect 758 198 764 199
rect 902 203 908 204
rect 916 203 918 274
rect 1014 268 1020 269
rect 1014 264 1015 268
rect 1019 264 1020 268
rect 1014 263 1020 264
rect 1016 255 1018 263
rect 1112 255 1114 278
rect 1015 254 1019 255
rect 1015 249 1019 250
rect 1111 254 1115 255
rect 1111 249 1115 250
rect 1014 248 1020 249
rect 1014 244 1015 248
rect 1019 244 1020 248
rect 1014 243 1020 244
rect 1112 234 1114 249
rect 1110 233 1116 234
rect 1110 229 1111 233
rect 1115 229 1116 233
rect 1110 228 1116 229
rect 1014 223 1020 224
rect 1002 219 1008 220
rect 1002 215 1003 219
rect 1007 215 1008 219
rect 1014 219 1015 223
rect 1019 219 1020 223
rect 1014 218 1020 219
rect 1002 214 1008 215
rect 902 199 903 203
rect 907 199 908 203
rect 902 198 908 199
rect 912 201 918 203
rect 694 187 700 188
rect 694 183 695 187
rect 699 183 700 187
rect 694 182 700 183
rect 760 179 762 198
rect 826 187 832 188
rect 826 183 827 187
rect 831 183 832 187
rect 826 182 832 183
rect 111 178 115 179
rect 111 173 115 174
rect 207 178 211 179
rect 207 173 211 174
rect 231 178 235 179
rect 319 178 323 179
rect 231 173 235 174
rect 290 175 296 176
rect 112 154 114 173
rect 232 166 234 173
rect 290 171 291 175
rect 295 171 296 175
rect 319 173 323 174
rect 351 178 355 179
rect 407 178 411 179
rect 351 173 355 174
rect 378 175 384 176
rect 290 170 296 171
rect 230 165 236 166
rect 230 161 231 165
rect 235 161 236 165
rect 230 160 236 161
rect 110 153 116 154
rect 110 149 111 153
rect 115 149 116 153
rect 292 152 294 170
rect 320 166 322 173
rect 378 171 379 175
rect 383 171 384 175
rect 487 178 491 179
rect 407 173 411 174
rect 466 175 472 176
rect 378 170 384 171
rect 318 165 324 166
rect 318 161 319 165
rect 323 161 324 165
rect 318 160 324 161
rect 380 152 382 170
rect 408 166 410 173
rect 466 171 467 175
rect 471 171 472 175
rect 487 173 491 174
rect 495 178 499 179
rect 583 178 587 179
rect 495 173 499 174
rect 554 175 560 176
rect 466 170 472 171
rect 406 165 412 166
rect 406 161 407 165
rect 411 161 412 165
rect 406 160 412 161
rect 468 152 470 170
rect 496 166 498 173
rect 554 171 555 175
rect 559 171 560 175
rect 583 173 587 174
rect 623 178 627 179
rect 671 178 675 179
rect 623 173 627 174
rect 642 175 648 176
rect 554 170 560 171
rect 494 165 500 166
rect 494 161 495 165
rect 499 161 500 165
rect 494 160 500 161
rect 556 152 558 170
rect 584 166 586 173
rect 642 171 643 175
rect 647 171 648 175
rect 759 178 763 179
rect 671 173 675 174
rect 730 175 736 176
rect 642 170 648 171
rect 582 165 588 166
rect 582 161 583 165
rect 587 161 588 165
rect 582 160 588 161
rect 644 152 646 170
rect 672 166 674 173
rect 730 171 731 175
rect 735 171 736 175
rect 759 173 763 174
rect 818 175 824 176
rect 730 170 736 171
rect 670 165 676 166
rect 670 161 671 165
rect 675 161 676 165
rect 670 160 676 161
rect 732 152 734 170
rect 760 166 762 173
rect 818 171 819 175
rect 823 171 824 175
rect 818 170 824 171
rect 758 165 764 166
rect 758 161 759 165
rect 763 161 764 165
rect 758 160 764 161
rect 820 152 822 170
rect 110 148 116 149
rect 290 151 296 152
rect 290 147 291 151
rect 295 147 296 151
rect 290 146 296 147
rect 378 151 384 152
rect 378 147 379 151
rect 383 147 384 151
rect 378 146 384 147
rect 466 151 472 152
rect 466 147 467 151
rect 471 147 472 151
rect 466 146 472 147
rect 554 151 560 152
rect 554 147 555 151
rect 559 147 560 151
rect 554 146 560 147
rect 642 151 648 152
rect 642 147 643 151
rect 647 147 648 151
rect 642 146 648 147
rect 730 151 736 152
rect 730 147 731 151
rect 735 147 736 151
rect 730 146 736 147
rect 818 151 824 152
rect 818 147 819 151
rect 823 147 824 151
rect 828 148 830 182
rect 904 179 906 198
rect 912 196 914 201
rect 1004 196 1006 214
rect 910 195 916 196
rect 910 191 911 195
rect 915 191 916 195
rect 910 190 916 191
rect 1002 195 1008 196
rect 1002 191 1003 195
rect 1007 191 1008 195
rect 1002 190 1008 191
rect 1002 183 1008 184
rect 1002 179 1003 183
rect 1007 179 1008 183
rect 847 178 851 179
rect 847 173 851 174
rect 903 178 907 179
rect 903 173 907 174
rect 935 178 939 179
rect 1002 178 1008 179
rect 935 173 939 174
rect 848 166 850 173
rect 936 166 938 173
rect 846 165 852 166
rect 846 161 847 165
rect 851 161 852 165
rect 846 160 852 161
rect 934 165 940 166
rect 934 161 935 165
rect 939 161 940 165
rect 934 160 940 161
rect 1004 148 1006 178
rect 1016 176 1018 218
rect 1110 215 1116 216
rect 1110 211 1111 215
rect 1115 211 1116 215
rect 1110 210 1116 211
rect 1022 203 1028 204
rect 1022 199 1023 203
rect 1027 199 1028 203
rect 1022 198 1028 199
rect 1024 179 1026 198
rect 1112 179 1114 210
rect 1023 178 1027 179
rect 1014 175 1020 176
rect 1014 171 1015 175
rect 1019 171 1020 175
rect 1023 173 1027 174
rect 1111 178 1115 179
rect 1111 173 1115 174
rect 1014 170 1020 171
rect 1024 166 1026 173
rect 1022 165 1028 166
rect 1022 161 1023 165
rect 1027 161 1028 165
rect 1022 160 1028 161
rect 1112 154 1114 173
rect 1110 153 1116 154
rect 1110 149 1111 153
rect 1115 149 1116 153
rect 1110 148 1116 149
rect 818 146 824 147
rect 826 147 832 148
rect 826 143 827 147
rect 831 143 832 147
rect 826 142 832 143
rect 1002 147 1008 148
rect 1002 143 1003 147
rect 1007 143 1008 147
rect 1002 142 1008 143
rect 110 135 116 136
rect 110 131 111 135
rect 115 131 116 135
rect 110 130 116 131
rect 1110 135 1116 136
rect 1110 131 1111 135
rect 1115 131 1116 135
rect 1110 130 1116 131
rect 112 115 114 130
rect 222 120 228 121
rect 222 116 223 120
rect 227 116 228 120
rect 222 115 228 116
rect 310 120 316 121
rect 310 116 311 120
rect 315 116 316 120
rect 310 115 316 116
rect 398 120 404 121
rect 398 116 399 120
rect 403 116 404 120
rect 398 115 404 116
rect 486 120 492 121
rect 486 116 487 120
rect 491 116 492 120
rect 486 115 492 116
rect 574 120 580 121
rect 574 116 575 120
rect 579 116 580 120
rect 574 115 580 116
rect 662 120 668 121
rect 662 116 663 120
rect 667 116 668 120
rect 662 115 668 116
rect 750 120 756 121
rect 750 116 751 120
rect 755 116 756 120
rect 750 115 756 116
rect 838 120 844 121
rect 838 116 839 120
rect 843 116 844 120
rect 838 115 844 116
rect 926 120 932 121
rect 926 116 927 120
rect 931 116 932 120
rect 926 115 932 116
rect 1014 120 1020 121
rect 1014 116 1015 120
rect 1019 116 1020 120
rect 1014 115 1020 116
rect 1112 115 1114 130
rect 111 114 115 115
rect 111 109 115 110
rect 223 114 227 115
rect 223 109 227 110
rect 311 114 315 115
rect 311 109 315 110
rect 399 114 403 115
rect 399 109 403 110
rect 487 114 491 115
rect 487 109 491 110
rect 575 114 579 115
rect 575 109 579 110
rect 663 114 667 115
rect 663 109 667 110
rect 751 114 755 115
rect 751 109 755 110
rect 839 114 843 115
rect 839 109 843 110
rect 927 114 931 115
rect 927 109 931 110
rect 1015 114 1019 115
rect 1015 109 1019 110
rect 1111 114 1115 115
rect 1111 109 1115 110
<< m4c >>
rect 111 1218 115 1222
rect 135 1218 139 1222
rect 223 1218 227 1222
rect 311 1218 315 1222
rect 399 1218 403 1222
rect 1111 1218 1115 1222
rect 151 1168 155 1172
rect 111 1154 115 1158
rect 143 1154 147 1158
rect 387 1168 391 1172
rect 231 1154 235 1158
rect 319 1154 323 1158
rect 407 1154 411 1158
rect 1111 1154 1115 1158
rect 111 1090 115 1094
rect 135 1090 139 1094
rect 223 1090 227 1094
rect 279 1090 283 1094
rect 311 1090 315 1094
rect 367 1090 371 1094
rect 399 1090 403 1094
rect 455 1090 459 1094
rect 543 1090 547 1094
rect 631 1090 635 1094
rect 1111 1090 1115 1094
rect 111 1018 115 1022
rect 287 1018 291 1022
rect 375 1018 379 1022
rect 463 1018 467 1022
rect 519 1018 523 1022
rect 551 1018 555 1022
rect 607 1018 611 1022
rect 639 1018 643 1022
rect 703 1018 707 1022
rect 807 1018 811 1022
rect 911 1018 915 1022
rect 1015 1018 1019 1022
rect 1111 1018 1115 1022
rect 111 954 115 958
rect 399 954 403 958
rect 487 954 491 958
rect 511 954 515 958
rect 575 954 579 958
rect 599 954 603 958
rect 663 954 667 958
rect 695 954 699 958
rect 751 954 755 958
rect 799 954 803 958
rect 415 920 419 924
rect 643 923 647 924
rect 643 920 647 923
rect 111 890 115 894
rect 143 890 147 894
rect 271 890 275 894
rect 407 890 411 894
rect 439 890 443 894
rect 495 890 499 894
rect 583 890 587 894
rect 631 890 635 894
rect 671 890 675 894
rect 759 890 763 894
rect 839 954 843 958
rect 903 954 907 958
rect 927 954 931 958
rect 839 890 843 894
rect 847 890 851 894
rect 935 890 939 894
rect 1007 954 1011 958
rect 1015 954 1019 958
rect 1111 954 1115 958
rect 447 872 451 876
rect 739 872 743 876
rect 1023 890 1027 894
rect 1111 890 1115 894
rect 111 822 115 826
rect 135 822 139 826
rect 263 822 267 826
rect 279 822 283 826
rect 431 822 435 826
rect 463 822 467 826
rect 623 822 627 826
rect 647 822 651 826
rect 831 822 835 826
rect 839 822 843 826
rect 1015 822 1019 826
rect 1111 822 1115 826
rect 191 784 195 788
rect 575 787 579 788
rect 111 746 115 750
rect 143 746 147 750
rect 183 746 187 750
rect 575 784 579 787
rect 287 746 291 750
rect 303 746 307 750
rect 431 746 435 750
rect 471 746 475 750
rect 567 746 571 750
rect 655 746 659 750
rect 719 746 723 750
rect 847 746 851 750
rect 879 746 883 750
rect 1023 746 1027 750
rect 1111 746 1115 750
rect 111 670 115 674
rect 175 670 179 674
rect 295 670 299 674
rect 343 670 347 674
rect 423 670 427 674
rect 455 670 459 674
rect 559 670 563 674
rect 583 670 587 674
rect 711 670 715 674
rect 719 670 723 674
rect 863 670 867 674
rect 871 670 875 674
rect 359 656 363 660
rect 635 656 639 660
rect 551 616 555 620
rect 111 598 115 602
rect 351 598 355 602
rect 463 598 467 602
rect 543 598 547 602
rect 811 616 815 620
rect 591 598 595 602
rect 631 598 635 602
rect 719 598 723 602
rect 727 598 731 602
rect 807 598 811 602
rect 871 598 875 602
rect 1015 670 1019 674
rect 1111 670 1115 674
rect 903 598 907 602
rect 1007 598 1011 602
rect 1023 598 1027 602
rect 1111 598 1115 602
rect 111 526 115 530
rect 479 526 483 530
rect 535 526 539 530
rect 567 526 571 530
rect 623 526 627 530
rect 655 526 659 530
rect 711 526 715 530
rect 743 526 747 530
rect 799 526 803 530
rect 831 526 835 530
rect 895 526 899 530
rect 919 526 923 530
rect 111 454 115 458
rect 271 454 275 458
rect 375 454 379 458
rect 487 454 491 458
rect 575 454 579 458
rect 599 454 603 458
rect 663 454 667 458
rect 719 454 723 458
rect 751 454 755 458
rect 839 454 843 458
rect 847 454 851 458
rect 111 386 115 390
rect 135 386 139 390
rect 263 386 267 390
rect 367 386 371 390
rect 431 386 435 390
rect 151 336 155 340
rect 203 336 207 340
rect 279 336 283 340
rect 479 386 483 390
rect 591 386 595 390
rect 607 386 611 390
rect 711 386 715 390
rect 791 386 795 390
rect 839 386 843 390
rect 927 454 931 458
rect 983 454 987 458
rect 999 526 1003 530
rect 1111 526 1115 530
rect 1111 454 1115 458
rect 975 386 979 390
rect 1111 386 1115 390
rect 539 336 543 340
rect 111 322 115 326
rect 143 322 147 326
rect 271 322 275 326
rect 303 322 307 326
rect 439 322 443 326
rect 487 322 491 326
rect 615 322 619 326
rect 671 322 675 326
rect 111 250 115 254
rect 135 250 139 254
rect 199 250 203 254
rect 295 250 299 254
rect 343 250 347 254
rect 479 250 483 254
rect 615 250 619 254
rect 663 250 667 254
rect 799 322 803 326
rect 855 322 859 326
rect 983 322 987 326
rect 1023 322 1027 326
rect 1111 322 1115 326
rect 751 250 755 254
rect 847 250 851 254
rect 895 250 899 254
rect 1015 250 1019 254
rect 1111 250 1115 254
rect 111 174 115 178
rect 207 174 211 178
rect 231 174 235 178
rect 319 174 323 178
rect 351 174 355 178
rect 407 174 411 178
rect 487 174 491 178
rect 495 174 499 178
rect 583 174 587 178
rect 623 174 627 178
rect 671 174 675 178
rect 759 174 763 178
rect 847 174 851 178
rect 903 174 907 178
rect 935 174 939 178
rect 1023 174 1027 178
rect 1111 174 1115 178
rect 111 110 115 114
rect 223 110 227 114
rect 311 110 315 114
rect 399 110 403 114
rect 487 110 491 114
rect 575 110 579 114
rect 663 110 667 114
rect 751 110 755 114
rect 839 110 843 114
rect 927 110 931 114
rect 1015 110 1019 114
rect 1111 110 1115 114
<< m4 >>
rect 84 1217 85 1223
rect 91 1222 1135 1223
rect 91 1218 111 1222
rect 115 1218 135 1222
rect 139 1218 223 1222
rect 227 1218 311 1222
rect 315 1218 399 1222
rect 403 1218 1111 1222
rect 1115 1218 1135 1222
rect 91 1217 1135 1218
rect 1141 1217 1142 1223
rect 150 1172 156 1173
rect 386 1172 392 1173
rect 150 1168 151 1172
rect 155 1168 387 1172
rect 391 1168 392 1172
rect 150 1167 156 1168
rect 386 1167 392 1168
rect 96 1153 97 1159
rect 103 1158 1147 1159
rect 103 1154 111 1158
rect 115 1154 143 1158
rect 147 1154 231 1158
rect 235 1154 319 1158
rect 323 1154 407 1158
rect 411 1154 1111 1158
rect 1115 1154 1147 1158
rect 103 1153 1147 1154
rect 1153 1153 1154 1159
rect 84 1089 85 1095
rect 91 1094 1135 1095
rect 91 1090 111 1094
rect 115 1090 135 1094
rect 139 1090 223 1094
rect 227 1090 279 1094
rect 283 1090 311 1094
rect 315 1090 367 1094
rect 371 1090 399 1094
rect 403 1090 455 1094
rect 459 1090 543 1094
rect 547 1090 631 1094
rect 635 1090 1111 1094
rect 1115 1090 1135 1094
rect 91 1089 1135 1090
rect 1141 1089 1142 1095
rect 96 1017 97 1023
rect 103 1022 1147 1023
rect 103 1018 111 1022
rect 115 1018 287 1022
rect 291 1018 375 1022
rect 379 1018 463 1022
rect 467 1018 519 1022
rect 523 1018 551 1022
rect 555 1018 607 1022
rect 611 1018 639 1022
rect 643 1018 703 1022
rect 707 1018 807 1022
rect 811 1018 911 1022
rect 915 1018 1015 1022
rect 1019 1018 1111 1022
rect 1115 1018 1147 1022
rect 103 1017 1147 1018
rect 1153 1017 1154 1023
rect 84 953 85 959
rect 91 958 1135 959
rect 91 954 111 958
rect 115 954 399 958
rect 403 954 487 958
rect 491 954 511 958
rect 515 954 575 958
rect 579 954 599 958
rect 603 954 663 958
rect 667 954 695 958
rect 699 954 751 958
rect 755 954 799 958
rect 803 954 839 958
rect 843 954 903 958
rect 907 954 927 958
rect 931 954 1007 958
rect 1011 954 1015 958
rect 1019 954 1111 958
rect 1115 954 1135 958
rect 91 953 1135 954
rect 1141 953 1142 959
rect 414 924 420 925
rect 642 924 648 925
rect 414 920 415 924
rect 419 920 643 924
rect 647 920 648 924
rect 414 919 420 920
rect 642 919 648 920
rect 96 889 97 895
rect 103 894 1147 895
rect 103 890 111 894
rect 115 890 143 894
rect 147 890 271 894
rect 275 890 407 894
rect 411 890 439 894
rect 443 890 495 894
rect 499 890 583 894
rect 587 890 631 894
rect 635 890 671 894
rect 675 890 759 894
rect 763 890 839 894
rect 843 890 847 894
rect 851 890 935 894
rect 939 890 1023 894
rect 1027 890 1111 894
rect 1115 890 1147 894
rect 103 889 1147 890
rect 1153 889 1154 895
rect 446 876 452 877
rect 738 876 744 877
rect 446 872 447 876
rect 451 872 739 876
rect 743 872 744 876
rect 446 871 452 872
rect 738 871 744 872
rect 84 821 85 827
rect 91 826 1135 827
rect 91 822 111 826
rect 115 822 135 826
rect 139 822 263 826
rect 267 822 279 826
rect 283 822 431 826
rect 435 822 463 826
rect 467 822 623 826
rect 627 822 647 826
rect 651 822 831 826
rect 835 822 839 826
rect 843 822 1015 826
rect 1019 822 1111 826
rect 1115 822 1135 826
rect 91 821 1135 822
rect 1141 821 1142 827
rect 190 788 196 789
rect 574 788 580 789
rect 190 784 191 788
rect 195 784 575 788
rect 579 784 580 788
rect 190 783 196 784
rect 574 783 580 784
rect 96 745 97 751
rect 103 750 1147 751
rect 103 746 111 750
rect 115 746 143 750
rect 147 746 183 750
rect 187 746 287 750
rect 291 746 303 750
rect 307 746 431 750
rect 435 746 471 750
rect 475 746 567 750
rect 571 746 655 750
rect 659 746 719 750
rect 723 746 847 750
rect 851 746 879 750
rect 883 746 1023 750
rect 1027 746 1111 750
rect 1115 746 1147 750
rect 103 745 1147 746
rect 1153 745 1154 751
rect 84 669 85 675
rect 91 674 1135 675
rect 91 670 111 674
rect 115 670 175 674
rect 179 670 295 674
rect 299 670 343 674
rect 347 670 423 674
rect 427 670 455 674
rect 459 670 559 674
rect 563 670 583 674
rect 587 670 711 674
rect 715 670 719 674
rect 723 670 863 674
rect 867 670 871 674
rect 875 670 1015 674
rect 1019 670 1111 674
rect 1115 670 1135 674
rect 91 669 1135 670
rect 1141 669 1142 675
rect 358 660 364 661
rect 634 660 640 661
rect 358 656 359 660
rect 363 656 635 660
rect 639 656 640 660
rect 358 655 364 656
rect 634 655 640 656
rect 550 620 556 621
rect 810 620 816 621
rect 550 616 551 620
rect 555 616 811 620
rect 815 616 816 620
rect 550 615 556 616
rect 810 615 816 616
rect 96 597 97 603
rect 103 602 1147 603
rect 103 598 111 602
rect 115 598 351 602
rect 355 598 463 602
rect 467 598 543 602
rect 547 598 591 602
rect 595 598 631 602
rect 635 598 719 602
rect 723 598 727 602
rect 731 598 807 602
rect 811 598 871 602
rect 875 598 903 602
rect 907 598 1007 602
rect 1011 598 1023 602
rect 1027 598 1111 602
rect 1115 598 1147 602
rect 103 597 1147 598
rect 1153 597 1154 603
rect 84 525 85 531
rect 91 530 1135 531
rect 91 526 111 530
rect 115 526 479 530
rect 483 526 535 530
rect 539 526 567 530
rect 571 526 623 530
rect 627 526 655 530
rect 659 526 711 530
rect 715 526 743 530
rect 747 526 799 530
rect 803 526 831 530
rect 835 526 895 530
rect 899 526 919 530
rect 923 526 999 530
rect 1003 526 1111 530
rect 1115 526 1135 530
rect 91 525 1135 526
rect 1141 525 1142 531
rect 96 453 97 459
rect 103 458 1147 459
rect 103 454 111 458
rect 115 454 271 458
rect 275 454 375 458
rect 379 454 487 458
rect 491 454 575 458
rect 579 454 599 458
rect 603 454 663 458
rect 667 454 719 458
rect 723 454 751 458
rect 755 454 839 458
rect 843 454 847 458
rect 851 454 927 458
rect 931 454 983 458
rect 987 454 1111 458
rect 1115 454 1147 458
rect 103 453 1147 454
rect 1153 453 1154 459
rect 84 385 85 391
rect 91 390 1135 391
rect 91 386 111 390
rect 115 386 135 390
rect 139 386 263 390
rect 267 386 367 390
rect 371 386 431 390
rect 435 386 479 390
rect 483 386 591 390
rect 595 386 607 390
rect 611 386 711 390
rect 715 386 791 390
rect 795 386 839 390
rect 843 386 975 390
rect 979 386 1111 390
rect 1115 386 1135 390
rect 91 385 1135 386
rect 1141 385 1142 391
rect 150 340 156 341
rect 202 340 208 341
rect 150 336 151 340
rect 155 336 203 340
rect 207 336 208 340
rect 150 335 156 336
rect 202 335 208 336
rect 278 340 284 341
rect 538 340 544 341
rect 278 336 279 340
rect 283 336 539 340
rect 543 336 544 340
rect 278 335 284 336
rect 538 335 544 336
rect 96 321 97 327
rect 103 326 1147 327
rect 103 322 111 326
rect 115 322 143 326
rect 147 322 271 326
rect 275 322 303 326
rect 307 322 439 326
rect 443 322 487 326
rect 491 322 615 326
rect 619 322 671 326
rect 675 322 799 326
rect 803 322 855 326
rect 859 322 983 326
rect 987 322 1023 326
rect 1027 322 1111 326
rect 1115 322 1147 326
rect 103 321 1147 322
rect 1153 321 1154 327
rect 84 249 85 255
rect 91 254 1135 255
rect 91 250 111 254
rect 115 250 135 254
rect 139 250 199 254
rect 203 250 295 254
rect 299 250 343 254
rect 347 250 479 254
rect 483 250 615 254
rect 619 250 663 254
rect 667 250 751 254
rect 755 250 847 254
rect 851 250 895 254
rect 899 250 1015 254
rect 1019 250 1111 254
rect 1115 250 1135 254
rect 91 249 1135 250
rect 1141 249 1142 255
rect 96 173 97 179
rect 103 178 1147 179
rect 103 174 111 178
rect 115 174 207 178
rect 211 174 231 178
rect 235 174 319 178
rect 323 174 351 178
rect 355 174 407 178
rect 411 174 487 178
rect 491 174 495 178
rect 499 174 583 178
rect 587 174 623 178
rect 627 174 671 178
rect 675 174 759 178
rect 763 174 847 178
rect 851 174 903 178
rect 907 174 935 178
rect 939 174 1023 178
rect 1027 174 1111 178
rect 1115 174 1147 178
rect 103 173 1147 174
rect 1153 173 1154 179
rect 84 109 85 115
rect 91 114 1135 115
rect 91 110 111 114
rect 115 110 223 114
rect 227 110 311 114
rect 315 110 399 114
rect 403 110 487 114
rect 491 110 575 114
rect 579 110 663 114
rect 667 110 751 114
rect 755 110 839 114
rect 843 110 927 114
rect 931 110 1015 114
rect 1019 110 1111 114
rect 1115 110 1135 114
rect 91 109 1135 110
rect 1141 109 1142 115
<< m5c >>
rect 85 1217 91 1223
rect 1135 1217 1141 1223
rect 97 1153 103 1159
rect 1147 1153 1153 1159
rect 85 1089 91 1095
rect 1135 1089 1141 1095
rect 97 1017 103 1023
rect 1147 1017 1153 1023
rect 85 953 91 959
rect 1135 953 1141 959
rect 97 889 103 895
rect 1147 889 1153 895
rect 85 821 91 827
rect 1135 821 1141 827
rect 97 745 103 751
rect 1147 745 1153 751
rect 85 669 91 675
rect 1135 669 1141 675
rect 97 597 103 603
rect 1147 597 1153 603
rect 85 525 91 531
rect 1135 525 1141 531
rect 97 453 103 459
rect 1147 453 1153 459
rect 85 385 91 391
rect 1135 385 1141 391
rect 97 321 103 327
rect 1147 321 1153 327
rect 85 249 91 255
rect 1135 249 1141 255
rect 97 173 103 179
rect 1147 173 1153 179
rect 85 109 91 115
rect 1135 109 1141 115
<< m5 >>
rect 84 1223 92 1224
rect 84 1217 85 1223
rect 91 1217 92 1223
rect 84 1095 92 1217
rect 84 1089 85 1095
rect 91 1089 92 1095
rect 84 959 92 1089
rect 84 953 85 959
rect 91 953 92 959
rect 84 827 92 953
rect 84 821 85 827
rect 91 821 92 827
rect 84 675 92 821
rect 84 669 85 675
rect 91 669 92 675
rect 84 531 92 669
rect 84 525 85 531
rect 91 525 92 531
rect 84 391 92 525
rect 84 385 85 391
rect 91 385 92 391
rect 84 255 92 385
rect 84 249 85 255
rect 91 249 92 255
rect 84 115 92 249
rect 84 109 85 115
rect 91 109 92 115
rect 84 72 92 109
rect 96 1159 104 1224
rect 96 1153 97 1159
rect 103 1153 104 1159
rect 96 1023 104 1153
rect 96 1017 97 1023
rect 103 1017 104 1023
rect 96 895 104 1017
rect 96 889 97 895
rect 103 889 104 895
rect 96 751 104 889
rect 96 745 97 751
rect 103 745 104 751
rect 96 603 104 745
rect 96 597 97 603
rect 103 597 104 603
rect 96 459 104 597
rect 96 453 97 459
rect 103 453 104 459
rect 96 327 104 453
rect 96 321 97 327
rect 103 321 104 327
rect 96 179 104 321
rect 96 173 97 179
rect 103 173 104 179
rect 96 72 104 173
rect 1134 1223 1142 1224
rect 1134 1217 1135 1223
rect 1141 1217 1142 1223
rect 1134 1095 1142 1217
rect 1134 1089 1135 1095
rect 1141 1089 1142 1095
rect 1134 959 1142 1089
rect 1134 953 1135 959
rect 1141 953 1142 959
rect 1134 827 1142 953
rect 1134 821 1135 827
rect 1141 821 1142 827
rect 1134 675 1142 821
rect 1134 669 1135 675
rect 1141 669 1142 675
rect 1134 531 1142 669
rect 1134 525 1135 531
rect 1141 525 1142 531
rect 1134 391 1142 525
rect 1134 385 1135 391
rect 1141 385 1142 391
rect 1134 255 1142 385
rect 1134 249 1135 255
rect 1141 249 1142 255
rect 1134 115 1142 249
rect 1134 109 1135 115
rect 1141 109 1142 115
rect 1134 72 1142 109
rect 1146 1159 1154 1224
rect 1146 1153 1147 1159
rect 1153 1153 1154 1159
rect 1146 1023 1154 1153
rect 1146 1017 1147 1023
rect 1153 1017 1154 1023
rect 1146 895 1154 1017
rect 1146 889 1147 895
rect 1153 889 1154 895
rect 1146 751 1154 889
rect 1146 745 1147 751
rect 1153 745 1154 751
rect 1146 603 1154 745
rect 1146 597 1147 603
rect 1153 597 1154 603
rect 1146 459 1154 597
rect 1146 453 1147 459
rect 1153 453 1154 459
rect 1146 327 1154 453
rect 1146 321 1147 327
rect 1153 321 1154 327
rect 1146 179 1154 321
rect 1146 173 1147 179
rect 1153 173 1154 179
rect 1146 72 1154 173
use welltap_svt  __well_tap__0
timestamp 1731001050
transform 1 0 104 0 1 128
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1731001050
transform 1 0 104 0 1 128
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0MUX2X1  mux_564_6
timestamp 1731001050
transform 1 0 216 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_564_6
timestamp 1731001050
transform 1 0 216 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_565_6
timestamp 1731001050
transform 1 0 304 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_565_6
timestamp 1731001050
transform 1 0 304 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_566_6
timestamp 1731001050
transform 1 0 392 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_566_6
timestamp 1731001050
transform 1 0 392 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_567_6
timestamp 1731001050
transform 1 0 480 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_567_6
timestamp 1731001050
transform 1 0 480 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_568_6
timestamp 1731001050
transform 1 0 568 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_568_6
timestamp 1731001050
transform 1 0 568 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_569_6
timestamp 1731001050
transform 1 0 656 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_569_6
timestamp 1731001050
transform 1 0 656 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_570_6
timestamp 1731001050
transform 1 0 744 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_570_6
timestamp 1731001050
transform 1 0 744 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_571_6
timestamp 1731001050
transform 1 0 832 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_571_6
timestamp 1731001050
transform 1 0 832 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_599_6
timestamp 1731001050
transform 1 0 920 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_599_6
timestamp 1731001050
transform 1 0 920 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_598_6
timestamp 1731001050
transform 1 0 1008 0 1 112
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_598_6
timestamp 1731001050
transform 1 0 1008 0 1 112
box 8 2 80 63
use welltap_svt  __well_tap__1
timestamp 1731001050
transform 1 0 1104 0 1 128
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1731001050
transform 1 0 1104 0 1 128
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_563_6
timestamp 1731001050
transform 1 0 192 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_563_6
timestamp 1731001050
transform 1 0 192 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_562_6
timestamp 1731001050
transform 1 0 336 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_562_6
timestamp 1731001050
transform 1 0 336 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_561_6
timestamp 1731001050
transform 1 0 472 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_561_6
timestamp 1731001050
transform 1 0 472 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_573_6
timestamp 1731001050
transform 1 0 608 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_573_6
timestamp 1731001050
transform 1 0 608 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_572_6
timestamp 1731001050
transform 1 0 744 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_572_6
timestamp 1731001050
transform 1 0 744 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_596_6
timestamp 1731001050
transform 1 0 888 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_596_6
timestamp 1731001050
transform 1 0 888 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_597_6
timestamp 1731001050
transform 1 0 1008 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_597_6
timestamp 1731001050
transform 1 0 1008 0 -1 252
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_558_6
timestamp 1731001050
transform 1 0 128 0 1 260
box 8 2 80 63
use welltap_svt  __well_tap__2
timestamp 1731001050
transform 1 0 104 0 -1 236
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_558_6
timestamp 1731001050
transform 1 0 128 0 1 260
box 8 2 80 63
use welltap_svt  __well_tap__2
timestamp 1731001050
transform 1 0 104 0 -1 236
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_559_6
timestamp 1731001050
transform 1 0 288 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_559_6
timestamp 1731001050
transform 1 0 288 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_560_6
timestamp 1731001050
transform 1 0 472 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_560_6
timestamp 1731001050
transform 1 0 472 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_574_6
timestamp 1731001050
transform 1 0 656 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_574_6
timestamp 1731001050
transform 1 0 656 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_595_6
timestamp 1731001050
transform 1 0 840 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_595_6
timestamp 1731001050
transform 1 0 840 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_594_6
timestamp 1731001050
transform 1 0 1008 0 1 260
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_594_6
timestamp 1731001050
transform 1 0 1008 0 1 260
box 8 2 80 63
use welltap_svt  __well_tap__3
timestamp 1731001050
transform 1 0 1104 0 -1 236
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1731001050
transform 1 0 1104 0 -1 236
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_557_6
timestamp 1731001050
transform 1 0 128 0 -1 388
box 8 2 80 63
use welltap_svt  __well_tap__4
timestamp 1731001050
transform 1 0 104 0 1 276
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_557_6
timestamp 1731001050
transform 1 0 128 0 -1 388
box 8 2 80 63
use welltap_svt  __well_tap__4
timestamp 1731001050
transform 1 0 104 0 1 276
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_556_6
timestamp 1731001050
transform 1 0 256 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_556_6
timestamp 1731001050
transform 1 0 256 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_554_6
timestamp 1731001050
transform 1 0 424 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_554_6
timestamp 1731001050
transform 1 0 424 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_555_6
timestamp 1731001050
transform 1 0 600 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_555_6
timestamp 1731001050
transform 1 0 600 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_575_6
timestamp 1731001050
transform 1 0 784 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_575_6
timestamp 1731001050
transform 1 0 784 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_593_6
timestamp 1731001050
transform 1 0 968 0 -1 388
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_593_6
timestamp 1731001050
transform 1 0 968 0 -1 388
box 8 2 80 63
use welltap_svt  __well_tap__5
timestamp 1731001050
transform 1 0 1104 0 1 276
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1731001050
transform 1 0 1104 0 1 276
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1731001050
transform 1 0 104 0 -1 372
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1731001050
transform 1 0 104 0 -1 372
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_552_6
timestamp 1731001050
transform 1 0 256 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_552_6
timestamp 1731001050
transform 1 0 256 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_553_6
timestamp 1731001050
transform 1 0 360 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_553_6
timestamp 1731001050
transform 1 0 360 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_551_6
timestamp 1731001050
transform 1 0 472 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_551_6
timestamp 1731001050
transform 1 0 472 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_549_6
timestamp 1731001050
transform 1 0 584 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_549_6
timestamp 1731001050
transform 1 0 584 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_550_6
timestamp 1731001050
transform 1 0 704 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_550_6
timestamp 1731001050
transform 1 0 704 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_576_6
timestamp 1731001050
transform 1 0 832 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_576_6
timestamp 1731001050
transform 1 0 832 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_592_6
timestamp 1731001050
transform 1 0 968 0 1 392
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_592_6
timestamp 1731001050
transform 1 0 968 0 1 392
box 8 2 80 63
use welltap_svt  __well_tap__7
timestamp 1731001050
transform 1 0 1104 0 -1 372
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1731001050
transform 1 0 1104 0 -1 372
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1731001050
transform 1 0 104 0 1 408
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1731001050
transform 1 0 104 0 1 408
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_547_6
timestamp 1731001050
transform 1 0 472 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_547_6
timestamp 1731001050
transform 1 0 472 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_548_6
timestamp 1731001050
transform 1 0 560 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_548_6
timestamp 1731001050
transform 1 0 560 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_546_6
timestamp 1731001050
transform 1 0 648 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_546_6
timestamp 1731001050
transform 1 0 648 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_545_6
timestamp 1731001050
transform 1 0 736 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_545_6
timestamp 1731001050
transform 1 0 736 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_544_6
timestamp 1731001050
transform 1 0 824 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_544_6
timestamp 1731001050
transform 1 0 824 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_577_6
timestamp 1731001050
transform 1 0 912 0 -1 528
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_577_6
timestamp 1731001050
transform 1 0 912 0 -1 528
box 8 2 80 63
use welltap_svt  __well_tap__9
timestamp 1731001050
transform 1 0 1104 0 1 408
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1731001050
transform 1 0 1104 0 1 408
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1731001050
transform 1 0 104 0 -1 512
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1731001050
transform 1 0 104 0 -1 512
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_540_6
timestamp 1731001050
transform 1 0 528 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_540_6
timestamp 1731001050
transform 1 0 528 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_541_6
timestamp 1731001050
transform 1 0 616 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_541_6
timestamp 1731001050
transform 1 0 616 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_542_6
timestamp 1731001050
transform 1 0 704 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_542_6
timestamp 1731001050
transform 1 0 704 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_543_6
timestamp 1731001050
transform 1 0 792 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_543_6
timestamp 1731001050
transform 1 0 792 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_578_6
timestamp 1731001050
transform 1 0 888 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_578_6
timestamp 1731001050
transform 1 0 888 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_591_6
timestamp 1731001050
transform 1 0 992 0 1 536
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_591_6
timestamp 1731001050
transform 1 0 992 0 1 536
box 8 2 80 63
use welltap_svt  __well_tap__11
timestamp 1731001050
transform 1 0 1104 0 -1 512
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1731001050
transform 1 0 1104 0 -1 512
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1731001050
transform 1 0 104 0 1 552
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1731001050
transform 1 0 104 0 1 552
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1731001050
transform 1 0 1104 0 1 552
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1731001050
transform 1 0 1104 0 1 552
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1731001050
transform 1 0 104 0 -1 656
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1731001050
transform 1 0 104 0 -1 656
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_535_6
timestamp 1731001050
transform 1 0 336 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_535_6
timestamp 1731001050
transform 1 0 336 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_536_6
timestamp 1731001050
transform 1 0 448 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_536_6
timestamp 1731001050
transform 1 0 448 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_537_6
timestamp 1731001050
transform 1 0 576 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_537_6
timestamp 1731001050
transform 1 0 576 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_538_6
timestamp 1731001050
transform 1 0 712 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_538_6
timestamp 1731001050
transform 1 0 712 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_539_6
timestamp 1731001050
transform 1 0 856 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_539_6
timestamp 1731001050
transform 1 0 856 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_590_6
timestamp 1731001050
transform 1 0 1008 0 -1 672
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_590_6
timestamp 1731001050
transform 1 0 1008 0 -1 672
box 8 2 80 63
use welltap_svt  __well_tap__15
timestamp 1731001050
transform 1 0 1104 0 -1 656
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1731001050
transform 1 0 1104 0 -1 656
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1731001050
transform 1 0 104 0 1 700
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1731001050
transform 1 0 104 0 1 700
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_530_6
timestamp 1731001050
transform 1 0 168 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_530_6
timestamp 1731001050
transform 1 0 168 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_531_6
timestamp 1731001050
transform 1 0 288 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_531_6
timestamp 1731001050
transform 1 0 288 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_532_6
timestamp 1731001050
transform 1 0 416 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_532_6
timestamp 1731001050
transform 1 0 416 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_533_6
timestamp 1731001050
transform 1 0 552 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_533_6
timestamp 1731001050
transform 1 0 552 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_534_6
timestamp 1731001050
transform 1 0 704 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_534_6
timestamp 1731001050
transform 1 0 704 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_579_6
timestamp 1731001050
transform 1 0 864 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_579_6
timestamp 1731001050
transform 1 0 864 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_589_6
timestamp 1731001050
transform 1 0 1008 0 1 684
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_589_6
timestamp 1731001050
transform 1 0 1008 0 1 684
box 8 2 80 63
use welltap_svt  __well_tap__17
timestamp 1731001050
transform 1 0 1104 0 1 700
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1731001050
transform 1 0 1104 0 1 700
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_526_6
timestamp 1731001050
transform 1 0 128 0 -1 824
box 8 2 80 63
use welltap_svt  __well_tap__18
timestamp 1731001050
transform 1 0 104 0 -1 808
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_526_6
timestamp 1731001050
transform 1 0 128 0 -1 824
box 8 2 80 63
use welltap_svt  __well_tap__18
timestamp 1731001050
transform 1 0 104 0 -1 808
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_527_6
timestamp 1731001050
transform 1 0 272 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_527_6
timestamp 1731001050
transform 1 0 272 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_528_6
timestamp 1731001050
transform 1 0 456 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_528_6
timestamp 1731001050
transform 1 0 456 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_529_6
timestamp 1731001050
transform 1 0 640 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_529_6
timestamp 1731001050
transform 1 0 640 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_580_6
timestamp 1731001050
transform 1 0 832 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_580_6
timestamp 1731001050
transform 1 0 832 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_588_6
timestamp 1731001050
transform 1 0 1008 0 -1 824
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_588_6
timestamp 1731001050
transform 1 0 1008 0 -1 824
box 8 2 80 63
use welltap_svt  __well_tap__19
timestamp 1731001050
transform 1 0 1104 0 -1 808
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1731001050
transform 1 0 1104 0 -1 808
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_525_6
timestamp 1731001050
transform 1 0 128 0 1 828
box 8 2 80 63
use welltap_svt  __well_tap__20
timestamp 1731001050
transform 1 0 104 0 1 844
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_525_6
timestamp 1731001050
transform 1 0 128 0 1 828
box 8 2 80 63
use welltap_svt  __well_tap__20
timestamp 1731001050
transform 1 0 104 0 1 844
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_524_6
timestamp 1731001050
transform 1 0 256 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_524_6
timestamp 1731001050
transform 1 0 256 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_523_6
timestamp 1731001050
transform 1 0 424 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_523_6
timestamp 1731001050
transform 1 0 424 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_521_6
timestamp 1731001050
transform 1 0 616 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_521_6
timestamp 1731001050
transform 1 0 616 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_522_6
timestamp 1731001050
transform 1 0 824 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_522_6
timestamp 1731001050
transform 1 0 824 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_587_6
timestamp 1731001050
transform 1 0 1008 0 1 828
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_587_6
timestamp 1731001050
transform 1 0 1008 0 1 828
box 8 2 80 63
use welltap_svt  __well_tap__21
timestamp 1731001050
transform 1 0 1104 0 1 844
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1731001050
transform 1 0 1104 0 1 844
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1731001050
transform 1 0 104 0 -1 940
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1731001050
transform 1 0 104 0 -1 940
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_518_6
timestamp 1731001050
transform 1 0 392 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_518_6
timestamp 1731001050
transform 1 0 392 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_519_6
timestamp 1731001050
transform 1 0 480 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_519_6
timestamp 1731001050
transform 1 0 480 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_520_6
timestamp 1731001050
transform 1 0 568 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_520_6
timestamp 1731001050
transform 1 0 568 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_517_6
timestamp 1731001050
transform 1 0 656 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_517_6
timestamp 1731001050
transform 1 0 656 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_581_6
timestamp 1731001050
transform 1 0 744 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_581_6
timestamp 1731001050
transform 1 0 744 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_582_6
timestamp 1731001050
transform 1 0 832 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_582_6
timestamp 1731001050
transform 1 0 832 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_585_6
timestamp 1731001050
transform 1 0 920 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_585_6
timestamp 1731001050
transform 1 0 920 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_586_6
timestamp 1731001050
transform 1 0 1008 0 -1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_586_6
timestamp 1731001050
transform 1 0 1008 0 -1 956
box 8 2 80 63
use welltap_svt  __well_tap__23
timestamp 1731001050
transform 1 0 1104 0 -1 940
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1731001050
transform 1 0 1104 0 -1 940
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1731001050
transform 1 0 104 0 1 972
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1731001050
transform 1 0 104 0 1 972
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_513_6
timestamp 1731001050
transform 1 0 504 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_513_6
timestamp 1731001050
transform 1 0 504 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_514_6
timestamp 1731001050
transform 1 0 592 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_514_6
timestamp 1731001050
transform 1 0 592 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_515_6
timestamp 1731001050
transform 1 0 688 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_515_6
timestamp 1731001050
transform 1 0 688 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_516_6
timestamp 1731001050
transform 1 0 792 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_516_6
timestamp 1731001050
transform 1 0 792 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_583_6
timestamp 1731001050
transform 1 0 896 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_583_6
timestamp 1731001050
transform 1 0 896 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_584_6
timestamp 1731001050
transform 1 0 1000 0 1 956
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_584_6
timestamp 1731001050
transform 1 0 1000 0 1 956
box 8 2 80 63
use welltap_svt  __well_tap__25
timestamp 1731001050
transform 1 0 1104 0 1 972
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1731001050
transform 1 0 1104 0 1 972
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1731001050
transform 1 0 104 0 -1 1076
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1731001050
transform 1 0 104 0 -1 1076
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_58_6
timestamp 1731001050
transform 1 0 272 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_58_6
timestamp 1731001050
transform 1 0 272 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_59_6
timestamp 1731001050
transform 1 0 360 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_59_6
timestamp 1731001050
transform 1 0 360 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_510_6
timestamp 1731001050
transform 1 0 448 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_510_6
timestamp 1731001050
transform 1 0 448 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_511_6
timestamp 1731001050
transform 1 0 536 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_511_6
timestamp 1731001050
transform 1 0 536 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_512_6
timestamp 1731001050
transform 1 0 624 0 -1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_512_6
timestamp 1731001050
transform 1 0 624 0 -1 1092
box 8 2 80 63
use welltap_svt  __well_tap__27
timestamp 1731001050
transform 1 0 1104 0 -1 1076
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1731001050
transform 1 0 1104 0 -1 1076
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_54_6
timestamp 1731001050
transform 1 0 128 0 1 1092
box 8 2 80 63
use welltap_svt  __well_tap__28
timestamp 1731001050
transform 1 0 104 0 1 1108
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_54_6
timestamp 1731001050
transform 1 0 128 0 1 1092
box 8 2 80 63
use welltap_svt  __well_tap__28
timestamp 1731001050
transform 1 0 104 0 1 1108
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_55_6
timestamp 1731001050
transform 1 0 216 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_55_6
timestamp 1731001050
transform 1 0 216 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_56_6
timestamp 1731001050
transform 1 0 304 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_56_6
timestamp 1731001050
transform 1 0 304 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_57_6
timestamp 1731001050
transform 1 0 392 0 1 1092
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_57_6
timestamp 1731001050
transform 1 0 392 0 1 1092
box 8 2 80 63
use welltap_svt  __well_tap__29
timestamp 1731001050
transform 1 0 1104 0 1 1108
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1731001050
transform 1 0 1104 0 1 1108
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_50_6
timestamp 1731001050
transform 1 0 128 0 -1 1220
box 8 2 80 63
use welltap_svt  __well_tap__30
timestamp 1731001050
transform 1 0 104 0 -1 1204
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_50_6
timestamp 1731001050
transform 1 0 128 0 -1 1220
box 8 2 80 63
use welltap_svt  __well_tap__30
timestamp 1731001050
transform 1 0 104 0 -1 1204
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_51_6
timestamp 1731001050
transform 1 0 216 0 -1 1220
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_51_6
timestamp 1731001050
transform 1 0 216 0 -1 1220
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_52_6
timestamp 1731001050
transform 1 0 304 0 -1 1220
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_52_6
timestamp 1731001050
transform 1 0 304 0 -1 1220
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_53_6
timestamp 1731001050
transform 1 0 392 0 -1 1220
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_53_6
timestamp 1731001050
transform 1 0 392 0 -1 1220
box 8 2 80 63
use welltap_svt  __well_tap__31
timestamp 1731001050
transform 1 0 1104 0 -1 1204
box 8 4 12 24
use welltap_svt  __well_tap__31
timestamp 1731001050
transform 1 0 1104 0 -1 1204
box 8 4 12 24
<< end >>
