magic
tech sky130l
timestamp 1730591762
<< m1 >>
rect 704 483 708 527
rect 704 375 708 427
rect 392 267 396 319
rect 592 307 596 355
rect 696 267 700 319
rect 128 163 132 211
rect 704 163 708 211
<< m2c >>
rect 111 829 115 833
rect 775 829 779 833
rect 111 811 115 815
rect 775 811 779 815
rect 202 799 206 803
rect 256 799 260 803
rect 314 799 318 803
rect 368 799 372 803
rect 426 799 430 803
rect 480 799 484 803
rect 202 779 206 783
rect 258 775 262 779
rect 314 775 318 779
rect 370 775 374 779
rect 426 775 430 779
rect 111 765 115 769
rect 775 765 779 769
rect 111 747 115 751
rect 775 747 779 751
rect 111 721 115 725
rect 775 721 779 725
rect 111 703 115 707
rect 775 703 779 707
rect 336 691 340 695
rect 395 691 399 695
rect 450 691 454 695
rect 506 691 510 695
rect 562 691 566 695
rect 442 683 446 687
rect 218 679 222 683
rect 274 679 278 683
rect 330 679 334 683
rect 386 679 390 683
rect 498 679 502 683
rect 554 679 558 683
rect 610 679 614 683
rect 666 679 670 683
rect 722 679 726 683
rect 111 669 115 673
rect 775 669 779 673
rect 111 651 115 655
rect 775 651 779 655
rect 111 613 115 617
rect 775 613 779 617
rect 111 595 115 599
rect 775 595 779 599
rect 144 583 148 587
rect 200 583 204 587
rect 272 583 276 587
rect 360 583 364 587
rect 450 583 454 587
rect 547 583 551 587
rect 640 583 644 587
rect 722 583 726 587
rect 146 567 150 571
rect 722 567 726 571
rect 202 563 206 567
rect 298 563 302 567
rect 402 563 406 567
rect 514 563 518 567
rect 626 563 630 567
rect 111 553 115 557
rect 775 553 779 557
rect 111 535 115 539
rect 775 535 779 539
rect 704 527 708 531
rect 111 509 115 513
rect 111 491 115 495
rect 775 509 779 513
rect 775 491 779 495
rect 192 479 196 483
rect 280 479 284 483
rect 376 479 380 483
rect 488 479 492 483
rect 608 479 612 483
rect 704 479 708 483
rect 720 479 724 483
rect 314 467 318 471
rect 722 467 726 471
rect 370 463 374 467
rect 426 463 430 467
rect 490 463 494 467
rect 562 463 566 467
rect 642 463 646 467
rect 111 453 115 457
rect 775 453 779 457
rect 111 435 115 439
rect 775 435 779 439
rect 704 427 708 431
rect 111 401 115 405
rect 111 383 115 387
rect 775 401 779 405
rect 775 383 779 387
rect 384 371 388 375
rect 442 371 446 375
rect 496 371 500 375
rect 552 371 556 375
rect 608 371 612 375
rect 664 371 668 375
rect 704 371 708 375
rect 720 371 724 375
rect 474 359 478 363
rect 714 359 718 363
rect 298 355 302 359
rect 354 355 358 359
rect 410 355 414 359
rect 546 355 550 359
rect 592 355 596 359
rect 626 355 630 359
rect 111 345 115 349
rect 111 327 115 331
rect 392 319 396 323
rect 111 293 115 297
rect 111 275 115 279
rect 775 345 779 349
rect 775 327 779 331
rect 592 303 596 307
rect 696 319 700 323
rect 775 293 779 297
rect 775 275 779 279
rect 168 263 172 267
rect 250 263 254 267
rect 328 263 332 267
rect 392 263 396 267
rect 416 263 420 267
rect 512 263 516 267
rect 610 263 614 267
rect 696 263 700 267
rect 712 263 716 267
rect 362 251 366 255
rect 618 251 622 255
rect 146 247 150 251
rect 242 247 246 251
rect 490 247 494 251
rect 722 247 726 251
rect 111 237 115 241
rect 775 237 779 241
rect 111 219 115 223
rect 775 219 779 223
rect 128 211 132 215
rect 111 189 115 193
rect 111 171 115 175
rect 704 211 708 215
rect 775 189 779 193
rect 775 171 779 175
rect 128 159 132 163
rect 144 159 148 163
rect 208 159 212 163
rect 296 159 300 163
rect 400 159 404 163
rect 504 159 508 163
rect 616 159 620 163
rect 704 159 708 163
rect 720 159 724 163
rect 162 139 166 143
rect 722 139 726 143
rect 218 135 222 139
rect 274 135 278 139
rect 330 135 334 139
rect 386 135 390 139
rect 442 135 446 139
rect 498 135 502 139
rect 554 135 558 139
rect 610 135 614 139
rect 666 135 670 139
rect 111 125 115 129
rect 775 125 779 129
rect 111 107 115 111
rect 775 107 779 111
<< m2 >>
rect 146 841 152 842
rect 146 837 147 841
rect 151 837 152 841
rect 146 836 152 837
rect 202 841 208 842
rect 202 837 203 841
rect 207 837 208 841
rect 202 836 208 837
rect 258 841 264 842
rect 258 837 259 841
rect 263 837 264 841
rect 258 836 264 837
rect 314 841 320 842
rect 314 837 315 841
rect 319 837 320 841
rect 314 836 320 837
rect 370 841 376 842
rect 370 837 371 841
rect 375 837 376 841
rect 370 836 376 837
rect 426 841 432 842
rect 426 837 427 841
rect 431 837 432 841
rect 426 836 432 837
rect 482 841 488 842
rect 482 837 483 841
rect 487 837 488 841
rect 482 836 488 837
rect 110 833 116 834
rect 110 829 111 833
rect 115 829 116 833
rect 110 828 116 829
rect 774 833 780 834
rect 774 829 775 833
rect 779 829 780 833
rect 774 828 780 829
rect 110 815 116 816
rect 110 811 111 815
rect 115 811 116 815
rect 190 815 196 816
rect 190 814 191 815
rect 153 812 191 814
rect 110 810 116 811
rect 190 811 191 812
rect 195 811 196 815
rect 302 815 308 816
rect 302 814 303 815
rect 209 812 242 814
rect 265 812 303 814
rect 190 810 196 811
rect 170 803 176 804
rect 170 799 171 803
rect 175 799 176 803
rect 170 798 176 799
rect 198 803 207 804
rect 198 799 199 803
rect 206 799 207 803
rect 198 798 207 799
rect 226 803 232 804
rect 226 799 227 803
rect 231 799 232 803
rect 240 802 242 812
rect 302 811 303 812
rect 307 811 308 815
rect 414 815 420 816
rect 414 814 415 815
rect 321 812 350 814
rect 377 812 415 814
rect 302 810 308 811
rect 255 803 261 804
rect 255 802 256 803
rect 240 800 256 802
rect 226 798 232 799
rect 255 799 256 800
rect 260 799 261 803
rect 255 798 261 799
rect 282 803 288 804
rect 282 799 283 803
rect 287 799 288 803
rect 282 798 288 799
rect 310 803 319 804
rect 310 799 311 803
rect 318 799 319 803
rect 310 798 319 799
rect 338 803 344 804
rect 338 799 339 803
rect 343 799 344 803
rect 348 802 350 812
rect 414 811 415 812
rect 419 811 420 815
rect 478 815 484 816
rect 433 812 462 814
rect 414 810 420 811
rect 367 803 373 804
rect 367 802 368 803
rect 348 800 368 802
rect 338 798 344 799
rect 367 799 368 800
rect 372 799 373 803
rect 367 798 373 799
rect 394 803 400 804
rect 394 799 395 803
rect 399 799 400 803
rect 394 798 400 799
rect 422 803 431 804
rect 422 799 423 803
rect 430 799 431 803
rect 422 798 431 799
rect 450 803 456 804
rect 450 799 451 803
rect 455 799 456 803
rect 460 802 462 812
rect 478 811 479 815
rect 483 811 484 815
rect 478 810 484 811
rect 774 815 780 816
rect 774 811 775 815
rect 779 811 780 815
rect 774 810 780 811
rect 479 803 485 804
rect 479 802 480 803
rect 460 800 480 802
rect 450 798 456 799
rect 479 799 480 800
rect 484 799 485 803
rect 479 798 485 799
rect 506 803 512 804
rect 506 799 507 803
rect 511 799 512 803
rect 506 798 512 799
rect 478 787 484 788
rect 478 786 479 787
rect 220 784 479 786
rect 201 783 207 784
rect 201 779 202 783
rect 206 782 207 783
rect 220 782 222 784
rect 478 783 479 784
rect 483 783 484 787
rect 478 782 484 783
rect 206 780 222 782
rect 226 781 232 782
rect 206 779 207 780
rect 201 778 207 779
rect 226 777 227 781
rect 231 777 232 781
rect 282 781 288 782
rect 257 779 263 780
rect 257 778 258 779
rect 226 776 232 777
rect 236 776 258 778
rect 236 770 238 776
rect 257 775 258 776
rect 262 775 263 779
rect 282 777 283 781
rect 287 777 288 781
rect 338 781 344 782
rect 313 779 319 780
rect 313 778 314 779
rect 282 776 288 777
rect 292 776 314 778
rect 257 774 263 775
rect 292 770 294 776
rect 313 775 314 776
rect 318 775 319 779
rect 338 777 339 781
rect 343 777 344 781
rect 394 781 400 782
rect 369 779 375 780
rect 369 778 370 779
rect 338 776 344 777
rect 348 776 370 778
rect 313 774 319 775
rect 348 770 350 776
rect 369 775 370 776
rect 374 775 375 779
rect 394 777 395 781
rect 399 777 400 781
rect 450 781 456 782
rect 425 779 431 780
rect 425 778 426 779
rect 394 776 400 777
rect 404 776 426 778
rect 369 774 375 775
rect 404 770 406 776
rect 425 775 426 776
rect 430 775 431 779
rect 450 777 451 781
rect 455 777 456 781
rect 450 776 456 777
rect 425 774 431 775
rect 110 769 116 770
rect 110 765 111 769
rect 115 765 116 769
rect 209 768 238 770
rect 265 768 294 770
rect 321 768 350 770
rect 377 768 406 770
rect 774 769 780 770
rect 110 764 116 765
rect 774 765 775 769
rect 779 765 780 769
rect 774 764 780 765
rect 110 751 116 752
rect 110 747 111 751
rect 115 747 116 751
rect 110 746 116 747
rect 346 751 352 752
rect 346 747 347 751
rect 351 750 352 751
rect 774 751 780 752
rect 351 748 418 750
rect 351 747 352 748
rect 346 746 352 747
rect 202 743 208 744
rect 202 739 203 743
rect 207 739 208 743
rect 202 738 208 739
rect 258 743 264 744
rect 258 739 259 743
rect 263 739 264 743
rect 258 738 264 739
rect 314 743 320 744
rect 314 739 315 743
rect 319 739 320 743
rect 314 738 320 739
rect 370 743 376 744
rect 370 739 371 743
rect 375 739 376 743
rect 416 741 418 748
rect 774 747 775 751
rect 779 747 780 751
rect 774 746 780 747
rect 426 743 432 744
rect 370 738 376 739
rect 426 739 427 743
rect 431 739 432 743
rect 426 738 432 739
rect 338 733 344 734
rect 338 729 339 733
rect 343 729 344 733
rect 338 728 344 729
rect 394 733 400 734
rect 394 729 395 733
rect 399 729 400 733
rect 394 728 400 729
rect 450 733 456 734
rect 450 729 451 733
rect 455 729 456 733
rect 450 728 456 729
rect 506 733 512 734
rect 506 729 507 733
rect 511 729 512 733
rect 506 728 512 729
rect 562 733 568 734
rect 562 729 563 733
rect 567 729 568 733
rect 562 728 568 729
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 110 720 116 721
rect 774 725 780 726
rect 774 721 775 725
rect 779 721 780 725
rect 774 720 780 721
rect 442 715 448 716
rect 442 711 443 715
rect 447 714 448 715
rect 447 712 562 714
rect 447 711 448 712
rect 442 710 448 711
rect 110 707 116 708
rect 110 703 111 707
rect 115 703 116 707
rect 382 707 388 708
rect 382 706 383 707
rect 345 704 383 706
rect 110 702 116 703
rect 382 703 383 704
rect 387 703 388 707
rect 401 704 445 706
rect 457 704 501 706
rect 513 704 557 706
rect 560 705 562 712
rect 774 707 780 708
rect 382 702 388 703
rect 443 698 445 704
rect 499 698 501 704
rect 555 698 557 704
rect 774 703 775 707
rect 779 703 780 707
rect 774 702 780 703
rect 443 696 453 698
rect 499 696 507 698
rect 555 696 563 698
rect 335 695 341 696
rect 335 691 336 695
rect 340 694 341 695
rect 346 695 352 696
rect 346 694 347 695
rect 340 692 347 694
rect 340 691 341 692
rect 335 690 341 691
rect 346 691 347 692
rect 351 691 352 695
rect 346 690 352 691
rect 362 695 368 696
rect 362 691 363 695
rect 367 691 368 695
rect 362 690 368 691
rect 386 695 392 696
rect 386 691 387 695
rect 391 694 392 695
rect 394 695 400 696
rect 394 694 395 695
rect 391 692 395 694
rect 391 691 392 692
rect 386 690 392 691
rect 394 691 395 692
rect 399 691 400 695
rect 394 690 400 691
rect 418 695 424 696
rect 418 691 419 695
rect 423 691 424 695
rect 418 690 424 691
rect 449 695 455 696
rect 449 691 450 695
rect 454 691 455 695
rect 449 690 455 691
rect 474 695 480 696
rect 474 691 475 695
rect 479 691 480 695
rect 474 690 480 691
rect 505 695 511 696
rect 505 691 506 695
rect 510 691 511 695
rect 505 690 511 691
rect 530 695 536 696
rect 530 691 531 695
rect 535 691 536 695
rect 530 690 536 691
rect 561 695 567 696
rect 561 691 562 695
rect 566 691 567 695
rect 561 690 567 691
rect 586 695 592 696
rect 586 691 587 695
rect 591 691 592 695
rect 586 690 592 691
rect 441 687 448 688
rect 242 685 248 686
rect 217 683 223 684
rect 217 679 218 683
rect 222 682 223 683
rect 234 683 240 684
rect 234 682 235 683
rect 222 680 235 682
rect 222 679 223 680
rect 217 678 223 679
rect 234 679 235 680
rect 239 679 240 683
rect 242 681 243 685
rect 247 681 248 685
rect 298 685 304 686
rect 273 683 279 684
rect 273 682 274 683
rect 242 680 248 681
rect 252 680 274 682
rect 234 678 240 679
rect 252 674 254 680
rect 273 679 274 680
rect 278 679 279 683
rect 298 681 299 685
rect 303 681 304 685
rect 354 685 360 686
rect 329 683 335 684
rect 329 682 330 683
rect 298 680 304 681
rect 319 680 330 682
rect 273 678 279 679
rect 319 674 321 680
rect 329 679 330 680
rect 334 679 335 683
rect 354 681 355 685
rect 359 681 360 685
rect 410 685 416 686
rect 354 680 360 681
rect 385 683 391 684
rect 329 678 335 679
rect 385 679 386 683
rect 390 682 391 683
rect 390 680 406 682
rect 410 681 411 685
rect 415 681 416 685
rect 441 683 442 687
rect 447 683 448 687
rect 441 682 448 683
rect 466 685 472 686
rect 410 680 416 681
rect 466 681 467 685
rect 471 681 472 685
rect 522 685 528 686
rect 466 680 472 681
rect 497 683 503 684
rect 390 679 391 680
rect 385 678 391 679
rect 404 678 406 680
rect 497 679 498 683
rect 502 682 503 683
rect 506 683 512 684
rect 506 682 507 683
rect 502 680 507 682
rect 502 679 503 680
rect 497 678 503 679
rect 506 679 507 680
rect 511 679 512 683
rect 522 681 523 685
rect 527 681 528 685
rect 578 685 584 686
rect 553 683 559 684
rect 553 682 554 683
rect 522 680 528 681
rect 532 680 554 682
rect 506 678 512 679
rect 404 676 414 678
rect 110 673 116 674
rect 110 669 111 673
rect 115 669 116 673
rect 225 672 254 674
rect 281 672 321 674
rect 350 671 356 672
rect 350 670 351 671
rect 110 668 116 669
rect 337 668 351 670
rect 350 667 351 668
rect 355 667 356 671
rect 412 670 414 676
rect 532 674 534 680
rect 553 679 554 680
rect 558 679 559 683
rect 578 681 579 685
rect 583 681 584 685
rect 634 685 640 686
rect 609 683 615 684
rect 609 682 610 683
rect 578 680 584 681
rect 588 680 610 682
rect 553 678 559 679
rect 588 674 590 680
rect 609 679 610 680
rect 614 679 615 683
rect 634 681 635 685
rect 639 681 640 685
rect 690 685 696 686
rect 665 683 671 684
rect 665 682 666 683
rect 634 680 640 681
rect 644 680 666 682
rect 609 678 615 679
rect 644 674 646 680
rect 665 679 666 680
rect 670 679 671 683
rect 690 681 691 685
rect 695 681 696 685
rect 746 685 752 686
rect 690 680 696 681
rect 721 683 727 684
rect 665 678 671 679
rect 721 679 722 683
rect 726 679 727 683
rect 746 681 747 685
rect 751 681 752 685
rect 746 680 752 681
rect 721 678 727 679
rect 684 676 725 678
rect 684 674 686 676
rect 505 672 534 674
rect 561 672 590 674
rect 617 672 646 674
rect 673 672 686 674
rect 774 673 780 674
rect 350 666 356 667
rect 234 663 240 664
rect 234 659 235 663
rect 239 662 240 663
rect 384 662 386 669
rect 412 668 441 670
rect 774 669 775 673
rect 779 669 780 673
rect 774 668 780 669
rect 239 660 386 662
rect 239 659 240 660
rect 234 658 240 659
rect 110 655 116 656
rect 110 651 111 655
rect 115 651 116 655
rect 110 650 116 651
rect 774 655 780 656
rect 774 651 775 655
rect 779 651 780 655
rect 774 650 780 651
rect 218 647 224 648
rect 218 643 219 647
rect 223 643 224 647
rect 218 642 224 643
rect 274 647 280 648
rect 274 643 275 647
rect 279 643 280 647
rect 274 642 280 643
rect 330 647 336 648
rect 330 643 331 647
rect 335 643 336 647
rect 330 642 336 643
rect 386 647 392 648
rect 386 643 387 647
rect 391 643 392 647
rect 386 642 392 643
rect 442 647 448 648
rect 442 643 443 647
rect 447 643 448 647
rect 442 642 448 643
rect 498 647 504 648
rect 498 643 499 647
rect 503 643 504 647
rect 498 642 504 643
rect 554 647 560 648
rect 554 643 555 647
rect 559 643 560 647
rect 554 642 560 643
rect 610 647 616 648
rect 610 643 611 647
rect 615 643 616 647
rect 610 642 616 643
rect 666 647 672 648
rect 666 643 667 647
rect 671 643 672 647
rect 722 647 728 648
rect 666 642 672 643
rect 650 639 656 640
rect 650 635 651 639
rect 655 638 656 639
rect 712 638 714 645
rect 722 643 723 647
rect 727 643 728 647
rect 722 642 728 643
rect 655 636 714 638
rect 655 635 656 636
rect 650 634 656 635
rect 506 627 512 628
rect 146 625 152 626
rect 146 621 147 625
rect 151 621 152 625
rect 146 620 152 621
rect 202 625 208 626
rect 202 621 203 625
rect 207 621 208 625
rect 202 620 208 621
rect 274 625 280 626
rect 274 621 275 625
rect 279 621 280 625
rect 274 620 280 621
rect 362 625 368 626
rect 362 621 363 625
rect 367 621 368 625
rect 362 620 368 621
rect 450 625 456 626
rect 450 621 451 625
rect 455 621 456 625
rect 506 623 507 627
rect 511 626 512 627
rect 511 624 537 626
rect 546 625 552 626
rect 511 623 512 624
rect 506 622 512 623
rect 450 620 456 621
rect 546 621 547 625
rect 551 621 552 625
rect 546 620 552 621
rect 642 625 648 626
rect 642 621 643 625
rect 647 621 648 625
rect 642 620 648 621
rect 722 625 728 626
rect 722 621 723 625
rect 727 621 728 625
rect 722 620 728 621
rect 110 617 116 618
rect 110 613 111 617
rect 115 613 116 617
rect 110 612 116 613
rect 774 617 780 618
rect 774 613 775 617
rect 779 613 780 617
rect 774 612 780 613
rect 274 607 280 608
rect 274 603 275 607
rect 279 606 280 607
rect 279 604 450 606
rect 279 603 280 604
rect 274 602 280 603
rect 110 599 116 600
rect 110 595 111 599
rect 115 595 116 599
rect 110 594 116 595
rect 146 599 152 600
rect 146 595 147 599
rect 151 595 152 599
rect 146 594 152 595
rect 160 596 201 598
rect 216 596 273 598
rect 369 596 406 598
rect 448 597 450 604
rect 722 599 728 600
rect 649 596 681 598
rect 143 587 149 588
rect 143 583 144 587
rect 148 586 149 587
rect 160 586 162 596
rect 148 584 162 586
rect 170 587 176 588
rect 148 583 149 584
rect 143 582 149 583
rect 170 583 171 587
rect 175 583 176 587
rect 170 582 176 583
rect 199 587 205 588
rect 199 583 200 587
rect 204 586 205 587
rect 216 586 218 596
rect 204 584 218 586
rect 226 587 232 588
rect 204 583 205 584
rect 199 582 205 583
rect 226 583 227 587
rect 231 583 232 587
rect 226 582 232 583
rect 271 587 280 588
rect 271 583 272 587
rect 279 583 280 587
rect 271 582 280 583
rect 298 587 304 588
rect 298 583 299 587
rect 303 583 304 587
rect 298 582 304 583
rect 350 587 356 588
rect 350 583 351 587
rect 355 586 356 587
rect 359 587 365 588
rect 359 586 360 587
rect 355 584 360 586
rect 355 583 356 584
rect 350 582 356 583
rect 359 583 360 584
rect 364 583 365 587
rect 359 582 365 583
rect 386 587 392 588
rect 386 583 387 587
rect 391 583 392 587
rect 386 582 392 583
rect 404 582 406 596
rect 449 587 455 588
rect 449 583 450 587
rect 454 583 455 587
rect 449 582 455 583
rect 474 587 480 588
rect 474 583 475 587
rect 479 583 480 587
rect 474 582 480 583
rect 546 587 552 588
rect 546 583 547 587
rect 551 583 552 587
rect 546 582 552 583
rect 570 587 576 588
rect 570 583 571 587
rect 575 583 576 587
rect 570 582 576 583
rect 639 587 645 588
rect 639 583 640 587
rect 644 586 645 587
rect 650 587 656 588
rect 650 586 651 587
rect 644 584 651 586
rect 644 583 645 584
rect 639 582 645 583
rect 650 583 651 584
rect 655 583 656 587
rect 650 582 656 583
rect 666 587 672 588
rect 666 583 667 587
rect 671 583 672 587
rect 666 582 672 583
rect 679 582 681 596
rect 722 595 723 599
rect 727 595 728 599
rect 722 594 728 595
rect 774 599 780 600
rect 774 595 775 599
rect 779 595 780 599
rect 774 594 780 595
rect 721 587 727 588
rect 721 583 722 587
rect 726 583 727 587
rect 721 582 727 583
rect 746 587 752 588
rect 746 583 747 587
rect 751 583 752 587
rect 746 582 752 583
rect 404 580 451 582
rect 679 580 723 582
rect 145 571 152 572
rect 145 567 146 571
rect 151 567 152 571
rect 721 571 728 572
rect 145 566 152 567
rect 170 569 176 570
rect 170 565 171 569
rect 175 565 176 569
rect 226 569 232 570
rect 201 567 207 568
rect 201 566 202 567
rect 170 564 176 565
rect 180 564 202 566
rect 180 558 182 564
rect 201 563 202 564
rect 206 563 207 567
rect 226 565 227 569
rect 231 565 232 569
rect 322 569 328 570
rect 297 567 303 568
rect 297 566 298 567
rect 226 564 232 565
rect 244 564 298 566
rect 201 562 207 563
rect 244 558 246 564
rect 297 563 298 564
rect 302 563 303 567
rect 322 565 323 569
rect 327 565 328 569
rect 426 569 432 570
rect 401 567 407 568
rect 401 566 402 567
rect 322 564 328 565
rect 360 564 402 566
rect 297 562 303 563
rect 360 558 362 564
rect 401 563 402 564
rect 406 563 407 567
rect 426 565 427 569
rect 431 565 432 569
rect 538 569 544 570
rect 513 567 519 568
rect 513 566 514 567
rect 426 564 432 565
rect 452 564 514 566
rect 401 562 407 563
rect 452 558 454 564
rect 513 563 514 564
rect 518 563 519 567
rect 538 565 539 569
rect 543 565 544 569
rect 650 569 656 570
rect 538 564 544 565
rect 625 567 631 568
rect 513 562 519 563
rect 625 563 626 567
rect 630 566 631 567
rect 642 567 648 568
rect 642 566 643 567
rect 630 564 643 566
rect 630 563 631 564
rect 625 562 631 563
rect 642 563 643 564
rect 647 563 648 567
rect 650 565 651 569
rect 655 565 656 569
rect 721 567 722 571
rect 727 567 728 571
rect 721 566 728 567
rect 746 569 752 570
rect 650 564 656 565
rect 746 565 747 569
rect 751 565 752 569
rect 746 564 752 565
rect 642 562 648 563
rect 110 557 116 558
rect 110 553 111 557
rect 115 553 116 557
rect 153 556 182 558
rect 209 556 246 558
rect 305 556 362 558
rect 409 556 454 558
rect 774 557 780 558
rect 110 552 116 553
rect 546 555 552 556
rect 546 551 547 555
rect 551 554 552 555
rect 551 552 625 554
rect 774 553 775 557
rect 779 553 780 557
rect 774 552 780 553
rect 551 551 552 552
rect 546 550 552 551
rect 110 539 116 540
rect 110 535 111 539
rect 115 535 116 539
rect 110 534 116 535
rect 210 539 216 540
rect 210 535 211 539
rect 215 538 216 539
rect 774 539 780 540
rect 215 536 506 538
rect 215 535 216 536
rect 210 534 216 535
rect 146 531 152 532
rect 146 527 147 531
rect 151 527 152 531
rect 146 526 152 527
rect 202 531 208 532
rect 202 527 203 531
rect 207 527 208 531
rect 202 526 208 527
rect 298 531 304 532
rect 298 527 299 531
rect 303 527 304 531
rect 298 526 304 527
rect 402 531 408 532
rect 402 527 403 531
rect 407 527 408 531
rect 504 529 506 536
rect 774 535 775 539
rect 779 535 780 539
rect 774 534 780 535
rect 514 531 520 532
rect 402 526 408 527
rect 514 527 515 531
rect 519 527 520 531
rect 514 526 520 527
rect 626 531 632 532
rect 626 527 627 531
rect 631 527 632 531
rect 626 526 632 527
rect 703 531 709 532
rect 703 527 704 531
rect 708 530 709 531
rect 722 531 728 532
rect 708 528 713 530
rect 708 527 709 528
rect 703 526 709 527
rect 722 527 723 531
rect 727 527 728 531
rect 722 526 728 527
rect 194 521 200 522
rect 194 517 195 521
rect 199 517 200 521
rect 194 516 200 517
rect 282 521 288 522
rect 282 517 283 521
rect 287 517 288 521
rect 282 516 288 517
rect 378 521 384 522
rect 378 517 379 521
rect 383 517 384 521
rect 378 516 384 517
rect 490 521 496 522
rect 490 517 491 521
rect 495 517 496 521
rect 490 516 496 517
rect 610 521 616 522
rect 610 517 611 521
rect 615 517 616 521
rect 610 516 616 517
rect 722 521 728 522
rect 722 517 723 521
rect 727 517 728 521
rect 722 516 728 517
rect 110 513 116 514
rect 110 509 111 513
rect 115 509 116 513
rect 110 508 116 509
rect 774 513 780 514
rect 774 509 775 513
rect 779 509 780 513
rect 774 508 780 509
rect 110 495 116 496
rect 110 491 111 495
rect 115 491 116 495
rect 606 495 612 496
rect 201 492 238 494
rect 289 492 321 494
rect 385 492 434 494
rect 497 492 549 494
rect 110 490 116 491
rect 191 483 197 484
rect 191 479 192 483
rect 196 482 197 483
rect 210 483 216 484
rect 210 482 211 483
rect 196 480 211 482
rect 196 479 197 480
rect 191 478 197 479
rect 210 479 211 480
rect 215 479 216 483
rect 210 478 216 479
rect 218 483 224 484
rect 218 479 219 483
rect 223 479 224 483
rect 236 482 238 492
rect 279 483 285 484
rect 279 482 280 483
rect 236 480 280 482
rect 218 478 224 479
rect 279 479 280 480
rect 284 479 285 483
rect 279 478 285 479
rect 306 483 312 484
rect 306 479 307 483
rect 311 479 312 483
rect 319 482 321 492
rect 375 483 381 484
rect 375 482 376 483
rect 319 480 376 482
rect 306 478 312 479
rect 375 479 376 480
rect 380 479 381 483
rect 375 478 381 479
rect 402 483 408 484
rect 402 479 403 483
rect 407 479 408 483
rect 432 482 434 492
rect 487 483 493 484
rect 487 482 488 483
rect 432 480 488 482
rect 402 478 408 479
rect 487 479 488 480
rect 492 479 493 483
rect 487 478 493 479
rect 514 483 520 484
rect 514 479 515 483
rect 519 479 520 483
rect 547 482 549 492
rect 606 491 607 495
rect 611 491 612 495
rect 606 490 612 491
rect 722 495 728 496
rect 722 491 723 495
rect 727 491 728 495
rect 722 490 728 491
rect 774 495 780 496
rect 774 491 775 495
rect 779 491 780 495
rect 774 490 780 491
rect 607 483 613 484
rect 607 482 608 483
rect 547 480 608 482
rect 514 478 520 479
rect 607 479 608 480
rect 612 479 613 483
rect 607 478 613 479
rect 634 483 640 484
rect 634 479 635 483
rect 639 479 640 483
rect 634 478 640 479
rect 703 483 709 484
rect 703 479 704 483
rect 708 482 709 483
rect 719 483 725 484
rect 719 482 720 483
rect 708 480 720 482
rect 708 479 709 480
rect 703 478 709 479
rect 719 479 720 480
rect 724 479 725 483
rect 719 478 725 479
rect 746 483 752 484
rect 746 479 747 483
rect 751 479 752 483
rect 746 478 752 479
rect 606 475 612 476
rect 606 474 607 475
rect 319 472 607 474
rect 313 471 321 472
rect 313 467 314 471
rect 318 468 321 471
rect 606 471 607 472
rect 611 471 612 475
rect 606 470 612 471
rect 721 471 728 472
rect 338 469 344 470
rect 318 467 319 468
rect 313 466 319 467
rect 338 465 339 469
rect 343 465 344 469
rect 394 469 400 470
rect 369 467 375 468
rect 369 466 370 467
rect 338 464 344 465
rect 348 464 370 466
rect 348 458 350 464
rect 369 463 370 464
rect 374 463 375 467
rect 394 465 395 469
rect 399 465 400 469
rect 450 469 456 470
rect 425 467 431 468
rect 425 466 426 467
rect 394 464 400 465
rect 404 464 426 466
rect 369 462 375 463
rect 404 458 406 464
rect 425 463 426 464
rect 430 463 431 467
rect 450 465 451 469
rect 455 465 456 469
rect 514 469 520 470
rect 450 464 456 465
rect 489 467 495 468
rect 425 462 431 463
rect 489 463 490 467
rect 494 463 495 467
rect 514 465 515 469
rect 519 465 520 469
rect 586 469 592 470
rect 561 467 567 468
rect 561 466 562 467
rect 514 464 520 465
rect 524 464 562 466
rect 489 462 495 463
rect 452 460 493 462
rect 452 458 454 460
rect 524 458 526 464
rect 561 463 562 464
rect 566 463 567 467
rect 586 465 587 469
rect 591 465 592 469
rect 666 469 672 470
rect 586 464 592 465
rect 641 467 647 468
rect 561 462 567 463
rect 641 463 642 467
rect 646 466 647 467
rect 650 467 656 468
rect 650 466 651 467
rect 646 464 651 466
rect 646 463 647 464
rect 641 462 647 463
rect 650 463 651 464
rect 655 463 656 467
rect 666 465 667 469
rect 671 465 672 469
rect 721 467 722 471
rect 727 467 728 471
rect 721 466 728 467
rect 746 469 752 470
rect 666 464 672 465
rect 746 465 747 469
rect 751 465 752 469
rect 746 464 752 465
rect 650 462 656 463
rect 110 457 116 458
rect 110 453 111 457
rect 115 453 116 457
rect 321 456 350 458
rect 377 456 406 458
rect 433 456 454 458
rect 497 456 526 458
rect 642 459 648 460
rect 586 455 592 456
rect 586 454 587 455
rect 110 452 116 453
rect 569 452 587 454
rect 586 451 587 452
rect 591 451 592 455
rect 642 455 643 459
rect 647 455 648 459
rect 642 454 648 455
rect 774 457 780 458
rect 774 453 775 457
rect 779 453 780 457
rect 774 452 780 453
rect 586 450 592 451
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 110 434 116 435
rect 774 439 780 440
rect 774 435 775 439
rect 779 435 780 439
rect 774 434 780 435
rect 314 431 320 432
rect 314 427 315 431
rect 319 427 320 431
rect 314 426 320 427
rect 370 431 376 432
rect 370 427 371 431
rect 375 427 376 431
rect 370 426 376 427
rect 426 431 432 432
rect 426 427 427 431
rect 431 427 432 431
rect 426 426 432 427
rect 490 431 496 432
rect 490 427 491 431
rect 495 427 496 431
rect 490 426 496 427
rect 562 431 568 432
rect 562 427 563 431
rect 567 427 568 431
rect 562 426 568 427
rect 642 431 648 432
rect 642 427 643 431
rect 647 427 648 431
rect 642 426 648 427
rect 703 431 709 432
rect 703 427 704 431
rect 708 430 709 431
rect 722 431 728 432
rect 708 428 713 430
rect 708 427 709 428
rect 703 426 709 427
rect 722 427 723 431
rect 727 427 728 431
rect 722 426 728 427
rect 650 423 656 424
rect 650 419 651 423
rect 655 419 656 423
rect 650 418 656 419
rect 652 414 654 418
rect 386 413 392 414
rect 386 409 387 413
rect 391 409 392 413
rect 386 408 392 409
rect 442 413 448 414
rect 442 409 443 413
rect 447 409 448 413
rect 442 408 448 409
rect 498 413 504 414
rect 498 409 499 413
rect 503 409 504 413
rect 498 408 504 409
rect 554 413 560 414
rect 554 409 555 413
rect 559 409 560 413
rect 554 408 560 409
rect 610 413 616 414
rect 610 409 611 413
rect 615 409 616 413
rect 652 412 657 414
rect 666 413 672 414
rect 610 408 616 409
rect 666 409 667 413
rect 671 409 672 413
rect 666 408 672 409
rect 722 413 728 414
rect 722 409 723 413
rect 727 409 728 413
rect 722 408 728 409
rect 110 405 116 406
rect 110 401 111 405
rect 115 401 116 405
rect 110 400 116 401
rect 774 405 780 406
rect 774 401 775 405
rect 779 401 780 405
rect 774 400 780 401
rect 386 395 392 396
rect 386 391 387 395
rect 391 394 392 395
rect 391 392 498 394
rect 391 391 392 392
rect 386 390 392 391
rect 110 387 116 388
rect 110 383 111 387
rect 115 383 116 387
rect 430 387 436 388
rect 430 386 431 387
rect 393 384 431 386
rect 110 382 116 383
rect 430 383 431 384
rect 435 383 436 387
rect 458 387 464 388
rect 458 386 459 387
rect 449 384 459 386
rect 430 382 436 383
rect 458 383 459 384
rect 463 383 464 387
rect 496 385 498 392
rect 718 387 724 388
rect 458 382 464 383
rect 512 384 553 386
rect 568 384 609 386
rect 383 375 392 376
rect 383 371 384 375
rect 391 371 392 375
rect 383 370 392 371
rect 410 375 416 376
rect 410 371 411 375
rect 415 371 416 375
rect 410 370 416 371
rect 438 375 447 376
rect 438 371 439 375
rect 446 371 447 375
rect 438 370 447 371
rect 466 375 472 376
rect 466 371 467 375
rect 471 371 472 375
rect 466 370 472 371
rect 495 375 501 376
rect 495 371 496 375
rect 500 374 501 375
rect 512 374 514 384
rect 500 372 514 374
rect 522 375 528 376
rect 500 371 501 372
rect 495 370 501 371
rect 522 371 523 375
rect 527 371 528 375
rect 522 370 528 371
rect 551 375 557 376
rect 551 371 552 375
rect 556 374 557 375
rect 568 374 570 384
rect 718 383 719 387
rect 723 383 724 387
rect 718 382 724 383
rect 774 387 780 388
rect 774 383 775 387
rect 779 383 780 387
rect 774 382 780 383
rect 556 372 570 374
rect 578 375 584 376
rect 556 371 557 372
rect 551 370 557 371
rect 578 371 579 375
rect 583 371 584 375
rect 578 370 584 371
rect 586 375 592 376
rect 586 371 587 375
rect 591 374 592 375
rect 607 375 613 376
rect 607 374 608 375
rect 591 372 608 374
rect 591 371 592 372
rect 586 370 592 371
rect 607 371 608 372
rect 612 371 613 375
rect 607 370 613 371
rect 634 375 640 376
rect 634 371 635 375
rect 639 371 640 375
rect 634 370 640 371
rect 642 375 648 376
rect 642 371 643 375
rect 647 374 648 375
rect 663 375 669 376
rect 663 374 664 375
rect 647 372 664 374
rect 647 371 648 372
rect 642 370 648 371
rect 663 371 664 372
rect 668 371 669 375
rect 663 370 669 371
rect 690 375 696 376
rect 690 371 691 375
rect 695 371 696 375
rect 690 370 696 371
rect 703 375 709 376
rect 703 371 704 375
rect 708 374 709 375
rect 719 375 725 376
rect 719 374 720 375
rect 708 372 720 374
rect 708 371 709 372
rect 703 370 709 371
rect 719 371 720 372
rect 724 371 725 375
rect 719 370 725 371
rect 746 375 752 376
rect 746 371 747 375
rect 751 371 752 375
rect 746 370 752 371
rect 458 363 464 364
rect 322 361 328 362
rect 297 359 303 360
rect 297 355 298 359
rect 302 358 303 359
rect 310 359 316 360
rect 310 358 311 359
rect 302 356 311 358
rect 302 355 303 356
rect 297 354 303 355
rect 310 355 311 356
rect 315 355 316 359
rect 322 357 323 361
rect 327 357 328 361
rect 378 361 384 362
rect 353 359 359 360
rect 353 358 354 359
rect 322 356 328 357
rect 336 356 354 358
rect 310 354 316 355
rect 336 350 338 356
rect 353 355 354 356
rect 358 355 359 359
rect 378 357 379 361
rect 383 357 384 361
rect 434 361 440 362
rect 409 359 415 360
rect 409 358 410 359
rect 378 356 384 357
rect 388 356 410 358
rect 353 354 359 355
rect 388 350 390 356
rect 409 355 410 356
rect 414 355 415 359
rect 434 357 435 361
rect 439 357 440 361
rect 458 359 459 363
rect 463 362 464 363
rect 473 363 479 364
rect 473 362 474 363
rect 463 360 474 362
rect 463 359 464 360
rect 458 358 464 359
rect 473 359 474 360
rect 478 359 479 363
rect 713 363 724 364
rect 473 358 479 359
rect 498 361 504 362
rect 434 356 440 357
rect 498 357 499 361
rect 503 357 504 361
rect 570 361 576 362
rect 545 359 551 360
rect 545 358 546 359
rect 498 356 504 357
rect 508 356 546 358
rect 409 354 415 355
rect 508 350 510 356
rect 545 355 546 356
rect 550 355 551 359
rect 570 357 571 361
rect 575 357 576 361
rect 650 361 656 362
rect 570 356 576 357
rect 591 359 597 360
rect 545 354 551 355
rect 591 355 592 359
rect 596 358 597 359
rect 625 359 631 360
rect 625 358 626 359
rect 596 356 626 358
rect 596 355 597 356
rect 591 354 597 355
rect 625 355 626 356
rect 630 355 631 359
rect 650 357 651 361
rect 655 357 656 361
rect 713 359 714 363
rect 718 359 719 363
rect 723 359 724 363
rect 713 358 724 359
rect 738 361 744 362
rect 650 356 656 357
rect 738 357 739 361
rect 743 357 744 361
rect 738 356 744 357
rect 625 354 631 355
rect 642 351 648 352
rect 642 350 643 351
rect 110 349 116 350
rect 110 345 111 349
rect 115 345 116 349
rect 305 348 338 350
rect 361 348 390 350
rect 481 348 510 350
rect 633 348 643 350
rect 642 347 643 348
rect 647 347 648 351
rect 642 346 648 347
rect 774 349 780 350
rect 774 345 775 349
rect 779 345 780 349
rect 110 344 116 345
rect 310 343 316 344
rect 310 339 311 343
rect 315 342 316 343
rect 544 342 546 345
rect 774 344 780 345
rect 315 340 546 342
rect 315 339 316 340
rect 310 338 316 339
rect 110 331 116 332
rect 110 327 111 331
rect 115 327 116 331
rect 110 326 116 327
rect 774 331 780 332
rect 774 327 775 331
rect 779 327 780 331
rect 774 326 780 327
rect 298 323 304 324
rect 298 319 299 323
rect 303 319 304 323
rect 298 318 304 319
rect 354 323 360 324
rect 354 319 355 323
rect 359 319 360 323
rect 354 318 360 319
rect 391 323 397 324
rect 391 319 392 323
rect 396 322 397 323
rect 410 323 416 324
rect 396 320 401 322
rect 396 319 397 320
rect 391 318 397 319
rect 410 319 411 323
rect 415 319 416 323
rect 410 318 416 319
rect 474 323 480 324
rect 474 319 475 323
rect 479 319 480 323
rect 474 318 480 319
rect 546 323 552 324
rect 546 319 547 323
rect 551 319 552 323
rect 546 318 552 319
rect 626 323 632 324
rect 626 319 627 323
rect 631 319 632 323
rect 626 318 632 319
rect 695 323 701 324
rect 695 319 696 323
rect 700 322 701 323
rect 714 323 720 324
rect 700 320 705 322
rect 700 319 701 320
rect 695 318 701 319
rect 714 319 715 323
rect 719 319 720 323
rect 714 318 720 319
rect 591 307 597 308
rect 170 305 176 306
rect 170 301 171 305
rect 175 301 176 305
rect 170 300 176 301
rect 250 305 256 306
rect 250 301 251 305
rect 255 301 256 305
rect 250 300 256 301
rect 330 305 336 306
rect 330 301 331 305
rect 335 301 336 305
rect 330 300 336 301
rect 418 305 424 306
rect 418 301 419 305
rect 423 301 424 305
rect 418 300 424 301
rect 514 305 520 306
rect 514 301 515 305
rect 519 301 520 305
rect 591 303 592 307
rect 596 306 597 307
rect 596 304 601 306
rect 610 305 616 306
rect 596 303 597 304
rect 591 302 597 303
rect 514 300 520 301
rect 610 301 611 305
rect 615 301 616 305
rect 610 300 616 301
rect 714 305 720 306
rect 714 301 715 305
rect 719 301 720 305
rect 714 300 720 301
rect 110 297 116 298
rect 110 293 111 297
rect 115 293 116 297
rect 110 292 116 293
rect 774 297 780 298
rect 774 293 775 297
rect 779 293 780 297
rect 774 292 780 293
rect 186 287 192 288
rect 186 283 187 287
rect 191 286 192 287
rect 191 284 418 286
rect 191 283 192 284
rect 186 282 192 283
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 346 279 352 280
rect 346 278 347 279
rect 177 276 245 278
rect 257 276 321 278
rect 337 276 347 278
rect 110 274 116 275
rect 167 267 173 268
rect 167 263 168 267
rect 172 266 173 267
rect 186 267 192 268
rect 186 266 187 267
rect 172 264 187 266
rect 172 263 173 264
rect 167 262 173 263
rect 186 263 187 264
rect 191 263 192 267
rect 186 262 192 263
rect 194 267 200 268
rect 194 263 195 267
rect 199 263 200 267
rect 243 266 245 276
rect 249 267 255 268
rect 249 266 250 267
rect 243 264 250 266
rect 194 262 200 263
rect 249 263 250 264
rect 254 263 255 267
rect 249 262 255 263
rect 274 267 280 268
rect 274 263 275 267
rect 279 263 280 267
rect 319 266 321 276
rect 346 275 347 276
rect 351 275 352 279
rect 416 277 418 284
rect 622 279 628 280
rect 521 276 562 278
rect 346 274 352 275
rect 327 267 333 268
rect 327 266 328 267
rect 319 264 328 266
rect 274 262 280 263
rect 327 263 328 264
rect 332 263 333 267
rect 327 262 333 263
rect 354 267 360 268
rect 354 263 355 267
rect 359 263 360 267
rect 354 262 360 263
rect 391 267 397 268
rect 391 263 392 267
rect 396 266 397 267
rect 415 267 421 268
rect 415 266 416 267
rect 396 264 416 266
rect 396 263 397 264
rect 391 262 397 263
rect 415 263 416 264
rect 420 263 421 267
rect 415 262 421 263
rect 442 267 448 268
rect 442 263 443 267
rect 447 263 448 267
rect 442 262 448 263
rect 494 267 500 268
rect 494 263 495 267
rect 499 266 500 267
rect 511 267 517 268
rect 511 266 512 267
rect 499 264 512 266
rect 499 263 500 264
rect 494 262 500 263
rect 511 263 512 264
rect 516 263 517 267
rect 511 262 517 263
rect 538 267 544 268
rect 538 263 539 267
rect 543 263 544 267
rect 560 266 562 276
rect 622 275 623 279
rect 627 278 628 279
rect 774 279 780 280
rect 627 276 713 278
rect 627 275 628 276
rect 622 274 628 275
rect 774 275 775 279
rect 779 275 780 279
rect 774 274 780 275
rect 609 267 615 268
rect 609 266 610 267
rect 560 264 610 266
rect 538 262 544 263
rect 609 263 610 264
rect 614 263 615 267
rect 609 262 615 263
rect 634 267 640 268
rect 634 263 635 267
rect 639 263 640 267
rect 634 262 640 263
rect 695 267 701 268
rect 695 263 696 267
rect 700 266 701 267
rect 711 267 717 268
rect 711 266 712 267
rect 700 264 712 266
rect 700 263 701 264
rect 695 262 701 263
rect 711 263 712 264
rect 716 263 717 267
rect 711 262 717 263
rect 738 267 744 268
rect 738 263 739 267
rect 743 263 744 267
rect 738 262 744 263
rect 346 255 352 256
rect 170 253 176 254
rect 145 251 151 252
rect 145 247 146 251
rect 150 250 151 251
rect 150 248 166 250
rect 170 249 171 253
rect 175 249 176 253
rect 266 253 272 254
rect 170 248 176 249
rect 241 251 247 252
rect 150 247 151 248
rect 145 246 151 247
rect 110 241 116 242
rect 110 237 111 241
rect 115 237 116 241
rect 110 236 116 237
rect 164 238 166 248
rect 241 247 242 251
rect 246 250 247 251
rect 246 248 262 250
rect 266 249 267 253
rect 271 249 272 253
rect 346 251 347 255
rect 351 254 352 255
rect 361 255 367 256
rect 361 254 362 255
rect 351 252 362 254
rect 351 251 352 252
rect 346 250 352 251
rect 361 251 362 252
rect 366 251 367 255
rect 617 255 628 256
rect 361 250 367 251
rect 386 253 392 254
rect 266 248 272 249
rect 386 249 387 253
rect 391 249 392 253
rect 514 253 520 254
rect 386 248 392 249
rect 478 251 484 252
rect 246 247 247 248
rect 241 246 247 247
rect 260 238 262 248
rect 478 247 479 251
rect 483 250 484 251
rect 489 251 495 252
rect 489 250 490 251
rect 483 248 490 250
rect 483 247 484 248
rect 478 246 484 247
rect 489 247 490 248
rect 494 247 495 251
rect 514 249 515 253
rect 519 249 520 253
rect 617 251 618 255
rect 622 251 623 255
rect 627 251 628 255
rect 617 250 628 251
rect 642 253 648 254
rect 514 248 520 249
rect 642 249 643 253
rect 647 249 648 253
rect 746 253 752 254
rect 721 251 727 252
rect 721 250 722 251
rect 642 248 648 249
rect 656 248 722 250
rect 489 246 495 247
rect 494 243 500 244
rect 494 239 495 243
rect 499 239 500 243
rect 656 242 658 248
rect 721 247 722 248
rect 726 247 727 251
rect 746 249 747 253
rect 751 249 752 253
rect 746 248 752 249
rect 721 246 727 247
rect 625 240 658 242
rect 774 241 780 242
rect 494 238 500 239
rect 164 236 241 238
rect 260 236 361 238
rect 774 237 775 241
rect 779 237 780 241
rect 774 236 780 237
rect 110 223 116 224
rect 110 219 111 223
rect 115 219 116 223
rect 110 218 116 219
rect 774 223 780 224
rect 774 219 775 223
rect 779 219 780 223
rect 774 218 780 219
rect 127 215 133 216
rect 127 211 128 215
rect 132 214 133 215
rect 146 215 152 216
rect 132 212 137 214
rect 132 211 133 212
rect 127 210 133 211
rect 146 211 147 215
rect 151 211 152 215
rect 146 210 152 211
rect 242 215 248 216
rect 242 211 243 215
rect 247 211 248 215
rect 242 210 248 211
rect 362 215 368 216
rect 362 211 363 215
rect 367 211 368 215
rect 362 210 368 211
rect 490 215 496 216
rect 490 211 491 215
rect 495 211 496 215
rect 490 210 496 211
rect 618 215 624 216
rect 618 211 619 215
rect 623 211 624 215
rect 618 210 624 211
rect 703 215 709 216
rect 703 211 704 215
rect 708 214 709 215
rect 722 215 728 216
rect 708 212 713 214
rect 708 211 709 212
rect 703 210 709 211
rect 722 211 723 215
rect 727 211 728 215
rect 722 210 728 211
rect 478 203 484 204
rect 146 201 152 202
rect 146 197 147 201
rect 151 197 152 201
rect 146 196 152 197
rect 210 201 216 202
rect 210 197 211 201
rect 215 197 216 201
rect 210 196 216 197
rect 298 201 304 202
rect 298 197 299 201
rect 303 197 304 201
rect 298 196 304 197
rect 402 201 408 202
rect 402 197 403 201
rect 407 197 408 201
rect 478 199 479 203
rect 483 202 484 203
rect 483 200 497 202
rect 506 201 512 202
rect 483 199 484 200
rect 478 198 484 199
rect 402 196 408 197
rect 506 197 507 201
rect 511 197 512 201
rect 506 196 512 197
rect 618 201 624 202
rect 618 197 619 201
rect 623 197 624 201
rect 618 196 624 197
rect 722 201 728 202
rect 722 197 723 201
rect 727 197 728 201
rect 722 196 728 197
rect 110 193 116 194
rect 110 189 111 193
rect 115 189 116 193
rect 110 188 116 189
rect 774 193 780 194
rect 774 189 775 193
rect 779 189 780 193
rect 774 188 780 189
rect 110 175 116 176
rect 110 171 111 175
rect 115 171 116 175
rect 398 175 404 176
rect 153 172 182 174
rect 217 172 251 174
rect 305 172 362 174
rect 110 170 116 171
rect 127 163 133 164
rect 127 159 128 163
rect 132 162 133 163
rect 143 163 149 164
rect 143 162 144 163
rect 132 160 144 162
rect 132 159 133 160
rect 127 158 133 159
rect 143 159 144 160
rect 148 159 149 163
rect 143 158 149 159
rect 170 163 176 164
rect 170 159 171 163
rect 175 159 176 163
rect 180 162 182 172
rect 207 163 213 164
rect 207 162 208 163
rect 180 160 208 162
rect 170 158 176 159
rect 207 159 208 160
rect 212 159 213 163
rect 207 158 213 159
rect 234 163 240 164
rect 234 159 235 163
rect 239 159 240 163
rect 249 162 251 172
rect 295 163 301 164
rect 295 162 296 163
rect 249 160 296 162
rect 234 158 240 159
rect 295 159 296 160
rect 300 159 301 163
rect 295 158 301 159
rect 322 163 328 164
rect 322 159 323 163
rect 327 159 328 163
rect 360 162 362 172
rect 398 171 399 175
rect 403 171 404 175
rect 722 175 728 176
rect 398 170 404 171
rect 520 172 617 174
rect 399 163 405 164
rect 399 162 400 163
rect 360 160 400 162
rect 322 158 328 159
rect 399 159 400 160
rect 404 159 405 163
rect 399 158 405 159
rect 426 163 432 164
rect 426 159 427 163
rect 431 159 432 163
rect 426 158 432 159
rect 503 163 509 164
rect 503 159 504 163
rect 508 162 509 163
rect 520 162 522 172
rect 722 171 723 175
rect 727 171 728 175
rect 722 170 728 171
rect 774 175 780 176
rect 774 171 775 175
rect 779 171 780 175
rect 774 170 780 171
rect 508 160 522 162
rect 530 163 536 164
rect 508 159 509 160
rect 503 158 509 159
rect 530 159 531 163
rect 535 159 536 163
rect 530 158 536 159
rect 558 163 564 164
rect 558 159 559 163
rect 563 162 564 163
rect 615 163 621 164
rect 615 162 616 163
rect 563 160 616 162
rect 563 159 564 160
rect 558 158 564 159
rect 615 159 616 160
rect 620 159 621 163
rect 615 158 621 159
rect 642 163 648 164
rect 642 159 643 163
rect 647 159 648 163
rect 642 158 648 159
rect 703 163 709 164
rect 703 159 704 163
rect 708 162 709 163
rect 719 163 725 164
rect 719 162 720 163
rect 708 160 720 162
rect 708 159 709 160
rect 703 158 709 159
rect 719 159 720 160
rect 724 159 725 163
rect 719 158 725 159
rect 746 163 752 164
rect 746 159 747 163
rect 751 159 752 163
rect 746 158 752 159
rect 398 147 404 148
rect 398 146 399 147
rect 180 144 399 146
rect 161 143 167 144
rect 161 139 162 143
rect 166 142 167 143
rect 180 142 182 144
rect 398 143 399 144
rect 403 143 404 147
rect 398 142 404 143
rect 721 143 728 144
rect 166 140 182 142
rect 186 141 192 142
rect 166 139 167 140
rect 161 138 167 139
rect 186 137 187 141
rect 191 137 192 141
rect 242 141 248 142
rect 217 139 223 140
rect 217 138 218 139
rect 186 136 192 137
rect 196 136 218 138
rect 196 130 198 136
rect 217 135 218 136
rect 222 135 223 139
rect 242 137 243 141
rect 247 137 248 141
rect 298 141 304 142
rect 273 139 279 140
rect 273 138 274 139
rect 242 136 248 137
rect 252 136 274 138
rect 217 134 223 135
rect 252 130 254 136
rect 273 135 274 136
rect 278 135 279 139
rect 298 137 299 141
rect 303 137 304 141
rect 354 141 360 142
rect 329 139 335 140
rect 329 138 330 139
rect 298 136 304 137
rect 319 136 330 138
rect 273 134 279 135
rect 319 130 321 136
rect 329 135 330 136
rect 334 135 335 139
rect 354 137 355 141
rect 359 137 360 141
rect 410 141 416 142
rect 385 139 391 140
rect 385 138 386 139
rect 354 136 360 137
rect 363 136 386 138
rect 329 134 335 135
rect 363 130 365 136
rect 385 135 386 136
rect 390 135 391 139
rect 410 137 411 141
rect 415 137 416 141
rect 466 141 472 142
rect 441 139 447 140
rect 441 138 442 139
rect 410 136 416 137
rect 420 136 442 138
rect 385 134 391 135
rect 420 130 422 136
rect 441 135 442 136
rect 446 135 447 139
rect 466 137 467 141
rect 471 137 472 141
rect 522 141 528 142
rect 497 139 503 140
rect 497 138 498 139
rect 466 136 472 137
rect 476 136 498 138
rect 441 134 447 135
rect 476 130 478 136
rect 497 135 498 136
rect 502 135 503 139
rect 522 137 523 141
rect 527 137 528 141
rect 578 141 584 142
rect 553 139 559 140
rect 553 138 554 139
rect 522 136 528 137
rect 532 136 554 138
rect 497 134 503 135
rect 532 130 534 136
rect 553 135 554 136
rect 558 135 559 139
rect 578 137 579 141
rect 583 137 584 141
rect 634 141 640 142
rect 578 136 584 137
rect 609 139 615 140
rect 553 134 559 135
rect 609 135 610 139
rect 614 138 615 139
rect 614 136 630 138
rect 634 137 635 141
rect 639 137 640 141
rect 690 141 696 142
rect 634 136 640 137
rect 665 139 671 140
rect 614 135 615 136
rect 609 134 615 135
rect 110 129 116 130
rect 110 125 111 129
rect 115 125 116 129
rect 169 128 198 130
rect 225 128 254 130
rect 281 128 321 130
rect 337 128 365 130
rect 393 128 422 130
rect 449 128 478 130
rect 505 128 534 130
rect 558 131 564 132
rect 558 127 559 131
rect 563 127 564 131
rect 558 126 564 127
rect 628 126 630 136
rect 665 135 666 139
rect 670 138 671 139
rect 670 136 686 138
rect 690 137 691 141
rect 695 137 696 141
rect 721 139 722 143
rect 727 139 728 143
rect 721 138 728 139
rect 746 141 752 142
rect 690 136 696 137
rect 746 137 747 141
rect 751 137 752 141
rect 746 136 752 137
rect 670 135 671 136
rect 665 134 671 135
rect 684 126 686 136
rect 774 129 780 130
rect 110 124 116 125
rect 628 124 665 126
rect 684 124 721 126
rect 774 125 775 129
rect 779 125 780 129
rect 774 124 780 125
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 110 106 116 107
rect 774 111 780 112
rect 774 107 775 111
rect 779 107 780 111
rect 774 106 780 107
rect 162 103 168 104
rect 162 99 163 103
rect 167 99 168 103
rect 162 98 168 99
rect 218 103 224 104
rect 218 99 219 103
rect 223 99 224 103
rect 218 98 224 99
rect 274 103 280 104
rect 274 99 275 103
rect 279 99 280 103
rect 274 98 280 99
rect 330 103 336 104
rect 330 99 331 103
rect 335 99 336 103
rect 330 98 336 99
rect 386 103 392 104
rect 386 99 387 103
rect 391 99 392 103
rect 386 98 392 99
rect 442 103 448 104
rect 442 99 443 103
rect 447 99 448 103
rect 442 98 448 99
rect 498 103 504 104
rect 498 99 499 103
rect 503 99 504 103
rect 498 98 504 99
rect 554 103 560 104
rect 554 99 555 103
rect 559 99 560 103
rect 554 98 560 99
rect 610 103 616 104
rect 610 99 611 103
rect 615 99 616 103
rect 610 98 616 99
rect 666 103 672 104
rect 666 99 667 103
rect 671 99 672 103
rect 666 98 672 99
rect 722 103 728 104
rect 722 99 723 103
rect 727 99 728 103
rect 722 98 728 99
<< m3c >>
rect 147 837 151 841
rect 203 837 207 841
rect 259 837 263 841
rect 315 837 319 841
rect 371 837 375 841
rect 427 837 431 841
rect 483 837 487 841
rect 111 829 115 833
rect 775 829 779 833
rect 111 811 115 815
rect 191 811 195 815
rect 171 799 175 803
rect 199 799 202 803
rect 202 799 203 803
rect 227 799 231 803
rect 303 811 307 815
rect 283 799 287 803
rect 311 799 314 803
rect 314 799 315 803
rect 339 799 343 803
rect 415 811 419 815
rect 395 799 399 803
rect 423 799 426 803
rect 426 799 427 803
rect 451 799 455 803
rect 479 811 483 815
rect 775 811 779 815
rect 507 799 511 803
rect 479 783 483 787
rect 227 777 231 781
rect 283 777 287 781
rect 339 777 343 781
rect 395 777 399 781
rect 451 777 455 781
rect 111 765 115 769
rect 775 765 779 769
rect 111 747 115 751
rect 347 747 351 751
rect 203 739 207 743
rect 259 739 263 743
rect 315 739 319 743
rect 371 739 375 743
rect 775 747 779 751
rect 427 739 431 743
rect 339 729 343 733
rect 395 729 399 733
rect 451 729 455 733
rect 507 729 511 733
rect 563 729 567 733
rect 111 721 115 725
rect 775 721 779 725
rect 443 711 447 715
rect 111 703 115 707
rect 383 703 387 707
rect 775 703 779 707
rect 347 691 351 695
rect 363 691 367 695
rect 387 691 391 695
rect 419 691 423 695
rect 475 691 479 695
rect 531 691 535 695
rect 587 691 591 695
rect 235 679 239 683
rect 243 681 247 685
rect 299 681 303 685
rect 355 681 359 685
rect 411 681 415 685
rect 443 683 446 687
rect 446 683 447 687
rect 467 681 471 685
rect 507 679 511 683
rect 523 681 527 685
rect 111 669 115 673
rect 351 667 355 671
rect 579 681 583 685
rect 635 681 639 685
rect 691 681 695 685
rect 747 681 751 685
rect 235 659 239 663
rect 775 669 779 673
rect 111 651 115 655
rect 775 651 779 655
rect 219 643 223 647
rect 275 643 279 647
rect 331 643 335 647
rect 387 643 391 647
rect 443 643 447 647
rect 499 643 503 647
rect 555 643 559 647
rect 611 643 615 647
rect 667 643 671 647
rect 651 635 655 639
rect 723 643 727 647
rect 147 621 151 625
rect 203 621 207 625
rect 275 621 279 625
rect 363 621 367 625
rect 451 621 455 625
rect 507 623 511 627
rect 547 621 551 625
rect 643 621 647 625
rect 723 621 727 625
rect 111 613 115 617
rect 775 613 779 617
rect 275 603 279 607
rect 111 595 115 599
rect 147 595 151 599
rect 171 583 175 587
rect 227 583 231 587
rect 275 583 276 587
rect 276 583 279 587
rect 299 583 303 587
rect 351 583 355 587
rect 387 583 391 587
rect 475 583 479 587
rect 547 583 551 587
rect 571 583 575 587
rect 651 583 655 587
rect 667 583 671 587
rect 723 595 727 599
rect 775 595 779 599
rect 747 583 751 587
rect 147 567 150 571
rect 150 567 151 571
rect 171 565 175 569
rect 227 565 231 569
rect 323 565 327 569
rect 427 565 431 569
rect 539 565 543 569
rect 643 563 647 567
rect 651 565 655 569
rect 723 567 726 571
rect 726 567 727 571
rect 747 565 751 569
rect 111 553 115 557
rect 547 551 551 555
rect 775 553 779 557
rect 111 535 115 539
rect 211 535 215 539
rect 147 527 151 531
rect 203 527 207 531
rect 299 527 303 531
rect 403 527 407 531
rect 775 535 779 539
rect 515 527 519 531
rect 627 527 631 531
rect 723 527 727 531
rect 195 517 199 521
rect 283 517 287 521
rect 379 517 383 521
rect 491 517 495 521
rect 611 517 615 521
rect 723 517 727 521
rect 111 509 115 513
rect 775 509 779 513
rect 111 491 115 495
rect 211 479 215 483
rect 219 479 223 483
rect 307 479 311 483
rect 403 479 407 483
rect 515 479 519 483
rect 607 491 611 495
rect 723 491 727 495
rect 775 491 779 495
rect 635 479 639 483
rect 747 479 751 483
rect 607 471 611 475
rect 339 465 343 469
rect 395 465 399 469
rect 451 465 455 469
rect 515 465 519 469
rect 587 465 591 469
rect 651 463 655 467
rect 667 465 671 469
rect 723 467 726 471
rect 726 467 727 471
rect 747 465 751 469
rect 111 453 115 457
rect 587 451 591 455
rect 643 455 647 459
rect 775 453 779 457
rect 111 435 115 439
rect 775 435 779 439
rect 315 427 319 431
rect 371 427 375 431
rect 427 427 431 431
rect 491 427 495 431
rect 563 427 567 431
rect 643 427 647 431
rect 723 427 727 431
rect 651 419 655 423
rect 387 409 391 413
rect 443 409 447 413
rect 499 409 503 413
rect 555 409 559 413
rect 611 409 615 413
rect 667 409 671 413
rect 723 409 727 413
rect 111 401 115 405
rect 775 401 779 405
rect 387 391 391 395
rect 111 383 115 387
rect 431 383 435 387
rect 459 383 463 387
rect 387 371 388 375
rect 388 371 391 375
rect 411 371 415 375
rect 439 371 442 375
rect 442 371 443 375
rect 467 371 471 375
rect 523 371 527 375
rect 719 383 723 387
rect 775 383 779 387
rect 579 371 583 375
rect 587 371 591 375
rect 635 371 639 375
rect 643 371 647 375
rect 691 371 695 375
rect 747 371 751 375
rect 311 355 315 359
rect 323 357 327 361
rect 379 357 383 361
rect 435 357 439 361
rect 459 359 463 363
rect 499 357 503 361
rect 571 357 575 361
rect 651 357 655 361
rect 719 359 723 363
rect 739 357 743 361
rect 111 345 115 349
rect 643 347 647 351
rect 775 345 779 349
rect 311 339 315 343
rect 111 327 115 331
rect 775 327 779 331
rect 299 319 303 323
rect 355 319 359 323
rect 411 319 415 323
rect 475 319 479 323
rect 547 319 551 323
rect 627 319 631 323
rect 715 319 719 323
rect 171 301 175 305
rect 251 301 255 305
rect 331 301 335 305
rect 419 301 423 305
rect 515 301 519 305
rect 611 301 615 305
rect 715 301 719 305
rect 111 293 115 297
rect 775 293 779 297
rect 187 283 191 287
rect 111 275 115 279
rect 187 263 191 267
rect 195 263 199 267
rect 275 263 279 267
rect 347 275 351 279
rect 355 263 359 267
rect 443 263 447 267
rect 495 263 499 267
rect 539 263 543 267
rect 623 275 627 279
rect 775 275 779 279
rect 635 263 639 267
rect 739 263 743 267
rect 171 249 175 253
rect 111 237 115 241
rect 267 249 271 253
rect 347 251 351 255
rect 387 249 391 253
rect 479 247 483 251
rect 515 249 519 253
rect 623 251 627 255
rect 643 249 647 253
rect 495 239 499 243
rect 747 249 751 253
rect 775 237 779 241
rect 111 219 115 223
rect 775 219 779 223
rect 147 211 151 215
rect 243 211 247 215
rect 363 211 367 215
rect 491 211 495 215
rect 619 211 623 215
rect 723 211 727 215
rect 147 197 151 201
rect 211 197 215 201
rect 299 197 303 201
rect 403 197 407 201
rect 479 199 483 203
rect 507 197 511 201
rect 619 197 623 201
rect 723 197 727 201
rect 111 189 115 193
rect 775 189 779 193
rect 111 171 115 175
rect 171 159 175 163
rect 235 159 239 163
rect 323 159 327 163
rect 399 171 403 175
rect 427 159 431 163
rect 723 171 727 175
rect 775 171 779 175
rect 531 159 535 163
rect 559 159 563 163
rect 643 159 647 163
rect 747 159 751 163
rect 399 143 403 147
rect 187 137 191 141
rect 243 137 247 141
rect 299 137 303 141
rect 355 137 359 141
rect 411 137 415 141
rect 467 137 471 141
rect 523 137 527 141
rect 579 137 583 141
rect 635 137 639 141
rect 111 125 115 129
rect 559 127 563 131
rect 691 137 695 141
rect 723 139 726 143
rect 726 139 727 143
rect 747 137 751 141
rect 775 125 779 129
rect 111 107 115 111
rect 775 107 779 111
rect 163 99 167 103
rect 219 99 223 103
rect 275 99 279 103
rect 331 99 335 103
rect 387 99 391 103
rect 443 99 447 103
rect 499 99 503 103
rect 555 99 559 103
rect 611 99 615 103
rect 667 99 671 103
rect 723 99 727 103
<< m3 >>
rect 111 846 115 847
rect 147 846 151 847
rect 203 846 207 847
rect 259 846 263 847
rect 315 846 319 847
rect 371 846 375 847
rect 427 846 431 847
rect 483 846 487 847
rect 775 846 779 847
rect 111 841 115 842
rect 146 841 152 842
rect 112 834 114 841
rect 146 837 147 841
rect 151 837 152 841
rect 146 836 152 837
rect 202 841 208 842
rect 202 837 203 841
rect 207 837 208 841
rect 202 836 208 837
rect 258 841 264 842
rect 258 837 259 841
rect 263 837 264 841
rect 258 836 264 837
rect 314 841 320 842
rect 314 837 315 841
rect 319 837 320 841
rect 314 836 320 837
rect 370 841 376 842
rect 370 837 371 841
rect 375 837 376 841
rect 370 836 376 837
rect 426 841 432 842
rect 426 837 427 841
rect 431 837 432 841
rect 426 836 432 837
rect 482 841 488 842
rect 775 841 779 842
rect 482 837 483 841
rect 487 837 488 841
rect 482 836 488 837
rect 776 834 778 841
rect 110 833 116 834
rect 110 829 111 833
rect 115 829 116 833
rect 110 828 116 829
rect 774 833 780 834
rect 774 829 775 833
rect 779 829 780 833
rect 774 828 780 829
rect 110 815 116 816
rect 110 811 111 815
rect 115 811 116 815
rect 110 810 116 811
rect 190 815 196 816
rect 190 811 191 815
rect 195 814 196 815
rect 302 815 308 816
rect 195 812 202 814
rect 195 811 196 812
rect 190 810 196 811
rect 112 787 114 810
rect 200 804 202 812
rect 302 811 303 815
rect 307 814 308 815
rect 414 815 420 816
rect 307 812 314 814
rect 307 811 308 812
rect 302 810 308 811
rect 312 804 314 812
rect 414 811 415 815
rect 419 814 420 815
rect 478 815 484 816
rect 419 812 426 814
rect 419 811 420 812
rect 414 810 420 811
rect 424 804 426 812
rect 478 811 479 815
rect 483 811 484 815
rect 478 810 484 811
rect 774 815 780 816
rect 774 811 775 815
rect 779 811 780 815
rect 774 810 780 811
rect 170 803 176 804
rect 170 799 171 803
rect 175 799 176 803
rect 170 798 176 799
rect 198 803 204 804
rect 198 799 199 803
rect 203 799 204 803
rect 198 798 204 799
rect 226 803 232 804
rect 226 799 227 803
rect 231 799 232 803
rect 226 798 232 799
rect 282 803 288 804
rect 282 799 283 803
rect 287 799 288 803
rect 282 798 288 799
rect 310 803 316 804
rect 310 799 311 803
rect 315 799 316 803
rect 310 798 316 799
rect 338 803 344 804
rect 338 799 339 803
rect 343 799 344 803
rect 338 798 344 799
rect 394 803 400 804
rect 394 799 395 803
rect 399 799 400 803
rect 394 798 400 799
rect 422 803 428 804
rect 422 799 423 803
rect 427 799 428 803
rect 422 798 428 799
rect 450 803 456 804
rect 450 799 451 803
rect 455 799 456 803
rect 450 798 456 799
rect 172 787 174 798
rect 228 787 230 798
rect 284 787 286 798
rect 340 787 342 798
rect 396 787 398 798
rect 452 787 454 798
rect 480 788 482 810
rect 506 803 512 804
rect 506 799 507 803
rect 511 799 512 803
rect 506 798 512 799
rect 478 787 484 788
rect 508 787 510 798
rect 776 787 778 810
rect 111 786 115 787
rect 111 781 115 782
rect 171 786 175 787
rect 227 786 231 787
rect 283 786 287 787
rect 339 786 343 787
rect 395 786 399 787
rect 451 786 455 787
rect 478 783 479 787
rect 483 783 484 787
rect 478 782 484 783
rect 507 786 511 787
rect 171 781 175 782
rect 226 781 232 782
rect 112 770 114 781
rect 226 777 227 781
rect 231 777 232 781
rect 226 776 232 777
rect 282 781 288 782
rect 282 777 283 781
rect 287 777 288 781
rect 282 776 288 777
rect 338 781 344 782
rect 338 777 339 781
rect 343 777 344 781
rect 338 776 344 777
rect 394 781 400 782
rect 394 777 395 781
rect 399 777 400 781
rect 394 776 400 777
rect 450 781 456 782
rect 507 781 511 782
rect 775 786 779 787
rect 775 781 779 782
rect 450 777 451 781
rect 455 777 456 781
rect 450 776 456 777
rect 776 770 778 781
rect 110 769 116 770
rect 110 765 111 769
rect 115 765 116 769
rect 110 764 116 765
rect 774 769 780 770
rect 774 765 775 769
rect 779 765 780 769
rect 774 764 780 765
rect 110 751 116 752
rect 110 747 111 751
rect 115 747 116 751
rect 110 746 116 747
rect 346 751 352 752
rect 346 747 347 751
rect 351 747 352 751
rect 346 746 352 747
rect 774 751 780 752
rect 774 747 775 751
rect 779 747 780 751
rect 774 746 780 747
rect 112 739 114 746
rect 202 743 208 744
rect 202 739 203 743
rect 207 739 208 743
rect 111 738 115 739
rect 202 738 208 739
rect 258 743 264 744
rect 258 739 259 743
rect 263 739 264 743
rect 258 738 264 739
rect 314 743 320 744
rect 314 739 315 743
rect 319 739 320 743
rect 314 738 320 739
rect 339 738 343 739
rect 111 733 115 734
rect 203 733 207 734
rect 259 733 263 734
rect 315 733 319 734
rect 338 733 344 734
rect 112 726 114 733
rect 338 729 339 733
rect 343 729 344 733
rect 338 728 344 729
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 110 720 116 721
rect 110 707 116 708
rect 110 703 111 707
rect 115 703 116 707
rect 110 702 116 703
rect 112 691 114 702
rect 348 696 350 746
rect 370 743 376 744
rect 370 739 371 743
rect 375 739 376 743
rect 426 743 432 744
rect 426 739 427 743
rect 431 739 432 743
rect 776 739 778 746
rect 370 738 376 739
rect 395 738 399 739
rect 426 738 432 739
rect 451 738 455 739
rect 507 738 511 739
rect 563 738 567 739
rect 775 738 779 739
rect 371 733 375 734
rect 394 733 400 734
rect 427 733 431 734
rect 450 733 456 734
rect 394 729 395 733
rect 399 729 400 733
rect 394 728 400 729
rect 450 729 451 733
rect 455 729 456 733
rect 450 728 456 729
rect 506 733 512 734
rect 506 729 507 733
rect 511 729 512 733
rect 506 728 512 729
rect 562 733 568 734
rect 775 733 779 734
rect 562 729 563 733
rect 567 729 568 733
rect 562 728 568 729
rect 776 726 778 733
rect 774 725 780 726
rect 774 721 775 725
rect 779 721 780 725
rect 774 720 780 721
rect 442 715 448 716
rect 442 711 443 715
rect 447 711 448 715
rect 442 710 448 711
rect 382 707 388 708
rect 382 703 383 707
rect 387 703 388 707
rect 382 702 388 703
rect 384 696 386 702
rect 346 695 352 696
rect 346 691 347 695
rect 351 691 352 695
rect 362 695 368 696
rect 362 691 363 695
rect 367 691 368 695
rect 384 695 392 696
rect 384 692 387 695
rect 111 690 115 691
rect 243 690 247 691
rect 299 690 303 691
rect 346 690 352 691
rect 355 690 359 691
rect 362 690 368 691
rect 386 691 387 692
rect 391 691 392 695
rect 418 695 424 696
rect 418 691 419 695
rect 423 691 424 695
rect 386 690 392 691
rect 411 690 415 691
rect 418 690 424 691
rect 444 688 446 710
rect 774 707 780 708
rect 774 703 775 707
rect 779 703 780 707
rect 774 702 780 703
rect 474 695 480 696
rect 474 691 475 695
rect 479 691 480 695
rect 530 695 536 696
rect 530 691 531 695
rect 535 691 536 695
rect 586 695 592 696
rect 586 691 587 695
rect 591 691 592 695
rect 776 691 778 702
rect 467 690 471 691
rect 474 690 480 691
rect 523 690 527 691
rect 530 690 536 691
rect 579 690 583 691
rect 586 690 592 691
rect 635 690 639 691
rect 111 685 115 686
rect 242 685 248 686
rect 112 674 114 685
rect 234 683 240 684
rect 234 679 235 683
rect 239 679 240 683
rect 242 681 243 685
rect 247 681 248 685
rect 242 680 248 681
rect 298 685 304 686
rect 298 681 299 685
rect 303 681 304 685
rect 298 680 304 681
rect 354 685 360 686
rect 363 685 367 686
rect 410 685 416 686
rect 419 685 423 686
rect 442 687 448 688
rect 354 681 355 685
rect 359 681 360 685
rect 354 680 360 681
rect 410 681 411 685
rect 415 681 416 685
rect 442 683 443 687
rect 447 683 448 687
rect 691 690 695 691
rect 747 690 751 691
rect 775 690 779 691
rect 442 682 448 683
rect 466 685 472 686
rect 475 685 479 686
rect 522 685 528 686
rect 531 685 535 686
rect 578 685 584 686
rect 587 685 591 686
rect 634 685 640 686
rect 410 680 416 681
rect 466 681 467 685
rect 471 681 472 685
rect 466 680 472 681
rect 506 683 512 684
rect 234 678 240 679
rect 506 679 507 683
rect 511 679 512 683
rect 522 681 523 685
rect 527 681 528 685
rect 522 680 528 681
rect 578 681 579 685
rect 583 681 584 685
rect 578 680 584 681
rect 634 681 635 685
rect 639 681 640 685
rect 634 680 640 681
rect 690 685 696 686
rect 690 681 691 685
rect 695 681 696 685
rect 690 680 696 681
rect 746 685 752 686
rect 775 685 779 686
rect 746 681 747 685
rect 751 681 752 685
rect 746 680 752 681
rect 506 678 512 679
rect 110 673 116 674
rect 110 669 111 673
rect 115 669 116 673
rect 110 668 116 669
rect 236 664 238 678
rect 350 671 356 672
rect 350 667 351 671
rect 355 667 356 671
rect 350 666 356 667
rect 234 663 240 664
rect 234 659 235 663
rect 239 659 240 663
rect 234 658 240 659
rect 110 655 116 656
rect 110 651 111 655
rect 115 651 116 655
rect 110 650 116 651
rect 112 631 114 650
rect 218 647 224 648
rect 218 643 219 647
rect 223 643 224 647
rect 218 642 224 643
rect 274 647 280 648
rect 274 643 275 647
rect 279 643 280 647
rect 274 642 280 643
rect 330 647 336 648
rect 330 643 331 647
rect 335 643 336 647
rect 330 642 336 643
rect 220 631 222 642
rect 276 631 278 642
rect 332 631 334 642
rect 111 630 115 631
rect 147 630 151 631
rect 203 630 207 631
rect 219 630 223 631
rect 275 630 279 631
rect 331 630 335 631
rect 111 625 115 626
rect 146 625 152 626
rect 112 618 114 625
rect 146 621 147 625
rect 151 621 152 625
rect 146 620 152 621
rect 202 625 208 626
rect 219 625 223 626
rect 274 625 280 626
rect 331 625 335 626
rect 202 621 203 625
rect 207 621 208 625
rect 202 620 208 621
rect 274 621 275 625
rect 279 621 280 625
rect 274 620 280 621
rect 110 617 116 618
rect 110 613 111 617
rect 115 613 116 617
rect 110 612 116 613
rect 274 607 280 608
rect 274 603 275 607
rect 279 603 280 607
rect 274 602 280 603
rect 110 599 116 600
rect 110 595 111 599
rect 115 595 116 599
rect 110 594 116 595
rect 146 599 152 600
rect 146 595 147 599
rect 151 595 152 599
rect 146 594 152 595
rect 112 575 114 594
rect 111 574 115 575
rect 148 572 150 594
rect 276 588 278 602
rect 352 588 354 666
rect 386 647 392 648
rect 386 643 387 647
rect 391 643 392 647
rect 386 642 392 643
rect 442 647 448 648
rect 442 643 443 647
rect 447 643 448 647
rect 442 642 448 643
rect 498 647 504 648
rect 498 643 499 647
rect 503 643 504 647
rect 498 642 504 643
rect 388 631 390 642
rect 444 631 446 642
rect 500 631 502 642
rect 363 630 367 631
rect 387 630 391 631
rect 362 625 368 626
rect 387 625 391 626
rect 443 630 447 631
rect 451 630 455 631
rect 499 630 503 631
rect 508 628 510 678
rect 776 674 778 685
rect 774 673 780 674
rect 774 669 775 673
rect 779 669 780 673
rect 774 668 780 669
rect 774 655 780 656
rect 774 651 775 655
rect 779 651 780 655
rect 774 650 780 651
rect 554 647 560 648
rect 554 643 555 647
rect 559 643 560 647
rect 554 642 560 643
rect 610 647 616 648
rect 610 643 611 647
rect 615 643 616 647
rect 610 642 616 643
rect 666 647 672 648
rect 666 643 667 647
rect 671 643 672 647
rect 666 642 672 643
rect 722 647 728 648
rect 722 643 723 647
rect 727 643 728 647
rect 722 642 728 643
rect 556 631 558 642
rect 612 631 614 642
rect 650 639 656 640
rect 650 635 651 639
rect 655 635 656 639
rect 650 634 656 635
rect 547 630 551 631
rect 443 625 447 626
rect 450 625 456 626
rect 499 625 503 626
rect 506 627 512 628
rect 362 621 363 625
rect 367 621 368 625
rect 362 620 368 621
rect 450 621 451 625
rect 455 621 456 625
rect 506 623 507 627
rect 511 623 512 627
rect 555 630 559 631
rect 506 622 512 623
rect 546 625 552 626
rect 555 625 559 626
rect 611 630 615 631
rect 643 630 647 631
rect 611 625 615 626
rect 642 625 648 626
rect 450 620 456 621
rect 546 621 547 625
rect 551 621 552 625
rect 546 620 552 621
rect 642 621 643 625
rect 647 621 648 625
rect 642 620 648 621
rect 652 588 654 634
rect 668 631 670 642
rect 724 631 726 642
rect 776 631 778 650
rect 667 630 671 631
rect 723 630 727 631
rect 775 630 779 631
rect 667 625 671 626
rect 722 625 728 626
rect 775 625 779 626
rect 722 621 723 625
rect 727 621 728 625
rect 722 620 728 621
rect 776 618 778 625
rect 774 617 780 618
rect 774 613 775 617
rect 779 613 780 617
rect 774 612 780 613
rect 722 599 728 600
rect 722 595 723 599
rect 727 595 728 599
rect 722 594 728 595
rect 774 599 780 600
rect 774 595 775 599
rect 779 595 780 599
rect 774 594 780 595
rect 170 587 176 588
rect 170 583 171 587
rect 175 583 176 587
rect 170 582 176 583
rect 226 587 232 588
rect 226 583 227 587
rect 231 583 232 587
rect 226 582 232 583
rect 274 587 280 588
rect 274 583 275 587
rect 279 583 280 587
rect 274 582 280 583
rect 298 587 304 588
rect 298 583 299 587
rect 303 583 304 587
rect 298 582 304 583
rect 350 587 356 588
rect 350 583 351 587
rect 355 583 356 587
rect 350 582 356 583
rect 386 587 392 588
rect 386 583 387 587
rect 391 583 392 587
rect 386 582 392 583
rect 474 587 480 588
rect 474 583 475 587
rect 479 583 480 587
rect 474 582 480 583
rect 546 587 552 588
rect 546 583 547 587
rect 551 583 552 587
rect 546 582 552 583
rect 570 587 576 588
rect 570 583 571 587
rect 575 583 576 587
rect 570 582 576 583
rect 650 587 656 588
rect 650 583 651 587
rect 655 583 656 587
rect 650 582 656 583
rect 666 587 672 588
rect 666 583 667 587
rect 671 583 672 587
rect 666 582 672 583
rect 172 575 174 582
rect 228 575 230 582
rect 300 575 302 582
rect 388 575 390 582
rect 476 575 478 582
rect 171 574 175 575
rect 111 569 115 570
rect 146 571 152 572
rect 112 558 114 569
rect 146 567 147 571
rect 151 567 152 571
rect 227 574 231 575
rect 299 574 303 575
rect 323 574 327 575
rect 387 574 391 575
rect 427 574 431 575
rect 475 574 479 575
rect 539 574 543 575
rect 146 566 152 567
rect 170 569 176 570
rect 170 565 171 569
rect 175 565 176 569
rect 170 564 176 565
rect 226 569 232 570
rect 299 569 303 570
rect 322 569 328 570
rect 387 569 391 570
rect 426 569 432 570
rect 475 569 479 570
rect 538 569 544 570
rect 226 565 227 569
rect 231 565 232 569
rect 226 564 232 565
rect 322 565 323 569
rect 327 565 328 569
rect 322 564 328 565
rect 426 565 427 569
rect 431 565 432 569
rect 426 564 432 565
rect 538 565 539 569
rect 543 565 544 569
rect 538 564 544 565
rect 110 557 116 558
rect 110 553 111 557
rect 115 553 116 557
rect 548 556 550 582
rect 572 575 574 582
rect 668 575 670 582
rect 571 574 575 575
rect 651 574 655 575
rect 667 574 671 575
rect 724 572 726 594
rect 746 587 752 588
rect 746 583 747 587
rect 751 583 752 587
rect 746 582 752 583
rect 748 575 750 582
rect 776 575 778 594
rect 747 574 751 575
rect 571 569 575 570
rect 650 569 656 570
rect 667 569 671 570
rect 722 571 728 572
rect 642 567 648 568
rect 642 563 643 567
rect 647 563 648 567
rect 650 565 651 569
rect 655 565 656 569
rect 722 567 723 571
rect 727 567 728 571
rect 775 574 779 575
rect 722 566 728 567
rect 746 569 752 570
rect 775 569 779 570
rect 650 564 656 565
rect 746 565 747 569
rect 751 565 752 569
rect 746 564 752 565
rect 642 562 648 563
rect 110 552 116 553
rect 546 555 552 556
rect 546 551 547 555
rect 551 551 552 555
rect 546 550 552 551
rect 110 539 116 540
rect 110 535 111 539
rect 115 535 116 539
rect 110 534 116 535
rect 210 539 216 540
rect 210 535 211 539
rect 215 535 216 539
rect 210 534 216 535
rect 112 527 114 534
rect 146 531 152 532
rect 146 527 147 531
rect 151 527 152 531
rect 202 531 208 532
rect 202 527 203 531
rect 207 527 208 531
rect 111 526 115 527
rect 146 526 152 527
rect 195 526 199 527
rect 202 526 208 527
rect 111 521 115 522
rect 147 521 151 522
rect 194 521 200 522
rect 203 521 207 522
rect 112 514 114 521
rect 194 517 195 521
rect 199 517 200 521
rect 194 516 200 517
rect 110 513 116 514
rect 110 509 111 513
rect 115 509 116 513
rect 110 508 116 509
rect 110 495 116 496
rect 110 491 111 495
rect 115 491 116 495
rect 110 490 116 491
rect 112 475 114 490
rect 212 484 214 534
rect 298 531 304 532
rect 298 527 299 531
rect 303 527 304 531
rect 402 531 408 532
rect 402 527 403 531
rect 407 527 408 531
rect 514 531 520 532
rect 514 527 515 531
rect 519 527 520 531
rect 626 531 632 532
rect 626 527 627 531
rect 631 527 632 531
rect 283 526 287 527
rect 298 526 304 527
rect 379 526 383 527
rect 402 526 408 527
rect 491 526 495 527
rect 514 526 520 527
rect 611 526 615 527
rect 626 526 632 527
rect 282 521 288 522
rect 299 521 303 522
rect 378 521 384 522
rect 403 521 407 522
rect 490 521 496 522
rect 515 521 519 522
rect 610 521 616 522
rect 627 521 631 522
rect 282 517 283 521
rect 287 517 288 521
rect 282 516 288 517
rect 378 517 379 521
rect 383 517 384 521
rect 378 516 384 517
rect 490 517 491 521
rect 495 517 496 521
rect 490 516 496 517
rect 610 517 611 521
rect 615 517 616 521
rect 610 516 616 517
rect 606 495 612 496
rect 606 491 607 495
rect 611 491 612 495
rect 606 490 612 491
rect 210 483 216 484
rect 210 479 211 483
rect 215 479 216 483
rect 210 478 216 479
rect 218 483 224 484
rect 218 479 219 483
rect 223 479 224 483
rect 218 478 224 479
rect 306 483 312 484
rect 306 479 307 483
rect 311 479 312 483
rect 306 478 312 479
rect 402 483 408 484
rect 402 479 403 483
rect 407 479 408 483
rect 402 478 408 479
rect 514 483 520 484
rect 514 479 515 483
rect 519 479 520 483
rect 514 478 520 479
rect 220 475 222 478
rect 308 475 310 478
rect 404 475 406 478
rect 516 475 518 478
rect 608 476 610 490
rect 634 483 640 484
rect 634 479 635 483
rect 639 479 640 483
rect 634 478 640 479
rect 606 475 612 476
rect 636 475 638 478
rect 111 474 115 475
rect 111 469 115 470
rect 219 474 223 475
rect 219 469 223 470
rect 307 474 311 475
rect 339 474 343 475
rect 395 474 399 475
rect 403 474 407 475
rect 451 474 455 475
rect 515 474 519 475
rect 587 474 591 475
rect 606 471 607 475
rect 611 471 612 475
rect 606 470 612 471
rect 635 474 639 475
rect 307 469 311 470
rect 338 469 344 470
rect 112 458 114 469
rect 338 465 339 469
rect 343 465 344 469
rect 338 464 344 465
rect 394 469 400 470
rect 403 469 407 470
rect 450 469 456 470
rect 394 465 395 469
rect 399 465 400 469
rect 394 464 400 465
rect 450 465 451 469
rect 455 465 456 469
rect 450 464 456 465
rect 514 469 520 470
rect 514 465 515 469
rect 519 465 520 469
rect 514 464 520 465
rect 586 469 592 470
rect 635 469 639 470
rect 586 465 587 469
rect 591 465 592 469
rect 586 464 592 465
rect 644 460 646 562
rect 776 558 778 569
rect 774 557 780 558
rect 774 553 775 557
rect 779 553 780 557
rect 774 552 780 553
rect 774 539 780 540
rect 774 535 775 539
rect 779 535 780 539
rect 774 534 780 535
rect 722 531 728 532
rect 722 527 723 531
rect 727 527 728 531
rect 776 527 778 534
rect 722 526 728 527
rect 775 526 779 527
rect 722 521 728 522
rect 775 521 779 522
rect 722 517 723 521
rect 727 517 728 521
rect 722 516 728 517
rect 776 514 778 521
rect 774 513 780 514
rect 774 509 775 513
rect 779 509 780 513
rect 774 508 780 509
rect 722 495 728 496
rect 722 491 723 495
rect 727 491 728 495
rect 722 490 728 491
rect 774 495 780 496
rect 774 491 775 495
rect 779 491 780 495
rect 774 490 780 491
rect 667 474 671 475
rect 724 472 726 490
rect 746 483 752 484
rect 746 479 747 483
rect 751 479 752 483
rect 746 478 752 479
rect 748 475 750 478
rect 776 475 778 490
rect 747 474 751 475
rect 722 471 728 472
rect 666 469 672 470
rect 650 467 656 468
rect 650 463 651 467
rect 655 463 656 467
rect 666 465 667 469
rect 671 465 672 469
rect 722 467 723 471
rect 727 467 728 471
rect 775 474 779 475
rect 722 466 728 467
rect 746 469 752 470
rect 775 469 779 470
rect 666 464 672 465
rect 746 465 747 469
rect 751 465 752 469
rect 746 464 752 465
rect 650 462 656 463
rect 642 459 648 460
rect 110 457 116 458
rect 110 453 111 457
rect 115 453 116 457
rect 110 452 116 453
rect 586 455 592 456
rect 586 451 587 455
rect 591 451 592 455
rect 642 455 643 459
rect 647 455 648 459
rect 642 454 648 455
rect 586 450 592 451
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 110 434 116 435
rect 112 419 114 434
rect 314 431 320 432
rect 314 427 315 431
rect 319 427 320 431
rect 314 426 320 427
rect 370 431 376 432
rect 370 427 371 431
rect 375 427 376 431
rect 370 426 376 427
rect 426 431 432 432
rect 426 427 427 431
rect 431 427 432 431
rect 426 426 432 427
rect 490 431 496 432
rect 490 427 491 431
rect 495 427 496 431
rect 490 426 496 427
rect 562 431 568 432
rect 562 427 563 431
rect 567 427 568 431
rect 562 426 568 427
rect 316 419 318 426
rect 372 419 374 426
rect 428 419 430 426
rect 492 419 494 426
rect 564 419 566 426
rect 111 418 115 419
rect 111 413 115 414
rect 315 418 319 419
rect 315 413 319 414
rect 371 418 375 419
rect 387 418 391 419
rect 427 418 431 419
rect 443 418 447 419
rect 491 418 495 419
rect 499 418 503 419
rect 555 418 559 419
rect 563 418 567 419
rect 371 413 375 414
rect 386 413 392 414
rect 427 413 431 414
rect 442 413 448 414
rect 491 413 495 414
rect 498 413 504 414
rect 112 406 114 413
rect 386 409 387 413
rect 391 409 392 413
rect 386 408 392 409
rect 442 409 443 413
rect 447 409 448 413
rect 442 408 448 409
rect 498 409 499 413
rect 503 409 504 413
rect 498 408 504 409
rect 554 413 560 414
rect 563 413 567 414
rect 554 409 555 413
rect 559 409 560 413
rect 554 408 560 409
rect 110 405 116 406
rect 110 401 111 405
rect 115 401 116 405
rect 110 400 116 401
rect 386 395 392 396
rect 386 391 387 395
rect 391 391 392 395
rect 386 390 392 391
rect 110 387 116 388
rect 110 383 111 387
rect 115 383 116 387
rect 110 382 116 383
rect 112 367 114 382
rect 388 376 390 390
rect 430 387 436 388
rect 430 383 431 387
rect 435 383 436 387
rect 430 382 436 383
rect 458 387 464 388
rect 458 383 459 387
rect 463 383 464 387
rect 458 382 464 383
rect 386 375 392 376
rect 386 371 387 375
rect 391 371 392 375
rect 386 370 392 371
rect 410 375 416 376
rect 410 371 411 375
rect 415 371 416 375
rect 432 374 434 382
rect 438 375 444 376
rect 438 374 439 375
rect 432 372 439 374
rect 410 370 416 371
rect 438 371 439 372
rect 443 371 444 375
rect 438 370 444 371
rect 412 367 414 370
rect 111 366 115 367
rect 323 366 327 367
rect 379 366 383 367
rect 411 366 415 367
rect 435 366 439 367
rect 460 364 462 382
rect 588 376 590 450
rect 642 431 648 432
rect 642 427 643 431
rect 647 427 648 431
rect 642 426 648 427
rect 644 419 646 426
rect 652 424 654 462
rect 776 458 778 469
rect 774 457 780 458
rect 774 453 775 457
rect 779 453 780 457
rect 774 452 780 453
rect 774 439 780 440
rect 774 435 775 439
rect 779 435 780 439
rect 774 434 780 435
rect 722 431 728 432
rect 722 427 723 431
rect 727 427 728 431
rect 722 426 728 427
rect 650 423 656 424
rect 650 419 651 423
rect 655 419 656 423
rect 724 419 726 426
rect 776 419 778 434
rect 611 418 615 419
rect 643 418 647 419
rect 650 418 656 419
rect 667 418 671 419
rect 723 418 727 419
rect 775 418 779 419
rect 610 413 616 414
rect 643 413 647 414
rect 666 413 672 414
rect 610 409 611 413
rect 615 409 616 413
rect 610 408 616 409
rect 666 409 667 413
rect 671 409 672 413
rect 666 408 672 409
rect 722 413 728 414
rect 775 413 779 414
rect 722 409 723 413
rect 727 409 728 413
rect 722 408 728 409
rect 776 406 778 413
rect 774 405 780 406
rect 774 401 775 405
rect 779 401 780 405
rect 774 400 780 401
rect 718 387 724 388
rect 718 383 719 387
rect 723 383 724 387
rect 718 382 724 383
rect 774 387 780 388
rect 774 383 775 387
rect 779 383 780 387
rect 774 382 780 383
rect 466 375 472 376
rect 466 371 467 375
rect 471 371 472 375
rect 466 370 472 371
rect 522 375 528 376
rect 522 371 523 375
rect 527 371 528 375
rect 522 370 528 371
rect 578 375 584 376
rect 578 371 579 375
rect 583 371 584 375
rect 578 370 584 371
rect 586 375 592 376
rect 586 371 587 375
rect 591 371 592 375
rect 586 370 592 371
rect 634 375 640 376
rect 634 371 635 375
rect 639 371 640 375
rect 634 370 640 371
rect 642 375 648 376
rect 642 371 643 375
rect 647 371 648 375
rect 642 370 648 371
rect 690 375 696 376
rect 690 371 691 375
rect 695 371 696 375
rect 690 370 696 371
rect 468 367 470 370
rect 524 367 526 370
rect 580 367 582 370
rect 636 367 638 370
rect 467 366 471 367
rect 458 363 464 364
rect 111 361 115 362
rect 322 361 328 362
rect 112 350 114 361
rect 310 359 316 360
rect 310 355 311 359
rect 315 355 316 359
rect 322 357 323 361
rect 327 357 328 361
rect 322 356 328 357
rect 378 361 384 362
rect 411 361 415 362
rect 434 361 440 362
rect 378 357 379 361
rect 383 357 384 361
rect 378 356 384 357
rect 434 357 435 361
rect 439 357 440 361
rect 458 359 459 363
rect 463 359 464 363
rect 499 366 503 367
rect 523 366 527 367
rect 571 366 575 367
rect 579 366 583 367
rect 467 361 471 362
rect 498 361 504 362
rect 523 361 527 362
rect 570 361 576 362
rect 579 361 583 362
rect 635 366 639 367
rect 635 361 639 362
rect 458 358 464 359
rect 434 356 440 357
rect 498 357 499 361
rect 503 357 504 361
rect 498 356 504 357
rect 570 357 571 361
rect 575 357 576 361
rect 570 356 576 357
rect 310 354 316 355
rect 110 349 116 350
rect 110 345 111 349
rect 115 345 116 349
rect 110 344 116 345
rect 312 344 314 354
rect 644 352 646 370
rect 692 367 694 370
rect 651 366 655 367
rect 691 366 695 367
rect 720 364 722 382
rect 746 375 752 376
rect 746 371 747 375
rect 751 371 752 375
rect 746 370 752 371
rect 748 367 750 370
rect 776 367 778 382
rect 739 366 743 367
rect 650 361 656 362
rect 691 361 695 362
rect 718 363 724 364
rect 650 357 651 361
rect 655 357 656 361
rect 718 359 719 363
rect 723 359 724 363
rect 747 366 751 367
rect 718 358 724 359
rect 738 361 744 362
rect 747 361 751 362
rect 775 366 779 367
rect 775 361 779 362
rect 650 356 656 357
rect 738 357 739 361
rect 743 357 744 361
rect 738 356 744 357
rect 642 351 648 352
rect 642 347 643 351
rect 647 347 648 351
rect 776 350 778 361
rect 642 346 648 347
rect 774 349 780 350
rect 774 345 775 349
rect 779 345 780 349
rect 774 344 780 345
rect 310 343 316 344
rect 310 339 311 343
rect 315 339 316 343
rect 310 338 316 339
rect 110 331 116 332
rect 110 327 111 331
rect 115 327 116 331
rect 110 326 116 327
rect 774 331 780 332
rect 774 327 775 331
rect 779 327 780 331
rect 774 326 780 327
rect 112 311 114 326
rect 298 323 304 324
rect 298 319 299 323
rect 303 319 304 323
rect 298 318 304 319
rect 354 323 360 324
rect 354 319 355 323
rect 359 319 360 323
rect 354 318 360 319
rect 410 323 416 324
rect 410 319 411 323
rect 415 319 416 323
rect 410 318 416 319
rect 474 323 480 324
rect 474 319 475 323
rect 479 319 480 323
rect 474 318 480 319
rect 546 323 552 324
rect 546 319 547 323
rect 551 319 552 323
rect 546 318 552 319
rect 626 323 632 324
rect 626 319 627 323
rect 631 319 632 323
rect 626 318 632 319
rect 714 323 720 324
rect 714 319 715 323
rect 719 319 720 323
rect 714 318 720 319
rect 300 311 302 318
rect 356 311 358 318
rect 412 311 414 318
rect 476 311 478 318
rect 548 311 550 318
rect 628 311 630 318
rect 716 311 718 318
rect 776 311 778 326
rect 111 310 115 311
rect 171 310 175 311
rect 251 310 255 311
rect 299 310 303 311
rect 331 310 335 311
rect 355 310 359 311
rect 111 305 115 306
rect 170 305 176 306
rect 112 298 114 305
rect 170 301 171 305
rect 175 301 176 305
rect 170 300 176 301
rect 250 305 256 306
rect 299 305 303 306
rect 330 305 336 306
rect 355 305 359 306
rect 411 310 415 311
rect 419 310 423 311
rect 475 310 479 311
rect 515 310 519 311
rect 547 310 551 311
rect 611 310 615 311
rect 627 310 631 311
rect 715 310 719 311
rect 775 310 779 311
rect 411 305 415 306
rect 418 305 424 306
rect 475 305 479 306
rect 514 305 520 306
rect 547 305 551 306
rect 610 305 616 306
rect 627 305 631 306
rect 714 305 720 306
rect 775 305 779 306
rect 250 301 251 305
rect 255 301 256 305
rect 250 300 256 301
rect 330 301 331 305
rect 335 301 336 305
rect 330 300 336 301
rect 418 301 419 305
rect 423 301 424 305
rect 418 300 424 301
rect 514 301 515 305
rect 519 301 520 305
rect 514 300 520 301
rect 610 301 611 305
rect 615 301 616 305
rect 610 300 616 301
rect 714 301 715 305
rect 719 301 720 305
rect 714 300 720 301
rect 776 298 778 305
rect 110 297 116 298
rect 110 293 111 297
rect 115 293 116 297
rect 110 292 116 293
rect 774 297 780 298
rect 774 293 775 297
rect 779 293 780 297
rect 774 292 780 293
rect 186 287 192 288
rect 186 283 187 287
rect 191 283 192 287
rect 186 282 192 283
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 110 274 116 275
rect 112 259 114 274
rect 188 268 190 282
rect 346 279 352 280
rect 346 275 347 279
rect 351 275 352 279
rect 346 274 352 275
rect 622 279 628 280
rect 622 275 623 279
rect 627 275 628 279
rect 622 274 628 275
rect 774 279 780 280
rect 774 275 775 279
rect 779 275 780 279
rect 774 274 780 275
rect 186 267 192 268
rect 186 263 187 267
rect 191 263 192 267
rect 186 262 192 263
rect 194 267 200 268
rect 194 263 195 267
rect 199 263 200 267
rect 194 262 200 263
rect 274 267 280 268
rect 274 263 275 267
rect 279 263 280 267
rect 274 262 280 263
rect 196 259 198 262
rect 276 259 278 262
rect 111 258 115 259
rect 171 258 175 259
rect 195 258 199 259
rect 267 258 271 259
rect 275 258 279 259
rect 348 256 350 274
rect 354 267 360 268
rect 354 263 355 267
rect 359 263 360 267
rect 354 262 360 263
rect 442 267 448 268
rect 442 263 443 267
rect 447 263 448 267
rect 442 262 448 263
rect 494 267 500 268
rect 494 263 495 267
rect 499 263 500 267
rect 494 262 500 263
rect 538 267 544 268
rect 538 263 539 267
rect 543 263 544 267
rect 538 262 544 263
rect 356 259 358 262
rect 444 259 446 262
rect 355 258 359 259
rect 111 253 115 254
rect 170 253 176 254
rect 195 253 199 254
rect 266 253 272 254
rect 275 253 279 254
rect 346 255 352 256
rect 112 242 114 253
rect 170 249 171 253
rect 175 249 176 253
rect 170 248 176 249
rect 266 249 267 253
rect 271 249 272 253
rect 346 251 347 255
rect 351 251 352 255
rect 387 258 391 259
rect 443 258 447 259
rect 355 253 359 254
rect 386 253 392 254
rect 443 253 447 254
rect 346 250 352 251
rect 266 248 272 249
rect 386 249 387 253
rect 391 249 392 253
rect 386 248 392 249
rect 478 251 484 252
rect 478 247 479 251
rect 483 247 484 251
rect 478 246 484 247
rect 110 241 116 242
rect 110 237 111 241
rect 115 237 116 241
rect 110 236 116 237
rect 110 223 116 224
rect 110 219 111 223
rect 115 219 116 223
rect 110 218 116 219
rect 112 207 114 218
rect 146 215 152 216
rect 146 211 147 215
rect 151 211 152 215
rect 146 210 152 211
rect 242 215 248 216
rect 242 211 243 215
rect 247 211 248 215
rect 242 210 248 211
rect 362 215 368 216
rect 362 211 363 215
rect 367 211 368 215
rect 362 210 368 211
rect 148 207 150 210
rect 244 207 246 210
rect 364 207 366 210
rect 111 206 115 207
rect 147 206 151 207
rect 211 206 215 207
rect 243 206 247 207
rect 299 206 303 207
rect 363 206 367 207
rect 403 206 407 207
rect 480 204 482 246
rect 496 244 498 262
rect 540 259 542 262
rect 515 258 519 259
rect 539 258 543 259
rect 624 256 626 274
rect 634 267 640 268
rect 634 263 635 267
rect 639 263 640 267
rect 634 262 640 263
rect 738 267 744 268
rect 738 263 739 267
rect 743 263 744 267
rect 738 262 744 263
rect 636 259 638 262
rect 740 259 742 262
rect 776 259 778 274
rect 635 258 639 259
rect 514 253 520 254
rect 539 253 543 254
rect 622 255 628 256
rect 514 249 515 253
rect 519 249 520 253
rect 622 251 623 255
rect 627 251 628 255
rect 643 258 647 259
rect 739 258 743 259
rect 747 258 751 259
rect 775 258 779 259
rect 635 253 639 254
rect 642 253 648 254
rect 739 253 743 254
rect 746 253 752 254
rect 775 253 779 254
rect 622 250 628 251
rect 514 248 520 249
rect 642 249 643 253
rect 647 249 648 253
rect 642 248 648 249
rect 746 249 747 253
rect 751 249 752 253
rect 746 248 752 249
rect 494 243 500 244
rect 494 239 495 243
rect 499 239 500 243
rect 776 242 778 253
rect 494 238 500 239
rect 774 241 780 242
rect 774 237 775 241
rect 779 237 780 241
rect 774 236 780 237
rect 774 223 780 224
rect 774 219 775 223
rect 779 219 780 223
rect 774 218 780 219
rect 490 215 496 216
rect 490 211 491 215
rect 495 211 496 215
rect 490 210 496 211
rect 618 215 624 216
rect 618 211 619 215
rect 623 211 624 215
rect 618 210 624 211
rect 722 215 728 216
rect 722 211 723 215
rect 727 211 728 215
rect 722 210 728 211
rect 492 207 494 210
rect 620 207 622 210
rect 724 207 726 210
rect 776 207 778 218
rect 491 206 495 207
rect 478 203 484 204
rect 111 201 115 202
rect 146 201 152 202
rect 112 194 114 201
rect 146 197 147 201
rect 151 197 152 201
rect 146 196 152 197
rect 210 201 216 202
rect 243 201 247 202
rect 298 201 304 202
rect 363 201 367 202
rect 402 201 408 202
rect 210 197 211 201
rect 215 197 216 201
rect 210 196 216 197
rect 298 197 299 201
rect 303 197 304 201
rect 298 196 304 197
rect 402 197 403 201
rect 407 197 408 201
rect 478 199 479 203
rect 483 199 484 203
rect 507 206 511 207
rect 619 206 623 207
rect 723 206 727 207
rect 775 206 779 207
rect 491 201 495 202
rect 506 201 512 202
rect 478 198 484 199
rect 402 196 408 197
rect 506 197 507 201
rect 511 197 512 201
rect 506 196 512 197
rect 618 201 624 202
rect 618 197 619 201
rect 623 197 624 201
rect 618 196 624 197
rect 722 201 728 202
rect 775 201 779 202
rect 722 197 723 201
rect 727 197 728 201
rect 722 196 728 197
rect 776 194 778 201
rect 110 193 116 194
rect 110 189 111 193
rect 115 189 116 193
rect 110 188 116 189
rect 774 193 780 194
rect 774 189 775 193
rect 779 189 780 193
rect 774 188 780 189
rect 110 175 116 176
rect 110 171 111 175
rect 115 171 116 175
rect 110 170 116 171
rect 398 175 404 176
rect 398 171 399 175
rect 403 171 404 175
rect 398 170 404 171
rect 722 175 728 176
rect 722 171 723 175
rect 727 171 728 175
rect 722 170 728 171
rect 774 175 780 176
rect 774 171 775 175
rect 779 171 780 175
rect 774 170 780 171
rect 112 147 114 170
rect 170 163 176 164
rect 170 159 171 163
rect 175 159 176 163
rect 170 158 176 159
rect 234 163 240 164
rect 234 159 235 163
rect 239 159 240 163
rect 234 158 240 159
rect 322 163 328 164
rect 322 159 323 163
rect 327 159 328 163
rect 322 158 328 159
rect 172 147 174 158
rect 236 147 238 158
rect 324 147 326 158
rect 400 148 402 170
rect 426 163 432 164
rect 426 159 427 163
rect 431 159 432 163
rect 426 158 432 159
rect 530 163 536 164
rect 530 159 531 163
rect 535 159 536 163
rect 530 158 536 159
rect 558 163 564 164
rect 558 159 559 163
rect 563 159 564 163
rect 558 158 564 159
rect 642 163 648 164
rect 642 159 643 163
rect 647 159 648 163
rect 642 158 648 159
rect 398 147 404 148
rect 428 147 430 158
rect 532 147 534 158
rect 111 146 115 147
rect 111 141 115 142
rect 171 146 175 147
rect 187 146 191 147
rect 235 146 239 147
rect 243 146 247 147
rect 299 146 303 147
rect 323 146 327 147
rect 355 146 359 147
rect 398 143 399 147
rect 403 143 404 147
rect 398 142 404 143
rect 411 146 415 147
rect 427 146 431 147
rect 467 146 471 147
rect 523 146 527 147
rect 531 146 535 147
rect 171 141 175 142
rect 186 141 192 142
rect 235 141 239 142
rect 242 141 248 142
rect 112 130 114 141
rect 186 137 187 141
rect 191 137 192 141
rect 186 136 192 137
rect 242 137 243 141
rect 247 137 248 141
rect 242 136 248 137
rect 298 141 304 142
rect 323 141 327 142
rect 354 141 360 142
rect 298 137 299 141
rect 303 137 304 141
rect 298 136 304 137
rect 354 137 355 141
rect 359 137 360 141
rect 354 136 360 137
rect 410 141 416 142
rect 427 141 431 142
rect 466 141 472 142
rect 410 137 411 141
rect 415 137 416 141
rect 410 136 416 137
rect 466 137 467 141
rect 471 137 472 141
rect 466 136 472 137
rect 522 141 528 142
rect 531 141 535 142
rect 522 137 523 141
rect 527 137 528 141
rect 522 136 528 137
rect 560 132 562 158
rect 644 147 646 158
rect 579 146 583 147
rect 635 146 639 147
rect 643 146 647 147
rect 691 146 695 147
rect 724 144 726 170
rect 746 163 752 164
rect 746 159 747 163
rect 751 159 752 163
rect 746 158 752 159
rect 748 147 750 158
rect 776 147 778 170
rect 747 146 751 147
rect 722 143 728 144
rect 578 141 584 142
rect 578 137 579 141
rect 583 137 584 141
rect 578 136 584 137
rect 634 141 640 142
rect 643 141 647 142
rect 690 141 696 142
rect 634 137 635 141
rect 639 137 640 141
rect 634 136 640 137
rect 690 137 691 141
rect 695 137 696 141
rect 722 139 723 143
rect 727 139 728 143
rect 775 146 779 147
rect 722 138 728 139
rect 746 141 752 142
rect 775 141 779 142
rect 690 136 696 137
rect 746 137 747 141
rect 751 137 752 141
rect 746 136 752 137
rect 558 131 564 132
rect 110 129 116 130
rect 110 125 111 129
rect 115 125 116 129
rect 558 127 559 131
rect 563 127 564 131
rect 776 130 778 141
rect 558 126 564 127
rect 774 129 780 130
rect 110 124 116 125
rect 774 125 775 129
rect 779 125 780 129
rect 774 124 780 125
rect 110 111 116 112
rect 110 107 111 111
rect 115 107 116 111
rect 110 106 116 107
rect 774 111 780 112
rect 774 107 775 111
rect 779 107 780 111
rect 774 106 780 107
rect 112 99 114 106
rect 162 103 168 104
rect 162 99 163 103
rect 167 99 168 103
rect 111 98 115 99
rect 162 98 168 99
rect 218 103 224 104
rect 218 99 219 103
rect 223 99 224 103
rect 218 98 224 99
rect 274 103 280 104
rect 274 99 275 103
rect 279 99 280 103
rect 274 98 280 99
rect 330 103 336 104
rect 330 99 331 103
rect 335 99 336 103
rect 330 98 336 99
rect 386 103 392 104
rect 386 99 387 103
rect 391 99 392 103
rect 386 98 392 99
rect 442 103 448 104
rect 442 99 443 103
rect 447 99 448 103
rect 442 98 448 99
rect 498 103 504 104
rect 498 99 499 103
rect 503 99 504 103
rect 498 98 504 99
rect 554 103 560 104
rect 554 99 555 103
rect 559 99 560 103
rect 554 98 560 99
rect 610 103 616 104
rect 610 99 611 103
rect 615 99 616 103
rect 610 98 616 99
rect 666 103 672 104
rect 666 99 667 103
rect 671 99 672 103
rect 666 98 672 99
rect 722 103 728 104
rect 722 99 723 103
rect 727 99 728 103
rect 776 99 778 106
rect 722 98 728 99
rect 775 98 779 99
rect 111 93 115 94
rect 163 93 167 94
rect 219 93 223 94
rect 275 93 279 94
rect 331 93 335 94
rect 387 93 391 94
rect 443 93 447 94
rect 499 93 503 94
rect 555 93 559 94
rect 611 93 615 94
rect 667 93 671 94
rect 723 93 727 94
rect 775 93 779 94
<< m4c >>
rect 111 842 115 846
rect 147 842 151 846
rect 203 842 207 846
rect 259 842 263 846
rect 315 842 319 846
rect 371 842 375 846
rect 427 842 431 846
rect 483 842 487 846
rect 775 842 779 846
rect 111 782 115 786
rect 171 782 175 786
rect 227 782 231 786
rect 283 782 287 786
rect 339 782 343 786
rect 395 782 399 786
rect 451 782 455 786
rect 507 782 511 786
rect 775 782 779 786
rect 111 734 115 738
rect 203 734 207 738
rect 259 734 263 738
rect 315 734 319 738
rect 339 734 343 738
rect 371 734 375 738
rect 395 734 399 738
rect 427 734 431 738
rect 451 734 455 738
rect 507 734 511 738
rect 563 734 567 738
rect 775 734 779 738
rect 111 686 115 690
rect 243 686 247 690
rect 299 686 303 690
rect 355 686 359 690
rect 363 686 367 690
rect 411 686 415 690
rect 419 686 423 690
rect 467 686 471 690
rect 475 686 479 690
rect 523 686 527 690
rect 531 686 535 690
rect 579 686 583 690
rect 587 686 591 690
rect 635 686 639 690
rect 691 686 695 690
rect 747 686 751 690
rect 775 686 779 690
rect 111 626 115 630
rect 147 626 151 630
rect 203 626 207 630
rect 219 626 223 630
rect 275 626 279 630
rect 331 626 335 630
rect 111 570 115 574
rect 363 626 367 630
rect 387 626 391 630
rect 443 626 447 630
rect 451 626 455 630
rect 499 626 503 630
rect 547 626 551 630
rect 555 626 559 630
rect 611 626 615 630
rect 643 626 647 630
rect 667 626 671 630
rect 723 626 727 630
rect 775 626 779 630
rect 171 570 175 574
rect 227 570 231 574
rect 299 570 303 574
rect 323 570 327 574
rect 387 570 391 574
rect 427 570 431 574
rect 475 570 479 574
rect 539 570 543 574
rect 571 570 575 574
rect 651 570 655 574
rect 667 570 671 574
rect 747 570 751 574
rect 775 570 779 574
rect 111 522 115 526
rect 147 522 151 526
rect 195 522 199 526
rect 203 522 207 526
rect 283 522 287 526
rect 299 522 303 526
rect 379 522 383 526
rect 403 522 407 526
rect 491 522 495 526
rect 515 522 519 526
rect 611 522 615 526
rect 627 522 631 526
rect 111 470 115 474
rect 219 470 223 474
rect 307 470 311 474
rect 339 470 343 474
rect 395 470 399 474
rect 403 470 407 474
rect 451 470 455 474
rect 515 470 519 474
rect 587 470 591 474
rect 635 470 639 474
rect 723 522 727 526
rect 775 522 779 526
rect 667 470 671 474
rect 747 470 751 474
rect 775 470 779 474
rect 111 414 115 418
rect 315 414 319 418
rect 371 414 375 418
rect 387 414 391 418
rect 427 414 431 418
rect 443 414 447 418
rect 491 414 495 418
rect 499 414 503 418
rect 555 414 559 418
rect 563 414 567 418
rect 111 362 115 366
rect 323 362 327 366
rect 379 362 383 366
rect 411 362 415 366
rect 435 362 439 366
rect 611 414 615 418
rect 643 414 647 418
rect 667 414 671 418
rect 723 414 727 418
rect 775 414 779 418
rect 467 362 471 366
rect 499 362 503 366
rect 523 362 527 366
rect 571 362 575 366
rect 579 362 583 366
rect 635 362 639 366
rect 651 362 655 366
rect 691 362 695 366
rect 739 362 743 366
rect 747 362 751 366
rect 775 362 779 366
rect 111 306 115 310
rect 171 306 175 310
rect 251 306 255 310
rect 299 306 303 310
rect 331 306 335 310
rect 355 306 359 310
rect 411 306 415 310
rect 419 306 423 310
rect 475 306 479 310
rect 515 306 519 310
rect 547 306 551 310
rect 611 306 615 310
rect 627 306 631 310
rect 715 306 719 310
rect 775 306 779 310
rect 111 254 115 258
rect 171 254 175 258
rect 195 254 199 258
rect 267 254 271 258
rect 275 254 279 258
rect 355 254 359 258
rect 387 254 391 258
rect 443 254 447 258
rect 111 202 115 206
rect 147 202 151 206
rect 211 202 215 206
rect 243 202 247 206
rect 299 202 303 206
rect 363 202 367 206
rect 403 202 407 206
rect 515 254 519 258
rect 539 254 543 258
rect 635 254 639 258
rect 643 254 647 258
rect 739 254 743 258
rect 747 254 751 258
rect 775 254 779 258
rect 491 202 495 206
rect 507 202 511 206
rect 619 202 623 206
rect 723 202 727 206
rect 775 202 779 206
rect 111 142 115 146
rect 171 142 175 146
rect 187 142 191 146
rect 235 142 239 146
rect 243 142 247 146
rect 299 142 303 146
rect 323 142 327 146
rect 355 142 359 146
rect 411 142 415 146
rect 427 142 431 146
rect 467 142 471 146
rect 523 142 527 146
rect 531 142 535 146
rect 579 142 583 146
rect 635 142 639 146
rect 643 142 647 146
rect 691 142 695 146
rect 747 142 751 146
rect 775 142 779 146
rect 111 94 115 98
rect 163 94 167 98
rect 219 94 223 98
rect 275 94 279 98
rect 331 94 335 98
rect 387 94 391 98
rect 443 94 447 98
rect 499 94 503 98
rect 555 94 559 98
rect 611 94 615 98
rect 667 94 671 98
rect 723 94 727 98
rect 775 94 779 98
<< m4 >>
rect 84 841 85 847
rect 91 846 799 847
rect 91 842 111 846
rect 115 842 147 846
rect 151 842 203 846
rect 207 842 259 846
rect 263 842 315 846
rect 319 842 371 846
rect 375 842 427 846
rect 431 842 483 846
rect 487 842 775 846
rect 779 842 799 846
rect 91 841 799 842
rect 805 841 806 847
rect 96 781 97 787
rect 103 786 811 787
rect 103 782 111 786
rect 115 782 171 786
rect 175 782 227 786
rect 231 782 283 786
rect 287 782 339 786
rect 343 782 395 786
rect 399 782 451 786
rect 455 782 507 786
rect 511 782 775 786
rect 779 782 811 786
rect 103 781 811 782
rect 817 781 818 787
rect 84 733 85 739
rect 91 738 799 739
rect 91 734 111 738
rect 115 734 203 738
rect 207 734 259 738
rect 263 734 315 738
rect 319 734 339 738
rect 343 734 371 738
rect 375 734 395 738
rect 399 734 427 738
rect 431 734 451 738
rect 455 734 507 738
rect 511 734 563 738
rect 567 734 775 738
rect 779 734 799 738
rect 91 733 799 734
rect 805 733 806 739
rect 96 685 97 691
rect 103 690 811 691
rect 103 686 111 690
rect 115 686 243 690
rect 247 686 299 690
rect 303 686 355 690
rect 359 686 363 690
rect 367 686 411 690
rect 415 686 419 690
rect 423 686 467 690
rect 471 686 475 690
rect 479 686 523 690
rect 527 686 531 690
rect 535 686 579 690
rect 583 686 587 690
rect 591 686 635 690
rect 639 686 691 690
rect 695 686 747 690
rect 751 686 775 690
rect 779 686 811 690
rect 103 685 811 686
rect 817 685 818 691
rect 84 625 85 631
rect 91 630 799 631
rect 91 626 111 630
rect 115 626 147 630
rect 151 626 203 630
rect 207 626 219 630
rect 223 626 275 630
rect 279 626 331 630
rect 335 626 363 630
rect 367 626 387 630
rect 391 626 443 630
rect 447 626 451 630
rect 455 626 499 630
rect 503 626 547 630
rect 551 626 555 630
rect 559 626 611 630
rect 615 626 643 630
rect 647 626 667 630
rect 671 626 723 630
rect 727 626 775 630
rect 779 626 799 630
rect 91 625 799 626
rect 805 625 806 631
rect 96 569 97 575
rect 103 574 811 575
rect 103 570 111 574
rect 115 570 171 574
rect 175 570 227 574
rect 231 570 299 574
rect 303 570 323 574
rect 327 570 387 574
rect 391 570 427 574
rect 431 570 475 574
rect 479 570 539 574
rect 543 570 571 574
rect 575 570 651 574
rect 655 570 667 574
rect 671 570 747 574
rect 751 570 775 574
rect 779 570 811 574
rect 103 569 811 570
rect 817 569 818 575
rect 84 521 85 527
rect 91 526 799 527
rect 91 522 111 526
rect 115 522 147 526
rect 151 522 195 526
rect 199 522 203 526
rect 207 522 283 526
rect 287 522 299 526
rect 303 522 379 526
rect 383 522 403 526
rect 407 522 491 526
rect 495 522 515 526
rect 519 522 611 526
rect 615 522 627 526
rect 631 522 723 526
rect 727 522 775 526
rect 779 522 799 526
rect 91 521 799 522
rect 805 521 806 527
rect 96 469 97 475
rect 103 474 811 475
rect 103 470 111 474
rect 115 470 219 474
rect 223 470 307 474
rect 311 470 339 474
rect 343 470 395 474
rect 399 470 403 474
rect 407 470 451 474
rect 455 470 515 474
rect 519 470 587 474
rect 591 470 635 474
rect 639 470 667 474
rect 671 470 747 474
rect 751 470 775 474
rect 779 470 811 474
rect 103 469 811 470
rect 817 469 818 475
rect 84 413 85 419
rect 91 418 799 419
rect 91 414 111 418
rect 115 414 315 418
rect 319 414 371 418
rect 375 414 387 418
rect 391 414 427 418
rect 431 414 443 418
rect 447 414 491 418
rect 495 414 499 418
rect 503 414 555 418
rect 559 414 563 418
rect 567 414 611 418
rect 615 414 643 418
rect 647 414 667 418
rect 671 414 723 418
rect 727 414 775 418
rect 779 414 799 418
rect 91 413 799 414
rect 805 413 806 419
rect 96 361 97 367
rect 103 366 811 367
rect 103 362 111 366
rect 115 362 323 366
rect 327 362 379 366
rect 383 362 411 366
rect 415 362 435 366
rect 439 362 467 366
rect 471 362 499 366
rect 503 362 523 366
rect 527 362 571 366
rect 575 362 579 366
rect 583 362 635 366
rect 639 362 651 366
rect 655 362 691 366
rect 695 362 739 366
rect 743 362 747 366
rect 751 362 775 366
rect 779 362 811 366
rect 103 361 811 362
rect 817 361 818 367
rect 84 305 85 311
rect 91 310 799 311
rect 91 306 111 310
rect 115 306 171 310
rect 175 306 251 310
rect 255 306 299 310
rect 303 306 331 310
rect 335 306 355 310
rect 359 306 411 310
rect 415 306 419 310
rect 423 306 475 310
rect 479 306 515 310
rect 519 306 547 310
rect 551 306 611 310
rect 615 306 627 310
rect 631 306 715 310
rect 719 306 775 310
rect 779 306 799 310
rect 91 305 799 306
rect 805 305 806 311
rect 96 253 97 259
rect 103 258 811 259
rect 103 254 111 258
rect 115 254 171 258
rect 175 254 195 258
rect 199 254 267 258
rect 271 254 275 258
rect 279 254 355 258
rect 359 254 387 258
rect 391 254 443 258
rect 447 254 515 258
rect 519 254 539 258
rect 543 254 635 258
rect 639 254 643 258
rect 647 254 739 258
rect 743 254 747 258
rect 751 254 775 258
rect 779 254 811 258
rect 103 253 811 254
rect 817 253 818 259
rect 84 201 85 207
rect 91 206 799 207
rect 91 202 111 206
rect 115 202 147 206
rect 151 202 211 206
rect 215 202 243 206
rect 247 202 299 206
rect 303 202 363 206
rect 367 202 403 206
rect 407 202 491 206
rect 495 202 507 206
rect 511 202 619 206
rect 623 202 723 206
rect 727 202 775 206
rect 779 202 799 206
rect 91 201 799 202
rect 805 201 806 207
rect 96 141 97 147
rect 103 146 811 147
rect 103 142 111 146
rect 115 142 171 146
rect 175 142 187 146
rect 191 142 235 146
rect 239 142 243 146
rect 247 142 299 146
rect 303 142 323 146
rect 327 142 355 146
rect 359 142 411 146
rect 415 142 427 146
rect 431 142 467 146
rect 471 142 523 146
rect 527 142 531 146
rect 535 142 579 146
rect 583 142 635 146
rect 639 142 643 146
rect 647 142 691 146
rect 695 142 747 146
rect 751 142 775 146
rect 779 142 811 146
rect 103 141 811 142
rect 817 141 818 147
rect 84 93 85 99
rect 91 98 799 99
rect 91 94 111 98
rect 115 94 163 98
rect 167 94 219 98
rect 223 94 275 98
rect 279 94 331 98
rect 335 94 387 98
rect 391 94 443 98
rect 447 94 499 98
rect 503 94 555 98
rect 559 94 611 98
rect 615 94 667 98
rect 671 94 723 98
rect 727 94 775 98
rect 779 94 799 98
rect 91 93 799 94
rect 805 93 806 99
<< m5c >>
rect 85 841 91 847
rect 799 841 805 847
rect 97 781 103 787
rect 811 781 817 787
rect 85 733 91 739
rect 799 733 805 739
rect 97 685 103 691
rect 811 685 817 691
rect 85 625 91 631
rect 799 625 805 631
rect 97 569 103 575
rect 811 569 817 575
rect 85 521 91 527
rect 799 521 805 527
rect 97 469 103 475
rect 811 469 817 475
rect 85 413 91 419
rect 799 413 805 419
rect 97 361 103 367
rect 811 361 817 367
rect 85 305 91 311
rect 799 305 805 311
rect 97 253 103 259
rect 811 253 817 259
rect 85 201 91 207
rect 799 201 805 207
rect 97 141 103 147
rect 811 141 817 147
rect 85 93 91 99
rect 799 93 805 99
<< m5 >>
rect 84 847 92 864
rect 84 841 85 847
rect 91 841 92 847
rect 84 739 92 841
rect 84 733 85 739
rect 91 733 92 739
rect 84 631 92 733
rect 84 625 85 631
rect 91 625 92 631
rect 84 527 92 625
rect 84 521 85 527
rect 91 521 92 527
rect 84 419 92 521
rect 84 413 85 419
rect 91 413 92 419
rect 84 311 92 413
rect 84 305 85 311
rect 91 305 92 311
rect 84 207 92 305
rect 84 201 85 207
rect 91 201 92 207
rect 84 99 92 201
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 787 104 864
rect 96 781 97 787
rect 103 781 104 787
rect 96 691 104 781
rect 96 685 97 691
rect 103 685 104 691
rect 96 575 104 685
rect 96 569 97 575
rect 103 569 104 575
rect 96 475 104 569
rect 96 469 97 475
rect 103 469 104 475
rect 96 367 104 469
rect 96 361 97 367
rect 103 361 104 367
rect 96 259 104 361
rect 96 253 97 259
rect 103 253 104 259
rect 96 147 104 253
rect 96 141 97 147
rect 103 141 104 147
rect 96 72 104 141
rect 798 847 806 864
rect 798 841 799 847
rect 805 841 806 847
rect 798 739 806 841
rect 798 733 799 739
rect 805 733 806 739
rect 798 631 806 733
rect 798 625 799 631
rect 805 625 806 631
rect 798 527 806 625
rect 798 521 799 527
rect 805 521 806 527
rect 798 419 806 521
rect 798 413 799 419
rect 805 413 806 419
rect 798 311 806 413
rect 798 305 799 311
rect 805 305 806 311
rect 798 207 806 305
rect 798 201 799 207
rect 805 201 806 207
rect 798 99 806 201
rect 798 93 799 99
rect 805 93 806 99
rect 798 72 806 93
rect 810 787 818 864
rect 810 781 811 787
rect 817 781 818 787
rect 810 691 818 781
rect 810 685 811 691
rect 817 685 818 691
rect 810 575 818 685
rect 810 569 811 575
rect 817 569 818 575
rect 810 475 818 569
rect 810 469 811 475
rect 817 469 818 475
rect 810 367 818 469
rect 810 361 811 367
rect 817 361 818 367
rect 810 259 818 361
rect 810 253 811 259
rect 817 253 818 259
rect 810 147 818 253
rect 810 141 811 147
rect 817 141 818 147
rect 810 72 818 141
use welltap_svt  __well_tap__0
timestamp 1730591762
transform 1 0 104 0 1 104
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730591762
transform 1 0 104 0 1 104
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0NOR2X1  nor_563_6
timestamp 1730591762
transform 1 0 144 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_563_6
timestamp 1730591762
transform 1 0 144 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_564_6
timestamp 1730591762
transform 1 0 200 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_564_6
timestamp 1730591762
transform 1 0 200 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_565_6
timestamp 1730591762
transform 1 0 256 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_565_6
timestamp 1730591762
transform 1 0 256 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_566_6
timestamp 1730591762
transform 1 0 312 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_566_6
timestamp 1730591762
transform 1 0 312 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_567_6
timestamp 1730591762
transform 1 0 368 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_567_6
timestamp 1730591762
transform 1 0 368 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_568_6
timestamp 1730591762
transform 1 0 424 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_568_6
timestamp 1730591762
transform 1 0 424 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_569_6
timestamp 1730591762
transform 1 0 480 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_569_6
timestamp 1730591762
transform 1 0 480 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_570_6
timestamp 1730591762
transform 1 0 536 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_570_6
timestamp 1730591762
transform 1 0 536 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_599_6
timestamp 1730591762
transform 1 0 592 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_599_6
timestamp 1730591762
transform 1 0 592 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_598_6
timestamp 1730591762
transform 1 0 648 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_598_6
timestamp 1730591762
transform 1 0 648 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_597_6
timestamp 1730591762
transform 1 0 704 0 1 96
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_597_6
timestamp 1730591762
transform 1 0 704 0 1 96
box 9 2 47 46
use welltap_svt  __well_tap__1
timestamp 1730591762
transform 1 0 768 0 1 104
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730591762
transform 1 0 768 0 1 104
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_559_6
timestamp 1730591762
transform 1 0 128 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_559_6
timestamp 1730591762
transform 1 0 128 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_560_6
timestamp 1730591762
transform 1 0 192 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_560_6
timestamp 1730591762
transform 1 0 192 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_561_6
timestamp 1730591762
transform 1 0 280 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_561_6
timestamp 1730591762
transform 1 0 280 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_562_6
timestamp 1730591762
transform 1 0 384 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_562_6
timestamp 1730591762
transform 1 0 384 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_572_6
timestamp 1730591762
transform 1 0 488 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_572_6
timestamp 1730591762
transform 1 0 488 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_571_6
timestamp 1730591762
transform 1 0 600 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_571_6
timestamp 1730591762
transform 1 0 600 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_596_6
timestamp 1730591762
transform 1 0 704 0 -1 204
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_596_6
timestamp 1730591762
transform 1 0 704 0 -1 204
box 9 2 47 46
use welltap_svt  __well_tap__2
timestamp 1730591762
transform 1 0 104 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730591762
transform 1 0 104 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730591762
transform 1 0 768 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730591762
transform 1 0 768 0 -1 196
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730591762
transform 1 0 104 0 1 216
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730591762
transform 1 0 104 0 1 216
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_558_6
timestamp 1730591762
transform 1 0 128 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_558_6
timestamp 1730591762
transform 1 0 128 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_557_6
timestamp 1730591762
transform 1 0 224 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_557_6
timestamp 1730591762
transform 1 0 224 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_556_6
timestamp 1730591762
transform 1 0 344 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_556_6
timestamp 1730591762
transform 1 0 344 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_573_6
timestamp 1730591762
transform 1 0 472 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_573_6
timestamp 1730591762
transform 1 0 472 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_594_6
timestamp 1730591762
transform 1 0 600 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_594_6
timestamp 1730591762
transform 1 0 600 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_595_6
timestamp 1730591762
transform 1 0 704 0 1 208
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_595_6
timestamp 1730591762
transform 1 0 704 0 1 208
box 9 2 47 46
use welltap_svt  __well_tap__5
timestamp 1730591762
transform 1 0 768 0 1 216
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730591762
transform 1 0 768 0 1 216
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730591762
transform 1 0 104 0 -1 300
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730591762
transform 1 0 104 0 -1 300
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_553_6
timestamp 1730591762
transform 1 0 152 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_553_6
timestamp 1730591762
transform 1 0 152 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_554_6
timestamp 1730591762
transform 1 0 232 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_554_6
timestamp 1730591762
transform 1 0 232 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_555_6
timestamp 1730591762
transform 1 0 312 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_555_6
timestamp 1730591762
transform 1 0 312 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_552_6
timestamp 1730591762
transform 1 0 400 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_552_6
timestamp 1730591762
transform 1 0 400 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_574_6
timestamp 1730591762
transform 1 0 496 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_574_6
timestamp 1730591762
transform 1 0 496 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_575_6
timestamp 1730591762
transform 1 0 592 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_575_6
timestamp 1730591762
transform 1 0 592 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_593_6
timestamp 1730591762
transform 1 0 696 0 -1 308
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_593_6
timestamp 1730591762
transform 1 0 696 0 -1 308
box 9 2 47 46
use welltap_svt  __well_tap__7
timestamp 1730591762
transform 1 0 768 0 -1 300
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730591762
transform 1 0 768 0 -1 300
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730591762
transform 1 0 104 0 1 324
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730591762
transform 1 0 104 0 1 324
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_549_6
timestamp 1730591762
transform 1 0 280 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_549_6
timestamp 1730591762
transform 1 0 280 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_550_6
timestamp 1730591762
transform 1 0 336 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_550_6
timestamp 1730591762
transform 1 0 336 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_551_6
timestamp 1730591762
transform 1 0 392 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_551_6
timestamp 1730591762
transform 1 0 392 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_547_6
timestamp 1730591762
transform 1 0 456 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_547_6
timestamp 1730591762
transform 1 0 456 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_548_6
timestamp 1730591762
transform 1 0 528 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_548_6
timestamp 1730591762
transform 1 0 528 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_576_6
timestamp 1730591762
transform 1 0 608 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_576_6
timestamp 1730591762
transform 1 0 608 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_592_6
timestamp 1730591762
transform 1 0 696 0 1 316
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_592_6
timestamp 1730591762
transform 1 0 696 0 1 316
box 9 2 47 46
use welltap_svt  __well_tap__9
timestamp 1730591762
transform 1 0 768 0 1 324
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730591762
transform 1 0 768 0 1 324
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730591762
transform 1 0 104 0 -1 408
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730591762
transform 1 0 104 0 -1 408
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_545_6
timestamp 1730591762
transform 1 0 368 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_545_6
timestamp 1730591762
transform 1 0 368 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_546_6
timestamp 1730591762
transform 1 0 424 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_546_6
timestamp 1730591762
transform 1 0 424 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_544_6
timestamp 1730591762
transform 1 0 480 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_544_6
timestamp 1730591762
transform 1 0 480 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_543_6
timestamp 1730591762
transform 1 0 536 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_543_6
timestamp 1730591762
transform 1 0 536 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_542_6
timestamp 1730591762
transform 1 0 592 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_542_6
timestamp 1730591762
transform 1 0 592 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_577_6
timestamp 1730591762
transform 1 0 648 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_577_6
timestamp 1730591762
transform 1 0 648 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_591_6
timestamp 1730591762
transform 1 0 704 0 -1 416
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_591_6
timestamp 1730591762
transform 1 0 704 0 -1 416
box 9 2 47 46
use welltap_svt  __well_tap__11
timestamp 1730591762
transform 1 0 768 0 -1 408
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730591762
transform 1 0 768 0 -1 408
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_537_6
timestamp 1730591762
transform 1 0 296 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_537_6
timestamp 1730591762
transform 1 0 296 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_538_6
timestamp 1730591762
transform 1 0 352 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_538_6
timestamp 1730591762
transform 1 0 352 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_539_6
timestamp 1730591762
transform 1 0 408 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_539_6
timestamp 1730591762
transform 1 0 408 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_540_6
timestamp 1730591762
transform 1 0 472 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_540_6
timestamp 1730591762
transform 1 0 472 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_541_6
timestamp 1730591762
transform 1 0 544 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_541_6
timestamp 1730591762
transform 1 0 544 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_578_6
timestamp 1730591762
transform 1 0 624 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_578_6
timestamp 1730591762
transform 1 0 624 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_590_6
timestamp 1730591762
transform 1 0 704 0 1 424
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_590_6
timestamp 1730591762
transform 1 0 704 0 1 424
box 9 2 47 46
use welltap_svt  __well_tap__12
timestamp 1730591762
transform 1 0 104 0 1 432
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730591762
transform 1 0 104 0 1 432
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730591762
transform 1 0 768 0 1 432
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730591762
transform 1 0 768 0 1 432
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730591762
transform 1 0 104 0 -1 516
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730591762
transform 1 0 104 0 -1 516
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_532_6
timestamp 1730591762
transform 1 0 176 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_532_6
timestamp 1730591762
transform 1 0 176 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_533_6
timestamp 1730591762
transform 1 0 264 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_533_6
timestamp 1730591762
transform 1 0 264 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_534_6
timestamp 1730591762
transform 1 0 360 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_534_6
timestamp 1730591762
transform 1 0 360 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_535_6
timestamp 1730591762
transform 1 0 472 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_535_6
timestamp 1730591762
transform 1 0 472 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_536_6
timestamp 1730591762
transform 1 0 592 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_536_6
timestamp 1730591762
transform 1 0 592 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_589_6
timestamp 1730591762
transform 1 0 704 0 -1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_589_6
timestamp 1730591762
transform 1 0 704 0 -1 524
box 9 2 47 46
use welltap_svt  __well_tap__15
timestamp 1730591762
transform 1 0 768 0 -1 516
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730591762
transform 1 0 768 0 -1 516
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730591762
transform 1 0 104 0 1 532
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730591762
transform 1 0 104 0 1 532
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_527_6
timestamp 1730591762
transform 1 0 128 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_527_6
timestamp 1730591762
transform 1 0 128 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_528_6
timestamp 1730591762
transform 1 0 184 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_528_6
timestamp 1730591762
transform 1 0 184 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_529_6
timestamp 1730591762
transform 1 0 280 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_529_6
timestamp 1730591762
transform 1 0 280 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_530_6
timestamp 1730591762
transform 1 0 384 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_530_6
timestamp 1730591762
transform 1 0 384 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_531_6
timestamp 1730591762
transform 1 0 496 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_531_6
timestamp 1730591762
transform 1 0 496 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_579_6
timestamp 1730591762
transform 1 0 608 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_579_6
timestamp 1730591762
transform 1 0 608 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_588_6
timestamp 1730591762
transform 1 0 704 0 1 524
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_588_6
timestamp 1730591762
transform 1 0 704 0 1 524
box 9 2 47 46
use welltap_svt  __well_tap__17
timestamp 1730591762
transform 1 0 768 0 1 532
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730591762
transform 1 0 768 0 1 532
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730591762
transform 1 0 104 0 -1 620
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730591762
transform 1 0 104 0 -1 620
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_526_6
timestamp 1730591762
transform 1 0 128 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_526_6
timestamp 1730591762
transform 1 0 128 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_525_6
timestamp 1730591762
transform 1 0 184 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_525_6
timestamp 1730591762
transform 1 0 184 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_524_6
timestamp 1730591762
transform 1 0 256 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_524_6
timestamp 1730591762
transform 1 0 256 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_522_6
timestamp 1730591762
transform 1 0 344 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_522_6
timestamp 1730591762
transform 1 0 344 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_523_6
timestamp 1730591762
transform 1 0 432 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_523_6
timestamp 1730591762
transform 1 0 432 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_580_6
timestamp 1730591762
transform 1 0 528 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_580_6
timestamp 1730591762
transform 1 0 528 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_586_6
timestamp 1730591762
transform 1 0 624 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_586_6
timestamp 1730591762
transform 1 0 624 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_587_6
timestamp 1730591762
transform 1 0 704 0 -1 628
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_587_6
timestamp 1730591762
transform 1 0 704 0 -1 628
box 9 2 47 46
use welltap_svt  __well_tap__19
timestamp 1730591762
transform 1 0 768 0 -1 620
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730591762
transform 1 0 768 0 -1 620
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730591762
transform 1 0 104 0 1 648
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730591762
transform 1 0 104 0 1 648
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_519_6
timestamp 1730591762
transform 1 0 200 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_519_6
timestamp 1730591762
transform 1 0 200 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_520_6
timestamp 1730591762
transform 1 0 256 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_520_6
timestamp 1730591762
transform 1 0 256 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_521_6
timestamp 1730591762
transform 1 0 312 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_521_6
timestamp 1730591762
transform 1 0 312 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_518_6
timestamp 1730591762
transform 1 0 368 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_518_6
timestamp 1730591762
transform 1 0 368 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_517_6
timestamp 1730591762
transform 1 0 424 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_517_6
timestamp 1730591762
transform 1 0 424 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_581_6
timestamp 1730591762
transform 1 0 480 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_581_6
timestamp 1730591762
transform 1 0 480 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_582_6
timestamp 1730591762
transform 1 0 536 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_582_6
timestamp 1730591762
transform 1 0 536 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_583_6
timestamp 1730591762
transform 1 0 592 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_583_6
timestamp 1730591762
transform 1 0 592 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_584_6
timestamp 1730591762
transform 1 0 648 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_584_6
timestamp 1730591762
transform 1 0 648 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_585_6
timestamp 1730591762
transform 1 0 704 0 1 640
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_585_6
timestamp 1730591762
transform 1 0 704 0 1 640
box 9 2 47 46
use welltap_svt  __well_tap__21
timestamp 1730591762
transform 1 0 768 0 1 648
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730591762
transform 1 0 768 0 1 648
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_512_6
timestamp 1730591762
transform 1 0 320 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_512_6
timestamp 1730591762
transform 1 0 320 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_513_6
timestamp 1730591762
transform 1 0 376 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_513_6
timestamp 1730591762
transform 1 0 376 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_514_6
timestamp 1730591762
transform 1 0 432 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_514_6
timestamp 1730591762
transform 1 0 432 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_515_6
timestamp 1730591762
transform 1 0 488 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_515_6
timestamp 1730591762
transform 1 0 488 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_516_6
timestamp 1730591762
transform 1 0 544 0 -1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_516_6
timestamp 1730591762
transform 1 0 544 0 -1 736
box 9 2 47 46
use welltap_svt  __well_tap__22
timestamp 1730591762
transform 1 0 104 0 -1 728
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730591762
transform 1 0 104 0 -1 728
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_57_6
timestamp 1730591762
transform 1 0 184 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_57_6
timestamp 1730591762
transform 1 0 184 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_58_6
timestamp 1730591762
transform 1 0 240 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_58_6
timestamp 1730591762
transform 1 0 240 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_59_6
timestamp 1730591762
transform 1 0 296 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_59_6
timestamp 1730591762
transform 1 0 296 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_510_6
timestamp 1730591762
transform 1 0 352 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_510_6
timestamp 1730591762
transform 1 0 352 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_511_6
timestamp 1730591762
transform 1 0 408 0 1 736
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_511_6
timestamp 1730591762
transform 1 0 408 0 1 736
box 9 2 47 46
use welltap_svt  __well_tap__23
timestamp 1730591762
transform 1 0 768 0 -1 728
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730591762
transform 1 0 768 0 -1 728
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730591762
transform 1 0 104 0 1 744
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730591762
transform 1 0 104 0 1 744
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730591762
transform 1 0 768 0 1 744
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730591762
transform 1 0 768 0 1 744
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730591762
transform 1 0 104 0 -1 836
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730591762
transform 1 0 104 0 -1 836
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_50_6
timestamp 1730591762
transform 1 0 128 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_50_6
timestamp 1730591762
transform 1 0 128 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_51_6
timestamp 1730591762
transform 1 0 184 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_51_6
timestamp 1730591762
transform 1 0 184 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_52_6
timestamp 1730591762
transform 1 0 240 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_52_6
timestamp 1730591762
transform 1 0 240 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_53_6
timestamp 1730591762
transform 1 0 296 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_53_6
timestamp 1730591762
transform 1 0 296 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_54_6
timestamp 1730591762
transform 1 0 352 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_54_6
timestamp 1730591762
transform 1 0 352 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_55_6
timestamp 1730591762
transform 1 0 408 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_55_6
timestamp 1730591762
transform 1 0 408 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_56_6
timestamp 1730591762
transform 1 0 464 0 -1 844
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_56_6
timestamp 1730591762
transform 1 0 464 0 -1 844
box 9 2 47 46
use welltap_svt  __well_tap__27
timestamp 1730591762
transform 1 0 768 0 -1 836
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730591762
transform 1 0 768 0 -1 836
box 8 4 12 24
<< end >>
