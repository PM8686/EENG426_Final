magic
tech sky130l
timestamp 1730589202
<< m1 >>
rect 424 1463 428 1507
rect 832 1431 836 1467
rect 1232 1431 1236 1463
rect 512 1351 516 1391
rect 520 1367 524 1415
rect 640 1351 644 1371
rect 248 1319 252 1347
rect 272 1267 276 1283
rect 1120 1263 1132 1267
rect 1116 1259 1124 1263
rect 400 1215 404 1231
rect 1328 1227 1332 1255
rect 1432 1183 1436 1203
rect 176 1107 180 1123
rect 400 1083 404 1103
rect 1072 1099 1076 1123
rect 1432 1119 1436 1131
rect 1376 1087 1380 1111
rect 352 947 356 967
rect 1432 939 1436 959
rect 1376 891 1380 931
rect 656 867 660 887
rect 880 867 884 879
rect 656 863 668 867
rect 664 859 668 863
rect 248 787 252 819
rect 560 759 564 783
rect 1008 783 1012 799
rect 1400 787 1404 799
rect 736 743 740 771
rect 176 699 180 715
rect 728 703 732 715
rect 992 703 996 739
rect 1304 679 1308 703
rect 1368 703 1372 715
rect 344 643 352 647
rect 232 619 236 635
rect 344 623 348 643
rect 772 607 780 611
rect 776 599 780 607
rect 776 595 784 599
rect 1176 567 1180 607
rect 1024 383 1028 463
rect 728 379 744 383
rect 1432 371 1436 395
rect 216 295 220 311
rect 264 299 268 331
rect 1120 299 1124 339
rect 1400 299 1404 311
rect 1384 227 1388 271
rect 1072 155 1076 203
rect 1200 127 1204 151
<< m2c >>
rect 424 1507 428 1511
rect 111 1493 115 1497
rect 304 1495 308 1499
rect 328 1495 332 1499
rect 352 1495 356 1499
rect 376 1495 380 1499
rect 416 1495 420 1499
rect 328 1487 332 1491
rect 352 1487 356 1491
rect 376 1487 380 1491
rect 416 1487 420 1491
rect 111 1475 115 1479
rect 304 1471 308 1475
rect 656 1499 660 1503
rect 896 1499 900 1503
rect 464 1495 468 1499
rect 520 1495 524 1499
rect 584 1495 588 1499
rect 816 1495 820 1499
rect 968 1495 972 1499
rect 1040 1495 1044 1499
rect 1112 1495 1116 1499
rect 1184 1495 1188 1499
rect 1256 1495 1260 1499
rect 1447 1493 1451 1497
rect 464 1487 468 1491
rect 520 1487 524 1491
rect 584 1487 588 1491
rect 656 1487 660 1491
rect 736 1487 740 1491
rect 896 1487 900 1491
rect 1040 1487 1044 1491
rect 1112 1483 1116 1487
rect 816 1479 820 1483
rect 1184 1475 1188 1479
rect 1447 1475 1451 1479
rect 968 1471 972 1475
rect 1256 1471 1260 1475
rect 111 1457 115 1461
rect 416 1459 420 1463
rect 424 1459 428 1463
rect 832 1467 836 1471
rect 160 1451 164 1455
rect 768 1451 772 1455
rect 184 1443 188 1447
rect 208 1443 212 1447
rect 240 1443 244 1447
rect 280 1443 284 1447
rect 328 1443 332 1447
rect 376 1443 380 1447
rect 464 1443 468 1447
rect 512 1443 516 1447
rect 560 1443 564 1447
rect 616 1443 620 1447
rect 672 1443 676 1447
rect 720 1443 724 1447
rect 824 1443 828 1447
rect 111 1439 115 1443
rect 160 1435 164 1439
rect 184 1435 188 1439
rect 208 1435 212 1439
rect 240 1435 244 1439
rect 280 1435 284 1439
rect 328 1435 332 1439
rect 416 1435 420 1439
rect 464 1435 468 1439
rect 512 1435 516 1439
rect 560 1435 564 1439
rect 616 1435 620 1439
rect 672 1435 676 1439
rect 824 1435 828 1439
rect 376 1431 380 1435
rect 720 1431 724 1435
rect 768 1431 772 1435
rect 1232 1463 1236 1467
rect 1080 1459 1084 1463
rect 936 1451 940 1455
rect 1176 1451 1180 1455
rect 880 1443 884 1447
rect 984 1443 988 1447
rect 1032 1443 1036 1447
rect 1128 1443 1132 1447
rect 1224 1443 1228 1447
rect 936 1435 940 1439
rect 984 1435 988 1439
rect 1080 1435 1084 1439
rect 1224 1435 1228 1439
rect 880 1431 884 1435
rect 1032 1431 1036 1435
rect 1128 1431 1132 1435
rect 1176 1431 1180 1435
rect 1447 1457 1451 1461
rect 1272 1451 1276 1455
rect 1320 1443 1324 1447
rect 1447 1439 1451 1443
rect 1320 1435 1324 1439
rect 1272 1431 1276 1435
rect 832 1427 836 1431
rect 1232 1427 1236 1431
rect 424 1419 428 1423
rect 1032 1419 1036 1423
rect 1272 1419 1276 1423
rect 1400 1419 1404 1423
rect 111 1413 115 1417
rect 144 1415 148 1419
rect 168 1415 172 1419
rect 192 1415 196 1419
rect 232 1415 236 1419
rect 296 1415 300 1419
rect 360 1415 364 1419
rect 488 1415 492 1419
rect 520 1415 524 1419
rect 544 1415 548 1419
rect 592 1415 596 1419
rect 640 1415 644 1419
rect 696 1415 700 1419
rect 752 1415 756 1419
rect 808 1415 812 1419
rect 864 1415 868 1419
rect 920 1415 924 1419
rect 976 1415 980 1419
rect 1080 1415 1084 1419
rect 1128 1415 1132 1419
rect 1176 1415 1180 1419
rect 1224 1415 1228 1419
rect 1312 1415 1316 1419
rect 1352 1415 1356 1419
rect 1424 1415 1428 1419
rect 192 1407 196 1411
rect 232 1407 236 1411
rect 296 1407 300 1411
rect 360 1407 364 1411
rect 424 1407 428 1411
rect 168 1399 172 1403
rect 111 1395 115 1399
rect 144 1391 148 1395
rect 488 1391 492 1395
rect 512 1391 516 1395
rect 111 1377 115 1381
rect 144 1371 148 1375
rect 240 1371 244 1375
rect 344 1371 348 1375
rect 400 1371 404 1375
rect 496 1371 500 1375
rect 168 1363 172 1367
rect 192 1363 196 1367
rect 288 1363 292 1367
rect 448 1363 452 1367
rect 111 1359 115 1363
rect 144 1355 148 1359
rect 168 1355 172 1359
rect 192 1355 196 1359
rect 288 1355 292 1359
rect 344 1355 348 1359
rect 448 1355 452 1359
rect 496 1355 500 1359
rect 240 1351 244 1355
rect 400 1351 404 1355
rect 1447 1413 1451 1417
rect 544 1407 548 1411
rect 640 1407 644 1411
rect 696 1407 700 1411
rect 752 1407 756 1411
rect 808 1407 812 1411
rect 864 1407 868 1411
rect 976 1407 980 1411
rect 1032 1407 1036 1411
rect 1128 1407 1132 1411
rect 1224 1407 1228 1411
rect 1272 1407 1276 1411
rect 1312 1407 1316 1411
rect 1400 1407 1404 1411
rect 1080 1403 1084 1407
rect 592 1399 596 1403
rect 1352 1399 1356 1403
rect 1447 1395 1451 1399
rect 920 1391 924 1395
rect 1176 1391 1180 1395
rect 1424 1391 1428 1395
rect 888 1379 892 1383
rect 1056 1379 1060 1383
rect 1296 1379 1300 1383
rect 1447 1377 1451 1381
rect 576 1371 580 1375
rect 640 1371 644 1375
rect 672 1371 676 1375
rect 776 1371 780 1375
rect 944 1371 948 1375
rect 520 1363 524 1367
rect 536 1363 540 1367
rect 624 1363 628 1367
rect 536 1355 540 1359
rect 624 1355 628 1359
rect 576 1351 580 1355
rect 720 1363 724 1367
rect 832 1363 836 1367
rect 1000 1363 1004 1367
rect 1104 1363 1108 1367
rect 1152 1363 1156 1367
rect 1200 1363 1204 1367
rect 1248 1363 1252 1367
rect 1344 1363 1348 1367
rect 1392 1363 1396 1367
rect 1424 1363 1428 1367
rect 1447 1359 1451 1363
rect 720 1355 724 1359
rect 832 1355 836 1359
rect 888 1355 892 1359
rect 944 1355 948 1359
rect 1000 1355 1004 1359
rect 1056 1355 1060 1359
rect 1152 1355 1156 1359
rect 1200 1355 1204 1359
rect 1296 1355 1300 1359
rect 1392 1355 1396 1359
rect 672 1351 676 1355
rect 776 1351 780 1355
rect 1104 1351 1108 1355
rect 1248 1351 1252 1355
rect 1344 1351 1348 1355
rect 1424 1351 1428 1355
rect 248 1347 252 1351
rect 512 1347 516 1351
rect 640 1347 644 1351
rect 176 1339 180 1343
rect 111 1333 115 1337
rect 200 1335 204 1339
rect 240 1335 244 1339
rect 176 1327 180 1331
rect 200 1319 204 1323
rect 288 1339 292 1343
rect 344 1339 348 1343
rect 584 1339 588 1343
rect 1016 1339 1020 1343
rect 1168 1339 1172 1343
rect 1424 1339 1428 1343
rect 400 1335 404 1339
rect 464 1335 468 1339
rect 528 1335 532 1339
rect 640 1335 644 1339
rect 688 1335 692 1339
rect 736 1335 740 1339
rect 776 1335 780 1339
rect 808 1335 812 1339
rect 840 1335 844 1339
rect 872 1335 876 1339
rect 904 1335 908 1339
rect 936 1335 940 1339
rect 976 1335 980 1339
rect 1064 1335 1068 1339
rect 1112 1335 1116 1339
rect 1224 1335 1228 1339
rect 1280 1335 1284 1339
rect 1336 1335 1340 1339
rect 1392 1335 1396 1339
rect 1447 1333 1451 1337
rect 400 1327 404 1331
rect 584 1327 588 1331
rect 688 1327 692 1331
rect 736 1327 740 1331
rect 808 1327 812 1331
rect 872 1327 876 1331
rect 904 1327 908 1331
rect 936 1327 940 1331
rect 976 1327 980 1331
rect 1016 1327 1020 1331
rect 1112 1327 1116 1331
rect 1168 1327 1172 1331
rect 1280 1327 1284 1331
rect 288 1323 292 1327
rect 344 1323 348 1327
rect 464 1319 468 1323
rect 776 1319 780 1323
rect 840 1319 844 1323
rect 1336 1319 1340 1323
rect 111 1315 115 1319
rect 240 1315 244 1319
rect 248 1315 252 1319
rect 1447 1315 1451 1319
rect 528 1311 532 1315
rect 640 1311 644 1315
rect 1064 1311 1068 1315
rect 1224 1311 1228 1315
rect 1392 1311 1396 1315
rect 1424 1311 1428 1315
rect 111 1297 115 1301
rect 1120 1299 1124 1303
rect 1312 1299 1316 1303
rect 1447 1297 1451 1301
rect 240 1291 244 1295
rect 312 1291 316 1295
rect 384 1291 388 1295
rect 704 1291 708 1295
rect 800 1291 804 1295
rect 264 1283 268 1287
rect 272 1283 276 1287
rect 288 1283 292 1287
rect 336 1283 340 1287
rect 360 1283 364 1287
rect 408 1283 412 1287
rect 432 1283 436 1287
rect 456 1283 460 1287
rect 480 1283 484 1287
rect 512 1283 516 1287
rect 552 1283 556 1287
rect 600 1283 604 1287
rect 656 1283 660 1287
rect 752 1283 756 1287
rect 848 1283 852 1287
rect 888 1283 892 1287
rect 920 1283 924 1287
rect 960 1283 964 1287
rect 1000 1283 1004 1287
rect 1040 1283 1044 1287
rect 1080 1283 1084 1287
rect 1160 1283 1164 1287
rect 1208 1283 1212 1287
rect 1256 1283 1260 1287
rect 1376 1283 1380 1287
rect 1424 1283 1428 1287
rect 111 1279 115 1283
rect 240 1275 244 1279
rect 264 1275 268 1279
rect 1447 1279 1451 1283
rect 312 1275 316 1279
rect 336 1275 340 1279
rect 360 1275 364 1279
rect 384 1275 388 1279
rect 408 1275 412 1279
rect 432 1275 436 1279
rect 456 1275 460 1279
rect 480 1275 484 1279
rect 512 1275 516 1279
rect 552 1275 556 1279
rect 600 1275 604 1279
rect 704 1275 708 1279
rect 752 1275 756 1279
rect 800 1275 804 1279
rect 848 1275 852 1279
rect 888 1275 892 1279
rect 920 1275 924 1279
rect 960 1275 964 1279
rect 1000 1275 1004 1279
rect 1040 1275 1044 1279
rect 1080 1275 1084 1279
rect 1120 1275 1124 1279
rect 1160 1275 1164 1279
rect 1208 1275 1212 1279
rect 1256 1275 1260 1279
rect 1312 1275 1316 1279
rect 1424 1275 1428 1279
rect 288 1271 292 1275
rect 656 1271 660 1275
rect 1376 1271 1380 1275
rect 1128 1267 1132 1271
rect 272 1263 276 1267
rect 320 1259 324 1263
rect 368 1259 372 1263
rect 488 1259 492 1263
rect 920 1259 924 1263
rect 1072 1259 1076 1263
rect 1112 1259 1116 1263
rect 1136 1259 1140 1263
rect 1384 1259 1388 1263
rect 111 1253 115 1257
rect 344 1255 348 1259
rect 392 1255 396 1259
rect 424 1255 428 1259
rect 456 1255 460 1259
rect 528 1255 532 1259
rect 568 1255 572 1259
rect 624 1255 628 1259
rect 688 1255 692 1259
rect 760 1255 764 1259
rect 840 1255 844 1259
rect 1000 1255 1004 1259
rect 1200 1255 1204 1259
rect 1256 1255 1260 1259
rect 1320 1255 1324 1259
rect 1328 1255 1332 1259
rect 1424 1255 1428 1259
rect 320 1247 324 1251
rect 368 1247 372 1251
rect 456 1247 460 1251
rect 488 1247 492 1251
rect 568 1247 572 1251
rect 624 1247 628 1251
rect 688 1247 692 1251
rect 920 1247 924 1251
rect 1000 1247 1004 1251
rect 1072 1247 1076 1251
rect 1136 1247 1140 1251
rect 1320 1247 1324 1251
rect 344 1239 348 1243
rect 424 1239 428 1243
rect 528 1239 532 1243
rect 840 1239 844 1243
rect 1200 1239 1204 1243
rect 111 1235 115 1239
rect 392 1231 396 1235
rect 400 1231 404 1235
rect 760 1231 764 1235
rect 1256 1231 1260 1235
rect 111 1217 115 1221
rect 1447 1253 1451 1257
rect 1384 1247 1388 1251
rect 1447 1235 1451 1239
rect 1424 1231 1428 1235
rect 1328 1223 1332 1227
rect 1447 1217 1451 1221
rect 400 1211 404 1215
rect 496 1211 500 1215
rect 760 1211 764 1215
rect 856 1211 860 1215
rect 952 1211 956 1215
rect 1048 1211 1052 1215
rect 1184 1211 1188 1215
rect 1352 1211 1356 1215
rect 336 1203 340 1207
rect 376 1203 380 1207
rect 416 1203 420 1207
rect 456 1203 460 1207
rect 536 1203 540 1207
rect 576 1203 580 1207
rect 616 1203 620 1207
rect 664 1203 668 1207
rect 712 1203 716 1207
rect 808 1203 812 1207
rect 904 1203 908 1207
rect 1000 1203 1004 1207
rect 1112 1203 1116 1207
rect 1264 1203 1268 1207
rect 1424 1203 1428 1207
rect 1432 1203 1436 1207
rect 111 1199 115 1203
rect 336 1195 340 1199
rect 376 1195 380 1199
rect 416 1195 420 1199
rect 456 1195 460 1199
rect 496 1195 500 1199
rect 536 1195 540 1199
rect 576 1195 580 1199
rect 616 1195 620 1199
rect 664 1195 668 1199
rect 760 1195 764 1199
rect 808 1195 812 1199
rect 904 1195 908 1199
rect 1000 1195 1004 1199
rect 1048 1195 1052 1199
rect 1112 1195 1116 1199
rect 1264 1195 1268 1199
rect 1424 1195 1428 1199
rect 712 1191 716 1195
rect 856 1191 860 1195
rect 952 1191 956 1195
rect 1184 1191 1188 1195
rect 1352 1191 1356 1195
rect 1447 1199 1451 1203
rect 144 1179 148 1183
rect 344 1179 348 1183
rect 432 1179 436 1183
rect 472 1179 476 1183
rect 920 1179 924 1183
rect 1240 1179 1244 1183
rect 1424 1179 1428 1183
rect 1432 1179 1436 1183
rect 111 1173 115 1177
rect 168 1175 172 1179
rect 192 1175 196 1179
rect 216 1175 220 1179
rect 240 1175 244 1179
rect 264 1175 268 1179
rect 288 1175 292 1179
rect 312 1175 316 1179
rect 392 1175 396 1179
rect 512 1175 516 1179
rect 552 1175 556 1179
rect 592 1175 596 1179
rect 632 1175 636 1179
rect 680 1175 684 1179
rect 728 1175 732 1179
rect 776 1175 780 1179
rect 824 1175 828 1179
rect 872 1175 876 1179
rect 968 1175 972 1179
rect 1016 1175 1020 1179
rect 1064 1175 1068 1179
rect 1112 1175 1116 1179
rect 1160 1175 1164 1179
rect 1200 1175 1204 1179
rect 1280 1175 1284 1179
rect 1320 1175 1324 1179
rect 1360 1175 1364 1179
rect 1400 1175 1404 1179
rect 1447 1173 1451 1177
rect 216 1167 220 1171
rect 240 1167 244 1171
rect 288 1167 292 1171
rect 312 1167 316 1171
rect 344 1167 348 1171
rect 472 1167 476 1171
rect 872 1167 876 1171
rect 920 1167 924 1171
rect 968 1167 972 1171
rect 1360 1167 1364 1171
rect 1424 1167 1428 1171
rect 432 1163 436 1167
rect 192 1159 196 1163
rect 264 1159 268 1163
rect 512 1159 516 1163
rect 1016 1159 1020 1163
rect 1240 1159 1244 1163
rect 1320 1159 1324 1163
rect 111 1155 115 1159
rect 392 1155 396 1159
rect 552 1155 556 1159
rect 592 1155 596 1159
rect 632 1155 636 1159
rect 680 1155 684 1159
rect 728 1155 732 1159
rect 776 1155 780 1159
rect 1064 1155 1068 1159
rect 1112 1155 1116 1159
rect 1200 1155 1204 1159
rect 1447 1155 1451 1159
rect 144 1151 148 1155
rect 168 1151 172 1155
rect 824 1151 828 1155
rect 1160 1151 1164 1155
rect 1280 1151 1284 1155
rect 1400 1151 1404 1155
rect 111 1137 115 1141
rect 1447 1137 1451 1141
rect 144 1131 148 1135
rect 224 1131 228 1135
rect 384 1131 388 1135
rect 472 1131 476 1135
rect 592 1131 596 1135
rect 720 1131 724 1135
rect 840 1131 844 1135
rect 952 1131 956 1135
rect 1064 1131 1068 1135
rect 1280 1131 1284 1135
rect 1400 1131 1404 1135
rect 1432 1131 1436 1135
rect 168 1123 172 1127
rect 176 1123 180 1127
rect 192 1123 196 1127
rect 264 1123 268 1127
rect 304 1123 308 1127
rect 344 1123 348 1127
rect 424 1123 428 1127
rect 528 1123 532 1127
rect 656 1123 660 1127
rect 776 1123 780 1127
rect 896 1123 900 1127
rect 1008 1123 1012 1127
rect 1072 1123 1076 1127
rect 1112 1123 1116 1127
rect 1160 1123 1164 1127
rect 1200 1123 1204 1127
rect 1240 1123 1244 1127
rect 1320 1123 1324 1127
rect 1360 1123 1364 1127
rect 1424 1123 1428 1127
rect 111 1119 115 1123
rect 144 1115 148 1119
rect 168 1115 172 1119
rect 224 1115 228 1119
rect 264 1115 268 1119
rect 304 1115 308 1119
rect 344 1115 348 1119
rect 424 1115 428 1119
rect 528 1115 532 1119
rect 656 1115 660 1119
rect 776 1115 780 1119
rect 840 1115 844 1119
rect 896 1115 900 1119
rect 1008 1115 1012 1119
rect 192 1111 196 1115
rect 384 1111 388 1115
rect 472 1111 476 1115
rect 592 1111 596 1115
rect 720 1111 724 1115
rect 952 1111 956 1115
rect 1064 1111 1068 1115
rect 176 1103 180 1107
rect 400 1103 404 1107
rect 192 1095 196 1099
rect 336 1095 340 1099
rect 111 1089 115 1093
rect 144 1091 148 1095
rect 168 1091 172 1095
rect 216 1091 220 1095
rect 256 1091 260 1095
rect 296 1091 300 1095
rect 376 1091 380 1095
rect 192 1083 196 1087
rect 216 1083 220 1087
rect 376 1083 380 1087
rect 1447 1119 1451 1123
rect 1112 1115 1116 1119
rect 1160 1115 1164 1119
rect 1200 1115 1204 1119
rect 1280 1115 1284 1119
rect 1320 1115 1324 1119
rect 1400 1115 1404 1119
rect 1424 1115 1428 1119
rect 1432 1115 1436 1119
rect 1240 1111 1244 1115
rect 1360 1111 1364 1115
rect 1376 1111 1380 1115
rect 1064 1095 1068 1099
rect 1072 1095 1076 1099
rect 1176 1095 1180 1099
rect 416 1091 420 1095
rect 464 1091 468 1095
rect 512 1091 516 1095
rect 568 1091 572 1095
rect 616 1091 620 1095
rect 664 1091 668 1095
rect 712 1091 716 1095
rect 752 1091 756 1095
rect 800 1091 804 1095
rect 848 1091 852 1095
rect 896 1091 900 1095
rect 952 1091 956 1095
rect 1008 1091 1012 1095
rect 1120 1091 1124 1095
rect 1224 1091 1228 1095
rect 1280 1091 1284 1095
rect 1336 1091 1340 1095
rect 1392 1095 1396 1099
rect 1424 1095 1428 1099
rect 1447 1089 1451 1093
rect 464 1083 468 1087
rect 512 1083 516 1087
rect 568 1083 572 1087
rect 616 1083 620 1087
rect 712 1083 716 1087
rect 752 1083 756 1087
rect 800 1083 804 1087
rect 848 1083 852 1087
rect 896 1083 900 1087
rect 952 1083 956 1087
rect 1008 1083 1012 1087
rect 1064 1083 1068 1087
rect 1224 1083 1228 1087
rect 1376 1083 1380 1087
rect 1392 1083 1396 1087
rect 336 1079 340 1083
rect 400 1079 404 1083
rect 1176 1079 1180 1083
rect 168 1075 172 1079
rect 256 1075 260 1079
rect 416 1075 420 1079
rect 1120 1075 1124 1079
rect 1280 1075 1284 1079
rect 111 1071 115 1075
rect 144 1071 148 1075
rect 1336 1071 1340 1075
rect 1447 1071 1451 1075
rect 296 1067 300 1071
rect 664 1067 668 1071
rect 1424 1067 1428 1071
rect 111 1053 115 1057
rect 984 1055 988 1059
rect 1447 1053 1451 1057
rect 144 1047 148 1051
rect 280 1047 284 1051
rect 360 1047 364 1051
rect 640 1047 644 1051
rect 832 1047 836 1051
rect 1184 1047 1188 1051
rect 1280 1047 1284 1051
rect 168 1039 172 1043
rect 192 1039 196 1043
rect 216 1039 220 1043
rect 240 1039 244 1043
rect 320 1039 324 1043
rect 400 1039 404 1043
rect 440 1039 444 1043
rect 480 1039 484 1043
rect 520 1039 524 1043
rect 560 1039 564 1043
rect 600 1039 604 1043
rect 680 1039 684 1043
rect 720 1039 724 1043
rect 752 1039 756 1043
rect 792 1039 796 1043
rect 880 1039 884 1043
rect 928 1039 932 1043
rect 1040 1039 1044 1043
rect 1088 1039 1092 1043
rect 1136 1039 1140 1043
rect 1232 1039 1236 1043
rect 1336 1039 1340 1043
rect 1392 1039 1396 1043
rect 1424 1039 1428 1043
rect 111 1035 115 1039
rect 1447 1035 1451 1039
rect 144 1031 148 1035
rect 168 1031 172 1035
rect 192 1031 196 1035
rect 216 1031 220 1035
rect 240 1031 244 1035
rect 280 1031 284 1035
rect 320 1031 324 1035
rect 360 1031 364 1035
rect 400 1031 404 1035
rect 440 1031 444 1035
rect 480 1031 484 1035
rect 520 1031 524 1035
rect 560 1031 564 1035
rect 640 1031 644 1035
rect 680 1031 684 1035
rect 720 1031 724 1035
rect 752 1031 756 1035
rect 792 1031 796 1035
rect 880 1031 884 1035
rect 984 1031 988 1035
rect 1040 1031 1044 1035
rect 1088 1031 1092 1035
rect 1136 1031 1140 1035
rect 1232 1031 1236 1035
rect 1336 1031 1340 1035
rect 1392 1031 1396 1035
rect 1424 1031 1428 1035
rect 600 1027 604 1031
rect 832 1027 836 1031
rect 928 1027 932 1031
rect 1184 1027 1188 1031
rect 1280 1027 1284 1031
rect 168 1015 172 1019
rect 584 1015 588 1019
rect 776 1015 780 1019
rect 1000 1015 1004 1019
rect 1392 1015 1396 1019
rect 111 1009 115 1013
rect 192 1011 196 1015
rect 216 1011 220 1015
rect 240 1011 244 1015
rect 272 1011 276 1015
rect 312 1011 316 1015
rect 352 1011 356 1015
rect 392 1011 396 1015
rect 440 1011 444 1015
rect 488 1011 492 1015
rect 536 1011 540 1015
rect 632 1011 636 1015
rect 680 1011 684 1015
rect 728 1011 732 1015
rect 832 1011 836 1015
rect 888 1011 892 1015
rect 944 1011 948 1015
rect 1056 1011 1060 1015
rect 1112 1011 1116 1015
rect 1168 1011 1172 1015
rect 1224 1011 1228 1015
rect 1280 1011 1284 1015
rect 1336 1011 1340 1015
rect 1424 1011 1428 1015
rect 1447 1009 1451 1013
rect 168 1003 172 1007
rect 392 1003 396 1007
rect 584 1003 588 1007
rect 680 1003 684 1007
rect 728 1003 732 1007
rect 776 1003 780 1007
rect 832 1003 836 1007
rect 1000 1003 1004 1007
rect 1168 1003 1172 1007
rect 1224 1003 1228 1007
rect 1336 1003 1340 1007
rect 1392 1003 1396 1007
rect 192 995 196 999
rect 440 995 444 999
rect 944 995 948 999
rect 1056 995 1060 999
rect 1280 995 1284 999
rect 111 991 115 995
rect 216 991 220 995
rect 240 991 244 995
rect 272 991 276 995
rect 312 991 316 995
rect 352 991 356 995
rect 488 991 492 995
rect 536 991 540 995
rect 1447 991 1451 995
rect 632 987 636 991
rect 888 987 892 991
rect 1112 987 1116 991
rect 1424 987 1428 991
rect 111 973 115 977
rect 896 975 900 979
rect 1447 973 1451 977
rect 216 967 220 971
rect 296 967 300 971
rect 352 967 356 971
rect 384 967 388 971
rect 432 967 436 971
rect 576 967 580 971
rect 784 967 788 971
rect 1152 967 1156 971
rect 240 959 244 963
rect 264 959 268 963
rect 336 959 340 963
rect 111 955 115 959
rect 216 951 220 955
rect 240 951 244 955
rect 264 951 268 955
rect 296 951 300 955
rect 336 951 340 955
rect 480 959 484 963
rect 528 959 532 963
rect 632 959 636 963
rect 688 959 692 963
rect 736 959 740 963
rect 840 959 844 963
rect 952 959 956 963
rect 1008 959 1012 963
rect 1056 959 1060 963
rect 1104 959 1108 963
rect 1200 959 1204 963
rect 1248 959 1252 963
rect 1296 959 1300 963
rect 1344 959 1348 963
rect 1392 959 1396 963
rect 1424 959 1428 963
rect 1432 959 1436 963
rect 432 951 436 955
rect 480 951 484 955
rect 576 951 580 955
rect 632 951 636 955
rect 688 951 692 955
rect 840 951 844 955
rect 896 951 900 955
rect 952 951 956 955
rect 1008 951 1012 955
rect 1056 951 1060 955
rect 1104 951 1108 955
rect 1152 951 1156 955
rect 1200 951 1204 955
rect 1248 951 1252 955
rect 1296 951 1300 955
rect 1344 951 1348 955
rect 1424 951 1428 955
rect 384 947 388 951
rect 528 947 532 951
rect 736 947 740 951
rect 784 947 788 951
rect 1392 947 1396 951
rect 352 943 356 947
rect 1447 955 1451 959
rect 296 935 300 939
rect 736 935 740 939
rect 928 935 932 939
rect 1424 935 1428 939
rect 1432 935 1436 939
rect 111 929 115 933
rect 224 931 228 935
rect 248 931 252 935
rect 272 931 276 935
rect 328 931 332 935
rect 360 931 364 935
rect 400 931 404 935
rect 440 931 444 935
rect 480 931 484 935
rect 528 931 532 935
rect 576 931 580 935
rect 624 931 628 935
rect 680 931 684 935
rect 792 931 796 935
rect 856 931 860 935
rect 1000 931 1004 935
rect 1064 931 1068 935
rect 1128 931 1132 935
rect 1184 931 1188 935
rect 1232 931 1236 935
rect 1272 931 1276 935
rect 1304 931 1308 935
rect 1336 931 1340 935
rect 1368 931 1372 935
rect 1376 931 1380 935
rect 1400 931 1404 935
rect 224 923 228 927
rect 440 923 444 927
rect 480 923 484 927
rect 528 923 532 927
rect 624 923 628 927
rect 680 923 684 927
rect 736 923 740 927
rect 792 923 796 927
rect 856 923 860 927
rect 1000 923 1004 927
rect 1128 923 1132 927
rect 1184 923 1188 927
rect 1232 923 1236 927
rect 1272 923 1276 927
rect 1304 923 1308 927
rect 1368 923 1372 927
rect 296 919 300 923
rect 928 919 932 923
rect 248 915 252 919
rect 1336 915 1340 919
rect 111 911 115 915
rect 272 911 276 915
rect 328 911 332 915
rect 360 911 364 915
rect 400 907 404 911
rect 576 907 580 911
rect 1064 907 1068 911
rect 111 893 115 897
rect 504 895 508 899
rect 816 895 820 899
rect 1447 929 1451 933
rect 1424 923 1428 927
rect 1447 911 1451 915
rect 1400 907 1404 911
rect 1447 893 1451 897
rect 432 887 436 891
rect 544 887 548 891
rect 656 887 660 891
rect 712 887 716 891
rect 1128 887 1132 891
rect 1240 887 1244 891
rect 1376 887 1380 891
rect 1392 887 1396 891
rect 240 883 244 887
rect 264 879 268 883
rect 288 879 292 883
rect 312 879 316 883
rect 336 879 340 883
rect 368 879 372 883
rect 400 879 404 883
rect 464 879 468 883
rect 584 879 588 883
rect 632 879 636 883
rect 111 875 115 879
rect 240 871 244 875
rect 264 871 268 875
rect 288 871 292 875
rect 312 871 316 875
rect 336 871 340 875
rect 368 871 372 875
rect 400 871 404 875
rect 464 871 468 875
rect 504 871 508 875
rect 544 871 548 875
rect 584 871 588 875
rect 632 871 636 875
rect 432 867 436 871
rect 672 879 676 883
rect 760 879 764 883
rect 872 879 876 883
rect 880 879 884 883
rect 936 879 940 883
rect 1000 879 1004 883
rect 1064 879 1068 883
rect 1184 879 1188 883
rect 1288 879 1292 883
rect 1336 879 1340 883
rect 1424 879 1428 883
rect 760 871 764 875
rect 816 871 820 875
rect 872 871 876 875
rect 672 867 676 871
rect 712 867 716 871
rect 1447 875 1451 879
rect 936 871 940 875
rect 1000 871 1004 875
rect 1064 871 1068 875
rect 1128 871 1132 875
rect 1184 871 1188 875
rect 1240 871 1244 875
rect 1288 871 1292 875
rect 1392 871 1396 875
rect 1336 867 1340 871
rect 1424 867 1428 871
rect 880 863 884 867
rect 360 855 364 859
rect 656 855 660 859
rect 664 855 668 859
rect 992 855 996 859
rect 1056 855 1060 859
rect 1216 855 1220 859
rect 1424 855 1428 859
rect 111 849 115 853
rect 216 851 220 855
rect 240 851 244 855
rect 264 851 268 855
rect 296 851 300 855
rect 328 851 332 855
rect 392 851 396 855
rect 424 851 428 855
rect 456 851 460 855
rect 488 851 492 855
rect 520 851 524 855
rect 560 851 564 855
rect 608 851 612 855
rect 712 851 716 855
rect 776 851 780 855
rect 848 851 852 855
rect 920 851 924 855
rect 1112 851 1116 855
rect 1168 851 1172 855
rect 1256 851 1260 855
rect 1304 851 1308 855
rect 1352 851 1356 855
rect 1400 851 1404 855
rect 1447 849 1451 853
rect 264 843 268 847
rect 296 843 300 847
rect 328 843 332 847
rect 360 843 364 847
rect 392 843 396 847
rect 424 843 428 847
rect 456 843 460 847
rect 488 843 492 847
rect 560 843 564 847
rect 608 843 612 847
rect 656 843 660 847
rect 920 843 924 847
rect 992 843 996 847
rect 1056 843 1060 847
rect 1216 843 1220 847
rect 1424 843 1428 847
rect 240 835 244 839
rect 712 835 716 839
rect 1112 835 1116 839
rect 1256 835 1260 839
rect 111 831 115 835
rect 776 831 780 835
rect 1168 831 1172 835
rect 1304 831 1308 835
rect 1447 831 1451 835
rect 216 827 220 831
rect 520 827 524 831
rect 848 827 852 831
rect 1352 827 1356 831
rect 1400 827 1404 831
rect 248 819 252 823
rect 111 813 115 817
rect 144 807 148 811
rect 168 799 172 803
rect 192 799 196 803
rect 224 799 228 803
rect 111 795 115 799
rect 144 791 148 795
rect 168 791 172 795
rect 192 791 196 795
rect 224 791 228 795
rect 664 815 668 819
rect 1447 813 1451 817
rect 440 807 444 811
rect 720 807 724 811
rect 824 807 828 811
rect 912 807 916 811
rect 976 807 980 811
rect 1024 807 1028 811
rect 1136 807 1140 811
rect 1216 807 1220 811
rect 1320 807 1324 811
rect 1104 803 1108 807
rect 272 799 276 803
rect 320 799 324 803
rect 376 799 380 803
rect 496 799 500 803
rect 552 799 556 803
rect 608 799 612 803
rect 776 799 780 803
rect 872 799 876 803
rect 944 799 948 803
rect 1000 799 1004 803
rect 1008 799 1012 803
rect 1048 799 1052 803
rect 1072 799 1076 803
rect 1176 799 1180 803
rect 1264 799 1268 803
rect 1384 799 1388 803
rect 1400 799 1404 803
rect 1424 799 1428 803
rect 272 791 276 795
rect 320 791 324 795
rect 440 791 444 795
rect 496 791 500 795
rect 608 791 612 795
rect 664 791 668 795
rect 776 791 780 795
rect 824 791 828 795
rect 912 791 916 795
rect 944 791 948 795
rect 976 791 980 795
rect 1000 791 1004 795
rect 376 787 380 791
rect 552 787 556 791
rect 720 787 724 791
rect 872 787 876 791
rect 248 783 252 787
rect 560 783 564 787
rect 416 775 420 779
rect 111 769 115 773
rect 144 771 148 775
rect 168 771 172 775
rect 192 771 196 775
rect 232 771 236 775
rect 288 771 292 775
rect 352 771 356 775
rect 472 771 476 775
rect 528 771 532 775
rect 192 763 196 767
rect 232 763 236 767
rect 288 763 292 767
rect 416 763 420 767
rect 472 763 476 767
rect 1048 791 1052 795
rect 1072 791 1076 795
rect 1176 791 1180 795
rect 1264 791 1268 795
rect 1384 791 1388 795
rect 1024 787 1028 791
rect 1104 787 1108 791
rect 1136 787 1140 791
rect 1216 787 1220 791
rect 1320 787 1324 791
rect 1447 795 1451 799
rect 1424 787 1428 791
rect 1400 783 1404 787
rect 1008 779 1012 783
rect 584 775 588 779
rect 808 775 812 779
rect 968 775 972 779
rect 1424 775 1428 779
rect 632 771 636 775
rect 680 771 684 775
rect 728 771 732 775
rect 736 771 740 775
rect 768 771 772 775
rect 848 771 852 775
rect 888 771 892 775
rect 928 771 932 775
rect 1000 771 1004 775
rect 1032 771 1036 775
rect 1064 771 1068 775
rect 1096 771 1100 775
rect 1136 771 1140 775
rect 1184 771 1188 775
rect 1240 771 1244 775
rect 1304 771 1308 775
rect 1376 771 1380 775
rect 728 763 732 767
rect 584 759 588 763
rect 632 759 636 763
rect 168 755 172 759
rect 352 755 356 759
rect 528 755 532 759
rect 560 755 564 759
rect 111 751 115 755
rect 144 747 148 751
rect 680 747 684 751
rect 1447 769 1451 773
rect 808 763 812 767
rect 848 763 852 767
rect 968 763 972 767
rect 1000 763 1004 767
rect 1424 763 1428 767
rect 888 755 892 759
rect 1032 755 1036 759
rect 928 751 932 755
rect 1064 751 1068 755
rect 1096 751 1100 755
rect 1136 751 1140 755
rect 1184 751 1188 755
rect 1240 751 1244 755
rect 1447 751 1451 755
rect 768 747 772 751
rect 1304 747 1308 751
rect 1376 747 1380 751
rect 736 739 740 743
rect 992 739 996 743
rect 111 729 115 733
rect 384 731 388 735
rect 672 731 676 735
rect 144 723 148 727
rect 192 723 196 727
rect 272 723 276 727
rect 432 723 436 727
rect 528 723 532 727
rect 624 723 628 727
rect 816 723 820 727
rect 952 723 956 727
rect 168 715 172 719
rect 176 715 180 719
rect 224 715 228 719
rect 328 715 332 719
rect 480 715 484 719
rect 576 715 580 719
rect 712 715 716 719
rect 728 715 732 719
rect 760 715 764 719
rect 880 715 884 719
rect 111 711 115 715
rect 144 707 148 711
rect 168 707 172 711
rect 224 707 228 711
rect 272 707 276 711
rect 328 707 332 711
rect 480 707 484 711
rect 576 707 580 711
rect 672 707 676 711
rect 712 707 716 711
rect 192 703 196 707
rect 384 703 388 707
rect 432 703 436 707
rect 528 703 532 707
rect 624 703 628 707
rect 760 707 764 711
rect 880 707 884 711
rect 816 703 820 707
rect 952 703 956 707
rect 1447 729 1451 733
rect 1096 723 1100 727
rect 1160 723 1164 727
rect 1024 715 1028 719
rect 1224 715 1228 719
rect 1280 715 1284 719
rect 1336 715 1340 719
rect 1368 715 1372 719
rect 1392 715 1396 719
rect 1424 715 1428 719
rect 1024 707 1028 711
rect 1160 707 1164 711
rect 1224 707 1228 711
rect 1336 707 1340 711
rect 1096 703 1100 707
rect 1280 703 1284 707
rect 1304 703 1308 707
rect 728 699 732 703
rect 992 699 996 703
rect 176 695 180 699
rect 144 691 148 695
rect 768 691 772 695
rect 976 691 980 695
rect 1288 691 1292 695
rect 111 685 115 689
rect 168 687 172 691
rect 208 687 212 691
rect 248 687 252 691
rect 296 687 300 691
rect 344 687 348 691
rect 400 687 404 691
rect 448 687 452 691
rect 496 687 500 691
rect 544 687 548 691
rect 592 687 596 691
rect 648 687 652 691
rect 704 687 708 691
rect 840 687 844 691
rect 912 687 916 691
rect 1040 687 1044 691
rect 1096 687 1100 691
rect 1144 687 1148 691
rect 1184 687 1188 691
rect 1224 687 1228 691
rect 1256 687 1260 691
rect 144 679 148 683
rect 400 679 404 683
rect 448 679 452 683
rect 704 679 708 683
rect 768 679 772 683
rect 840 679 844 683
rect 912 679 916 683
rect 976 679 980 683
rect 1096 679 1100 683
rect 1144 679 1148 683
rect 1184 679 1188 683
rect 1224 679 1228 683
rect 1288 679 1292 683
rect 1447 711 1451 715
rect 1392 703 1396 707
rect 1424 703 1428 707
rect 1368 699 1372 703
rect 1424 691 1428 695
rect 1320 687 1324 691
rect 1352 687 1356 691
rect 1376 687 1380 691
rect 1400 687 1404 691
rect 1447 685 1451 689
rect 1352 679 1356 683
rect 1424 679 1428 683
rect 1304 675 1308 679
rect 168 671 172 675
rect 1256 671 1260 675
rect 1320 671 1324 675
rect 1400 671 1404 675
rect 111 667 115 671
rect 208 667 212 671
rect 248 667 252 671
rect 296 667 300 671
rect 496 667 500 671
rect 544 667 548 671
rect 1447 667 1451 671
rect 344 663 348 667
rect 592 663 596 667
rect 648 663 652 667
rect 1040 663 1044 667
rect 1376 663 1380 667
rect 111 649 115 653
rect 824 651 828 655
rect 1447 649 1451 653
rect 200 643 204 647
rect 248 643 252 647
rect 304 643 308 647
rect 352 643 356 647
rect 376 643 380 647
rect 416 643 420 647
rect 512 643 516 647
rect 616 643 620 647
rect 872 643 876 647
rect 1200 643 1204 647
rect 1272 643 1276 647
rect 1352 643 1356 647
rect 224 635 228 639
rect 232 635 236 639
rect 272 635 276 639
rect 336 635 340 639
rect 111 631 115 635
rect 200 627 204 631
rect 224 627 228 631
rect 272 627 276 631
rect 304 627 308 631
rect 336 627 340 631
rect 248 623 252 627
rect 464 635 468 639
rect 560 635 564 639
rect 672 635 676 639
rect 728 635 732 639
rect 776 635 780 639
rect 912 635 916 639
rect 944 635 948 639
rect 976 635 980 639
rect 1016 635 1020 639
rect 1056 635 1060 639
rect 1096 635 1100 639
rect 1136 635 1140 639
rect 1168 635 1172 639
rect 1232 635 1236 639
rect 1312 635 1316 639
rect 1447 631 1451 635
rect 416 627 420 631
rect 464 627 468 631
rect 560 627 564 631
rect 616 627 620 631
rect 672 627 676 631
rect 824 627 828 631
rect 872 627 876 631
rect 912 627 916 631
rect 944 627 948 631
rect 976 627 980 631
rect 1016 627 1020 631
rect 1056 627 1060 631
rect 1096 627 1100 631
rect 1168 627 1172 631
rect 1232 627 1236 631
rect 1312 627 1316 631
rect 376 623 380 627
rect 512 623 516 627
rect 728 623 732 627
rect 776 623 780 627
rect 1136 623 1140 627
rect 1200 623 1204 627
rect 1272 623 1276 627
rect 1352 623 1356 627
rect 344 619 348 623
rect 232 615 236 619
rect 280 611 284 615
rect 424 611 428 615
rect 448 611 452 615
rect 688 611 692 615
rect 984 611 988 615
rect 1200 611 1204 615
rect 111 605 115 609
rect 304 607 308 611
rect 328 607 332 611
rect 352 607 356 611
rect 376 607 380 611
rect 400 607 404 611
rect 488 607 492 611
rect 528 607 532 611
rect 576 607 580 611
rect 632 607 636 611
rect 744 607 748 611
rect 768 607 772 611
rect 792 607 796 611
rect 840 607 844 611
rect 888 607 892 611
rect 936 607 940 611
rect 1032 607 1036 611
rect 1080 607 1084 611
rect 1120 607 1124 611
rect 1160 607 1164 611
rect 1176 607 1180 611
rect 1248 607 1252 611
rect 1296 607 1300 611
rect 1344 607 1348 611
rect 280 599 284 603
rect 632 599 636 603
rect 688 599 692 603
rect 744 599 748 603
rect 888 599 892 603
rect 936 599 940 603
rect 984 599 988 603
rect 1032 599 1036 603
rect 1080 599 1084 603
rect 1120 599 1124 603
rect 1160 599 1164 603
rect 304 595 308 599
rect 400 595 404 599
rect 784 595 788 599
rect 792 595 796 599
rect 448 591 452 595
rect 111 587 115 591
rect 328 587 332 591
rect 352 587 356 591
rect 376 587 380 591
rect 488 587 492 591
rect 528 587 532 591
rect 424 583 428 587
rect 576 583 580 587
rect 840 583 844 587
rect 111 569 115 573
rect 784 571 788 575
rect 440 567 444 571
rect 1447 605 1451 609
rect 1200 599 1204 603
rect 1248 591 1252 595
rect 1296 587 1300 591
rect 1447 587 1451 591
rect 1344 583 1348 587
rect 1447 569 1451 573
rect 272 563 276 567
rect 560 563 564 567
rect 616 563 620 567
rect 840 563 844 567
rect 1080 563 1084 567
rect 1176 563 1180 567
rect 1192 563 1196 567
rect 296 555 300 559
rect 320 555 324 559
rect 344 555 348 559
rect 368 555 372 559
rect 392 555 396 559
rect 416 555 420 559
rect 472 555 476 559
rect 512 555 516 559
rect 672 555 676 559
rect 728 555 732 559
rect 896 555 900 559
rect 952 555 956 559
rect 1016 555 1020 559
rect 1136 555 1140 559
rect 1256 555 1260 559
rect 1320 555 1324 559
rect 1384 555 1388 559
rect 111 551 115 555
rect 1447 551 1451 555
rect 272 547 276 551
rect 296 547 300 551
rect 320 547 324 551
rect 344 547 348 551
rect 368 547 372 551
rect 392 547 396 551
rect 416 547 420 551
rect 440 547 444 551
rect 472 547 476 551
rect 560 547 564 551
rect 616 547 620 551
rect 672 547 676 551
rect 784 547 788 551
rect 840 547 844 551
rect 896 547 900 551
rect 952 547 956 551
rect 1136 547 1140 551
rect 1256 547 1260 551
rect 1320 547 1324 551
rect 1384 547 1388 551
rect 512 543 516 547
rect 728 543 732 547
rect 1016 543 1020 547
rect 1080 543 1084 547
rect 1192 543 1196 547
rect 400 531 404 535
rect 536 531 540 535
rect 632 531 636 535
rect 1032 531 1036 535
rect 1280 531 1284 535
rect 1400 531 1404 535
rect 111 525 115 529
rect 232 527 236 531
rect 256 527 260 531
rect 280 527 284 531
rect 304 527 308 531
rect 336 527 340 531
rect 368 527 372 531
rect 432 527 436 531
rect 464 527 468 531
rect 496 527 500 531
rect 584 527 588 531
rect 680 527 684 531
rect 720 527 724 531
rect 768 527 772 531
rect 816 527 820 531
rect 864 527 868 531
rect 920 527 924 531
rect 976 527 980 531
rect 1088 527 1092 531
rect 1136 527 1140 531
rect 1184 527 1188 531
rect 1232 527 1236 531
rect 1320 527 1324 531
rect 1360 527 1364 531
rect 1424 527 1428 531
rect 1447 525 1451 529
rect 304 519 308 523
rect 336 519 340 523
rect 368 519 372 523
rect 400 519 404 523
rect 432 519 436 523
rect 464 519 468 523
rect 496 519 500 523
rect 536 519 540 523
rect 720 519 724 523
rect 816 519 820 523
rect 864 519 868 523
rect 920 519 924 523
rect 1032 519 1036 523
rect 1088 519 1092 523
rect 1136 519 1140 523
rect 1184 519 1188 523
rect 1232 519 1236 523
rect 1280 519 1284 523
rect 1400 519 1404 523
rect 632 515 636 519
rect 280 511 284 515
rect 584 511 588 515
rect 768 511 772 515
rect 976 511 980 515
rect 1320 511 1324 515
rect 111 507 115 511
rect 1360 507 1364 511
rect 1447 507 1451 511
rect 232 503 236 507
rect 256 503 260 507
rect 680 503 684 507
rect 1424 503 1428 507
rect 111 489 115 493
rect 1447 489 1451 493
rect 144 483 148 487
rect 440 483 444 487
rect 552 483 556 487
rect 640 483 644 487
rect 672 483 676 487
rect 696 483 700 487
rect 768 483 772 487
rect 912 483 916 487
rect 1008 483 1012 487
rect 1104 483 1108 487
rect 1208 483 1212 487
rect 1320 483 1324 487
rect 1384 479 1388 483
rect 168 475 172 479
rect 192 475 196 479
rect 232 475 236 479
rect 280 475 284 479
rect 328 475 332 479
rect 384 475 388 479
rect 496 475 500 479
rect 600 475 604 479
rect 728 475 732 479
rect 808 475 812 479
rect 856 475 860 479
rect 960 475 964 479
rect 1056 475 1060 479
rect 1152 475 1156 479
rect 1264 475 1268 479
rect 1424 475 1428 479
rect 111 471 115 475
rect 1447 471 1451 475
rect 144 467 148 471
rect 168 467 172 471
rect 192 467 196 471
rect 232 467 236 471
rect 280 467 284 471
rect 328 467 332 471
rect 496 467 500 471
rect 600 467 604 471
rect 640 467 644 471
rect 696 467 700 471
rect 728 467 732 471
rect 808 467 812 471
rect 912 467 916 471
rect 960 467 964 471
rect 1056 467 1060 471
rect 1152 467 1156 471
rect 1264 467 1268 471
rect 1384 467 1388 471
rect 1424 467 1428 471
rect 384 463 388 467
rect 440 463 444 467
rect 552 463 556 467
rect 672 463 676 467
rect 768 463 772 467
rect 856 463 860 467
rect 1008 463 1012 467
rect 1024 463 1028 467
rect 1104 463 1108 467
rect 1208 463 1212 467
rect 1320 463 1324 467
rect 360 451 364 455
rect 800 451 804 455
rect 952 451 956 455
rect 111 445 115 449
rect 144 447 148 451
rect 168 447 172 451
rect 200 447 204 451
rect 248 447 252 451
rect 304 447 308 451
rect 424 447 428 451
rect 488 447 492 451
rect 552 447 556 451
rect 616 447 620 451
rect 680 447 684 451
rect 744 447 748 451
rect 848 447 852 451
rect 888 447 892 451
rect 920 447 924 451
rect 976 447 980 451
rect 1008 447 1012 451
rect 168 439 172 443
rect 200 439 204 443
rect 248 439 252 443
rect 304 439 308 443
rect 360 439 364 443
rect 424 439 428 443
rect 488 439 492 443
rect 552 439 556 443
rect 616 439 620 443
rect 680 439 684 443
rect 800 439 804 443
rect 848 439 852 443
rect 888 439 892 443
rect 952 439 956 443
rect 1008 439 1012 443
rect 144 431 148 435
rect 744 431 748 435
rect 920 431 924 435
rect 111 427 115 431
rect 976 423 980 427
rect 111 409 115 413
rect 144 403 148 407
rect 280 403 284 407
rect 400 403 404 407
rect 456 403 460 407
rect 984 403 988 407
rect 168 395 172 399
rect 192 395 196 399
rect 224 395 228 399
rect 336 395 340 399
rect 512 395 516 399
rect 560 395 564 399
rect 608 395 612 399
rect 656 395 660 399
rect 712 395 716 399
rect 776 395 780 399
rect 840 395 844 399
rect 912 395 916 399
rect 111 391 115 395
rect 144 387 148 391
rect 168 387 172 391
rect 192 387 196 391
rect 280 387 284 391
rect 336 387 340 391
rect 456 387 460 391
rect 512 387 516 391
rect 560 387 564 391
rect 608 387 612 391
rect 656 387 660 391
rect 776 387 780 391
rect 840 387 844 391
rect 984 387 988 391
rect 224 383 228 387
rect 400 383 404 387
rect 712 383 716 387
rect 912 383 916 387
rect 1040 447 1044 451
rect 1080 447 1084 451
rect 1128 447 1132 451
rect 1184 447 1188 451
rect 1248 447 1252 451
rect 1312 447 1316 451
rect 1376 447 1380 451
rect 1424 447 1428 451
rect 1447 445 1451 449
rect 1376 439 1380 443
rect 1040 431 1044 435
rect 1080 427 1084 431
rect 1128 427 1132 431
rect 1184 427 1188 431
rect 1447 427 1451 431
rect 1248 423 1252 427
rect 1312 423 1316 427
rect 1424 423 1428 427
rect 1328 411 1332 415
rect 1447 409 1451 413
rect 1112 403 1116 407
rect 1048 395 1052 399
rect 1168 395 1172 399
rect 1216 395 1220 399
rect 1256 395 1260 399
rect 1288 395 1292 399
rect 1368 395 1372 399
rect 1400 395 1404 399
rect 1424 395 1428 399
rect 1432 395 1436 399
rect 1048 387 1052 391
rect 1112 387 1116 391
rect 1168 387 1172 391
rect 1216 387 1220 391
rect 1256 387 1260 391
rect 1288 387 1292 391
rect 1328 387 1332 391
rect 1368 387 1372 391
rect 1424 387 1428 391
rect 1400 383 1404 387
rect 744 379 748 383
rect 1024 379 1028 383
rect 728 375 732 379
rect 1447 391 1451 395
rect 144 367 148 371
rect 736 367 740 371
rect 1240 367 1244 371
rect 1424 367 1428 371
rect 1432 367 1436 371
rect 111 361 115 365
rect 168 363 172 367
rect 192 363 196 367
rect 216 363 220 367
rect 240 363 244 367
rect 264 363 268 367
rect 304 363 308 367
rect 344 363 348 367
rect 384 363 388 367
rect 424 363 428 367
rect 464 363 468 367
rect 504 363 508 367
rect 544 363 548 367
rect 584 363 588 367
rect 624 363 628 367
rect 664 363 668 367
rect 696 363 700 367
rect 784 363 788 367
rect 840 363 844 367
rect 896 363 900 367
rect 960 363 964 367
rect 1024 363 1028 367
rect 1088 363 1092 367
rect 1144 363 1148 367
rect 1192 363 1196 367
rect 1280 363 1284 367
rect 1320 363 1324 367
rect 1360 363 1364 367
rect 1400 363 1404 367
rect 1447 361 1451 365
rect 144 355 148 359
rect 424 355 428 359
rect 464 355 468 359
rect 504 355 508 359
rect 584 355 588 359
rect 624 355 628 359
rect 664 355 668 359
rect 696 355 700 359
rect 784 355 788 359
rect 896 355 900 359
rect 960 355 964 359
rect 1024 355 1028 359
rect 1192 355 1196 359
rect 1240 355 1244 359
rect 1280 355 1284 359
rect 1424 355 1428 359
rect 168 347 172 351
rect 544 347 548 351
rect 736 347 740 351
rect 840 347 844 351
rect 1144 347 1148 351
rect 1320 347 1324 351
rect 1360 347 1364 351
rect 111 343 115 347
rect 192 343 196 347
rect 216 343 220 347
rect 240 343 244 347
rect 264 343 268 347
rect 304 343 308 347
rect 1447 343 1451 347
rect 344 339 348 343
rect 384 339 388 343
rect 1088 339 1092 343
rect 1120 339 1124 343
rect 1400 339 1404 343
rect 264 331 268 335
rect 111 325 115 329
rect 184 319 188 323
rect 232 319 236 323
rect 208 311 212 315
rect 216 311 220 315
rect 256 311 260 315
rect 111 307 115 311
rect 184 303 188 307
rect 208 303 212 307
rect 256 303 260 307
rect 232 299 236 303
rect 288 319 292 323
rect 368 319 372 323
rect 408 319 412 323
rect 536 319 540 323
rect 744 319 748 323
rect 1048 319 1052 323
rect 328 311 332 315
rect 448 311 452 315
rect 488 311 492 315
rect 592 311 596 315
rect 648 311 652 315
rect 696 311 700 315
rect 800 311 804 315
rect 856 311 860 315
rect 904 311 908 315
rect 952 311 956 315
rect 1000 311 1004 315
rect 1096 311 1100 315
rect 288 303 292 307
rect 328 303 332 307
rect 408 303 412 307
rect 448 303 452 307
rect 536 303 540 307
rect 592 303 596 307
rect 648 303 652 307
rect 744 303 748 307
rect 800 303 804 307
rect 856 303 860 307
rect 904 303 908 307
rect 952 303 956 307
rect 1048 303 1052 307
rect 1096 303 1100 307
rect 368 299 372 303
rect 488 299 492 303
rect 696 299 700 303
rect 1000 299 1004 303
rect 1288 327 1292 331
rect 1447 325 1451 329
rect 1144 311 1148 315
rect 1192 311 1196 315
rect 1240 311 1244 315
rect 1336 311 1340 315
rect 1392 311 1396 315
rect 1400 311 1404 315
rect 1424 311 1428 315
rect 1144 303 1148 307
rect 1192 303 1196 307
rect 1288 303 1292 307
rect 1392 303 1396 307
rect 1240 299 1244 303
rect 1336 299 1340 303
rect 1447 307 1451 311
rect 1424 299 1428 303
rect 264 295 268 299
rect 1120 295 1124 299
rect 1400 295 1404 299
rect 216 291 220 295
rect 256 287 260 291
rect 520 287 524 291
rect 1256 287 1260 291
rect 1424 287 1428 291
rect 111 281 115 285
rect 280 283 284 287
rect 304 283 308 287
rect 328 283 332 287
rect 352 283 356 287
rect 376 283 380 287
rect 408 283 412 287
rect 440 283 444 287
rect 480 283 484 287
rect 568 283 572 287
rect 624 283 628 287
rect 672 283 676 287
rect 720 283 724 287
rect 768 283 772 287
rect 816 283 820 287
rect 856 283 860 287
rect 888 283 892 287
rect 912 283 916 287
rect 936 283 940 287
rect 960 283 964 287
rect 984 283 988 287
rect 1008 283 1012 287
rect 1032 283 1036 287
rect 1056 283 1060 287
rect 1080 283 1084 287
rect 1104 283 1108 287
rect 1136 283 1140 287
rect 1168 283 1172 287
rect 1208 283 1212 287
rect 1312 283 1316 287
rect 1376 283 1380 287
rect 1447 281 1451 285
rect 256 275 260 279
rect 480 275 484 279
rect 520 275 524 279
rect 568 275 572 279
rect 624 275 628 279
rect 672 275 676 279
rect 720 275 724 279
rect 768 275 772 279
rect 816 275 820 279
rect 888 275 892 279
rect 912 275 916 279
rect 936 275 940 279
rect 960 275 964 279
rect 984 275 988 279
rect 1008 275 1012 279
rect 1032 275 1036 279
rect 1056 275 1060 279
rect 1080 275 1084 279
rect 1104 275 1108 279
rect 1136 275 1140 279
rect 1168 275 1172 279
rect 1208 275 1212 279
rect 1256 275 1260 279
rect 1312 275 1316 279
rect 304 271 308 275
rect 440 271 444 275
rect 1384 271 1388 275
rect 1424 271 1428 275
rect 280 267 284 271
rect 856 267 860 271
rect 111 263 115 267
rect 328 263 332 267
rect 352 263 356 267
rect 376 263 380 267
rect 408 263 412 267
rect 1376 263 1380 267
rect 111 245 115 249
rect 1288 247 1292 251
rect 296 239 300 243
rect 368 239 372 243
rect 440 239 444 243
rect 512 239 516 243
rect 632 239 636 243
rect 1048 239 1052 243
rect 592 235 596 239
rect 272 231 276 235
rect 320 231 324 235
rect 344 231 348 235
rect 392 231 396 235
rect 416 231 420 235
rect 472 231 476 235
rect 552 231 556 235
rect 688 231 692 235
rect 752 231 756 235
rect 816 231 820 235
rect 888 231 892 235
rect 968 231 972 235
rect 1128 231 1132 235
rect 1208 231 1212 235
rect 1368 231 1372 235
rect 111 227 115 231
rect 1447 263 1451 267
rect 1447 245 1451 249
rect 1424 231 1428 235
rect 1447 227 1451 231
rect 272 223 276 227
rect 296 223 300 227
rect 320 223 324 227
rect 344 223 348 227
rect 368 223 372 227
rect 392 223 396 227
rect 416 223 420 227
rect 472 223 476 227
rect 552 223 556 227
rect 632 223 636 227
rect 688 223 692 227
rect 752 223 756 227
rect 816 223 820 227
rect 888 223 892 227
rect 1128 223 1132 227
rect 1288 223 1292 227
rect 1368 223 1372 227
rect 1384 223 1388 227
rect 440 219 444 223
rect 512 219 516 223
rect 592 219 596 223
rect 968 219 972 223
rect 1048 219 1052 223
rect 1208 219 1212 223
rect 1424 219 1428 223
rect 392 207 396 211
rect 1424 207 1428 211
rect 111 201 115 205
rect 248 203 252 207
rect 272 203 276 207
rect 296 203 300 207
rect 320 203 324 207
rect 344 203 348 207
rect 368 203 372 207
rect 416 203 420 207
rect 440 203 444 207
rect 472 203 476 207
rect 520 203 524 207
rect 568 203 572 207
rect 624 203 628 207
rect 680 203 684 207
rect 728 203 732 207
rect 776 203 780 207
rect 824 203 828 207
rect 872 203 876 207
rect 928 203 932 207
rect 984 203 988 207
rect 1040 203 1044 207
rect 1072 203 1076 207
rect 1096 203 1100 207
rect 1144 203 1148 207
rect 1192 203 1196 207
rect 1240 203 1244 207
rect 1288 203 1292 207
rect 1336 203 1340 207
rect 1392 203 1396 207
rect 272 195 276 199
rect 296 195 300 199
rect 320 195 324 199
rect 344 195 348 199
rect 392 195 396 199
rect 416 195 420 199
rect 728 195 732 199
rect 776 195 780 199
rect 824 195 828 199
rect 872 195 876 199
rect 928 195 932 199
rect 984 195 988 199
rect 1040 195 1044 199
rect 368 187 372 191
rect 440 187 444 191
rect 111 183 115 187
rect 472 183 476 187
rect 520 183 524 187
rect 568 183 572 187
rect 624 183 628 187
rect 248 179 252 183
rect 680 179 684 183
rect 111 165 115 169
rect 192 159 196 163
rect 432 159 436 163
rect 536 159 540 163
rect 664 159 668 163
rect 832 159 836 163
rect 928 159 932 163
rect 1040 159 1044 163
rect 1447 201 1451 205
rect 1096 195 1100 199
rect 1144 195 1148 199
rect 1192 195 1196 199
rect 1336 195 1340 199
rect 1288 187 1292 191
rect 1392 187 1396 191
rect 1447 183 1451 187
rect 1240 179 1244 183
rect 1424 179 1428 183
rect 1368 167 1372 171
rect 1447 165 1451 169
rect 1136 159 1140 163
rect 1400 155 1404 159
rect 216 151 220 155
rect 248 151 252 155
rect 288 151 292 155
rect 336 151 340 155
rect 384 151 388 155
rect 480 151 484 155
rect 600 151 604 155
rect 720 151 724 155
rect 776 151 780 155
rect 880 151 884 155
rect 984 151 988 155
rect 1072 151 1076 155
rect 1088 151 1092 155
rect 1184 151 1188 155
rect 1200 151 1204 155
rect 1232 151 1236 155
rect 1272 151 1276 155
rect 1304 151 1308 155
rect 1336 151 1340 155
rect 1424 151 1428 155
rect 111 147 115 151
rect 192 143 196 147
rect 216 143 220 147
rect 248 143 252 147
rect 288 143 292 147
rect 336 143 340 147
rect 480 143 484 147
rect 600 143 604 147
rect 664 143 668 147
rect 720 143 724 147
rect 832 143 836 147
rect 880 143 884 147
rect 984 143 988 147
rect 1040 143 1044 147
rect 1088 143 1092 147
rect 1184 143 1188 147
rect 384 139 388 143
rect 432 139 436 143
rect 536 139 540 143
rect 776 139 780 143
rect 928 139 932 143
rect 1136 139 1140 143
rect 1447 147 1451 151
rect 1232 143 1236 147
rect 1272 143 1276 147
rect 1368 143 1372 147
rect 1400 143 1404 147
rect 1424 143 1428 147
rect 1304 139 1308 143
rect 1336 139 1340 143
rect 1200 123 1204 127
rect 408 115 412 119
rect 440 115 444 119
rect 1344 115 1348 119
rect 1424 115 1428 119
rect 111 109 115 113
rect 144 111 148 115
rect 168 111 172 115
rect 192 111 196 115
rect 216 111 220 115
rect 240 111 244 115
rect 264 111 268 115
rect 288 111 292 115
rect 312 111 316 115
rect 336 111 340 115
rect 360 111 364 115
rect 384 111 388 115
rect 472 111 476 115
rect 496 111 500 115
rect 520 111 524 115
rect 544 111 548 115
rect 568 111 572 115
rect 592 111 596 115
rect 616 111 620 115
rect 640 111 644 115
rect 664 111 668 115
rect 688 111 692 115
rect 712 111 716 115
rect 736 111 740 115
rect 760 111 764 115
rect 784 111 788 115
rect 808 111 812 115
rect 832 111 836 115
rect 864 111 868 115
rect 896 111 900 115
rect 928 111 932 115
rect 960 111 964 115
rect 992 111 996 115
rect 1024 111 1028 115
rect 1056 111 1060 115
rect 1080 111 1084 115
rect 1104 111 1108 115
rect 1128 111 1132 115
rect 1152 111 1156 115
rect 1184 111 1188 115
rect 1216 111 1220 115
rect 1248 111 1252 115
rect 1280 111 1284 115
rect 1312 111 1316 115
rect 1376 111 1380 115
rect 1400 111 1404 115
rect 1447 109 1451 113
rect 168 103 172 107
rect 192 103 196 107
rect 240 103 244 107
rect 312 103 316 107
rect 336 103 340 107
rect 360 103 364 107
rect 384 103 388 107
rect 408 103 412 107
rect 440 103 444 107
rect 472 103 476 107
rect 1056 103 1060 107
rect 1080 103 1084 107
rect 1104 103 1108 107
rect 1128 103 1132 107
rect 1152 103 1156 107
rect 1184 103 1188 107
rect 1216 103 1220 107
rect 1248 103 1252 107
rect 1280 103 1284 107
rect 1312 103 1316 107
rect 1344 103 1348 107
rect 1376 103 1380 107
rect 1424 103 1428 107
rect 216 95 220 99
rect 288 95 292 99
rect 496 95 500 99
rect 1400 95 1404 99
rect 111 91 115 95
rect 520 91 524 95
rect 544 91 548 95
rect 568 91 572 95
rect 592 91 596 95
rect 616 91 620 95
rect 640 91 644 95
rect 664 91 668 95
rect 688 91 692 95
rect 712 91 716 95
rect 736 91 740 95
rect 760 91 764 95
rect 784 91 788 95
rect 808 91 812 95
rect 832 91 836 95
rect 864 91 868 95
rect 896 91 900 95
rect 928 91 932 95
rect 960 91 964 95
rect 992 91 996 95
rect 1024 91 1028 95
rect 1447 91 1451 95
rect 264 87 268 91
<< m2 >>
rect 423 1511 429 1512
rect 423 1507 424 1511
rect 428 1510 429 1511
rect 818 1511 824 1512
rect 428 1508 659 1510
rect 428 1507 429 1508
rect 423 1506 429 1507
rect 657 1504 659 1508
rect 818 1507 819 1511
rect 823 1510 824 1511
rect 823 1508 899 1510
rect 823 1507 824 1508
rect 818 1506 824 1507
rect 897 1504 899 1508
rect 655 1503 661 1504
rect 895 1503 901 1504
rect 294 1502 300 1503
rect 294 1498 295 1502
rect 299 1498 300 1502
rect 318 1502 324 1503
rect 110 1497 116 1498
rect 294 1497 300 1498
rect 303 1499 309 1500
rect 110 1493 111 1497
rect 115 1493 116 1497
rect 303 1495 304 1499
rect 308 1495 309 1499
rect 318 1498 319 1502
rect 323 1498 324 1502
rect 342 1502 348 1503
rect 318 1497 324 1498
rect 327 1499 333 1500
rect 303 1494 309 1495
rect 327 1495 328 1499
rect 332 1498 333 1499
rect 342 1498 343 1502
rect 347 1498 348 1502
rect 366 1502 372 1503
rect 332 1496 338 1498
rect 342 1497 348 1498
rect 351 1499 357 1500
rect 332 1495 333 1496
rect 327 1494 333 1495
rect 110 1492 116 1493
rect 305 1490 307 1494
rect 327 1491 333 1492
rect 327 1490 328 1491
rect 305 1488 328 1490
rect 327 1487 328 1488
rect 332 1487 333 1491
rect 336 1490 338 1496
rect 351 1495 352 1499
rect 356 1498 357 1499
rect 366 1498 367 1502
rect 371 1498 372 1502
rect 406 1502 412 1503
rect 356 1496 362 1498
rect 366 1497 372 1498
rect 375 1499 381 1500
rect 356 1495 357 1496
rect 351 1494 357 1495
rect 351 1491 357 1492
rect 351 1490 352 1491
rect 336 1488 352 1490
rect 327 1486 333 1487
rect 351 1487 352 1488
rect 356 1487 357 1491
rect 360 1490 362 1496
rect 375 1495 376 1499
rect 380 1498 381 1499
rect 406 1498 407 1502
rect 411 1498 412 1502
rect 454 1502 460 1503
rect 380 1496 398 1498
rect 406 1497 412 1498
rect 415 1499 421 1500
rect 380 1495 381 1496
rect 375 1494 381 1495
rect 375 1491 381 1492
rect 375 1490 376 1491
rect 360 1488 376 1490
rect 351 1486 357 1487
rect 375 1487 376 1488
rect 380 1487 381 1491
rect 396 1490 398 1496
rect 415 1495 416 1499
rect 420 1498 421 1499
rect 454 1498 455 1502
rect 459 1498 460 1502
rect 510 1502 516 1503
rect 420 1496 442 1498
rect 454 1497 460 1498
rect 463 1499 469 1500
rect 420 1495 421 1496
rect 415 1494 421 1495
rect 415 1491 421 1492
rect 415 1490 416 1491
rect 396 1488 416 1490
rect 375 1486 381 1487
rect 415 1487 416 1488
rect 420 1487 421 1491
rect 440 1490 442 1496
rect 463 1495 464 1499
rect 468 1498 469 1499
rect 510 1498 511 1502
rect 515 1498 516 1502
rect 574 1502 580 1503
rect 468 1496 494 1498
rect 510 1497 516 1498
rect 519 1499 525 1500
rect 468 1495 469 1496
rect 463 1494 469 1495
rect 463 1491 469 1492
rect 463 1490 464 1491
rect 440 1488 464 1490
rect 415 1486 421 1487
rect 463 1487 464 1488
rect 468 1487 469 1491
rect 492 1490 494 1496
rect 519 1495 520 1499
rect 524 1498 525 1499
rect 574 1498 575 1502
rect 579 1498 580 1502
rect 646 1502 652 1503
rect 524 1496 554 1498
rect 574 1497 580 1498
rect 583 1499 589 1500
rect 524 1495 525 1496
rect 519 1494 525 1495
rect 519 1491 525 1492
rect 519 1490 520 1491
rect 492 1488 520 1490
rect 463 1486 469 1487
rect 519 1487 520 1488
rect 524 1487 525 1491
rect 552 1490 554 1496
rect 583 1495 584 1499
rect 588 1498 589 1499
rect 646 1498 647 1502
rect 651 1498 652 1502
rect 655 1499 656 1503
rect 660 1499 661 1503
rect 655 1498 661 1499
rect 726 1502 732 1503
rect 726 1498 727 1502
rect 731 1498 732 1502
rect 588 1496 622 1498
rect 646 1497 652 1498
rect 726 1497 732 1498
rect 806 1502 812 1503
rect 806 1498 807 1502
rect 811 1498 812 1502
rect 886 1502 892 1503
rect 806 1497 812 1498
rect 815 1499 821 1500
rect 588 1495 589 1496
rect 583 1494 589 1495
rect 583 1491 589 1492
rect 583 1490 584 1491
rect 552 1488 584 1490
rect 519 1486 525 1487
rect 583 1487 584 1488
rect 588 1487 589 1491
rect 620 1490 622 1496
rect 815 1495 816 1499
rect 820 1495 821 1499
rect 886 1498 887 1502
rect 891 1498 892 1502
rect 895 1499 896 1503
rect 900 1499 901 1503
rect 895 1498 901 1499
rect 958 1502 964 1503
rect 958 1498 959 1502
rect 963 1498 964 1502
rect 1030 1502 1036 1503
rect 886 1497 892 1498
rect 958 1497 964 1498
rect 967 1499 973 1500
rect 815 1494 821 1495
rect 967 1495 968 1499
rect 972 1495 973 1499
rect 1030 1498 1031 1502
rect 1035 1498 1036 1502
rect 1102 1502 1108 1503
rect 1030 1497 1036 1498
rect 1039 1499 1045 1500
rect 967 1494 973 1495
rect 1039 1495 1040 1499
rect 1044 1498 1045 1499
rect 1082 1499 1088 1500
rect 1082 1498 1083 1499
rect 1044 1496 1083 1498
rect 1044 1495 1045 1496
rect 1039 1494 1045 1495
rect 1082 1495 1083 1496
rect 1087 1495 1088 1499
rect 1102 1498 1103 1502
rect 1107 1498 1108 1502
rect 1174 1502 1180 1503
rect 1102 1497 1108 1498
rect 1111 1499 1120 1500
rect 1082 1494 1088 1495
rect 1111 1495 1112 1499
rect 1119 1495 1120 1499
rect 1174 1498 1175 1502
rect 1179 1498 1180 1502
rect 1246 1502 1252 1503
rect 1174 1497 1180 1498
rect 1183 1499 1189 1500
rect 1111 1494 1120 1495
rect 1183 1495 1184 1499
rect 1188 1495 1189 1499
rect 1246 1498 1247 1502
rect 1251 1498 1252 1502
rect 1246 1497 1252 1498
rect 1255 1499 1261 1500
rect 1183 1494 1189 1495
rect 1255 1495 1256 1499
rect 1260 1495 1261 1499
rect 1255 1494 1261 1495
rect 1446 1497 1452 1498
rect 655 1491 661 1492
rect 655 1490 656 1491
rect 620 1488 656 1490
rect 583 1486 589 1487
rect 655 1487 656 1488
rect 660 1487 661 1491
rect 655 1486 661 1487
rect 735 1491 741 1492
rect 735 1487 736 1491
rect 740 1490 741 1491
rect 816 1490 818 1494
rect 740 1488 818 1490
rect 895 1491 901 1492
rect 740 1487 741 1488
rect 735 1486 741 1487
rect 895 1487 896 1491
rect 900 1490 901 1491
rect 968 1490 970 1494
rect 900 1488 970 1490
rect 1039 1491 1045 1492
rect 900 1487 901 1488
rect 895 1486 901 1487
rect 1039 1487 1040 1491
rect 1044 1490 1045 1491
rect 1102 1491 1108 1492
rect 1102 1490 1103 1491
rect 1044 1488 1103 1490
rect 1044 1487 1045 1488
rect 1039 1486 1045 1487
rect 1102 1487 1103 1488
rect 1107 1487 1108 1491
rect 1102 1486 1108 1487
rect 1111 1487 1117 1488
rect 815 1483 824 1484
rect 110 1479 116 1480
rect 110 1475 111 1479
rect 115 1475 116 1479
rect 815 1479 816 1483
rect 823 1479 824 1483
rect 1111 1483 1112 1487
rect 1116 1486 1117 1487
rect 1184 1486 1186 1494
rect 1256 1486 1258 1494
rect 1446 1493 1447 1497
rect 1451 1493 1452 1497
rect 1446 1492 1452 1493
rect 1116 1484 1186 1486
rect 1220 1484 1258 1486
rect 1116 1483 1117 1484
rect 1111 1482 1117 1483
rect 815 1478 824 1479
rect 1183 1479 1189 1480
rect 110 1474 116 1475
rect 294 1476 300 1477
rect 318 1476 324 1477
rect 294 1472 295 1476
rect 299 1472 300 1476
rect 294 1471 300 1472
rect 303 1475 312 1476
rect 303 1471 304 1475
rect 311 1471 312 1475
rect 318 1472 319 1476
rect 323 1472 324 1476
rect 318 1471 324 1472
rect 342 1476 348 1477
rect 342 1472 343 1476
rect 347 1472 348 1476
rect 342 1471 348 1472
rect 366 1476 372 1477
rect 366 1472 367 1476
rect 371 1472 372 1476
rect 366 1471 372 1472
rect 406 1476 412 1477
rect 406 1472 407 1476
rect 411 1472 412 1476
rect 406 1471 412 1472
rect 454 1476 460 1477
rect 454 1472 455 1476
rect 459 1472 460 1476
rect 454 1471 460 1472
rect 510 1476 516 1477
rect 510 1472 511 1476
rect 515 1472 516 1476
rect 510 1471 516 1472
rect 574 1476 580 1477
rect 574 1472 575 1476
rect 579 1472 580 1476
rect 574 1471 580 1472
rect 646 1476 652 1477
rect 646 1472 647 1476
rect 651 1472 652 1476
rect 646 1471 652 1472
rect 726 1476 732 1477
rect 726 1472 727 1476
rect 731 1472 732 1476
rect 726 1471 732 1472
rect 806 1476 812 1477
rect 806 1472 807 1476
rect 811 1472 812 1476
rect 886 1476 892 1477
rect 886 1472 887 1476
rect 891 1472 892 1476
rect 806 1471 812 1472
rect 831 1471 837 1472
rect 886 1471 892 1472
rect 958 1476 964 1477
rect 1030 1476 1036 1477
rect 958 1472 959 1476
rect 963 1472 964 1476
rect 958 1471 964 1472
rect 967 1475 973 1476
rect 967 1471 968 1475
rect 972 1471 973 1475
rect 1030 1472 1031 1476
rect 1035 1472 1036 1476
rect 1030 1471 1036 1472
rect 1102 1476 1108 1477
rect 1102 1472 1103 1476
rect 1107 1472 1108 1476
rect 1102 1471 1108 1472
rect 1174 1476 1180 1477
rect 1174 1472 1175 1476
rect 1179 1472 1180 1476
rect 1183 1475 1184 1479
rect 1188 1478 1189 1479
rect 1220 1478 1222 1484
rect 1188 1476 1222 1478
rect 1446 1479 1452 1480
rect 1246 1476 1252 1477
rect 1188 1475 1189 1476
rect 1183 1474 1189 1475
rect 1174 1471 1180 1472
rect 1246 1472 1247 1476
rect 1251 1472 1252 1476
rect 1246 1471 1252 1472
rect 1255 1475 1261 1476
rect 1255 1471 1256 1475
rect 1260 1471 1261 1475
rect 1446 1475 1447 1479
rect 1451 1475 1452 1479
rect 1446 1474 1452 1475
rect 303 1470 312 1471
rect 831 1467 832 1471
rect 836 1470 837 1471
rect 967 1470 973 1471
rect 1255 1470 1261 1471
rect 836 1468 882 1470
rect 836 1467 837 1468
rect 831 1466 837 1467
rect 880 1466 882 1468
rect 896 1468 938 1470
rect 896 1466 898 1468
rect 150 1464 156 1465
rect 110 1461 116 1462
rect 110 1457 111 1461
rect 115 1457 116 1461
rect 150 1460 151 1464
rect 155 1460 156 1464
rect 150 1459 156 1460
rect 174 1464 180 1465
rect 174 1460 175 1464
rect 179 1460 180 1464
rect 174 1459 180 1460
rect 198 1464 204 1465
rect 198 1460 199 1464
rect 203 1460 204 1464
rect 198 1459 204 1460
rect 230 1464 236 1465
rect 230 1460 231 1464
rect 235 1460 236 1464
rect 230 1459 236 1460
rect 270 1464 276 1465
rect 270 1460 271 1464
rect 275 1460 276 1464
rect 270 1459 276 1460
rect 318 1464 324 1465
rect 318 1460 319 1464
rect 323 1460 324 1464
rect 318 1459 324 1460
rect 366 1464 372 1465
rect 366 1460 367 1464
rect 371 1460 372 1464
rect 366 1459 372 1460
rect 406 1464 412 1465
rect 454 1464 460 1465
rect 406 1460 407 1464
rect 411 1460 412 1464
rect 406 1459 412 1460
rect 415 1463 421 1464
rect 415 1459 416 1463
rect 420 1462 421 1463
rect 423 1463 429 1464
rect 423 1462 424 1463
rect 420 1460 424 1462
rect 420 1459 421 1460
rect 415 1458 421 1459
rect 423 1459 424 1460
rect 428 1459 429 1463
rect 454 1460 455 1464
rect 459 1460 460 1464
rect 454 1459 460 1460
rect 502 1464 508 1465
rect 502 1460 503 1464
rect 507 1460 508 1464
rect 502 1459 508 1460
rect 550 1464 556 1465
rect 550 1460 551 1464
rect 555 1460 556 1464
rect 550 1459 556 1460
rect 606 1464 612 1465
rect 606 1460 607 1464
rect 611 1460 612 1464
rect 606 1459 612 1460
rect 662 1464 668 1465
rect 662 1460 663 1464
rect 667 1460 668 1464
rect 662 1459 668 1460
rect 710 1464 716 1465
rect 710 1460 711 1464
rect 715 1460 716 1464
rect 710 1459 716 1460
rect 758 1464 764 1465
rect 758 1460 759 1464
rect 763 1460 764 1464
rect 758 1459 764 1460
rect 814 1464 820 1465
rect 814 1460 815 1464
rect 819 1460 820 1464
rect 814 1459 820 1460
rect 870 1464 876 1465
rect 880 1464 898 1466
rect 936 1466 938 1468
rect 968 1466 970 1470
rect 926 1464 932 1465
rect 936 1464 970 1466
rect 1231 1467 1237 1468
rect 974 1464 980 1465
rect 870 1460 871 1464
rect 875 1460 876 1464
rect 870 1459 876 1460
rect 926 1460 927 1464
rect 931 1460 932 1464
rect 926 1459 932 1460
rect 974 1460 975 1464
rect 979 1460 980 1464
rect 974 1459 980 1460
rect 1022 1464 1028 1465
rect 1022 1460 1023 1464
rect 1027 1460 1028 1464
rect 1022 1459 1028 1460
rect 1070 1464 1076 1465
rect 1118 1464 1124 1465
rect 1070 1460 1071 1464
rect 1075 1460 1076 1464
rect 1070 1459 1076 1460
rect 1079 1463 1088 1464
rect 1079 1459 1080 1463
rect 1087 1459 1088 1463
rect 1118 1460 1119 1464
rect 1123 1460 1124 1464
rect 1118 1459 1124 1460
rect 1166 1464 1172 1465
rect 1166 1460 1167 1464
rect 1171 1460 1172 1464
rect 1166 1459 1172 1460
rect 1214 1464 1220 1465
rect 1214 1460 1215 1464
rect 1219 1460 1220 1464
rect 1231 1463 1232 1467
rect 1236 1466 1237 1467
rect 1257 1466 1259 1470
rect 1236 1464 1259 1466
rect 1262 1464 1268 1465
rect 1236 1463 1237 1464
rect 1231 1462 1237 1463
rect 1214 1459 1220 1460
rect 1262 1460 1263 1464
rect 1267 1460 1268 1464
rect 1262 1459 1268 1460
rect 1310 1464 1316 1465
rect 1310 1460 1311 1464
rect 1315 1460 1316 1464
rect 1310 1459 1316 1460
rect 1446 1461 1452 1462
rect 423 1458 429 1459
rect 1079 1458 1088 1459
rect 110 1456 116 1457
rect 1446 1457 1447 1461
rect 1451 1457 1452 1461
rect 1446 1456 1452 1457
rect 159 1455 165 1456
rect 159 1451 160 1455
rect 164 1454 165 1455
rect 426 1455 432 1456
rect 426 1454 427 1455
rect 164 1452 427 1454
rect 164 1451 165 1452
rect 159 1450 165 1451
rect 426 1451 427 1452
rect 431 1451 432 1455
rect 426 1450 432 1451
rect 767 1455 773 1456
rect 767 1451 768 1455
rect 772 1454 773 1455
rect 826 1455 832 1456
rect 826 1454 827 1455
rect 772 1452 827 1454
rect 772 1451 773 1452
rect 767 1450 773 1451
rect 826 1451 827 1452
rect 831 1451 832 1455
rect 826 1450 832 1451
rect 935 1455 941 1456
rect 935 1451 936 1455
rect 940 1454 941 1455
rect 986 1455 992 1456
rect 986 1454 987 1455
rect 940 1452 987 1454
rect 940 1451 941 1452
rect 935 1450 941 1451
rect 986 1451 987 1452
rect 991 1451 992 1455
rect 986 1450 992 1451
rect 1175 1455 1181 1456
rect 1175 1451 1176 1455
rect 1180 1454 1181 1455
rect 1226 1455 1232 1456
rect 1226 1454 1227 1455
rect 1180 1452 1227 1454
rect 1180 1451 1181 1452
rect 1175 1450 1181 1451
rect 1226 1451 1227 1452
rect 1231 1451 1232 1455
rect 1226 1450 1232 1451
rect 1271 1455 1277 1456
rect 1271 1451 1272 1455
rect 1276 1454 1277 1455
rect 1322 1455 1328 1456
rect 1322 1454 1323 1455
rect 1276 1452 1323 1454
rect 1276 1451 1277 1452
rect 1271 1450 1277 1451
rect 1322 1451 1323 1452
rect 1327 1451 1328 1455
rect 1322 1450 1328 1451
rect 183 1447 189 1448
rect 183 1446 184 1447
rect 169 1444 184 1446
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 159 1439 165 1440
rect 110 1438 116 1439
rect 150 1438 156 1439
rect 150 1434 151 1438
rect 155 1434 156 1438
rect 159 1435 160 1439
rect 164 1438 165 1439
rect 169 1438 171 1444
rect 183 1443 184 1444
rect 188 1443 189 1447
rect 207 1447 213 1448
rect 207 1446 208 1447
rect 183 1442 189 1443
rect 193 1444 208 1446
rect 183 1439 189 1440
rect 164 1436 171 1438
rect 174 1438 180 1439
rect 164 1435 165 1436
rect 159 1434 165 1435
rect 174 1434 175 1438
rect 179 1434 180 1438
rect 183 1435 184 1439
rect 188 1438 189 1439
rect 193 1438 195 1444
rect 207 1443 208 1444
rect 212 1443 213 1447
rect 239 1447 245 1448
rect 239 1446 240 1447
rect 207 1442 213 1443
rect 225 1444 240 1446
rect 207 1439 213 1440
rect 188 1436 195 1438
rect 198 1438 204 1439
rect 188 1435 189 1436
rect 183 1434 189 1435
rect 198 1434 199 1438
rect 203 1434 204 1438
rect 207 1435 208 1439
rect 212 1438 213 1439
rect 225 1438 227 1444
rect 239 1443 240 1444
rect 244 1443 245 1447
rect 279 1447 285 1448
rect 279 1446 280 1447
rect 239 1442 245 1443
rect 260 1444 280 1446
rect 239 1439 245 1440
rect 212 1436 227 1438
rect 230 1438 236 1439
rect 212 1435 213 1436
rect 207 1434 213 1435
rect 230 1434 231 1438
rect 235 1434 236 1438
rect 239 1435 240 1439
rect 244 1438 245 1439
rect 260 1438 262 1444
rect 279 1443 280 1444
rect 284 1443 285 1447
rect 327 1447 333 1448
rect 327 1446 328 1447
rect 279 1442 285 1443
rect 300 1444 328 1446
rect 279 1439 285 1440
rect 244 1436 262 1438
rect 270 1438 276 1439
rect 244 1435 245 1436
rect 239 1434 245 1435
rect 270 1434 271 1438
rect 275 1434 276 1438
rect 279 1435 280 1439
rect 284 1438 285 1439
rect 300 1438 302 1444
rect 327 1443 328 1444
rect 332 1443 333 1447
rect 375 1447 381 1448
rect 375 1446 376 1447
rect 327 1442 333 1443
rect 352 1444 376 1446
rect 327 1439 333 1440
rect 284 1436 302 1438
rect 318 1438 324 1439
rect 284 1435 285 1436
rect 279 1434 285 1435
rect 318 1434 319 1438
rect 323 1434 324 1438
rect 327 1435 328 1439
rect 332 1438 333 1439
rect 352 1438 354 1444
rect 375 1443 376 1444
rect 380 1443 381 1447
rect 463 1447 469 1448
rect 463 1446 464 1447
rect 375 1442 381 1443
rect 424 1444 464 1446
rect 415 1439 421 1440
rect 332 1436 354 1438
rect 366 1438 372 1439
rect 332 1435 333 1436
rect 327 1434 333 1435
rect 366 1434 367 1438
rect 371 1434 372 1438
rect 406 1438 412 1439
rect 150 1433 156 1434
rect 174 1433 180 1434
rect 198 1433 204 1434
rect 230 1433 236 1434
rect 270 1433 276 1434
rect 318 1433 324 1434
rect 366 1433 372 1434
rect 375 1435 381 1436
rect 206 1431 212 1432
rect 206 1427 207 1431
rect 211 1430 212 1431
rect 298 1431 304 1432
rect 298 1430 299 1431
rect 211 1428 299 1430
rect 211 1427 212 1428
rect 206 1426 212 1427
rect 298 1427 299 1428
rect 303 1427 304 1431
rect 298 1426 304 1427
rect 306 1431 312 1432
rect 306 1427 307 1431
rect 311 1430 312 1431
rect 375 1431 376 1435
rect 380 1431 381 1435
rect 406 1434 407 1438
rect 411 1434 412 1438
rect 415 1435 416 1439
rect 420 1438 421 1439
rect 424 1438 426 1444
rect 463 1443 464 1444
rect 468 1443 469 1447
rect 511 1447 517 1448
rect 511 1446 512 1447
rect 463 1442 469 1443
rect 488 1444 512 1446
rect 463 1439 469 1440
rect 420 1436 426 1438
rect 454 1438 460 1439
rect 420 1435 421 1436
rect 415 1434 421 1435
rect 454 1434 455 1438
rect 459 1434 460 1438
rect 463 1435 464 1439
rect 468 1438 469 1439
rect 488 1438 490 1444
rect 511 1443 512 1444
rect 516 1443 517 1447
rect 559 1447 565 1448
rect 559 1446 560 1447
rect 511 1442 517 1443
rect 536 1444 560 1446
rect 511 1439 517 1440
rect 468 1436 490 1438
rect 502 1438 508 1439
rect 468 1435 469 1436
rect 463 1434 469 1435
rect 502 1434 503 1438
rect 507 1434 508 1438
rect 511 1435 512 1439
rect 516 1438 517 1439
rect 536 1438 538 1444
rect 559 1443 560 1444
rect 564 1443 565 1447
rect 615 1447 621 1448
rect 615 1446 616 1447
rect 559 1442 565 1443
rect 588 1444 616 1446
rect 559 1439 565 1440
rect 516 1436 538 1438
rect 550 1438 556 1439
rect 516 1435 517 1436
rect 511 1434 517 1435
rect 550 1434 551 1438
rect 555 1434 556 1438
rect 559 1435 560 1439
rect 564 1438 565 1439
rect 588 1438 590 1444
rect 615 1443 616 1444
rect 620 1443 621 1447
rect 671 1447 677 1448
rect 671 1446 672 1447
rect 615 1442 621 1443
rect 644 1444 672 1446
rect 615 1439 621 1440
rect 564 1436 590 1438
rect 606 1438 612 1439
rect 564 1435 565 1436
rect 559 1434 565 1435
rect 606 1434 607 1438
rect 611 1434 612 1438
rect 615 1435 616 1439
rect 620 1438 621 1439
rect 644 1438 646 1444
rect 671 1443 672 1444
rect 676 1443 677 1447
rect 719 1447 725 1448
rect 719 1446 720 1447
rect 671 1442 677 1443
rect 696 1444 720 1446
rect 671 1439 677 1440
rect 620 1436 646 1438
rect 662 1438 668 1439
rect 620 1435 621 1436
rect 615 1434 621 1435
rect 662 1434 663 1438
rect 667 1434 668 1438
rect 671 1435 672 1439
rect 676 1438 677 1439
rect 696 1438 698 1444
rect 719 1443 720 1444
rect 724 1443 725 1447
rect 719 1442 725 1443
rect 823 1447 829 1448
rect 823 1443 824 1447
rect 828 1446 829 1447
rect 879 1447 885 1448
rect 828 1444 854 1446
rect 828 1443 829 1444
rect 823 1442 829 1443
rect 823 1439 832 1440
rect 676 1436 698 1438
rect 710 1438 716 1439
rect 676 1435 677 1436
rect 671 1434 677 1435
rect 710 1434 711 1438
rect 715 1434 716 1438
rect 758 1438 764 1439
rect 406 1433 412 1434
rect 454 1433 460 1434
rect 502 1433 508 1434
rect 550 1433 556 1434
rect 606 1433 612 1434
rect 662 1433 668 1434
rect 710 1433 716 1434
rect 719 1435 725 1436
rect 375 1430 381 1431
rect 558 1431 564 1432
rect 311 1428 321 1430
rect 311 1427 312 1428
rect 306 1426 312 1427
rect 319 1426 321 1428
rect 336 1428 378 1430
rect 336 1426 338 1428
rect 558 1427 559 1431
rect 563 1430 564 1431
rect 719 1431 720 1435
rect 724 1431 725 1435
rect 758 1434 759 1438
rect 763 1434 764 1438
rect 814 1438 820 1439
rect 758 1433 764 1434
rect 767 1435 773 1436
rect 719 1430 725 1431
rect 767 1431 768 1435
rect 772 1434 773 1435
rect 814 1434 815 1438
rect 819 1434 820 1438
rect 823 1435 824 1439
rect 831 1435 832 1439
rect 823 1434 832 1435
rect 772 1432 810 1434
rect 814 1433 820 1434
rect 772 1431 773 1432
rect 767 1430 773 1431
rect 808 1430 810 1432
rect 831 1431 837 1432
rect 831 1430 832 1431
rect 563 1428 723 1430
rect 808 1428 832 1430
rect 563 1427 564 1428
rect 558 1426 564 1427
rect 831 1427 832 1428
rect 836 1427 837 1431
rect 852 1430 854 1444
rect 879 1443 880 1447
rect 884 1446 885 1447
rect 983 1447 989 1448
rect 884 1444 938 1446
rect 884 1443 885 1444
rect 879 1442 885 1443
rect 936 1440 938 1444
rect 983 1443 984 1447
rect 988 1446 989 1447
rect 1031 1447 1040 1448
rect 988 1444 1011 1446
rect 988 1443 989 1444
rect 983 1442 989 1443
rect 935 1439 941 1440
rect 983 1439 992 1440
rect 870 1438 876 1439
rect 870 1434 871 1438
rect 875 1434 876 1438
rect 926 1438 932 1439
rect 870 1433 876 1434
rect 879 1435 885 1436
rect 879 1431 880 1435
rect 884 1431 885 1435
rect 926 1434 927 1438
rect 931 1434 932 1438
rect 935 1435 936 1439
rect 940 1435 941 1439
rect 935 1434 941 1435
rect 974 1438 980 1439
rect 974 1434 975 1438
rect 979 1434 980 1438
rect 983 1435 984 1439
rect 991 1435 992 1439
rect 983 1434 992 1435
rect 926 1433 932 1434
rect 974 1433 980 1434
rect 879 1430 885 1431
rect 1009 1430 1011 1444
rect 1031 1443 1032 1447
rect 1039 1443 1040 1447
rect 1127 1447 1133 1448
rect 1127 1446 1128 1447
rect 1031 1442 1040 1443
rect 1104 1444 1128 1446
rect 1079 1439 1085 1440
rect 1022 1438 1028 1439
rect 1022 1434 1023 1438
rect 1027 1434 1028 1438
rect 1070 1438 1076 1439
rect 1022 1433 1028 1434
rect 1031 1435 1037 1436
rect 1031 1431 1032 1435
rect 1036 1431 1037 1435
rect 1070 1434 1071 1438
rect 1075 1434 1076 1438
rect 1079 1435 1080 1439
rect 1084 1438 1085 1439
rect 1104 1438 1106 1444
rect 1127 1443 1128 1444
rect 1132 1443 1133 1447
rect 1127 1442 1133 1443
rect 1223 1447 1229 1448
rect 1223 1443 1224 1447
rect 1228 1446 1229 1447
rect 1274 1447 1280 1448
rect 1228 1444 1250 1446
rect 1228 1443 1229 1444
rect 1223 1442 1229 1443
rect 1223 1439 1232 1440
rect 1084 1436 1106 1438
rect 1118 1438 1124 1439
rect 1084 1435 1085 1436
rect 1079 1434 1085 1435
rect 1118 1434 1119 1438
rect 1123 1434 1124 1438
rect 1166 1438 1172 1439
rect 1070 1433 1076 1434
rect 1118 1433 1124 1434
rect 1127 1435 1136 1436
rect 1031 1430 1037 1431
rect 1127 1431 1128 1435
rect 1135 1431 1136 1435
rect 1166 1434 1167 1438
rect 1171 1434 1172 1438
rect 1214 1438 1220 1439
rect 1166 1433 1172 1434
rect 1175 1435 1181 1436
rect 1127 1430 1136 1431
rect 1175 1431 1176 1435
rect 1180 1431 1181 1435
rect 1214 1434 1215 1438
rect 1219 1434 1220 1438
rect 1223 1435 1224 1439
rect 1231 1435 1232 1439
rect 1223 1434 1232 1435
rect 1214 1433 1220 1434
rect 1175 1430 1181 1431
rect 1231 1431 1237 1432
rect 1231 1430 1232 1431
rect 852 1428 882 1430
rect 1009 1428 1034 1430
rect 1177 1428 1232 1430
rect 831 1426 837 1427
rect 1231 1427 1232 1428
rect 1236 1427 1237 1431
rect 1248 1430 1250 1444
rect 1274 1443 1275 1447
rect 1279 1446 1280 1447
rect 1319 1447 1325 1448
rect 1319 1446 1320 1447
rect 1279 1444 1320 1446
rect 1279 1443 1280 1444
rect 1274 1442 1280 1443
rect 1319 1443 1320 1444
rect 1324 1443 1325 1447
rect 1319 1442 1325 1443
rect 1446 1443 1452 1444
rect 1319 1439 1328 1440
rect 1262 1438 1268 1439
rect 1262 1434 1263 1438
rect 1267 1434 1268 1438
rect 1310 1438 1316 1439
rect 1262 1433 1268 1434
rect 1271 1435 1277 1436
rect 1271 1431 1272 1435
rect 1276 1431 1277 1435
rect 1310 1434 1311 1438
rect 1315 1434 1316 1438
rect 1319 1435 1320 1439
rect 1327 1435 1328 1439
rect 1446 1439 1447 1443
rect 1451 1439 1452 1443
rect 1446 1438 1452 1439
rect 1319 1434 1328 1435
rect 1310 1433 1316 1434
rect 1271 1430 1277 1431
rect 1354 1431 1360 1432
rect 1248 1428 1274 1430
rect 1231 1426 1237 1427
rect 1354 1427 1355 1431
rect 1359 1430 1360 1431
rect 1359 1428 1403 1430
rect 1359 1427 1360 1428
rect 1354 1426 1360 1427
rect 319 1424 338 1426
rect 1401 1424 1403 1428
rect 423 1423 432 1424
rect 1031 1423 1040 1424
rect 1271 1423 1280 1424
rect 1399 1423 1405 1424
rect 134 1422 140 1423
rect 134 1418 135 1422
rect 139 1418 140 1422
rect 158 1422 164 1423
rect 110 1417 116 1418
rect 134 1417 140 1418
rect 143 1419 149 1420
rect 110 1413 111 1417
rect 115 1413 116 1417
rect 143 1415 144 1419
rect 148 1415 149 1419
rect 158 1418 159 1422
rect 163 1418 164 1422
rect 182 1422 188 1423
rect 158 1417 164 1418
rect 167 1419 173 1420
rect 143 1414 149 1415
rect 167 1415 168 1419
rect 172 1415 173 1419
rect 182 1418 183 1422
rect 187 1418 188 1422
rect 222 1422 228 1423
rect 182 1417 188 1418
rect 191 1419 197 1420
rect 167 1414 173 1415
rect 191 1415 192 1419
rect 196 1418 197 1419
rect 222 1418 223 1422
rect 227 1418 228 1422
rect 286 1422 292 1423
rect 196 1416 214 1418
rect 222 1417 228 1418
rect 231 1419 237 1420
rect 196 1415 197 1416
rect 191 1414 197 1415
rect 110 1412 116 1413
rect 145 1406 147 1414
rect 169 1410 171 1414
rect 191 1411 197 1412
rect 191 1410 192 1411
rect 169 1408 192 1410
rect 191 1407 192 1408
rect 196 1407 197 1411
rect 212 1410 214 1416
rect 231 1415 232 1419
rect 236 1418 237 1419
rect 286 1418 287 1422
rect 291 1418 292 1422
rect 350 1422 356 1423
rect 236 1416 270 1418
rect 286 1417 292 1418
rect 295 1419 301 1420
rect 236 1415 237 1416
rect 231 1414 237 1415
rect 231 1411 237 1412
rect 231 1410 232 1411
rect 212 1408 232 1410
rect 191 1406 197 1407
rect 231 1407 232 1408
rect 236 1407 237 1411
rect 268 1410 270 1416
rect 295 1415 296 1419
rect 300 1418 301 1419
rect 350 1418 351 1422
rect 355 1418 356 1422
rect 414 1422 420 1423
rect 300 1416 321 1418
rect 350 1417 356 1418
rect 359 1419 365 1420
rect 300 1415 301 1416
rect 295 1414 301 1415
rect 295 1411 301 1412
rect 295 1410 296 1411
rect 268 1408 296 1410
rect 231 1406 237 1407
rect 295 1407 296 1408
rect 300 1407 301 1411
rect 319 1410 321 1416
rect 359 1415 360 1419
rect 364 1418 365 1419
rect 414 1418 415 1422
rect 419 1418 420 1422
rect 423 1419 424 1423
rect 431 1419 432 1423
rect 423 1418 432 1419
rect 478 1422 484 1423
rect 478 1418 479 1422
rect 483 1418 484 1422
rect 534 1422 540 1423
rect 364 1416 394 1418
rect 414 1417 420 1418
rect 478 1417 484 1418
rect 487 1419 493 1420
rect 364 1415 365 1416
rect 359 1414 365 1415
rect 359 1411 365 1412
rect 359 1410 360 1411
rect 319 1408 360 1410
rect 295 1406 301 1407
rect 359 1407 360 1408
rect 364 1407 365 1411
rect 392 1410 394 1416
rect 487 1415 488 1419
rect 492 1418 493 1419
rect 519 1419 525 1420
rect 519 1418 520 1419
rect 492 1416 520 1418
rect 492 1415 493 1416
rect 487 1414 493 1415
rect 519 1415 520 1416
rect 524 1415 525 1419
rect 534 1418 535 1422
rect 539 1418 540 1422
rect 582 1422 588 1423
rect 534 1417 540 1418
rect 543 1419 549 1420
rect 519 1414 525 1415
rect 543 1415 544 1419
rect 548 1418 549 1419
rect 582 1418 583 1422
rect 587 1418 588 1422
rect 630 1422 636 1423
rect 548 1416 570 1418
rect 582 1417 588 1418
rect 591 1419 597 1420
rect 548 1415 549 1416
rect 543 1414 549 1415
rect 423 1411 429 1412
rect 423 1410 424 1411
rect 392 1408 424 1410
rect 359 1406 365 1407
rect 423 1407 424 1408
rect 428 1407 429 1411
rect 423 1406 429 1407
rect 543 1411 549 1412
rect 543 1407 544 1411
rect 548 1410 549 1411
rect 558 1411 564 1412
rect 558 1410 559 1411
rect 548 1408 559 1410
rect 548 1407 549 1408
rect 543 1406 549 1407
rect 558 1407 559 1408
rect 563 1407 564 1411
rect 558 1406 564 1407
rect 568 1406 570 1416
rect 591 1415 592 1419
rect 596 1415 597 1419
rect 630 1418 631 1422
rect 635 1418 636 1422
rect 686 1422 692 1423
rect 630 1417 636 1418
rect 639 1419 645 1420
rect 591 1414 597 1415
rect 639 1415 640 1419
rect 644 1418 645 1419
rect 686 1418 687 1422
rect 691 1418 692 1422
rect 742 1422 748 1423
rect 644 1416 670 1418
rect 686 1417 692 1418
rect 695 1419 701 1420
rect 644 1415 645 1416
rect 639 1414 645 1415
rect 593 1410 595 1414
rect 639 1411 645 1412
rect 639 1410 640 1411
rect 593 1408 640 1410
rect 639 1407 640 1408
rect 644 1407 645 1411
rect 668 1410 670 1416
rect 695 1415 696 1419
rect 700 1418 701 1419
rect 742 1418 743 1422
rect 747 1418 748 1422
rect 798 1422 804 1423
rect 700 1416 726 1418
rect 742 1417 748 1418
rect 751 1419 757 1420
rect 700 1415 701 1416
rect 695 1414 701 1415
rect 695 1411 701 1412
rect 695 1410 696 1411
rect 668 1408 696 1410
rect 639 1406 645 1407
rect 695 1407 696 1408
rect 700 1407 701 1411
rect 724 1410 726 1416
rect 751 1415 752 1419
rect 756 1418 757 1419
rect 798 1418 799 1422
rect 803 1418 804 1422
rect 854 1422 860 1423
rect 756 1416 782 1418
rect 798 1417 804 1418
rect 807 1419 813 1420
rect 756 1415 757 1416
rect 751 1414 757 1415
rect 751 1411 757 1412
rect 751 1410 752 1411
rect 724 1408 752 1410
rect 695 1406 701 1407
rect 751 1407 752 1408
rect 756 1407 757 1411
rect 780 1410 782 1416
rect 807 1415 808 1419
rect 812 1418 813 1419
rect 854 1418 855 1422
rect 859 1418 860 1422
rect 910 1422 916 1423
rect 812 1416 838 1418
rect 854 1417 860 1418
rect 863 1419 869 1420
rect 812 1415 813 1416
rect 807 1414 813 1415
rect 807 1411 813 1412
rect 807 1410 808 1411
rect 780 1408 808 1410
rect 751 1406 757 1407
rect 807 1407 808 1408
rect 812 1407 813 1411
rect 836 1410 838 1416
rect 863 1415 864 1419
rect 868 1418 869 1419
rect 890 1419 896 1420
rect 890 1418 891 1419
rect 868 1416 891 1418
rect 868 1415 869 1416
rect 863 1414 869 1415
rect 890 1415 891 1416
rect 895 1415 896 1419
rect 910 1418 911 1422
rect 915 1418 916 1422
rect 966 1422 972 1423
rect 910 1417 916 1418
rect 919 1419 925 1420
rect 890 1414 896 1415
rect 919 1415 920 1419
rect 924 1418 925 1419
rect 966 1418 967 1422
rect 971 1418 972 1422
rect 1022 1422 1028 1423
rect 924 1416 950 1418
rect 966 1417 972 1418
rect 975 1419 981 1420
rect 924 1415 925 1416
rect 919 1414 925 1415
rect 863 1411 869 1412
rect 863 1410 864 1411
rect 836 1408 864 1410
rect 807 1406 813 1407
rect 863 1407 864 1408
rect 868 1407 869 1411
rect 948 1410 950 1416
rect 975 1415 976 1419
rect 980 1418 981 1419
rect 1022 1418 1023 1422
rect 1027 1418 1028 1422
rect 1031 1419 1032 1423
rect 1039 1419 1040 1423
rect 1031 1418 1040 1419
rect 1070 1422 1076 1423
rect 1070 1418 1071 1422
rect 1075 1418 1076 1422
rect 1118 1422 1124 1423
rect 980 1416 1006 1418
rect 1022 1417 1028 1418
rect 1070 1417 1076 1418
rect 1079 1419 1088 1420
rect 980 1415 981 1416
rect 975 1414 981 1415
rect 975 1411 981 1412
rect 975 1410 976 1411
rect 948 1408 976 1410
rect 863 1406 869 1407
rect 975 1407 976 1408
rect 980 1407 981 1411
rect 1004 1410 1006 1416
rect 1079 1415 1080 1419
rect 1087 1415 1088 1419
rect 1118 1418 1119 1422
rect 1123 1418 1124 1422
rect 1166 1422 1172 1423
rect 1118 1417 1124 1418
rect 1127 1419 1133 1420
rect 1079 1414 1088 1415
rect 1127 1415 1128 1419
rect 1132 1418 1133 1419
rect 1138 1419 1144 1420
rect 1138 1418 1139 1419
rect 1132 1416 1139 1418
rect 1132 1415 1133 1416
rect 1127 1414 1133 1415
rect 1138 1415 1139 1416
rect 1143 1415 1144 1419
rect 1166 1418 1167 1422
rect 1171 1418 1172 1422
rect 1214 1422 1220 1423
rect 1166 1417 1172 1418
rect 1175 1419 1181 1420
rect 1138 1414 1144 1415
rect 1175 1415 1176 1419
rect 1180 1418 1181 1419
rect 1214 1418 1215 1422
rect 1219 1418 1220 1422
rect 1262 1422 1268 1423
rect 1180 1416 1202 1418
rect 1214 1417 1220 1418
rect 1223 1419 1229 1420
rect 1180 1415 1181 1416
rect 1175 1414 1181 1415
rect 1031 1411 1037 1412
rect 1031 1410 1032 1411
rect 1004 1408 1032 1410
rect 975 1406 981 1407
rect 1031 1407 1032 1408
rect 1036 1407 1037 1411
rect 1127 1411 1136 1412
rect 1031 1406 1037 1407
rect 1079 1407 1085 1408
rect 145 1404 171 1406
rect 568 1404 595 1406
rect 167 1403 173 1404
rect 110 1399 116 1400
rect 110 1395 111 1399
rect 115 1395 116 1399
rect 167 1399 168 1403
rect 172 1399 173 1403
rect 167 1398 173 1399
rect 591 1403 597 1404
rect 591 1399 592 1403
rect 596 1399 597 1403
rect 1079 1403 1080 1407
rect 1084 1406 1085 1407
rect 1118 1407 1124 1408
rect 1118 1406 1119 1407
rect 1084 1404 1119 1406
rect 1084 1403 1085 1404
rect 1079 1402 1085 1403
rect 1118 1403 1119 1404
rect 1123 1403 1124 1407
rect 1127 1407 1128 1411
rect 1135 1407 1136 1411
rect 1200 1410 1202 1416
rect 1223 1415 1224 1419
rect 1228 1418 1229 1419
rect 1262 1418 1263 1422
rect 1267 1418 1268 1422
rect 1271 1419 1272 1423
rect 1279 1419 1280 1423
rect 1271 1418 1280 1419
rect 1302 1422 1308 1423
rect 1302 1418 1303 1422
rect 1307 1418 1308 1422
rect 1342 1422 1348 1423
rect 1228 1416 1250 1418
rect 1262 1417 1268 1418
rect 1302 1417 1308 1418
rect 1311 1419 1320 1420
rect 1228 1415 1229 1416
rect 1223 1414 1229 1415
rect 1223 1411 1229 1412
rect 1223 1410 1224 1411
rect 1200 1408 1224 1410
rect 1127 1406 1136 1407
rect 1223 1407 1224 1408
rect 1228 1407 1229 1411
rect 1248 1410 1250 1416
rect 1311 1415 1312 1419
rect 1319 1415 1320 1419
rect 1342 1418 1343 1422
rect 1347 1418 1348 1422
rect 1390 1422 1396 1423
rect 1342 1417 1348 1418
rect 1351 1419 1357 1420
rect 1311 1414 1320 1415
rect 1351 1415 1352 1419
rect 1356 1415 1357 1419
rect 1390 1418 1391 1422
rect 1395 1418 1396 1422
rect 1399 1419 1400 1423
rect 1404 1419 1405 1423
rect 1399 1418 1405 1419
rect 1414 1422 1420 1423
rect 1414 1418 1415 1422
rect 1419 1418 1420 1422
rect 1390 1417 1396 1418
rect 1414 1417 1420 1418
rect 1423 1419 1429 1420
rect 1351 1414 1357 1415
rect 1423 1415 1424 1419
rect 1428 1415 1429 1419
rect 1423 1414 1429 1415
rect 1446 1417 1452 1418
rect 1271 1411 1277 1412
rect 1271 1410 1272 1411
rect 1248 1408 1272 1410
rect 1223 1406 1229 1407
rect 1271 1407 1272 1408
rect 1276 1407 1277 1411
rect 1271 1406 1277 1407
rect 1311 1411 1317 1412
rect 1311 1407 1312 1411
rect 1316 1410 1317 1411
rect 1352 1410 1354 1414
rect 1316 1408 1354 1410
rect 1399 1411 1405 1412
rect 1316 1407 1317 1408
rect 1311 1406 1317 1407
rect 1399 1407 1400 1411
rect 1404 1410 1405 1411
rect 1425 1410 1427 1414
rect 1446 1413 1447 1417
rect 1451 1413 1452 1417
rect 1446 1412 1452 1413
rect 1404 1408 1427 1410
rect 1404 1407 1405 1408
rect 1399 1406 1405 1407
rect 1118 1402 1124 1403
rect 1351 1403 1360 1404
rect 591 1398 597 1399
rect 1351 1399 1352 1403
rect 1359 1399 1360 1403
rect 1351 1398 1360 1399
rect 1446 1399 1452 1400
rect 110 1394 116 1395
rect 134 1396 140 1397
rect 158 1396 164 1397
rect 134 1392 135 1396
rect 139 1392 140 1396
rect 134 1391 140 1392
rect 143 1395 152 1396
rect 143 1391 144 1395
rect 151 1391 152 1395
rect 158 1392 159 1396
rect 163 1392 164 1396
rect 158 1391 164 1392
rect 182 1396 188 1397
rect 182 1392 183 1396
rect 187 1392 188 1396
rect 182 1391 188 1392
rect 222 1396 228 1397
rect 222 1392 223 1396
rect 227 1392 228 1396
rect 222 1391 228 1392
rect 286 1396 292 1397
rect 286 1392 287 1396
rect 291 1392 292 1396
rect 286 1391 292 1392
rect 350 1396 356 1397
rect 350 1392 351 1396
rect 355 1392 356 1396
rect 350 1391 356 1392
rect 414 1396 420 1397
rect 414 1392 415 1396
rect 419 1392 420 1396
rect 414 1391 420 1392
rect 478 1396 484 1397
rect 534 1396 540 1397
rect 478 1392 479 1396
rect 483 1392 484 1396
rect 478 1391 484 1392
rect 487 1395 493 1396
rect 487 1391 488 1395
rect 492 1394 493 1395
rect 511 1395 517 1396
rect 511 1394 512 1395
rect 492 1392 512 1394
rect 492 1391 493 1392
rect 143 1390 152 1391
rect 487 1390 493 1391
rect 511 1391 512 1392
rect 516 1391 517 1395
rect 534 1392 535 1396
rect 539 1392 540 1396
rect 534 1391 540 1392
rect 582 1396 588 1397
rect 582 1392 583 1396
rect 587 1392 588 1396
rect 582 1391 588 1392
rect 630 1396 636 1397
rect 630 1392 631 1396
rect 635 1392 636 1396
rect 630 1391 636 1392
rect 686 1396 692 1397
rect 686 1392 687 1396
rect 691 1392 692 1396
rect 686 1391 692 1392
rect 742 1396 748 1397
rect 742 1392 743 1396
rect 747 1392 748 1396
rect 742 1391 748 1392
rect 798 1396 804 1397
rect 798 1392 799 1396
rect 803 1392 804 1396
rect 798 1391 804 1392
rect 854 1396 860 1397
rect 854 1392 855 1396
rect 859 1392 860 1396
rect 854 1391 860 1392
rect 910 1396 916 1397
rect 966 1396 972 1397
rect 910 1392 911 1396
rect 915 1392 916 1396
rect 910 1391 916 1392
rect 919 1395 925 1396
rect 919 1391 920 1395
rect 924 1394 925 1395
rect 946 1395 952 1396
rect 946 1394 947 1395
rect 924 1392 947 1394
rect 924 1391 925 1392
rect 511 1390 517 1391
rect 919 1390 925 1391
rect 946 1391 947 1392
rect 951 1391 952 1395
rect 966 1392 967 1396
rect 971 1392 972 1396
rect 966 1391 972 1392
rect 1022 1396 1028 1397
rect 1022 1392 1023 1396
rect 1027 1392 1028 1396
rect 1022 1391 1028 1392
rect 1070 1396 1076 1397
rect 1070 1392 1071 1396
rect 1075 1392 1076 1396
rect 1070 1391 1076 1392
rect 1118 1396 1124 1397
rect 1118 1392 1119 1396
rect 1123 1392 1124 1396
rect 1118 1391 1124 1392
rect 1166 1396 1172 1397
rect 1214 1396 1220 1397
rect 1166 1392 1167 1396
rect 1171 1392 1172 1396
rect 1166 1391 1172 1392
rect 1175 1395 1181 1396
rect 1175 1391 1176 1395
rect 1180 1394 1181 1395
rect 1206 1395 1212 1396
rect 1206 1394 1207 1395
rect 1180 1392 1207 1394
rect 1180 1391 1181 1392
rect 946 1390 952 1391
rect 1175 1390 1181 1391
rect 1206 1391 1207 1392
rect 1211 1391 1212 1395
rect 1214 1392 1215 1396
rect 1219 1392 1220 1396
rect 1214 1391 1220 1392
rect 1262 1396 1268 1397
rect 1262 1392 1263 1396
rect 1267 1392 1268 1396
rect 1262 1391 1268 1392
rect 1302 1396 1308 1397
rect 1302 1392 1303 1396
rect 1307 1392 1308 1396
rect 1302 1391 1308 1392
rect 1342 1396 1348 1397
rect 1342 1392 1343 1396
rect 1347 1392 1348 1396
rect 1342 1391 1348 1392
rect 1390 1396 1396 1397
rect 1390 1392 1391 1396
rect 1395 1392 1396 1396
rect 1390 1391 1396 1392
rect 1414 1396 1420 1397
rect 1414 1392 1415 1396
rect 1419 1392 1420 1396
rect 1414 1391 1420 1392
rect 1423 1395 1432 1396
rect 1423 1391 1424 1395
rect 1431 1391 1432 1395
rect 1446 1395 1447 1399
rect 1451 1395 1452 1399
rect 1446 1394 1452 1395
rect 1206 1390 1212 1391
rect 1423 1390 1432 1391
rect 134 1384 140 1385
rect 110 1381 116 1382
rect 110 1377 111 1381
rect 115 1377 116 1381
rect 134 1380 135 1384
rect 139 1380 140 1384
rect 134 1379 140 1380
rect 158 1384 164 1385
rect 158 1380 159 1384
rect 163 1380 164 1384
rect 158 1379 164 1380
rect 182 1384 188 1385
rect 182 1380 183 1384
rect 187 1380 188 1384
rect 182 1379 188 1380
rect 230 1384 236 1385
rect 230 1380 231 1384
rect 235 1380 236 1384
rect 230 1379 236 1380
rect 278 1384 284 1385
rect 278 1380 279 1384
rect 283 1380 284 1384
rect 278 1379 284 1380
rect 334 1384 340 1385
rect 334 1380 335 1384
rect 339 1380 340 1384
rect 334 1379 340 1380
rect 390 1384 396 1385
rect 390 1380 391 1384
rect 395 1380 396 1384
rect 390 1379 396 1380
rect 438 1384 444 1385
rect 438 1380 439 1384
rect 443 1380 444 1384
rect 438 1379 444 1380
rect 486 1384 492 1385
rect 486 1380 487 1384
rect 491 1380 492 1384
rect 486 1379 492 1380
rect 526 1384 532 1385
rect 526 1380 527 1384
rect 531 1380 532 1384
rect 526 1379 532 1380
rect 566 1384 572 1385
rect 566 1380 567 1384
rect 571 1380 572 1384
rect 566 1379 572 1380
rect 614 1384 620 1385
rect 614 1380 615 1384
rect 619 1380 620 1384
rect 614 1379 620 1380
rect 662 1384 668 1385
rect 662 1380 663 1384
rect 667 1380 668 1384
rect 662 1379 668 1380
rect 710 1384 716 1385
rect 710 1380 711 1384
rect 715 1380 716 1384
rect 710 1379 716 1380
rect 766 1384 772 1385
rect 766 1380 767 1384
rect 771 1380 772 1384
rect 766 1379 772 1380
rect 822 1384 828 1385
rect 822 1380 823 1384
rect 827 1380 828 1384
rect 822 1379 828 1380
rect 878 1384 884 1385
rect 934 1384 940 1385
rect 878 1380 879 1384
rect 883 1380 884 1384
rect 878 1379 884 1380
rect 887 1383 896 1384
rect 887 1379 888 1383
rect 895 1379 896 1383
rect 934 1380 935 1384
rect 939 1380 940 1384
rect 934 1379 940 1380
rect 990 1384 996 1385
rect 990 1380 991 1384
rect 995 1380 996 1384
rect 990 1379 996 1380
rect 1046 1384 1052 1385
rect 1094 1384 1100 1385
rect 1046 1380 1047 1384
rect 1051 1380 1052 1384
rect 1046 1379 1052 1380
rect 1055 1383 1061 1384
rect 1055 1379 1056 1383
rect 1060 1382 1061 1383
rect 1082 1383 1088 1384
rect 1082 1382 1083 1383
rect 1060 1380 1083 1382
rect 1060 1379 1061 1380
rect 887 1378 896 1379
rect 1055 1378 1061 1379
rect 1082 1379 1083 1380
rect 1087 1379 1088 1383
rect 1094 1380 1095 1384
rect 1099 1380 1100 1384
rect 1094 1379 1100 1380
rect 1142 1384 1148 1385
rect 1142 1380 1143 1384
rect 1147 1380 1148 1384
rect 1142 1379 1148 1380
rect 1190 1384 1196 1385
rect 1190 1380 1191 1384
rect 1195 1380 1196 1384
rect 1190 1379 1196 1380
rect 1238 1384 1244 1385
rect 1238 1380 1239 1384
rect 1243 1380 1244 1384
rect 1238 1379 1244 1380
rect 1286 1384 1292 1385
rect 1334 1384 1340 1385
rect 1286 1380 1287 1384
rect 1291 1380 1292 1384
rect 1286 1379 1292 1380
rect 1295 1383 1301 1384
rect 1295 1379 1296 1383
rect 1300 1382 1301 1383
rect 1314 1383 1320 1384
rect 1314 1382 1315 1383
rect 1300 1380 1315 1382
rect 1300 1379 1301 1380
rect 1082 1378 1088 1379
rect 1295 1378 1301 1379
rect 1314 1379 1315 1380
rect 1319 1379 1320 1383
rect 1334 1380 1335 1384
rect 1339 1380 1340 1384
rect 1334 1379 1340 1380
rect 1382 1384 1388 1385
rect 1382 1380 1383 1384
rect 1387 1380 1388 1384
rect 1382 1379 1388 1380
rect 1414 1384 1420 1385
rect 1414 1380 1415 1384
rect 1419 1380 1420 1384
rect 1414 1379 1420 1380
rect 1446 1381 1452 1382
rect 1314 1378 1320 1379
rect 110 1376 116 1377
rect 1446 1377 1447 1381
rect 1451 1377 1452 1381
rect 1446 1376 1452 1377
rect 143 1375 149 1376
rect 143 1371 144 1375
rect 148 1374 149 1375
rect 170 1375 176 1376
rect 170 1374 171 1375
rect 148 1372 171 1374
rect 148 1371 149 1372
rect 143 1370 149 1371
rect 170 1371 171 1372
rect 175 1371 176 1375
rect 194 1375 200 1376
rect 194 1374 195 1375
rect 170 1370 176 1371
rect 184 1372 195 1374
rect 167 1367 173 1368
rect 110 1363 116 1364
rect 110 1359 111 1363
rect 115 1359 116 1363
rect 167 1363 168 1367
rect 172 1366 173 1367
rect 184 1366 186 1372
rect 194 1371 195 1372
rect 199 1371 200 1375
rect 194 1370 200 1371
rect 239 1375 245 1376
rect 239 1371 240 1375
rect 244 1374 245 1375
rect 290 1375 296 1376
rect 290 1374 291 1375
rect 244 1372 291 1374
rect 244 1371 245 1372
rect 239 1370 245 1371
rect 290 1371 291 1372
rect 295 1371 296 1375
rect 290 1370 296 1371
rect 298 1375 304 1376
rect 298 1371 299 1375
rect 303 1374 304 1375
rect 343 1375 349 1376
rect 343 1374 344 1375
rect 303 1372 344 1374
rect 303 1371 304 1372
rect 298 1370 304 1371
rect 343 1371 344 1372
rect 348 1371 349 1375
rect 343 1370 349 1371
rect 399 1375 405 1376
rect 399 1371 400 1375
rect 404 1374 405 1375
rect 450 1375 456 1376
rect 450 1374 451 1375
rect 404 1372 451 1374
rect 404 1371 405 1372
rect 399 1370 405 1371
rect 450 1371 451 1372
rect 455 1371 456 1375
rect 450 1370 456 1371
rect 495 1375 501 1376
rect 495 1371 496 1375
rect 500 1374 501 1375
rect 538 1375 544 1376
rect 538 1374 539 1375
rect 500 1372 539 1374
rect 500 1371 501 1372
rect 495 1370 501 1371
rect 538 1371 539 1372
rect 543 1371 544 1375
rect 538 1370 544 1371
rect 575 1375 581 1376
rect 575 1371 576 1375
rect 580 1374 581 1375
rect 626 1375 632 1376
rect 626 1374 627 1375
rect 580 1372 627 1374
rect 580 1371 581 1372
rect 575 1370 581 1371
rect 626 1371 627 1372
rect 631 1371 632 1375
rect 626 1370 632 1371
rect 639 1375 645 1376
rect 639 1371 640 1375
rect 644 1374 645 1375
rect 671 1375 677 1376
rect 644 1372 666 1374
rect 644 1371 645 1372
rect 639 1370 645 1371
rect 172 1364 186 1366
rect 191 1367 197 1368
rect 172 1363 173 1364
rect 167 1362 173 1363
rect 191 1363 192 1367
rect 196 1366 197 1367
rect 287 1367 293 1368
rect 196 1364 227 1366
rect 196 1363 197 1364
rect 191 1362 197 1363
rect 143 1359 152 1360
rect 167 1359 176 1360
rect 191 1359 200 1360
rect 110 1358 116 1359
rect 134 1358 140 1359
rect 134 1354 135 1358
rect 139 1354 140 1358
rect 143 1355 144 1359
rect 151 1355 152 1359
rect 143 1354 152 1355
rect 158 1358 164 1359
rect 158 1354 159 1358
rect 163 1354 164 1358
rect 167 1355 168 1359
rect 175 1355 176 1359
rect 167 1354 176 1355
rect 182 1358 188 1359
rect 182 1354 183 1358
rect 187 1354 188 1358
rect 191 1355 192 1359
rect 199 1355 200 1359
rect 191 1354 200 1355
rect 134 1353 140 1354
rect 158 1353 164 1354
rect 182 1353 188 1354
rect 206 1351 212 1352
rect 206 1350 207 1351
rect 177 1348 207 1350
rect 177 1344 179 1348
rect 206 1347 207 1348
rect 211 1347 212 1351
rect 225 1350 227 1364
rect 287 1363 288 1367
rect 292 1366 293 1367
rect 447 1367 453 1368
rect 292 1364 347 1366
rect 292 1363 293 1364
rect 287 1362 293 1363
rect 345 1360 347 1364
rect 447 1363 448 1367
rect 452 1366 453 1367
rect 519 1367 525 1368
rect 452 1364 498 1366
rect 452 1363 453 1364
rect 447 1362 453 1363
rect 496 1360 498 1364
rect 519 1363 520 1367
rect 524 1366 525 1367
rect 535 1367 541 1368
rect 535 1366 536 1367
rect 524 1364 536 1366
rect 524 1363 525 1364
rect 519 1362 525 1363
rect 535 1363 536 1364
rect 540 1363 541 1367
rect 535 1362 541 1363
rect 623 1367 629 1368
rect 623 1363 624 1367
rect 628 1366 629 1367
rect 664 1366 666 1372
rect 671 1371 672 1375
rect 676 1374 677 1375
rect 722 1375 728 1376
rect 722 1374 723 1375
rect 676 1372 723 1374
rect 676 1371 677 1372
rect 671 1370 677 1371
rect 722 1371 723 1372
rect 727 1371 728 1375
rect 722 1370 728 1371
rect 775 1375 781 1376
rect 775 1371 776 1375
rect 780 1374 781 1375
rect 834 1375 840 1376
rect 834 1374 835 1375
rect 780 1372 835 1374
rect 780 1371 781 1372
rect 775 1370 781 1371
rect 834 1371 835 1372
rect 839 1371 840 1375
rect 834 1370 840 1371
rect 943 1375 949 1376
rect 943 1371 944 1375
rect 948 1374 949 1375
rect 1002 1375 1008 1376
rect 1002 1374 1003 1375
rect 948 1372 1003 1374
rect 948 1371 949 1372
rect 943 1370 949 1371
rect 1002 1371 1003 1372
rect 1007 1371 1008 1375
rect 1002 1370 1008 1371
rect 1394 1375 1400 1376
rect 1394 1371 1395 1375
rect 1399 1374 1400 1375
rect 1426 1375 1432 1376
rect 1426 1374 1427 1375
rect 1399 1372 1427 1374
rect 1399 1371 1400 1372
rect 1394 1370 1400 1371
rect 1426 1371 1427 1372
rect 1431 1371 1432 1375
rect 1426 1370 1432 1371
rect 719 1367 725 1368
rect 719 1366 720 1367
rect 628 1364 659 1366
rect 664 1364 720 1366
rect 628 1363 629 1364
rect 623 1362 629 1363
rect 287 1359 296 1360
rect 343 1359 349 1360
rect 447 1359 456 1360
rect 495 1359 501 1360
rect 535 1359 544 1360
rect 623 1359 632 1360
rect 230 1358 236 1359
rect 230 1354 231 1358
rect 235 1354 236 1358
rect 278 1358 284 1359
rect 230 1353 236 1354
rect 239 1355 245 1356
rect 239 1351 240 1355
rect 244 1351 245 1355
rect 278 1354 279 1358
rect 283 1354 284 1358
rect 287 1355 288 1359
rect 295 1355 296 1359
rect 287 1354 296 1355
rect 334 1358 340 1359
rect 334 1354 335 1358
rect 339 1354 340 1358
rect 343 1355 344 1359
rect 348 1355 349 1359
rect 343 1354 349 1355
rect 390 1358 396 1359
rect 390 1354 391 1358
rect 395 1354 396 1358
rect 438 1358 444 1359
rect 278 1353 284 1354
rect 334 1353 340 1354
rect 390 1353 396 1354
rect 399 1355 405 1356
rect 239 1350 245 1351
rect 247 1351 253 1352
rect 225 1348 242 1350
rect 206 1346 212 1347
rect 247 1347 248 1351
rect 252 1350 253 1351
rect 318 1351 324 1352
rect 252 1348 290 1350
rect 252 1347 253 1348
rect 247 1346 253 1347
rect 288 1344 290 1348
rect 318 1347 319 1351
rect 323 1350 324 1351
rect 399 1351 400 1355
rect 404 1354 405 1355
rect 438 1354 439 1358
rect 443 1354 444 1358
rect 447 1355 448 1359
rect 455 1355 456 1359
rect 447 1354 456 1355
rect 486 1358 492 1359
rect 486 1354 487 1358
rect 491 1354 492 1358
rect 495 1355 496 1359
rect 500 1355 501 1359
rect 495 1354 501 1355
rect 526 1358 532 1359
rect 526 1354 527 1358
rect 531 1354 532 1358
rect 535 1355 536 1359
rect 543 1355 544 1359
rect 535 1354 544 1355
rect 566 1358 572 1359
rect 566 1354 567 1358
rect 571 1354 572 1358
rect 614 1358 620 1359
rect 404 1352 434 1354
rect 438 1353 444 1354
rect 486 1353 492 1354
rect 526 1353 532 1354
rect 566 1353 572 1354
rect 575 1355 581 1356
rect 404 1351 405 1352
rect 399 1350 405 1351
rect 432 1350 434 1352
rect 494 1351 500 1352
rect 494 1350 495 1351
rect 323 1348 347 1350
rect 432 1348 495 1350
rect 323 1347 324 1348
rect 318 1346 324 1347
rect 345 1344 347 1348
rect 494 1347 495 1348
rect 499 1347 500 1351
rect 494 1346 500 1347
rect 511 1351 517 1352
rect 511 1347 512 1351
rect 516 1350 517 1351
rect 575 1351 576 1355
rect 580 1351 581 1355
rect 614 1354 615 1358
rect 619 1354 620 1358
rect 623 1355 624 1359
rect 631 1355 632 1359
rect 623 1354 632 1355
rect 614 1353 620 1354
rect 575 1350 581 1351
rect 639 1351 645 1352
rect 639 1350 640 1351
rect 516 1348 578 1350
rect 624 1348 640 1350
rect 516 1347 517 1348
rect 511 1346 517 1347
rect 175 1343 181 1344
rect 287 1343 293 1344
rect 343 1343 349 1344
rect 583 1343 589 1344
rect 166 1342 172 1343
rect 166 1338 167 1342
rect 171 1338 172 1342
rect 175 1339 176 1343
rect 180 1339 181 1343
rect 175 1338 181 1339
rect 190 1342 196 1343
rect 190 1338 191 1342
rect 195 1338 196 1342
rect 230 1342 236 1343
rect 110 1337 116 1338
rect 166 1337 172 1338
rect 190 1337 196 1338
rect 199 1339 205 1340
rect 110 1333 111 1337
rect 115 1333 116 1337
rect 199 1335 200 1339
rect 204 1335 205 1339
rect 230 1338 231 1342
rect 235 1338 236 1342
rect 278 1342 284 1343
rect 230 1337 236 1338
rect 239 1339 245 1340
rect 199 1334 205 1335
rect 239 1335 240 1339
rect 244 1335 245 1339
rect 278 1338 279 1342
rect 283 1338 284 1342
rect 287 1339 288 1343
rect 292 1339 293 1343
rect 287 1338 293 1339
rect 334 1342 340 1343
rect 334 1338 335 1342
rect 339 1338 340 1342
rect 343 1339 344 1343
rect 348 1339 349 1343
rect 343 1338 349 1339
rect 390 1342 396 1343
rect 390 1338 391 1342
rect 395 1338 396 1342
rect 454 1342 460 1343
rect 278 1337 284 1338
rect 334 1337 340 1338
rect 390 1337 396 1338
rect 399 1339 405 1340
rect 239 1334 245 1335
rect 399 1335 400 1339
rect 404 1338 405 1339
rect 410 1339 416 1340
rect 410 1338 411 1339
rect 404 1336 411 1338
rect 404 1335 405 1336
rect 399 1334 405 1335
rect 410 1335 411 1336
rect 415 1335 416 1339
rect 454 1338 455 1342
rect 459 1338 460 1342
rect 518 1342 524 1343
rect 454 1337 460 1338
rect 463 1339 469 1340
rect 410 1334 416 1335
rect 463 1335 464 1339
rect 468 1335 469 1339
rect 518 1338 519 1342
rect 523 1338 524 1342
rect 574 1342 580 1343
rect 518 1337 524 1338
rect 527 1339 533 1340
rect 463 1334 469 1335
rect 527 1335 528 1339
rect 532 1335 533 1339
rect 574 1338 575 1342
rect 579 1338 580 1342
rect 583 1339 584 1343
rect 588 1342 589 1343
rect 624 1342 626 1348
rect 639 1347 640 1348
rect 644 1347 645 1351
rect 657 1350 659 1364
rect 719 1363 720 1364
rect 724 1363 725 1367
rect 719 1362 725 1363
rect 831 1367 837 1368
rect 831 1363 832 1367
rect 836 1366 837 1367
rect 999 1367 1005 1368
rect 836 1364 890 1366
rect 836 1363 837 1364
rect 831 1362 837 1363
rect 888 1360 890 1364
rect 999 1363 1000 1367
rect 1004 1366 1005 1367
rect 1018 1367 1024 1368
rect 1018 1366 1019 1367
rect 1004 1364 1019 1366
rect 1004 1363 1005 1364
rect 999 1362 1005 1363
rect 1018 1363 1019 1364
rect 1023 1363 1024 1367
rect 1103 1367 1109 1368
rect 1103 1366 1104 1367
rect 1018 1362 1024 1363
rect 1080 1364 1104 1366
rect 719 1359 728 1360
rect 831 1359 840 1360
rect 887 1359 893 1360
rect 943 1359 952 1360
rect 999 1359 1008 1360
rect 1055 1359 1061 1360
rect 662 1358 668 1359
rect 662 1354 663 1358
rect 667 1354 668 1358
rect 710 1358 716 1359
rect 662 1353 668 1354
rect 671 1355 677 1356
rect 671 1351 672 1355
rect 676 1351 677 1355
rect 710 1354 711 1358
rect 715 1354 716 1358
rect 719 1355 720 1359
rect 727 1355 728 1359
rect 719 1354 728 1355
rect 766 1358 772 1359
rect 766 1354 767 1358
rect 771 1354 772 1358
rect 822 1358 828 1359
rect 710 1353 716 1354
rect 766 1353 772 1354
rect 775 1355 781 1356
rect 671 1350 677 1351
rect 690 1351 696 1352
rect 657 1348 674 1350
rect 639 1346 645 1347
rect 690 1347 691 1351
rect 695 1350 696 1351
rect 775 1351 776 1355
rect 780 1351 781 1355
rect 822 1354 823 1358
rect 827 1354 828 1358
rect 831 1355 832 1359
rect 839 1355 840 1359
rect 831 1354 840 1355
rect 878 1358 884 1359
rect 878 1354 879 1358
rect 883 1354 884 1358
rect 887 1355 888 1359
rect 892 1355 893 1359
rect 887 1354 893 1355
rect 934 1358 940 1359
rect 934 1354 935 1358
rect 939 1354 940 1358
rect 943 1355 944 1359
rect 951 1355 952 1359
rect 943 1354 952 1355
rect 990 1358 996 1359
rect 990 1354 991 1358
rect 995 1354 996 1358
rect 999 1355 1000 1359
rect 1007 1355 1008 1359
rect 999 1354 1008 1355
rect 1046 1358 1052 1359
rect 1046 1354 1047 1358
rect 1051 1354 1052 1358
rect 1055 1355 1056 1359
rect 1060 1358 1061 1359
rect 1080 1358 1082 1364
rect 1103 1363 1104 1364
rect 1108 1363 1109 1367
rect 1103 1362 1109 1363
rect 1151 1367 1157 1368
rect 1151 1363 1152 1367
rect 1156 1366 1157 1367
rect 1170 1367 1176 1368
rect 1170 1366 1171 1367
rect 1156 1364 1171 1366
rect 1156 1363 1157 1364
rect 1151 1362 1157 1363
rect 1170 1363 1171 1364
rect 1175 1363 1176 1367
rect 1199 1367 1205 1368
rect 1199 1366 1200 1367
rect 1170 1362 1176 1363
rect 1180 1364 1200 1366
rect 1151 1359 1157 1360
rect 1060 1356 1082 1358
rect 1094 1358 1100 1359
rect 1060 1355 1061 1356
rect 1055 1354 1061 1355
rect 1094 1354 1095 1358
rect 1099 1354 1100 1358
rect 1142 1358 1148 1359
rect 822 1353 828 1354
rect 878 1353 884 1354
rect 934 1353 940 1354
rect 990 1353 996 1354
rect 1046 1353 1052 1354
rect 1094 1353 1100 1354
rect 1103 1355 1109 1356
rect 775 1350 781 1351
rect 1103 1351 1104 1355
rect 1108 1354 1109 1355
rect 1114 1355 1120 1356
rect 1114 1354 1115 1355
rect 1108 1352 1115 1354
rect 1108 1351 1109 1352
rect 1103 1350 1109 1351
rect 1114 1351 1115 1352
rect 1119 1351 1120 1355
rect 1142 1354 1143 1358
rect 1147 1354 1148 1358
rect 1151 1355 1152 1359
rect 1156 1358 1157 1359
rect 1180 1358 1182 1364
rect 1199 1363 1200 1364
rect 1204 1363 1205 1367
rect 1247 1367 1253 1368
rect 1247 1366 1248 1367
rect 1199 1362 1205 1363
rect 1224 1364 1248 1366
rect 1199 1359 1205 1360
rect 1156 1356 1182 1358
rect 1190 1358 1196 1359
rect 1156 1355 1157 1356
rect 1151 1354 1157 1355
rect 1190 1354 1191 1358
rect 1195 1354 1196 1358
rect 1199 1355 1200 1359
rect 1204 1358 1205 1359
rect 1224 1358 1226 1364
rect 1247 1363 1248 1364
rect 1252 1363 1253 1367
rect 1343 1367 1349 1368
rect 1343 1366 1344 1367
rect 1247 1362 1253 1363
rect 1321 1364 1344 1366
rect 1295 1359 1301 1360
rect 1204 1356 1226 1358
rect 1238 1358 1244 1359
rect 1204 1355 1205 1356
rect 1199 1354 1205 1355
rect 1238 1354 1239 1358
rect 1243 1354 1244 1358
rect 1286 1358 1292 1359
rect 1142 1353 1148 1354
rect 1190 1353 1196 1354
rect 1238 1353 1244 1354
rect 1247 1355 1253 1356
rect 1114 1350 1120 1351
rect 1206 1351 1212 1352
rect 695 1348 779 1350
rect 695 1347 696 1348
rect 690 1346 696 1347
rect 1206 1347 1207 1351
rect 1211 1350 1212 1351
rect 1247 1351 1248 1355
rect 1252 1351 1253 1355
rect 1286 1354 1287 1358
rect 1291 1354 1292 1358
rect 1295 1355 1296 1359
rect 1300 1358 1301 1359
rect 1321 1358 1323 1364
rect 1343 1363 1344 1364
rect 1348 1363 1349 1367
rect 1343 1362 1349 1363
rect 1391 1367 1397 1368
rect 1391 1363 1392 1367
rect 1396 1366 1397 1367
rect 1423 1367 1432 1368
rect 1396 1364 1410 1366
rect 1396 1363 1397 1364
rect 1391 1362 1397 1363
rect 1391 1359 1400 1360
rect 1300 1356 1323 1358
rect 1334 1358 1340 1359
rect 1300 1355 1301 1356
rect 1295 1354 1301 1355
rect 1334 1354 1335 1358
rect 1339 1354 1340 1358
rect 1382 1358 1388 1359
rect 1286 1353 1292 1354
rect 1334 1353 1340 1354
rect 1343 1355 1349 1356
rect 1247 1350 1253 1351
rect 1343 1351 1344 1355
rect 1348 1354 1349 1355
rect 1374 1355 1380 1356
rect 1374 1354 1375 1355
rect 1348 1352 1375 1354
rect 1348 1351 1349 1352
rect 1343 1350 1349 1351
rect 1374 1351 1375 1352
rect 1379 1351 1380 1355
rect 1382 1354 1383 1358
rect 1387 1354 1388 1358
rect 1391 1355 1392 1359
rect 1399 1355 1400 1359
rect 1391 1354 1400 1355
rect 1382 1353 1388 1354
rect 1374 1350 1380 1351
rect 1408 1350 1410 1364
rect 1423 1363 1424 1367
rect 1431 1363 1432 1367
rect 1423 1362 1432 1363
rect 1446 1363 1452 1364
rect 1446 1359 1447 1363
rect 1451 1359 1452 1363
rect 1414 1358 1420 1359
rect 1446 1358 1452 1359
rect 1414 1354 1415 1358
rect 1419 1354 1420 1358
rect 1414 1353 1420 1354
rect 1423 1355 1429 1356
rect 1423 1351 1424 1355
rect 1428 1351 1429 1355
rect 1423 1350 1429 1351
rect 1211 1348 1250 1350
rect 1408 1348 1427 1350
rect 1211 1347 1212 1348
rect 1206 1346 1212 1347
rect 1015 1343 1024 1344
rect 1167 1343 1176 1344
rect 1423 1343 1432 1344
rect 588 1340 626 1342
rect 630 1342 636 1343
rect 588 1339 589 1340
rect 583 1338 589 1339
rect 630 1338 631 1342
rect 635 1338 636 1342
rect 678 1342 684 1343
rect 574 1337 580 1338
rect 630 1337 636 1338
rect 639 1339 645 1340
rect 527 1334 533 1335
rect 639 1335 640 1339
rect 644 1335 645 1339
rect 678 1338 679 1342
rect 683 1338 684 1342
rect 726 1342 732 1343
rect 678 1337 684 1338
rect 687 1339 693 1340
rect 639 1334 645 1335
rect 687 1335 688 1339
rect 692 1338 693 1339
rect 726 1338 727 1342
rect 731 1338 732 1342
rect 766 1342 772 1343
rect 692 1336 714 1338
rect 726 1337 732 1338
rect 735 1339 741 1340
rect 692 1335 693 1336
rect 687 1334 693 1335
rect 110 1332 116 1333
rect 175 1331 181 1332
rect 175 1327 176 1331
rect 180 1330 181 1331
rect 200 1330 202 1334
rect 180 1328 202 1330
rect 180 1327 181 1328
rect 175 1326 181 1327
rect 240 1326 242 1334
rect 399 1331 405 1332
rect 220 1324 242 1326
rect 287 1327 293 1328
rect 199 1323 205 1324
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 199 1319 200 1323
rect 204 1322 205 1323
rect 220 1322 222 1324
rect 287 1323 288 1327
rect 292 1326 293 1327
rect 318 1327 324 1328
rect 318 1326 319 1327
rect 292 1324 319 1326
rect 292 1323 293 1324
rect 287 1322 293 1323
rect 318 1323 319 1324
rect 323 1323 324 1327
rect 318 1322 324 1323
rect 326 1327 332 1328
rect 326 1323 327 1327
rect 331 1326 332 1327
rect 343 1327 349 1328
rect 343 1326 344 1327
rect 331 1324 344 1326
rect 331 1323 332 1324
rect 326 1322 332 1323
rect 343 1323 344 1324
rect 348 1323 349 1327
rect 399 1327 400 1331
rect 404 1330 405 1331
rect 464 1330 466 1334
rect 404 1328 466 1330
rect 404 1327 405 1328
rect 399 1326 405 1327
rect 529 1326 531 1334
rect 583 1331 589 1332
rect 583 1327 584 1331
rect 588 1330 589 1331
rect 640 1330 642 1334
rect 588 1328 642 1330
rect 687 1331 696 1332
rect 588 1327 589 1328
rect 583 1326 589 1327
rect 687 1327 688 1331
rect 695 1327 696 1331
rect 712 1330 714 1336
rect 735 1335 736 1339
rect 740 1338 741 1339
rect 766 1338 767 1342
rect 771 1338 772 1342
rect 798 1342 804 1343
rect 740 1336 758 1338
rect 766 1337 772 1338
rect 775 1339 781 1340
rect 740 1335 741 1336
rect 735 1334 741 1335
rect 735 1331 741 1332
rect 735 1330 736 1331
rect 712 1328 736 1330
rect 687 1326 696 1327
rect 735 1327 736 1328
rect 740 1327 741 1331
rect 735 1326 741 1327
rect 756 1326 758 1336
rect 775 1335 776 1339
rect 780 1335 781 1339
rect 798 1338 799 1342
rect 803 1338 804 1342
rect 830 1342 836 1343
rect 798 1337 804 1338
rect 807 1339 813 1340
rect 775 1334 781 1335
rect 807 1335 808 1339
rect 812 1338 813 1339
rect 830 1338 831 1342
rect 835 1338 836 1342
rect 862 1342 868 1343
rect 812 1336 826 1338
rect 830 1337 836 1338
rect 839 1339 845 1340
rect 812 1335 813 1336
rect 807 1334 813 1335
rect 777 1330 779 1334
rect 807 1331 813 1332
rect 807 1330 808 1331
rect 777 1328 808 1330
rect 807 1327 808 1328
rect 812 1327 813 1331
rect 807 1326 813 1327
rect 824 1326 826 1336
rect 839 1335 840 1339
rect 844 1335 845 1339
rect 862 1338 863 1342
rect 867 1338 868 1342
rect 894 1342 900 1343
rect 862 1337 868 1338
rect 871 1339 877 1340
rect 839 1334 845 1335
rect 871 1335 872 1339
rect 876 1338 877 1339
rect 894 1338 895 1342
rect 899 1338 900 1342
rect 926 1342 932 1343
rect 876 1336 890 1338
rect 894 1337 900 1338
rect 903 1339 909 1340
rect 876 1335 877 1336
rect 871 1334 877 1335
rect 841 1330 843 1334
rect 871 1331 877 1332
rect 871 1330 872 1331
rect 841 1328 872 1330
rect 871 1327 872 1328
rect 876 1327 877 1331
rect 888 1330 890 1336
rect 903 1335 904 1339
rect 908 1338 909 1339
rect 926 1338 927 1342
rect 931 1338 932 1342
rect 966 1342 972 1343
rect 908 1336 922 1338
rect 926 1337 932 1338
rect 935 1339 941 1340
rect 908 1335 909 1336
rect 903 1334 909 1335
rect 903 1331 909 1332
rect 903 1330 904 1331
rect 888 1328 904 1330
rect 871 1326 877 1327
rect 903 1327 904 1328
rect 908 1327 909 1331
rect 920 1330 922 1336
rect 935 1335 936 1339
rect 940 1338 941 1339
rect 966 1338 967 1342
rect 971 1338 972 1342
rect 1006 1342 1012 1343
rect 940 1336 958 1338
rect 966 1337 972 1338
rect 975 1339 984 1340
rect 940 1335 941 1336
rect 935 1334 941 1335
rect 935 1331 941 1332
rect 935 1330 936 1331
rect 920 1328 936 1330
rect 903 1326 909 1327
rect 935 1327 936 1328
rect 940 1327 941 1331
rect 956 1330 958 1336
rect 975 1335 976 1339
rect 983 1335 984 1339
rect 1006 1338 1007 1342
rect 1011 1338 1012 1342
rect 1015 1339 1016 1343
rect 1023 1339 1024 1343
rect 1015 1338 1024 1339
rect 1054 1342 1060 1343
rect 1054 1338 1055 1342
rect 1059 1338 1060 1342
rect 1102 1342 1108 1343
rect 1006 1337 1012 1338
rect 1054 1337 1060 1338
rect 1063 1339 1069 1340
rect 975 1334 984 1335
rect 1063 1335 1064 1339
rect 1068 1335 1069 1339
rect 1102 1338 1103 1342
rect 1107 1338 1108 1342
rect 1158 1342 1164 1343
rect 1102 1337 1108 1338
rect 1111 1339 1117 1340
rect 1063 1334 1069 1335
rect 1111 1335 1112 1339
rect 1116 1338 1117 1339
rect 1122 1339 1128 1340
rect 1122 1338 1123 1339
rect 1116 1336 1123 1338
rect 1116 1335 1117 1336
rect 1111 1334 1117 1335
rect 1122 1335 1123 1336
rect 1127 1335 1128 1339
rect 1158 1338 1159 1342
rect 1163 1338 1164 1342
rect 1167 1339 1168 1343
rect 1175 1339 1176 1343
rect 1167 1338 1176 1339
rect 1214 1342 1220 1343
rect 1214 1338 1215 1342
rect 1219 1338 1220 1342
rect 1270 1342 1276 1343
rect 1158 1337 1164 1338
rect 1214 1337 1220 1338
rect 1223 1339 1229 1340
rect 1122 1334 1128 1335
rect 1223 1335 1224 1339
rect 1228 1335 1229 1339
rect 1270 1338 1271 1342
rect 1275 1338 1276 1342
rect 1326 1342 1332 1343
rect 1270 1337 1276 1338
rect 1279 1339 1285 1340
rect 1223 1334 1229 1335
rect 1279 1335 1280 1339
rect 1284 1338 1285 1339
rect 1314 1339 1320 1340
rect 1314 1338 1315 1339
rect 1284 1336 1315 1338
rect 1284 1335 1285 1336
rect 1279 1334 1285 1335
rect 1314 1335 1315 1336
rect 1319 1335 1320 1339
rect 1326 1338 1327 1342
rect 1331 1338 1332 1342
rect 1382 1342 1388 1343
rect 1326 1337 1332 1338
rect 1335 1339 1341 1340
rect 1314 1334 1320 1335
rect 1335 1335 1336 1339
rect 1340 1335 1341 1339
rect 1382 1338 1383 1342
rect 1387 1338 1388 1342
rect 1414 1342 1420 1343
rect 1382 1337 1388 1338
rect 1391 1339 1397 1340
rect 1335 1334 1341 1335
rect 1391 1335 1392 1339
rect 1396 1335 1397 1339
rect 1414 1338 1415 1342
rect 1419 1338 1420 1342
rect 1423 1339 1424 1343
rect 1431 1339 1432 1343
rect 1423 1338 1432 1339
rect 1414 1337 1420 1338
rect 1446 1337 1452 1338
rect 1391 1334 1397 1335
rect 975 1331 981 1332
rect 975 1330 976 1331
rect 956 1328 976 1330
rect 935 1326 941 1327
rect 975 1327 976 1328
rect 980 1327 981 1331
rect 975 1326 981 1327
rect 1015 1331 1021 1332
rect 1015 1327 1016 1331
rect 1020 1330 1021 1331
rect 1065 1330 1067 1334
rect 1020 1328 1067 1330
rect 1111 1331 1120 1332
rect 1020 1327 1021 1328
rect 1015 1326 1021 1327
rect 1111 1327 1112 1331
rect 1119 1327 1120 1331
rect 1111 1326 1120 1327
rect 1167 1331 1173 1332
rect 1167 1327 1168 1331
rect 1172 1330 1173 1331
rect 1224 1330 1226 1334
rect 1172 1328 1226 1330
rect 1279 1331 1285 1332
rect 1172 1327 1173 1328
rect 1167 1326 1173 1327
rect 1279 1327 1280 1331
rect 1284 1330 1285 1331
rect 1336 1330 1338 1334
rect 1284 1328 1338 1330
rect 1284 1327 1285 1328
rect 1279 1326 1285 1327
rect 1392 1326 1394 1334
rect 1446 1333 1447 1337
rect 1451 1333 1452 1337
rect 1446 1332 1452 1333
rect 496 1324 531 1326
rect 756 1324 779 1326
rect 824 1324 843 1326
rect 1344 1324 1394 1326
rect 343 1322 349 1323
rect 463 1323 469 1324
rect 204 1320 222 1322
rect 204 1319 205 1320
rect 199 1318 205 1319
rect 239 1319 245 1320
rect 110 1314 116 1315
rect 166 1316 172 1317
rect 166 1312 167 1316
rect 171 1312 172 1316
rect 166 1311 172 1312
rect 190 1316 196 1317
rect 190 1312 191 1316
rect 195 1312 196 1316
rect 190 1311 196 1312
rect 230 1316 236 1317
rect 230 1312 231 1316
rect 235 1312 236 1316
rect 239 1315 240 1319
rect 244 1318 245 1319
rect 247 1319 253 1320
rect 247 1318 248 1319
rect 244 1316 248 1318
rect 244 1315 245 1316
rect 239 1314 245 1315
rect 247 1315 248 1316
rect 252 1315 253 1319
rect 463 1319 464 1323
rect 468 1322 469 1323
rect 496 1322 498 1324
rect 468 1320 498 1322
rect 775 1323 781 1324
rect 468 1319 469 1320
rect 463 1318 469 1319
rect 775 1319 776 1323
rect 780 1319 781 1323
rect 775 1318 781 1319
rect 839 1323 845 1324
rect 839 1319 840 1323
rect 844 1319 845 1323
rect 839 1318 845 1319
rect 1335 1323 1341 1324
rect 1335 1319 1336 1323
rect 1340 1322 1341 1323
rect 1344 1322 1346 1324
rect 1340 1320 1346 1322
rect 1340 1319 1341 1320
rect 1335 1318 1341 1319
rect 1446 1319 1452 1320
rect 247 1314 253 1315
rect 278 1316 284 1317
rect 230 1311 236 1312
rect 278 1312 279 1316
rect 283 1312 284 1316
rect 278 1311 284 1312
rect 334 1316 340 1317
rect 334 1312 335 1316
rect 339 1312 340 1316
rect 334 1311 340 1312
rect 390 1316 396 1317
rect 390 1312 391 1316
rect 395 1312 396 1316
rect 390 1311 396 1312
rect 454 1316 460 1317
rect 454 1312 455 1316
rect 459 1312 460 1316
rect 518 1316 524 1317
rect 574 1316 580 1317
rect 518 1312 519 1316
rect 523 1312 524 1316
rect 454 1311 460 1312
rect 494 1311 500 1312
rect 518 1311 524 1312
rect 527 1315 533 1316
rect 527 1311 528 1315
rect 532 1311 533 1315
rect 574 1312 575 1316
rect 579 1312 580 1316
rect 574 1311 580 1312
rect 630 1316 636 1317
rect 678 1316 684 1317
rect 630 1312 631 1316
rect 635 1312 636 1316
rect 630 1311 636 1312
rect 639 1315 645 1316
rect 639 1311 640 1315
rect 644 1314 645 1315
rect 670 1315 676 1316
rect 670 1314 671 1315
rect 644 1312 671 1314
rect 644 1311 645 1312
rect 494 1307 495 1311
rect 499 1310 500 1311
rect 527 1310 533 1311
rect 639 1310 645 1311
rect 670 1311 671 1312
rect 675 1311 676 1315
rect 678 1312 679 1316
rect 683 1312 684 1316
rect 678 1311 684 1312
rect 726 1316 732 1317
rect 726 1312 727 1316
rect 731 1312 732 1316
rect 726 1311 732 1312
rect 766 1316 772 1317
rect 766 1312 767 1316
rect 771 1312 772 1316
rect 766 1311 772 1312
rect 798 1316 804 1317
rect 798 1312 799 1316
rect 803 1312 804 1316
rect 798 1311 804 1312
rect 830 1316 836 1317
rect 830 1312 831 1316
rect 835 1312 836 1316
rect 830 1311 836 1312
rect 862 1316 868 1317
rect 862 1312 863 1316
rect 867 1312 868 1316
rect 862 1311 868 1312
rect 894 1316 900 1317
rect 894 1312 895 1316
rect 899 1312 900 1316
rect 894 1311 900 1312
rect 926 1316 932 1317
rect 926 1312 927 1316
rect 931 1312 932 1316
rect 926 1311 932 1312
rect 966 1316 972 1317
rect 966 1312 967 1316
rect 971 1312 972 1316
rect 966 1311 972 1312
rect 1006 1316 1012 1317
rect 1006 1312 1007 1316
rect 1011 1312 1012 1316
rect 1006 1311 1012 1312
rect 1054 1316 1060 1317
rect 1102 1316 1108 1317
rect 1054 1312 1055 1316
rect 1059 1312 1060 1316
rect 1054 1311 1060 1312
rect 1063 1315 1069 1316
rect 1063 1311 1064 1315
rect 1068 1314 1069 1315
rect 1082 1315 1088 1316
rect 1082 1314 1083 1315
rect 1068 1312 1083 1314
rect 1068 1311 1069 1312
rect 670 1310 676 1311
rect 1063 1310 1069 1311
rect 1082 1311 1083 1312
rect 1087 1311 1088 1315
rect 1102 1312 1103 1316
rect 1107 1312 1108 1316
rect 1102 1311 1108 1312
rect 1158 1316 1164 1317
rect 1158 1312 1159 1316
rect 1163 1312 1164 1316
rect 1158 1311 1164 1312
rect 1214 1316 1220 1317
rect 1270 1316 1276 1317
rect 1214 1312 1215 1316
rect 1219 1312 1220 1316
rect 1214 1311 1220 1312
rect 1223 1315 1229 1316
rect 1223 1311 1224 1315
rect 1228 1314 1229 1315
rect 1258 1315 1264 1316
rect 1258 1314 1259 1315
rect 1228 1312 1259 1314
rect 1228 1311 1229 1312
rect 1082 1310 1088 1311
rect 1223 1310 1229 1311
rect 1258 1311 1259 1312
rect 1263 1311 1264 1315
rect 1270 1312 1271 1316
rect 1275 1312 1276 1316
rect 1270 1311 1276 1312
rect 1326 1316 1332 1317
rect 1326 1312 1327 1316
rect 1331 1312 1332 1316
rect 1382 1316 1388 1317
rect 1414 1316 1420 1317
rect 1382 1312 1383 1316
rect 1387 1312 1388 1316
rect 1326 1311 1332 1312
rect 1374 1311 1380 1312
rect 1382 1311 1388 1312
rect 1391 1315 1397 1316
rect 1391 1311 1392 1315
rect 1396 1311 1397 1315
rect 1414 1312 1415 1316
rect 1419 1312 1420 1316
rect 1414 1311 1420 1312
rect 1423 1315 1432 1316
rect 1423 1311 1424 1315
rect 1431 1311 1432 1315
rect 1446 1315 1447 1319
rect 1451 1315 1452 1319
rect 1446 1314 1452 1315
rect 1258 1310 1264 1311
rect 499 1308 514 1310
rect 499 1307 500 1308
rect 494 1306 500 1307
rect 512 1306 514 1308
rect 529 1306 531 1310
rect 1374 1307 1375 1311
rect 1379 1307 1380 1311
rect 1391 1310 1397 1311
rect 1423 1310 1432 1311
rect 1374 1306 1380 1307
rect 1392 1306 1394 1310
rect 230 1304 236 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 230 1300 231 1304
rect 235 1300 236 1304
rect 230 1299 236 1300
rect 254 1304 260 1305
rect 254 1300 255 1304
rect 259 1300 260 1304
rect 254 1299 260 1300
rect 278 1304 284 1305
rect 278 1300 279 1304
rect 283 1300 284 1304
rect 278 1299 284 1300
rect 302 1304 308 1305
rect 302 1300 303 1304
rect 307 1300 308 1304
rect 302 1299 308 1300
rect 326 1304 332 1305
rect 326 1300 327 1304
rect 331 1300 332 1304
rect 326 1299 332 1300
rect 350 1304 356 1305
rect 350 1300 351 1304
rect 355 1300 356 1304
rect 350 1299 356 1300
rect 374 1304 380 1305
rect 374 1300 375 1304
rect 379 1300 380 1304
rect 374 1299 380 1300
rect 398 1304 404 1305
rect 398 1300 399 1304
rect 403 1300 404 1304
rect 398 1299 404 1300
rect 422 1304 428 1305
rect 422 1300 423 1304
rect 427 1300 428 1304
rect 422 1299 428 1300
rect 446 1304 452 1305
rect 446 1300 447 1304
rect 451 1300 452 1304
rect 446 1299 452 1300
rect 470 1304 476 1305
rect 470 1300 471 1304
rect 475 1300 476 1304
rect 470 1299 476 1300
rect 502 1304 508 1305
rect 512 1304 531 1306
rect 542 1304 548 1305
rect 502 1300 503 1304
rect 507 1300 508 1304
rect 502 1299 508 1300
rect 542 1300 543 1304
rect 547 1300 548 1304
rect 542 1299 548 1300
rect 590 1304 596 1305
rect 590 1300 591 1304
rect 595 1300 596 1304
rect 590 1299 596 1300
rect 646 1304 652 1305
rect 646 1300 647 1304
rect 651 1300 652 1304
rect 646 1299 652 1300
rect 694 1304 700 1305
rect 694 1300 695 1304
rect 699 1300 700 1304
rect 694 1299 700 1300
rect 742 1304 748 1305
rect 742 1300 743 1304
rect 747 1300 748 1304
rect 742 1299 748 1300
rect 790 1304 796 1305
rect 790 1300 791 1304
rect 795 1300 796 1304
rect 790 1299 796 1300
rect 838 1304 844 1305
rect 838 1300 839 1304
rect 843 1300 844 1304
rect 838 1299 844 1300
rect 878 1304 884 1305
rect 878 1300 879 1304
rect 883 1300 884 1304
rect 878 1299 884 1300
rect 910 1304 916 1305
rect 910 1300 911 1304
rect 915 1300 916 1304
rect 910 1299 916 1300
rect 950 1304 956 1305
rect 950 1300 951 1304
rect 955 1300 956 1304
rect 950 1299 956 1300
rect 990 1304 996 1305
rect 990 1300 991 1304
rect 995 1300 996 1304
rect 990 1299 996 1300
rect 1030 1304 1036 1305
rect 1030 1300 1031 1304
rect 1035 1300 1036 1304
rect 1030 1299 1036 1300
rect 1070 1304 1076 1305
rect 1070 1300 1071 1304
rect 1075 1300 1076 1304
rect 1070 1299 1076 1300
rect 1110 1304 1116 1305
rect 1150 1304 1156 1305
rect 1110 1300 1111 1304
rect 1115 1300 1116 1304
rect 1110 1299 1116 1300
rect 1119 1303 1128 1304
rect 1119 1299 1120 1303
rect 1127 1299 1128 1303
rect 1150 1300 1151 1304
rect 1155 1300 1156 1304
rect 1150 1299 1156 1300
rect 1198 1304 1204 1305
rect 1198 1300 1199 1304
rect 1203 1300 1204 1304
rect 1198 1299 1204 1300
rect 1246 1304 1252 1305
rect 1246 1300 1247 1304
rect 1251 1300 1252 1304
rect 1246 1299 1252 1300
rect 1302 1304 1308 1305
rect 1366 1304 1372 1305
rect 1376 1304 1394 1306
rect 1414 1304 1420 1305
rect 1302 1300 1303 1304
rect 1307 1300 1308 1304
rect 1302 1299 1308 1300
rect 1311 1303 1320 1304
rect 1311 1299 1312 1303
rect 1319 1299 1320 1303
rect 1366 1300 1367 1304
rect 1371 1300 1372 1304
rect 1366 1299 1372 1300
rect 1414 1300 1415 1304
rect 1419 1300 1420 1304
rect 1414 1299 1420 1300
rect 1446 1301 1452 1302
rect 1119 1298 1128 1299
rect 1311 1298 1320 1299
rect 110 1296 116 1297
rect 1446 1297 1447 1301
rect 1451 1297 1452 1301
rect 1446 1296 1452 1297
rect 239 1295 245 1296
rect 239 1291 240 1295
rect 244 1294 245 1295
rect 266 1295 272 1296
rect 266 1294 267 1295
rect 244 1292 267 1294
rect 244 1291 245 1292
rect 239 1290 245 1291
rect 266 1291 267 1292
rect 271 1291 272 1295
rect 266 1290 272 1291
rect 311 1295 317 1296
rect 311 1291 312 1295
rect 316 1294 317 1295
rect 338 1295 344 1296
rect 338 1294 339 1295
rect 316 1292 339 1294
rect 316 1291 317 1292
rect 311 1290 317 1291
rect 338 1291 339 1292
rect 343 1291 344 1295
rect 338 1290 344 1291
rect 383 1295 389 1296
rect 383 1291 384 1295
rect 388 1294 389 1295
rect 410 1295 416 1296
rect 410 1294 411 1295
rect 388 1292 411 1294
rect 388 1291 389 1292
rect 383 1290 389 1291
rect 410 1291 411 1292
rect 415 1291 416 1295
rect 410 1290 416 1291
rect 703 1295 709 1296
rect 703 1291 704 1295
rect 708 1294 709 1295
rect 754 1295 760 1296
rect 754 1294 755 1295
rect 708 1292 755 1294
rect 708 1291 709 1292
rect 703 1290 709 1291
rect 754 1291 755 1292
rect 759 1291 760 1295
rect 754 1290 760 1291
rect 799 1295 805 1296
rect 799 1291 800 1295
rect 804 1294 805 1295
rect 978 1295 984 1296
rect 978 1294 979 1295
rect 804 1292 979 1294
rect 804 1291 805 1292
rect 799 1290 805 1291
rect 978 1291 979 1292
rect 983 1291 984 1295
rect 978 1290 984 1291
rect 263 1287 269 1288
rect 110 1283 116 1284
rect 110 1279 111 1283
rect 115 1279 116 1283
rect 263 1283 264 1287
rect 268 1286 269 1287
rect 271 1287 277 1288
rect 271 1286 272 1287
rect 268 1284 272 1286
rect 268 1283 269 1284
rect 263 1282 269 1283
rect 271 1283 272 1284
rect 276 1283 277 1287
rect 271 1282 277 1283
rect 287 1287 293 1288
rect 287 1283 288 1287
rect 292 1286 293 1287
rect 318 1287 324 1288
rect 292 1284 314 1286
rect 292 1283 293 1284
rect 287 1282 293 1283
rect 312 1280 314 1284
rect 318 1283 319 1287
rect 323 1286 324 1287
rect 335 1287 341 1288
rect 335 1286 336 1287
rect 323 1284 336 1286
rect 323 1283 324 1284
rect 318 1282 324 1283
rect 335 1283 336 1284
rect 340 1283 341 1287
rect 335 1282 341 1283
rect 359 1287 365 1288
rect 359 1283 360 1287
rect 364 1286 365 1287
rect 407 1287 413 1288
rect 407 1286 408 1287
rect 364 1284 387 1286
rect 364 1283 365 1284
rect 359 1282 365 1283
rect 385 1280 387 1284
rect 392 1284 408 1286
rect 239 1279 248 1280
rect 263 1279 272 1280
rect 311 1279 317 1280
rect 335 1279 344 1280
rect 359 1279 368 1280
rect 383 1279 389 1280
rect 110 1278 116 1279
rect 230 1278 236 1279
rect 230 1274 231 1278
rect 235 1274 236 1278
rect 239 1275 240 1279
rect 247 1275 248 1279
rect 239 1274 248 1275
rect 254 1278 260 1279
rect 254 1274 255 1278
rect 259 1274 260 1278
rect 263 1275 264 1279
rect 271 1275 272 1279
rect 263 1274 272 1275
rect 278 1278 284 1279
rect 278 1274 279 1278
rect 283 1274 284 1278
rect 302 1278 308 1279
rect 230 1273 236 1274
rect 254 1273 260 1274
rect 278 1273 284 1274
rect 287 1275 293 1276
rect 287 1271 288 1275
rect 292 1271 293 1275
rect 302 1274 303 1278
rect 307 1274 308 1278
rect 311 1275 312 1279
rect 316 1275 317 1279
rect 311 1274 317 1275
rect 326 1278 332 1279
rect 326 1274 327 1278
rect 331 1274 332 1278
rect 335 1275 336 1279
rect 343 1275 344 1279
rect 335 1274 344 1275
rect 350 1278 356 1279
rect 350 1274 351 1278
rect 355 1274 356 1278
rect 359 1275 360 1279
rect 367 1275 368 1279
rect 359 1274 368 1275
rect 374 1278 380 1279
rect 374 1274 375 1278
rect 379 1274 380 1278
rect 383 1275 384 1279
rect 388 1275 389 1279
rect 383 1274 389 1275
rect 302 1273 308 1274
rect 326 1273 332 1274
rect 350 1273 356 1274
rect 374 1273 380 1274
rect 287 1270 293 1271
rect 342 1271 348 1272
rect 271 1267 277 1268
rect 271 1263 272 1267
rect 276 1266 277 1267
rect 288 1266 290 1270
rect 276 1264 290 1266
rect 318 1267 324 1268
rect 276 1263 277 1264
rect 318 1263 319 1267
rect 323 1264 324 1267
rect 342 1267 343 1271
rect 347 1270 348 1271
rect 392 1270 394 1284
rect 407 1283 408 1284
rect 412 1283 413 1287
rect 431 1287 437 1288
rect 431 1286 432 1287
rect 407 1282 413 1283
rect 416 1284 432 1286
rect 407 1279 413 1280
rect 398 1278 404 1279
rect 398 1274 399 1278
rect 403 1274 404 1278
rect 407 1275 408 1279
rect 412 1278 413 1279
rect 416 1278 418 1284
rect 431 1283 432 1284
rect 436 1283 437 1287
rect 455 1287 461 1288
rect 455 1286 456 1287
rect 431 1282 437 1283
rect 440 1284 456 1286
rect 431 1279 437 1280
rect 412 1276 418 1278
rect 422 1278 428 1279
rect 412 1275 413 1276
rect 407 1274 413 1275
rect 422 1274 423 1278
rect 427 1274 428 1278
rect 431 1275 432 1279
rect 436 1278 437 1279
rect 440 1278 442 1284
rect 455 1283 456 1284
rect 460 1283 461 1287
rect 479 1287 485 1288
rect 479 1286 480 1287
rect 455 1282 461 1283
rect 464 1284 480 1286
rect 455 1279 461 1280
rect 436 1276 442 1278
rect 446 1278 452 1279
rect 436 1275 437 1276
rect 431 1274 437 1275
rect 446 1274 447 1278
rect 451 1274 452 1278
rect 455 1275 456 1279
rect 460 1278 461 1279
rect 464 1278 466 1284
rect 479 1283 480 1284
rect 484 1283 485 1287
rect 511 1287 517 1288
rect 511 1286 512 1287
rect 479 1282 485 1283
rect 496 1284 512 1286
rect 479 1279 485 1280
rect 460 1276 466 1278
rect 470 1278 476 1279
rect 460 1275 461 1276
rect 455 1274 461 1275
rect 470 1274 471 1278
rect 475 1274 476 1278
rect 479 1275 480 1279
rect 484 1278 485 1279
rect 496 1278 498 1284
rect 511 1283 512 1284
rect 516 1283 517 1287
rect 551 1287 557 1288
rect 551 1286 552 1287
rect 511 1282 517 1283
rect 532 1284 552 1286
rect 511 1279 517 1280
rect 484 1276 498 1278
rect 502 1278 508 1279
rect 484 1275 485 1276
rect 479 1274 485 1275
rect 502 1274 503 1278
rect 507 1274 508 1278
rect 511 1275 512 1279
rect 516 1278 517 1279
rect 532 1278 534 1284
rect 551 1283 552 1284
rect 556 1283 557 1287
rect 599 1287 605 1288
rect 599 1286 600 1287
rect 551 1282 557 1283
rect 576 1284 600 1286
rect 551 1279 557 1280
rect 516 1276 534 1278
rect 542 1278 548 1279
rect 516 1275 517 1276
rect 511 1274 517 1275
rect 542 1274 543 1278
rect 547 1274 548 1278
rect 551 1275 552 1279
rect 556 1278 557 1279
rect 576 1278 578 1284
rect 599 1283 600 1284
rect 604 1283 605 1287
rect 655 1287 661 1288
rect 655 1286 656 1287
rect 599 1282 605 1283
rect 628 1284 656 1286
rect 599 1279 605 1280
rect 556 1276 578 1278
rect 590 1278 596 1279
rect 556 1275 557 1276
rect 551 1274 557 1275
rect 590 1274 591 1278
rect 595 1274 596 1278
rect 599 1275 600 1279
rect 604 1278 605 1279
rect 628 1278 630 1284
rect 655 1283 656 1284
rect 660 1283 661 1287
rect 655 1282 661 1283
rect 670 1287 676 1288
rect 670 1283 671 1287
rect 675 1286 676 1287
rect 751 1287 757 1288
rect 675 1284 706 1286
rect 675 1283 676 1284
rect 670 1282 676 1283
rect 704 1280 706 1284
rect 751 1283 752 1287
rect 756 1286 757 1287
rect 847 1287 853 1288
rect 847 1286 848 1287
rect 756 1284 786 1286
rect 756 1283 757 1284
rect 751 1282 757 1283
rect 703 1279 709 1280
rect 751 1279 760 1280
rect 604 1276 630 1278
rect 646 1278 652 1279
rect 604 1275 605 1276
rect 599 1274 605 1275
rect 646 1274 647 1278
rect 651 1274 652 1278
rect 694 1278 700 1279
rect 398 1273 404 1274
rect 422 1273 428 1274
rect 446 1273 452 1274
rect 470 1273 476 1274
rect 502 1273 508 1274
rect 542 1273 548 1274
rect 590 1273 596 1274
rect 646 1273 652 1274
rect 655 1275 661 1276
rect 530 1271 536 1272
rect 347 1268 370 1270
rect 392 1268 490 1270
rect 347 1267 348 1268
rect 342 1266 348 1267
rect 368 1264 370 1268
rect 488 1264 490 1268
rect 530 1267 531 1271
rect 535 1270 536 1271
rect 655 1271 656 1275
rect 660 1271 661 1275
rect 694 1274 695 1278
rect 699 1274 700 1278
rect 703 1275 704 1279
rect 708 1275 709 1279
rect 703 1274 709 1275
rect 742 1278 748 1279
rect 742 1274 743 1278
rect 747 1274 748 1278
rect 751 1275 752 1279
rect 759 1275 760 1279
rect 751 1274 760 1275
rect 694 1273 700 1274
rect 742 1273 748 1274
rect 655 1270 661 1271
rect 784 1270 786 1284
rect 824 1284 848 1286
rect 799 1279 805 1280
rect 790 1278 796 1279
rect 790 1274 791 1278
rect 795 1274 796 1278
rect 799 1275 800 1279
rect 804 1278 805 1279
rect 824 1278 826 1284
rect 847 1283 848 1284
rect 852 1283 853 1287
rect 887 1287 893 1288
rect 887 1286 888 1287
rect 847 1282 853 1283
rect 868 1284 888 1286
rect 847 1279 853 1280
rect 804 1276 826 1278
rect 838 1278 844 1279
rect 804 1275 805 1276
rect 799 1274 805 1275
rect 838 1274 839 1278
rect 843 1274 844 1278
rect 847 1275 848 1279
rect 852 1278 853 1279
rect 868 1278 870 1284
rect 887 1283 888 1284
rect 892 1283 893 1287
rect 919 1287 925 1288
rect 919 1286 920 1287
rect 887 1282 893 1283
rect 904 1284 920 1286
rect 887 1279 893 1280
rect 852 1276 870 1278
rect 878 1278 884 1279
rect 852 1275 853 1276
rect 847 1274 853 1275
rect 878 1274 879 1278
rect 883 1274 884 1278
rect 887 1275 888 1279
rect 892 1278 893 1279
rect 904 1278 906 1284
rect 919 1283 920 1284
rect 924 1283 925 1287
rect 959 1287 965 1288
rect 959 1286 960 1287
rect 919 1282 925 1283
rect 940 1284 960 1286
rect 919 1279 925 1280
rect 892 1276 906 1278
rect 910 1278 916 1279
rect 892 1275 893 1276
rect 887 1274 893 1275
rect 910 1274 911 1278
rect 915 1274 916 1278
rect 919 1275 920 1279
rect 924 1278 925 1279
rect 940 1278 942 1284
rect 959 1283 960 1284
rect 964 1283 965 1287
rect 999 1287 1005 1288
rect 999 1286 1000 1287
rect 959 1282 965 1283
rect 980 1284 1000 1286
rect 959 1279 965 1280
rect 924 1276 942 1278
rect 950 1278 956 1279
rect 924 1275 925 1276
rect 919 1274 925 1275
rect 950 1274 951 1278
rect 955 1274 956 1278
rect 959 1275 960 1279
rect 964 1278 965 1279
rect 980 1278 982 1284
rect 999 1283 1000 1284
rect 1004 1283 1005 1287
rect 1039 1287 1045 1288
rect 1039 1286 1040 1287
rect 999 1282 1005 1283
rect 1020 1284 1040 1286
rect 999 1279 1005 1280
rect 964 1276 982 1278
rect 990 1278 996 1279
rect 964 1275 965 1276
rect 959 1274 965 1275
rect 990 1274 991 1278
rect 995 1274 996 1278
rect 999 1275 1000 1279
rect 1004 1278 1005 1279
rect 1020 1278 1022 1284
rect 1039 1283 1040 1284
rect 1044 1283 1045 1287
rect 1079 1287 1085 1288
rect 1079 1286 1080 1287
rect 1039 1282 1045 1283
rect 1060 1284 1080 1286
rect 1039 1279 1045 1280
rect 1004 1276 1022 1278
rect 1030 1278 1036 1279
rect 1004 1275 1005 1276
rect 999 1274 1005 1275
rect 1030 1274 1031 1278
rect 1035 1274 1036 1278
rect 1039 1275 1040 1279
rect 1044 1278 1045 1279
rect 1060 1278 1062 1284
rect 1079 1283 1080 1284
rect 1084 1283 1085 1287
rect 1079 1282 1085 1283
rect 1138 1287 1144 1288
rect 1138 1283 1139 1287
rect 1143 1286 1144 1287
rect 1159 1287 1165 1288
rect 1159 1286 1160 1287
rect 1143 1284 1160 1286
rect 1143 1283 1144 1284
rect 1138 1282 1144 1283
rect 1159 1283 1160 1284
rect 1164 1283 1165 1287
rect 1207 1287 1213 1288
rect 1207 1286 1208 1287
rect 1159 1282 1165 1283
rect 1184 1284 1208 1286
rect 1079 1279 1088 1280
rect 1119 1279 1125 1280
rect 1159 1279 1165 1280
rect 1044 1276 1062 1278
rect 1070 1278 1076 1279
rect 1044 1275 1045 1276
rect 1039 1274 1045 1275
rect 1070 1274 1071 1278
rect 1075 1274 1076 1278
rect 1079 1275 1080 1279
rect 1087 1275 1088 1279
rect 1079 1274 1088 1275
rect 1110 1278 1116 1279
rect 1110 1274 1111 1278
rect 1115 1274 1116 1278
rect 1119 1275 1120 1279
rect 1124 1275 1125 1279
rect 1119 1274 1125 1275
rect 1150 1278 1156 1279
rect 1150 1274 1151 1278
rect 1155 1274 1156 1278
rect 1159 1275 1160 1279
rect 1164 1278 1165 1279
rect 1184 1278 1186 1284
rect 1207 1283 1208 1284
rect 1212 1283 1213 1287
rect 1255 1287 1261 1288
rect 1255 1286 1256 1287
rect 1207 1282 1213 1283
rect 1232 1284 1256 1286
rect 1207 1279 1213 1280
rect 1164 1276 1186 1278
rect 1198 1278 1204 1279
rect 1164 1275 1165 1276
rect 1159 1274 1165 1275
rect 1198 1274 1199 1278
rect 1203 1274 1204 1278
rect 1207 1275 1208 1279
rect 1212 1278 1213 1279
rect 1232 1278 1234 1284
rect 1255 1283 1256 1284
rect 1260 1283 1261 1287
rect 1375 1287 1381 1288
rect 1375 1286 1376 1287
rect 1255 1282 1261 1283
rect 1344 1284 1376 1286
rect 1255 1279 1264 1280
rect 1311 1279 1317 1280
rect 1212 1276 1234 1278
rect 1246 1278 1252 1279
rect 1212 1275 1213 1276
rect 1207 1274 1213 1275
rect 1246 1274 1247 1278
rect 1251 1274 1252 1278
rect 1255 1275 1256 1279
rect 1263 1275 1264 1279
rect 1255 1274 1264 1275
rect 1302 1278 1308 1279
rect 1302 1274 1303 1278
rect 1307 1274 1308 1278
rect 1311 1275 1312 1279
rect 1316 1278 1317 1279
rect 1344 1278 1346 1284
rect 1375 1283 1376 1284
rect 1380 1283 1381 1287
rect 1375 1282 1381 1283
rect 1386 1287 1392 1288
rect 1386 1283 1387 1287
rect 1391 1286 1392 1287
rect 1423 1287 1429 1288
rect 1423 1286 1424 1287
rect 1391 1284 1424 1286
rect 1391 1283 1392 1284
rect 1386 1282 1392 1283
rect 1423 1283 1424 1284
rect 1428 1283 1429 1287
rect 1423 1282 1429 1283
rect 1446 1283 1452 1284
rect 1423 1279 1432 1280
rect 1316 1276 1346 1278
rect 1366 1278 1372 1279
rect 1316 1275 1317 1276
rect 1311 1274 1317 1275
rect 1366 1274 1367 1278
rect 1371 1274 1372 1278
rect 1414 1278 1420 1279
rect 790 1273 796 1274
rect 838 1273 844 1274
rect 878 1273 884 1274
rect 910 1273 916 1274
rect 950 1273 956 1274
rect 990 1273 996 1274
rect 1030 1273 1036 1274
rect 1070 1273 1076 1274
rect 1110 1273 1116 1274
rect 1002 1271 1008 1272
rect 535 1268 659 1270
rect 784 1268 922 1270
rect 535 1267 536 1268
rect 530 1266 536 1267
rect 920 1264 922 1268
rect 1002 1267 1003 1271
rect 1007 1270 1008 1271
rect 1120 1270 1122 1274
rect 1150 1273 1156 1274
rect 1198 1273 1204 1274
rect 1246 1273 1252 1274
rect 1302 1273 1308 1274
rect 1366 1273 1372 1274
rect 1375 1275 1381 1276
rect 1007 1268 1122 1270
rect 1127 1271 1133 1272
rect 1007 1267 1008 1268
rect 1002 1266 1008 1267
rect 1127 1267 1128 1271
rect 1132 1270 1133 1271
rect 1294 1271 1300 1272
rect 1294 1270 1295 1271
rect 1132 1268 1295 1270
rect 1132 1267 1133 1268
rect 1127 1266 1133 1267
rect 1294 1267 1295 1268
rect 1299 1267 1300 1271
rect 1294 1266 1300 1267
rect 1322 1271 1328 1272
rect 1322 1267 1323 1271
rect 1327 1270 1328 1271
rect 1375 1271 1376 1275
rect 1380 1271 1381 1275
rect 1414 1274 1415 1278
rect 1419 1274 1420 1278
rect 1423 1275 1424 1279
rect 1431 1275 1432 1279
rect 1446 1279 1447 1283
rect 1451 1279 1452 1283
rect 1446 1278 1452 1279
rect 1423 1274 1432 1275
rect 1414 1273 1420 1274
rect 1375 1270 1381 1271
rect 1327 1268 1378 1270
rect 1327 1267 1328 1268
rect 1322 1266 1328 1267
rect 323 1263 325 1264
rect 367 1263 373 1264
rect 487 1263 493 1264
rect 919 1263 925 1264
rect 1071 1263 1077 1264
rect 271 1262 277 1263
rect 310 1262 316 1263
rect 318 1262 320 1263
rect 310 1258 311 1262
rect 315 1258 316 1262
rect 319 1259 320 1262
rect 324 1259 325 1263
rect 319 1258 325 1259
rect 334 1262 340 1263
rect 334 1258 335 1262
rect 339 1258 340 1262
rect 358 1262 364 1263
rect 110 1257 116 1258
rect 310 1257 316 1258
rect 334 1257 340 1258
rect 343 1259 349 1260
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 343 1255 344 1259
rect 348 1255 349 1259
rect 358 1258 359 1262
rect 363 1258 364 1262
rect 367 1259 368 1263
rect 372 1259 373 1263
rect 367 1258 373 1259
rect 382 1262 388 1263
rect 382 1258 383 1262
rect 387 1258 388 1262
rect 414 1262 420 1263
rect 358 1257 364 1258
rect 382 1257 388 1258
rect 391 1259 397 1260
rect 343 1254 349 1255
rect 391 1255 392 1259
rect 396 1258 397 1259
rect 414 1258 415 1262
rect 419 1258 420 1262
rect 446 1262 452 1263
rect 396 1256 410 1258
rect 414 1257 420 1258
rect 423 1259 429 1260
rect 396 1255 397 1256
rect 391 1254 397 1255
rect 110 1252 116 1253
rect 319 1251 325 1252
rect 319 1247 320 1251
rect 324 1250 325 1251
rect 345 1250 347 1254
rect 324 1248 347 1250
rect 366 1251 373 1252
rect 324 1247 325 1248
rect 319 1246 325 1247
rect 366 1247 367 1251
rect 372 1247 373 1251
rect 366 1246 373 1247
rect 408 1246 410 1256
rect 423 1255 424 1259
rect 428 1255 429 1259
rect 446 1258 447 1262
rect 451 1258 452 1262
rect 478 1262 484 1263
rect 446 1257 452 1258
rect 455 1259 461 1260
rect 423 1254 429 1255
rect 455 1255 456 1259
rect 460 1258 461 1259
rect 478 1258 479 1262
rect 483 1258 484 1262
rect 487 1259 488 1263
rect 492 1259 493 1263
rect 487 1258 493 1259
rect 518 1262 524 1263
rect 518 1258 519 1262
rect 523 1258 524 1262
rect 558 1262 564 1263
rect 460 1256 474 1258
rect 478 1257 484 1258
rect 518 1257 524 1258
rect 527 1259 533 1260
rect 460 1255 461 1256
rect 455 1254 461 1255
rect 425 1250 427 1254
rect 455 1251 461 1252
rect 455 1250 456 1251
rect 425 1248 456 1250
rect 455 1247 456 1248
rect 460 1247 461 1251
rect 472 1250 474 1256
rect 527 1255 528 1259
rect 532 1255 533 1259
rect 558 1258 559 1262
rect 563 1258 564 1262
rect 614 1262 620 1263
rect 558 1257 564 1258
rect 567 1259 573 1260
rect 527 1254 533 1255
rect 567 1255 568 1259
rect 572 1258 573 1259
rect 614 1258 615 1262
rect 619 1258 620 1262
rect 678 1262 684 1263
rect 572 1256 598 1258
rect 614 1257 620 1258
rect 623 1259 629 1260
rect 572 1255 573 1256
rect 567 1254 573 1255
rect 487 1251 493 1252
rect 487 1250 488 1251
rect 472 1248 488 1250
rect 455 1246 461 1247
rect 487 1247 488 1248
rect 492 1247 493 1251
rect 529 1250 531 1254
rect 567 1251 573 1252
rect 567 1250 568 1251
rect 529 1248 568 1250
rect 487 1246 493 1247
rect 567 1247 568 1248
rect 572 1247 573 1251
rect 596 1250 598 1256
rect 623 1255 624 1259
rect 628 1258 629 1259
rect 678 1258 679 1262
rect 683 1258 684 1262
rect 750 1262 756 1263
rect 628 1256 662 1258
rect 678 1257 684 1258
rect 687 1259 696 1260
rect 628 1255 629 1256
rect 623 1254 629 1255
rect 623 1251 629 1252
rect 623 1250 624 1251
rect 596 1248 624 1250
rect 567 1246 573 1247
rect 623 1247 624 1248
rect 628 1247 629 1251
rect 660 1250 662 1256
rect 687 1255 688 1259
rect 695 1255 696 1259
rect 750 1258 751 1262
rect 755 1258 756 1262
rect 830 1262 836 1263
rect 750 1257 756 1258
rect 759 1259 765 1260
rect 687 1254 696 1255
rect 759 1255 760 1259
rect 764 1258 765 1259
rect 830 1258 831 1262
rect 835 1258 836 1262
rect 910 1262 916 1263
rect 764 1256 802 1258
rect 830 1257 836 1258
rect 839 1259 845 1260
rect 764 1255 765 1256
rect 759 1254 765 1255
rect 687 1251 693 1252
rect 687 1250 688 1251
rect 660 1248 688 1250
rect 623 1246 629 1247
rect 687 1247 688 1248
rect 692 1247 693 1251
rect 687 1246 693 1247
rect 800 1246 802 1256
rect 839 1255 840 1259
rect 844 1255 845 1259
rect 910 1258 911 1262
rect 915 1258 916 1262
rect 919 1259 920 1263
rect 924 1259 925 1263
rect 919 1258 925 1259
rect 990 1262 996 1263
rect 990 1258 991 1262
rect 995 1258 996 1262
rect 1062 1262 1068 1263
rect 910 1257 916 1258
rect 990 1257 996 1258
rect 999 1259 1005 1260
rect 839 1254 845 1255
rect 999 1255 1000 1259
rect 1004 1258 1005 1259
rect 1062 1258 1063 1262
rect 1067 1258 1068 1262
rect 1071 1259 1072 1263
rect 1076 1262 1077 1263
rect 1111 1263 1117 1264
rect 1135 1263 1144 1264
rect 1383 1263 1392 1264
rect 1111 1262 1112 1263
rect 1076 1260 1112 1262
rect 1076 1259 1077 1260
rect 1071 1258 1077 1259
rect 1111 1259 1112 1260
rect 1116 1259 1117 1263
rect 1111 1258 1117 1259
rect 1126 1262 1132 1263
rect 1126 1258 1127 1262
rect 1131 1258 1132 1262
rect 1135 1259 1136 1263
rect 1143 1259 1144 1263
rect 1135 1258 1144 1259
rect 1190 1262 1196 1263
rect 1190 1258 1191 1262
rect 1195 1258 1196 1262
rect 1246 1262 1252 1263
rect 1004 1256 1038 1258
rect 1062 1257 1068 1258
rect 1126 1257 1132 1258
rect 1190 1257 1196 1258
rect 1199 1259 1205 1260
rect 1004 1255 1005 1256
rect 999 1254 1005 1255
rect 841 1250 843 1254
rect 919 1251 925 1252
rect 919 1250 920 1251
rect 841 1248 920 1250
rect 919 1247 920 1248
rect 924 1247 925 1251
rect 919 1246 925 1247
rect 999 1251 1008 1252
rect 999 1247 1000 1251
rect 1007 1247 1008 1251
rect 1036 1250 1038 1256
rect 1199 1255 1200 1259
rect 1204 1255 1205 1259
rect 1246 1258 1247 1262
rect 1251 1258 1252 1262
rect 1310 1262 1316 1263
rect 1246 1257 1252 1258
rect 1255 1259 1261 1260
rect 1199 1254 1205 1255
rect 1255 1255 1256 1259
rect 1260 1255 1261 1259
rect 1310 1258 1311 1262
rect 1315 1258 1316 1262
rect 1374 1262 1380 1263
rect 1310 1257 1316 1258
rect 1319 1259 1325 1260
rect 1255 1254 1261 1255
rect 1319 1255 1320 1259
rect 1324 1258 1325 1259
rect 1327 1259 1333 1260
rect 1327 1258 1328 1259
rect 1324 1256 1328 1258
rect 1324 1255 1325 1256
rect 1319 1254 1325 1255
rect 1327 1255 1328 1256
rect 1332 1255 1333 1259
rect 1374 1258 1375 1262
rect 1379 1258 1380 1262
rect 1383 1259 1384 1263
rect 1391 1259 1392 1263
rect 1383 1258 1392 1259
rect 1414 1262 1420 1263
rect 1414 1258 1415 1262
rect 1419 1258 1420 1262
rect 1374 1257 1380 1258
rect 1414 1257 1420 1258
rect 1423 1259 1429 1260
rect 1327 1254 1333 1255
rect 1423 1255 1424 1259
rect 1428 1255 1429 1259
rect 1423 1254 1429 1255
rect 1446 1257 1452 1258
rect 1071 1251 1077 1252
rect 1071 1250 1072 1251
rect 1036 1248 1072 1250
rect 999 1246 1008 1247
rect 1071 1247 1072 1248
rect 1076 1247 1077 1251
rect 1071 1246 1077 1247
rect 1135 1251 1141 1252
rect 1135 1247 1136 1251
rect 1140 1250 1141 1251
rect 1201 1250 1203 1254
rect 1140 1248 1203 1250
rect 1140 1247 1141 1248
rect 1135 1246 1141 1247
rect 1256 1246 1258 1254
rect 1319 1251 1328 1252
rect 1319 1247 1320 1251
rect 1327 1247 1328 1251
rect 1319 1246 1328 1247
rect 1383 1251 1389 1252
rect 1383 1247 1384 1251
rect 1388 1250 1389 1251
rect 1425 1250 1427 1254
rect 1446 1253 1447 1257
rect 1451 1253 1452 1257
rect 1446 1252 1452 1253
rect 1388 1248 1427 1250
rect 1388 1247 1389 1248
rect 1383 1246 1389 1247
rect 408 1244 427 1246
rect 800 1244 843 1246
rect 1201 1244 1258 1246
rect 343 1243 352 1244
rect 110 1239 116 1240
rect 110 1235 111 1239
rect 115 1235 116 1239
rect 343 1239 344 1243
rect 351 1239 352 1243
rect 343 1238 352 1239
rect 423 1243 429 1244
rect 423 1239 424 1243
rect 428 1239 429 1243
rect 423 1238 429 1239
rect 527 1243 536 1244
rect 527 1239 528 1243
rect 535 1239 536 1243
rect 527 1238 536 1239
rect 839 1243 845 1244
rect 839 1239 840 1243
rect 844 1239 845 1243
rect 839 1238 845 1239
rect 1199 1243 1205 1244
rect 1199 1239 1200 1243
rect 1204 1239 1205 1243
rect 1199 1238 1205 1239
rect 1446 1239 1452 1240
rect 110 1234 116 1235
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 334 1236 340 1237
rect 334 1232 335 1236
rect 339 1232 340 1236
rect 334 1231 340 1232
rect 358 1236 364 1237
rect 358 1232 359 1236
rect 363 1232 364 1236
rect 358 1231 364 1232
rect 382 1236 388 1237
rect 414 1236 420 1237
rect 382 1232 383 1236
rect 387 1232 388 1236
rect 382 1231 388 1232
rect 391 1235 397 1236
rect 391 1231 392 1235
rect 396 1234 397 1235
rect 399 1235 405 1236
rect 399 1234 400 1235
rect 396 1232 400 1234
rect 396 1231 397 1232
rect 391 1230 397 1231
rect 399 1231 400 1232
rect 404 1231 405 1235
rect 414 1232 415 1236
rect 419 1232 420 1236
rect 414 1231 420 1232
rect 446 1236 452 1237
rect 446 1232 447 1236
rect 451 1232 452 1236
rect 446 1231 452 1232
rect 478 1236 484 1237
rect 478 1232 479 1236
rect 483 1232 484 1236
rect 478 1231 484 1232
rect 518 1236 524 1237
rect 518 1232 519 1236
rect 523 1232 524 1236
rect 518 1231 524 1232
rect 558 1236 564 1237
rect 558 1232 559 1236
rect 563 1232 564 1236
rect 558 1231 564 1232
rect 614 1236 620 1237
rect 614 1232 615 1236
rect 619 1232 620 1236
rect 614 1231 620 1232
rect 678 1236 684 1237
rect 678 1232 679 1236
rect 683 1232 684 1236
rect 678 1231 684 1232
rect 750 1236 756 1237
rect 830 1236 836 1237
rect 750 1232 751 1236
rect 755 1232 756 1236
rect 750 1231 756 1232
rect 759 1235 768 1236
rect 759 1231 760 1235
rect 767 1231 768 1235
rect 830 1232 831 1236
rect 835 1232 836 1236
rect 830 1231 836 1232
rect 910 1236 916 1237
rect 910 1232 911 1236
rect 915 1232 916 1236
rect 910 1231 916 1232
rect 990 1236 996 1237
rect 990 1232 991 1236
rect 995 1232 996 1236
rect 990 1231 996 1232
rect 1062 1236 1068 1237
rect 1062 1232 1063 1236
rect 1067 1232 1068 1236
rect 1062 1231 1068 1232
rect 1126 1236 1132 1237
rect 1126 1232 1127 1236
rect 1131 1232 1132 1236
rect 1126 1231 1132 1232
rect 1190 1236 1196 1237
rect 1190 1232 1191 1236
rect 1195 1232 1196 1236
rect 1190 1231 1196 1232
rect 1246 1236 1252 1237
rect 1310 1236 1316 1237
rect 1246 1232 1247 1236
rect 1251 1232 1252 1236
rect 1246 1231 1252 1232
rect 1255 1235 1261 1236
rect 1255 1231 1256 1235
rect 1260 1234 1261 1235
rect 1260 1232 1290 1234
rect 1260 1231 1261 1232
rect 399 1230 405 1231
rect 759 1230 768 1231
rect 1255 1230 1261 1231
rect 1288 1226 1290 1232
rect 1310 1232 1311 1236
rect 1315 1232 1316 1236
rect 1310 1231 1316 1232
rect 1374 1236 1380 1237
rect 1374 1232 1375 1236
rect 1379 1232 1380 1236
rect 1374 1231 1380 1232
rect 1414 1236 1420 1237
rect 1414 1232 1415 1236
rect 1419 1232 1420 1236
rect 1414 1231 1420 1232
rect 1423 1235 1432 1236
rect 1423 1231 1424 1235
rect 1431 1231 1432 1235
rect 1446 1235 1447 1239
rect 1451 1235 1452 1239
rect 1446 1234 1452 1235
rect 1423 1230 1432 1231
rect 1327 1227 1333 1228
rect 1327 1226 1328 1227
rect 326 1224 332 1225
rect 110 1221 116 1222
rect 110 1217 111 1221
rect 115 1217 116 1221
rect 326 1220 327 1224
rect 331 1220 332 1224
rect 326 1219 332 1220
rect 366 1224 372 1225
rect 366 1220 367 1224
rect 371 1220 372 1224
rect 366 1219 372 1220
rect 406 1224 412 1225
rect 406 1220 407 1224
rect 411 1220 412 1224
rect 406 1219 412 1220
rect 446 1224 452 1225
rect 446 1220 447 1224
rect 451 1220 452 1224
rect 446 1219 452 1220
rect 486 1224 492 1225
rect 486 1220 487 1224
rect 491 1220 492 1224
rect 486 1219 492 1220
rect 526 1224 532 1225
rect 526 1220 527 1224
rect 531 1220 532 1224
rect 526 1219 532 1220
rect 566 1224 572 1225
rect 566 1220 567 1224
rect 571 1220 572 1224
rect 566 1219 572 1220
rect 606 1224 612 1225
rect 606 1220 607 1224
rect 611 1220 612 1224
rect 606 1219 612 1220
rect 654 1224 660 1225
rect 654 1220 655 1224
rect 659 1220 660 1224
rect 654 1219 660 1220
rect 702 1224 708 1225
rect 702 1220 703 1224
rect 707 1220 708 1224
rect 702 1219 708 1220
rect 750 1224 756 1225
rect 750 1220 751 1224
rect 755 1220 756 1224
rect 750 1219 756 1220
rect 798 1224 804 1225
rect 798 1220 799 1224
rect 803 1220 804 1224
rect 798 1219 804 1220
rect 846 1224 852 1225
rect 846 1220 847 1224
rect 851 1220 852 1224
rect 846 1219 852 1220
rect 894 1224 900 1225
rect 894 1220 895 1224
rect 899 1220 900 1224
rect 894 1219 900 1220
rect 942 1224 948 1225
rect 942 1220 943 1224
rect 947 1220 948 1224
rect 942 1219 948 1220
rect 990 1224 996 1225
rect 990 1220 991 1224
rect 995 1220 996 1224
rect 990 1219 996 1220
rect 1038 1224 1044 1225
rect 1038 1220 1039 1224
rect 1043 1220 1044 1224
rect 1038 1219 1044 1220
rect 1102 1224 1108 1225
rect 1102 1220 1103 1224
rect 1107 1220 1108 1224
rect 1102 1219 1108 1220
rect 1174 1224 1180 1225
rect 1174 1220 1175 1224
rect 1179 1220 1180 1224
rect 1174 1219 1180 1220
rect 1254 1224 1260 1225
rect 1288 1224 1328 1226
rect 1254 1220 1255 1224
rect 1259 1220 1260 1224
rect 1327 1223 1328 1224
rect 1332 1223 1333 1227
rect 1327 1222 1333 1223
rect 1342 1224 1348 1225
rect 1254 1219 1260 1220
rect 1342 1220 1343 1224
rect 1347 1220 1348 1224
rect 1342 1219 1348 1220
rect 1414 1224 1420 1225
rect 1414 1220 1415 1224
rect 1419 1220 1420 1224
rect 1414 1219 1420 1220
rect 1446 1221 1452 1222
rect 110 1216 116 1217
rect 1446 1217 1447 1221
rect 1451 1217 1452 1221
rect 1446 1216 1452 1217
rect 399 1215 405 1216
rect 399 1211 400 1215
rect 404 1214 405 1215
rect 458 1215 464 1216
rect 458 1214 459 1215
rect 404 1212 459 1214
rect 404 1211 405 1212
rect 399 1210 405 1211
rect 458 1211 459 1212
rect 463 1211 464 1215
rect 458 1210 464 1211
rect 495 1215 501 1216
rect 495 1211 496 1215
rect 500 1214 501 1215
rect 690 1215 696 1216
rect 690 1214 691 1215
rect 500 1212 691 1214
rect 500 1211 501 1212
rect 495 1210 501 1211
rect 690 1211 691 1212
rect 695 1211 696 1215
rect 690 1210 696 1211
rect 759 1215 765 1216
rect 759 1211 760 1215
rect 764 1214 765 1215
rect 810 1215 816 1216
rect 810 1214 811 1215
rect 764 1212 811 1214
rect 764 1211 765 1212
rect 759 1210 765 1211
rect 810 1211 811 1212
rect 815 1211 816 1215
rect 810 1210 816 1211
rect 855 1215 861 1216
rect 855 1211 856 1215
rect 860 1214 861 1215
rect 906 1215 912 1216
rect 906 1214 907 1215
rect 860 1212 907 1214
rect 860 1211 861 1212
rect 855 1210 861 1211
rect 906 1211 907 1212
rect 911 1211 912 1215
rect 906 1210 912 1211
rect 951 1215 957 1216
rect 951 1211 952 1215
rect 956 1214 957 1215
rect 1002 1215 1008 1216
rect 1002 1214 1003 1215
rect 956 1212 1003 1214
rect 956 1211 957 1212
rect 951 1210 957 1211
rect 1002 1211 1003 1212
rect 1007 1211 1008 1215
rect 1002 1210 1008 1211
rect 1047 1215 1053 1216
rect 1047 1211 1048 1215
rect 1052 1214 1053 1215
rect 1114 1215 1120 1216
rect 1114 1214 1115 1215
rect 1052 1212 1115 1214
rect 1052 1211 1053 1212
rect 1047 1210 1053 1211
rect 1114 1211 1115 1212
rect 1119 1211 1120 1215
rect 1114 1210 1120 1211
rect 1183 1215 1189 1216
rect 1183 1211 1184 1215
rect 1188 1214 1189 1215
rect 1266 1215 1272 1216
rect 1266 1214 1267 1215
rect 1188 1212 1267 1214
rect 1188 1211 1189 1212
rect 1183 1210 1189 1211
rect 1266 1211 1267 1212
rect 1271 1211 1272 1215
rect 1266 1210 1272 1211
rect 1294 1215 1300 1216
rect 1294 1211 1295 1215
rect 1299 1214 1300 1215
rect 1351 1215 1357 1216
rect 1351 1214 1352 1215
rect 1299 1212 1352 1214
rect 1299 1211 1300 1212
rect 1294 1210 1300 1211
rect 1351 1211 1352 1212
rect 1356 1211 1357 1215
rect 1351 1210 1357 1211
rect 335 1207 341 1208
rect 110 1203 116 1204
rect 110 1199 111 1203
rect 115 1199 116 1203
rect 335 1203 336 1207
rect 340 1206 341 1207
rect 346 1207 352 1208
rect 346 1206 347 1207
rect 340 1204 347 1206
rect 340 1203 341 1204
rect 335 1202 341 1203
rect 346 1203 347 1204
rect 351 1203 352 1207
rect 375 1207 381 1208
rect 375 1206 376 1207
rect 346 1202 352 1203
rect 356 1204 376 1206
rect 335 1199 341 1200
rect 110 1198 116 1199
rect 326 1198 332 1199
rect 326 1194 327 1198
rect 331 1194 332 1198
rect 335 1195 336 1199
rect 340 1198 341 1199
rect 356 1198 358 1204
rect 375 1203 376 1204
rect 380 1203 381 1207
rect 415 1207 421 1208
rect 415 1206 416 1207
rect 375 1202 381 1203
rect 396 1204 416 1206
rect 375 1199 381 1200
rect 340 1196 358 1198
rect 366 1198 372 1199
rect 340 1195 341 1196
rect 335 1194 341 1195
rect 366 1194 367 1198
rect 371 1194 372 1198
rect 375 1195 376 1199
rect 380 1198 381 1199
rect 396 1198 398 1204
rect 415 1203 416 1204
rect 420 1203 421 1207
rect 455 1207 461 1208
rect 455 1206 456 1207
rect 415 1202 421 1203
rect 436 1204 456 1206
rect 415 1199 421 1200
rect 380 1196 398 1198
rect 406 1198 412 1199
rect 380 1195 381 1196
rect 375 1194 381 1195
rect 406 1194 407 1198
rect 411 1194 412 1198
rect 415 1195 416 1199
rect 420 1198 421 1199
rect 436 1198 438 1204
rect 455 1203 456 1204
rect 460 1203 461 1207
rect 535 1207 541 1208
rect 535 1206 536 1207
rect 455 1202 461 1203
rect 516 1204 536 1206
rect 455 1199 464 1200
rect 495 1199 501 1200
rect 420 1196 438 1198
rect 446 1198 452 1199
rect 420 1195 421 1196
rect 415 1194 421 1195
rect 446 1194 447 1198
rect 451 1194 452 1198
rect 455 1195 456 1199
rect 463 1195 464 1199
rect 455 1194 464 1195
rect 486 1198 492 1199
rect 486 1194 487 1198
rect 491 1194 492 1198
rect 495 1195 496 1199
rect 500 1198 501 1199
rect 516 1198 518 1204
rect 535 1203 536 1204
rect 540 1203 541 1207
rect 575 1207 581 1208
rect 575 1206 576 1207
rect 535 1202 541 1203
rect 556 1204 576 1206
rect 535 1199 541 1200
rect 500 1196 518 1198
rect 526 1198 532 1199
rect 500 1195 501 1196
rect 495 1194 501 1195
rect 526 1194 527 1198
rect 531 1194 532 1198
rect 535 1195 536 1199
rect 540 1198 541 1199
rect 556 1198 558 1204
rect 575 1203 576 1204
rect 580 1203 581 1207
rect 615 1207 621 1208
rect 615 1206 616 1207
rect 575 1202 581 1203
rect 596 1204 616 1206
rect 575 1199 581 1200
rect 540 1196 558 1198
rect 566 1198 572 1199
rect 540 1195 541 1196
rect 535 1194 541 1195
rect 566 1194 567 1198
rect 571 1194 572 1198
rect 575 1195 576 1199
rect 580 1198 581 1199
rect 596 1198 598 1204
rect 615 1203 616 1204
rect 620 1203 621 1207
rect 663 1207 669 1208
rect 663 1206 664 1207
rect 615 1202 621 1203
rect 640 1204 664 1206
rect 615 1199 621 1200
rect 580 1196 598 1198
rect 606 1198 612 1199
rect 580 1195 581 1196
rect 575 1194 581 1195
rect 606 1194 607 1198
rect 611 1194 612 1198
rect 615 1195 616 1199
rect 620 1198 621 1199
rect 640 1198 642 1204
rect 663 1203 664 1204
rect 668 1203 669 1207
rect 711 1207 717 1208
rect 711 1206 712 1207
rect 663 1202 669 1203
rect 688 1204 712 1206
rect 663 1199 669 1200
rect 620 1196 642 1198
rect 654 1198 660 1199
rect 620 1195 621 1196
rect 615 1194 621 1195
rect 654 1194 655 1198
rect 659 1194 660 1198
rect 663 1195 664 1199
rect 668 1198 669 1199
rect 688 1198 690 1204
rect 711 1203 712 1204
rect 716 1203 717 1207
rect 711 1202 717 1203
rect 807 1207 813 1208
rect 807 1203 808 1207
rect 812 1206 813 1207
rect 903 1207 909 1208
rect 812 1204 843 1206
rect 812 1203 813 1204
rect 807 1202 813 1203
rect 759 1199 768 1200
rect 807 1199 816 1200
rect 668 1196 690 1198
rect 702 1198 708 1199
rect 668 1195 669 1196
rect 663 1194 669 1195
rect 702 1194 703 1198
rect 707 1194 708 1198
rect 750 1198 756 1199
rect 326 1193 332 1194
rect 366 1193 372 1194
rect 406 1193 412 1194
rect 446 1193 452 1194
rect 486 1193 492 1194
rect 526 1193 532 1194
rect 566 1193 572 1194
rect 606 1193 612 1194
rect 654 1193 660 1194
rect 702 1193 708 1194
rect 711 1195 717 1196
rect 170 1191 176 1192
rect 170 1190 171 1191
rect 145 1188 171 1190
rect 145 1184 147 1188
rect 170 1187 171 1188
rect 175 1187 176 1191
rect 170 1186 176 1187
rect 414 1191 420 1192
rect 414 1187 415 1191
rect 419 1190 420 1191
rect 694 1191 700 1192
rect 694 1190 695 1191
rect 419 1188 434 1190
rect 419 1187 420 1188
rect 414 1186 420 1187
rect 432 1184 434 1188
rect 473 1188 695 1190
rect 473 1184 475 1188
rect 694 1187 695 1188
rect 699 1187 700 1191
rect 711 1191 712 1195
rect 716 1194 717 1195
rect 750 1194 751 1198
rect 755 1194 756 1198
rect 759 1195 760 1199
rect 767 1195 768 1199
rect 759 1194 768 1195
rect 798 1198 804 1199
rect 798 1194 799 1198
rect 803 1194 804 1198
rect 807 1195 808 1199
rect 815 1195 816 1199
rect 807 1194 816 1195
rect 716 1192 746 1194
rect 750 1193 756 1194
rect 798 1193 804 1194
rect 716 1191 717 1192
rect 711 1190 717 1191
rect 744 1190 746 1192
rect 778 1191 784 1192
rect 778 1190 779 1191
rect 744 1188 779 1190
rect 694 1186 700 1187
rect 778 1187 779 1188
rect 783 1187 784 1191
rect 841 1190 843 1204
rect 903 1203 904 1207
rect 908 1206 909 1207
rect 922 1207 928 1208
rect 922 1206 923 1207
rect 908 1204 923 1206
rect 908 1203 909 1204
rect 903 1202 909 1203
rect 922 1203 923 1204
rect 927 1203 928 1207
rect 922 1202 928 1203
rect 999 1207 1005 1208
rect 999 1203 1000 1207
rect 1004 1206 1005 1207
rect 1111 1207 1117 1208
rect 1004 1204 1050 1206
rect 1004 1203 1005 1204
rect 999 1202 1005 1203
rect 1048 1200 1050 1204
rect 1111 1203 1112 1207
rect 1116 1206 1117 1207
rect 1263 1207 1269 1208
rect 1116 1204 1161 1206
rect 1116 1203 1117 1204
rect 1111 1202 1117 1203
rect 903 1199 912 1200
rect 999 1199 1008 1200
rect 1047 1199 1053 1200
rect 1111 1199 1120 1200
rect 846 1198 852 1199
rect 846 1194 847 1198
rect 851 1194 852 1198
rect 894 1198 900 1199
rect 846 1193 852 1194
rect 855 1195 861 1196
rect 855 1191 856 1195
rect 860 1191 861 1195
rect 894 1194 895 1198
rect 899 1194 900 1198
rect 903 1195 904 1199
rect 911 1195 912 1199
rect 903 1194 912 1195
rect 942 1198 948 1199
rect 942 1194 943 1198
rect 947 1194 948 1198
rect 990 1198 996 1199
rect 894 1193 900 1194
rect 942 1193 948 1194
rect 951 1195 957 1196
rect 855 1190 861 1191
rect 951 1191 952 1195
rect 956 1191 957 1195
rect 990 1194 991 1198
rect 995 1194 996 1198
rect 999 1195 1000 1199
rect 1007 1195 1008 1199
rect 999 1194 1008 1195
rect 1038 1198 1044 1199
rect 1038 1194 1039 1198
rect 1043 1194 1044 1198
rect 1047 1195 1048 1199
rect 1052 1195 1053 1199
rect 1047 1194 1053 1195
rect 1102 1198 1108 1199
rect 1102 1194 1103 1198
rect 1107 1194 1108 1198
rect 1111 1195 1112 1199
rect 1119 1195 1120 1199
rect 1111 1194 1120 1195
rect 990 1193 996 1194
rect 1038 1193 1044 1194
rect 1102 1193 1108 1194
rect 951 1190 957 1191
rect 1114 1191 1120 1192
rect 1114 1190 1115 1191
rect 841 1188 858 1190
rect 953 1188 1022 1190
rect 778 1186 784 1187
rect 1020 1186 1022 1188
rect 1048 1188 1115 1190
rect 1048 1186 1050 1188
rect 1114 1187 1115 1188
rect 1119 1187 1120 1191
rect 1159 1190 1161 1204
rect 1263 1203 1264 1207
rect 1268 1206 1269 1207
rect 1423 1207 1429 1208
rect 1268 1204 1310 1206
rect 1268 1203 1269 1204
rect 1263 1202 1269 1203
rect 1263 1199 1272 1200
rect 1174 1198 1180 1199
rect 1174 1194 1175 1198
rect 1179 1194 1180 1198
rect 1254 1198 1260 1199
rect 1174 1193 1180 1194
rect 1183 1195 1189 1196
rect 1183 1191 1184 1195
rect 1188 1191 1189 1195
rect 1254 1194 1255 1198
rect 1259 1194 1260 1198
rect 1263 1195 1264 1199
rect 1271 1195 1272 1199
rect 1263 1194 1272 1195
rect 1254 1193 1260 1194
rect 1183 1190 1189 1191
rect 1282 1191 1288 1192
rect 1282 1190 1283 1191
rect 1159 1188 1186 1190
rect 1241 1188 1283 1190
rect 1114 1186 1120 1187
rect 1020 1184 1050 1186
rect 1241 1184 1243 1188
rect 1282 1187 1283 1188
rect 1287 1187 1288 1191
rect 1308 1190 1310 1204
rect 1423 1203 1424 1207
rect 1428 1206 1429 1207
rect 1431 1207 1437 1208
rect 1431 1206 1432 1207
rect 1428 1204 1432 1206
rect 1428 1203 1429 1204
rect 1423 1202 1429 1203
rect 1431 1203 1432 1204
rect 1436 1203 1437 1207
rect 1431 1202 1437 1203
rect 1446 1203 1452 1204
rect 1423 1199 1432 1200
rect 1342 1198 1348 1199
rect 1342 1194 1343 1198
rect 1347 1194 1348 1198
rect 1414 1198 1420 1199
rect 1342 1193 1348 1194
rect 1351 1195 1357 1196
rect 1351 1191 1352 1195
rect 1356 1191 1357 1195
rect 1414 1194 1415 1198
rect 1419 1194 1420 1198
rect 1423 1195 1424 1199
rect 1431 1195 1432 1199
rect 1446 1199 1447 1203
rect 1451 1199 1452 1203
rect 1446 1198 1452 1199
rect 1423 1194 1432 1195
rect 1414 1193 1420 1194
rect 1351 1190 1357 1191
rect 1308 1188 1354 1190
rect 1282 1186 1288 1187
rect 143 1183 149 1184
rect 343 1183 352 1184
rect 431 1183 437 1184
rect 471 1183 477 1184
rect 919 1183 928 1184
rect 1239 1183 1245 1184
rect 1423 1183 1429 1184
rect 134 1182 140 1183
rect 134 1178 135 1182
rect 139 1178 140 1182
rect 143 1179 144 1183
rect 148 1179 149 1183
rect 143 1178 149 1179
rect 158 1182 164 1183
rect 158 1178 159 1182
rect 163 1178 164 1182
rect 182 1182 188 1183
rect 110 1177 116 1178
rect 134 1177 140 1178
rect 158 1177 164 1178
rect 167 1179 173 1180
rect 110 1173 111 1177
rect 115 1173 116 1177
rect 167 1175 168 1179
rect 172 1175 173 1179
rect 182 1178 183 1182
rect 187 1178 188 1182
rect 206 1182 212 1183
rect 182 1177 188 1178
rect 191 1179 197 1180
rect 167 1174 173 1175
rect 191 1175 192 1179
rect 196 1175 197 1179
rect 206 1178 207 1182
rect 211 1178 212 1182
rect 230 1182 236 1183
rect 206 1177 212 1178
rect 215 1179 221 1180
rect 191 1174 197 1175
rect 215 1175 216 1179
rect 220 1178 221 1179
rect 230 1178 231 1182
rect 235 1178 236 1182
rect 254 1182 260 1183
rect 220 1176 227 1178
rect 230 1177 236 1178
rect 239 1179 245 1180
rect 220 1175 221 1176
rect 215 1174 221 1175
rect 110 1172 116 1173
rect 169 1166 171 1174
rect 193 1170 195 1174
rect 215 1171 221 1172
rect 215 1170 216 1171
rect 193 1168 216 1170
rect 215 1167 216 1168
rect 220 1167 221 1171
rect 225 1170 227 1176
rect 239 1175 240 1179
rect 244 1178 245 1179
rect 254 1178 255 1182
rect 259 1178 260 1182
rect 278 1182 284 1183
rect 244 1176 250 1178
rect 254 1177 260 1178
rect 263 1179 269 1180
rect 244 1175 245 1176
rect 239 1174 245 1175
rect 239 1171 245 1172
rect 239 1170 240 1171
rect 225 1168 240 1170
rect 215 1166 221 1167
rect 239 1167 240 1168
rect 244 1167 245 1171
rect 239 1166 245 1167
rect 248 1166 250 1176
rect 263 1175 264 1179
rect 268 1175 269 1179
rect 278 1178 279 1182
rect 283 1178 284 1182
rect 302 1182 308 1183
rect 278 1177 284 1178
rect 287 1179 293 1180
rect 263 1174 269 1175
rect 287 1175 288 1179
rect 292 1178 293 1179
rect 302 1178 303 1182
rect 307 1178 308 1182
rect 334 1182 340 1183
rect 292 1176 298 1178
rect 302 1177 308 1178
rect 311 1179 320 1180
rect 292 1175 293 1176
rect 287 1174 293 1175
rect 265 1170 267 1174
rect 287 1171 293 1172
rect 287 1170 288 1171
rect 265 1168 288 1170
rect 287 1167 288 1168
rect 292 1167 293 1171
rect 296 1170 298 1176
rect 311 1175 312 1179
rect 319 1175 320 1179
rect 334 1178 335 1182
rect 339 1178 340 1182
rect 343 1179 344 1183
rect 351 1179 352 1183
rect 343 1178 352 1179
rect 382 1182 388 1183
rect 382 1178 383 1182
rect 387 1178 388 1182
rect 422 1182 428 1183
rect 334 1177 340 1178
rect 382 1177 388 1178
rect 391 1179 397 1180
rect 311 1174 320 1175
rect 391 1175 392 1179
rect 396 1175 397 1179
rect 422 1178 423 1182
rect 427 1178 428 1182
rect 431 1179 432 1183
rect 436 1179 437 1183
rect 431 1178 437 1179
rect 462 1182 468 1183
rect 462 1178 463 1182
rect 467 1178 468 1182
rect 471 1179 472 1183
rect 476 1179 477 1183
rect 471 1178 477 1179
rect 502 1182 508 1183
rect 502 1178 503 1182
rect 507 1178 508 1182
rect 542 1182 548 1183
rect 422 1177 428 1178
rect 462 1177 468 1178
rect 502 1177 508 1178
rect 511 1179 517 1180
rect 391 1174 397 1175
rect 511 1175 512 1179
rect 516 1175 517 1179
rect 542 1178 543 1182
rect 547 1178 548 1182
rect 582 1182 588 1183
rect 542 1177 548 1178
rect 551 1179 557 1180
rect 511 1174 517 1175
rect 551 1175 552 1179
rect 556 1175 557 1179
rect 582 1178 583 1182
rect 587 1178 588 1182
rect 622 1182 628 1183
rect 582 1177 588 1178
rect 591 1179 597 1180
rect 551 1174 557 1175
rect 591 1175 592 1179
rect 596 1175 597 1179
rect 622 1178 623 1182
rect 627 1178 628 1182
rect 670 1182 676 1183
rect 622 1177 628 1178
rect 631 1179 637 1180
rect 591 1174 597 1175
rect 631 1175 632 1179
rect 636 1175 637 1179
rect 670 1178 671 1182
rect 675 1178 676 1182
rect 718 1182 724 1183
rect 670 1177 676 1178
rect 679 1179 685 1180
rect 631 1174 637 1175
rect 679 1175 680 1179
rect 684 1175 685 1179
rect 718 1178 719 1182
rect 723 1178 724 1182
rect 766 1182 772 1183
rect 718 1177 724 1178
rect 727 1179 733 1180
rect 679 1174 685 1175
rect 727 1175 728 1179
rect 732 1175 733 1179
rect 766 1178 767 1182
rect 771 1178 772 1182
rect 814 1182 820 1183
rect 766 1177 772 1178
rect 775 1179 781 1180
rect 727 1174 733 1175
rect 775 1175 776 1179
rect 780 1175 781 1179
rect 814 1178 815 1182
rect 819 1178 820 1182
rect 862 1182 868 1183
rect 814 1177 820 1178
rect 823 1179 829 1180
rect 775 1174 781 1175
rect 823 1175 824 1179
rect 828 1178 829 1179
rect 862 1178 863 1182
rect 867 1178 868 1182
rect 910 1182 916 1183
rect 828 1176 850 1178
rect 862 1177 868 1178
rect 871 1179 877 1180
rect 828 1175 829 1176
rect 823 1174 829 1175
rect 311 1171 317 1172
rect 311 1170 312 1171
rect 296 1168 312 1170
rect 287 1166 293 1167
rect 311 1167 312 1168
rect 316 1167 317 1171
rect 311 1166 317 1167
rect 343 1171 349 1172
rect 343 1167 344 1171
rect 348 1170 349 1171
rect 392 1170 394 1174
rect 348 1168 394 1170
rect 471 1171 477 1172
rect 348 1167 349 1168
rect 343 1166 349 1167
rect 398 1167 404 1168
rect 169 1164 195 1166
rect 248 1164 267 1166
rect 191 1163 197 1164
rect 110 1159 116 1160
rect 110 1155 111 1159
rect 115 1155 116 1159
rect 191 1159 192 1163
rect 196 1159 197 1163
rect 191 1158 197 1159
rect 263 1163 269 1164
rect 263 1159 264 1163
rect 268 1159 269 1163
rect 398 1163 399 1167
rect 403 1166 404 1167
rect 431 1167 437 1168
rect 431 1166 432 1167
rect 403 1164 432 1166
rect 403 1163 404 1164
rect 398 1162 404 1163
rect 431 1163 432 1164
rect 436 1163 437 1167
rect 471 1167 472 1171
rect 476 1170 477 1171
rect 512 1170 514 1174
rect 476 1168 514 1170
rect 476 1167 477 1168
rect 471 1166 477 1167
rect 552 1166 554 1174
rect 593 1166 595 1174
rect 632 1166 634 1174
rect 679 1166 681 1174
rect 728 1166 730 1174
rect 777 1166 779 1174
rect 848 1170 850 1176
rect 871 1175 872 1179
rect 876 1178 877 1179
rect 910 1178 911 1182
rect 915 1178 916 1182
rect 919 1179 920 1183
rect 927 1179 928 1183
rect 919 1178 928 1179
rect 958 1182 964 1183
rect 958 1178 959 1182
rect 963 1178 964 1182
rect 1006 1182 1012 1183
rect 876 1176 898 1178
rect 910 1177 916 1178
rect 958 1177 964 1178
rect 967 1179 973 1180
rect 876 1175 877 1176
rect 871 1174 877 1175
rect 871 1171 877 1172
rect 871 1170 872 1171
rect 848 1168 872 1170
rect 871 1167 872 1168
rect 876 1167 877 1171
rect 896 1170 898 1176
rect 967 1175 968 1179
rect 972 1178 973 1179
rect 998 1179 1004 1180
rect 998 1178 999 1179
rect 972 1176 999 1178
rect 972 1175 973 1176
rect 967 1174 973 1175
rect 998 1175 999 1176
rect 1003 1175 1004 1179
rect 1006 1178 1007 1182
rect 1011 1178 1012 1182
rect 1054 1182 1060 1183
rect 1006 1177 1012 1178
rect 1015 1179 1021 1180
rect 998 1174 1004 1175
rect 1015 1175 1016 1179
rect 1020 1175 1021 1179
rect 1054 1178 1055 1182
rect 1059 1178 1060 1182
rect 1102 1182 1108 1183
rect 1054 1177 1060 1178
rect 1063 1179 1069 1180
rect 1015 1174 1021 1175
rect 1063 1175 1064 1179
rect 1068 1175 1069 1179
rect 1102 1178 1103 1182
rect 1107 1178 1108 1182
rect 1150 1182 1156 1183
rect 1102 1177 1108 1178
rect 1111 1179 1117 1180
rect 1063 1174 1069 1175
rect 1111 1175 1112 1179
rect 1116 1175 1117 1179
rect 1150 1178 1151 1182
rect 1155 1178 1156 1182
rect 1190 1182 1196 1183
rect 1150 1177 1156 1178
rect 1159 1179 1165 1180
rect 1111 1174 1117 1175
rect 1159 1175 1160 1179
rect 1164 1178 1165 1179
rect 1182 1179 1188 1180
rect 1182 1178 1183 1179
rect 1164 1176 1183 1178
rect 1164 1175 1165 1176
rect 1159 1174 1165 1175
rect 1182 1175 1183 1176
rect 1187 1175 1188 1179
rect 1190 1178 1191 1182
rect 1195 1178 1196 1182
rect 1230 1182 1236 1183
rect 1190 1177 1196 1178
rect 1199 1179 1205 1180
rect 1182 1174 1188 1175
rect 1199 1175 1200 1179
rect 1204 1175 1205 1179
rect 1230 1178 1231 1182
rect 1235 1178 1236 1182
rect 1239 1179 1240 1183
rect 1244 1179 1245 1183
rect 1239 1178 1245 1179
rect 1270 1182 1276 1183
rect 1270 1178 1271 1182
rect 1275 1178 1276 1182
rect 1310 1182 1316 1183
rect 1230 1177 1236 1178
rect 1270 1177 1276 1178
rect 1279 1179 1285 1180
rect 1199 1174 1205 1175
rect 1279 1175 1280 1179
rect 1284 1175 1285 1179
rect 1310 1178 1311 1182
rect 1315 1178 1316 1182
rect 1350 1182 1356 1183
rect 1310 1177 1316 1178
rect 1319 1179 1325 1180
rect 1279 1174 1285 1175
rect 1319 1175 1320 1179
rect 1324 1175 1325 1179
rect 1350 1178 1351 1182
rect 1355 1178 1356 1182
rect 1390 1182 1396 1183
rect 1350 1177 1356 1178
rect 1359 1179 1368 1180
rect 1319 1174 1325 1175
rect 1359 1175 1360 1179
rect 1367 1175 1368 1179
rect 1390 1178 1391 1182
rect 1395 1178 1396 1182
rect 1414 1182 1420 1183
rect 1390 1177 1396 1178
rect 1399 1179 1405 1180
rect 1359 1174 1368 1175
rect 1399 1175 1400 1179
rect 1404 1175 1405 1179
rect 1414 1178 1415 1182
rect 1419 1178 1420 1182
rect 1423 1179 1424 1183
rect 1428 1182 1429 1183
rect 1431 1183 1437 1184
rect 1431 1182 1432 1183
rect 1428 1180 1432 1182
rect 1428 1179 1429 1180
rect 1423 1178 1429 1179
rect 1431 1179 1432 1180
rect 1436 1179 1437 1183
rect 1431 1178 1437 1179
rect 1414 1177 1420 1178
rect 1446 1177 1452 1178
rect 1399 1174 1405 1175
rect 919 1171 925 1172
rect 919 1170 920 1171
rect 896 1168 920 1170
rect 871 1166 877 1167
rect 919 1167 920 1168
rect 924 1167 925 1171
rect 919 1166 925 1167
rect 967 1171 973 1172
rect 967 1167 968 1171
rect 972 1170 973 1171
rect 1016 1170 1018 1174
rect 972 1168 1018 1170
rect 972 1167 973 1168
rect 967 1166 973 1167
rect 1065 1166 1067 1174
rect 1113 1166 1115 1174
rect 532 1164 554 1166
rect 572 1164 595 1166
rect 612 1164 634 1166
rect 657 1164 681 1166
rect 704 1164 730 1166
rect 752 1164 779 1166
rect 1040 1164 1067 1166
rect 1088 1164 1115 1166
rect 1201 1166 1203 1174
rect 1281 1166 1283 1174
rect 1321 1170 1323 1174
rect 1359 1171 1365 1172
rect 1359 1170 1360 1171
rect 1321 1168 1360 1170
rect 1359 1167 1360 1168
rect 1364 1167 1365 1171
rect 1401 1170 1403 1174
rect 1446 1173 1447 1177
rect 1451 1173 1452 1177
rect 1446 1172 1452 1173
rect 1423 1171 1429 1172
rect 1423 1170 1424 1171
rect 1401 1168 1424 1170
rect 1359 1166 1365 1167
rect 1423 1167 1424 1168
rect 1428 1167 1429 1171
rect 1423 1166 1429 1167
rect 1201 1164 1243 1166
rect 1281 1164 1323 1166
rect 431 1162 437 1163
rect 511 1163 517 1164
rect 263 1158 269 1159
rect 391 1159 397 1160
rect 110 1154 116 1155
rect 134 1156 140 1157
rect 158 1156 164 1157
rect 182 1156 188 1157
rect 134 1152 135 1156
rect 139 1152 140 1156
rect 134 1151 140 1152
rect 143 1155 152 1156
rect 143 1151 144 1155
rect 151 1151 152 1155
rect 158 1152 159 1156
rect 163 1152 164 1156
rect 158 1151 164 1152
rect 167 1155 176 1156
rect 167 1151 168 1155
rect 175 1151 176 1155
rect 182 1152 183 1156
rect 187 1152 188 1156
rect 182 1151 188 1152
rect 206 1156 212 1157
rect 206 1152 207 1156
rect 211 1152 212 1156
rect 206 1151 212 1152
rect 230 1156 236 1157
rect 230 1152 231 1156
rect 235 1152 236 1156
rect 230 1151 236 1152
rect 254 1156 260 1157
rect 254 1152 255 1156
rect 259 1152 260 1156
rect 254 1151 260 1152
rect 278 1156 284 1157
rect 278 1152 279 1156
rect 283 1152 284 1156
rect 278 1151 284 1152
rect 302 1156 308 1157
rect 302 1152 303 1156
rect 307 1152 308 1156
rect 302 1151 308 1152
rect 334 1156 340 1157
rect 334 1152 335 1156
rect 339 1152 340 1156
rect 334 1151 340 1152
rect 382 1156 388 1157
rect 382 1152 383 1156
rect 387 1152 388 1156
rect 391 1155 392 1159
rect 396 1158 397 1159
rect 414 1159 420 1160
rect 414 1158 415 1159
rect 396 1156 415 1158
rect 396 1155 397 1156
rect 391 1154 397 1155
rect 414 1155 415 1156
rect 419 1155 420 1159
rect 511 1159 512 1163
rect 516 1162 517 1163
rect 532 1162 534 1164
rect 516 1160 534 1162
rect 516 1159 517 1160
rect 511 1158 517 1159
rect 551 1159 557 1160
rect 414 1154 420 1155
rect 422 1156 428 1157
rect 382 1151 388 1152
rect 422 1152 423 1156
rect 427 1152 428 1156
rect 422 1151 428 1152
rect 462 1156 468 1157
rect 462 1152 463 1156
rect 467 1152 468 1156
rect 462 1151 468 1152
rect 502 1156 508 1157
rect 502 1152 503 1156
rect 507 1152 508 1156
rect 502 1151 508 1152
rect 542 1156 548 1157
rect 542 1152 543 1156
rect 547 1152 548 1156
rect 551 1155 552 1159
rect 556 1158 557 1159
rect 572 1158 574 1164
rect 556 1156 574 1158
rect 591 1159 597 1160
rect 582 1156 588 1157
rect 556 1155 557 1156
rect 551 1154 557 1155
rect 542 1151 548 1152
rect 582 1152 583 1156
rect 587 1152 588 1156
rect 591 1155 592 1159
rect 596 1158 597 1159
rect 612 1158 614 1164
rect 596 1156 614 1158
rect 631 1159 637 1160
rect 622 1156 628 1157
rect 596 1155 597 1156
rect 591 1154 597 1155
rect 582 1151 588 1152
rect 622 1152 623 1156
rect 627 1152 628 1156
rect 631 1155 632 1159
rect 636 1158 637 1159
rect 657 1158 659 1164
rect 636 1156 659 1158
rect 679 1159 685 1160
rect 670 1156 676 1157
rect 636 1155 637 1156
rect 631 1154 637 1155
rect 622 1151 628 1152
rect 670 1152 671 1156
rect 675 1152 676 1156
rect 679 1155 680 1159
rect 684 1158 685 1159
rect 704 1158 706 1164
rect 684 1156 706 1158
rect 727 1159 733 1160
rect 718 1156 724 1157
rect 684 1155 685 1156
rect 679 1154 685 1155
rect 670 1151 676 1152
rect 718 1152 719 1156
rect 723 1152 724 1156
rect 727 1155 728 1159
rect 732 1158 733 1159
rect 752 1158 754 1164
rect 1015 1163 1021 1164
rect 732 1156 754 1158
rect 775 1159 784 1160
rect 766 1156 772 1157
rect 732 1155 733 1156
rect 727 1154 733 1155
rect 718 1151 724 1152
rect 766 1152 767 1156
rect 771 1152 772 1156
rect 775 1155 776 1159
rect 783 1155 784 1159
rect 1015 1159 1016 1163
rect 1020 1162 1021 1163
rect 1040 1162 1042 1164
rect 1020 1160 1042 1162
rect 1020 1159 1021 1160
rect 1015 1158 1021 1159
rect 1063 1159 1069 1160
rect 775 1154 784 1155
rect 814 1156 820 1157
rect 862 1156 868 1157
rect 766 1151 772 1152
rect 814 1152 815 1156
rect 819 1152 820 1156
rect 823 1155 829 1156
rect 823 1152 824 1155
rect 814 1151 820 1152
rect 822 1151 824 1152
rect 828 1151 829 1155
rect 862 1152 863 1156
rect 867 1152 868 1156
rect 862 1151 868 1152
rect 910 1156 916 1157
rect 910 1152 911 1156
rect 915 1152 916 1156
rect 910 1151 916 1152
rect 958 1156 964 1157
rect 958 1152 959 1156
rect 963 1152 964 1156
rect 958 1151 964 1152
rect 1006 1156 1012 1157
rect 1006 1152 1007 1156
rect 1011 1152 1012 1156
rect 1006 1151 1012 1152
rect 1054 1156 1060 1157
rect 1054 1152 1055 1156
rect 1059 1152 1060 1156
rect 1063 1155 1064 1159
rect 1068 1158 1069 1159
rect 1088 1158 1090 1164
rect 1239 1163 1245 1164
rect 1068 1156 1090 1158
rect 1111 1159 1120 1160
rect 1102 1156 1108 1157
rect 1068 1155 1069 1156
rect 1063 1154 1069 1155
rect 1054 1151 1060 1152
rect 1102 1152 1103 1156
rect 1107 1152 1108 1156
rect 1111 1155 1112 1159
rect 1119 1155 1120 1159
rect 1199 1159 1208 1160
rect 1111 1154 1120 1155
rect 1150 1156 1156 1157
rect 1190 1156 1196 1157
rect 1102 1151 1108 1152
rect 1150 1152 1151 1156
rect 1155 1152 1156 1156
rect 1150 1151 1156 1152
rect 1159 1155 1165 1156
rect 1159 1151 1160 1155
rect 1164 1154 1165 1155
rect 1182 1155 1188 1156
rect 1182 1154 1183 1155
rect 1164 1152 1183 1154
rect 1164 1151 1165 1152
rect 143 1150 152 1151
rect 167 1150 176 1151
rect 822 1147 823 1151
rect 827 1150 829 1151
rect 1159 1150 1165 1151
rect 1182 1151 1183 1152
rect 1187 1151 1188 1155
rect 1190 1152 1191 1156
rect 1195 1152 1196 1156
rect 1199 1155 1200 1159
rect 1207 1155 1208 1159
rect 1239 1159 1240 1163
rect 1244 1159 1245 1163
rect 1239 1158 1245 1159
rect 1319 1163 1325 1164
rect 1319 1159 1320 1163
rect 1324 1159 1325 1163
rect 1319 1158 1325 1159
rect 1446 1159 1452 1160
rect 1199 1154 1208 1155
rect 1230 1156 1236 1157
rect 1190 1151 1196 1152
rect 1230 1152 1231 1156
rect 1235 1152 1236 1156
rect 1230 1151 1236 1152
rect 1270 1156 1276 1157
rect 1310 1156 1316 1157
rect 1270 1152 1271 1156
rect 1275 1152 1276 1156
rect 1270 1151 1276 1152
rect 1279 1155 1288 1156
rect 1279 1151 1280 1155
rect 1287 1151 1288 1155
rect 1310 1152 1311 1156
rect 1315 1152 1316 1156
rect 1310 1151 1316 1152
rect 1350 1156 1356 1157
rect 1350 1152 1351 1156
rect 1355 1152 1356 1156
rect 1350 1151 1356 1152
rect 1390 1156 1396 1157
rect 1414 1156 1420 1157
rect 1390 1152 1391 1156
rect 1395 1152 1396 1156
rect 1390 1151 1396 1152
rect 1399 1155 1408 1156
rect 1399 1151 1400 1155
rect 1407 1151 1408 1155
rect 1414 1152 1415 1156
rect 1419 1152 1420 1156
rect 1446 1155 1447 1159
rect 1451 1155 1452 1159
rect 1446 1154 1452 1155
rect 1414 1151 1420 1152
rect 1182 1150 1188 1151
rect 1279 1150 1288 1151
rect 1399 1150 1408 1151
rect 827 1147 828 1150
rect 822 1146 828 1147
rect 134 1144 140 1145
rect 110 1141 116 1142
rect 110 1137 111 1141
rect 115 1137 116 1141
rect 134 1140 135 1144
rect 139 1140 140 1144
rect 134 1139 140 1140
rect 158 1144 164 1145
rect 158 1140 159 1144
rect 163 1140 164 1144
rect 158 1139 164 1140
rect 182 1144 188 1145
rect 182 1140 183 1144
rect 187 1140 188 1144
rect 182 1139 188 1140
rect 214 1144 220 1145
rect 214 1140 215 1144
rect 219 1140 220 1144
rect 214 1139 220 1140
rect 254 1144 260 1145
rect 254 1140 255 1144
rect 259 1140 260 1144
rect 254 1139 260 1140
rect 294 1144 300 1145
rect 294 1140 295 1144
rect 299 1140 300 1144
rect 294 1139 300 1140
rect 334 1144 340 1145
rect 334 1140 335 1144
rect 339 1140 340 1144
rect 334 1139 340 1140
rect 374 1144 380 1145
rect 374 1140 375 1144
rect 379 1140 380 1144
rect 374 1139 380 1140
rect 414 1144 420 1145
rect 414 1140 415 1144
rect 419 1140 420 1144
rect 414 1139 420 1140
rect 462 1144 468 1145
rect 462 1140 463 1144
rect 467 1140 468 1144
rect 462 1139 468 1140
rect 518 1144 524 1145
rect 518 1140 519 1144
rect 523 1140 524 1144
rect 518 1139 524 1140
rect 582 1144 588 1145
rect 582 1140 583 1144
rect 587 1140 588 1144
rect 582 1139 588 1140
rect 646 1144 652 1145
rect 646 1140 647 1144
rect 651 1140 652 1144
rect 646 1139 652 1140
rect 710 1144 716 1145
rect 710 1140 711 1144
rect 715 1140 716 1144
rect 710 1139 716 1140
rect 766 1144 772 1145
rect 766 1140 767 1144
rect 771 1140 772 1144
rect 766 1139 772 1140
rect 830 1144 836 1145
rect 830 1140 831 1144
rect 835 1140 836 1144
rect 830 1139 836 1140
rect 886 1144 892 1145
rect 886 1140 887 1144
rect 891 1140 892 1144
rect 886 1139 892 1140
rect 942 1144 948 1145
rect 942 1140 943 1144
rect 947 1140 948 1144
rect 942 1139 948 1140
rect 998 1144 1004 1145
rect 998 1140 999 1144
rect 1003 1140 1004 1144
rect 998 1139 1004 1140
rect 1054 1144 1060 1145
rect 1054 1140 1055 1144
rect 1059 1140 1060 1144
rect 1054 1139 1060 1140
rect 1102 1144 1108 1145
rect 1102 1140 1103 1144
rect 1107 1140 1108 1144
rect 1102 1139 1108 1140
rect 1150 1144 1156 1145
rect 1150 1140 1151 1144
rect 1155 1140 1156 1144
rect 1150 1139 1156 1140
rect 1190 1144 1196 1145
rect 1190 1140 1191 1144
rect 1195 1140 1196 1144
rect 1190 1139 1196 1140
rect 1230 1144 1236 1145
rect 1230 1140 1231 1144
rect 1235 1140 1236 1144
rect 1230 1139 1236 1140
rect 1270 1144 1276 1145
rect 1270 1140 1271 1144
rect 1275 1140 1276 1144
rect 1270 1139 1276 1140
rect 1310 1144 1316 1145
rect 1310 1140 1311 1144
rect 1315 1140 1316 1144
rect 1310 1139 1316 1140
rect 1350 1144 1356 1145
rect 1350 1140 1351 1144
rect 1355 1140 1356 1144
rect 1350 1139 1356 1140
rect 1390 1144 1396 1145
rect 1390 1140 1391 1144
rect 1395 1140 1396 1144
rect 1390 1139 1396 1140
rect 1414 1144 1420 1145
rect 1414 1140 1415 1144
rect 1419 1140 1420 1144
rect 1414 1139 1420 1140
rect 1446 1141 1452 1142
rect 110 1136 116 1137
rect 1446 1137 1447 1141
rect 1451 1137 1452 1141
rect 1446 1136 1452 1137
rect 143 1135 149 1136
rect 143 1131 144 1135
rect 148 1134 149 1135
rect 170 1135 176 1136
rect 170 1134 171 1135
rect 148 1132 171 1134
rect 148 1131 149 1132
rect 143 1130 149 1131
rect 170 1131 171 1132
rect 175 1131 176 1135
rect 170 1130 176 1131
rect 223 1135 229 1136
rect 223 1131 224 1135
rect 228 1134 229 1135
rect 314 1135 320 1136
rect 314 1134 315 1135
rect 228 1132 315 1134
rect 228 1131 229 1132
rect 223 1130 229 1131
rect 314 1131 315 1132
rect 319 1131 320 1135
rect 314 1130 320 1131
rect 383 1135 389 1136
rect 383 1131 384 1135
rect 388 1134 389 1135
rect 426 1135 432 1136
rect 426 1134 427 1135
rect 388 1132 427 1134
rect 388 1131 389 1132
rect 383 1130 389 1131
rect 426 1131 427 1132
rect 431 1131 432 1135
rect 426 1130 432 1131
rect 471 1135 477 1136
rect 471 1131 472 1135
rect 476 1134 477 1135
rect 530 1135 536 1136
rect 530 1134 531 1135
rect 476 1132 531 1134
rect 476 1131 477 1132
rect 471 1130 477 1131
rect 530 1131 531 1132
rect 535 1131 536 1135
rect 530 1130 536 1131
rect 591 1135 597 1136
rect 591 1131 592 1135
rect 596 1134 597 1135
rect 658 1135 664 1136
rect 658 1134 659 1135
rect 596 1132 659 1134
rect 596 1131 597 1132
rect 591 1130 597 1131
rect 658 1131 659 1132
rect 663 1131 664 1135
rect 658 1130 664 1131
rect 694 1135 700 1136
rect 694 1131 695 1135
rect 699 1134 700 1135
rect 719 1135 725 1136
rect 719 1134 720 1135
rect 699 1132 720 1134
rect 699 1131 700 1132
rect 694 1130 700 1131
rect 719 1131 720 1132
rect 724 1131 725 1135
rect 719 1130 725 1131
rect 839 1135 845 1136
rect 839 1131 840 1135
rect 844 1134 845 1135
rect 898 1135 904 1136
rect 898 1134 899 1135
rect 844 1132 899 1134
rect 844 1131 845 1132
rect 839 1130 845 1131
rect 898 1131 899 1132
rect 903 1131 904 1135
rect 898 1130 904 1131
rect 951 1135 957 1136
rect 951 1131 952 1135
rect 956 1134 957 1135
rect 1010 1135 1016 1136
rect 1010 1134 1011 1135
rect 956 1132 1011 1134
rect 956 1131 957 1132
rect 951 1130 957 1131
rect 1010 1131 1011 1132
rect 1015 1131 1016 1135
rect 1010 1130 1016 1131
rect 1018 1135 1024 1136
rect 1018 1131 1019 1135
rect 1023 1134 1024 1135
rect 1063 1135 1069 1136
rect 1063 1134 1064 1135
rect 1023 1132 1064 1134
rect 1023 1131 1024 1132
rect 1018 1130 1024 1131
rect 1063 1131 1064 1132
rect 1068 1131 1069 1135
rect 1063 1130 1069 1131
rect 1279 1135 1285 1136
rect 1279 1131 1280 1135
rect 1284 1134 1285 1135
rect 1362 1135 1368 1136
rect 1362 1134 1363 1135
rect 1284 1132 1363 1134
rect 1284 1131 1285 1132
rect 1279 1130 1285 1131
rect 1362 1131 1363 1132
rect 1367 1131 1368 1135
rect 1362 1130 1368 1131
rect 1399 1135 1405 1136
rect 1399 1131 1400 1135
rect 1404 1134 1405 1135
rect 1431 1135 1437 1136
rect 1431 1134 1432 1135
rect 1404 1132 1432 1134
rect 1404 1131 1405 1132
rect 1399 1130 1405 1131
rect 1431 1131 1432 1132
rect 1436 1131 1437 1135
rect 1431 1130 1437 1131
rect 167 1127 173 1128
rect 110 1123 116 1124
rect 110 1119 111 1123
rect 115 1119 116 1123
rect 167 1123 168 1127
rect 172 1126 173 1127
rect 175 1127 181 1128
rect 175 1126 176 1127
rect 172 1124 176 1126
rect 172 1123 173 1124
rect 167 1122 173 1123
rect 175 1123 176 1124
rect 180 1123 181 1127
rect 175 1122 181 1123
rect 191 1127 200 1128
rect 191 1123 192 1127
rect 199 1123 200 1127
rect 263 1127 269 1128
rect 263 1126 264 1127
rect 191 1122 200 1123
rect 244 1124 264 1126
rect 143 1119 152 1120
rect 167 1119 176 1120
rect 223 1119 229 1120
rect 110 1118 116 1119
rect 134 1118 140 1119
rect 134 1114 135 1118
rect 139 1114 140 1118
rect 143 1115 144 1119
rect 151 1115 152 1119
rect 143 1114 152 1115
rect 158 1118 164 1119
rect 158 1114 159 1118
rect 163 1114 164 1118
rect 167 1115 168 1119
rect 175 1115 176 1119
rect 167 1114 176 1115
rect 182 1118 188 1119
rect 182 1114 183 1118
rect 187 1114 188 1118
rect 214 1118 220 1119
rect 134 1113 140 1114
rect 158 1113 164 1114
rect 182 1113 188 1114
rect 191 1115 197 1116
rect 191 1111 192 1115
rect 196 1111 197 1115
rect 214 1114 215 1118
rect 219 1114 220 1118
rect 223 1115 224 1119
rect 228 1118 229 1119
rect 244 1118 246 1124
rect 263 1123 264 1124
rect 268 1123 269 1127
rect 303 1127 309 1128
rect 303 1126 304 1127
rect 263 1122 269 1123
rect 284 1124 304 1126
rect 263 1119 269 1120
rect 228 1116 246 1118
rect 254 1118 260 1119
rect 228 1115 229 1116
rect 223 1114 229 1115
rect 254 1114 255 1118
rect 259 1114 260 1118
rect 263 1115 264 1119
rect 268 1118 269 1119
rect 284 1118 286 1124
rect 303 1123 304 1124
rect 308 1123 309 1127
rect 343 1127 349 1128
rect 343 1126 344 1127
rect 303 1122 309 1123
rect 324 1124 344 1126
rect 303 1119 309 1120
rect 268 1116 286 1118
rect 294 1118 300 1119
rect 268 1115 269 1116
rect 263 1114 269 1115
rect 294 1114 295 1118
rect 299 1114 300 1118
rect 303 1115 304 1119
rect 308 1118 309 1119
rect 324 1118 326 1124
rect 343 1123 344 1124
rect 348 1123 349 1127
rect 398 1127 404 1128
rect 398 1126 399 1127
rect 343 1122 349 1123
rect 368 1124 399 1126
rect 343 1119 349 1120
rect 308 1116 326 1118
rect 334 1118 340 1119
rect 308 1115 309 1116
rect 303 1114 309 1115
rect 334 1114 335 1118
rect 339 1114 340 1118
rect 343 1115 344 1119
rect 348 1118 349 1119
rect 368 1118 370 1124
rect 398 1123 399 1124
rect 403 1123 404 1127
rect 398 1122 404 1123
rect 423 1127 429 1128
rect 423 1123 424 1127
rect 428 1126 429 1127
rect 527 1127 533 1128
rect 428 1124 451 1126
rect 428 1123 429 1124
rect 423 1122 429 1123
rect 423 1119 432 1120
rect 348 1116 370 1118
rect 374 1118 380 1119
rect 348 1115 349 1116
rect 343 1114 349 1115
rect 374 1114 375 1118
rect 379 1114 380 1118
rect 414 1118 420 1119
rect 214 1113 220 1114
rect 254 1113 260 1114
rect 294 1113 300 1114
rect 334 1113 340 1114
rect 374 1113 380 1114
rect 383 1115 392 1116
rect 191 1110 197 1111
rect 383 1111 384 1115
rect 391 1111 392 1115
rect 414 1114 415 1118
rect 419 1114 420 1118
rect 423 1115 424 1119
rect 431 1115 432 1119
rect 423 1114 432 1115
rect 414 1113 420 1114
rect 383 1110 392 1111
rect 449 1110 451 1124
rect 527 1123 528 1127
rect 532 1126 533 1127
rect 655 1127 661 1128
rect 532 1124 562 1126
rect 532 1123 533 1124
rect 527 1122 533 1123
rect 527 1119 536 1120
rect 462 1118 468 1119
rect 462 1114 463 1118
rect 467 1114 468 1118
rect 518 1118 524 1119
rect 462 1113 468 1114
rect 471 1115 477 1116
rect 471 1111 472 1115
rect 476 1111 477 1115
rect 518 1114 519 1118
rect 523 1114 524 1118
rect 527 1115 528 1119
rect 535 1115 536 1119
rect 527 1114 536 1115
rect 518 1113 524 1114
rect 471 1110 477 1111
rect 560 1110 562 1124
rect 655 1123 656 1127
rect 660 1126 661 1127
rect 775 1127 781 1128
rect 660 1124 681 1126
rect 660 1123 661 1124
rect 655 1122 661 1123
rect 655 1119 664 1120
rect 582 1118 588 1119
rect 582 1114 583 1118
rect 587 1114 588 1118
rect 646 1118 652 1119
rect 582 1113 588 1114
rect 591 1115 597 1116
rect 591 1111 592 1115
rect 596 1111 597 1115
rect 646 1114 647 1118
rect 651 1114 652 1118
rect 655 1115 656 1119
rect 663 1115 664 1119
rect 655 1114 664 1115
rect 646 1113 652 1114
rect 591 1110 597 1111
rect 679 1110 681 1124
rect 775 1123 776 1127
rect 780 1126 781 1127
rect 895 1127 901 1128
rect 780 1124 842 1126
rect 780 1123 781 1124
rect 775 1122 781 1123
rect 840 1120 842 1124
rect 895 1123 896 1127
rect 900 1126 901 1127
rect 1007 1127 1013 1128
rect 900 1124 926 1126
rect 900 1123 901 1124
rect 895 1122 901 1123
rect 775 1119 781 1120
rect 710 1118 716 1119
rect 710 1114 711 1118
rect 715 1114 716 1118
rect 766 1118 772 1119
rect 710 1113 716 1114
rect 719 1115 725 1116
rect 719 1111 720 1115
rect 724 1111 725 1115
rect 766 1114 767 1118
rect 771 1114 772 1118
rect 775 1115 776 1119
rect 780 1118 781 1119
rect 822 1119 828 1120
rect 839 1119 845 1120
rect 895 1119 904 1120
rect 822 1118 823 1119
rect 780 1116 823 1118
rect 780 1115 781 1116
rect 775 1114 781 1115
rect 822 1115 823 1116
rect 827 1115 828 1119
rect 822 1114 828 1115
rect 830 1118 836 1119
rect 830 1114 831 1118
rect 835 1114 836 1118
rect 839 1115 840 1119
rect 844 1115 845 1119
rect 839 1114 845 1115
rect 886 1118 892 1119
rect 886 1114 887 1118
rect 891 1114 892 1118
rect 895 1115 896 1119
rect 903 1115 904 1119
rect 895 1114 904 1115
rect 766 1113 772 1114
rect 830 1113 836 1114
rect 886 1113 892 1114
rect 719 1110 725 1111
rect 924 1110 926 1124
rect 1007 1123 1008 1127
rect 1012 1126 1013 1127
rect 1071 1127 1077 1128
rect 1012 1124 1038 1126
rect 1012 1123 1013 1124
rect 1007 1122 1013 1123
rect 1007 1119 1016 1120
rect 942 1118 948 1119
rect 942 1114 943 1118
rect 947 1114 948 1118
rect 998 1118 1004 1119
rect 942 1113 948 1114
rect 951 1115 957 1116
rect 951 1111 952 1115
rect 956 1111 957 1115
rect 998 1114 999 1118
rect 1003 1114 1004 1118
rect 1007 1115 1008 1119
rect 1015 1115 1016 1119
rect 1007 1114 1016 1115
rect 998 1113 1004 1114
rect 951 1110 957 1111
rect 1036 1110 1038 1124
rect 1071 1123 1072 1127
rect 1076 1126 1077 1127
rect 1111 1127 1117 1128
rect 1111 1126 1112 1127
rect 1076 1124 1112 1126
rect 1076 1123 1077 1124
rect 1071 1122 1077 1123
rect 1111 1123 1112 1124
rect 1116 1123 1117 1127
rect 1159 1127 1165 1128
rect 1159 1126 1160 1127
rect 1111 1122 1117 1123
rect 1136 1124 1160 1126
rect 1111 1119 1117 1120
rect 1054 1118 1060 1119
rect 1054 1114 1055 1118
rect 1059 1114 1060 1118
rect 1102 1118 1108 1119
rect 1054 1113 1060 1114
rect 1063 1115 1069 1116
rect 1063 1111 1064 1115
rect 1068 1111 1069 1115
rect 1102 1114 1103 1118
rect 1107 1114 1108 1118
rect 1111 1115 1112 1119
rect 1116 1118 1117 1119
rect 1136 1118 1138 1124
rect 1159 1123 1160 1124
rect 1164 1123 1165 1127
rect 1199 1127 1205 1128
rect 1199 1126 1200 1127
rect 1159 1122 1165 1123
rect 1180 1124 1200 1126
rect 1159 1119 1165 1120
rect 1116 1116 1138 1118
rect 1150 1118 1156 1119
rect 1116 1115 1117 1116
rect 1111 1114 1117 1115
rect 1150 1114 1151 1118
rect 1155 1114 1156 1118
rect 1159 1115 1160 1119
rect 1164 1118 1165 1119
rect 1180 1118 1182 1124
rect 1199 1123 1200 1124
rect 1204 1123 1205 1127
rect 1239 1127 1245 1128
rect 1239 1126 1240 1127
rect 1199 1122 1205 1123
rect 1220 1124 1240 1126
rect 1199 1119 1205 1120
rect 1164 1116 1182 1118
rect 1190 1118 1196 1119
rect 1164 1115 1165 1116
rect 1159 1114 1165 1115
rect 1190 1114 1191 1118
rect 1195 1114 1196 1118
rect 1199 1115 1200 1119
rect 1204 1118 1205 1119
rect 1220 1118 1222 1124
rect 1239 1123 1240 1124
rect 1244 1123 1245 1127
rect 1319 1127 1325 1128
rect 1319 1126 1320 1127
rect 1239 1122 1245 1123
rect 1300 1124 1320 1126
rect 1279 1119 1285 1120
rect 1204 1116 1222 1118
rect 1230 1118 1236 1119
rect 1204 1115 1205 1116
rect 1199 1114 1205 1115
rect 1230 1114 1231 1118
rect 1235 1114 1236 1118
rect 1270 1118 1276 1119
rect 1102 1113 1108 1114
rect 1150 1113 1156 1114
rect 1190 1113 1196 1114
rect 1230 1113 1236 1114
rect 1239 1115 1245 1116
rect 1063 1110 1069 1111
rect 1182 1111 1188 1112
rect 175 1107 181 1108
rect 175 1103 176 1107
rect 180 1106 181 1107
rect 193 1106 195 1110
rect 449 1108 474 1110
rect 560 1108 595 1110
rect 679 1108 722 1110
rect 924 1108 954 1110
rect 1036 1108 1066 1110
rect 399 1107 405 1108
rect 399 1106 400 1107
rect 180 1104 195 1106
rect 360 1104 400 1106
rect 180 1103 181 1104
rect 175 1102 181 1103
rect 191 1099 200 1100
rect 335 1099 341 1100
rect 134 1098 140 1099
rect 134 1094 135 1098
rect 139 1094 140 1098
rect 158 1098 164 1099
rect 110 1093 116 1094
rect 134 1093 140 1094
rect 143 1095 149 1096
rect 110 1089 111 1093
rect 115 1089 116 1093
rect 143 1091 144 1095
rect 148 1091 149 1095
rect 158 1094 159 1098
rect 163 1094 164 1098
rect 182 1098 188 1099
rect 158 1093 164 1094
rect 167 1095 173 1096
rect 143 1090 149 1091
rect 167 1091 168 1095
rect 172 1091 173 1095
rect 182 1094 183 1098
rect 187 1094 188 1098
rect 191 1095 192 1099
rect 199 1095 200 1099
rect 191 1094 200 1095
rect 206 1098 212 1099
rect 206 1094 207 1098
rect 211 1094 212 1098
rect 246 1098 252 1099
rect 182 1093 188 1094
rect 206 1093 212 1094
rect 215 1095 224 1096
rect 167 1090 173 1091
rect 215 1091 216 1095
rect 223 1091 224 1095
rect 246 1094 247 1098
rect 251 1094 252 1098
rect 286 1098 292 1099
rect 246 1093 252 1094
rect 255 1095 261 1096
rect 215 1090 224 1091
rect 255 1091 256 1095
rect 260 1091 261 1095
rect 286 1094 287 1098
rect 291 1094 292 1098
rect 326 1098 332 1099
rect 286 1093 292 1094
rect 295 1095 301 1096
rect 255 1090 261 1091
rect 295 1091 296 1095
rect 300 1091 301 1095
rect 326 1094 327 1098
rect 331 1094 332 1098
rect 335 1095 336 1099
rect 340 1098 341 1099
rect 360 1098 362 1104
rect 399 1103 400 1104
rect 404 1103 405 1107
rect 399 1102 405 1103
rect 1122 1107 1128 1108
rect 1122 1103 1123 1107
rect 1127 1106 1128 1107
rect 1182 1107 1183 1111
rect 1187 1110 1188 1111
rect 1239 1111 1240 1115
rect 1244 1111 1245 1115
rect 1270 1114 1271 1118
rect 1275 1114 1276 1118
rect 1279 1115 1280 1119
rect 1284 1118 1285 1119
rect 1300 1118 1302 1124
rect 1319 1123 1320 1124
rect 1324 1123 1325 1127
rect 1359 1127 1365 1128
rect 1359 1126 1360 1127
rect 1319 1122 1325 1123
rect 1340 1124 1360 1126
rect 1319 1119 1325 1120
rect 1284 1116 1302 1118
rect 1310 1118 1316 1119
rect 1284 1115 1285 1116
rect 1279 1114 1285 1115
rect 1310 1114 1311 1118
rect 1315 1114 1316 1118
rect 1319 1115 1320 1119
rect 1324 1118 1325 1119
rect 1340 1118 1342 1124
rect 1359 1123 1360 1124
rect 1364 1123 1365 1127
rect 1359 1122 1365 1123
rect 1423 1127 1432 1128
rect 1423 1123 1424 1127
rect 1431 1123 1432 1127
rect 1423 1122 1432 1123
rect 1446 1123 1452 1124
rect 1399 1119 1408 1120
rect 1423 1119 1429 1120
rect 1324 1116 1342 1118
rect 1350 1118 1356 1119
rect 1324 1115 1325 1116
rect 1319 1114 1325 1115
rect 1350 1114 1351 1118
rect 1355 1114 1356 1118
rect 1390 1118 1396 1119
rect 1270 1113 1276 1114
rect 1310 1113 1316 1114
rect 1350 1113 1356 1114
rect 1359 1115 1365 1116
rect 1239 1110 1245 1111
rect 1359 1111 1360 1115
rect 1364 1114 1365 1115
rect 1375 1115 1381 1116
rect 1375 1114 1376 1115
rect 1364 1112 1376 1114
rect 1364 1111 1365 1112
rect 1359 1110 1365 1111
rect 1375 1111 1376 1112
rect 1380 1111 1381 1115
rect 1390 1114 1391 1118
rect 1395 1114 1396 1118
rect 1399 1115 1400 1119
rect 1407 1115 1408 1119
rect 1399 1114 1408 1115
rect 1414 1118 1420 1119
rect 1414 1114 1415 1118
rect 1419 1114 1420 1118
rect 1423 1115 1424 1119
rect 1428 1118 1429 1119
rect 1431 1119 1437 1120
rect 1431 1118 1432 1119
rect 1428 1116 1432 1118
rect 1428 1115 1429 1116
rect 1423 1114 1429 1115
rect 1431 1115 1432 1116
rect 1436 1115 1437 1119
rect 1446 1119 1447 1123
rect 1451 1119 1452 1123
rect 1446 1118 1452 1119
rect 1431 1114 1437 1115
rect 1390 1113 1396 1114
rect 1414 1113 1420 1114
rect 1375 1110 1381 1111
rect 1187 1108 1243 1110
rect 1187 1107 1188 1108
rect 1182 1106 1188 1107
rect 1338 1107 1344 1108
rect 1127 1104 1178 1106
rect 1127 1103 1128 1104
rect 1122 1102 1128 1103
rect 1176 1100 1178 1104
rect 1338 1103 1339 1107
rect 1343 1106 1344 1107
rect 1343 1104 1395 1106
rect 1343 1103 1344 1104
rect 1338 1102 1344 1103
rect 1393 1100 1395 1104
rect 1063 1099 1069 1100
rect 340 1096 362 1098
rect 366 1098 372 1099
rect 340 1095 341 1096
rect 335 1094 341 1095
rect 366 1094 367 1098
rect 371 1094 372 1098
rect 406 1098 412 1099
rect 326 1093 332 1094
rect 366 1093 372 1094
rect 375 1095 384 1096
rect 295 1090 301 1091
rect 375 1091 376 1095
rect 383 1091 384 1095
rect 406 1094 407 1098
rect 411 1094 412 1098
rect 454 1098 460 1099
rect 406 1093 412 1094
rect 415 1095 421 1096
rect 375 1090 384 1091
rect 415 1091 416 1095
rect 420 1091 421 1095
rect 454 1094 455 1098
rect 459 1094 460 1098
rect 502 1098 508 1099
rect 454 1093 460 1094
rect 463 1095 469 1096
rect 415 1090 421 1091
rect 463 1091 464 1095
rect 468 1094 469 1095
rect 502 1094 503 1098
rect 507 1094 508 1098
rect 558 1098 564 1099
rect 468 1092 490 1094
rect 502 1093 508 1094
rect 511 1095 517 1096
rect 468 1091 469 1092
rect 463 1090 469 1091
rect 110 1088 116 1089
rect 145 1086 147 1090
rect 169 1086 171 1090
rect 191 1087 197 1088
rect 191 1086 192 1087
rect 145 1084 163 1086
rect 169 1084 192 1086
rect 161 1082 163 1084
rect 191 1083 192 1084
rect 196 1083 197 1087
rect 191 1082 197 1083
rect 215 1087 221 1088
rect 215 1083 216 1087
rect 220 1086 221 1087
rect 257 1086 259 1090
rect 220 1084 259 1086
rect 220 1083 221 1084
rect 215 1082 221 1083
rect 296 1082 298 1090
rect 375 1087 381 1088
rect 161 1080 171 1082
rect 257 1080 298 1082
rect 335 1083 341 1084
rect 167 1079 173 1080
rect 110 1075 116 1076
rect 110 1071 111 1075
rect 115 1071 116 1075
rect 143 1075 149 1076
rect 110 1070 116 1071
rect 134 1072 140 1073
rect 134 1068 135 1072
rect 139 1068 140 1072
rect 143 1071 144 1075
rect 148 1071 149 1075
rect 167 1075 168 1079
rect 172 1075 173 1079
rect 167 1074 173 1075
rect 255 1079 261 1080
rect 255 1075 256 1079
rect 260 1075 261 1079
rect 335 1079 336 1083
rect 340 1082 341 1083
rect 366 1083 372 1084
rect 366 1082 367 1083
rect 340 1080 367 1082
rect 340 1079 341 1080
rect 335 1078 341 1079
rect 366 1079 367 1080
rect 371 1079 372 1083
rect 375 1083 376 1087
rect 380 1086 381 1087
rect 386 1087 392 1088
rect 386 1086 387 1087
rect 380 1084 387 1086
rect 380 1083 381 1084
rect 375 1082 381 1083
rect 386 1083 387 1084
rect 391 1083 392 1087
rect 417 1086 419 1090
rect 463 1087 469 1088
rect 463 1086 464 1087
rect 417 1084 464 1086
rect 386 1082 392 1083
rect 399 1083 405 1084
rect 366 1078 372 1079
rect 399 1079 400 1083
rect 404 1082 405 1083
rect 463 1083 464 1084
rect 468 1083 469 1087
rect 488 1086 490 1092
rect 511 1091 512 1095
rect 516 1094 517 1095
rect 558 1094 559 1098
rect 563 1094 564 1098
rect 606 1098 612 1099
rect 516 1092 542 1094
rect 558 1093 564 1094
rect 567 1095 573 1096
rect 516 1091 517 1092
rect 511 1090 517 1091
rect 511 1087 517 1088
rect 511 1086 512 1087
rect 488 1084 512 1086
rect 463 1082 469 1083
rect 511 1083 512 1084
rect 516 1083 517 1087
rect 540 1086 542 1092
rect 567 1091 568 1095
rect 572 1094 573 1095
rect 606 1094 607 1098
rect 611 1094 612 1098
rect 654 1098 660 1099
rect 572 1092 594 1094
rect 606 1093 612 1094
rect 615 1095 624 1096
rect 572 1091 573 1092
rect 567 1090 573 1091
rect 567 1087 573 1088
rect 567 1086 568 1087
rect 540 1084 568 1086
rect 511 1082 517 1083
rect 567 1083 568 1084
rect 572 1083 573 1087
rect 592 1086 594 1092
rect 615 1091 616 1095
rect 623 1091 624 1095
rect 654 1094 655 1098
rect 659 1094 660 1098
rect 702 1098 708 1099
rect 654 1093 660 1094
rect 663 1095 669 1096
rect 615 1090 624 1091
rect 663 1091 664 1095
rect 668 1094 669 1095
rect 702 1094 703 1098
rect 707 1094 708 1098
rect 742 1098 748 1099
rect 668 1092 681 1094
rect 702 1093 708 1094
rect 711 1095 717 1096
rect 668 1091 669 1092
rect 663 1090 669 1091
rect 615 1087 621 1088
rect 615 1086 616 1087
rect 592 1084 616 1086
rect 567 1082 573 1083
rect 615 1083 616 1084
rect 620 1083 621 1087
rect 679 1086 681 1092
rect 711 1091 712 1095
rect 716 1094 717 1095
rect 742 1094 743 1098
rect 747 1094 748 1098
rect 790 1098 796 1099
rect 716 1092 734 1094
rect 742 1093 748 1094
rect 751 1095 757 1096
rect 716 1091 717 1092
rect 711 1090 717 1091
rect 711 1087 717 1088
rect 711 1086 712 1087
rect 679 1084 712 1086
rect 615 1082 621 1083
rect 711 1083 712 1084
rect 716 1083 717 1087
rect 732 1086 734 1092
rect 751 1091 752 1095
rect 756 1094 757 1095
rect 790 1094 791 1098
rect 795 1094 796 1098
rect 838 1098 844 1099
rect 756 1092 778 1094
rect 790 1093 796 1094
rect 799 1095 805 1096
rect 756 1091 757 1092
rect 751 1090 757 1091
rect 751 1087 757 1088
rect 751 1086 752 1087
rect 732 1084 752 1086
rect 711 1082 717 1083
rect 751 1083 752 1084
rect 756 1083 757 1087
rect 776 1086 778 1092
rect 799 1091 800 1095
rect 804 1094 805 1095
rect 838 1094 839 1098
rect 843 1094 844 1098
rect 886 1098 892 1099
rect 804 1092 826 1094
rect 838 1093 844 1094
rect 847 1095 853 1096
rect 804 1091 805 1092
rect 799 1090 805 1091
rect 799 1087 805 1088
rect 799 1086 800 1087
rect 776 1084 800 1086
rect 751 1082 757 1083
rect 799 1083 800 1084
rect 804 1083 805 1087
rect 824 1086 826 1092
rect 847 1091 848 1095
rect 852 1094 853 1095
rect 886 1094 887 1098
rect 891 1094 892 1098
rect 942 1098 948 1099
rect 852 1092 874 1094
rect 886 1093 892 1094
rect 895 1095 901 1096
rect 852 1091 853 1092
rect 847 1090 853 1091
rect 847 1087 853 1088
rect 847 1086 848 1087
rect 824 1084 848 1086
rect 799 1082 805 1083
rect 847 1083 848 1084
rect 852 1083 853 1087
rect 872 1086 874 1092
rect 895 1091 896 1095
rect 900 1094 901 1095
rect 942 1094 943 1098
rect 947 1094 948 1098
rect 998 1098 1004 1099
rect 900 1092 926 1094
rect 942 1093 948 1094
rect 951 1095 957 1096
rect 900 1091 901 1092
rect 895 1090 901 1091
rect 895 1087 901 1088
rect 895 1086 896 1087
rect 872 1084 896 1086
rect 847 1082 853 1083
rect 895 1083 896 1084
rect 900 1083 901 1087
rect 924 1086 926 1092
rect 951 1091 952 1095
rect 956 1094 957 1095
rect 998 1094 999 1098
rect 1003 1094 1004 1098
rect 1054 1098 1060 1099
rect 956 1092 982 1094
rect 998 1093 1004 1094
rect 1007 1095 1016 1096
rect 956 1091 957 1092
rect 951 1090 957 1091
rect 951 1087 957 1088
rect 951 1086 952 1087
rect 924 1084 952 1086
rect 895 1082 901 1083
rect 951 1083 952 1084
rect 956 1083 957 1087
rect 980 1086 982 1092
rect 1007 1091 1008 1095
rect 1015 1091 1016 1095
rect 1054 1094 1055 1098
rect 1059 1094 1060 1098
rect 1063 1095 1064 1099
rect 1068 1098 1069 1099
rect 1071 1099 1077 1100
rect 1175 1099 1181 1100
rect 1391 1099 1397 1100
rect 1423 1099 1432 1100
rect 1071 1098 1072 1099
rect 1068 1096 1072 1098
rect 1068 1095 1069 1096
rect 1063 1094 1069 1095
rect 1071 1095 1072 1096
rect 1076 1095 1077 1099
rect 1071 1094 1077 1095
rect 1110 1098 1116 1099
rect 1110 1094 1111 1098
rect 1115 1094 1116 1098
rect 1166 1098 1172 1099
rect 1054 1093 1060 1094
rect 1110 1093 1116 1094
rect 1119 1095 1125 1096
rect 1007 1090 1016 1091
rect 1119 1091 1120 1095
rect 1124 1091 1125 1095
rect 1166 1094 1167 1098
rect 1171 1094 1172 1098
rect 1175 1095 1176 1099
rect 1180 1095 1181 1099
rect 1175 1094 1181 1095
rect 1214 1098 1220 1099
rect 1214 1094 1215 1098
rect 1219 1094 1220 1098
rect 1270 1098 1276 1099
rect 1166 1093 1172 1094
rect 1214 1093 1220 1094
rect 1223 1095 1229 1096
rect 1119 1090 1125 1091
rect 1223 1091 1224 1095
rect 1228 1094 1229 1095
rect 1262 1095 1268 1096
rect 1262 1094 1263 1095
rect 1228 1092 1263 1094
rect 1228 1091 1229 1092
rect 1223 1090 1229 1091
rect 1262 1091 1263 1092
rect 1267 1091 1268 1095
rect 1270 1094 1271 1098
rect 1275 1094 1276 1098
rect 1326 1098 1332 1099
rect 1270 1093 1276 1094
rect 1279 1095 1285 1096
rect 1262 1090 1268 1091
rect 1279 1091 1280 1095
rect 1284 1091 1285 1095
rect 1326 1094 1327 1098
rect 1331 1094 1332 1098
rect 1382 1098 1388 1099
rect 1326 1093 1332 1094
rect 1335 1095 1341 1096
rect 1279 1090 1285 1091
rect 1335 1091 1336 1095
rect 1340 1091 1341 1095
rect 1382 1094 1383 1098
rect 1387 1094 1388 1098
rect 1391 1095 1392 1099
rect 1396 1095 1397 1099
rect 1391 1094 1397 1095
rect 1414 1098 1420 1099
rect 1414 1094 1415 1098
rect 1419 1094 1420 1098
rect 1423 1095 1424 1099
rect 1431 1095 1432 1099
rect 1423 1094 1432 1095
rect 1382 1093 1388 1094
rect 1414 1093 1420 1094
rect 1446 1093 1452 1094
rect 1335 1090 1341 1091
rect 1007 1087 1013 1088
rect 1007 1086 1008 1087
rect 980 1084 1008 1086
rect 951 1082 957 1083
rect 1007 1083 1008 1084
rect 1012 1083 1013 1087
rect 1007 1082 1013 1083
rect 1063 1087 1069 1088
rect 1063 1083 1064 1087
rect 1068 1086 1069 1087
rect 1120 1086 1122 1090
rect 1068 1084 1122 1086
rect 1223 1087 1229 1088
rect 1068 1083 1069 1084
rect 1063 1082 1069 1083
rect 1138 1083 1144 1084
rect 404 1080 419 1082
rect 404 1079 405 1080
rect 399 1078 405 1079
rect 415 1079 421 1080
rect 255 1074 261 1075
rect 415 1075 416 1079
rect 420 1075 421 1079
rect 415 1074 421 1075
rect 1119 1079 1128 1080
rect 1119 1075 1120 1079
rect 1127 1075 1128 1079
rect 1138 1079 1139 1083
rect 1143 1082 1144 1083
rect 1175 1083 1181 1084
rect 1175 1082 1176 1083
rect 1143 1080 1176 1082
rect 1143 1079 1144 1080
rect 1138 1078 1144 1079
rect 1175 1079 1176 1080
rect 1180 1079 1181 1083
rect 1223 1083 1224 1087
rect 1228 1086 1229 1087
rect 1281 1086 1283 1090
rect 1228 1084 1283 1086
rect 1228 1083 1229 1084
rect 1223 1082 1229 1083
rect 1337 1082 1339 1090
rect 1446 1089 1447 1093
rect 1451 1089 1452 1093
rect 1446 1088 1452 1089
rect 1375 1087 1381 1088
rect 1375 1083 1376 1087
rect 1380 1086 1381 1087
rect 1391 1087 1397 1088
rect 1391 1086 1392 1087
rect 1380 1084 1392 1086
rect 1380 1083 1381 1084
rect 1375 1082 1381 1083
rect 1391 1083 1392 1084
rect 1396 1083 1397 1087
rect 1391 1082 1397 1083
rect 1281 1080 1339 1082
rect 1175 1078 1181 1079
rect 1279 1079 1285 1080
rect 1119 1074 1128 1075
rect 1279 1075 1280 1079
rect 1284 1075 1285 1079
rect 1279 1074 1285 1075
rect 1335 1075 1344 1076
rect 143 1070 149 1071
rect 158 1072 164 1073
rect 134 1067 140 1068
rect 158 1068 159 1072
rect 163 1068 164 1072
rect 158 1067 164 1068
rect 182 1072 188 1073
rect 182 1068 183 1072
rect 187 1068 188 1072
rect 182 1067 188 1068
rect 206 1072 212 1073
rect 206 1068 207 1072
rect 211 1068 212 1072
rect 206 1067 212 1068
rect 246 1072 252 1073
rect 246 1068 247 1072
rect 251 1068 252 1072
rect 246 1067 252 1068
rect 286 1072 292 1073
rect 326 1072 332 1073
rect 286 1068 287 1072
rect 291 1068 292 1072
rect 286 1067 292 1068
rect 295 1071 304 1072
rect 295 1067 296 1071
rect 303 1067 304 1071
rect 326 1068 327 1072
rect 331 1068 332 1072
rect 326 1067 332 1068
rect 366 1072 372 1073
rect 366 1068 367 1072
rect 371 1068 372 1072
rect 366 1067 372 1068
rect 406 1072 412 1073
rect 406 1068 407 1072
rect 411 1068 412 1072
rect 406 1067 412 1068
rect 454 1072 460 1073
rect 454 1068 455 1072
rect 459 1068 460 1072
rect 454 1067 460 1068
rect 502 1072 508 1073
rect 502 1068 503 1072
rect 507 1068 508 1072
rect 502 1067 508 1068
rect 558 1072 564 1073
rect 558 1068 559 1072
rect 563 1068 564 1072
rect 558 1067 564 1068
rect 606 1072 612 1073
rect 606 1068 607 1072
rect 611 1068 612 1072
rect 606 1067 612 1068
rect 654 1072 660 1073
rect 702 1072 708 1073
rect 654 1068 655 1072
rect 659 1068 660 1072
rect 654 1067 660 1068
rect 663 1071 669 1072
rect 663 1067 664 1071
rect 668 1070 669 1071
rect 694 1071 700 1072
rect 694 1070 695 1071
rect 668 1068 695 1070
rect 668 1067 669 1068
rect 295 1066 304 1067
rect 663 1066 669 1067
rect 694 1067 695 1068
rect 699 1067 700 1071
rect 702 1068 703 1072
rect 707 1068 708 1072
rect 702 1067 708 1068
rect 742 1072 748 1073
rect 742 1068 743 1072
rect 747 1068 748 1072
rect 742 1067 748 1068
rect 790 1072 796 1073
rect 790 1068 791 1072
rect 795 1068 796 1072
rect 790 1067 796 1068
rect 838 1072 844 1073
rect 838 1068 839 1072
rect 843 1068 844 1072
rect 838 1067 844 1068
rect 886 1072 892 1073
rect 886 1068 887 1072
rect 891 1068 892 1072
rect 886 1067 892 1068
rect 942 1072 948 1073
rect 942 1068 943 1072
rect 947 1068 948 1072
rect 942 1067 948 1068
rect 998 1072 1004 1073
rect 998 1068 999 1072
rect 1003 1068 1004 1072
rect 998 1067 1004 1068
rect 1054 1072 1060 1073
rect 1054 1068 1055 1072
rect 1059 1068 1060 1072
rect 1054 1067 1060 1068
rect 1110 1072 1116 1073
rect 1110 1068 1111 1072
rect 1115 1068 1116 1072
rect 1110 1067 1116 1068
rect 1166 1072 1172 1073
rect 1166 1068 1167 1072
rect 1171 1068 1172 1072
rect 1166 1067 1172 1068
rect 1214 1072 1220 1073
rect 1214 1068 1215 1072
rect 1219 1068 1220 1072
rect 1214 1067 1220 1068
rect 1270 1072 1276 1073
rect 1270 1068 1271 1072
rect 1275 1068 1276 1072
rect 1270 1067 1276 1068
rect 1326 1072 1332 1073
rect 1326 1068 1327 1072
rect 1331 1068 1332 1072
rect 1335 1071 1336 1075
rect 1343 1071 1344 1075
rect 1446 1075 1452 1076
rect 1335 1070 1344 1071
rect 1382 1072 1388 1073
rect 1326 1067 1332 1068
rect 1382 1068 1383 1072
rect 1387 1068 1388 1072
rect 1382 1067 1388 1068
rect 1414 1072 1420 1073
rect 1414 1068 1415 1072
rect 1419 1068 1420 1072
rect 1414 1067 1420 1068
rect 1423 1071 1432 1072
rect 1423 1067 1424 1071
rect 1431 1067 1432 1071
rect 1446 1071 1447 1075
rect 1451 1071 1452 1075
rect 1446 1070 1452 1071
rect 694 1066 700 1067
rect 1423 1066 1432 1067
rect 134 1060 140 1061
rect 110 1057 116 1058
rect 110 1053 111 1057
rect 115 1053 116 1057
rect 134 1056 135 1060
rect 139 1056 140 1060
rect 134 1055 140 1056
rect 158 1060 164 1061
rect 158 1056 159 1060
rect 163 1056 164 1060
rect 158 1055 164 1056
rect 182 1060 188 1061
rect 182 1056 183 1060
rect 187 1056 188 1060
rect 182 1055 188 1056
rect 206 1060 212 1061
rect 206 1056 207 1060
rect 211 1056 212 1060
rect 206 1055 212 1056
rect 230 1060 236 1061
rect 230 1056 231 1060
rect 235 1056 236 1060
rect 230 1055 236 1056
rect 270 1060 276 1061
rect 270 1056 271 1060
rect 275 1056 276 1060
rect 270 1055 276 1056
rect 310 1060 316 1061
rect 310 1056 311 1060
rect 315 1056 316 1060
rect 310 1055 316 1056
rect 350 1060 356 1061
rect 350 1056 351 1060
rect 355 1056 356 1060
rect 350 1055 356 1056
rect 390 1060 396 1061
rect 390 1056 391 1060
rect 395 1056 396 1060
rect 390 1055 396 1056
rect 430 1060 436 1061
rect 430 1056 431 1060
rect 435 1056 436 1060
rect 430 1055 436 1056
rect 470 1060 476 1061
rect 470 1056 471 1060
rect 475 1056 476 1060
rect 470 1055 476 1056
rect 510 1060 516 1061
rect 510 1056 511 1060
rect 515 1056 516 1060
rect 510 1055 516 1056
rect 550 1060 556 1061
rect 550 1056 551 1060
rect 555 1056 556 1060
rect 550 1055 556 1056
rect 590 1060 596 1061
rect 590 1056 591 1060
rect 595 1056 596 1060
rect 590 1055 596 1056
rect 630 1060 636 1061
rect 630 1056 631 1060
rect 635 1056 636 1060
rect 630 1055 636 1056
rect 670 1060 676 1061
rect 670 1056 671 1060
rect 675 1056 676 1060
rect 670 1055 676 1056
rect 710 1060 716 1061
rect 710 1056 711 1060
rect 715 1056 716 1060
rect 710 1055 716 1056
rect 742 1060 748 1061
rect 742 1056 743 1060
rect 747 1056 748 1060
rect 742 1055 748 1056
rect 782 1060 788 1061
rect 782 1056 783 1060
rect 787 1056 788 1060
rect 782 1055 788 1056
rect 822 1060 828 1061
rect 822 1056 823 1060
rect 827 1056 828 1060
rect 822 1055 828 1056
rect 870 1060 876 1061
rect 870 1056 871 1060
rect 875 1056 876 1060
rect 870 1055 876 1056
rect 918 1060 924 1061
rect 918 1056 919 1060
rect 923 1056 924 1060
rect 918 1055 924 1056
rect 974 1060 980 1061
rect 1030 1060 1036 1061
rect 974 1056 975 1060
rect 979 1056 980 1060
rect 974 1055 980 1056
rect 983 1059 989 1060
rect 983 1055 984 1059
rect 988 1058 989 1059
rect 1010 1059 1016 1060
rect 1010 1058 1011 1059
rect 988 1056 1011 1058
rect 988 1055 989 1056
rect 983 1054 989 1055
rect 1010 1055 1011 1056
rect 1015 1055 1016 1059
rect 1030 1056 1031 1060
rect 1035 1056 1036 1060
rect 1030 1055 1036 1056
rect 1078 1060 1084 1061
rect 1078 1056 1079 1060
rect 1083 1056 1084 1060
rect 1078 1055 1084 1056
rect 1126 1060 1132 1061
rect 1126 1056 1127 1060
rect 1131 1056 1132 1060
rect 1126 1055 1132 1056
rect 1174 1060 1180 1061
rect 1174 1056 1175 1060
rect 1179 1056 1180 1060
rect 1174 1055 1180 1056
rect 1222 1060 1228 1061
rect 1222 1056 1223 1060
rect 1227 1056 1228 1060
rect 1222 1055 1228 1056
rect 1270 1060 1276 1061
rect 1270 1056 1271 1060
rect 1275 1056 1276 1060
rect 1270 1055 1276 1056
rect 1326 1060 1332 1061
rect 1326 1056 1327 1060
rect 1331 1056 1332 1060
rect 1326 1055 1332 1056
rect 1382 1060 1388 1061
rect 1382 1056 1383 1060
rect 1387 1056 1388 1060
rect 1382 1055 1388 1056
rect 1414 1060 1420 1061
rect 1414 1056 1415 1060
rect 1419 1056 1420 1060
rect 1414 1055 1420 1056
rect 1446 1057 1452 1058
rect 1010 1054 1016 1055
rect 110 1052 116 1053
rect 1446 1053 1447 1057
rect 1451 1053 1452 1057
rect 1446 1052 1452 1053
rect 143 1051 149 1052
rect 143 1047 144 1051
rect 148 1050 149 1051
rect 170 1051 176 1052
rect 170 1050 171 1051
rect 148 1048 171 1050
rect 148 1047 149 1048
rect 143 1046 149 1047
rect 170 1047 171 1048
rect 175 1047 176 1051
rect 194 1051 200 1052
rect 194 1050 195 1051
rect 170 1046 176 1047
rect 185 1048 195 1050
rect 167 1043 173 1044
rect 110 1039 116 1040
rect 110 1035 111 1039
rect 115 1035 116 1039
rect 167 1039 168 1043
rect 172 1042 173 1043
rect 185 1042 187 1048
rect 194 1047 195 1048
rect 199 1047 200 1051
rect 218 1051 224 1052
rect 218 1050 219 1051
rect 194 1046 200 1047
rect 209 1048 219 1050
rect 172 1040 187 1042
rect 191 1043 197 1044
rect 172 1039 173 1040
rect 167 1038 173 1039
rect 191 1039 192 1043
rect 196 1042 197 1043
rect 209 1042 211 1048
rect 218 1047 219 1048
rect 223 1047 224 1051
rect 242 1051 248 1052
rect 242 1050 243 1051
rect 218 1046 224 1047
rect 233 1048 243 1050
rect 196 1040 211 1042
rect 215 1043 221 1044
rect 196 1039 197 1040
rect 191 1038 197 1039
rect 215 1039 216 1043
rect 220 1042 221 1043
rect 233 1042 235 1048
rect 242 1047 243 1048
rect 247 1047 248 1051
rect 242 1046 248 1047
rect 279 1051 285 1052
rect 279 1047 280 1051
rect 284 1050 285 1051
rect 322 1051 328 1052
rect 322 1050 323 1051
rect 284 1048 323 1050
rect 284 1047 285 1048
rect 279 1046 285 1047
rect 322 1047 323 1048
rect 327 1047 328 1051
rect 322 1046 328 1047
rect 359 1051 365 1052
rect 359 1047 360 1051
rect 364 1050 365 1051
rect 618 1051 624 1052
rect 618 1050 619 1051
rect 364 1048 619 1050
rect 364 1047 365 1048
rect 359 1046 365 1047
rect 618 1047 619 1048
rect 623 1047 624 1051
rect 618 1046 624 1047
rect 639 1051 645 1052
rect 639 1047 640 1051
rect 644 1050 645 1051
rect 774 1051 780 1052
rect 774 1050 775 1051
rect 644 1048 775 1050
rect 644 1047 645 1048
rect 639 1046 645 1047
rect 774 1047 775 1048
rect 779 1047 780 1051
rect 774 1046 780 1047
rect 831 1051 837 1052
rect 831 1047 832 1051
rect 836 1050 837 1051
rect 882 1051 888 1052
rect 882 1050 883 1051
rect 836 1048 883 1050
rect 836 1047 837 1048
rect 831 1046 837 1047
rect 882 1047 883 1048
rect 887 1047 888 1051
rect 882 1046 888 1047
rect 1183 1051 1189 1052
rect 1183 1047 1184 1051
rect 1188 1050 1189 1051
rect 1234 1051 1240 1052
rect 1234 1050 1235 1051
rect 1188 1048 1235 1050
rect 1188 1047 1189 1048
rect 1183 1046 1189 1047
rect 1234 1047 1235 1048
rect 1239 1047 1240 1051
rect 1234 1046 1240 1047
rect 1279 1051 1285 1052
rect 1279 1047 1280 1051
rect 1284 1050 1285 1051
rect 1338 1051 1344 1052
rect 1338 1050 1339 1051
rect 1284 1048 1339 1050
rect 1284 1047 1285 1048
rect 1279 1046 1285 1047
rect 1338 1047 1339 1048
rect 1343 1047 1344 1051
rect 1338 1046 1344 1047
rect 220 1040 235 1042
rect 239 1043 245 1044
rect 220 1039 221 1040
rect 215 1038 221 1039
rect 239 1039 240 1043
rect 244 1042 245 1043
rect 319 1043 325 1044
rect 319 1042 320 1043
rect 244 1040 283 1042
rect 244 1039 245 1040
rect 239 1038 245 1039
rect 281 1036 283 1040
rect 288 1040 320 1042
rect 143 1035 152 1036
rect 167 1035 176 1036
rect 191 1035 200 1036
rect 215 1035 224 1036
rect 239 1035 248 1036
rect 279 1035 285 1036
rect 110 1034 116 1035
rect 134 1034 140 1035
rect 134 1030 135 1034
rect 139 1030 140 1034
rect 143 1031 144 1035
rect 151 1031 152 1035
rect 143 1030 152 1031
rect 158 1034 164 1035
rect 158 1030 159 1034
rect 163 1030 164 1034
rect 167 1031 168 1035
rect 175 1031 176 1035
rect 167 1030 176 1031
rect 182 1034 188 1035
rect 182 1030 183 1034
rect 187 1030 188 1034
rect 191 1031 192 1035
rect 199 1031 200 1035
rect 191 1030 200 1031
rect 206 1034 212 1035
rect 206 1030 207 1034
rect 211 1030 212 1034
rect 215 1031 216 1035
rect 223 1031 224 1035
rect 215 1030 224 1031
rect 230 1034 236 1035
rect 230 1030 231 1034
rect 235 1030 236 1034
rect 239 1031 240 1035
rect 247 1031 248 1035
rect 239 1030 248 1031
rect 270 1034 276 1035
rect 270 1030 271 1034
rect 275 1030 276 1034
rect 279 1031 280 1035
rect 284 1031 285 1035
rect 279 1030 285 1031
rect 134 1029 140 1030
rect 158 1029 164 1030
rect 182 1029 188 1030
rect 206 1029 212 1030
rect 230 1029 236 1030
rect 270 1029 276 1030
rect 288 1026 290 1040
rect 319 1039 320 1040
rect 324 1039 325 1043
rect 399 1043 405 1044
rect 399 1042 400 1043
rect 319 1038 325 1039
rect 380 1040 400 1042
rect 319 1035 328 1036
rect 359 1035 365 1036
rect 310 1034 316 1035
rect 310 1030 311 1034
rect 315 1030 316 1034
rect 319 1031 320 1035
rect 327 1031 328 1035
rect 319 1030 328 1031
rect 350 1034 356 1035
rect 350 1030 351 1034
rect 355 1030 356 1034
rect 359 1031 360 1035
rect 364 1034 365 1035
rect 380 1034 382 1040
rect 399 1039 400 1040
rect 404 1039 405 1043
rect 439 1043 445 1044
rect 439 1042 440 1043
rect 399 1038 405 1039
rect 420 1040 440 1042
rect 399 1035 405 1036
rect 364 1032 382 1034
rect 390 1034 396 1035
rect 364 1031 365 1032
rect 359 1030 365 1031
rect 390 1030 391 1034
rect 395 1030 396 1034
rect 399 1031 400 1035
rect 404 1034 405 1035
rect 420 1034 422 1040
rect 439 1039 440 1040
rect 444 1039 445 1043
rect 479 1043 485 1044
rect 479 1042 480 1043
rect 439 1038 445 1039
rect 460 1040 480 1042
rect 439 1035 445 1036
rect 404 1032 422 1034
rect 430 1034 436 1035
rect 404 1031 405 1032
rect 399 1030 405 1031
rect 430 1030 431 1034
rect 435 1030 436 1034
rect 439 1031 440 1035
rect 444 1034 445 1035
rect 460 1034 462 1040
rect 479 1039 480 1040
rect 484 1039 485 1043
rect 519 1043 525 1044
rect 519 1042 520 1043
rect 479 1038 485 1039
rect 500 1040 520 1042
rect 479 1035 485 1036
rect 444 1032 462 1034
rect 470 1034 476 1035
rect 444 1031 445 1032
rect 439 1030 445 1031
rect 470 1030 471 1034
rect 475 1030 476 1034
rect 479 1031 480 1035
rect 484 1034 485 1035
rect 500 1034 502 1040
rect 519 1039 520 1040
rect 524 1039 525 1043
rect 559 1043 565 1044
rect 559 1042 560 1043
rect 519 1038 525 1039
rect 544 1040 560 1042
rect 519 1035 525 1036
rect 484 1032 502 1034
rect 510 1034 516 1035
rect 484 1031 485 1032
rect 479 1030 485 1031
rect 510 1030 511 1034
rect 515 1030 516 1034
rect 519 1031 520 1035
rect 524 1034 525 1035
rect 544 1034 546 1040
rect 559 1039 560 1040
rect 564 1039 565 1043
rect 599 1043 605 1044
rect 599 1042 600 1043
rect 559 1038 565 1039
rect 580 1040 600 1042
rect 559 1035 565 1036
rect 524 1032 546 1034
rect 550 1034 556 1035
rect 524 1031 525 1032
rect 519 1030 525 1031
rect 550 1030 551 1034
rect 555 1030 556 1034
rect 559 1031 560 1035
rect 564 1034 565 1035
rect 580 1034 582 1040
rect 599 1039 600 1040
rect 604 1039 605 1043
rect 679 1043 685 1044
rect 679 1042 680 1043
rect 599 1038 605 1039
rect 660 1040 680 1042
rect 639 1035 645 1036
rect 564 1032 582 1034
rect 590 1034 596 1035
rect 564 1031 565 1032
rect 559 1030 565 1031
rect 590 1030 591 1034
rect 595 1030 596 1034
rect 630 1034 636 1035
rect 310 1029 316 1030
rect 350 1029 356 1030
rect 390 1029 396 1030
rect 430 1029 436 1030
rect 470 1029 476 1030
rect 510 1029 516 1030
rect 550 1029 556 1030
rect 590 1029 596 1030
rect 599 1031 608 1032
rect 169 1024 290 1026
rect 538 1027 544 1028
rect 169 1020 171 1024
rect 538 1023 539 1027
rect 543 1026 544 1027
rect 599 1027 600 1031
rect 607 1027 608 1031
rect 630 1030 631 1034
rect 635 1030 636 1034
rect 639 1031 640 1035
rect 644 1034 645 1035
rect 660 1034 662 1040
rect 679 1039 680 1040
rect 684 1039 685 1043
rect 719 1043 725 1044
rect 719 1042 720 1043
rect 679 1038 685 1039
rect 700 1040 720 1042
rect 679 1035 685 1036
rect 644 1032 662 1034
rect 670 1034 676 1035
rect 644 1031 645 1032
rect 639 1030 645 1031
rect 670 1030 671 1034
rect 675 1030 676 1034
rect 679 1031 680 1035
rect 684 1034 685 1035
rect 700 1034 702 1040
rect 719 1039 720 1040
rect 724 1039 725 1043
rect 751 1043 757 1044
rect 751 1042 752 1043
rect 719 1038 725 1039
rect 736 1040 752 1042
rect 719 1035 725 1036
rect 684 1032 702 1034
rect 710 1034 716 1035
rect 684 1031 685 1032
rect 679 1030 685 1031
rect 710 1030 711 1034
rect 715 1030 716 1034
rect 719 1031 720 1035
rect 724 1034 725 1035
rect 736 1034 738 1040
rect 751 1039 752 1040
rect 756 1039 757 1043
rect 791 1043 797 1044
rect 791 1042 792 1043
rect 751 1038 757 1039
rect 772 1040 792 1042
rect 751 1035 757 1036
rect 724 1032 738 1034
rect 742 1034 748 1035
rect 724 1031 725 1032
rect 719 1030 725 1031
rect 742 1030 743 1034
rect 747 1030 748 1034
rect 751 1031 752 1035
rect 756 1034 757 1035
rect 772 1034 774 1040
rect 791 1039 792 1040
rect 796 1039 797 1043
rect 791 1038 797 1039
rect 879 1043 885 1044
rect 879 1039 880 1043
rect 884 1042 885 1043
rect 927 1043 933 1044
rect 884 1040 906 1042
rect 884 1039 885 1040
rect 879 1038 885 1039
rect 791 1035 800 1036
rect 879 1035 888 1036
rect 756 1032 774 1034
rect 782 1034 788 1035
rect 756 1031 757 1032
rect 751 1030 757 1031
rect 782 1030 783 1034
rect 787 1030 788 1034
rect 791 1031 792 1035
rect 799 1031 800 1035
rect 791 1030 800 1031
rect 822 1034 828 1035
rect 822 1030 823 1034
rect 827 1030 828 1034
rect 870 1034 876 1035
rect 630 1029 636 1030
rect 670 1029 676 1030
rect 710 1029 716 1030
rect 742 1029 748 1030
rect 782 1029 788 1030
rect 822 1029 828 1030
rect 831 1031 840 1032
rect 599 1026 608 1027
rect 831 1027 832 1031
rect 839 1027 840 1031
rect 870 1030 871 1034
rect 875 1030 876 1034
rect 879 1031 880 1035
rect 887 1031 888 1035
rect 879 1030 888 1031
rect 870 1029 876 1030
rect 831 1026 840 1027
rect 904 1026 906 1040
rect 927 1039 928 1043
rect 932 1042 933 1043
rect 1002 1043 1008 1044
rect 932 1040 986 1042
rect 932 1039 933 1040
rect 927 1038 933 1039
rect 984 1036 986 1040
rect 1002 1039 1003 1043
rect 1007 1042 1008 1043
rect 1039 1043 1045 1044
rect 1039 1042 1040 1043
rect 1007 1040 1040 1042
rect 1007 1039 1008 1040
rect 1002 1038 1008 1039
rect 1039 1039 1040 1040
rect 1044 1039 1045 1043
rect 1087 1043 1093 1044
rect 1087 1042 1088 1043
rect 1039 1038 1045 1039
rect 1064 1040 1088 1042
rect 983 1035 989 1036
rect 1039 1035 1045 1036
rect 918 1034 924 1035
rect 918 1030 919 1034
rect 923 1030 924 1034
rect 974 1034 980 1035
rect 918 1029 924 1030
rect 927 1031 933 1032
rect 927 1027 928 1031
rect 932 1027 933 1031
rect 974 1030 975 1034
rect 979 1030 980 1034
rect 983 1031 984 1035
rect 988 1031 989 1035
rect 983 1030 989 1031
rect 1030 1034 1036 1035
rect 1030 1030 1031 1034
rect 1035 1030 1036 1034
rect 1039 1031 1040 1035
rect 1044 1034 1045 1035
rect 1064 1034 1066 1040
rect 1087 1039 1088 1040
rect 1092 1039 1093 1043
rect 1135 1043 1141 1044
rect 1135 1042 1136 1043
rect 1087 1038 1093 1039
rect 1112 1040 1136 1042
rect 1087 1035 1093 1036
rect 1044 1032 1066 1034
rect 1078 1034 1084 1035
rect 1044 1031 1045 1032
rect 1039 1030 1045 1031
rect 1078 1030 1079 1034
rect 1083 1030 1084 1034
rect 1087 1031 1088 1035
rect 1092 1034 1093 1035
rect 1112 1034 1114 1040
rect 1135 1039 1136 1040
rect 1140 1039 1141 1043
rect 1135 1038 1141 1039
rect 1231 1043 1237 1044
rect 1231 1039 1232 1043
rect 1236 1042 1237 1043
rect 1262 1043 1268 1044
rect 1236 1040 1258 1042
rect 1236 1039 1237 1040
rect 1231 1038 1237 1039
rect 1135 1035 1144 1036
rect 1231 1035 1240 1036
rect 1092 1032 1114 1034
rect 1126 1034 1132 1035
rect 1092 1031 1093 1032
rect 1087 1030 1093 1031
rect 1126 1030 1127 1034
rect 1131 1030 1132 1034
rect 1135 1031 1136 1035
rect 1143 1031 1144 1035
rect 1135 1030 1144 1031
rect 1174 1034 1180 1035
rect 1174 1030 1175 1034
rect 1179 1030 1180 1034
rect 1222 1034 1228 1035
rect 974 1029 980 1030
rect 1030 1029 1036 1030
rect 1078 1029 1084 1030
rect 1126 1029 1132 1030
rect 1174 1029 1180 1030
rect 1183 1031 1192 1032
rect 927 1026 933 1027
rect 1183 1027 1184 1031
rect 1191 1027 1192 1031
rect 1222 1030 1223 1034
rect 1227 1030 1228 1034
rect 1231 1031 1232 1035
rect 1239 1031 1240 1035
rect 1231 1030 1240 1031
rect 1222 1029 1228 1030
rect 1183 1026 1192 1027
rect 1256 1026 1258 1040
rect 1262 1039 1263 1043
rect 1267 1042 1268 1043
rect 1335 1043 1341 1044
rect 1335 1042 1336 1043
rect 1267 1040 1336 1042
rect 1267 1039 1268 1040
rect 1262 1038 1268 1039
rect 1335 1039 1336 1040
rect 1340 1039 1341 1043
rect 1335 1038 1341 1039
rect 1391 1043 1400 1044
rect 1391 1039 1392 1043
rect 1399 1039 1400 1043
rect 1423 1043 1429 1044
rect 1423 1042 1424 1043
rect 1391 1038 1400 1039
rect 1408 1040 1424 1042
rect 1335 1035 1344 1036
rect 1391 1035 1397 1036
rect 1270 1034 1276 1035
rect 1270 1030 1271 1034
rect 1275 1030 1276 1034
rect 1326 1034 1332 1035
rect 1270 1029 1276 1030
rect 1279 1031 1285 1032
rect 1279 1027 1280 1031
rect 1284 1027 1285 1031
rect 1326 1030 1327 1034
rect 1331 1030 1332 1034
rect 1335 1031 1336 1035
rect 1343 1031 1344 1035
rect 1335 1030 1344 1031
rect 1382 1034 1388 1035
rect 1382 1030 1383 1034
rect 1387 1030 1388 1034
rect 1391 1031 1392 1035
rect 1396 1034 1397 1035
rect 1408 1034 1410 1040
rect 1423 1039 1424 1040
rect 1428 1039 1429 1043
rect 1423 1038 1429 1039
rect 1446 1039 1452 1040
rect 1423 1035 1432 1036
rect 1396 1032 1410 1034
rect 1414 1034 1420 1035
rect 1396 1031 1397 1032
rect 1391 1030 1397 1031
rect 1414 1030 1415 1034
rect 1419 1030 1420 1034
rect 1423 1031 1424 1035
rect 1431 1031 1432 1035
rect 1446 1035 1447 1039
rect 1451 1035 1452 1039
rect 1446 1034 1452 1035
rect 1423 1030 1432 1031
rect 1326 1029 1332 1030
rect 1382 1029 1388 1030
rect 1414 1029 1420 1030
rect 1279 1026 1285 1027
rect 543 1024 586 1026
rect 904 1024 930 1026
rect 1256 1024 1283 1026
rect 543 1023 544 1024
rect 538 1022 544 1023
rect 584 1020 586 1024
rect 774 1023 780 1024
rect 167 1019 173 1020
rect 583 1019 589 1020
rect 774 1019 775 1023
rect 779 1020 780 1023
rect 779 1019 781 1020
rect 999 1019 1008 1020
rect 1391 1019 1400 1020
rect 158 1018 164 1019
rect 158 1014 159 1018
rect 163 1014 164 1018
rect 167 1015 168 1019
rect 172 1015 173 1019
rect 167 1014 173 1015
rect 182 1018 188 1019
rect 182 1014 183 1018
rect 187 1014 188 1018
rect 206 1018 212 1019
rect 110 1013 116 1014
rect 158 1013 164 1014
rect 182 1013 188 1014
rect 191 1015 197 1016
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 191 1011 192 1015
rect 196 1011 197 1015
rect 206 1014 207 1018
rect 211 1014 212 1018
rect 230 1018 236 1019
rect 206 1013 212 1014
rect 215 1015 221 1016
rect 191 1010 197 1011
rect 215 1011 216 1015
rect 220 1011 221 1015
rect 230 1014 231 1018
rect 235 1014 236 1018
rect 262 1018 268 1019
rect 230 1013 236 1014
rect 239 1015 245 1016
rect 215 1010 221 1011
rect 239 1011 240 1015
rect 244 1011 245 1015
rect 262 1014 263 1018
rect 267 1014 268 1018
rect 302 1018 308 1019
rect 262 1013 268 1014
rect 271 1015 277 1016
rect 239 1010 245 1011
rect 271 1011 272 1015
rect 276 1011 277 1015
rect 302 1014 303 1018
rect 307 1014 308 1018
rect 342 1018 348 1019
rect 302 1013 308 1014
rect 311 1015 317 1016
rect 271 1010 277 1011
rect 311 1011 312 1015
rect 316 1011 317 1015
rect 342 1014 343 1018
rect 347 1014 348 1018
rect 382 1018 388 1019
rect 342 1013 348 1014
rect 351 1015 357 1016
rect 311 1010 317 1011
rect 351 1011 352 1015
rect 356 1011 357 1015
rect 382 1014 383 1018
rect 387 1014 388 1018
rect 430 1018 436 1019
rect 382 1013 388 1014
rect 391 1015 397 1016
rect 351 1010 357 1011
rect 391 1011 392 1015
rect 396 1014 397 1015
rect 410 1015 416 1016
rect 410 1014 411 1015
rect 396 1012 411 1014
rect 396 1011 397 1012
rect 391 1010 397 1011
rect 410 1011 411 1012
rect 415 1011 416 1015
rect 430 1014 431 1018
rect 435 1014 436 1018
rect 478 1018 484 1019
rect 430 1013 436 1014
rect 439 1015 445 1016
rect 410 1010 416 1011
rect 439 1011 440 1015
rect 444 1011 445 1015
rect 478 1014 479 1018
rect 483 1014 484 1018
rect 526 1018 532 1019
rect 478 1013 484 1014
rect 487 1015 493 1016
rect 439 1010 445 1011
rect 487 1011 488 1015
rect 492 1011 493 1015
rect 526 1014 527 1018
rect 531 1014 532 1018
rect 574 1018 580 1019
rect 526 1013 532 1014
rect 535 1015 541 1016
rect 487 1010 493 1011
rect 535 1011 536 1015
rect 540 1011 541 1015
rect 574 1014 575 1018
rect 579 1014 580 1018
rect 583 1015 584 1019
rect 588 1015 589 1019
rect 583 1014 589 1015
rect 622 1018 628 1019
rect 622 1014 623 1018
rect 627 1014 628 1018
rect 670 1018 676 1019
rect 574 1013 580 1014
rect 622 1013 628 1014
rect 631 1015 637 1016
rect 535 1010 541 1011
rect 631 1011 632 1015
rect 636 1014 637 1015
rect 670 1014 671 1018
rect 675 1014 676 1018
rect 718 1018 724 1019
rect 636 1012 658 1014
rect 670 1013 676 1014
rect 679 1015 685 1016
rect 636 1011 637 1012
rect 631 1010 637 1011
rect 110 1008 116 1009
rect 167 1007 173 1008
rect 167 1003 168 1007
rect 172 1006 173 1007
rect 193 1006 195 1010
rect 172 1004 195 1006
rect 172 1003 173 1004
rect 167 1002 173 1003
rect 217 1002 219 1010
rect 241 1002 243 1010
rect 272 1002 274 1010
rect 313 1002 315 1010
rect 353 1002 355 1010
rect 391 1007 397 1008
rect 391 1003 392 1007
rect 396 1006 397 1007
rect 440 1006 442 1010
rect 396 1004 442 1006
rect 396 1003 397 1004
rect 391 1002 397 1003
rect 488 1002 490 1010
rect 536 1002 538 1010
rect 583 1007 589 1008
rect 583 1003 584 1007
rect 588 1006 589 1007
rect 602 1007 608 1008
rect 602 1006 603 1007
rect 588 1004 603 1006
rect 588 1003 589 1004
rect 583 1002 589 1003
rect 602 1003 603 1004
rect 607 1003 608 1007
rect 656 1006 658 1012
rect 679 1011 680 1015
rect 684 1014 685 1015
rect 718 1014 719 1018
rect 723 1014 724 1018
rect 766 1018 772 1019
rect 774 1018 776 1019
rect 684 1012 706 1014
rect 718 1013 724 1014
rect 727 1015 733 1016
rect 684 1011 685 1012
rect 679 1010 685 1011
rect 679 1007 685 1008
rect 679 1006 680 1007
rect 656 1004 680 1006
rect 602 1002 608 1003
rect 679 1003 680 1004
rect 684 1003 685 1007
rect 704 1006 706 1012
rect 727 1011 728 1015
rect 732 1014 733 1015
rect 766 1014 767 1018
rect 771 1014 772 1018
rect 775 1015 776 1018
rect 780 1015 781 1019
rect 775 1014 781 1015
rect 822 1018 828 1019
rect 822 1014 823 1018
rect 827 1014 828 1018
rect 878 1018 884 1019
rect 732 1012 754 1014
rect 766 1013 772 1014
rect 822 1013 828 1014
rect 831 1015 837 1016
rect 732 1011 733 1012
rect 727 1010 733 1011
rect 727 1007 733 1008
rect 727 1006 728 1007
rect 704 1004 728 1006
rect 679 1002 685 1003
rect 727 1003 728 1004
rect 732 1003 733 1007
rect 752 1006 754 1012
rect 831 1011 832 1015
rect 836 1014 837 1015
rect 878 1014 879 1018
rect 883 1014 884 1018
rect 934 1018 940 1019
rect 836 1012 862 1014
rect 878 1013 884 1014
rect 887 1015 893 1016
rect 836 1011 837 1012
rect 831 1010 837 1011
rect 775 1007 781 1008
rect 775 1006 776 1007
rect 752 1004 776 1006
rect 727 1002 733 1003
rect 775 1003 776 1004
rect 780 1003 781 1007
rect 775 1002 781 1003
rect 831 1007 840 1008
rect 831 1003 832 1007
rect 839 1003 840 1007
rect 831 1002 840 1003
rect 860 1002 862 1012
rect 887 1011 888 1015
rect 892 1014 893 1015
rect 934 1014 935 1018
rect 939 1014 940 1018
rect 990 1018 996 1019
rect 892 1011 894 1014
rect 934 1013 940 1014
rect 943 1015 949 1016
rect 887 1010 894 1011
rect 943 1011 944 1015
rect 948 1011 949 1015
rect 990 1014 991 1018
rect 995 1014 996 1018
rect 999 1015 1000 1019
rect 1007 1015 1008 1019
rect 999 1014 1008 1015
rect 1046 1018 1052 1019
rect 1046 1014 1047 1018
rect 1051 1014 1052 1018
rect 1102 1018 1108 1019
rect 990 1013 996 1014
rect 1046 1013 1052 1014
rect 1055 1015 1061 1016
rect 943 1010 949 1011
rect 1055 1011 1056 1015
rect 1060 1011 1061 1015
rect 1102 1014 1103 1018
rect 1107 1014 1108 1018
rect 1158 1018 1164 1019
rect 1102 1013 1108 1014
rect 1111 1015 1117 1016
rect 1055 1010 1061 1011
rect 1111 1011 1112 1015
rect 1116 1011 1117 1015
rect 1158 1014 1159 1018
rect 1163 1014 1164 1018
rect 1214 1018 1220 1019
rect 1158 1013 1164 1014
rect 1167 1015 1173 1016
rect 1111 1010 1117 1011
rect 1167 1011 1168 1015
rect 1172 1014 1173 1015
rect 1214 1014 1215 1018
rect 1219 1014 1220 1018
rect 1270 1018 1276 1019
rect 1172 1012 1211 1014
rect 1214 1013 1220 1014
rect 1223 1015 1229 1016
rect 1172 1011 1173 1012
rect 1167 1010 1173 1011
rect 193 1000 219 1002
rect 228 1000 243 1002
rect 257 1000 274 1002
rect 292 1000 315 1002
rect 332 1000 355 1002
rect 464 1000 490 1002
rect 513 1000 538 1002
rect 860 1000 890 1002
rect 191 999 197 1000
rect 110 995 116 996
rect 110 991 111 995
rect 115 991 116 995
rect 191 995 192 999
rect 196 995 197 999
rect 228 998 230 1000
rect 217 996 230 998
rect 191 994 197 995
rect 215 995 221 996
rect 110 990 116 991
rect 158 992 164 993
rect 158 988 159 992
rect 163 988 164 992
rect 158 987 164 988
rect 182 992 188 993
rect 182 988 183 992
rect 187 988 188 992
rect 182 987 188 988
rect 206 992 212 993
rect 206 988 207 992
rect 211 988 212 992
rect 215 991 216 995
rect 220 991 221 995
rect 239 995 245 996
rect 215 990 221 991
rect 230 992 236 993
rect 206 987 212 988
rect 230 988 231 992
rect 235 988 236 992
rect 239 991 240 995
rect 244 994 245 995
rect 257 994 259 1000
rect 244 992 259 994
rect 271 995 277 996
rect 262 992 268 993
rect 244 991 245 992
rect 239 990 245 991
rect 230 987 236 988
rect 262 988 263 992
rect 267 988 268 992
rect 271 991 272 995
rect 276 994 277 995
rect 292 994 294 1000
rect 276 992 294 994
rect 311 995 317 996
rect 302 992 308 993
rect 276 991 277 992
rect 271 990 277 991
rect 262 987 268 988
rect 302 988 303 992
rect 307 988 308 992
rect 311 991 312 995
rect 316 994 317 995
rect 332 994 334 1000
rect 439 999 445 1000
rect 316 992 334 994
rect 351 995 360 996
rect 342 992 348 993
rect 316 991 317 992
rect 311 990 317 991
rect 302 987 308 988
rect 342 988 343 992
rect 347 988 348 992
rect 351 991 352 995
rect 359 991 360 995
rect 439 995 440 999
rect 444 998 445 999
rect 464 998 466 1000
rect 444 996 466 998
rect 444 995 445 996
rect 439 994 445 995
rect 487 995 493 996
rect 351 990 360 991
rect 382 992 388 993
rect 342 987 348 988
rect 382 988 383 992
rect 387 988 388 992
rect 382 987 388 988
rect 430 992 436 993
rect 430 988 431 992
rect 435 988 436 992
rect 430 987 436 988
rect 478 992 484 993
rect 478 988 479 992
rect 483 988 484 992
rect 487 991 488 995
rect 492 994 493 995
rect 513 994 515 1000
rect 492 992 515 994
rect 535 995 544 996
rect 526 992 532 993
rect 492 991 493 992
rect 487 990 493 991
rect 478 987 484 988
rect 526 988 527 992
rect 531 988 532 992
rect 535 991 536 995
rect 543 991 544 995
rect 535 990 544 991
rect 574 992 580 993
rect 526 987 532 988
rect 574 988 575 992
rect 579 988 580 992
rect 574 987 580 988
rect 622 992 628 993
rect 670 992 676 993
rect 622 988 623 992
rect 627 988 628 992
rect 622 987 628 988
rect 631 991 637 992
rect 631 987 632 991
rect 636 990 637 991
rect 662 991 668 992
rect 662 990 663 991
rect 636 988 663 990
rect 636 987 637 988
rect 631 986 637 987
rect 662 987 663 988
rect 667 987 668 991
rect 670 988 671 992
rect 675 988 676 992
rect 670 987 676 988
rect 718 992 724 993
rect 718 988 719 992
rect 723 988 724 992
rect 718 987 724 988
rect 766 992 772 993
rect 766 988 767 992
rect 771 988 772 992
rect 766 987 772 988
rect 822 992 828 993
rect 822 988 823 992
rect 827 988 828 992
rect 822 987 828 988
rect 878 992 884 993
rect 888 992 890 1000
rect 892 998 894 1010
rect 898 1007 904 1008
rect 898 1003 899 1007
rect 903 1006 904 1007
rect 944 1006 946 1010
rect 903 1004 946 1006
rect 999 1007 1005 1008
rect 903 1003 904 1004
rect 898 1002 904 1003
rect 999 1003 1000 1007
rect 1004 1006 1005 1007
rect 1056 1006 1058 1010
rect 1004 1004 1058 1006
rect 1004 1003 1005 1004
rect 999 1002 1005 1003
rect 1112 1002 1114 1010
rect 1167 1007 1173 1008
rect 1167 1003 1168 1007
rect 1172 1006 1173 1007
rect 1186 1007 1192 1008
rect 1186 1006 1187 1007
rect 1172 1004 1187 1006
rect 1172 1003 1173 1004
rect 1167 1002 1173 1003
rect 1186 1003 1187 1004
rect 1191 1003 1192 1007
rect 1209 1006 1211 1012
rect 1223 1011 1224 1015
rect 1228 1014 1229 1015
rect 1270 1014 1271 1018
rect 1275 1014 1276 1018
rect 1326 1018 1332 1019
rect 1228 1012 1254 1014
rect 1270 1013 1276 1014
rect 1279 1015 1285 1016
rect 1228 1011 1229 1012
rect 1223 1010 1229 1011
rect 1223 1007 1229 1008
rect 1223 1006 1224 1007
rect 1209 1004 1224 1006
rect 1186 1002 1192 1003
rect 1223 1003 1224 1004
rect 1228 1003 1229 1007
rect 1223 1002 1229 1003
rect 1252 1002 1254 1012
rect 1279 1011 1280 1015
rect 1284 1011 1285 1015
rect 1326 1014 1327 1018
rect 1331 1014 1332 1018
rect 1382 1018 1388 1019
rect 1326 1013 1332 1014
rect 1335 1015 1341 1016
rect 1279 1010 1285 1011
rect 1335 1011 1336 1015
rect 1340 1014 1341 1015
rect 1346 1015 1352 1016
rect 1346 1014 1347 1015
rect 1340 1012 1347 1014
rect 1340 1011 1341 1012
rect 1335 1010 1341 1011
rect 1346 1011 1347 1012
rect 1351 1011 1352 1015
rect 1382 1014 1383 1018
rect 1387 1014 1388 1018
rect 1391 1015 1392 1019
rect 1399 1015 1400 1019
rect 1391 1014 1400 1015
rect 1414 1018 1420 1019
rect 1414 1014 1415 1018
rect 1419 1014 1420 1018
rect 1382 1013 1388 1014
rect 1414 1013 1420 1014
rect 1423 1015 1429 1016
rect 1346 1010 1352 1011
rect 1423 1011 1424 1015
rect 1428 1011 1429 1015
rect 1423 1010 1429 1011
rect 1446 1013 1452 1014
rect 1281 1006 1283 1010
rect 1335 1007 1341 1008
rect 1335 1006 1336 1007
rect 1281 1004 1336 1006
rect 1335 1003 1336 1004
rect 1340 1003 1341 1007
rect 1335 1002 1341 1003
rect 1391 1007 1397 1008
rect 1391 1003 1392 1007
rect 1396 1006 1397 1007
rect 1425 1006 1427 1010
rect 1446 1009 1447 1013
rect 1451 1009 1452 1013
rect 1446 1008 1452 1009
rect 1396 1004 1427 1006
rect 1396 1003 1397 1004
rect 1391 1002 1397 1003
rect 916 1000 946 1002
rect 1084 1000 1114 1002
rect 1252 1000 1283 1002
rect 916 998 918 1000
rect 892 996 918 998
rect 943 999 949 1000
rect 943 995 944 999
rect 948 995 949 999
rect 943 994 949 995
rect 1055 999 1061 1000
rect 1055 995 1056 999
rect 1060 998 1061 999
rect 1084 998 1086 1000
rect 1060 996 1086 998
rect 1279 999 1285 1000
rect 1060 995 1061 996
rect 1055 994 1061 995
rect 1279 995 1280 999
rect 1284 995 1285 999
rect 1279 994 1285 995
rect 1446 995 1452 996
rect 934 992 940 993
rect 878 988 879 992
rect 883 988 884 992
rect 878 987 884 988
rect 887 991 893 992
rect 887 987 888 991
rect 892 987 893 991
rect 934 988 935 992
rect 939 988 940 992
rect 934 987 940 988
rect 990 992 996 993
rect 990 988 991 992
rect 995 988 996 992
rect 990 987 996 988
rect 1046 992 1052 993
rect 1046 988 1047 992
rect 1051 988 1052 992
rect 1046 987 1052 988
rect 1102 992 1108 993
rect 1158 992 1164 993
rect 1102 988 1103 992
rect 1107 988 1108 992
rect 1102 987 1108 988
rect 1111 991 1120 992
rect 1111 987 1112 991
rect 1119 987 1120 991
rect 1158 988 1159 992
rect 1163 988 1164 992
rect 1158 987 1164 988
rect 1214 992 1220 993
rect 1214 988 1215 992
rect 1219 988 1220 992
rect 1214 987 1220 988
rect 1270 992 1276 993
rect 1270 988 1271 992
rect 1275 988 1276 992
rect 1270 987 1276 988
rect 1326 992 1332 993
rect 1326 988 1327 992
rect 1331 988 1332 992
rect 1326 987 1332 988
rect 1382 992 1388 993
rect 1382 988 1383 992
rect 1387 988 1388 992
rect 1382 987 1388 988
rect 1414 992 1420 993
rect 1414 988 1415 992
rect 1419 988 1420 992
rect 1414 987 1420 988
rect 1423 991 1432 992
rect 1423 987 1424 991
rect 1431 987 1432 991
rect 1446 991 1447 995
rect 1451 991 1452 995
rect 1446 990 1452 991
rect 662 986 668 987
rect 887 986 893 987
rect 1111 986 1120 987
rect 1423 986 1432 987
rect 206 980 212 981
rect 110 977 116 978
rect 110 973 111 977
rect 115 973 116 977
rect 206 976 207 980
rect 211 976 212 980
rect 206 975 212 976
rect 230 980 236 981
rect 230 976 231 980
rect 235 976 236 980
rect 230 975 236 976
rect 254 980 260 981
rect 254 976 255 980
rect 259 976 260 980
rect 254 975 260 976
rect 286 980 292 981
rect 286 976 287 980
rect 291 976 292 980
rect 286 975 292 976
rect 326 980 332 981
rect 326 976 327 980
rect 331 976 332 980
rect 326 975 332 976
rect 374 980 380 981
rect 374 976 375 980
rect 379 976 380 980
rect 374 975 380 976
rect 422 980 428 981
rect 422 976 423 980
rect 427 976 428 980
rect 422 975 428 976
rect 470 980 476 981
rect 470 976 471 980
rect 475 976 476 980
rect 470 975 476 976
rect 518 980 524 981
rect 518 976 519 980
rect 523 976 524 980
rect 518 975 524 976
rect 566 980 572 981
rect 566 976 567 980
rect 571 976 572 980
rect 566 975 572 976
rect 622 980 628 981
rect 622 976 623 980
rect 627 976 628 980
rect 622 975 628 976
rect 678 980 684 981
rect 678 976 679 980
rect 683 976 684 980
rect 678 975 684 976
rect 726 980 732 981
rect 726 976 727 980
rect 731 976 732 980
rect 726 975 732 976
rect 774 980 780 981
rect 774 976 775 980
rect 779 976 780 980
rect 774 975 780 976
rect 830 980 836 981
rect 830 976 831 980
rect 835 976 836 980
rect 830 975 836 976
rect 886 980 892 981
rect 942 980 948 981
rect 886 976 887 980
rect 891 976 892 980
rect 886 975 892 976
rect 895 979 904 980
rect 895 975 896 979
rect 903 975 904 979
rect 942 976 943 980
rect 947 976 948 980
rect 942 975 948 976
rect 998 980 1004 981
rect 998 976 999 980
rect 1003 976 1004 980
rect 998 975 1004 976
rect 1046 980 1052 981
rect 1046 976 1047 980
rect 1051 976 1052 980
rect 1046 975 1052 976
rect 1094 980 1100 981
rect 1094 976 1095 980
rect 1099 976 1100 980
rect 1094 975 1100 976
rect 1142 980 1148 981
rect 1142 976 1143 980
rect 1147 976 1148 980
rect 1142 975 1148 976
rect 1190 980 1196 981
rect 1190 976 1191 980
rect 1195 976 1196 980
rect 1190 975 1196 976
rect 1238 980 1244 981
rect 1238 976 1239 980
rect 1243 976 1244 980
rect 1238 975 1244 976
rect 1286 980 1292 981
rect 1286 976 1287 980
rect 1291 976 1292 980
rect 1286 975 1292 976
rect 1334 980 1340 981
rect 1334 976 1335 980
rect 1339 976 1340 980
rect 1334 975 1340 976
rect 1382 980 1388 981
rect 1382 976 1383 980
rect 1387 976 1388 980
rect 1382 975 1388 976
rect 1414 980 1420 981
rect 1414 976 1415 980
rect 1419 976 1420 980
rect 1414 975 1420 976
rect 1446 977 1452 978
rect 895 974 904 975
rect 110 972 116 973
rect 1446 973 1447 977
rect 1451 973 1452 977
rect 1446 972 1452 973
rect 215 971 221 972
rect 215 967 216 971
rect 220 970 221 971
rect 242 971 248 972
rect 242 970 243 971
rect 220 968 243 970
rect 220 967 221 968
rect 215 966 221 967
rect 242 967 243 968
rect 247 967 248 971
rect 266 971 272 972
rect 266 970 267 971
rect 242 966 248 967
rect 257 968 267 970
rect 239 963 245 964
rect 110 959 116 960
rect 110 955 111 959
rect 115 955 116 959
rect 239 959 240 963
rect 244 962 245 963
rect 257 962 259 968
rect 266 967 267 968
rect 271 967 272 971
rect 266 966 272 967
rect 295 971 301 972
rect 295 967 296 971
rect 300 970 301 971
rect 338 971 344 972
rect 338 970 339 971
rect 300 968 339 970
rect 300 967 301 968
rect 295 966 301 967
rect 338 967 339 968
rect 343 967 344 971
rect 338 966 344 967
rect 351 971 357 972
rect 351 967 352 971
rect 356 970 357 971
rect 383 971 389 972
rect 383 970 384 971
rect 356 968 384 970
rect 356 967 357 968
rect 351 966 357 967
rect 383 967 384 968
rect 388 967 389 971
rect 383 966 389 967
rect 410 971 416 972
rect 410 967 411 971
rect 415 970 416 971
rect 431 971 437 972
rect 431 970 432 971
rect 415 968 432 970
rect 415 967 416 968
rect 410 966 416 967
rect 431 967 432 968
rect 436 967 437 971
rect 431 966 437 967
rect 575 971 581 972
rect 575 967 576 971
rect 580 970 581 971
rect 738 971 744 972
rect 738 970 739 971
rect 580 968 739 970
rect 580 967 581 968
rect 575 966 581 967
rect 738 967 739 968
rect 743 967 744 971
rect 738 966 744 967
rect 783 971 789 972
rect 783 967 784 971
rect 788 970 789 971
rect 842 971 848 972
rect 842 970 843 971
rect 788 968 843 970
rect 788 967 789 968
rect 783 966 789 967
rect 842 967 843 968
rect 847 967 848 971
rect 842 966 848 967
rect 1151 971 1157 972
rect 1151 967 1152 971
rect 1156 970 1157 971
rect 1346 971 1352 972
rect 1346 970 1347 971
rect 1156 968 1347 970
rect 1156 967 1157 968
rect 1151 966 1157 967
rect 1346 967 1347 968
rect 1351 967 1352 971
rect 1346 966 1352 967
rect 244 960 259 962
rect 263 963 269 964
rect 244 959 245 960
rect 239 958 245 959
rect 263 959 264 963
rect 268 962 269 963
rect 335 963 341 964
rect 268 960 298 962
rect 268 959 269 960
rect 263 958 269 959
rect 296 956 298 960
rect 335 959 336 963
rect 340 962 341 963
rect 479 963 485 964
rect 479 962 480 963
rect 340 960 362 962
rect 340 959 341 960
rect 335 958 341 959
rect 215 955 224 956
rect 239 955 248 956
rect 263 955 272 956
rect 295 955 301 956
rect 335 955 344 956
rect 110 954 116 955
rect 206 954 212 955
rect 206 950 207 954
rect 211 950 212 954
rect 215 951 216 955
rect 223 951 224 955
rect 215 950 224 951
rect 230 954 236 955
rect 230 950 231 954
rect 235 950 236 954
rect 239 951 240 955
rect 247 951 248 955
rect 239 950 248 951
rect 254 954 260 955
rect 254 950 255 954
rect 259 950 260 954
rect 263 951 264 955
rect 271 951 272 955
rect 263 950 272 951
rect 286 954 292 955
rect 286 950 287 954
rect 291 950 292 954
rect 295 951 296 955
rect 300 951 301 955
rect 295 950 301 951
rect 326 954 332 955
rect 326 950 327 954
rect 331 950 332 954
rect 335 951 336 955
rect 343 951 344 955
rect 335 950 344 951
rect 206 949 212 950
rect 230 949 236 950
rect 254 949 260 950
rect 286 949 292 950
rect 326 949 332 950
rect 274 947 280 948
rect 274 943 275 947
rect 279 946 280 947
rect 302 947 308 948
rect 279 944 298 946
rect 279 943 280 944
rect 274 942 280 943
rect 296 940 298 944
rect 302 943 303 947
rect 307 946 308 947
rect 351 947 357 948
rect 351 946 352 947
rect 307 944 352 946
rect 307 943 308 944
rect 302 942 308 943
rect 351 943 352 944
rect 356 943 357 947
rect 360 946 362 960
rect 456 960 480 962
rect 431 955 437 956
rect 374 954 380 955
rect 374 950 375 954
rect 379 950 380 954
rect 422 954 428 955
rect 374 949 380 950
rect 383 951 389 952
rect 383 947 384 951
rect 388 947 389 951
rect 422 950 423 954
rect 427 950 428 954
rect 431 951 432 955
rect 436 954 437 955
rect 456 954 458 960
rect 479 959 480 960
rect 484 959 485 963
rect 527 963 533 964
rect 527 962 528 963
rect 479 958 485 959
rect 504 960 528 962
rect 479 955 485 956
rect 436 952 458 954
rect 470 954 476 955
rect 436 951 437 952
rect 431 950 437 951
rect 470 950 471 954
rect 475 950 476 954
rect 479 951 480 955
rect 484 954 485 955
rect 504 954 506 960
rect 527 959 528 960
rect 532 959 533 963
rect 631 963 637 964
rect 631 962 632 963
rect 527 958 533 959
rect 604 960 632 962
rect 575 955 581 956
rect 484 952 506 954
rect 518 954 524 955
rect 484 951 485 952
rect 479 950 485 951
rect 518 950 519 954
rect 523 950 524 954
rect 566 954 572 955
rect 422 949 428 950
rect 470 949 476 950
rect 518 949 524 950
rect 527 951 536 952
rect 383 946 389 947
rect 527 947 528 951
rect 535 947 536 951
rect 566 950 567 954
rect 571 950 572 954
rect 575 951 576 955
rect 580 954 581 955
rect 604 954 606 960
rect 631 959 632 960
rect 636 959 637 963
rect 687 963 693 964
rect 687 962 688 963
rect 631 958 637 959
rect 656 960 688 962
rect 631 955 637 956
rect 580 952 606 954
rect 622 954 628 955
rect 580 951 581 952
rect 575 950 581 951
rect 622 950 623 954
rect 627 950 628 954
rect 631 951 632 955
rect 636 954 637 955
rect 656 954 658 960
rect 687 959 688 960
rect 692 959 693 963
rect 735 963 741 964
rect 735 962 736 963
rect 687 958 693 959
rect 712 960 736 962
rect 687 955 693 956
rect 636 952 658 954
rect 678 954 684 955
rect 636 951 637 952
rect 631 950 637 951
rect 678 950 679 954
rect 683 950 684 954
rect 687 951 688 955
rect 692 954 693 955
rect 712 954 714 960
rect 735 959 736 960
rect 740 959 741 963
rect 735 958 741 959
rect 839 963 845 964
rect 839 959 840 963
rect 844 962 845 963
rect 930 963 936 964
rect 844 960 898 962
rect 844 959 845 960
rect 839 958 845 959
rect 896 956 898 960
rect 930 959 931 963
rect 935 962 936 963
rect 951 963 957 964
rect 951 962 952 963
rect 935 960 952 962
rect 935 959 936 960
rect 930 958 936 959
rect 951 959 952 960
rect 956 959 957 963
rect 1007 963 1013 964
rect 1007 962 1008 963
rect 951 958 957 959
rect 980 960 1008 962
rect 839 955 848 956
rect 895 955 901 956
rect 951 955 957 956
rect 692 952 714 954
rect 726 954 732 955
rect 692 951 693 952
rect 687 950 693 951
rect 726 950 727 954
rect 731 950 732 954
rect 774 954 780 955
rect 566 949 572 950
rect 622 949 628 950
rect 678 949 684 950
rect 726 949 732 950
rect 735 951 741 952
rect 527 946 536 947
rect 662 947 668 948
rect 360 944 386 946
rect 351 942 357 943
rect 662 943 663 947
rect 667 946 668 947
rect 735 947 736 951
rect 740 947 741 951
rect 774 950 775 954
rect 779 950 780 954
rect 830 954 836 955
rect 774 949 780 950
rect 783 951 789 952
rect 735 946 741 947
rect 783 947 784 951
rect 788 950 789 951
rect 794 951 800 952
rect 794 950 795 951
rect 788 948 795 950
rect 788 947 789 948
rect 783 946 789 947
rect 794 947 795 948
rect 799 947 800 951
rect 830 950 831 954
rect 835 950 836 954
rect 839 951 840 955
rect 847 951 848 955
rect 839 950 848 951
rect 886 954 892 955
rect 886 950 887 954
rect 891 950 892 954
rect 895 951 896 955
rect 900 951 901 955
rect 895 950 901 951
rect 942 954 948 955
rect 942 950 943 954
rect 947 950 948 954
rect 951 951 952 955
rect 956 954 957 955
rect 980 954 982 960
rect 1007 959 1008 960
rect 1012 959 1013 963
rect 1055 963 1061 964
rect 1055 962 1056 963
rect 1007 958 1013 959
rect 1032 960 1056 962
rect 1007 955 1013 956
rect 956 952 982 954
rect 998 954 1004 955
rect 956 951 957 952
rect 951 950 957 951
rect 998 950 999 954
rect 1003 950 1004 954
rect 1007 951 1008 955
rect 1012 954 1013 955
rect 1032 954 1034 960
rect 1055 959 1056 960
rect 1060 959 1061 963
rect 1103 963 1109 964
rect 1103 962 1104 963
rect 1055 958 1061 959
rect 1080 960 1104 962
rect 1055 955 1061 956
rect 1012 952 1034 954
rect 1046 954 1052 955
rect 1012 951 1013 952
rect 1007 950 1013 951
rect 1046 950 1047 954
rect 1051 950 1052 954
rect 1055 951 1056 955
rect 1060 954 1061 955
rect 1080 954 1082 960
rect 1103 959 1104 960
rect 1108 959 1109 963
rect 1199 963 1205 964
rect 1199 962 1200 963
rect 1103 958 1109 959
rect 1159 960 1200 962
rect 1103 955 1109 956
rect 1060 952 1082 954
rect 1094 954 1100 955
rect 1060 951 1061 952
rect 1055 950 1061 951
rect 1094 950 1095 954
rect 1099 950 1100 954
rect 1103 951 1104 955
rect 1108 954 1109 955
rect 1114 955 1120 956
rect 1151 955 1157 956
rect 1114 954 1115 955
rect 1108 952 1115 954
rect 1108 951 1109 952
rect 1103 950 1109 951
rect 1114 951 1115 952
rect 1119 951 1120 955
rect 1114 950 1120 951
rect 1142 954 1148 955
rect 1142 950 1143 954
rect 1147 950 1148 954
rect 1151 951 1152 955
rect 1156 954 1157 955
rect 1159 954 1161 960
rect 1199 959 1200 960
rect 1204 959 1205 963
rect 1247 963 1253 964
rect 1247 962 1248 963
rect 1199 958 1205 959
rect 1224 960 1248 962
rect 1199 955 1205 956
rect 1156 952 1161 954
rect 1190 954 1196 955
rect 1156 951 1157 952
rect 1151 950 1157 951
rect 1190 950 1191 954
rect 1195 950 1196 954
rect 1199 951 1200 955
rect 1204 954 1205 955
rect 1224 954 1226 960
rect 1247 959 1248 960
rect 1252 959 1253 963
rect 1295 963 1301 964
rect 1295 962 1296 963
rect 1247 958 1253 959
rect 1272 960 1296 962
rect 1247 955 1253 956
rect 1204 952 1226 954
rect 1238 954 1244 955
rect 1204 951 1205 952
rect 1199 950 1205 951
rect 1238 950 1239 954
rect 1243 950 1244 954
rect 1247 951 1248 955
rect 1252 954 1253 955
rect 1272 954 1274 960
rect 1295 959 1296 960
rect 1300 959 1301 963
rect 1343 963 1349 964
rect 1343 962 1344 963
rect 1295 958 1301 959
rect 1321 960 1344 962
rect 1295 955 1301 956
rect 1252 952 1274 954
rect 1286 954 1292 955
rect 1252 951 1253 952
rect 1247 950 1253 951
rect 1286 950 1287 954
rect 1291 950 1292 954
rect 1295 951 1296 955
rect 1300 954 1301 955
rect 1321 954 1323 960
rect 1343 959 1344 960
rect 1348 959 1349 963
rect 1391 963 1397 964
rect 1391 962 1392 963
rect 1343 958 1349 959
rect 1368 960 1392 962
rect 1343 955 1349 956
rect 1300 952 1323 954
rect 1334 954 1340 955
rect 1300 951 1301 952
rect 1295 950 1301 951
rect 1334 950 1335 954
rect 1339 950 1340 954
rect 1343 951 1344 955
rect 1348 954 1349 955
rect 1368 954 1370 960
rect 1391 959 1392 960
rect 1396 959 1397 963
rect 1391 958 1397 959
rect 1423 963 1429 964
rect 1423 959 1424 963
rect 1428 962 1429 963
rect 1431 963 1437 964
rect 1431 962 1432 963
rect 1428 960 1432 962
rect 1428 959 1429 960
rect 1423 958 1429 959
rect 1431 959 1432 960
rect 1436 959 1437 963
rect 1431 958 1437 959
rect 1446 959 1452 960
rect 1423 955 1432 956
rect 1348 952 1370 954
rect 1382 954 1388 955
rect 1348 951 1349 952
rect 1343 950 1349 951
rect 1382 950 1383 954
rect 1387 950 1388 954
rect 1414 954 1420 955
rect 830 949 836 950
rect 886 949 892 950
rect 942 949 948 950
rect 998 949 1004 950
rect 1046 949 1052 950
rect 1094 949 1100 950
rect 1142 949 1148 950
rect 1190 949 1196 950
rect 1238 949 1244 950
rect 1286 949 1292 950
rect 1334 949 1340 950
rect 1382 949 1388 950
rect 1391 951 1397 952
rect 794 946 800 947
rect 1130 947 1136 948
rect 667 944 681 946
rect 667 943 668 944
rect 662 942 668 943
rect 679 942 681 944
rect 696 944 738 946
rect 696 942 698 944
rect 1130 943 1131 947
rect 1135 946 1136 947
rect 1391 947 1392 951
rect 1396 947 1397 951
rect 1414 950 1415 954
rect 1419 950 1420 954
rect 1423 951 1424 955
rect 1431 951 1432 955
rect 1446 955 1447 959
rect 1451 955 1452 959
rect 1446 954 1452 955
rect 1423 950 1432 951
rect 1414 949 1420 950
rect 1391 946 1397 947
rect 1135 944 1395 946
rect 1135 943 1136 944
rect 1130 942 1136 943
rect 679 940 698 942
rect 295 939 301 940
rect 735 939 744 940
rect 927 939 936 940
rect 1423 939 1429 940
rect 214 938 220 939
rect 214 934 215 938
rect 219 934 220 938
rect 238 938 244 939
rect 110 933 116 934
rect 214 933 220 934
rect 223 935 232 936
rect 110 929 111 933
rect 115 929 116 933
rect 223 931 224 935
rect 231 931 232 935
rect 238 934 239 938
rect 243 934 244 938
rect 262 938 268 939
rect 238 933 244 934
rect 247 935 253 936
rect 223 930 232 931
rect 247 931 248 935
rect 252 931 253 935
rect 262 934 263 938
rect 267 934 268 938
rect 286 938 292 939
rect 262 933 268 934
rect 271 935 277 936
rect 247 930 253 931
rect 271 931 272 935
rect 276 931 277 935
rect 286 934 287 938
rect 291 934 292 938
rect 295 935 296 939
rect 300 935 301 939
rect 295 934 301 935
rect 318 938 324 939
rect 318 934 319 938
rect 323 934 324 938
rect 350 938 356 939
rect 286 933 292 934
rect 318 933 324 934
rect 327 935 333 936
rect 271 930 277 931
rect 327 931 328 935
rect 332 931 333 935
rect 350 934 351 938
rect 355 934 356 938
rect 390 938 396 939
rect 350 933 356 934
rect 359 935 365 936
rect 327 930 333 931
rect 359 931 360 935
rect 364 931 365 935
rect 390 934 391 938
rect 395 934 396 938
rect 430 938 436 939
rect 390 933 396 934
rect 399 935 405 936
rect 359 930 365 931
rect 399 931 400 935
rect 404 931 405 935
rect 430 934 431 938
rect 435 934 436 938
rect 470 938 476 939
rect 430 933 436 934
rect 439 935 445 936
rect 399 930 405 931
rect 439 931 440 935
rect 444 934 445 935
rect 470 934 471 938
rect 475 934 476 938
rect 518 938 524 939
rect 444 932 462 934
rect 470 933 476 934
rect 479 935 485 936
rect 444 931 445 932
rect 439 930 445 931
rect 110 928 116 929
rect 223 927 229 928
rect 223 923 224 927
rect 228 926 229 927
rect 248 926 250 930
rect 228 924 250 926
rect 228 923 229 924
rect 223 922 229 923
rect 272 922 274 930
rect 260 920 274 922
rect 295 923 301 924
rect 247 919 253 920
rect 110 915 116 916
rect 110 911 111 915
rect 115 911 116 915
rect 247 915 248 919
rect 252 918 253 919
rect 260 918 262 920
rect 295 919 296 923
rect 300 922 301 923
rect 328 922 330 930
rect 360 922 362 930
rect 400 922 402 930
rect 439 927 448 928
rect 439 923 440 927
rect 447 923 448 927
rect 460 926 462 932
rect 479 931 480 935
rect 484 934 485 935
rect 506 935 512 936
rect 506 934 507 935
rect 484 932 507 934
rect 484 931 485 932
rect 479 930 485 931
rect 506 931 507 932
rect 511 931 512 935
rect 518 934 519 938
rect 523 934 524 938
rect 566 938 572 939
rect 518 933 524 934
rect 527 935 533 936
rect 506 930 512 931
rect 527 931 528 935
rect 532 934 533 935
rect 538 935 544 936
rect 538 934 539 935
rect 532 932 539 934
rect 532 931 533 932
rect 527 930 533 931
rect 538 931 539 932
rect 543 931 544 935
rect 566 934 567 938
rect 571 934 572 938
rect 614 938 620 939
rect 566 933 572 934
rect 575 935 581 936
rect 538 930 544 931
rect 575 931 576 935
rect 580 934 581 935
rect 614 934 615 938
rect 619 934 620 938
rect 670 938 676 939
rect 580 932 602 934
rect 614 933 620 934
rect 623 935 629 936
rect 580 931 581 932
rect 575 930 581 931
rect 479 927 485 928
rect 479 926 480 927
rect 460 924 480 926
rect 439 922 448 923
rect 479 923 480 924
rect 484 923 485 927
rect 479 922 485 923
rect 527 927 536 928
rect 527 923 528 927
rect 535 923 536 927
rect 600 926 602 932
rect 623 931 624 935
rect 628 934 629 935
rect 670 934 671 938
rect 675 934 676 938
rect 726 938 732 939
rect 628 932 654 934
rect 670 933 676 934
rect 679 935 685 936
rect 628 931 629 932
rect 623 930 629 931
rect 623 927 629 928
rect 623 926 624 927
rect 600 924 624 926
rect 527 922 536 923
rect 623 923 624 924
rect 628 923 629 927
rect 652 926 654 932
rect 679 931 680 935
rect 684 934 685 935
rect 726 934 727 938
rect 731 934 732 938
rect 735 935 736 939
rect 743 935 744 939
rect 735 934 744 935
rect 782 938 788 939
rect 782 934 783 938
rect 787 934 788 938
rect 846 938 852 939
rect 684 932 710 934
rect 726 933 732 934
rect 782 933 788 934
rect 791 935 797 936
rect 684 931 685 932
rect 679 930 685 931
rect 679 927 685 928
rect 679 926 680 927
rect 652 924 680 926
rect 623 922 629 923
rect 679 923 680 924
rect 684 923 685 927
rect 708 926 710 932
rect 791 931 792 935
rect 796 934 797 935
rect 846 934 847 938
rect 851 934 852 938
rect 918 938 924 939
rect 796 932 827 934
rect 846 933 852 934
rect 855 935 864 936
rect 796 931 797 932
rect 791 930 797 931
rect 735 927 741 928
rect 735 926 736 927
rect 708 924 736 926
rect 679 922 685 923
rect 735 923 736 924
rect 740 923 741 927
rect 735 922 741 923
rect 791 927 800 928
rect 791 923 792 927
rect 799 923 800 927
rect 825 926 827 932
rect 855 931 856 935
rect 863 931 864 935
rect 918 934 919 938
rect 923 934 924 938
rect 927 935 928 939
rect 935 935 936 939
rect 927 934 936 935
rect 990 938 996 939
rect 990 934 991 938
rect 995 934 996 938
rect 1054 938 1060 939
rect 918 933 924 934
rect 990 933 996 934
rect 999 935 1008 936
rect 855 930 864 931
rect 999 931 1000 935
rect 1007 931 1008 935
rect 1054 934 1055 938
rect 1059 934 1060 938
rect 1118 938 1124 939
rect 1054 933 1060 934
rect 1063 935 1069 936
rect 999 930 1008 931
rect 1063 931 1064 935
rect 1068 931 1069 935
rect 1118 934 1119 938
rect 1123 934 1124 938
rect 1174 938 1180 939
rect 1118 933 1124 934
rect 1127 935 1133 936
rect 1063 930 1069 931
rect 1127 931 1128 935
rect 1132 934 1133 935
rect 1174 934 1175 938
rect 1179 934 1180 938
rect 1222 938 1228 939
rect 1132 932 1161 934
rect 1174 933 1180 934
rect 1183 935 1189 936
rect 1132 931 1133 932
rect 1127 930 1133 931
rect 855 927 861 928
rect 855 926 856 927
rect 825 924 856 926
rect 791 922 800 923
rect 855 923 856 924
rect 860 923 861 927
rect 999 927 1005 928
rect 855 922 861 923
rect 927 923 933 924
rect 300 920 330 922
rect 345 920 362 922
rect 380 920 402 922
rect 300 919 301 920
rect 295 918 301 919
rect 252 916 262 918
rect 252 915 253 916
rect 247 914 253 915
rect 271 915 280 916
rect 110 910 116 911
rect 214 912 220 913
rect 214 908 215 912
rect 219 908 220 912
rect 214 907 220 908
rect 238 912 244 913
rect 238 908 239 912
rect 243 908 244 912
rect 238 907 244 908
rect 262 912 268 913
rect 262 908 263 912
rect 267 908 268 912
rect 271 911 272 915
rect 279 911 280 915
rect 327 915 333 916
rect 271 910 280 911
rect 286 912 292 913
rect 262 907 268 908
rect 286 908 287 912
rect 291 908 292 912
rect 286 907 292 908
rect 318 912 324 913
rect 318 908 319 912
rect 323 908 324 912
rect 327 911 328 915
rect 332 914 333 915
rect 345 914 347 920
rect 332 912 347 914
rect 359 915 365 916
rect 350 912 356 913
rect 332 911 333 912
rect 327 910 333 911
rect 318 907 324 908
rect 350 908 351 912
rect 355 908 356 912
rect 359 911 360 915
rect 364 914 365 915
rect 380 914 382 920
rect 927 919 928 923
rect 932 922 933 923
rect 990 923 996 924
rect 990 922 991 923
rect 932 920 991 922
rect 932 919 933 920
rect 927 918 933 919
rect 990 919 991 920
rect 995 919 996 923
rect 999 923 1000 927
rect 1004 926 1005 927
rect 1064 926 1066 930
rect 1004 924 1066 926
rect 1127 927 1136 928
rect 1004 923 1005 924
rect 999 922 1005 923
rect 1127 923 1128 927
rect 1135 923 1136 927
rect 1159 926 1161 932
rect 1183 931 1184 935
rect 1188 934 1189 935
rect 1222 934 1223 938
rect 1227 934 1228 938
rect 1262 938 1268 939
rect 1188 932 1210 934
rect 1222 933 1228 934
rect 1231 935 1237 936
rect 1188 931 1189 932
rect 1183 930 1189 931
rect 1183 927 1189 928
rect 1183 926 1184 927
rect 1159 924 1184 926
rect 1127 922 1136 923
rect 1183 923 1184 924
rect 1188 923 1189 927
rect 1208 926 1210 932
rect 1231 931 1232 935
rect 1236 934 1237 935
rect 1262 934 1263 938
rect 1267 934 1268 938
rect 1294 938 1300 939
rect 1236 932 1259 934
rect 1262 933 1268 934
rect 1271 935 1277 936
rect 1236 931 1237 932
rect 1231 930 1237 931
rect 1231 927 1237 928
rect 1231 926 1232 927
rect 1208 924 1232 926
rect 1183 922 1189 923
rect 1231 923 1232 924
rect 1236 923 1237 927
rect 1257 926 1259 932
rect 1271 931 1272 935
rect 1276 934 1277 935
rect 1294 934 1295 938
rect 1299 934 1300 938
rect 1326 938 1332 939
rect 1276 932 1291 934
rect 1294 933 1300 934
rect 1303 935 1309 936
rect 1276 931 1277 932
rect 1271 930 1277 931
rect 1271 927 1277 928
rect 1271 926 1272 927
rect 1257 924 1272 926
rect 1231 922 1237 923
rect 1271 923 1272 924
rect 1276 923 1277 927
rect 1289 926 1291 932
rect 1303 931 1304 935
rect 1308 934 1309 935
rect 1326 934 1327 938
rect 1331 934 1332 938
rect 1358 938 1364 939
rect 1308 932 1323 934
rect 1326 933 1332 934
rect 1335 935 1341 936
rect 1308 931 1309 932
rect 1303 930 1309 931
rect 1303 927 1309 928
rect 1303 926 1304 927
rect 1289 924 1304 926
rect 1271 922 1277 923
rect 1303 923 1304 924
rect 1308 923 1309 927
rect 1303 922 1309 923
rect 1321 922 1323 932
rect 1335 931 1336 935
rect 1340 931 1341 935
rect 1358 934 1359 938
rect 1363 934 1364 938
rect 1390 938 1396 939
rect 1358 933 1364 934
rect 1367 935 1373 936
rect 1335 930 1341 931
rect 1367 931 1368 935
rect 1372 934 1373 935
rect 1375 935 1381 936
rect 1375 934 1376 935
rect 1372 932 1376 934
rect 1372 931 1373 932
rect 1367 930 1373 931
rect 1375 931 1376 932
rect 1380 931 1381 935
rect 1390 934 1391 938
rect 1395 934 1396 938
rect 1414 938 1420 939
rect 1390 933 1396 934
rect 1399 935 1405 936
rect 1375 930 1381 931
rect 1399 931 1400 935
rect 1404 931 1405 935
rect 1414 934 1415 938
rect 1419 934 1420 938
rect 1423 935 1424 939
rect 1428 938 1429 939
rect 1431 939 1437 940
rect 1431 938 1432 939
rect 1428 936 1432 938
rect 1428 935 1429 936
rect 1423 934 1429 935
rect 1431 935 1432 936
rect 1436 935 1437 939
rect 1431 934 1437 935
rect 1414 933 1420 934
rect 1446 933 1452 934
rect 1399 930 1405 931
rect 1337 926 1339 930
rect 1367 927 1373 928
rect 1367 926 1368 927
rect 1337 924 1368 926
rect 1367 923 1368 924
rect 1372 923 1373 927
rect 1401 926 1403 930
rect 1446 929 1447 933
rect 1451 929 1452 933
rect 1446 928 1452 929
rect 1423 927 1429 928
rect 1423 926 1424 927
rect 1401 924 1424 926
rect 1367 922 1373 923
rect 1423 923 1424 924
rect 1428 923 1429 927
rect 1423 922 1429 923
rect 1321 920 1339 922
rect 990 918 996 919
rect 1335 919 1341 920
rect 1335 915 1336 919
rect 1340 915 1341 919
rect 1335 914 1341 915
rect 1446 915 1452 916
rect 364 912 382 914
rect 390 912 396 913
rect 430 912 436 913
rect 364 911 365 912
rect 359 910 365 911
rect 350 907 356 908
rect 390 908 391 912
rect 395 908 396 912
rect 390 907 396 908
rect 399 911 408 912
rect 399 907 400 911
rect 407 907 408 911
rect 430 908 431 912
rect 435 908 436 912
rect 430 907 436 908
rect 470 912 476 913
rect 470 908 471 912
rect 475 908 476 912
rect 470 907 476 908
rect 518 912 524 913
rect 518 908 519 912
rect 523 908 524 912
rect 518 907 524 908
rect 566 912 572 913
rect 614 912 620 913
rect 566 908 567 912
rect 571 908 572 912
rect 566 907 572 908
rect 575 911 581 912
rect 575 907 576 911
rect 580 910 581 911
rect 606 911 612 912
rect 606 910 607 911
rect 580 908 607 910
rect 580 907 581 908
rect 399 906 408 907
rect 575 906 581 907
rect 606 907 607 908
rect 611 907 612 911
rect 614 908 615 912
rect 619 908 620 912
rect 614 907 620 908
rect 670 912 676 913
rect 670 908 671 912
rect 675 908 676 912
rect 670 907 676 908
rect 726 912 732 913
rect 726 908 727 912
rect 731 908 732 912
rect 726 907 732 908
rect 782 912 788 913
rect 782 908 783 912
rect 787 908 788 912
rect 782 907 788 908
rect 846 912 852 913
rect 846 908 847 912
rect 851 908 852 912
rect 846 907 852 908
rect 918 912 924 913
rect 918 908 919 912
rect 923 908 924 912
rect 918 907 924 908
rect 990 912 996 913
rect 990 908 991 912
rect 995 908 996 912
rect 990 907 996 908
rect 1054 912 1060 913
rect 1118 912 1124 913
rect 1054 908 1055 912
rect 1059 908 1060 912
rect 1054 907 1060 908
rect 1063 911 1072 912
rect 1063 907 1064 911
rect 1071 907 1072 911
rect 1118 908 1119 912
rect 1123 908 1124 912
rect 1118 907 1124 908
rect 1174 912 1180 913
rect 1174 908 1175 912
rect 1179 908 1180 912
rect 1174 907 1180 908
rect 1222 912 1228 913
rect 1222 908 1223 912
rect 1227 908 1228 912
rect 1222 907 1228 908
rect 1262 912 1268 913
rect 1262 908 1263 912
rect 1267 908 1268 912
rect 1262 907 1268 908
rect 1294 912 1300 913
rect 1294 908 1295 912
rect 1299 908 1300 912
rect 1294 907 1300 908
rect 1326 912 1332 913
rect 1326 908 1327 912
rect 1331 908 1332 912
rect 1326 907 1332 908
rect 1358 912 1364 913
rect 1358 908 1359 912
rect 1363 908 1364 912
rect 1358 907 1364 908
rect 1390 912 1396 913
rect 1414 912 1420 913
rect 1390 908 1391 912
rect 1395 908 1396 912
rect 1390 907 1396 908
rect 1399 911 1408 912
rect 1399 907 1400 911
rect 1407 907 1408 911
rect 1414 908 1415 912
rect 1419 908 1420 912
rect 1446 911 1447 915
rect 1451 911 1452 915
rect 1446 910 1452 911
rect 1414 907 1420 908
rect 606 906 612 907
rect 1063 906 1072 907
rect 1399 906 1408 907
rect 230 900 236 901
rect 110 897 116 898
rect 110 893 111 897
rect 115 893 116 897
rect 230 896 231 900
rect 235 896 236 900
rect 230 895 236 896
rect 254 900 260 901
rect 254 896 255 900
rect 259 896 260 900
rect 254 895 260 896
rect 278 900 284 901
rect 278 896 279 900
rect 283 896 284 900
rect 278 895 284 896
rect 302 900 308 901
rect 302 896 303 900
rect 307 896 308 900
rect 302 895 308 896
rect 326 900 332 901
rect 326 896 327 900
rect 331 896 332 900
rect 326 895 332 896
rect 358 900 364 901
rect 358 896 359 900
rect 363 896 364 900
rect 358 895 364 896
rect 390 900 396 901
rect 390 896 391 900
rect 395 896 396 900
rect 390 895 396 896
rect 422 900 428 901
rect 422 896 423 900
rect 427 896 428 900
rect 422 895 428 896
rect 454 900 460 901
rect 454 896 455 900
rect 459 896 460 900
rect 454 895 460 896
rect 494 900 500 901
rect 534 900 540 901
rect 494 896 495 900
rect 499 896 500 900
rect 494 895 500 896
rect 503 899 512 900
rect 503 895 504 899
rect 511 895 512 899
rect 534 896 535 900
rect 539 896 540 900
rect 534 895 540 896
rect 574 900 580 901
rect 574 896 575 900
rect 579 896 580 900
rect 574 895 580 896
rect 622 900 628 901
rect 622 896 623 900
rect 627 896 628 900
rect 622 895 628 896
rect 662 900 668 901
rect 662 896 663 900
rect 667 896 668 900
rect 662 895 668 896
rect 702 900 708 901
rect 702 896 703 900
rect 707 896 708 900
rect 702 895 708 896
rect 750 900 756 901
rect 750 896 751 900
rect 755 896 756 900
rect 750 895 756 896
rect 806 900 812 901
rect 862 900 868 901
rect 806 896 807 900
rect 811 896 812 900
rect 806 895 812 896
rect 815 899 821 900
rect 815 895 816 899
rect 820 898 821 899
rect 854 899 860 900
rect 854 898 855 899
rect 820 896 855 898
rect 820 895 821 896
rect 503 894 512 895
rect 815 894 821 895
rect 854 895 855 896
rect 859 895 860 899
rect 862 896 863 900
rect 867 896 868 900
rect 862 895 868 896
rect 926 900 932 901
rect 926 896 927 900
rect 931 896 932 900
rect 926 895 932 896
rect 990 900 996 901
rect 990 896 991 900
rect 995 896 996 900
rect 990 895 996 896
rect 1054 900 1060 901
rect 1054 896 1055 900
rect 1059 896 1060 900
rect 1054 895 1060 896
rect 1118 900 1124 901
rect 1118 896 1119 900
rect 1123 896 1124 900
rect 1118 895 1124 896
rect 1174 900 1180 901
rect 1174 896 1175 900
rect 1179 896 1180 900
rect 1174 895 1180 896
rect 1230 900 1236 901
rect 1230 896 1231 900
rect 1235 896 1236 900
rect 1230 895 1236 896
rect 1278 900 1284 901
rect 1278 896 1279 900
rect 1283 896 1284 900
rect 1278 895 1284 896
rect 1326 900 1332 901
rect 1326 896 1327 900
rect 1331 896 1332 900
rect 1326 895 1332 896
rect 1382 900 1388 901
rect 1382 896 1383 900
rect 1387 896 1388 900
rect 1382 895 1388 896
rect 1414 900 1420 901
rect 1414 896 1415 900
rect 1419 896 1420 900
rect 1414 895 1420 896
rect 1446 897 1452 898
rect 854 894 860 895
rect 110 892 116 893
rect 1446 893 1447 897
rect 1451 893 1452 897
rect 1446 892 1452 893
rect 431 891 437 892
rect 238 887 245 888
rect 238 883 239 887
rect 244 883 245 887
rect 431 887 432 891
rect 436 890 437 891
rect 466 891 472 892
rect 466 890 467 891
rect 436 888 467 890
rect 436 887 437 888
rect 431 886 437 887
rect 466 887 467 888
rect 471 887 472 891
rect 466 886 472 887
rect 543 891 549 892
rect 543 887 544 891
rect 548 890 549 891
rect 655 891 661 892
rect 655 890 656 891
rect 548 888 656 890
rect 548 887 549 888
rect 543 886 549 887
rect 655 887 656 888
rect 660 887 661 891
rect 655 886 661 887
rect 711 891 717 892
rect 711 887 712 891
rect 716 890 717 891
rect 762 891 768 892
rect 762 890 763 891
rect 716 888 763 890
rect 716 887 717 888
rect 711 886 717 887
rect 762 887 763 888
rect 767 887 768 891
rect 762 886 768 887
rect 1127 891 1133 892
rect 1127 887 1128 891
rect 1132 890 1133 891
rect 1186 891 1192 892
rect 1186 890 1187 891
rect 1132 888 1187 890
rect 1132 887 1133 888
rect 1127 886 1133 887
rect 1186 887 1187 888
rect 1191 887 1192 891
rect 1186 886 1192 887
rect 1239 891 1245 892
rect 1239 887 1240 891
rect 1244 890 1245 891
rect 1290 891 1296 892
rect 1290 890 1291 891
rect 1244 888 1291 890
rect 1244 887 1245 888
rect 1239 886 1245 887
rect 1290 887 1291 888
rect 1295 887 1296 891
rect 1290 886 1296 887
rect 1375 891 1381 892
rect 1375 887 1376 891
rect 1380 890 1381 891
rect 1391 891 1397 892
rect 1391 890 1392 891
rect 1380 888 1392 890
rect 1380 887 1381 888
rect 1375 886 1381 887
rect 1391 887 1392 888
rect 1396 887 1397 891
rect 1391 886 1397 887
rect 238 882 245 883
rect 263 883 269 884
rect 263 882 264 883
rect 248 880 264 882
rect 110 879 116 880
rect 110 875 111 879
rect 115 875 116 879
rect 239 875 245 876
rect 110 874 116 875
rect 230 874 236 875
rect 230 870 231 874
rect 235 870 236 874
rect 239 871 240 875
rect 244 874 245 875
rect 248 874 250 880
rect 263 879 264 880
rect 268 879 269 883
rect 287 883 293 884
rect 287 882 288 883
rect 263 878 269 879
rect 272 880 288 882
rect 263 875 269 876
rect 244 872 250 874
rect 254 874 260 875
rect 244 871 245 872
rect 239 870 245 871
rect 254 870 255 874
rect 259 870 260 874
rect 263 871 264 875
rect 268 874 269 875
rect 272 874 274 880
rect 287 879 288 880
rect 292 879 293 883
rect 311 883 317 884
rect 311 882 312 883
rect 287 878 293 879
rect 296 880 312 882
rect 287 875 293 876
rect 268 872 274 874
rect 278 874 284 875
rect 268 871 269 872
rect 263 870 269 871
rect 278 870 279 874
rect 283 870 284 874
rect 287 871 288 875
rect 292 874 293 875
rect 296 874 298 880
rect 311 879 312 880
rect 316 879 317 883
rect 335 883 341 884
rect 335 882 336 883
rect 311 878 317 879
rect 320 880 336 882
rect 311 875 317 876
rect 292 872 298 874
rect 302 874 308 875
rect 292 871 293 872
rect 287 870 293 871
rect 302 870 303 874
rect 307 870 308 874
rect 311 871 312 875
rect 316 874 317 875
rect 320 874 322 880
rect 335 879 336 880
rect 340 879 341 883
rect 367 883 373 884
rect 367 882 368 883
rect 335 878 341 879
rect 353 880 368 882
rect 335 875 341 876
rect 316 872 322 874
rect 326 874 332 875
rect 316 871 317 872
rect 311 870 317 871
rect 326 870 327 874
rect 331 870 332 874
rect 335 871 336 875
rect 340 874 341 875
rect 353 874 355 880
rect 367 879 368 880
rect 372 879 373 883
rect 399 883 405 884
rect 399 882 400 883
rect 367 878 373 879
rect 384 880 400 882
rect 367 875 373 876
rect 340 872 355 874
rect 358 874 364 875
rect 340 871 341 872
rect 335 870 341 871
rect 358 870 359 874
rect 363 870 364 874
rect 367 871 368 875
rect 372 874 373 875
rect 384 874 386 880
rect 399 879 400 880
rect 404 879 405 883
rect 399 878 405 879
rect 463 883 469 884
rect 463 879 464 883
rect 468 882 469 883
rect 583 883 589 884
rect 583 882 584 883
rect 468 880 506 882
rect 468 879 469 880
rect 463 878 469 879
rect 504 876 506 880
rect 564 880 584 882
rect 399 875 408 876
rect 463 875 472 876
rect 503 875 509 876
rect 543 875 549 876
rect 372 872 386 874
rect 390 874 396 875
rect 372 871 373 872
rect 367 870 373 871
rect 390 870 391 874
rect 395 870 396 874
rect 399 871 400 875
rect 407 871 408 875
rect 399 870 408 871
rect 422 874 428 875
rect 422 870 423 874
rect 427 870 428 874
rect 454 874 460 875
rect 230 869 236 870
rect 254 869 260 870
rect 278 869 284 870
rect 302 869 308 870
rect 326 869 332 870
rect 358 869 364 870
rect 390 869 396 870
rect 422 869 428 870
rect 431 871 437 872
rect 238 867 244 868
rect 238 863 239 867
rect 243 866 244 867
rect 398 867 404 868
rect 243 864 362 866
rect 243 863 244 864
rect 238 862 244 863
rect 360 860 362 864
rect 398 863 399 867
rect 403 866 404 867
rect 431 867 432 871
rect 436 867 437 871
rect 454 870 455 874
rect 459 870 460 874
rect 463 871 464 875
rect 471 871 472 875
rect 463 870 472 871
rect 494 874 500 875
rect 494 870 495 874
rect 499 870 500 874
rect 503 871 504 875
rect 508 871 509 875
rect 503 870 509 871
rect 534 874 540 875
rect 534 870 535 874
rect 539 870 540 874
rect 543 871 544 875
rect 548 874 549 875
rect 564 874 566 880
rect 583 879 584 880
rect 588 879 589 883
rect 631 883 637 884
rect 631 882 632 883
rect 583 878 589 879
rect 608 880 632 882
rect 583 875 589 876
rect 548 872 566 874
rect 574 874 580 875
rect 548 871 549 872
rect 543 870 549 871
rect 574 870 575 874
rect 579 870 580 874
rect 583 871 584 875
rect 588 874 589 875
rect 608 874 610 880
rect 631 879 632 880
rect 636 879 637 883
rect 671 883 677 884
rect 671 882 672 883
rect 631 878 637 879
rect 652 880 672 882
rect 631 875 637 876
rect 588 872 610 874
rect 622 874 628 875
rect 588 871 589 872
rect 583 870 589 871
rect 622 870 623 874
rect 627 870 628 874
rect 631 871 632 875
rect 636 874 637 875
rect 652 874 654 880
rect 671 879 672 880
rect 676 879 677 883
rect 671 878 677 879
rect 759 883 765 884
rect 759 879 760 883
rect 764 882 765 883
rect 871 883 877 884
rect 764 880 818 882
rect 764 879 765 880
rect 759 878 765 879
rect 816 876 818 880
rect 871 879 872 883
rect 876 882 877 883
rect 879 883 885 884
rect 879 882 880 883
rect 876 880 880 882
rect 876 879 877 880
rect 871 878 877 879
rect 879 879 880 880
rect 884 879 885 883
rect 935 883 941 884
rect 935 882 936 883
rect 879 878 885 879
rect 888 880 936 882
rect 759 875 768 876
rect 815 875 821 876
rect 871 875 877 876
rect 636 872 654 874
rect 662 874 668 875
rect 636 871 637 872
rect 631 870 637 871
rect 662 870 663 874
rect 667 870 668 874
rect 702 874 708 875
rect 454 869 460 870
rect 494 869 500 870
rect 534 869 540 870
rect 574 869 580 870
rect 622 869 628 870
rect 662 869 668 870
rect 671 871 677 872
rect 431 866 437 867
rect 606 867 612 868
rect 403 864 435 866
rect 403 863 404 864
rect 398 862 404 863
rect 606 863 607 867
rect 611 866 612 867
rect 671 867 672 871
rect 676 867 677 871
rect 702 870 703 874
rect 707 870 708 874
rect 750 874 756 875
rect 702 869 708 870
rect 711 871 717 872
rect 671 866 677 867
rect 711 867 712 871
rect 716 870 717 871
rect 750 870 751 874
rect 755 870 756 874
rect 759 871 760 875
rect 767 871 768 875
rect 759 870 768 871
rect 806 874 812 875
rect 806 870 807 874
rect 811 870 812 874
rect 815 871 816 875
rect 820 871 821 875
rect 815 870 821 871
rect 862 874 868 875
rect 862 870 863 874
rect 867 870 868 874
rect 871 871 872 875
rect 876 874 877 875
rect 888 874 890 880
rect 935 879 936 880
rect 940 879 941 883
rect 999 883 1005 884
rect 999 882 1000 883
rect 935 878 941 879
rect 968 880 1000 882
rect 935 875 941 876
rect 876 872 890 874
rect 926 874 932 875
rect 876 871 877 872
rect 871 870 877 871
rect 926 870 927 874
rect 931 870 932 874
rect 935 871 936 875
rect 940 874 941 875
rect 968 874 970 880
rect 999 879 1000 880
rect 1004 879 1005 883
rect 1063 883 1069 884
rect 1063 882 1064 883
rect 999 878 1005 879
rect 1032 880 1064 882
rect 999 875 1005 876
rect 940 872 970 874
rect 990 874 996 875
rect 940 871 941 872
rect 935 870 941 871
rect 990 870 991 874
rect 995 870 996 874
rect 999 871 1000 875
rect 1004 874 1005 875
rect 1032 874 1034 880
rect 1063 879 1064 880
rect 1068 879 1069 883
rect 1063 878 1069 879
rect 1183 883 1189 884
rect 1183 879 1184 883
rect 1188 882 1189 883
rect 1287 883 1293 884
rect 1188 880 1243 882
rect 1188 879 1189 880
rect 1183 878 1189 879
rect 1241 876 1243 880
rect 1287 879 1288 883
rect 1292 882 1293 883
rect 1335 883 1341 884
rect 1292 880 1323 882
rect 1292 879 1293 880
rect 1287 878 1293 879
rect 1063 875 1072 876
rect 1127 875 1133 876
rect 1183 875 1192 876
rect 1004 872 1034 874
rect 1054 874 1060 875
rect 1004 871 1005 872
rect 999 870 1005 871
rect 1054 870 1055 874
rect 1059 870 1060 874
rect 1063 871 1064 875
rect 1071 871 1072 875
rect 1063 870 1072 871
rect 1118 874 1124 875
rect 1118 870 1119 874
rect 1123 870 1124 874
rect 1127 871 1128 875
rect 1132 874 1133 875
rect 1174 874 1180 875
rect 1132 872 1161 874
rect 1132 871 1133 872
rect 1127 870 1133 871
rect 716 868 746 870
rect 750 869 756 870
rect 806 869 812 870
rect 862 869 868 870
rect 926 869 932 870
rect 990 869 996 870
rect 1054 869 1060 870
rect 1118 869 1124 870
rect 716 867 717 868
rect 711 866 717 867
rect 744 866 746 868
rect 778 867 784 868
rect 778 866 779 867
rect 611 864 674 866
rect 744 864 779 866
rect 611 863 612 864
rect 606 862 612 863
rect 778 863 779 864
rect 783 863 784 867
rect 778 862 784 863
rect 879 867 885 868
rect 879 863 880 867
rect 884 866 885 867
rect 1159 866 1161 872
rect 1174 870 1175 874
rect 1179 870 1180 874
rect 1183 871 1184 875
rect 1191 871 1192 875
rect 1183 870 1192 871
rect 1198 875 1204 876
rect 1239 875 1245 876
rect 1287 875 1296 876
rect 1198 871 1199 875
rect 1203 871 1204 875
rect 1198 870 1204 871
rect 1230 874 1236 875
rect 1230 870 1231 874
rect 1235 870 1236 874
rect 1239 871 1240 875
rect 1244 871 1245 875
rect 1239 870 1245 871
rect 1278 874 1284 875
rect 1278 870 1279 874
rect 1283 870 1284 874
rect 1287 871 1288 875
rect 1295 871 1296 875
rect 1287 870 1296 871
rect 1174 869 1180 870
rect 1200 868 1226 870
rect 1230 869 1236 870
rect 1278 869 1284 870
rect 1182 867 1188 868
rect 884 864 994 866
rect 884 863 885 864
rect 879 862 885 863
rect 992 860 994 864
rect 1096 864 1130 866
rect 1159 864 1178 866
rect 359 859 365 860
rect 655 859 661 860
rect 206 858 212 859
rect 206 854 207 858
rect 211 854 212 858
rect 230 858 236 859
rect 110 853 116 854
rect 206 853 212 854
rect 215 855 221 856
rect 110 849 111 853
rect 115 849 116 853
rect 215 851 216 855
rect 220 851 221 855
rect 230 854 231 858
rect 235 854 236 858
rect 254 858 260 859
rect 230 853 236 854
rect 239 855 245 856
rect 215 850 221 851
rect 239 851 240 855
rect 244 851 245 855
rect 254 854 255 858
rect 259 854 260 858
rect 286 858 292 859
rect 254 853 260 854
rect 263 855 269 856
rect 239 850 245 851
rect 263 851 264 855
rect 268 854 269 855
rect 286 854 287 858
rect 291 854 292 858
rect 318 858 324 859
rect 268 852 283 854
rect 286 853 292 854
rect 295 855 301 856
rect 268 851 269 852
rect 263 850 269 851
rect 110 848 116 849
rect 217 842 219 850
rect 241 846 243 850
rect 263 847 269 848
rect 263 846 264 847
rect 241 844 264 846
rect 263 843 264 844
rect 268 843 269 847
rect 281 846 283 852
rect 295 851 296 855
rect 300 854 301 855
rect 318 854 319 858
rect 323 854 324 858
rect 350 858 356 859
rect 300 852 307 854
rect 318 853 324 854
rect 327 855 333 856
rect 300 851 301 852
rect 295 850 301 851
rect 295 847 301 848
rect 295 846 296 847
rect 281 844 296 846
rect 263 842 269 843
rect 295 843 296 844
rect 300 843 301 847
rect 305 846 307 852
rect 327 851 328 855
rect 332 854 333 855
rect 350 854 351 858
rect 355 854 356 858
rect 359 855 360 859
rect 364 855 365 859
rect 359 854 365 855
rect 382 858 388 859
rect 382 854 383 858
rect 387 854 388 858
rect 414 858 420 859
rect 332 852 346 854
rect 350 853 356 854
rect 382 853 388 854
rect 391 855 397 856
rect 332 851 333 852
rect 327 850 333 851
rect 327 847 333 848
rect 327 846 328 847
rect 305 844 328 846
rect 295 842 301 843
rect 327 843 328 844
rect 332 843 333 847
rect 344 846 346 852
rect 391 851 392 855
rect 396 854 397 855
rect 414 854 415 858
rect 419 854 420 858
rect 446 858 452 859
rect 396 852 410 854
rect 414 853 420 854
rect 423 855 429 856
rect 396 851 397 852
rect 391 850 397 851
rect 359 847 365 848
rect 359 846 360 847
rect 344 844 360 846
rect 327 842 333 843
rect 359 843 360 844
rect 364 843 365 847
rect 359 842 365 843
rect 391 847 397 848
rect 391 843 392 847
rect 396 843 397 847
rect 408 846 410 852
rect 423 851 424 855
rect 428 854 429 855
rect 446 854 447 858
rect 451 854 452 858
rect 478 858 484 859
rect 428 852 442 854
rect 446 853 452 854
rect 455 855 461 856
rect 428 851 429 852
rect 423 850 429 851
rect 423 847 429 848
rect 423 846 424 847
rect 408 844 424 846
rect 391 842 397 843
rect 423 843 424 844
rect 428 843 429 847
rect 440 846 442 852
rect 455 851 456 855
rect 460 854 461 855
rect 478 854 479 858
rect 483 854 484 858
rect 510 858 516 859
rect 460 852 474 854
rect 478 853 484 854
rect 487 855 493 856
rect 460 851 461 852
rect 455 850 461 851
rect 455 847 461 848
rect 455 846 456 847
rect 440 844 456 846
rect 423 842 429 843
rect 455 843 456 844
rect 460 843 461 847
rect 472 846 474 852
rect 487 851 488 855
rect 492 854 493 855
rect 498 855 504 856
rect 498 854 499 855
rect 492 852 499 854
rect 492 851 493 852
rect 487 850 493 851
rect 498 851 499 852
rect 503 851 504 855
rect 510 854 511 858
rect 515 854 516 858
rect 550 858 556 859
rect 510 853 516 854
rect 519 855 525 856
rect 498 850 504 851
rect 519 851 520 855
rect 524 854 525 855
rect 550 854 551 858
rect 555 854 556 858
rect 598 858 604 859
rect 524 852 547 854
rect 550 853 556 854
rect 559 855 565 856
rect 524 851 525 852
rect 519 850 525 851
rect 487 847 493 848
rect 487 846 488 847
rect 472 844 488 846
rect 455 842 461 843
rect 487 843 488 844
rect 492 843 493 847
rect 545 846 547 852
rect 559 851 560 855
rect 564 854 565 855
rect 598 854 599 858
rect 603 854 604 858
rect 646 858 652 859
rect 564 852 586 854
rect 598 853 604 854
rect 607 855 613 856
rect 564 851 565 852
rect 559 850 565 851
rect 559 847 565 848
rect 559 846 560 847
rect 545 844 560 846
rect 487 842 493 843
rect 559 843 560 844
rect 564 843 565 847
rect 584 846 586 852
rect 607 851 608 855
rect 612 854 613 855
rect 646 854 647 858
rect 651 854 652 858
rect 655 855 656 859
rect 660 858 661 859
rect 663 859 669 860
rect 991 859 997 860
rect 1055 859 1061 860
rect 663 858 664 859
rect 660 856 664 858
rect 660 855 661 856
rect 655 854 661 855
rect 663 855 664 856
rect 668 855 669 859
rect 663 854 669 855
rect 702 858 708 859
rect 702 854 703 858
rect 707 854 708 858
rect 766 858 772 859
rect 612 852 634 854
rect 646 853 652 854
rect 702 853 708 854
rect 711 855 717 856
rect 612 851 613 852
rect 607 850 613 851
rect 607 847 613 848
rect 607 846 608 847
rect 584 844 608 846
rect 559 842 565 843
rect 607 843 608 844
rect 612 843 613 847
rect 632 846 634 852
rect 711 851 712 855
rect 716 851 717 855
rect 766 854 767 858
rect 771 854 772 858
rect 838 858 844 859
rect 766 853 772 854
rect 775 855 781 856
rect 711 850 717 851
rect 775 851 776 855
rect 780 851 781 855
rect 838 854 839 858
rect 843 854 844 858
rect 910 858 916 859
rect 838 853 844 854
rect 847 855 853 856
rect 775 850 781 851
rect 847 851 848 855
rect 852 854 853 855
rect 910 854 911 858
rect 915 854 916 858
rect 982 858 988 859
rect 852 852 886 854
rect 910 853 916 854
rect 919 855 925 856
rect 852 851 853 852
rect 847 850 853 851
rect 655 847 661 848
rect 655 846 656 847
rect 632 844 656 846
rect 607 842 613 843
rect 655 843 656 844
rect 660 843 661 847
rect 655 842 661 843
rect 666 847 672 848
rect 666 843 667 847
rect 671 846 672 847
rect 712 846 714 850
rect 671 844 714 846
rect 671 843 672 844
rect 666 842 672 843
rect 776 842 778 850
rect 884 846 886 852
rect 919 851 920 855
rect 924 854 925 855
rect 982 854 983 858
rect 987 854 988 858
rect 991 855 992 859
rect 996 855 997 859
rect 991 854 997 855
rect 1046 858 1052 859
rect 1046 854 1047 858
rect 1051 854 1052 858
rect 1055 855 1056 859
rect 1060 858 1061 859
rect 1096 858 1098 864
rect 1060 856 1098 858
rect 1102 858 1108 859
rect 1060 855 1061 856
rect 1055 854 1061 855
rect 1102 854 1103 858
rect 1107 854 1108 858
rect 1128 858 1130 864
rect 1150 859 1156 860
rect 1150 858 1151 859
rect 1128 856 1151 858
rect 924 852 958 854
rect 982 853 988 854
rect 1046 853 1052 854
rect 1102 853 1108 854
rect 1111 855 1117 856
rect 924 851 925 852
rect 919 850 925 851
rect 919 847 925 848
rect 919 846 920 847
rect 884 844 920 846
rect 919 843 920 844
rect 924 843 925 847
rect 956 846 958 852
rect 1111 851 1112 855
rect 1116 851 1117 855
rect 1150 855 1151 856
rect 1155 855 1156 859
rect 1150 854 1156 855
rect 1158 858 1164 859
rect 1158 854 1159 858
rect 1163 854 1164 858
rect 1176 858 1178 864
rect 1182 863 1183 867
rect 1187 866 1188 867
rect 1224 866 1226 868
rect 1302 867 1308 868
rect 1302 866 1303 867
rect 1187 864 1218 866
rect 1224 864 1303 866
rect 1187 863 1188 864
rect 1182 862 1188 863
rect 1216 860 1218 864
rect 1302 863 1303 864
rect 1307 863 1308 867
rect 1321 866 1323 880
rect 1335 879 1336 883
rect 1340 882 1341 883
rect 1423 883 1432 884
rect 1340 880 1395 882
rect 1340 879 1341 880
rect 1335 878 1341 879
rect 1393 876 1395 880
rect 1423 879 1424 883
rect 1431 879 1432 883
rect 1423 878 1432 879
rect 1446 879 1452 880
rect 1391 875 1397 876
rect 1446 875 1447 879
rect 1451 875 1452 879
rect 1326 874 1332 875
rect 1326 870 1327 874
rect 1331 870 1332 874
rect 1382 874 1388 875
rect 1326 869 1332 870
rect 1335 871 1341 872
rect 1335 867 1336 871
rect 1340 867 1341 871
rect 1382 870 1383 874
rect 1387 870 1388 874
rect 1391 871 1392 875
rect 1396 871 1397 875
rect 1391 870 1397 871
rect 1414 874 1420 875
rect 1446 874 1452 875
rect 1414 870 1415 874
rect 1419 870 1420 874
rect 1382 869 1388 870
rect 1414 869 1420 870
rect 1423 871 1429 872
rect 1335 866 1341 867
rect 1402 867 1408 868
rect 1321 864 1339 866
rect 1302 862 1308 863
rect 1402 863 1403 867
rect 1407 866 1408 867
rect 1423 867 1424 871
rect 1428 867 1429 871
rect 1423 866 1429 867
rect 1407 864 1427 866
rect 1407 863 1408 864
rect 1402 862 1408 863
rect 1198 859 1204 860
rect 1215 859 1221 860
rect 1423 859 1432 860
rect 1198 858 1199 859
rect 1176 856 1199 858
rect 1158 853 1164 854
rect 1167 855 1173 856
rect 1111 850 1117 851
rect 1167 851 1168 855
rect 1172 851 1173 855
rect 1198 855 1199 856
rect 1203 855 1204 859
rect 1198 854 1204 855
rect 1206 858 1212 859
rect 1206 854 1207 858
rect 1211 854 1212 858
rect 1215 855 1216 859
rect 1220 855 1221 859
rect 1215 854 1221 855
rect 1246 858 1252 859
rect 1246 854 1247 858
rect 1251 854 1252 858
rect 1294 858 1300 859
rect 1206 853 1212 854
rect 1246 853 1252 854
rect 1255 855 1261 856
rect 1167 850 1173 851
rect 1255 851 1256 855
rect 1260 851 1261 855
rect 1294 854 1295 858
rect 1299 854 1300 858
rect 1342 858 1348 859
rect 1294 853 1300 854
rect 1303 855 1309 856
rect 1255 850 1261 851
rect 1303 851 1304 855
rect 1308 851 1309 855
rect 1342 854 1343 858
rect 1347 854 1348 858
rect 1390 858 1396 859
rect 1342 853 1348 854
rect 1351 855 1357 856
rect 1303 850 1309 851
rect 1351 851 1352 855
rect 1356 851 1357 855
rect 1390 854 1391 858
rect 1395 854 1396 858
rect 1414 858 1420 859
rect 1390 853 1396 854
rect 1399 855 1405 856
rect 1351 850 1357 851
rect 1399 851 1400 855
rect 1404 851 1405 855
rect 1414 854 1415 858
rect 1419 854 1420 858
rect 1423 855 1424 859
rect 1431 855 1432 859
rect 1423 854 1432 855
rect 1414 853 1420 854
rect 1446 853 1452 854
rect 1399 850 1405 851
rect 991 847 997 848
rect 991 846 992 847
rect 956 844 992 846
rect 919 842 925 843
rect 991 843 992 844
rect 996 843 997 847
rect 991 842 997 843
rect 1055 847 1061 848
rect 1055 843 1056 847
rect 1060 846 1061 847
rect 1112 846 1114 850
rect 1060 844 1114 846
rect 1060 843 1061 844
rect 1055 842 1061 843
rect 1169 842 1171 850
rect 1215 847 1221 848
rect 1215 843 1216 847
rect 1220 846 1221 847
rect 1257 846 1259 850
rect 1220 844 1259 846
rect 1220 843 1221 844
rect 1215 842 1221 843
rect 1304 842 1306 850
rect 1352 842 1354 850
rect 1401 846 1403 850
rect 1446 849 1447 853
rect 1451 849 1452 853
rect 1446 848 1452 849
rect 1423 847 1429 848
rect 1423 846 1424 847
rect 1401 844 1424 846
rect 1423 843 1424 844
rect 1428 843 1429 847
rect 1423 842 1429 843
rect 217 840 243 842
rect 744 840 778 842
rect 1140 840 1171 842
rect 1257 840 1306 842
rect 1328 840 1354 842
rect 239 839 245 840
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 239 835 240 839
rect 244 835 245 839
rect 239 834 245 835
rect 711 839 717 840
rect 711 835 712 839
rect 716 838 717 839
rect 744 838 746 840
rect 716 836 746 838
rect 1111 839 1117 840
rect 716 835 717 836
rect 711 834 717 835
rect 775 835 784 836
rect 110 830 116 831
rect 206 832 212 833
rect 230 832 236 833
rect 206 828 207 832
rect 211 828 212 832
rect 206 827 212 828
rect 215 831 221 832
rect 215 827 216 831
rect 220 830 221 831
rect 220 828 227 830
rect 220 827 221 828
rect 215 826 221 827
rect 225 822 227 828
rect 230 828 231 832
rect 235 828 236 832
rect 230 827 236 828
rect 254 832 260 833
rect 254 828 255 832
rect 259 828 260 832
rect 254 827 260 828
rect 286 832 292 833
rect 286 828 287 832
rect 291 828 292 832
rect 286 827 292 828
rect 318 832 324 833
rect 318 828 319 832
rect 323 828 324 832
rect 318 827 324 828
rect 350 832 356 833
rect 350 828 351 832
rect 355 828 356 832
rect 350 827 356 828
rect 382 832 388 833
rect 382 828 383 832
rect 387 828 388 832
rect 382 827 388 828
rect 414 832 420 833
rect 414 828 415 832
rect 419 828 420 832
rect 414 827 420 828
rect 446 832 452 833
rect 446 828 447 832
rect 451 828 452 832
rect 446 827 452 828
rect 478 832 484 833
rect 478 828 479 832
rect 483 828 484 832
rect 478 827 484 828
rect 510 832 516 833
rect 550 832 556 833
rect 510 828 511 832
rect 515 828 516 832
rect 510 827 516 828
rect 519 831 525 832
rect 519 827 520 831
rect 524 830 525 831
rect 534 831 540 832
rect 534 830 535 831
rect 524 828 535 830
rect 524 827 525 828
rect 519 826 525 827
rect 534 827 535 828
rect 539 827 540 831
rect 550 828 551 832
rect 555 828 556 832
rect 550 827 556 828
rect 598 832 604 833
rect 598 828 599 832
rect 603 828 604 832
rect 598 827 604 828
rect 646 832 652 833
rect 646 828 647 832
rect 651 828 652 832
rect 646 827 652 828
rect 702 832 708 833
rect 702 828 703 832
rect 707 828 708 832
rect 702 827 708 828
rect 766 832 772 833
rect 766 828 767 832
rect 771 828 772 832
rect 775 831 776 835
rect 783 831 784 835
rect 1111 835 1112 839
rect 1116 838 1117 839
rect 1140 838 1142 840
rect 1116 836 1142 838
rect 1255 839 1261 840
rect 1116 835 1117 836
rect 1111 834 1117 835
rect 1167 835 1173 836
rect 775 830 784 831
rect 838 832 844 833
rect 910 832 916 833
rect 766 827 772 828
rect 838 828 839 832
rect 843 828 844 832
rect 838 827 844 828
rect 847 831 856 832
rect 847 827 848 831
rect 855 827 856 831
rect 910 828 911 832
rect 915 828 916 832
rect 910 827 916 828
rect 982 832 988 833
rect 982 828 983 832
rect 987 828 988 832
rect 982 827 988 828
rect 1046 832 1052 833
rect 1046 828 1047 832
rect 1051 828 1052 832
rect 1046 827 1052 828
rect 1102 832 1108 833
rect 1102 828 1103 832
rect 1107 828 1108 832
rect 1102 827 1108 828
rect 1158 832 1164 833
rect 1158 828 1159 832
rect 1163 828 1164 832
rect 1167 831 1168 835
rect 1172 834 1173 835
rect 1182 835 1188 836
rect 1182 834 1183 835
rect 1172 832 1183 834
rect 1172 831 1173 832
rect 1167 830 1173 831
rect 1182 831 1183 832
rect 1187 831 1188 835
rect 1255 835 1256 839
rect 1260 835 1261 839
rect 1255 834 1261 835
rect 1303 835 1309 836
rect 1182 830 1188 831
rect 1206 832 1212 833
rect 1158 827 1164 828
rect 1206 828 1207 832
rect 1211 828 1212 832
rect 1206 827 1212 828
rect 1246 832 1252 833
rect 1246 828 1247 832
rect 1251 828 1252 832
rect 1246 827 1252 828
rect 1294 832 1300 833
rect 1294 828 1295 832
rect 1299 828 1300 832
rect 1303 831 1304 835
rect 1308 834 1309 835
rect 1328 834 1330 840
rect 1308 832 1330 834
rect 1446 835 1452 836
rect 1342 832 1348 833
rect 1390 832 1396 833
rect 1414 832 1420 833
rect 1308 831 1309 832
rect 1303 830 1309 831
rect 1342 828 1343 832
rect 1347 828 1348 832
rect 1294 827 1300 828
rect 1302 827 1308 828
rect 1342 827 1348 828
rect 1351 831 1357 832
rect 1351 827 1352 831
rect 1356 827 1357 831
rect 1390 828 1391 832
rect 1395 828 1396 832
rect 1390 827 1396 828
rect 1399 831 1408 832
rect 1399 827 1400 831
rect 1407 827 1408 831
rect 1414 828 1415 832
rect 1419 828 1420 832
rect 1446 831 1447 835
rect 1451 831 1452 835
rect 1446 830 1452 831
rect 1414 827 1420 828
rect 534 826 540 827
rect 847 826 856 827
rect 247 823 253 824
rect 247 822 248 823
rect 134 820 140 821
rect 110 817 116 818
rect 110 813 111 817
rect 115 813 116 817
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 158 820 164 821
rect 158 816 159 820
rect 163 816 164 820
rect 158 815 164 816
rect 182 820 188 821
rect 182 816 183 820
rect 187 816 188 820
rect 182 815 188 816
rect 214 820 220 821
rect 225 820 248 822
rect 214 816 215 820
rect 219 816 220 820
rect 247 819 248 820
rect 252 819 253 823
rect 1302 823 1303 827
rect 1307 826 1308 827
rect 1351 826 1357 827
rect 1399 826 1408 827
rect 1307 824 1339 826
rect 1307 823 1308 824
rect 1302 822 1308 823
rect 1337 822 1339 824
rect 1352 822 1354 826
rect 247 818 253 819
rect 262 820 268 821
rect 214 815 220 816
rect 262 816 263 820
rect 267 816 268 820
rect 262 815 268 816
rect 310 820 316 821
rect 310 816 311 820
rect 315 816 316 820
rect 310 815 316 816
rect 366 820 372 821
rect 366 816 367 820
rect 371 816 372 820
rect 366 815 372 816
rect 430 820 436 821
rect 430 816 431 820
rect 435 816 436 820
rect 430 815 436 816
rect 486 820 492 821
rect 486 816 487 820
rect 491 816 492 820
rect 486 815 492 816
rect 542 820 548 821
rect 542 816 543 820
rect 547 816 548 820
rect 542 815 548 816
rect 598 820 604 821
rect 598 816 599 820
rect 603 816 604 820
rect 598 815 604 816
rect 654 820 660 821
rect 710 820 716 821
rect 654 816 655 820
rect 659 816 660 820
rect 654 815 660 816
rect 663 819 672 820
rect 663 815 664 819
rect 671 815 672 819
rect 710 816 711 820
rect 715 816 716 820
rect 710 815 716 816
rect 766 820 772 821
rect 766 816 767 820
rect 771 816 772 820
rect 766 815 772 816
rect 814 820 820 821
rect 814 816 815 820
rect 819 816 820 820
rect 814 815 820 816
rect 862 820 868 821
rect 862 816 863 820
rect 867 816 868 820
rect 862 815 868 816
rect 902 820 908 821
rect 902 816 903 820
rect 907 816 908 820
rect 902 815 908 816
rect 934 820 940 821
rect 934 816 935 820
rect 939 816 940 820
rect 934 815 940 816
rect 966 820 972 821
rect 966 816 967 820
rect 971 816 972 820
rect 966 815 972 816
rect 990 820 996 821
rect 990 816 991 820
rect 995 816 996 820
rect 990 815 996 816
rect 1014 820 1020 821
rect 1014 816 1015 820
rect 1019 816 1020 820
rect 1014 815 1020 816
rect 1038 820 1044 821
rect 1038 816 1039 820
rect 1043 816 1044 820
rect 1038 815 1044 816
rect 1062 820 1068 821
rect 1062 816 1063 820
rect 1067 816 1068 820
rect 1062 815 1068 816
rect 1094 820 1100 821
rect 1094 816 1095 820
rect 1099 816 1100 820
rect 1094 815 1100 816
rect 1126 820 1132 821
rect 1126 816 1127 820
rect 1131 816 1132 820
rect 1126 815 1132 816
rect 1166 820 1172 821
rect 1166 816 1167 820
rect 1171 816 1172 820
rect 1166 815 1172 816
rect 1206 820 1212 821
rect 1206 816 1207 820
rect 1211 816 1212 820
rect 1206 815 1212 816
rect 1254 820 1260 821
rect 1254 816 1255 820
rect 1259 816 1260 820
rect 1254 815 1260 816
rect 1310 820 1316 821
rect 1337 820 1354 822
rect 1374 820 1380 821
rect 1310 816 1311 820
rect 1315 816 1316 820
rect 1310 815 1316 816
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1414 820 1420 821
rect 1414 816 1415 820
rect 1419 816 1420 820
rect 1414 815 1420 816
rect 1446 817 1452 818
rect 663 814 672 815
rect 110 812 116 813
rect 1446 813 1447 817
rect 1451 813 1452 817
rect 1446 812 1452 813
rect 143 811 149 812
rect 143 807 144 811
rect 148 810 149 811
rect 418 811 424 812
rect 418 810 419 811
rect 148 808 419 810
rect 148 807 149 808
rect 143 806 149 807
rect 418 807 419 808
rect 423 807 424 811
rect 418 806 424 807
rect 439 811 445 812
rect 439 807 440 811
rect 444 810 445 811
rect 498 811 504 812
rect 498 810 499 811
rect 444 808 499 810
rect 444 807 445 808
rect 439 806 445 807
rect 498 807 499 808
rect 503 807 504 811
rect 498 806 504 807
rect 610 811 616 812
rect 610 807 611 811
rect 615 810 616 811
rect 719 811 725 812
rect 719 810 720 811
rect 615 808 720 810
rect 615 807 616 808
rect 610 806 616 807
rect 719 807 720 808
rect 724 807 725 811
rect 719 806 725 807
rect 778 811 784 812
rect 778 807 779 811
rect 783 810 784 811
rect 823 811 829 812
rect 823 810 824 811
rect 783 808 824 810
rect 783 807 784 808
rect 778 806 784 807
rect 823 807 824 808
rect 828 807 829 811
rect 823 806 829 807
rect 911 811 917 812
rect 911 807 912 811
rect 916 810 917 811
rect 946 811 952 812
rect 946 810 947 811
rect 916 808 947 810
rect 916 807 917 808
rect 911 806 917 807
rect 946 807 947 808
rect 951 807 952 811
rect 946 806 952 807
rect 975 811 981 812
rect 975 807 976 811
rect 980 810 981 811
rect 1002 811 1008 812
rect 1002 810 1003 811
rect 980 808 1003 810
rect 980 807 981 808
rect 975 806 981 807
rect 1002 807 1003 808
rect 1007 807 1008 811
rect 1002 806 1008 807
rect 1023 811 1029 812
rect 1023 807 1024 811
rect 1028 810 1029 811
rect 1050 811 1056 812
rect 1050 810 1051 811
rect 1028 808 1051 810
rect 1028 807 1029 808
rect 1023 806 1029 807
rect 1050 807 1051 808
rect 1055 807 1056 811
rect 1074 811 1080 812
rect 1074 810 1075 811
rect 1050 806 1056 807
rect 1064 808 1075 810
rect 167 803 173 804
rect 167 802 168 803
rect 152 800 168 802
rect 110 799 116 800
rect 110 795 111 799
rect 115 795 116 799
rect 143 795 149 796
rect 110 794 116 795
rect 134 794 140 795
rect 134 790 135 794
rect 139 790 140 794
rect 143 791 144 795
rect 148 794 149 795
rect 152 794 154 800
rect 167 799 168 800
rect 172 799 173 803
rect 191 803 197 804
rect 191 802 192 803
rect 167 798 173 799
rect 176 800 192 802
rect 167 795 173 796
rect 148 792 154 794
rect 158 794 164 795
rect 148 791 149 792
rect 143 790 149 791
rect 158 790 159 794
rect 163 790 164 794
rect 167 791 168 795
rect 172 794 173 795
rect 176 794 178 800
rect 191 799 192 800
rect 196 799 197 803
rect 223 803 229 804
rect 223 802 224 803
rect 191 798 197 799
rect 209 800 224 802
rect 191 795 197 796
rect 172 792 178 794
rect 182 794 188 795
rect 172 791 173 792
rect 167 790 173 791
rect 182 790 183 794
rect 187 790 188 794
rect 191 791 192 795
rect 196 794 197 795
rect 209 794 211 800
rect 223 799 224 800
rect 228 799 229 803
rect 271 803 277 804
rect 271 802 272 803
rect 223 798 229 799
rect 248 800 272 802
rect 223 795 229 796
rect 196 792 211 794
rect 214 794 220 795
rect 196 791 197 792
rect 191 790 197 791
rect 214 790 215 794
rect 219 790 220 794
rect 223 791 224 795
rect 228 794 229 795
rect 248 794 250 800
rect 271 799 272 800
rect 276 799 277 803
rect 319 803 325 804
rect 319 802 320 803
rect 271 798 277 799
rect 296 800 320 802
rect 271 795 277 796
rect 228 792 250 794
rect 262 794 268 795
rect 228 791 229 792
rect 223 790 229 791
rect 262 790 263 794
rect 267 790 268 794
rect 271 791 272 795
rect 276 794 277 795
rect 296 794 298 800
rect 319 799 320 800
rect 324 799 325 803
rect 375 803 381 804
rect 375 802 376 803
rect 319 798 325 799
rect 348 800 376 802
rect 319 795 325 796
rect 276 792 298 794
rect 310 794 316 795
rect 276 791 277 792
rect 271 790 277 791
rect 310 790 311 794
rect 315 790 316 794
rect 319 791 320 795
rect 324 794 325 795
rect 348 794 350 800
rect 375 799 376 800
rect 380 799 381 803
rect 495 803 501 804
rect 495 802 496 803
rect 375 798 381 799
rect 468 800 496 802
rect 439 795 445 796
rect 324 792 350 794
rect 366 794 372 795
rect 324 791 325 792
rect 319 790 325 791
rect 366 790 367 794
rect 371 790 372 794
rect 430 794 436 795
rect 134 789 140 790
rect 158 789 164 790
rect 182 789 188 790
rect 214 789 220 790
rect 262 789 268 790
rect 310 789 316 790
rect 366 789 372 790
rect 375 791 381 792
rect 247 787 253 788
rect 247 783 248 787
rect 252 786 253 787
rect 375 787 376 791
rect 380 787 381 791
rect 430 790 431 794
rect 435 790 436 794
rect 439 791 440 795
rect 444 794 445 795
rect 468 794 470 800
rect 495 799 496 800
rect 500 799 501 803
rect 551 803 557 804
rect 551 802 552 803
rect 495 798 501 799
rect 524 800 552 802
rect 495 795 501 796
rect 444 792 470 794
rect 486 794 492 795
rect 444 791 445 792
rect 439 790 445 791
rect 486 790 487 794
rect 491 790 492 794
rect 495 791 496 795
rect 500 794 501 795
rect 524 794 526 800
rect 551 799 552 800
rect 556 799 557 803
rect 551 798 557 799
rect 607 803 613 804
rect 607 799 608 803
rect 612 802 613 803
rect 775 803 781 804
rect 612 800 666 802
rect 612 799 613 800
rect 607 798 613 799
rect 664 796 666 800
rect 775 799 776 803
rect 780 802 781 803
rect 806 803 812 804
rect 806 802 807 803
rect 780 800 807 802
rect 780 799 781 800
rect 775 798 781 799
rect 806 799 807 800
rect 811 799 812 803
rect 806 798 812 799
rect 871 803 877 804
rect 871 799 872 803
rect 876 802 877 803
rect 943 803 949 804
rect 876 800 914 802
rect 876 799 877 800
rect 871 798 877 799
rect 912 796 914 800
rect 943 799 944 803
rect 948 802 949 803
rect 999 803 1005 804
rect 948 800 978 802
rect 948 799 949 800
rect 943 798 949 799
rect 976 796 978 800
rect 999 799 1000 803
rect 1004 802 1005 803
rect 1007 803 1013 804
rect 1007 802 1008 803
rect 1004 800 1008 802
rect 1004 799 1005 800
rect 999 798 1005 799
rect 1007 799 1008 800
rect 1012 799 1013 803
rect 1007 798 1013 799
rect 1047 803 1053 804
rect 1047 799 1048 803
rect 1052 802 1053 803
rect 1064 802 1066 808
rect 1074 807 1075 808
rect 1079 807 1080 811
rect 1135 811 1141 812
rect 1074 806 1080 807
rect 1102 807 1109 808
rect 1052 800 1066 802
rect 1071 803 1077 804
rect 1052 799 1053 800
rect 1047 798 1053 799
rect 1071 799 1072 803
rect 1076 802 1077 803
rect 1102 803 1103 807
rect 1108 803 1109 807
rect 1135 807 1136 811
rect 1140 810 1141 811
rect 1178 811 1184 812
rect 1178 810 1179 811
rect 1140 808 1179 810
rect 1140 807 1141 808
rect 1135 806 1141 807
rect 1178 807 1179 808
rect 1183 807 1184 811
rect 1178 806 1184 807
rect 1215 811 1221 812
rect 1215 807 1216 811
rect 1220 810 1221 811
rect 1266 811 1272 812
rect 1266 810 1267 811
rect 1220 808 1267 810
rect 1220 807 1221 808
rect 1215 806 1221 807
rect 1266 807 1267 808
rect 1271 807 1272 811
rect 1266 806 1272 807
rect 1274 811 1280 812
rect 1274 807 1275 811
rect 1279 810 1280 811
rect 1319 811 1325 812
rect 1319 810 1320 811
rect 1279 808 1320 810
rect 1279 807 1280 808
rect 1274 806 1280 807
rect 1319 807 1320 808
rect 1324 807 1325 811
rect 1319 806 1325 807
rect 1102 802 1109 803
rect 1175 803 1181 804
rect 1076 800 1090 802
rect 1076 799 1077 800
rect 1071 798 1077 799
rect 607 795 616 796
rect 663 795 669 796
rect 775 795 784 796
rect 823 795 829 796
rect 500 792 526 794
rect 542 794 548 795
rect 500 791 501 792
rect 495 790 501 791
rect 542 790 543 794
rect 547 790 548 794
rect 598 794 604 795
rect 430 789 436 790
rect 486 789 492 790
rect 542 789 548 790
rect 551 791 557 792
rect 375 786 381 787
rect 534 787 540 788
rect 252 784 379 786
rect 252 783 253 784
rect 247 782 253 783
rect 534 783 535 787
rect 539 786 540 787
rect 551 787 552 791
rect 556 787 557 791
rect 598 790 599 794
rect 603 790 604 794
rect 607 791 608 795
rect 615 791 616 795
rect 607 790 616 791
rect 654 794 660 795
rect 654 790 655 794
rect 659 790 660 794
rect 663 791 664 795
rect 668 791 669 795
rect 663 790 669 791
rect 710 794 716 795
rect 710 790 711 794
rect 715 790 716 794
rect 766 794 772 795
rect 598 789 604 790
rect 654 789 660 790
rect 710 789 716 790
rect 719 791 725 792
rect 551 786 557 787
rect 559 787 565 788
rect 539 784 554 786
rect 539 783 540 784
rect 534 782 540 783
rect 559 783 560 787
rect 564 786 565 787
rect 719 787 720 791
rect 724 790 725 791
rect 730 791 736 792
rect 730 790 731 791
rect 724 788 731 790
rect 724 787 725 788
rect 719 786 725 787
rect 730 787 731 788
rect 735 787 736 791
rect 766 790 767 794
rect 771 790 772 794
rect 775 791 776 795
rect 783 791 784 795
rect 775 790 784 791
rect 814 794 820 795
rect 814 790 815 794
rect 819 790 820 794
rect 823 791 824 795
rect 828 794 829 795
rect 850 795 856 796
rect 911 795 917 796
rect 943 795 952 796
rect 975 795 981 796
rect 999 795 1008 796
rect 1047 795 1056 796
rect 1071 795 1080 796
rect 850 794 851 795
rect 828 792 851 794
rect 828 791 829 792
rect 823 790 829 791
rect 850 791 851 792
rect 855 791 856 795
rect 850 790 856 791
rect 862 794 868 795
rect 862 790 863 794
rect 867 790 868 794
rect 902 794 908 795
rect 766 789 772 790
rect 814 789 820 790
rect 862 789 868 790
rect 871 791 877 792
rect 730 786 736 787
rect 871 787 872 791
rect 876 787 877 791
rect 902 790 903 794
rect 907 790 908 794
rect 911 791 912 795
rect 916 791 917 795
rect 911 790 917 791
rect 934 794 940 795
rect 934 790 935 794
rect 939 790 940 794
rect 943 791 944 795
rect 951 791 952 795
rect 943 790 952 791
rect 966 794 972 795
rect 966 790 967 794
rect 971 790 972 794
rect 975 791 976 795
rect 980 791 981 795
rect 975 790 981 791
rect 990 794 996 795
rect 990 790 991 794
rect 995 790 996 794
rect 999 791 1000 795
rect 1007 791 1008 795
rect 999 790 1008 791
rect 1014 794 1020 795
rect 1014 790 1015 794
rect 1019 790 1020 794
rect 1038 794 1044 795
rect 902 789 908 790
rect 934 789 940 790
rect 966 789 972 790
rect 990 789 996 790
rect 1014 789 1020 790
rect 1023 791 1029 792
rect 871 786 877 787
rect 950 787 956 788
rect 564 784 586 786
rect 873 784 946 786
rect 564 783 565 784
rect 559 782 565 783
rect 584 780 586 784
rect 806 783 812 784
rect 415 779 424 780
rect 583 779 589 780
rect 806 779 807 783
rect 811 780 812 783
rect 811 779 813 780
rect 134 778 140 779
rect 134 774 135 778
rect 139 774 140 778
rect 158 778 164 779
rect 110 773 116 774
rect 134 773 140 774
rect 143 775 149 776
rect 110 769 111 773
rect 115 769 116 773
rect 143 771 144 775
rect 148 771 149 775
rect 158 774 159 778
rect 163 774 164 778
rect 182 778 188 779
rect 158 773 164 774
rect 167 775 173 776
rect 143 770 149 771
rect 167 771 168 775
rect 172 771 173 775
rect 182 774 183 778
rect 187 774 188 778
rect 222 778 228 779
rect 182 773 188 774
rect 191 775 197 776
rect 167 770 173 771
rect 191 771 192 775
rect 196 774 197 775
rect 222 774 223 778
rect 227 774 228 778
rect 278 778 284 779
rect 196 772 214 774
rect 222 773 228 774
rect 231 775 237 776
rect 196 771 197 772
rect 191 770 197 771
rect 110 768 116 769
rect 145 762 147 770
rect 169 766 171 770
rect 191 767 197 768
rect 191 766 192 767
rect 169 764 192 766
rect 191 763 192 764
rect 196 763 197 767
rect 212 766 214 772
rect 231 771 232 775
rect 236 774 237 775
rect 278 774 279 778
rect 283 774 284 778
rect 342 778 348 779
rect 236 772 262 774
rect 278 773 284 774
rect 287 775 293 776
rect 236 771 237 772
rect 231 770 237 771
rect 231 767 237 768
rect 231 766 232 767
rect 212 764 232 766
rect 191 762 197 763
rect 231 763 232 764
rect 236 763 237 767
rect 260 766 262 772
rect 287 771 288 775
rect 292 774 293 775
rect 342 774 343 778
rect 347 774 348 778
rect 406 778 412 779
rect 292 772 322 774
rect 342 773 348 774
rect 351 775 357 776
rect 292 771 293 772
rect 287 770 293 771
rect 287 767 293 768
rect 287 766 288 767
rect 260 764 288 766
rect 231 762 237 763
rect 287 763 288 764
rect 292 763 293 767
rect 287 762 293 763
rect 320 762 322 772
rect 351 771 352 775
rect 356 771 357 775
rect 406 774 407 778
rect 411 774 412 778
rect 415 775 416 779
rect 423 775 424 779
rect 415 774 424 775
rect 462 778 468 779
rect 462 774 463 778
rect 467 774 468 778
rect 518 778 524 779
rect 406 773 412 774
rect 462 773 468 774
rect 471 775 477 776
rect 351 770 357 771
rect 471 771 472 775
rect 476 774 477 775
rect 510 775 516 776
rect 510 774 511 775
rect 476 772 511 774
rect 476 771 477 772
rect 471 770 477 771
rect 510 771 511 772
rect 515 771 516 775
rect 518 774 519 778
rect 523 774 524 778
rect 574 778 580 779
rect 518 773 524 774
rect 527 775 533 776
rect 510 770 516 771
rect 527 771 528 775
rect 532 771 533 775
rect 574 774 575 778
rect 579 774 580 778
rect 583 775 584 779
rect 588 775 589 779
rect 583 774 589 775
rect 622 778 628 779
rect 622 774 623 778
rect 627 774 628 778
rect 670 778 676 779
rect 574 773 580 774
rect 622 773 628 774
rect 631 775 640 776
rect 527 770 533 771
rect 631 771 632 775
rect 639 771 640 775
rect 670 774 671 778
rect 675 774 676 778
rect 718 778 724 779
rect 670 773 676 774
rect 679 775 685 776
rect 631 770 640 771
rect 679 771 680 775
rect 684 771 685 775
rect 718 774 719 778
rect 723 774 724 778
rect 758 778 764 779
rect 718 773 724 774
rect 727 775 733 776
rect 679 770 685 771
rect 727 771 728 775
rect 732 774 733 775
rect 735 775 741 776
rect 735 774 736 775
rect 732 772 736 774
rect 732 771 733 772
rect 727 770 733 771
rect 735 771 736 772
rect 740 771 741 775
rect 758 774 759 778
rect 763 774 764 778
rect 798 778 804 779
rect 806 778 808 779
rect 758 773 764 774
rect 767 775 773 776
rect 735 770 741 771
rect 767 771 768 775
rect 772 774 773 775
rect 798 774 799 778
rect 803 774 804 778
rect 807 775 808 778
rect 812 775 813 779
rect 807 774 813 775
rect 838 778 844 779
rect 838 774 839 778
rect 843 774 844 778
rect 878 778 884 779
rect 772 772 790 774
rect 798 773 804 774
rect 838 773 844 774
rect 847 775 853 776
rect 772 771 773 772
rect 767 770 773 771
rect 353 766 355 770
rect 415 767 421 768
rect 415 766 416 767
rect 353 764 416 766
rect 415 763 416 764
rect 420 763 421 767
rect 415 762 421 763
rect 471 767 477 768
rect 471 763 472 767
rect 476 766 477 767
rect 528 766 530 770
rect 476 764 530 766
rect 476 763 477 764
rect 471 762 477 763
rect 583 763 589 764
rect 145 760 171 762
rect 320 760 355 762
rect 167 759 173 760
rect 110 755 116 756
rect 110 751 111 755
rect 115 751 116 755
rect 167 755 168 759
rect 172 755 173 759
rect 167 754 173 755
rect 351 759 357 760
rect 351 755 352 759
rect 356 755 357 759
rect 351 754 357 755
rect 527 759 533 760
rect 527 755 528 759
rect 532 758 533 759
rect 559 759 565 760
rect 559 758 560 759
rect 532 756 560 758
rect 532 755 533 756
rect 527 754 533 755
rect 559 755 560 756
rect 564 755 565 759
rect 583 759 584 763
rect 588 762 589 763
rect 622 763 628 764
rect 622 762 623 763
rect 588 760 623 762
rect 588 759 589 760
rect 583 758 589 759
rect 622 759 623 760
rect 627 759 628 763
rect 622 758 628 759
rect 631 763 637 764
rect 631 759 632 763
rect 636 762 637 763
rect 679 762 681 770
rect 727 767 736 768
rect 727 763 728 767
rect 735 763 736 767
rect 788 766 790 772
rect 847 771 848 775
rect 852 774 853 775
rect 862 775 868 776
rect 862 774 863 775
rect 852 772 863 774
rect 852 771 853 772
rect 847 770 853 771
rect 862 771 863 772
rect 867 771 868 775
rect 878 774 879 778
rect 883 774 884 778
rect 918 778 924 779
rect 878 773 884 774
rect 887 775 893 776
rect 862 770 868 771
rect 887 771 888 775
rect 892 771 893 775
rect 918 774 919 778
rect 923 774 924 778
rect 918 773 924 774
rect 927 775 933 776
rect 887 770 893 771
rect 927 771 928 775
rect 932 771 933 775
rect 927 770 933 771
rect 807 767 813 768
rect 807 766 808 767
rect 788 764 808 766
rect 727 762 736 763
rect 807 763 808 764
rect 812 763 813 767
rect 807 762 813 763
rect 847 767 853 768
rect 847 763 848 767
rect 852 766 853 767
rect 888 766 890 770
rect 852 764 890 766
rect 852 763 853 764
rect 847 762 853 763
rect 928 762 930 770
rect 944 766 946 784
rect 950 783 951 787
rect 955 786 956 787
rect 1023 787 1024 791
rect 1028 787 1029 791
rect 1038 790 1039 794
rect 1043 790 1044 794
rect 1047 791 1048 795
rect 1055 791 1056 795
rect 1047 790 1056 791
rect 1062 794 1068 795
rect 1062 790 1063 794
rect 1067 790 1068 794
rect 1071 791 1072 795
rect 1079 791 1080 795
rect 1071 790 1080 791
rect 1038 789 1044 790
rect 1062 789 1068 790
rect 1023 786 1029 787
rect 1088 786 1090 800
rect 1175 799 1176 803
rect 1180 802 1181 803
rect 1263 803 1269 804
rect 1180 800 1203 802
rect 1180 799 1181 800
rect 1175 798 1181 799
rect 1158 795 1164 796
rect 1175 795 1184 796
rect 1094 794 1100 795
rect 1094 790 1095 794
rect 1099 790 1100 794
rect 1126 794 1132 795
rect 1094 789 1100 790
rect 1103 791 1109 792
rect 1103 787 1104 791
rect 1108 787 1109 791
rect 1126 790 1127 794
rect 1131 790 1132 794
rect 1126 789 1132 790
rect 1135 791 1141 792
rect 1103 786 1109 787
rect 1135 787 1136 791
rect 1140 790 1141 791
rect 1158 791 1159 795
rect 1163 791 1164 795
rect 1158 790 1164 791
rect 1166 794 1172 795
rect 1166 790 1167 794
rect 1171 790 1172 794
rect 1175 791 1176 795
rect 1183 791 1184 795
rect 1175 790 1184 791
rect 1140 788 1161 790
rect 1166 789 1172 790
rect 1140 787 1141 788
rect 1135 786 1141 787
rect 1201 786 1203 800
rect 1263 799 1264 803
rect 1268 802 1269 803
rect 1383 803 1389 804
rect 1268 800 1294 802
rect 1268 799 1269 800
rect 1263 798 1269 799
rect 1263 795 1272 796
rect 1206 794 1212 795
rect 1206 790 1207 794
rect 1211 790 1212 794
rect 1254 794 1260 795
rect 1206 789 1212 790
rect 1215 791 1221 792
rect 1215 787 1216 791
rect 1220 787 1221 791
rect 1254 790 1255 794
rect 1259 790 1260 794
rect 1263 791 1264 795
rect 1271 791 1272 795
rect 1263 790 1272 791
rect 1254 789 1260 790
rect 1215 786 1221 787
rect 1274 787 1280 788
rect 1274 786 1275 787
rect 955 784 971 786
rect 1016 784 1026 786
rect 1088 784 1106 786
rect 1159 784 1186 786
rect 1201 784 1218 786
rect 1224 784 1275 786
rect 955 783 956 784
rect 950 782 956 783
rect 969 780 971 784
rect 1007 783 1013 784
rect 967 779 973 780
rect 1007 779 1008 783
rect 1012 782 1013 783
rect 1016 782 1018 784
rect 1012 780 1018 782
rect 1150 783 1156 784
rect 1012 779 1013 780
rect 1150 779 1151 783
rect 1155 782 1156 783
rect 1159 782 1161 784
rect 1155 780 1161 782
rect 1184 782 1186 784
rect 1224 782 1226 784
rect 1274 783 1275 784
rect 1279 783 1280 787
rect 1292 786 1294 800
rect 1383 799 1384 803
rect 1388 802 1389 803
rect 1399 803 1405 804
rect 1399 802 1400 803
rect 1388 800 1400 802
rect 1388 799 1389 800
rect 1383 798 1389 799
rect 1399 799 1400 800
rect 1404 799 1405 803
rect 1399 798 1405 799
rect 1423 803 1432 804
rect 1423 799 1424 803
rect 1431 799 1432 803
rect 1423 798 1432 799
rect 1446 799 1452 800
rect 1383 795 1389 796
rect 1310 794 1316 795
rect 1310 790 1311 794
rect 1315 790 1316 794
rect 1374 794 1380 795
rect 1310 789 1316 790
rect 1319 791 1325 792
rect 1319 787 1320 791
rect 1324 787 1325 791
rect 1374 790 1375 794
rect 1379 790 1380 794
rect 1383 791 1384 795
rect 1388 794 1389 795
rect 1402 795 1408 796
rect 1446 795 1447 799
rect 1451 795 1452 799
rect 1402 794 1403 795
rect 1388 792 1403 794
rect 1388 791 1389 792
rect 1383 790 1389 791
rect 1402 791 1403 792
rect 1407 791 1408 795
rect 1402 790 1408 791
rect 1414 794 1420 795
rect 1446 794 1452 795
rect 1414 790 1415 794
rect 1419 790 1420 794
rect 1374 789 1380 790
rect 1414 789 1420 790
rect 1423 791 1429 792
rect 1319 786 1325 787
rect 1399 787 1405 788
rect 1292 784 1323 786
rect 1274 782 1280 783
rect 1399 783 1400 787
rect 1404 786 1405 787
rect 1423 787 1424 791
rect 1428 787 1429 791
rect 1423 786 1429 787
rect 1404 784 1427 786
rect 1404 783 1405 784
rect 1399 782 1405 783
rect 1184 780 1226 782
rect 1155 779 1156 780
rect 1423 779 1432 780
rect 958 778 964 779
rect 958 774 959 778
rect 963 774 964 778
rect 967 775 968 779
rect 972 775 973 779
rect 967 774 973 775
rect 990 778 996 779
rect 1007 778 1013 779
rect 1022 778 1028 779
rect 990 774 991 778
rect 995 774 996 778
rect 958 773 964 774
rect 990 773 996 774
rect 999 775 1008 776
rect 999 771 1000 775
rect 1007 771 1008 775
rect 1022 774 1023 778
rect 1027 774 1028 778
rect 1054 778 1060 779
rect 1022 773 1028 774
rect 1031 775 1037 776
rect 999 770 1008 771
rect 1031 771 1032 775
rect 1036 771 1037 775
rect 1054 774 1055 778
rect 1059 774 1060 778
rect 1086 778 1092 779
rect 1054 773 1060 774
rect 1063 775 1069 776
rect 1031 770 1037 771
rect 1063 771 1064 775
rect 1068 771 1069 775
rect 1086 774 1087 778
rect 1091 774 1092 778
rect 1126 778 1132 779
rect 1150 778 1156 779
rect 1174 778 1180 779
rect 1086 773 1092 774
rect 1095 775 1101 776
rect 1063 770 1069 771
rect 1095 771 1096 775
rect 1100 771 1101 775
rect 1126 774 1127 778
rect 1131 774 1132 778
rect 1126 773 1132 774
rect 1135 775 1141 776
rect 1095 770 1101 771
rect 1135 771 1136 775
rect 1140 771 1141 775
rect 1174 774 1175 778
rect 1179 774 1180 778
rect 1230 778 1236 779
rect 1174 773 1180 774
rect 1183 775 1189 776
rect 1135 770 1141 771
rect 1183 771 1184 775
rect 1188 771 1189 775
rect 1230 774 1231 778
rect 1235 774 1236 778
rect 1294 778 1300 779
rect 1230 773 1236 774
rect 1239 775 1245 776
rect 1183 770 1189 771
rect 1239 771 1240 775
rect 1244 771 1245 775
rect 1294 774 1295 778
rect 1299 774 1300 778
rect 1366 778 1372 779
rect 1294 773 1300 774
rect 1303 775 1309 776
rect 1239 770 1245 771
rect 1303 771 1304 775
rect 1308 771 1309 775
rect 1366 774 1367 778
rect 1371 774 1372 778
rect 1414 778 1420 779
rect 1366 773 1372 774
rect 1375 775 1381 776
rect 1303 770 1309 771
rect 1375 771 1376 775
rect 1380 771 1381 775
rect 1414 774 1415 778
rect 1419 774 1420 778
rect 1423 775 1424 779
rect 1431 775 1432 779
rect 1423 774 1432 775
rect 1414 773 1420 774
rect 1446 773 1452 774
rect 1375 770 1381 771
rect 967 767 973 768
rect 967 766 968 767
rect 944 764 968 766
rect 967 763 968 764
rect 972 763 973 767
rect 967 762 973 763
rect 999 767 1005 768
rect 999 763 1000 767
rect 1004 766 1005 767
rect 1032 766 1034 770
rect 1004 764 1034 766
rect 1004 763 1005 764
rect 999 762 1005 763
rect 1064 762 1066 770
rect 1096 762 1098 770
rect 1136 762 1138 770
rect 1184 762 1186 770
rect 1241 762 1243 770
rect 1304 762 1306 770
rect 1377 766 1379 770
rect 1446 769 1447 773
rect 1451 769 1452 773
rect 1446 768 1452 769
rect 1423 767 1429 768
rect 1423 766 1424 767
rect 1377 764 1424 766
rect 1423 763 1424 764
rect 1428 763 1429 767
rect 1423 762 1429 763
rect 636 760 681 762
rect 908 760 930 762
rect 1048 760 1066 762
rect 1080 760 1098 762
rect 1116 760 1138 762
rect 1159 760 1186 762
rect 1212 760 1243 762
rect 1272 760 1306 762
rect 636 759 637 760
rect 631 758 637 759
rect 887 759 893 760
rect 559 754 565 755
rect 887 755 888 759
rect 892 758 893 759
rect 908 758 910 760
rect 892 756 910 758
rect 1031 759 1037 760
rect 892 755 893 756
rect 887 754 893 755
rect 927 755 933 756
rect 110 750 116 751
rect 134 752 140 753
rect 158 752 164 753
rect 134 748 135 752
rect 139 748 140 752
rect 134 747 140 748
rect 143 751 152 752
rect 143 747 144 751
rect 151 747 152 751
rect 158 748 159 752
rect 163 748 164 752
rect 158 747 164 748
rect 182 752 188 753
rect 182 748 183 752
rect 187 748 188 752
rect 182 747 188 748
rect 222 752 228 753
rect 222 748 223 752
rect 227 748 228 752
rect 222 747 228 748
rect 278 752 284 753
rect 278 748 279 752
rect 283 748 284 752
rect 278 747 284 748
rect 342 752 348 753
rect 342 748 343 752
rect 347 748 348 752
rect 342 747 348 748
rect 406 752 412 753
rect 406 748 407 752
rect 411 748 412 752
rect 406 747 412 748
rect 462 752 468 753
rect 462 748 463 752
rect 467 748 468 752
rect 462 747 468 748
rect 518 752 524 753
rect 518 748 519 752
rect 523 748 524 752
rect 518 747 524 748
rect 574 752 580 753
rect 574 748 575 752
rect 579 748 580 752
rect 574 747 580 748
rect 622 752 628 753
rect 622 748 623 752
rect 627 748 628 752
rect 622 747 628 748
rect 670 752 676 753
rect 718 752 724 753
rect 670 748 671 752
rect 675 748 676 752
rect 670 747 676 748
rect 679 751 685 752
rect 679 747 680 751
rect 684 750 685 751
rect 684 748 706 750
rect 684 747 685 748
rect 143 746 152 747
rect 679 746 685 747
rect 126 743 132 744
rect 126 739 127 743
rect 131 742 132 743
rect 510 743 516 744
rect 131 740 386 742
rect 131 739 132 740
rect 126 738 132 739
rect 134 736 140 737
rect 110 733 116 734
rect 110 729 111 733
rect 115 729 116 733
rect 134 732 135 736
rect 139 732 140 736
rect 134 731 140 732
rect 158 736 164 737
rect 158 732 159 736
rect 163 732 164 736
rect 158 731 164 732
rect 182 736 188 737
rect 182 732 183 736
rect 187 732 188 736
rect 182 731 188 732
rect 214 736 220 737
rect 214 732 215 736
rect 219 732 220 736
rect 214 731 220 732
rect 262 736 268 737
rect 262 732 263 736
rect 267 732 268 736
rect 262 731 268 732
rect 318 736 324 737
rect 318 732 319 736
rect 323 732 324 736
rect 318 731 324 732
rect 374 736 380 737
rect 384 736 386 740
rect 510 739 511 743
rect 515 742 516 743
rect 704 742 706 748
rect 718 748 719 752
rect 723 748 724 752
rect 718 747 724 748
rect 758 752 764 753
rect 798 752 804 753
rect 758 748 759 752
rect 763 748 764 752
rect 758 747 764 748
rect 767 751 776 752
rect 767 747 768 751
rect 775 747 776 751
rect 798 748 799 752
rect 803 748 804 752
rect 798 747 804 748
rect 838 752 844 753
rect 838 748 839 752
rect 843 748 844 752
rect 838 747 844 748
rect 878 752 884 753
rect 878 748 879 752
rect 883 748 884 752
rect 878 747 884 748
rect 918 752 924 753
rect 918 748 919 752
rect 923 748 924 752
rect 927 751 928 755
rect 932 754 933 755
rect 950 755 956 756
rect 950 754 951 755
rect 932 752 951 754
rect 932 751 933 752
rect 927 750 933 751
rect 950 751 951 752
rect 955 751 956 755
rect 1031 755 1032 759
rect 1036 758 1037 759
rect 1048 758 1050 760
rect 1036 756 1050 758
rect 1036 755 1037 756
rect 1031 754 1037 755
rect 1063 755 1069 756
rect 950 750 956 751
rect 958 752 964 753
rect 918 747 924 748
rect 958 748 959 752
rect 963 748 964 752
rect 958 747 964 748
rect 990 752 996 753
rect 990 748 991 752
rect 995 748 996 752
rect 990 747 996 748
rect 1022 752 1028 753
rect 1022 748 1023 752
rect 1027 748 1028 752
rect 1022 747 1028 748
rect 1054 752 1060 753
rect 1054 748 1055 752
rect 1059 748 1060 752
rect 1063 751 1064 755
rect 1068 754 1069 755
rect 1080 754 1082 760
rect 1068 752 1082 754
rect 1095 755 1101 756
rect 1086 752 1092 753
rect 1068 751 1069 752
rect 1063 750 1069 751
rect 1054 747 1060 748
rect 1086 748 1087 752
rect 1091 748 1092 752
rect 1095 751 1096 755
rect 1100 754 1101 755
rect 1116 754 1118 760
rect 1100 752 1118 754
rect 1135 755 1141 756
rect 1126 752 1132 753
rect 1100 751 1101 752
rect 1095 750 1101 751
rect 1086 747 1092 748
rect 1126 748 1127 752
rect 1131 748 1132 752
rect 1135 751 1136 755
rect 1140 754 1141 755
rect 1159 754 1161 760
rect 1140 752 1161 754
rect 1183 755 1189 756
rect 1174 752 1180 753
rect 1140 751 1141 752
rect 1135 750 1141 751
rect 1126 747 1132 748
rect 1174 748 1175 752
rect 1179 748 1180 752
rect 1183 751 1184 755
rect 1188 754 1189 755
rect 1212 754 1214 760
rect 1188 752 1214 754
rect 1239 755 1245 756
rect 1230 752 1236 753
rect 1188 751 1189 752
rect 1183 750 1189 751
rect 1174 747 1180 748
rect 1230 748 1231 752
rect 1235 748 1236 752
rect 1239 751 1240 755
rect 1244 754 1245 755
rect 1272 754 1274 760
rect 1244 752 1274 754
rect 1446 755 1452 756
rect 1294 752 1300 753
rect 1366 752 1372 753
rect 1414 752 1420 753
rect 1244 751 1245 752
rect 1239 750 1245 751
rect 1230 747 1236 748
rect 1294 748 1295 752
rect 1299 748 1300 752
rect 1294 747 1300 748
rect 1303 751 1309 752
rect 1303 747 1304 751
rect 1308 747 1309 751
rect 1366 748 1367 752
rect 1371 748 1372 752
rect 1375 751 1381 752
rect 1375 748 1376 751
rect 1366 747 1372 748
rect 1374 747 1376 748
rect 1380 747 1381 751
rect 1414 748 1415 752
rect 1419 748 1420 752
rect 1446 751 1447 755
rect 1451 751 1452 755
rect 1446 750 1452 751
rect 1414 747 1420 748
rect 767 746 776 747
rect 1303 746 1309 747
rect 735 743 741 744
rect 735 742 736 743
rect 515 740 674 742
rect 704 740 736 742
rect 515 739 516 740
rect 510 738 516 739
rect 422 736 428 737
rect 374 732 375 736
rect 379 732 380 736
rect 374 731 380 732
rect 383 735 389 736
rect 383 731 384 735
rect 388 731 389 735
rect 422 732 423 736
rect 427 732 428 736
rect 422 731 428 732
rect 470 736 476 737
rect 470 732 471 736
rect 475 732 476 736
rect 470 731 476 732
rect 518 736 524 737
rect 518 732 519 736
rect 523 732 524 736
rect 518 731 524 732
rect 566 736 572 737
rect 566 732 567 736
rect 571 732 572 736
rect 566 731 572 732
rect 614 736 620 737
rect 614 732 615 736
rect 619 732 620 736
rect 614 731 620 732
rect 662 736 668 737
rect 672 736 674 740
rect 735 739 736 740
rect 740 739 741 743
rect 735 738 741 739
rect 862 743 868 744
rect 862 739 863 743
rect 867 742 868 743
rect 991 743 997 744
rect 991 742 992 743
rect 867 740 992 742
rect 867 739 868 740
rect 862 738 868 739
rect 991 739 992 740
rect 996 739 997 743
rect 991 738 997 739
rect 1002 743 1008 744
rect 1002 739 1003 743
rect 1007 742 1008 743
rect 1102 743 1108 744
rect 1102 742 1103 743
rect 1007 740 1103 742
rect 1007 739 1008 740
rect 1002 738 1008 739
rect 1102 739 1103 740
rect 1107 739 1108 743
rect 1102 738 1108 739
rect 1158 743 1164 744
rect 1158 739 1159 743
rect 1163 742 1164 743
rect 1304 742 1306 746
rect 1374 743 1375 747
rect 1379 746 1381 747
rect 1379 743 1380 746
rect 1374 742 1380 743
rect 1163 740 1306 742
rect 1163 739 1164 740
rect 1158 738 1164 739
rect 702 736 708 737
rect 662 732 663 736
rect 667 732 668 736
rect 662 731 668 732
rect 671 735 677 736
rect 671 731 672 735
rect 676 731 677 735
rect 702 732 703 736
rect 707 732 708 736
rect 702 731 708 732
rect 750 736 756 737
rect 750 732 751 736
rect 755 732 756 736
rect 750 731 756 732
rect 806 736 812 737
rect 806 732 807 736
rect 811 732 812 736
rect 806 731 812 732
rect 870 736 876 737
rect 870 732 871 736
rect 875 732 876 736
rect 870 731 876 732
rect 942 736 948 737
rect 942 732 943 736
rect 947 732 948 736
rect 942 731 948 732
rect 1014 736 1020 737
rect 1014 732 1015 736
rect 1019 732 1020 736
rect 1014 731 1020 732
rect 1086 736 1092 737
rect 1086 732 1087 736
rect 1091 732 1092 736
rect 1086 731 1092 732
rect 1150 736 1156 737
rect 1150 732 1151 736
rect 1155 732 1156 736
rect 1150 731 1156 732
rect 1214 736 1220 737
rect 1214 732 1215 736
rect 1219 732 1220 736
rect 1214 731 1220 732
rect 1270 736 1276 737
rect 1270 732 1271 736
rect 1275 732 1276 736
rect 1270 731 1276 732
rect 1326 736 1332 737
rect 1326 732 1327 736
rect 1331 732 1332 736
rect 1326 731 1332 732
rect 1382 736 1388 737
rect 1382 732 1383 736
rect 1387 732 1388 736
rect 1382 731 1388 732
rect 1414 736 1420 737
rect 1414 732 1415 736
rect 1419 732 1420 736
rect 1414 731 1420 732
rect 1446 733 1452 734
rect 383 730 389 731
rect 671 730 677 731
rect 110 728 116 729
rect 1446 729 1447 733
rect 1451 729 1452 733
rect 1446 728 1452 729
rect 143 727 149 728
rect 143 723 144 727
rect 148 726 149 727
rect 170 727 176 728
rect 170 726 171 727
rect 148 724 171 726
rect 148 723 149 724
rect 143 722 149 723
rect 170 723 171 724
rect 175 723 176 727
rect 170 722 176 723
rect 191 727 197 728
rect 191 723 192 727
rect 196 726 197 727
rect 226 727 232 728
rect 226 726 227 727
rect 196 724 227 726
rect 196 723 197 724
rect 191 722 197 723
rect 226 723 227 724
rect 231 723 232 727
rect 226 722 232 723
rect 271 727 277 728
rect 271 723 272 727
rect 276 726 277 727
rect 330 727 336 728
rect 330 726 331 727
rect 276 724 331 726
rect 276 723 277 724
rect 271 722 277 723
rect 330 723 331 724
rect 335 723 336 727
rect 330 722 336 723
rect 431 727 437 728
rect 431 723 432 727
rect 436 726 437 727
rect 482 727 488 728
rect 482 726 483 727
rect 436 724 483 726
rect 436 723 437 724
rect 431 722 437 723
rect 482 723 483 724
rect 487 723 488 727
rect 482 722 488 723
rect 527 727 533 728
rect 527 723 528 727
rect 532 726 533 727
rect 578 727 584 728
rect 578 726 579 727
rect 532 724 579 726
rect 532 723 533 724
rect 527 722 533 723
rect 578 723 579 724
rect 583 723 584 727
rect 578 722 584 723
rect 623 727 629 728
rect 623 723 624 727
rect 628 726 629 727
rect 674 727 680 728
rect 674 726 675 727
rect 628 724 675 726
rect 628 723 629 724
rect 623 722 629 723
rect 674 723 675 724
rect 679 723 680 727
rect 674 722 680 723
rect 815 727 821 728
rect 815 723 816 727
rect 820 726 821 727
rect 882 727 888 728
rect 882 726 883 727
rect 820 724 883 726
rect 820 723 821 724
rect 815 722 821 723
rect 882 723 883 724
rect 887 723 888 727
rect 882 722 888 723
rect 951 727 957 728
rect 951 723 952 727
rect 956 726 957 727
rect 1026 727 1032 728
rect 1026 726 1027 727
rect 956 724 1027 726
rect 956 723 957 724
rect 951 722 957 723
rect 1026 723 1027 724
rect 1031 723 1032 727
rect 1026 722 1032 723
rect 1050 727 1056 728
rect 1050 723 1051 727
rect 1055 726 1056 727
rect 1095 727 1101 728
rect 1095 726 1096 727
rect 1055 724 1096 726
rect 1055 723 1056 724
rect 1050 722 1056 723
rect 1095 723 1096 724
rect 1100 723 1101 727
rect 1095 722 1101 723
rect 1159 727 1165 728
rect 1159 723 1160 727
rect 1164 726 1165 727
rect 1290 727 1296 728
rect 1290 726 1291 727
rect 1164 724 1291 726
rect 1164 723 1165 724
rect 1159 722 1165 723
rect 1290 723 1291 724
rect 1295 723 1296 727
rect 1290 722 1296 723
rect 167 719 173 720
rect 110 715 116 716
rect 110 711 111 715
rect 115 711 116 715
rect 167 715 168 719
rect 172 718 173 719
rect 175 719 181 720
rect 175 718 176 719
rect 172 716 176 718
rect 172 715 173 716
rect 167 714 173 715
rect 175 715 176 716
rect 180 715 181 719
rect 175 714 181 715
rect 223 719 229 720
rect 223 715 224 719
rect 228 718 229 719
rect 327 719 333 720
rect 228 716 274 718
rect 228 715 229 716
rect 223 714 229 715
rect 272 712 274 716
rect 327 715 328 719
rect 332 718 333 719
rect 479 719 485 720
rect 332 716 358 718
rect 332 715 333 716
rect 327 714 333 715
rect 143 711 152 712
rect 167 711 176 712
rect 223 711 232 712
rect 271 711 277 712
rect 327 711 336 712
rect 110 710 116 711
rect 134 710 140 711
rect 134 706 135 710
rect 139 706 140 710
rect 143 707 144 711
rect 151 707 152 711
rect 143 706 152 707
rect 158 710 164 711
rect 158 706 159 710
rect 163 706 164 710
rect 167 707 168 711
rect 175 707 176 711
rect 167 706 176 707
rect 182 710 188 711
rect 182 706 183 710
rect 187 706 188 710
rect 214 710 220 711
rect 134 705 140 706
rect 158 705 164 706
rect 182 705 188 706
rect 191 707 197 708
rect 126 703 132 704
rect 126 699 127 703
rect 131 702 132 703
rect 191 703 192 707
rect 196 703 197 707
rect 214 706 215 710
rect 219 706 220 710
rect 223 707 224 711
rect 231 707 232 711
rect 223 706 232 707
rect 262 710 268 711
rect 262 706 263 710
rect 267 706 268 710
rect 271 707 272 711
rect 276 707 277 711
rect 271 706 277 707
rect 318 710 324 711
rect 318 706 319 710
rect 323 706 324 710
rect 327 707 328 711
rect 335 707 336 711
rect 327 706 336 707
rect 214 705 220 706
rect 262 705 268 706
rect 318 705 324 706
rect 191 702 197 703
rect 356 702 358 716
rect 479 715 480 719
rect 484 718 485 719
rect 575 719 581 720
rect 484 716 515 718
rect 484 715 485 716
rect 479 714 485 715
rect 479 711 488 712
rect 374 710 380 711
rect 374 706 375 710
rect 379 706 380 710
rect 422 710 428 711
rect 374 705 380 706
rect 383 707 389 708
rect 383 703 384 707
rect 388 703 389 707
rect 422 706 423 710
rect 427 706 428 710
rect 470 710 476 711
rect 422 705 428 706
rect 431 707 437 708
rect 383 702 389 703
rect 431 703 432 707
rect 436 706 437 707
rect 470 706 471 710
rect 475 706 476 710
rect 479 707 480 711
rect 487 707 488 711
rect 479 706 488 707
rect 436 704 466 706
rect 470 705 476 706
rect 436 703 437 704
rect 431 702 437 703
rect 464 702 466 704
rect 494 703 500 704
rect 494 702 495 703
rect 131 700 147 702
rect 131 699 132 700
rect 126 698 132 699
rect 145 696 147 700
rect 175 699 181 700
rect 143 695 149 696
rect 175 695 176 699
rect 180 698 181 699
rect 192 698 194 702
rect 356 700 386 702
rect 464 700 495 702
rect 494 699 495 700
rect 499 699 500 703
rect 513 702 515 716
rect 575 715 576 719
rect 580 718 581 719
rect 711 719 717 720
rect 580 716 602 718
rect 580 715 581 716
rect 575 714 581 715
rect 575 711 584 712
rect 518 710 524 711
rect 518 706 519 710
rect 523 706 524 710
rect 566 710 572 711
rect 518 705 524 706
rect 527 707 533 708
rect 527 703 528 707
rect 532 703 533 707
rect 566 706 567 710
rect 571 706 572 710
rect 575 707 576 711
rect 583 707 584 711
rect 575 706 584 707
rect 566 705 572 706
rect 527 702 533 703
rect 600 702 602 716
rect 711 715 712 719
rect 716 718 717 719
rect 727 719 733 720
rect 727 718 728 719
rect 716 716 728 718
rect 716 715 717 716
rect 711 714 717 715
rect 727 715 728 716
rect 732 715 733 719
rect 759 719 765 720
rect 759 718 760 719
rect 727 714 733 715
rect 736 716 760 718
rect 671 711 680 712
rect 711 711 717 712
rect 614 710 620 711
rect 614 706 615 710
rect 619 706 620 710
rect 662 710 668 711
rect 614 705 620 706
rect 623 707 629 708
rect 623 703 624 707
rect 628 703 629 707
rect 662 706 663 710
rect 667 706 668 710
rect 671 707 672 711
rect 679 707 680 711
rect 671 706 680 707
rect 702 710 708 711
rect 702 706 703 710
rect 707 706 708 710
rect 711 707 712 711
rect 716 710 717 711
rect 736 710 738 716
rect 759 715 760 716
rect 764 715 765 719
rect 759 714 765 715
rect 879 719 885 720
rect 879 715 880 719
rect 884 718 885 719
rect 1023 719 1029 720
rect 884 716 918 718
rect 884 715 885 716
rect 879 714 885 715
rect 759 711 765 712
rect 716 708 738 710
rect 750 710 756 711
rect 716 707 717 708
rect 711 706 717 707
rect 750 706 751 710
rect 755 706 756 710
rect 759 707 760 711
rect 764 710 765 711
rect 770 711 776 712
rect 879 711 888 712
rect 770 710 771 711
rect 764 708 771 710
rect 764 707 765 708
rect 759 706 765 707
rect 770 707 771 708
rect 775 707 776 711
rect 770 706 776 707
rect 806 710 812 711
rect 806 706 807 710
rect 811 706 812 710
rect 870 710 876 711
rect 662 705 668 706
rect 702 705 708 706
rect 750 705 756 706
rect 806 705 812 706
rect 815 707 821 708
rect 623 702 629 703
rect 727 703 733 704
rect 513 700 530 702
rect 600 700 626 702
rect 494 698 500 699
rect 727 699 728 703
rect 732 702 733 703
rect 815 703 816 707
rect 820 706 821 707
rect 838 707 844 708
rect 838 706 839 707
rect 820 704 839 706
rect 820 703 821 704
rect 815 702 821 703
rect 838 703 839 704
rect 843 703 844 707
rect 870 706 871 710
rect 875 706 876 710
rect 879 707 880 711
rect 887 707 888 711
rect 879 706 888 707
rect 870 705 876 706
rect 838 702 844 703
rect 846 703 852 704
rect 732 700 770 702
rect 732 699 733 700
rect 727 698 733 699
rect 180 696 194 698
rect 768 696 770 700
rect 846 699 847 703
rect 851 702 852 703
rect 916 702 918 716
rect 1023 715 1024 719
rect 1028 718 1029 719
rect 1223 719 1229 720
rect 1223 718 1224 719
rect 1028 716 1062 718
rect 1028 715 1029 716
rect 1023 714 1029 715
rect 1023 711 1032 712
rect 942 710 948 711
rect 942 706 943 710
rect 947 706 948 710
rect 1014 710 1020 711
rect 942 705 948 706
rect 951 707 957 708
rect 951 703 952 707
rect 956 703 957 707
rect 1014 706 1015 710
rect 1019 706 1020 710
rect 1023 707 1024 711
rect 1031 707 1032 711
rect 1023 706 1032 707
rect 1014 705 1020 706
rect 951 702 957 703
rect 991 703 997 704
rect 851 700 914 702
rect 916 700 954 702
rect 960 700 978 702
rect 851 699 852 700
rect 846 698 852 699
rect 912 698 914 700
rect 960 698 962 700
rect 912 696 962 698
rect 976 696 978 700
rect 991 699 992 703
rect 996 702 997 703
rect 1050 703 1056 704
rect 1050 702 1051 703
rect 996 700 1051 702
rect 996 699 997 700
rect 991 698 997 699
rect 1050 699 1051 700
rect 1055 699 1056 703
rect 1060 702 1062 716
rect 1193 716 1224 718
rect 1159 711 1165 712
rect 1086 710 1092 711
rect 1086 706 1087 710
rect 1091 706 1092 710
rect 1150 710 1156 711
rect 1086 705 1092 706
rect 1095 707 1101 708
rect 1095 703 1096 707
rect 1100 703 1101 707
rect 1150 706 1151 710
rect 1155 706 1156 710
rect 1159 707 1160 711
rect 1164 710 1165 711
rect 1193 710 1195 716
rect 1223 715 1224 716
rect 1228 715 1229 719
rect 1279 719 1285 720
rect 1279 718 1280 719
rect 1223 714 1229 715
rect 1252 716 1280 718
rect 1223 711 1229 712
rect 1164 708 1195 710
rect 1214 710 1220 711
rect 1164 707 1165 708
rect 1159 706 1165 707
rect 1214 706 1215 710
rect 1219 706 1220 710
rect 1223 707 1224 711
rect 1228 710 1229 711
rect 1252 710 1254 716
rect 1279 715 1280 716
rect 1284 715 1285 719
rect 1279 714 1285 715
rect 1335 719 1341 720
rect 1335 715 1336 719
rect 1340 718 1341 719
rect 1367 719 1373 720
rect 1367 718 1368 719
rect 1340 716 1368 718
rect 1340 715 1341 716
rect 1335 714 1341 715
rect 1367 715 1368 716
rect 1372 715 1373 719
rect 1367 714 1373 715
rect 1391 719 1397 720
rect 1391 715 1392 719
rect 1396 715 1397 719
rect 1391 714 1397 715
rect 1423 719 1432 720
rect 1423 715 1424 719
rect 1431 715 1432 719
rect 1423 714 1432 715
rect 1446 715 1452 716
rect 1393 712 1410 714
rect 1335 711 1341 712
rect 1228 708 1254 710
rect 1270 710 1276 711
rect 1228 707 1229 708
rect 1223 706 1229 707
rect 1270 706 1271 710
rect 1275 706 1276 710
rect 1326 710 1332 711
rect 1150 705 1156 706
rect 1214 705 1220 706
rect 1270 705 1276 706
rect 1279 707 1285 708
rect 1095 702 1101 703
rect 1279 703 1280 707
rect 1284 706 1285 707
rect 1303 707 1309 708
rect 1303 706 1304 707
rect 1284 704 1304 706
rect 1284 703 1285 704
rect 1279 702 1285 703
rect 1303 703 1304 704
rect 1308 703 1309 707
rect 1326 706 1327 710
rect 1331 706 1332 710
rect 1335 707 1336 711
rect 1340 710 1341 711
rect 1374 711 1380 712
rect 1374 710 1375 711
rect 1340 708 1375 710
rect 1340 707 1341 708
rect 1335 706 1341 707
rect 1374 707 1375 708
rect 1379 707 1380 711
rect 1374 706 1380 707
rect 1382 710 1388 711
rect 1382 706 1383 710
rect 1387 706 1388 710
rect 1326 705 1332 706
rect 1382 705 1388 706
rect 1391 707 1397 708
rect 1303 702 1309 703
rect 1367 703 1373 704
rect 1060 700 1098 702
rect 1050 698 1056 699
rect 1367 699 1368 703
rect 1372 702 1373 703
rect 1391 703 1392 707
rect 1396 703 1397 707
rect 1391 702 1397 703
rect 1408 702 1410 712
rect 1446 711 1447 715
rect 1451 711 1452 715
rect 1414 710 1420 711
rect 1446 710 1452 711
rect 1414 706 1415 710
rect 1419 706 1420 710
rect 1414 705 1420 706
rect 1423 707 1429 708
rect 1423 703 1424 707
rect 1428 703 1429 707
rect 1423 702 1429 703
rect 1372 700 1395 702
rect 1408 700 1427 702
rect 1372 699 1373 700
rect 1367 698 1373 699
rect 180 695 181 696
rect 767 695 773 696
rect 975 695 981 696
rect 1287 695 1296 696
rect 1423 695 1432 696
rect 134 694 140 695
rect 134 690 135 694
rect 139 690 140 694
rect 143 691 144 695
rect 148 691 149 695
rect 143 690 149 691
rect 158 694 164 695
rect 175 694 181 695
rect 198 694 204 695
rect 158 690 159 694
rect 163 690 164 694
rect 110 689 116 690
rect 134 689 140 690
rect 158 689 164 690
rect 167 691 173 692
rect 110 685 111 689
rect 115 685 116 689
rect 167 687 168 691
rect 172 687 173 691
rect 198 690 199 694
rect 203 690 204 694
rect 238 694 244 695
rect 198 689 204 690
rect 207 691 213 692
rect 167 686 173 687
rect 207 687 208 691
rect 212 687 213 691
rect 238 690 239 694
rect 243 690 244 694
rect 286 694 292 695
rect 238 689 244 690
rect 247 691 253 692
rect 207 686 213 687
rect 247 687 248 691
rect 252 687 253 691
rect 286 690 287 694
rect 291 690 292 694
rect 334 694 340 695
rect 286 689 292 690
rect 295 691 301 692
rect 247 686 253 687
rect 295 687 296 691
rect 300 687 301 691
rect 334 690 335 694
rect 339 690 340 694
rect 390 694 396 695
rect 334 689 340 690
rect 343 691 349 692
rect 295 686 301 687
rect 343 687 344 691
rect 348 687 349 691
rect 390 690 391 694
rect 395 690 396 694
rect 438 694 444 695
rect 390 689 396 690
rect 399 691 405 692
rect 343 686 349 687
rect 399 687 400 691
rect 404 690 405 691
rect 430 691 436 692
rect 430 690 431 691
rect 404 688 431 690
rect 404 687 405 688
rect 399 686 405 687
rect 430 687 431 688
rect 435 687 436 691
rect 438 690 439 694
rect 443 690 444 694
rect 486 694 492 695
rect 438 689 444 690
rect 447 691 456 692
rect 430 686 436 687
rect 447 687 448 691
rect 455 687 456 691
rect 486 690 487 694
rect 491 690 492 694
rect 534 694 540 695
rect 486 689 492 690
rect 495 691 501 692
rect 447 686 456 687
rect 495 687 496 691
rect 500 687 501 691
rect 534 690 535 694
rect 539 690 540 694
rect 582 694 588 695
rect 534 689 540 690
rect 543 691 549 692
rect 495 686 501 687
rect 543 687 544 691
rect 548 687 549 691
rect 582 690 583 694
rect 587 690 588 694
rect 638 694 644 695
rect 582 689 588 690
rect 591 691 597 692
rect 543 686 549 687
rect 591 687 592 691
rect 596 687 597 691
rect 638 690 639 694
rect 643 690 644 694
rect 694 694 700 695
rect 638 689 644 690
rect 647 691 653 692
rect 591 686 597 687
rect 647 687 648 691
rect 652 690 653 691
rect 694 690 695 694
rect 699 690 700 694
rect 758 694 764 695
rect 652 688 681 690
rect 694 689 700 690
rect 703 691 709 692
rect 652 687 653 688
rect 647 686 653 687
rect 110 684 116 685
rect 143 683 149 684
rect 143 679 144 683
rect 148 682 149 683
rect 169 682 171 686
rect 148 680 171 682
rect 148 679 149 680
rect 143 678 149 679
rect 209 678 211 686
rect 248 678 250 686
rect 296 678 298 686
rect 345 682 347 686
rect 169 676 211 678
rect 228 676 250 678
rect 272 676 298 678
rect 320 680 347 682
rect 399 683 405 684
rect 167 675 173 676
rect 110 671 116 672
rect 110 667 111 671
rect 115 667 116 671
rect 167 671 168 675
rect 172 671 173 675
rect 167 670 173 671
rect 207 671 213 672
rect 110 666 116 667
rect 134 668 140 669
rect 134 664 135 668
rect 139 664 140 668
rect 134 663 140 664
rect 158 668 164 669
rect 158 664 159 668
rect 163 664 164 668
rect 158 663 164 664
rect 198 668 204 669
rect 198 664 199 668
rect 203 664 204 668
rect 207 667 208 671
rect 212 670 213 671
rect 228 670 230 676
rect 212 668 230 670
rect 247 671 253 672
rect 238 668 244 669
rect 212 667 213 668
rect 207 666 213 667
rect 198 663 204 664
rect 238 664 239 668
rect 243 664 244 668
rect 247 667 248 671
rect 252 670 253 671
rect 272 670 274 676
rect 252 668 274 670
rect 295 671 301 672
rect 286 668 292 669
rect 252 667 253 668
rect 247 666 253 667
rect 238 663 244 664
rect 286 664 287 668
rect 291 664 292 668
rect 295 667 296 671
rect 300 670 301 671
rect 320 670 322 680
rect 399 679 400 683
rect 404 682 405 683
rect 438 683 444 684
rect 438 682 439 683
rect 404 680 439 682
rect 404 679 405 680
rect 399 678 405 679
rect 438 679 439 680
rect 443 679 444 683
rect 438 678 444 679
rect 447 683 453 684
rect 447 679 448 683
rect 452 682 453 683
rect 497 682 499 686
rect 545 682 547 686
rect 593 682 595 686
rect 452 680 499 682
rect 520 680 547 682
rect 568 680 595 682
rect 679 682 681 688
rect 703 687 704 691
rect 708 690 709 691
rect 758 690 759 694
rect 763 690 764 694
rect 767 691 768 695
rect 772 691 773 695
rect 767 690 773 691
rect 830 694 836 695
rect 830 690 831 694
rect 835 690 836 694
rect 902 694 908 695
rect 708 688 738 690
rect 758 689 764 690
rect 830 689 836 690
rect 839 691 845 692
rect 708 687 709 688
rect 703 686 709 687
rect 703 683 709 684
rect 703 682 704 683
rect 679 680 704 682
rect 452 679 453 680
rect 447 678 453 679
rect 300 668 322 670
rect 495 671 501 672
rect 334 668 340 669
rect 390 668 396 669
rect 300 667 301 668
rect 295 666 301 667
rect 286 663 292 664
rect 334 664 335 668
rect 339 664 340 668
rect 334 663 340 664
rect 343 667 352 668
rect 343 663 344 667
rect 351 663 352 667
rect 390 664 391 668
rect 395 664 396 668
rect 390 663 396 664
rect 438 668 444 669
rect 438 664 439 668
rect 443 664 444 668
rect 438 663 444 664
rect 486 668 492 669
rect 486 664 487 668
rect 491 664 492 668
rect 495 667 496 671
rect 500 670 501 671
rect 520 670 522 680
rect 500 668 522 670
rect 543 671 549 672
rect 534 668 540 669
rect 500 667 501 668
rect 495 666 501 667
rect 534 664 535 668
rect 539 664 540 668
rect 543 667 544 671
rect 548 670 549 671
rect 568 670 570 680
rect 703 679 704 680
rect 708 679 709 683
rect 736 682 738 688
rect 839 687 840 691
rect 844 690 845 691
rect 902 690 903 694
rect 907 690 908 694
rect 966 694 972 695
rect 844 688 878 690
rect 902 689 908 690
rect 911 691 917 692
rect 844 687 845 688
rect 839 686 845 687
rect 767 683 773 684
rect 767 682 768 683
rect 736 680 768 682
rect 703 678 709 679
rect 767 679 768 680
rect 772 679 773 683
rect 767 678 773 679
rect 838 683 845 684
rect 838 679 839 683
rect 844 679 845 683
rect 876 682 878 688
rect 911 687 912 691
rect 916 690 917 691
rect 966 690 967 694
rect 971 690 972 694
rect 975 691 976 695
rect 980 691 981 695
rect 975 690 981 691
rect 1030 694 1036 695
rect 1030 690 1031 694
rect 1035 690 1036 694
rect 1086 694 1092 695
rect 916 688 946 690
rect 966 689 972 690
rect 1030 689 1036 690
rect 1039 691 1045 692
rect 916 687 917 688
rect 911 686 917 687
rect 911 683 917 684
rect 911 682 912 683
rect 876 680 912 682
rect 838 678 845 679
rect 911 679 912 680
rect 916 679 917 683
rect 944 682 946 688
rect 1039 687 1040 691
rect 1044 687 1045 691
rect 1086 690 1087 694
rect 1091 690 1092 694
rect 1134 694 1140 695
rect 1086 689 1092 690
rect 1095 691 1101 692
rect 1039 686 1045 687
rect 1095 687 1096 691
rect 1100 690 1101 691
rect 1134 690 1135 694
rect 1139 690 1140 694
rect 1174 694 1180 695
rect 1100 688 1122 690
rect 1134 689 1140 690
rect 1143 691 1149 692
rect 1100 687 1101 688
rect 1095 686 1101 687
rect 975 683 981 684
rect 975 682 976 683
rect 944 680 976 682
rect 911 678 917 679
rect 975 679 976 680
rect 980 679 981 683
rect 1041 682 1043 686
rect 1095 683 1101 684
rect 1095 682 1096 683
rect 1041 680 1096 682
rect 975 678 981 679
rect 1095 679 1096 680
rect 1100 679 1101 683
rect 1120 682 1122 688
rect 1143 687 1144 691
rect 1148 690 1149 691
rect 1174 690 1175 694
rect 1179 690 1180 694
rect 1214 694 1220 695
rect 1148 688 1161 690
rect 1174 689 1180 690
rect 1183 691 1189 692
rect 1148 687 1149 688
rect 1143 686 1149 687
rect 1143 683 1149 684
rect 1143 682 1144 683
rect 1120 680 1144 682
rect 1095 678 1101 679
rect 1143 679 1144 680
rect 1148 679 1149 683
rect 1159 682 1161 688
rect 1183 687 1184 691
rect 1188 690 1189 691
rect 1214 690 1215 694
rect 1219 690 1220 694
rect 1246 694 1252 695
rect 1188 688 1206 690
rect 1214 689 1220 690
rect 1223 691 1229 692
rect 1188 687 1189 688
rect 1183 686 1189 687
rect 1183 683 1189 684
rect 1183 682 1184 683
rect 1159 680 1184 682
rect 1143 678 1149 679
rect 1183 679 1184 680
rect 1188 679 1189 683
rect 1204 682 1206 688
rect 1223 687 1224 691
rect 1228 690 1229 691
rect 1246 690 1247 694
rect 1251 690 1252 694
rect 1278 694 1284 695
rect 1228 688 1242 690
rect 1246 689 1252 690
rect 1255 691 1261 692
rect 1228 687 1229 688
rect 1223 686 1229 687
rect 1223 683 1229 684
rect 1223 682 1224 683
rect 1204 680 1224 682
rect 1183 678 1189 679
rect 1223 679 1224 680
rect 1228 679 1229 683
rect 1223 678 1229 679
rect 1240 678 1242 688
rect 1255 687 1256 691
rect 1260 687 1261 691
rect 1278 690 1279 694
rect 1283 690 1284 694
rect 1287 691 1288 695
rect 1295 691 1296 695
rect 1287 690 1296 691
rect 1310 694 1316 695
rect 1310 690 1311 694
rect 1315 690 1316 694
rect 1342 694 1348 695
rect 1278 689 1284 690
rect 1310 689 1316 690
rect 1319 691 1325 692
rect 1255 686 1261 687
rect 1319 687 1320 691
rect 1324 687 1325 691
rect 1342 690 1343 694
rect 1347 690 1348 694
rect 1366 694 1372 695
rect 1342 689 1348 690
rect 1351 691 1360 692
rect 1319 686 1325 687
rect 1351 687 1352 691
rect 1359 687 1360 691
rect 1366 690 1367 694
rect 1371 690 1372 694
rect 1390 694 1396 695
rect 1366 689 1372 690
rect 1375 691 1381 692
rect 1351 686 1360 687
rect 1375 687 1376 691
rect 1380 687 1381 691
rect 1390 690 1391 694
rect 1395 690 1396 694
rect 1414 694 1420 695
rect 1390 689 1396 690
rect 1399 691 1405 692
rect 1375 686 1381 687
rect 1399 687 1400 691
rect 1404 687 1405 691
rect 1414 690 1415 694
rect 1419 690 1420 694
rect 1423 691 1424 695
rect 1431 691 1432 695
rect 1423 690 1432 691
rect 1414 689 1420 690
rect 1446 689 1452 690
rect 1399 686 1405 687
rect 1257 682 1259 686
rect 1287 683 1293 684
rect 1287 682 1288 683
rect 1257 680 1288 682
rect 1287 679 1288 680
rect 1292 679 1293 683
rect 1321 682 1323 686
rect 1351 683 1357 684
rect 1351 682 1352 683
rect 1321 680 1352 682
rect 1287 678 1293 679
rect 1303 679 1309 680
rect 1240 676 1259 678
rect 1255 675 1261 676
rect 1255 671 1256 675
rect 1260 671 1261 675
rect 1303 675 1304 679
rect 1308 678 1309 679
rect 1351 679 1352 680
rect 1356 679 1357 683
rect 1351 678 1357 679
rect 1377 678 1379 686
rect 1401 682 1403 686
rect 1446 685 1447 689
rect 1451 685 1452 689
rect 1446 684 1452 685
rect 1423 683 1429 684
rect 1423 682 1424 683
rect 1401 680 1424 682
rect 1423 679 1424 680
rect 1428 679 1429 683
rect 1423 678 1429 679
rect 1308 676 1323 678
rect 1377 676 1403 678
rect 1308 675 1309 676
rect 1303 674 1309 675
rect 1319 675 1325 676
rect 1255 670 1261 671
rect 1319 671 1320 675
rect 1324 671 1325 675
rect 1319 670 1325 671
rect 1399 675 1405 676
rect 1399 671 1400 675
rect 1404 671 1405 675
rect 1399 670 1405 671
rect 1446 671 1452 672
rect 548 668 570 670
rect 582 668 588 669
rect 638 668 644 669
rect 694 668 700 669
rect 548 667 549 668
rect 543 666 549 667
rect 486 663 492 664
rect 494 663 500 664
rect 534 663 540 664
rect 582 664 583 668
rect 587 664 588 668
rect 582 663 588 664
rect 591 667 597 668
rect 591 663 592 667
rect 596 663 597 667
rect 638 664 639 668
rect 643 664 644 668
rect 638 663 644 664
rect 647 667 656 668
rect 647 663 648 667
rect 655 663 656 667
rect 694 664 695 668
rect 699 664 700 668
rect 694 663 700 664
rect 758 668 764 669
rect 758 664 759 668
rect 763 664 764 668
rect 758 663 764 664
rect 830 668 836 669
rect 830 664 831 668
rect 835 664 836 668
rect 830 663 836 664
rect 902 668 908 669
rect 902 664 903 668
rect 907 664 908 668
rect 902 663 908 664
rect 966 668 972 669
rect 966 664 967 668
rect 971 664 972 668
rect 966 663 972 664
rect 1030 668 1036 669
rect 1086 668 1092 669
rect 1030 664 1031 668
rect 1035 664 1036 668
rect 1030 663 1036 664
rect 1039 667 1045 668
rect 1039 663 1040 667
rect 1044 666 1045 667
rect 1078 667 1084 668
rect 1078 666 1079 667
rect 1044 664 1079 666
rect 1044 663 1045 664
rect 343 662 352 663
rect 449 660 482 662
rect 430 659 436 660
rect 190 656 196 657
rect 110 653 116 654
rect 110 649 111 653
rect 115 649 116 653
rect 190 652 191 656
rect 195 652 196 656
rect 190 651 196 652
rect 214 656 220 657
rect 214 652 215 656
rect 219 652 220 656
rect 214 651 220 652
rect 238 656 244 657
rect 238 652 239 656
rect 243 652 244 656
rect 238 651 244 652
rect 262 656 268 657
rect 262 652 263 656
rect 267 652 268 656
rect 262 651 268 652
rect 294 656 300 657
rect 294 652 295 656
rect 299 652 300 656
rect 294 651 300 652
rect 326 656 332 657
rect 326 652 327 656
rect 331 652 332 656
rect 326 651 332 652
rect 366 656 372 657
rect 366 652 367 656
rect 371 652 372 656
rect 366 651 372 652
rect 406 656 412 657
rect 406 652 407 656
rect 411 652 412 656
rect 430 655 431 659
rect 435 658 436 659
rect 449 658 451 660
rect 435 656 451 658
rect 454 656 460 657
rect 435 655 436 656
rect 430 654 436 655
rect 406 651 412 652
rect 454 652 455 656
rect 459 652 460 656
rect 454 651 460 652
rect 110 648 116 649
rect 199 647 205 648
rect 199 643 200 647
rect 204 646 205 647
rect 226 647 232 648
rect 226 646 227 647
rect 204 644 227 646
rect 204 643 205 644
rect 199 642 205 643
rect 226 643 227 644
rect 231 643 232 647
rect 226 642 232 643
rect 247 647 253 648
rect 247 643 248 647
rect 252 646 253 647
rect 274 647 280 648
rect 274 646 275 647
rect 252 644 275 646
rect 252 643 253 644
rect 247 642 253 643
rect 274 643 275 644
rect 279 643 280 647
rect 274 642 280 643
rect 303 647 309 648
rect 303 643 304 647
rect 308 646 309 647
rect 338 647 344 648
rect 338 646 339 647
rect 308 644 339 646
rect 308 643 309 644
rect 303 642 309 643
rect 338 643 339 644
rect 343 643 344 647
rect 338 642 344 643
rect 351 647 357 648
rect 351 643 352 647
rect 356 646 357 647
rect 375 647 381 648
rect 375 646 376 647
rect 356 644 376 646
rect 356 643 357 644
rect 351 642 357 643
rect 375 643 376 644
rect 380 643 381 647
rect 375 642 381 643
rect 415 647 421 648
rect 415 643 416 647
rect 420 646 421 647
rect 466 647 472 648
rect 466 646 467 647
rect 420 644 467 646
rect 420 643 421 644
rect 415 642 421 643
rect 466 643 467 644
rect 471 643 472 647
rect 466 642 472 643
rect 480 642 482 660
rect 494 659 495 663
rect 499 662 500 663
rect 591 662 597 663
rect 647 662 656 663
rect 1039 662 1045 663
rect 1078 663 1079 664
rect 1083 663 1084 667
rect 1086 664 1087 668
rect 1091 664 1092 668
rect 1086 663 1092 664
rect 1134 668 1140 669
rect 1134 664 1135 668
rect 1139 664 1140 668
rect 1134 663 1140 664
rect 1174 668 1180 669
rect 1174 664 1175 668
rect 1179 664 1180 668
rect 1174 663 1180 664
rect 1214 668 1220 669
rect 1214 664 1215 668
rect 1219 664 1220 668
rect 1214 663 1220 664
rect 1246 668 1252 669
rect 1246 664 1247 668
rect 1251 664 1252 668
rect 1246 663 1252 664
rect 1278 668 1284 669
rect 1278 664 1279 668
rect 1283 664 1284 668
rect 1278 663 1284 664
rect 1310 668 1316 669
rect 1310 664 1311 668
rect 1315 664 1316 668
rect 1310 663 1316 664
rect 1342 668 1348 669
rect 1342 664 1343 668
rect 1347 664 1348 668
rect 1342 663 1348 664
rect 1366 668 1372 669
rect 1390 668 1396 669
rect 1366 664 1367 668
rect 1371 664 1372 668
rect 1366 663 1372 664
rect 1375 667 1381 668
rect 1375 663 1376 667
rect 1380 663 1381 667
rect 1390 664 1391 668
rect 1395 664 1396 668
rect 1390 663 1396 664
rect 1414 668 1420 669
rect 1414 664 1415 668
rect 1419 664 1420 668
rect 1446 667 1447 671
rect 1451 667 1452 671
rect 1446 666 1452 667
rect 1414 663 1420 664
rect 1078 662 1084 663
rect 1375 662 1381 663
rect 499 660 530 662
rect 499 659 500 660
rect 494 658 500 659
rect 528 658 530 660
rect 545 660 578 662
rect 545 658 547 660
rect 502 656 508 657
rect 528 656 547 658
rect 576 658 578 660
rect 593 658 595 662
rect 550 656 556 657
rect 576 656 595 658
rect 1354 659 1360 660
rect 606 656 612 657
rect 502 652 503 656
rect 507 652 508 656
rect 502 651 508 652
rect 550 652 551 656
rect 555 652 556 656
rect 550 651 556 652
rect 606 652 607 656
rect 611 652 612 656
rect 606 651 612 652
rect 662 656 668 657
rect 662 652 663 656
rect 667 652 668 656
rect 662 651 668 652
rect 718 656 724 657
rect 718 652 719 656
rect 723 652 724 656
rect 718 651 724 652
rect 766 656 772 657
rect 766 652 767 656
rect 771 652 772 656
rect 766 651 772 652
rect 814 656 820 657
rect 862 656 868 657
rect 814 652 815 656
rect 819 652 820 656
rect 814 651 820 652
rect 823 655 829 656
rect 823 651 824 655
rect 828 654 829 655
rect 846 655 852 656
rect 846 654 847 655
rect 828 652 847 654
rect 828 651 829 652
rect 823 650 829 651
rect 846 651 847 652
rect 851 651 852 655
rect 862 652 863 656
rect 867 652 868 656
rect 862 651 868 652
rect 902 656 908 657
rect 902 652 903 656
rect 907 652 908 656
rect 902 651 908 652
rect 934 656 940 657
rect 934 652 935 656
rect 939 652 940 656
rect 934 651 940 652
rect 966 656 972 657
rect 966 652 967 656
rect 971 652 972 656
rect 966 651 972 652
rect 1006 656 1012 657
rect 1006 652 1007 656
rect 1011 652 1012 656
rect 1006 651 1012 652
rect 1046 656 1052 657
rect 1046 652 1047 656
rect 1051 652 1052 656
rect 1046 651 1052 652
rect 1086 656 1092 657
rect 1086 652 1087 656
rect 1091 652 1092 656
rect 1086 651 1092 652
rect 1126 656 1132 657
rect 1126 652 1127 656
rect 1131 652 1132 656
rect 1126 651 1132 652
rect 1158 656 1164 657
rect 1158 652 1159 656
rect 1163 652 1164 656
rect 1158 651 1164 652
rect 1190 656 1196 657
rect 1190 652 1191 656
rect 1195 652 1196 656
rect 1190 651 1196 652
rect 1222 656 1228 657
rect 1222 652 1223 656
rect 1227 652 1228 656
rect 1222 651 1228 652
rect 1262 656 1268 657
rect 1262 652 1263 656
rect 1267 652 1268 656
rect 1262 651 1268 652
rect 1302 656 1308 657
rect 1302 652 1303 656
rect 1307 652 1308 656
rect 1302 651 1308 652
rect 1342 656 1348 657
rect 1342 652 1343 656
rect 1347 652 1348 656
rect 1354 655 1355 659
rect 1359 658 1360 659
rect 1377 658 1379 662
rect 1359 656 1379 658
rect 1359 655 1360 656
rect 1354 654 1360 655
rect 1342 651 1348 652
rect 1446 653 1452 654
rect 846 650 852 651
rect 1446 649 1447 653
rect 1451 649 1452 653
rect 1446 648 1452 649
rect 511 647 517 648
rect 511 643 512 647
rect 516 646 517 647
rect 562 647 568 648
rect 562 646 563 647
rect 516 644 563 646
rect 516 643 517 644
rect 511 642 517 643
rect 562 643 563 644
rect 567 643 568 647
rect 562 642 568 643
rect 615 647 621 648
rect 615 643 616 647
rect 620 646 621 647
rect 674 647 680 648
rect 674 646 675 647
rect 620 644 675 646
rect 620 643 621 644
rect 615 642 621 643
rect 674 643 675 644
rect 679 643 680 647
rect 674 642 680 643
rect 871 647 877 648
rect 871 643 872 647
rect 876 646 877 647
rect 986 647 992 648
rect 986 646 987 647
rect 876 644 987 646
rect 876 643 877 644
rect 871 642 877 643
rect 986 643 987 644
rect 991 643 992 647
rect 986 642 992 643
rect 1078 647 1084 648
rect 1078 643 1079 647
rect 1083 646 1084 647
rect 1170 647 1176 648
rect 1170 646 1171 647
rect 1083 644 1171 646
rect 1083 643 1084 644
rect 1078 642 1084 643
rect 1170 643 1171 644
rect 1175 643 1176 647
rect 1170 642 1176 643
rect 1199 647 1205 648
rect 1199 643 1200 647
rect 1204 646 1205 647
rect 1234 647 1240 648
rect 1234 646 1235 647
rect 1204 644 1235 646
rect 1204 643 1205 644
rect 1199 642 1205 643
rect 1234 643 1235 644
rect 1239 643 1240 647
rect 1234 642 1240 643
rect 1271 647 1277 648
rect 1271 643 1272 647
rect 1276 646 1277 647
rect 1314 647 1320 648
rect 1314 646 1315 647
rect 1276 644 1315 646
rect 1276 643 1277 644
rect 1271 642 1277 643
rect 1314 643 1315 644
rect 1319 643 1320 647
rect 1314 642 1320 643
rect 1322 647 1328 648
rect 1322 643 1323 647
rect 1327 646 1328 647
rect 1351 647 1357 648
rect 1351 646 1352 647
rect 1327 644 1352 646
rect 1327 643 1328 644
rect 1322 642 1328 643
rect 1351 643 1352 644
rect 1356 643 1357 647
rect 1351 642 1357 643
rect 480 640 506 642
rect 223 639 229 640
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 223 635 224 639
rect 228 638 229 639
rect 231 639 237 640
rect 231 638 232 639
rect 228 636 232 638
rect 228 635 229 636
rect 223 634 229 635
rect 231 635 232 636
rect 236 635 237 639
rect 231 634 237 635
rect 271 639 277 640
rect 271 635 272 639
rect 276 638 277 639
rect 335 639 341 640
rect 276 636 307 638
rect 276 635 277 636
rect 271 634 277 635
rect 305 632 307 636
rect 335 635 336 639
rect 340 638 341 639
rect 463 639 469 640
rect 340 636 358 638
rect 340 635 341 636
rect 335 634 341 635
rect 199 631 208 632
rect 223 631 232 632
rect 271 631 280 632
rect 303 631 309 632
rect 335 631 344 632
rect 110 630 116 631
rect 190 630 196 631
rect 190 626 191 630
rect 195 626 196 630
rect 199 627 200 631
rect 207 627 208 631
rect 199 626 208 627
rect 214 630 220 631
rect 214 626 215 630
rect 219 626 220 630
rect 223 627 224 631
rect 231 627 232 631
rect 223 626 232 627
rect 238 630 244 631
rect 238 626 239 630
rect 243 626 244 630
rect 262 630 268 631
rect 190 625 196 626
rect 214 625 220 626
rect 238 625 244 626
rect 247 627 253 628
rect 247 623 248 627
rect 252 623 253 627
rect 262 626 263 630
rect 267 626 268 630
rect 271 627 272 631
rect 279 627 280 631
rect 271 626 280 627
rect 294 630 300 631
rect 294 626 295 630
rect 299 626 300 630
rect 303 627 304 631
rect 308 627 309 631
rect 303 626 309 627
rect 326 630 332 631
rect 326 626 327 630
rect 331 626 332 630
rect 335 627 336 631
rect 343 627 344 631
rect 335 626 344 627
rect 262 625 268 626
rect 294 625 300 626
rect 326 625 332 626
rect 247 622 253 623
rect 343 623 349 624
rect 343 622 344 623
rect 233 620 250 622
rect 281 620 344 622
rect 231 619 237 620
rect 231 615 232 619
rect 236 615 237 619
rect 281 616 283 620
rect 343 619 344 620
rect 348 619 349 623
rect 356 622 358 636
rect 463 635 464 639
rect 468 638 469 639
rect 504 638 506 640
rect 559 639 565 640
rect 559 638 560 639
rect 468 636 499 638
rect 504 636 560 638
rect 468 635 469 636
rect 463 634 469 635
rect 415 631 421 632
rect 366 630 372 631
rect 366 626 367 630
rect 371 626 372 630
rect 406 630 412 631
rect 366 625 372 626
rect 375 627 381 628
rect 375 623 376 627
rect 380 623 381 627
rect 406 626 407 630
rect 411 626 412 630
rect 415 627 416 631
rect 420 630 421 631
rect 446 631 452 632
rect 463 631 472 632
rect 446 630 447 631
rect 420 628 447 630
rect 420 627 421 628
rect 415 626 421 627
rect 446 627 447 628
rect 451 627 452 631
rect 446 626 452 627
rect 454 630 460 631
rect 454 626 455 630
rect 459 626 460 630
rect 463 627 464 631
rect 471 627 472 631
rect 463 626 472 627
rect 406 625 412 626
rect 454 625 460 626
rect 375 622 381 623
rect 497 622 499 636
rect 559 635 560 636
rect 564 635 565 639
rect 559 634 565 635
rect 671 639 677 640
rect 671 635 672 639
rect 676 638 677 639
rect 710 639 716 640
rect 676 636 706 638
rect 676 635 677 636
rect 671 634 677 635
rect 559 631 568 632
rect 615 631 621 632
rect 502 630 508 631
rect 502 626 503 630
rect 507 626 508 630
rect 550 630 556 631
rect 502 625 508 626
rect 511 627 517 628
rect 511 623 512 627
rect 516 623 517 627
rect 550 626 551 630
rect 555 626 556 630
rect 559 627 560 631
rect 567 627 568 631
rect 559 626 568 627
rect 606 630 612 631
rect 606 626 607 630
rect 611 626 612 630
rect 615 627 616 631
rect 620 630 621 631
rect 650 631 656 632
rect 671 631 680 632
rect 650 630 651 631
rect 620 628 651 630
rect 620 627 621 628
rect 615 626 621 627
rect 650 627 651 628
rect 655 627 656 631
rect 650 626 656 627
rect 662 630 668 631
rect 662 626 663 630
rect 667 626 668 630
rect 671 627 672 631
rect 679 627 680 631
rect 671 626 680 627
rect 550 625 556 626
rect 606 625 612 626
rect 662 625 668 626
rect 511 622 517 623
rect 704 622 706 636
rect 710 635 711 639
rect 715 638 716 639
rect 727 639 733 640
rect 727 638 728 639
rect 715 636 728 638
rect 715 635 716 636
rect 710 634 716 635
rect 727 635 728 636
rect 732 635 733 639
rect 727 634 733 635
rect 775 639 781 640
rect 775 635 776 639
rect 780 638 781 639
rect 911 639 917 640
rect 911 638 912 639
rect 780 636 826 638
rect 780 635 781 636
rect 775 634 781 635
rect 824 632 826 636
rect 892 636 912 638
rect 823 631 829 632
rect 871 631 877 632
rect 718 630 724 631
rect 718 626 719 630
rect 723 626 724 630
rect 766 630 772 631
rect 718 625 724 626
rect 727 627 733 628
rect 727 623 728 627
rect 732 623 733 627
rect 766 626 767 630
rect 771 626 772 630
rect 814 630 820 631
rect 766 625 772 626
rect 775 627 781 628
rect 775 624 776 627
rect 727 622 733 623
rect 774 623 776 624
rect 780 623 781 627
rect 814 626 815 630
rect 819 626 820 630
rect 823 627 824 631
rect 828 627 829 631
rect 823 626 829 627
rect 862 630 868 631
rect 862 626 863 630
rect 867 626 868 630
rect 871 627 872 631
rect 876 630 877 631
rect 892 630 894 636
rect 911 635 912 636
rect 916 635 917 639
rect 943 639 949 640
rect 943 638 944 639
rect 911 634 917 635
rect 928 636 944 638
rect 911 631 917 632
rect 876 628 894 630
rect 902 630 908 631
rect 876 627 877 628
rect 871 626 877 627
rect 902 626 903 630
rect 907 626 908 630
rect 911 627 912 631
rect 916 630 917 631
rect 928 630 930 636
rect 943 635 944 636
rect 948 635 949 639
rect 975 639 981 640
rect 975 638 976 639
rect 943 634 949 635
rect 960 636 976 638
rect 943 631 949 632
rect 916 628 930 630
rect 934 630 940 631
rect 916 627 917 628
rect 911 626 917 627
rect 934 626 935 630
rect 939 626 940 630
rect 943 627 944 631
rect 948 630 949 631
rect 960 630 962 636
rect 975 635 976 636
rect 980 635 981 639
rect 1015 639 1021 640
rect 1015 638 1016 639
rect 975 634 981 635
rect 996 636 1016 638
rect 975 631 981 632
rect 948 628 962 630
rect 966 630 972 631
rect 948 627 949 628
rect 943 626 949 627
rect 966 626 967 630
rect 971 626 972 630
rect 975 627 976 631
rect 980 630 981 631
rect 996 630 998 636
rect 1015 635 1016 636
rect 1020 635 1021 639
rect 1055 639 1061 640
rect 1055 638 1056 639
rect 1015 634 1021 635
rect 1040 636 1056 638
rect 1015 631 1021 632
rect 980 628 998 630
rect 1006 630 1012 631
rect 980 627 981 628
rect 975 626 981 627
rect 1006 626 1007 630
rect 1011 626 1012 630
rect 1015 627 1016 631
rect 1020 630 1021 631
rect 1040 630 1042 636
rect 1055 635 1056 636
rect 1060 635 1061 639
rect 1095 639 1101 640
rect 1095 638 1096 639
rect 1055 634 1061 635
rect 1076 636 1096 638
rect 1055 631 1061 632
rect 1020 628 1042 630
rect 1046 630 1052 631
rect 1020 627 1021 628
rect 1015 626 1021 627
rect 1046 626 1047 630
rect 1051 626 1052 630
rect 1055 627 1056 631
rect 1060 630 1061 631
rect 1076 630 1078 636
rect 1095 635 1096 636
rect 1100 635 1101 639
rect 1135 639 1141 640
rect 1135 638 1136 639
rect 1095 634 1101 635
rect 1116 636 1136 638
rect 1095 631 1101 632
rect 1060 628 1078 630
rect 1086 630 1092 631
rect 1060 627 1061 628
rect 1055 626 1061 627
rect 1086 626 1087 630
rect 1091 626 1092 630
rect 1095 627 1096 631
rect 1100 630 1101 631
rect 1116 630 1118 636
rect 1135 635 1136 636
rect 1140 635 1141 639
rect 1135 634 1141 635
rect 1167 639 1173 640
rect 1167 635 1168 639
rect 1172 638 1173 639
rect 1231 639 1237 640
rect 1172 636 1186 638
rect 1172 635 1173 636
rect 1167 634 1173 635
rect 1167 631 1176 632
rect 1100 628 1118 630
rect 1126 630 1132 631
rect 1100 627 1101 628
rect 1095 626 1101 627
rect 1126 626 1127 630
rect 1131 626 1132 630
rect 1158 630 1164 631
rect 814 625 820 626
rect 862 625 868 626
rect 902 625 908 626
rect 934 625 940 626
rect 966 625 972 626
rect 1006 625 1012 626
rect 1046 625 1052 626
rect 1086 625 1092 626
rect 1126 625 1132 626
rect 1135 627 1141 628
rect 356 620 378 622
rect 433 620 451 622
rect 497 620 514 622
rect 704 620 730 622
rect 343 618 349 619
rect 422 619 428 620
rect 279 615 285 616
rect 422 615 423 619
rect 427 616 428 619
rect 427 615 429 616
rect 231 614 237 615
rect 270 614 276 615
rect 270 610 271 614
rect 275 610 276 614
rect 279 611 280 615
rect 284 611 285 615
rect 279 610 285 611
rect 294 614 300 615
rect 294 610 295 614
rect 299 610 300 614
rect 318 614 324 615
rect 110 609 116 610
rect 270 609 276 610
rect 294 609 300 610
rect 303 611 312 612
rect 110 605 111 609
rect 115 605 116 609
rect 303 607 304 611
rect 311 607 312 611
rect 318 610 319 614
rect 323 610 324 614
rect 342 614 348 615
rect 318 609 324 610
rect 327 611 333 612
rect 303 606 312 607
rect 327 607 328 611
rect 332 607 333 611
rect 342 610 343 614
rect 347 610 348 614
rect 366 614 372 615
rect 342 609 348 610
rect 351 611 357 612
rect 327 606 333 607
rect 351 607 352 611
rect 356 607 357 611
rect 366 610 367 614
rect 371 610 372 614
rect 390 614 396 615
rect 366 609 372 610
rect 375 611 381 612
rect 351 606 357 607
rect 375 607 376 611
rect 380 607 381 611
rect 390 610 391 614
rect 395 610 396 614
rect 414 614 420 615
rect 422 614 424 615
rect 390 609 396 610
rect 399 611 408 612
rect 375 606 381 607
rect 399 607 400 611
rect 407 607 408 611
rect 414 610 415 614
rect 419 610 420 614
rect 423 611 424 614
rect 428 611 429 615
rect 423 610 429 611
rect 414 609 420 610
rect 399 606 408 607
rect 110 604 116 605
rect 279 603 285 604
rect 279 599 280 603
rect 284 602 285 603
rect 294 603 300 604
rect 294 602 295 603
rect 284 600 295 602
rect 284 599 285 600
rect 279 598 285 599
rect 294 599 295 600
rect 299 599 300 603
rect 294 598 300 599
rect 303 599 309 600
rect 303 595 304 599
rect 308 598 309 599
rect 328 598 330 606
rect 352 598 354 606
rect 376 598 378 606
rect 390 599 396 600
rect 390 598 391 599
rect 308 596 330 598
rect 340 596 354 598
rect 364 596 378 598
rect 308 595 309 596
rect 303 594 309 595
rect 340 594 342 596
rect 364 594 366 596
rect 388 595 391 598
rect 395 595 396 599
rect 388 594 396 595
rect 399 599 405 600
rect 399 595 400 599
rect 404 598 405 599
rect 414 599 420 600
rect 414 598 415 599
rect 404 596 415 598
rect 404 595 405 596
rect 399 594 405 595
rect 414 595 415 596
rect 419 595 420 599
rect 414 594 420 595
rect 336 592 342 594
rect 360 592 366 594
rect 376 592 390 594
rect 110 591 116 592
rect 110 587 111 591
rect 115 587 116 591
rect 327 591 333 592
rect 110 586 116 587
rect 270 588 276 589
rect 270 584 271 588
rect 275 584 276 588
rect 270 583 276 584
rect 294 588 300 589
rect 294 584 295 588
rect 299 584 300 588
rect 294 583 300 584
rect 318 588 324 589
rect 318 584 319 588
rect 323 584 324 588
rect 327 587 328 591
rect 332 590 333 591
rect 336 590 338 592
rect 332 588 338 590
rect 351 591 357 592
rect 342 588 348 589
rect 332 587 333 588
rect 327 586 333 587
rect 318 583 324 584
rect 342 584 343 588
rect 347 584 348 588
rect 351 587 352 591
rect 356 590 357 591
rect 360 590 362 592
rect 356 588 362 590
rect 375 591 381 592
rect 366 588 372 589
rect 356 587 357 588
rect 351 586 357 587
rect 342 583 348 584
rect 366 584 367 588
rect 371 584 372 588
rect 375 587 376 591
rect 380 587 381 591
rect 375 586 381 587
rect 390 588 396 589
rect 366 583 372 584
rect 390 584 391 588
rect 395 584 396 588
rect 390 583 396 584
rect 414 588 420 589
rect 414 584 415 588
rect 419 584 420 588
rect 414 583 420 584
rect 423 587 429 588
rect 423 583 424 587
rect 428 586 429 587
rect 433 586 435 620
rect 449 616 451 620
rect 774 619 775 623
rect 779 622 781 623
rect 1034 623 1040 624
rect 779 619 780 622
rect 774 618 780 619
rect 1034 619 1035 623
rect 1039 622 1040 623
rect 1135 623 1136 627
rect 1140 623 1141 627
rect 1158 626 1159 630
rect 1163 626 1164 630
rect 1167 627 1168 631
rect 1175 627 1176 631
rect 1167 626 1176 627
rect 1158 625 1164 626
rect 1135 622 1141 623
rect 1184 622 1186 636
rect 1231 635 1232 639
rect 1236 638 1237 639
rect 1311 639 1317 640
rect 1236 636 1254 638
rect 1236 635 1237 636
rect 1231 634 1237 635
rect 1231 631 1240 632
rect 1190 630 1196 631
rect 1190 626 1191 630
rect 1195 626 1196 630
rect 1222 630 1228 631
rect 1190 625 1196 626
rect 1199 627 1205 628
rect 1199 623 1200 627
rect 1204 623 1205 627
rect 1222 626 1223 630
rect 1227 626 1228 630
rect 1231 627 1232 631
rect 1239 627 1240 631
rect 1231 626 1240 627
rect 1222 625 1228 626
rect 1199 622 1205 623
rect 1252 622 1254 636
rect 1311 635 1312 639
rect 1316 638 1317 639
rect 1316 636 1339 638
rect 1316 635 1317 636
rect 1311 634 1317 635
rect 1311 631 1320 632
rect 1262 630 1268 631
rect 1262 626 1263 630
rect 1267 626 1268 630
rect 1302 630 1308 631
rect 1262 625 1268 626
rect 1271 627 1277 628
rect 1271 623 1272 627
rect 1276 623 1277 627
rect 1302 626 1303 630
rect 1307 626 1308 630
rect 1311 627 1312 631
rect 1319 627 1320 631
rect 1311 626 1320 627
rect 1302 625 1308 626
rect 1271 622 1277 623
rect 1322 623 1328 624
rect 1322 622 1323 623
rect 1039 620 1138 622
rect 1184 620 1203 622
rect 1232 620 1250 622
rect 1252 620 1274 622
rect 1280 620 1323 622
rect 1039 619 1040 620
rect 1034 618 1040 619
rect 447 615 453 616
rect 687 615 693 616
rect 438 614 444 615
rect 438 610 439 614
rect 443 610 444 614
rect 447 611 448 615
rect 452 611 453 615
rect 447 610 453 611
rect 478 614 484 615
rect 478 610 479 614
rect 483 610 484 614
rect 518 614 524 615
rect 438 609 444 610
rect 478 609 484 610
rect 487 611 493 612
rect 487 607 488 611
rect 492 607 493 611
rect 518 610 519 614
rect 523 610 524 614
rect 566 614 572 615
rect 518 609 524 610
rect 527 611 533 612
rect 487 606 493 607
rect 527 607 528 611
rect 532 607 533 611
rect 566 610 567 614
rect 571 610 572 614
rect 622 614 628 615
rect 566 609 572 610
rect 575 611 581 612
rect 527 606 533 607
rect 575 607 576 611
rect 580 610 581 611
rect 622 610 623 614
rect 627 610 628 614
rect 678 614 684 615
rect 580 608 606 610
rect 622 609 628 610
rect 631 611 637 612
rect 580 607 581 608
rect 575 606 581 607
rect 488 598 490 606
rect 528 598 530 606
rect 604 602 606 608
rect 631 607 632 611
rect 636 610 637 611
rect 678 610 679 614
rect 683 610 684 614
rect 687 611 688 615
rect 692 614 693 615
rect 710 615 716 616
rect 983 615 992 616
rect 1199 615 1205 616
rect 710 614 711 615
rect 692 612 711 614
rect 692 611 693 612
rect 687 610 693 611
rect 710 611 711 612
rect 715 611 716 615
rect 710 610 716 611
rect 734 614 740 615
rect 734 610 735 614
rect 739 610 740 614
rect 782 614 788 615
rect 636 608 670 610
rect 678 609 684 610
rect 734 609 740 610
rect 743 611 749 612
rect 636 607 637 608
rect 631 606 637 607
rect 631 603 637 604
rect 631 602 632 603
rect 604 600 632 602
rect 631 599 632 600
rect 636 599 637 603
rect 668 602 670 608
rect 743 607 744 611
rect 748 610 749 611
rect 767 611 773 612
rect 767 610 768 611
rect 748 608 768 610
rect 748 607 749 608
rect 743 606 749 607
rect 767 607 768 608
rect 772 607 773 611
rect 782 610 783 614
rect 787 610 788 614
rect 830 614 836 615
rect 782 609 788 610
rect 791 611 800 612
rect 767 606 773 607
rect 791 607 792 611
rect 799 607 800 611
rect 830 610 831 614
rect 835 610 836 614
rect 878 614 884 615
rect 830 609 836 610
rect 839 611 845 612
rect 791 606 800 607
rect 839 607 840 611
rect 844 607 845 611
rect 878 610 879 614
rect 883 610 884 614
rect 926 614 932 615
rect 878 609 884 610
rect 887 611 893 612
rect 839 606 845 607
rect 887 607 888 611
rect 892 610 893 611
rect 926 610 927 614
rect 931 610 932 614
rect 974 614 980 615
rect 892 608 914 610
rect 926 609 932 610
rect 935 611 941 612
rect 892 607 893 608
rect 887 606 893 607
rect 687 603 693 604
rect 687 602 688 603
rect 668 600 688 602
rect 631 598 637 599
rect 687 599 688 600
rect 692 599 693 603
rect 687 598 693 599
rect 743 603 749 604
rect 743 599 744 603
rect 748 602 749 603
rect 774 603 780 604
rect 774 602 775 603
rect 748 600 775 602
rect 748 599 749 600
rect 743 598 749 599
rect 774 599 775 600
rect 779 599 780 603
rect 841 602 843 606
rect 887 603 893 604
rect 887 602 888 603
rect 841 600 888 602
rect 774 598 780 599
rect 783 599 789 600
rect 468 596 490 598
rect 508 596 530 598
rect 447 595 453 596
rect 447 591 448 595
rect 452 594 453 595
rect 468 594 470 596
rect 452 592 470 594
rect 452 591 453 592
rect 447 590 453 591
rect 487 591 493 592
rect 428 584 435 586
rect 438 588 444 589
rect 438 584 439 588
rect 443 584 444 588
rect 428 583 429 584
rect 438 583 444 584
rect 478 588 484 589
rect 478 584 479 588
rect 483 584 484 588
rect 487 587 488 591
rect 492 590 493 591
rect 508 590 510 596
rect 783 595 784 599
rect 788 598 789 599
rect 791 599 797 600
rect 791 598 792 599
rect 788 596 792 598
rect 788 595 789 596
rect 783 594 789 595
rect 791 595 792 596
rect 796 595 797 599
rect 887 599 888 600
rect 892 599 893 603
rect 912 602 914 608
rect 935 607 936 611
rect 940 610 941 611
rect 974 610 975 614
rect 979 610 980 614
rect 983 611 984 615
rect 991 611 992 615
rect 983 610 992 611
rect 1022 614 1028 615
rect 1022 610 1023 614
rect 1027 610 1028 614
rect 1070 614 1076 615
rect 940 608 962 610
rect 974 609 980 610
rect 1022 609 1028 610
rect 1031 611 1037 612
rect 940 607 941 608
rect 935 606 941 607
rect 935 603 941 604
rect 935 602 936 603
rect 912 600 936 602
rect 887 598 893 599
rect 935 599 936 600
rect 940 599 941 603
rect 960 602 962 608
rect 1031 607 1032 611
rect 1036 610 1037 611
rect 1070 610 1071 614
rect 1075 610 1076 614
rect 1110 614 1116 615
rect 1036 608 1058 610
rect 1070 609 1076 610
rect 1079 611 1085 612
rect 1036 607 1037 608
rect 1031 606 1037 607
rect 983 603 989 604
rect 983 602 984 603
rect 960 600 984 602
rect 935 598 941 599
rect 983 599 984 600
rect 988 599 989 603
rect 983 598 989 599
rect 1031 603 1040 604
rect 1031 599 1032 603
rect 1039 599 1040 603
rect 1056 602 1058 608
rect 1079 607 1080 611
rect 1084 610 1085 611
rect 1110 610 1111 614
rect 1115 610 1116 614
rect 1150 614 1156 615
rect 1084 608 1102 610
rect 1110 609 1116 610
rect 1119 611 1125 612
rect 1084 607 1085 608
rect 1079 606 1085 607
rect 1079 603 1085 604
rect 1079 602 1080 603
rect 1056 600 1080 602
rect 1031 598 1040 599
rect 1079 599 1080 600
rect 1084 599 1085 603
rect 1100 602 1102 608
rect 1119 607 1120 611
rect 1124 610 1125 611
rect 1150 610 1151 614
rect 1155 610 1156 614
rect 1190 614 1196 615
rect 1124 608 1147 610
rect 1150 609 1156 610
rect 1159 611 1165 612
rect 1124 607 1125 608
rect 1119 606 1125 607
rect 1119 603 1125 604
rect 1119 602 1120 603
rect 1100 600 1120 602
rect 1079 598 1085 599
rect 1119 599 1120 600
rect 1124 599 1125 603
rect 1145 602 1147 608
rect 1159 607 1160 611
rect 1164 610 1165 611
rect 1175 611 1181 612
rect 1175 610 1176 611
rect 1164 608 1176 610
rect 1164 607 1165 608
rect 1159 606 1165 607
rect 1175 607 1176 608
rect 1180 607 1181 611
rect 1190 610 1191 614
rect 1195 610 1196 614
rect 1199 611 1200 615
rect 1204 614 1205 615
rect 1232 614 1234 620
rect 1248 618 1250 620
rect 1280 618 1282 620
rect 1322 619 1323 620
rect 1327 619 1328 623
rect 1337 622 1339 636
rect 1446 635 1452 636
rect 1446 631 1447 635
rect 1451 631 1452 635
rect 1342 630 1348 631
rect 1446 630 1452 631
rect 1342 626 1343 630
rect 1347 626 1348 630
rect 1342 625 1348 626
rect 1351 627 1357 628
rect 1351 623 1352 627
rect 1356 623 1357 627
rect 1351 622 1357 623
rect 1337 620 1354 622
rect 1322 618 1328 619
rect 1248 616 1282 618
rect 1204 612 1234 614
rect 1238 614 1244 615
rect 1204 611 1205 612
rect 1199 610 1205 611
rect 1238 610 1239 614
rect 1243 610 1244 614
rect 1286 614 1292 615
rect 1190 609 1196 610
rect 1238 609 1244 610
rect 1247 611 1253 612
rect 1175 606 1181 607
rect 1247 607 1248 611
rect 1252 607 1253 611
rect 1286 610 1287 614
rect 1291 610 1292 614
rect 1334 614 1340 615
rect 1286 609 1292 610
rect 1295 611 1301 612
rect 1247 606 1253 607
rect 1295 607 1296 611
rect 1300 607 1301 611
rect 1334 610 1335 614
rect 1339 610 1340 614
rect 1334 609 1340 610
rect 1343 611 1349 612
rect 1295 606 1301 607
rect 1343 607 1344 611
rect 1348 607 1349 611
rect 1343 606 1349 607
rect 1446 609 1452 610
rect 1159 603 1165 604
rect 1159 602 1160 603
rect 1145 600 1160 602
rect 1119 598 1125 599
rect 1159 599 1160 600
rect 1164 599 1165 603
rect 1159 598 1165 599
rect 1199 603 1205 604
rect 1199 599 1200 603
rect 1204 602 1205 603
rect 1248 602 1250 606
rect 1204 600 1250 602
rect 1204 599 1205 600
rect 1199 598 1205 599
rect 1296 598 1298 606
rect 1344 598 1346 606
rect 1446 605 1447 609
rect 1451 605 1452 609
rect 1446 604 1452 605
rect 1272 596 1298 598
rect 1321 596 1346 598
rect 791 594 797 595
rect 1247 595 1253 596
rect 492 588 510 590
rect 527 591 536 592
rect 518 588 524 589
rect 492 587 493 588
rect 487 586 493 587
rect 478 583 484 584
rect 518 584 519 588
rect 523 584 524 588
rect 527 587 528 591
rect 535 587 536 591
rect 1247 591 1248 595
rect 1252 594 1253 595
rect 1272 594 1274 596
rect 1252 592 1274 594
rect 1252 591 1253 592
rect 1247 590 1253 591
rect 1295 591 1301 592
rect 527 586 536 587
rect 566 588 572 589
rect 622 588 628 589
rect 518 583 524 584
rect 566 584 567 588
rect 571 584 572 588
rect 566 583 572 584
rect 575 587 581 588
rect 575 583 576 587
rect 580 586 581 587
rect 614 587 620 588
rect 614 586 615 587
rect 580 584 615 586
rect 580 583 581 584
rect 423 582 429 583
rect 575 582 581 583
rect 614 583 615 584
rect 619 583 620 587
rect 622 584 623 588
rect 627 584 628 588
rect 622 583 628 584
rect 678 588 684 589
rect 678 584 679 588
rect 683 584 684 588
rect 678 583 684 584
rect 734 588 740 589
rect 734 584 735 588
rect 739 584 740 588
rect 734 583 740 584
rect 782 588 788 589
rect 782 584 783 588
rect 787 584 788 588
rect 782 583 788 584
rect 830 588 836 589
rect 878 588 884 589
rect 830 584 831 588
rect 835 584 836 588
rect 830 583 836 584
rect 839 587 845 588
rect 839 583 840 587
rect 844 586 845 587
rect 870 587 876 588
rect 870 586 871 587
rect 844 584 871 586
rect 844 583 845 584
rect 614 582 620 583
rect 839 582 845 583
rect 870 583 871 584
rect 875 583 876 587
rect 878 584 879 588
rect 883 584 884 588
rect 878 583 884 584
rect 926 588 932 589
rect 926 584 927 588
rect 931 584 932 588
rect 926 583 932 584
rect 974 588 980 589
rect 974 584 975 588
rect 979 584 980 588
rect 974 583 980 584
rect 1022 588 1028 589
rect 1022 584 1023 588
rect 1027 584 1028 588
rect 1022 583 1028 584
rect 1070 588 1076 589
rect 1070 584 1071 588
rect 1075 584 1076 588
rect 1070 583 1076 584
rect 1110 588 1116 589
rect 1110 584 1111 588
rect 1115 584 1116 588
rect 1110 583 1116 584
rect 1150 588 1156 589
rect 1150 584 1151 588
rect 1155 584 1156 588
rect 1150 583 1156 584
rect 1190 588 1196 589
rect 1190 584 1191 588
rect 1195 584 1196 588
rect 1190 583 1196 584
rect 1238 588 1244 589
rect 1238 584 1239 588
rect 1243 584 1244 588
rect 1238 583 1244 584
rect 1286 588 1292 589
rect 1286 584 1287 588
rect 1291 584 1292 588
rect 1295 587 1296 591
rect 1300 590 1301 591
rect 1321 590 1323 596
rect 1300 588 1323 590
rect 1446 591 1452 592
rect 1334 588 1340 589
rect 1300 587 1301 588
rect 1295 586 1301 587
rect 1286 583 1292 584
rect 1334 584 1335 588
rect 1339 584 1340 588
rect 1334 583 1340 584
rect 1343 587 1349 588
rect 1343 583 1344 587
rect 1348 586 1349 587
rect 1386 587 1392 588
rect 1386 586 1387 587
rect 1348 584 1387 586
rect 1348 583 1349 584
rect 870 582 876 583
rect 1343 582 1349 583
rect 1386 583 1387 584
rect 1391 583 1392 587
rect 1446 587 1447 591
rect 1451 587 1452 591
rect 1446 586 1452 587
rect 1386 582 1392 583
rect 262 576 268 577
rect 110 573 116 574
rect 110 569 111 573
rect 115 569 116 573
rect 262 572 263 576
rect 267 572 268 576
rect 262 571 268 572
rect 286 576 292 577
rect 286 572 287 576
rect 291 572 292 576
rect 286 571 292 572
rect 310 576 316 577
rect 310 572 311 576
rect 315 572 316 576
rect 310 571 316 572
rect 334 576 340 577
rect 334 572 335 576
rect 339 572 340 576
rect 334 571 340 572
rect 358 576 364 577
rect 358 572 359 576
rect 363 572 364 576
rect 358 571 364 572
rect 382 576 388 577
rect 382 572 383 576
rect 387 572 388 576
rect 382 571 388 572
rect 406 576 412 577
rect 406 572 407 576
rect 411 572 412 576
rect 406 571 412 572
rect 430 576 436 577
rect 430 572 431 576
rect 435 572 436 576
rect 462 576 468 577
rect 462 572 463 576
rect 467 572 468 576
rect 430 571 436 572
rect 439 571 445 572
rect 462 571 468 572
rect 502 576 508 577
rect 502 572 503 576
rect 507 572 508 576
rect 502 571 508 572
rect 550 576 556 577
rect 550 572 551 576
rect 555 572 556 576
rect 550 571 556 572
rect 606 576 612 577
rect 606 572 607 576
rect 611 572 612 576
rect 606 571 612 572
rect 662 576 668 577
rect 662 572 663 576
rect 667 572 668 576
rect 662 571 668 572
rect 718 576 724 577
rect 718 572 719 576
rect 723 572 724 576
rect 718 571 724 572
rect 774 576 780 577
rect 830 576 836 577
rect 774 572 775 576
rect 779 572 780 576
rect 774 571 780 572
rect 783 575 789 576
rect 783 571 784 575
rect 788 574 789 575
rect 794 575 800 576
rect 794 574 795 575
rect 788 572 795 574
rect 788 571 789 572
rect 110 568 116 569
rect 271 567 277 568
rect 271 563 272 567
rect 276 566 277 567
rect 398 567 404 568
rect 398 566 399 567
rect 276 564 399 566
rect 276 563 277 564
rect 271 562 277 563
rect 398 563 399 564
rect 403 563 404 567
rect 439 567 440 571
rect 444 567 445 571
rect 783 570 789 571
rect 794 571 795 572
rect 799 571 800 575
rect 830 572 831 576
rect 835 572 836 576
rect 830 571 836 572
rect 886 576 892 577
rect 886 572 887 576
rect 891 572 892 576
rect 886 571 892 572
rect 942 576 948 577
rect 942 572 943 576
rect 947 572 948 576
rect 942 571 948 572
rect 1006 576 1012 577
rect 1006 572 1007 576
rect 1011 572 1012 576
rect 1006 571 1012 572
rect 1070 576 1076 577
rect 1070 572 1071 576
rect 1075 572 1076 576
rect 1070 571 1076 572
rect 1126 576 1132 577
rect 1126 572 1127 576
rect 1131 572 1132 576
rect 1126 571 1132 572
rect 1182 576 1188 577
rect 1182 572 1183 576
rect 1187 572 1188 576
rect 1182 571 1188 572
rect 1246 576 1252 577
rect 1246 572 1247 576
rect 1251 572 1252 576
rect 1246 571 1252 572
rect 1310 576 1316 577
rect 1310 572 1311 576
rect 1315 572 1316 576
rect 1310 571 1316 572
rect 1374 576 1380 577
rect 1374 572 1375 576
rect 1379 572 1380 576
rect 1374 571 1380 572
rect 1446 573 1452 574
rect 794 570 800 571
rect 1446 569 1447 573
rect 1451 569 1452 573
rect 1446 568 1452 569
rect 439 566 445 567
rect 559 567 565 568
rect 559 566 560 567
rect 398 562 404 563
rect 480 564 560 566
rect 295 559 301 560
rect 295 558 296 559
rect 281 556 296 558
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 271 551 277 552
rect 110 550 116 551
rect 262 550 268 551
rect 262 546 263 550
rect 267 546 268 550
rect 271 547 272 551
rect 276 550 277 551
rect 281 550 283 556
rect 295 555 296 556
rect 300 555 301 559
rect 319 559 325 560
rect 319 558 320 559
rect 295 554 301 555
rect 305 556 320 558
rect 295 551 301 552
rect 276 548 283 550
rect 286 550 292 551
rect 276 547 277 548
rect 271 546 277 547
rect 286 546 287 550
rect 291 546 292 550
rect 295 547 296 551
rect 300 550 301 551
rect 305 550 307 556
rect 319 555 320 556
rect 324 555 325 559
rect 343 559 349 560
rect 343 558 344 559
rect 319 554 325 555
rect 328 556 344 558
rect 319 551 325 552
rect 300 548 307 550
rect 310 550 316 551
rect 300 547 301 548
rect 295 546 301 547
rect 310 546 311 550
rect 315 546 316 550
rect 319 547 320 551
rect 324 550 325 551
rect 328 550 330 556
rect 343 555 344 556
rect 348 555 349 559
rect 367 559 373 560
rect 367 558 368 559
rect 343 554 349 555
rect 352 556 368 558
rect 343 551 349 552
rect 324 548 330 550
rect 334 550 340 551
rect 324 547 325 548
rect 319 546 325 547
rect 334 546 335 550
rect 339 546 340 550
rect 343 547 344 551
rect 348 550 349 551
rect 352 550 354 556
rect 367 555 368 556
rect 372 555 373 559
rect 391 559 397 560
rect 391 558 392 559
rect 367 554 373 555
rect 376 556 392 558
rect 367 551 373 552
rect 348 548 354 550
rect 358 550 364 551
rect 348 547 349 548
rect 343 546 349 547
rect 358 546 359 550
rect 363 546 364 550
rect 367 547 368 551
rect 372 550 373 551
rect 376 550 378 556
rect 391 555 392 556
rect 396 555 397 559
rect 415 559 421 560
rect 415 558 416 559
rect 391 554 397 555
rect 401 556 416 558
rect 391 551 397 552
rect 372 548 378 550
rect 382 550 388 551
rect 372 547 373 548
rect 367 546 373 547
rect 382 546 383 550
rect 387 546 388 550
rect 391 547 392 551
rect 396 550 397 551
rect 401 550 403 556
rect 415 555 416 556
rect 420 555 421 559
rect 471 559 477 560
rect 471 558 472 559
rect 415 554 421 555
rect 456 556 472 558
rect 415 551 421 552
rect 439 551 445 552
rect 396 548 403 550
rect 406 550 412 551
rect 396 547 397 548
rect 391 546 397 547
rect 406 546 407 550
rect 411 546 412 550
rect 415 547 416 551
rect 420 547 421 551
rect 415 546 421 547
rect 430 550 436 551
rect 430 546 431 550
rect 435 546 436 550
rect 439 547 440 551
rect 444 550 445 551
rect 456 550 458 556
rect 471 555 472 556
rect 476 555 477 559
rect 471 554 477 555
rect 471 551 477 552
rect 444 548 458 550
rect 462 550 468 551
rect 444 547 445 548
rect 439 546 445 547
rect 462 546 463 550
rect 467 546 468 550
rect 471 547 472 551
rect 476 550 477 551
rect 480 550 482 564
rect 559 563 560 564
rect 564 563 565 567
rect 559 562 565 563
rect 615 567 621 568
rect 615 563 616 567
rect 620 566 621 567
rect 674 567 680 568
rect 674 566 675 567
rect 620 564 675 566
rect 620 563 621 564
rect 615 562 621 563
rect 674 563 675 564
rect 679 563 680 567
rect 674 562 680 563
rect 839 567 845 568
rect 839 563 840 567
rect 844 566 845 567
rect 1034 567 1040 568
rect 1034 566 1035 567
rect 844 564 1035 566
rect 844 563 845 564
rect 839 562 845 563
rect 1034 563 1035 564
rect 1039 563 1040 567
rect 1034 562 1040 563
rect 1079 567 1085 568
rect 1079 563 1080 567
rect 1084 566 1085 567
rect 1138 567 1144 568
rect 1138 566 1139 567
rect 1084 564 1139 566
rect 1084 563 1085 564
rect 1079 562 1085 563
rect 1138 563 1139 564
rect 1143 563 1144 567
rect 1138 562 1144 563
rect 1175 567 1181 568
rect 1175 563 1176 567
rect 1180 566 1181 567
rect 1191 567 1197 568
rect 1191 566 1192 567
rect 1180 564 1192 566
rect 1180 563 1181 564
rect 1175 562 1181 563
rect 1191 563 1192 564
rect 1196 563 1197 567
rect 1191 562 1197 563
rect 511 559 517 560
rect 511 555 512 559
rect 516 558 517 559
rect 538 559 544 560
rect 538 558 539 559
rect 516 556 539 558
rect 516 555 517 556
rect 511 554 517 555
rect 538 555 539 556
rect 543 555 544 559
rect 671 559 677 560
rect 671 558 672 559
rect 538 554 544 555
rect 600 556 672 558
rect 559 551 565 552
rect 476 548 482 550
rect 502 550 508 551
rect 476 547 477 548
rect 471 546 477 547
rect 502 546 503 550
rect 507 546 508 550
rect 550 550 556 551
rect 262 545 268 546
rect 286 545 292 546
rect 310 545 316 546
rect 334 545 340 546
rect 358 545 364 546
rect 382 545 388 546
rect 406 545 412 546
rect 430 545 436 546
rect 462 545 468 546
rect 502 545 508 546
rect 511 547 520 548
rect 511 543 512 547
rect 519 543 520 547
rect 550 546 551 550
rect 555 546 556 550
rect 559 547 560 551
rect 564 550 565 551
rect 600 550 602 556
rect 671 555 672 556
rect 676 555 677 559
rect 671 554 677 555
rect 727 559 733 560
rect 727 555 728 559
rect 732 558 733 559
rect 895 559 901 560
rect 895 558 896 559
rect 732 556 786 558
rect 732 555 733 556
rect 727 554 733 555
rect 784 552 786 556
rect 864 556 896 558
rect 615 551 624 552
rect 671 551 680 552
rect 783 551 789 552
rect 839 551 845 552
rect 564 548 602 550
rect 606 550 612 551
rect 564 547 565 548
rect 559 546 565 547
rect 606 546 607 550
rect 611 546 612 550
rect 615 547 616 551
rect 623 547 624 551
rect 615 546 624 547
rect 662 550 668 551
rect 662 546 663 550
rect 667 546 668 550
rect 671 547 672 551
rect 679 547 680 551
rect 671 546 680 547
rect 718 550 724 551
rect 718 546 719 550
rect 723 546 724 550
rect 774 550 780 551
rect 550 545 556 546
rect 606 545 612 546
rect 662 545 668 546
rect 718 545 724 546
rect 727 547 736 548
rect 511 542 520 543
rect 586 543 592 544
rect 398 539 404 540
rect 398 535 399 539
rect 403 536 404 539
rect 586 539 587 543
rect 591 542 592 543
rect 727 543 728 547
rect 735 543 736 547
rect 774 546 775 550
rect 779 546 780 550
rect 783 547 784 551
rect 788 547 789 551
rect 783 546 789 547
rect 830 550 836 551
rect 830 546 831 550
rect 835 546 836 550
rect 839 547 840 551
rect 844 550 845 551
rect 864 550 866 556
rect 895 555 896 556
rect 900 555 901 559
rect 951 559 957 560
rect 951 558 952 559
rect 895 554 901 555
rect 924 556 952 558
rect 895 551 901 552
rect 844 548 866 550
rect 886 550 892 551
rect 844 547 845 548
rect 839 546 845 547
rect 886 546 887 550
rect 891 546 892 550
rect 895 547 896 551
rect 900 550 901 551
rect 924 550 926 556
rect 951 555 952 556
rect 956 555 957 559
rect 1015 559 1021 560
rect 1015 558 1016 559
rect 951 554 957 555
rect 984 556 1016 558
rect 951 551 957 552
rect 900 548 926 550
rect 942 550 948 551
rect 900 547 901 548
rect 895 546 901 547
rect 942 546 943 550
rect 947 546 948 550
rect 951 547 952 551
rect 956 550 957 551
rect 984 550 986 556
rect 1015 555 1016 556
rect 1020 555 1021 559
rect 1015 554 1021 555
rect 1135 559 1141 560
rect 1135 555 1136 559
rect 1140 558 1141 559
rect 1255 559 1261 560
rect 1140 556 1161 558
rect 1140 555 1141 556
rect 1135 554 1141 555
rect 1135 551 1144 552
rect 956 548 986 550
rect 1006 550 1012 551
rect 956 547 957 548
rect 951 546 957 547
rect 1006 546 1007 550
rect 1011 546 1012 550
rect 1070 550 1076 551
rect 774 545 780 546
rect 830 545 836 546
rect 886 545 892 546
rect 942 545 948 546
rect 1006 545 1012 546
rect 1015 547 1021 548
rect 727 542 736 543
rect 870 543 876 544
rect 591 540 634 542
rect 591 539 592 540
rect 586 538 592 539
rect 632 536 634 540
rect 870 539 871 543
rect 875 542 876 543
rect 1015 543 1016 547
rect 1020 543 1021 547
rect 1070 546 1071 550
rect 1075 546 1076 550
rect 1126 550 1132 551
rect 1070 545 1076 546
rect 1079 547 1085 548
rect 1015 542 1021 543
rect 1079 543 1080 547
rect 1084 546 1085 547
rect 1090 547 1096 548
rect 1090 546 1091 547
rect 1084 544 1091 546
rect 1084 543 1085 544
rect 1079 542 1085 543
rect 1090 543 1091 544
rect 1095 543 1096 547
rect 1126 546 1127 550
rect 1131 546 1132 550
rect 1135 547 1136 551
rect 1143 547 1144 551
rect 1135 546 1144 547
rect 1126 545 1132 546
rect 1090 542 1096 543
rect 1159 542 1161 556
rect 1255 555 1256 559
rect 1260 558 1261 559
rect 1282 559 1288 560
rect 1282 558 1283 559
rect 1260 556 1283 558
rect 1260 555 1261 556
rect 1255 554 1261 555
rect 1282 555 1283 556
rect 1287 555 1288 559
rect 1319 559 1325 560
rect 1319 558 1320 559
rect 1282 554 1288 555
rect 1292 556 1320 558
rect 1255 551 1261 552
rect 1182 550 1188 551
rect 1182 546 1183 550
rect 1187 546 1188 550
rect 1246 550 1252 551
rect 1182 545 1188 546
rect 1191 547 1197 548
rect 1191 543 1192 547
rect 1196 543 1197 547
rect 1246 546 1247 550
rect 1251 546 1252 550
rect 1255 547 1256 551
rect 1260 550 1261 551
rect 1292 550 1294 556
rect 1319 555 1320 556
rect 1324 555 1325 559
rect 1383 559 1389 560
rect 1383 558 1384 559
rect 1319 554 1325 555
rect 1352 556 1384 558
rect 1319 551 1325 552
rect 1260 548 1294 550
rect 1310 550 1316 551
rect 1260 547 1261 548
rect 1255 546 1261 547
rect 1310 546 1311 550
rect 1315 546 1316 550
rect 1319 547 1320 551
rect 1324 550 1325 551
rect 1352 550 1354 556
rect 1383 555 1384 556
rect 1388 555 1389 559
rect 1383 554 1389 555
rect 1446 555 1452 556
rect 1383 551 1392 552
rect 1324 548 1354 550
rect 1374 550 1380 551
rect 1324 547 1325 548
rect 1319 546 1325 547
rect 1374 546 1375 550
rect 1379 546 1380 550
rect 1383 547 1384 551
rect 1391 547 1392 551
rect 1446 551 1447 555
rect 1451 551 1452 555
rect 1446 550 1452 551
rect 1383 546 1392 547
rect 1246 545 1252 546
rect 1310 545 1316 546
rect 1374 545 1380 546
rect 1191 542 1197 543
rect 1362 543 1368 544
rect 875 540 1018 542
rect 1159 540 1195 542
rect 875 539 876 540
rect 870 538 876 539
rect 1362 539 1363 543
rect 1367 542 1368 543
rect 1367 540 1403 542
rect 1367 539 1368 540
rect 1362 538 1368 539
rect 1401 536 1403 540
rect 403 535 405 536
rect 535 535 544 536
rect 631 535 637 536
rect 1031 535 1040 536
rect 1279 535 1288 536
rect 1399 535 1405 536
rect 222 534 228 535
rect 222 530 223 534
rect 227 530 228 534
rect 246 534 252 535
rect 110 529 116 530
rect 222 529 228 530
rect 231 531 240 532
rect 110 525 111 529
rect 115 525 116 529
rect 231 527 232 531
rect 239 527 240 531
rect 246 530 247 534
rect 251 530 252 534
rect 270 534 276 535
rect 246 529 252 530
rect 255 531 261 532
rect 231 526 240 527
rect 255 527 256 531
rect 260 527 261 531
rect 270 530 271 534
rect 275 530 276 534
rect 294 534 300 535
rect 270 529 276 530
rect 279 531 285 532
rect 255 526 261 527
rect 279 527 280 531
rect 284 527 285 531
rect 294 530 295 534
rect 299 530 300 534
rect 326 534 332 535
rect 294 529 300 530
rect 303 531 309 532
rect 279 526 285 527
rect 303 527 304 531
rect 308 530 309 531
rect 326 530 327 534
rect 331 530 332 534
rect 358 534 364 535
rect 308 528 322 530
rect 326 529 332 530
rect 335 531 341 532
rect 308 527 309 528
rect 303 526 309 527
rect 110 524 116 525
rect 257 518 259 526
rect 281 522 283 526
rect 303 523 309 524
rect 303 522 304 523
rect 281 520 304 522
rect 303 519 304 520
rect 308 519 309 523
rect 320 522 322 528
rect 335 527 336 531
rect 340 530 341 531
rect 358 530 359 534
rect 363 530 364 534
rect 390 534 396 535
rect 398 534 400 535
rect 340 528 354 530
rect 358 529 364 530
rect 367 531 373 532
rect 340 527 341 528
rect 335 526 341 527
rect 335 523 341 524
rect 335 522 336 523
rect 320 520 336 522
rect 303 518 309 519
rect 335 519 336 520
rect 340 519 341 523
rect 352 522 354 528
rect 367 527 368 531
rect 372 530 373 531
rect 390 530 391 534
rect 395 530 396 534
rect 399 531 400 534
rect 404 531 405 535
rect 399 530 405 531
rect 422 534 428 535
rect 422 530 423 534
rect 427 530 428 534
rect 454 534 460 535
rect 372 528 386 530
rect 390 529 396 530
rect 422 529 428 530
rect 431 531 437 532
rect 372 527 373 528
rect 367 526 373 527
rect 367 523 373 524
rect 367 522 368 523
rect 352 520 368 522
rect 335 518 341 519
rect 367 519 368 520
rect 372 519 373 523
rect 384 522 386 528
rect 431 527 432 531
rect 436 530 437 531
rect 446 531 452 532
rect 446 530 447 531
rect 436 528 447 530
rect 436 527 437 528
rect 431 526 437 527
rect 446 527 447 528
rect 451 527 452 531
rect 454 530 455 534
rect 459 530 460 534
rect 486 534 492 535
rect 454 529 460 530
rect 463 531 472 532
rect 446 526 452 527
rect 463 527 464 531
rect 471 527 472 531
rect 486 530 487 534
rect 491 530 492 534
rect 526 534 532 535
rect 486 529 492 530
rect 495 531 504 532
rect 463 526 472 527
rect 495 527 496 531
rect 503 527 504 531
rect 526 530 527 534
rect 531 530 532 534
rect 535 531 536 535
rect 543 531 544 535
rect 535 530 544 531
rect 574 534 580 535
rect 574 530 575 534
rect 579 530 580 534
rect 622 534 628 535
rect 526 529 532 530
rect 574 529 580 530
rect 583 531 589 532
rect 495 526 504 527
rect 583 527 584 531
rect 588 527 589 531
rect 622 530 623 534
rect 627 530 628 534
rect 631 531 632 535
rect 636 531 637 535
rect 631 530 637 531
rect 670 534 676 535
rect 670 530 671 534
rect 675 530 676 534
rect 710 534 716 535
rect 622 529 628 530
rect 670 529 676 530
rect 679 531 685 532
rect 583 526 589 527
rect 679 527 680 531
rect 684 527 685 531
rect 710 530 711 534
rect 715 530 716 534
rect 758 534 764 535
rect 710 529 716 530
rect 719 531 725 532
rect 679 526 685 527
rect 719 527 720 531
rect 724 530 725 531
rect 758 530 759 534
rect 763 530 764 534
rect 806 534 812 535
rect 724 528 746 530
rect 758 529 764 530
rect 767 531 773 532
rect 724 527 725 528
rect 719 526 725 527
rect 399 523 405 524
rect 399 522 400 523
rect 384 520 400 522
rect 367 518 373 519
rect 399 519 400 520
rect 404 519 405 523
rect 399 518 405 519
rect 431 523 437 524
rect 431 519 432 523
rect 436 522 437 523
rect 454 523 460 524
rect 454 522 455 523
rect 436 520 455 522
rect 436 519 437 520
rect 431 518 437 519
rect 454 519 455 520
rect 459 519 460 523
rect 454 518 460 519
rect 463 523 469 524
rect 463 519 464 523
rect 468 522 469 523
rect 486 523 492 524
rect 486 522 487 523
rect 468 520 487 522
rect 468 519 469 520
rect 463 518 469 519
rect 486 519 487 520
rect 491 519 492 523
rect 486 518 492 519
rect 495 523 501 524
rect 495 519 496 523
rect 500 522 501 523
rect 514 523 520 524
rect 514 522 515 523
rect 500 520 515 522
rect 500 519 501 520
rect 495 518 501 519
rect 514 519 515 520
rect 519 519 520 523
rect 514 518 520 519
rect 535 523 541 524
rect 535 519 536 523
rect 540 522 541 523
rect 584 522 586 526
rect 540 520 586 522
rect 540 519 541 520
rect 535 518 541 519
rect 631 519 637 520
rect 257 516 283 518
rect 279 515 285 516
rect 110 511 116 512
rect 110 507 111 511
rect 115 507 116 511
rect 279 511 280 515
rect 284 511 285 515
rect 279 510 285 511
rect 583 515 592 516
rect 583 511 584 515
rect 591 511 592 515
rect 631 515 632 519
rect 636 518 637 519
rect 679 518 681 526
rect 719 523 725 524
rect 719 519 720 523
rect 724 522 725 523
rect 730 523 736 524
rect 730 522 731 523
rect 724 520 731 522
rect 724 519 725 520
rect 719 518 725 519
rect 730 519 731 520
rect 735 519 736 523
rect 730 518 736 519
rect 744 518 746 528
rect 767 527 768 531
rect 772 527 773 531
rect 806 530 807 534
rect 811 530 812 534
rect 854 534 860 535
rect 806 529 812 530
rect 815 531 821 532
rect 767 526 773 527
rect 815 527 816 531
rect 820 530 821 531
rect 854 530 855 534
rect 859 530 860 534
rect 910 534 916 535
rect 820 528 842 530
rect 854 529 860 530
rect 863 531 869 532
rect 820 527 821 528
rect 815 526 821 527
rect 769 522 771 526
rect 815 523 821 524
rect 815 522 816 523
rect 769 520 816 522
rect 815 519 816 520
rect 820 519 821 523
rect 840 522 842 528
rect 863 527 864 531
rect 868 530 869 531
rect 910 530 911 534
rect 915 530 916 534
rect 966 534 972 535
rect 868 528 894 530
rect 910 529 916 530
rect 919 531 925 532
rect 868 527 869 528
rect 863 526 869 527
rect 863 523 869 524
rect 863 522 864 523
rect 840 520 864 522
rect 815 518 821 519
rect 863 519 864 520
rect 868 519 869 523
rect 892 522 894 528
rect 919 527 920 531
rect 924 530 925 531
rect 966 530 967 534
rect 971 530 972 534
rect 1022 534 1028 535
rect 924 528 950 530
rect 966 529 972 530
rect 975 531 981 532
rect 924 527 925 528
rect 919 526 925 527
rect 919 523 925 524
rect 919 522 920 523
rect 892 520 920 522
rect 863 518 869 519
rect 919 519 920 520
rect 924 519 925 523
rect 919 518 925 519
rect 948 518 950 528
rect 975 527 976 531
rect 980 527 981 531
rect 1022 530 1023 534
rect 1027 530 1028 534
rect 1031 531 1032 535
rect 1039 531 1040 535
rect 1031 530 1040 531
rect 1078 534 1084 535
rect 1078 530 1079 534
rect 1083 530 1084 534
rect 1126 534 1132 535
rect 1022 529 1028 530
rect 1078 529 1084 530
rect 1087 531 1093 532
rect 975 526 981 527
rect 1087 527 1088 531
rect 1092 530 1093 531
rect 1126 530 1127 534
rect 1131 530 1132 534
rect 1174 534 1180 535
rect 1092 528 1114 530
rect 1126 529 1132 530
rect 1135 531 1141 532
rect 1092 527 1093 528
rect 1087 526 1093 527
rect 977 522 979 526
rect 1031 523 1037 524
rect 1031 522 1032 523
rect 977 520 1032 522
rect 1031 519 1032 520
rect 1036 519 1037 523
rect 1031 518 1037 519
rect 1087 523 1096 524
rect 1087 519 1088 523
rect 1095 519 1096 523
rect 1112 522 1114 528
rect 1135 527 1136 531
rect 1140 530 1141 531
rect 1174 530 1175 534
rect 1179 530 1180 534
rect 1222 534 1228 535
rect 1140 528 1161 530
rect 1174 529 1180 530
rect 1183 531 1189 532
rect 1140 527 1141 528
rect 1135 526 1141 527
rect 1135 523 1141 524
rect 1135 522 1136 523
rect 1112 520 1136 522
rect 1087 518 1096 519
rect 1135 519 1136 520
rect 1140 519 1141 523
rect 1159 522 1161 528
rect 1183 527 1184 531
rect 1188 530 1189 531
rect 1222 530 1223 534
rect 1227 530 1228 534
rect 1270 534 1276 535
rect 1188 528 1211 530
rect 1222 529 1228 530
rect 1231 531 1237 532
rect 1188 527 1189 528
rect 1183 526 1189 527
rect 1183 523 1189 524
rect 1183 522 1184 523
rect 1159 520 1184 522
rect 1135 518 1141 519
rect 1183 519 1184 520
rect 1188 519 1189 523
rect 1209 522 1211 528
rect 1231 527 1232 531
rect 1236 530 1237 531
rect 1262 531 1268 532
rect 1262 530 1263 531
rect 1236 528 1263 530
rect 1236 527 1237 528
rect 1231 526 1237 527
rect 1262 527 1263 528
rect 1267 527 1268 531
rect 1270 530 1271 534
rect 1275 530 1276 534
rect 1279 531 1280 535
rect 1287 531 1288 535
rect 1279 530 1288 531
rect 1310 534 1316 535
rect 1310 530 1311 534
rect 1315 530 1316 534
rect 1350 534 1356 535
rect 1270 529 1276 530
rect 1310 529 1316 530
rect 1319 531 1325 532
rect 1262 526 1268 527
rect 1319 527 1320 531
rect 1324 527 1325 531
rect 1350 530 1351 534
rect 1355 530 1356 534
rect 1390 534 1396 535
rect 1350 529 1356 530
rect 1359 531 1365 532
rect 1319 526 1325 527
rect 1359 527 1360 531
rect 1364 527 1365 531
rect 1390 530 1391 534
rect 1395 530 1396 534
rect 1399 531 1400 535
rect 1404 531 1405 535
rect 1399 530 1405 531
rect 1414 534 1420 535
rect 1414 530 1415 534
rect 1419 530 1420 534
rect 1390 529 1396 530
rect 1414 529 1420 530
rect 1423 531 1429 532
rect 1359 526 1365 527
rect 1423 527 1424 531
rect 1428 527 1429 531
rect 1423 526 1429 527
rect 1446 529 1452 530
rect 1231 523 1237 524
rect 1231 522 1232 523
rect 1209 520 1232 522
rect 1183 518 1189 519
rect 1231 519 1232 520
rect 1236 519 1237 523
rect 1231 518 1237 519
rect 1279 523 1285 524
rect 1279 519 1280 523
rect 1284 522 1285 523
rect 1321 522 1323 526
rect 1284 520 1323 522
rect 1284 519 1285 520
rect 1279 518 1285 519
rect 1361 518 1363 526
rect 1399 523 1405 524
rect 1399 519 1400 523
rect 1404 522 1405 523
rect 1425 522 1427 526
rect 1446 525 1447 529
rect 1451 525 1452 529
rect 1446 524 1452 525
rect 1404 520 1427 522
rect 1404 519 1405 520
rect 1399 518 1405 519
rect 636 516 681 518
rect 744 516 771 518
rect 948 516 979 518
rect 1321 516 1363 518
rect 636 515 637 516
rect 631 514 637 515
rect 767 515 773 516
rect 583 510 592 511
rect 767 511 768 515
rect 772 511 773 515
rect 767 510 773 511
rect 975 515 981 516
rect 975 511 976 515
rect 980 511 981 515
rect 975 510 981 511
rect 1319 515 1325 516
rect 1319 511 1320 515
rect 1324 511 1325 515
rect 1319 510 1325 511
rect 1359 511 1368 512
rect 110 506 116 507
rect 222 508 228 509
rect 246 508 252 509
rect 270 508 276 509
rect 222 504 223 508
rect 227 504 228 508
rect 231 507 237 508
rect 231 504 232 507
rect 222 503 228 504
rect 230 503 232 504
rect 236 503 237 507
rect 246 504 247 508
rect 251 504 252 508
rect 246 503 252 504
rect 255 507 261 508
rect 255 503 256 507
rect 260 503 261 507
rect 270 504 271 508
rect 275 504 276 508
rect 270 503 276 504
rect 294 508 300 509
rect 294 504 295 508
rect 299 504 300 508
rect 294 503 300 504
rect 326 508 332 509
rect 326 504 327 508
rect 331 504 332 508
rect 326 503 332 504
rect 358 508 364 509
rect 358 504 359 508
rect 363 504 364 508
rect 358 503 364 504
rect 390 508 396 509
rect 390 504 391 508
rect 395 504 396 508
rect 390 503 396 504
rect 422 508 428 509
rect 422 504 423 508
rect 427 504 428 508
rect 422 503 428 504
rect 454 508 460 509
rect 454 504 455 508
rect 459 504 460 508
rect 454 503 460 504
rect 486 508 492 509
rect 486 504 487 508
rect 491 504 492 508
rect 486 503 492 504
rect 526 508 532 509
rect 526 504 527 508
rect 531 504 532 508
rect 526 503 532 504
rect 574 508 580 509
rect 574 504 575 508
rect 579 504 580 508
rect 574 503 580 504
rect 622 508 628 509
rect 622 504 623 508
rect 627 504 628 508
rect 622 503 628 504
rect 670 508 676 509
rect 710 508 716 509
rect 670 504 671 508
rect 675 504 676 508
rect 679 507 685 508
rect 679 504 680 507
rect 670 503 676 504
rect 678 503 680 504
rect 684 503 685 507
rect 710 504 711 508
rect 715 504 716 508
rect 710 503 716 504
rect 758 508 764 509
rect 758 504 759 508
rect 763 504 764 508
rect 758 503 764 504
rect 806 508 812 509
rect 806 504 807 508
rect 811 504 812 508
rect 806 503 812 504
rect 854 508 860 509
rect 854 504 855 508
rect 859 504 860 508
rect 854 503 860 504
rect 910 508 916 509
rect 910 504 911 508
rect 915 504 916 508
rect 910 503 916 504
rect 966 508 972 509
rect 966 504 967 508
rect 971 504 972 508
rect 966 503 972 504
rect 1022 508 1028 509
rect 1022 504 1023 508
rect 1027 504 1028 508
rect 1022 503 1028 504
rect 1078 508 1084 509
rect 1078 504 1079 508
rect 1083 504 1084 508
rect 1078 503 1084 504
rect 1126 508 1132 509
rect 1126 504 1127 508
rect 1131 504 1132 508
rect 1126 503 1132 504
rect 1174 508 1180 509
rect 1174 504 1175 508
rect 1179 504 1180 508
rect 1174 503 1180 504
rect 1222 508 1228 509
rect 1222 504 1223 508
rect 1227 504 1228 508
rect 1222 503 1228 504
rect 1270 508 1276 509
rect 1270 504 1271 508
rect 1275 504 1276 508
rect 1270 503 1276 504
rect 1310 508 1316 509
rect 1310 504 1311 508
rect 1315 504 1316 508
rect 1310 503 1316 504
rect 1350 508 1356 509
rect 1350 504 1351 508
rect 1355 504 1356 508
rect 1359 507 1360 511
rect 1367 507 1368 511
rect 1446 511 1452 512
rect 1359 506 1368 507
rect 1390 508 1396 509
rect 1350 503 1356 504
rect 1390 504 1391 508
rect 1395 504 1396 508
rect 1390 503 1396 504
rect 1414 508 1420 509
rect 1414 504 1415 508
rect 1419 504 1420 508
rect 1414 503 1420 504
rect 1423 507 1432 508
rect 1423 503 1424 507
rect 1431 503 1432 507
rect 1446 507 1447 511
rect 1451 507 1452 511
rect 1446 506 1452 507
rect 230 499 231 503
rect 235 502 237 503
rect 255 502 261 503
rect 235 499 236 502
rect 230 498 236 499
rect 238 499 244 500
rect 134 496 140 497
rect 110 493 116 494
rect 110 489 111 493
rect 115 489 116 493
rect 134 492 135 496
rect 139 492 140 496
rect 134 491 140 492
rect 158 496 164 497
rect 158 492 159 496
rect 163 492 164 496
rect 158 491 164 492
rect 182 496 188 497
rect 182 492 183 496
rect 187 492 188 496
rect 182 491 188 492
rect 222 496 228 497
rect 222 492 223 496
rect 227 492 228 496
rect 238 495 239 499
rect 243 498 244 499
rect 257 498 259 502
rect 678 499 679 503
rect 683 502 685 503
rect 1423 502 1432 503
rect 683 499 684 502
rect 678 498 684 499
rect 243 496 259 498
rect 270 496 276 497
rect 243 495 244 496
rect 238 494 244 495
rect 222 491 228 492
rect 270 492 271 496
rect 275 492 276 496
rect 270 491 276 492
rect 318 496 324 497
rect 318 492 319 496
rect 323 492 324 496
rect 318 491 324 492
rect 374 496 380 497
rect 374 492 375 496
rect 379 492 380 496
rect 374 491 380 492
rect 430 496 436 497
rect 430 492 431 496
rect 435 492 436 496
rect 430 491 436 492
rect 486 496 492 497
rect 486 492 487 496
rect 491 492 492 496
rect 486 491 492 492
rect 542 496 548 497
rect 542 492 543 496
rect 547 492 548 496
rect 542 491 548 492
rect 590 496 596 497
rect 590 492 591 496
rect 595 492 596 496
rect 590 491 596 492
rect 630 496 636 497
rect 630 492 631 496
rect 635 492 636 496
rect 630 491 636 492
rect 662 496 668 497
rect 662 492 663 496
rect 667 492 668 496
rect 662 491 668 492
rect 686 496 692 497
rect 686 492 687 496
rect 691 492 692 496
rect 686 491 692 492
rect 718 496 724 497
rect 718 492 719 496
rect 723 492 724 496
rect 718 491 724 492
rect 758 496 764 497
rect 758 492 759 496
rect 763 492 764 496
rect 758 491 764 492
rect 798 496 804 497
rect 798 492 799 496
rect 803 492 804 496
rect 798 491 804 492
rect 846 496 852 497
rect 846 492 847 496
rect 851 492 852 496
rect 846 491 852 492
rect 902 496 908 497
rect 902 492 903 496
rect 907 492 908 496
rect 902 491 908 492
rect 950 496 956 497
rect 950 492 951 496
rect 955 492 956 496
rect 950 491 956 492
rect 998 496 1004 497
rect 998 492 999 496
rect 1003 492 1004 496
rect 998 491 1004 492
rect 1046 496 1052 497
rect 1046 492 1047 496
rect 1051 492 1052 496
rect 1046 491 1052 492
rect 1094 496 1100 497
rect 1094 492 1095 496
rect 1099 492 1100 496
rect 1094 491 1100 492
rect 1142 496 1148 497
rect 1142 492 1143 496
rect 1147 492 1148 496
rect 1142 491 1148 492
rect 1198 496 1204 497
rect 1198 492 1199 496
rect 1203 492 1204 496
rect 1198 491 1204 492
rect 1254 496 1260 497
rect 1254 492 1255 496
rect 1259 492 1260 496
rect 1254 491 1260 492
rect 1310 496 1316 497
rect 1310 492 1311 496
rect 1315 492 1316 496
rect 1310 491 1316 492
rect 1374 496 1380 497
rect 1374 492 1375 496
rect 1379 492 1380 496
rect 1374 491 1380 492
rect 1414 496 1420 497
rect 1414 492 1415 496
rect 1419 492 1420 496
rect 1414 491 1420 492
rect 1446 493 1452 494
rect 110 488 116 489
rect 1446 489 1447 493
rect 1451 489 1452 493
rect 1446 488 1452 489
rect 143 487 149 488
rect 143 483 144 487
rect 148 486 149 487
rect 362 487 368 488
rect 362 486 363 487
rect 148 484 363 486
rect 148 483 149 484
rect 143 482 149 483
rect 362 483 363 484
rect 367 483 368 487
rect 362 482 368 483
rect 439 487 445 488
rect 439 483 440 487
rect 444 486 445 487
rect 498 487 504 488
rect 498 486 499 487
rect 444 484 499 486
rect 444 483 445 484
rect 439 482 445 483
rect 498 483 499 484
rect 503 483 504 487
rect 498 482 504 483
rect 551 487 557 488
rect 551 483 552 487
rect 556 486 557 487
rect 602 487 608 488
rect 602 486 603 487
rect 556 484 603 486
rect 556 483 557 484
rect 551 482 557 483
rect 602 483 603 484
rect 607 483 608 487
rect 602 482 608 483
rect 639 487 645 488
rect 639 483 640 487
rect 644 486 645 487
rect 671 487 677 488
rect 644 484 662 486
rect 644 483 645 484
rect 639 482 645 483
rect 167 479 173 480
rect 167 478 168 479
rect 152 476 168 478
rect 110 475 116 476
rect 110 471 111 475
rect 115 471 116 475
rect 143 471 149 472
rect 110 470 116 471
rect 134 470 140 471
rect 134 466 135 470
rect 139 466 140 470
rect 143 467 144 471
rect 148 470 149 471
rect 152 470 154 476
rect 167 475 168 476
rect 172 475 173 479
rect 191 479 197 480
rect 191 478 192 479
rect 167 474 173 475
rect 176 476 192 478
rect 167 471 173 472
rect 148 468 154 470
rect 158 470 164 471
rect 148 467 149 468
rect 143 466 149 467
rect 158 466 159 470
rect 163 466 164 470
rect 167 467 168 471
rect 172 470 173 471
rect 176 470 178 476
rect 191 475 192 476
rect 196 475 197 479
rect 231 479 237 480
rect 231 478 232 479
rect 191 474 197 475
rect 212 476 232 478
rect 191 471 197 472
rect 172 468 178 470
rect 182 470 188 471
rect 172 467 173 468
rect 167 466 173 467
rect 182 466 183 470
rect 187 466 188 470
rect 191 467 192 471
rect 196 470 197 471
rect 212 470 214 476
rect 231 475 232 476
rect 236 475 237 479
rect 279 479 285 480
rect 279 478 280 479
rect 231 474 237 475
rect 257 476 280 478
rect 231 471 237 472
rect 196 468 214 470
rect 222 470 228 471
rect 196 467 197 468
rect 191 466 197 467
rect 222 466 223 470
rect 227 466 228 470
rect 231 467 232 471
rect 236 470 237 471
rect 257 470 259 476
rect 279 475 280 476
rect 284 475 285 479
rect 327 479 333 480
rect 327 478 328 479
rect 279 474 285 475
rect 300 476 328 478
rect 279 471 285 472
rect 236 468 259 470
rect 270 470 276 471
rect 236 467 237 468
rect 231 466 237 467
rect 270 466 271 470
rect 275 466 276 470
rect 279 467 280 471
rect 284 470 285 471
rect 300 470 302 476
rect 327 475 328 476
rect 332 475 333 479
rect 383 479 389 480
rect 383 478 384 479
rect 327 474 333 475
rect 356 476 384 478
rect 327 471 333 472
rect 284 468 302 470
rect 318 470 324 471
rect 284 467 285 468
rect 279 466 285 467
rect 318 466 319 470
rect 323 466 324 470
rect 327 467 328 471
rect 332 470 333 471
rect 356 470 358 476
rect 383 475 384 476
rect 388 475 389 479
rect 383 474 389 475
rect 446 479 452 480
rect 446 475 447 479
rect 451 478 452 479
rect 495 479 501 480
rect 495 478 496 479
rect 451 476 496 478
rect 451 475 452 476
rect 446 474 452 475
rect 495 475 496 476
rect 500 475 501 479
rect 495 474 501 475
rect 599 479 605 480
rect 599 475 600 479
rect 604 478 605 479
rect 660 478 662 484
rect 671 483 672 487
rect 676 486 677 487
rect 695 487 701 488
rect 676 484 690 486
rect 676 483 677 484
rect 671 482 677 483
rect 678 479 684 480
rect 678 478 679 479
rect 604 476 642 478
rect 660 476 679 478
rect 604 475 605 476
rect 599 474 605 475
rect 640 472 642 476
rect 678 475 679 476
rect 683 475 684 479
rect 688 478 690 484
rect 695 483 696 487
rect 700 486 701 487
rect 730 487 736 488
rect 730 486 731 487
rect 700 484 731 486
rect 700 483 701 484
rect 695 482 701 483
rect 730 483 731 484
rect 735 483 736 487
rect 730 482 736 483
rect 767 487 773 488
rect 767 483 768 487
rect 772 486 773 487
rect 810 487 816 488
rect 810 486 811 487
rect 772 484 811 486
rect 772 483 773 484
rect 767 482 773 483
rect 810 483 811 484
rect 815 483 816 487
rect 810 482 816 483
rect 818 487 824 488
rect 818 483 819 487
rect 823 486 824 487
rect 894 487 900 488
rect 894 486 895 487
rect 823 484 895 486
rect 823 483 824 484
rect 818 482 824 483
rect 894 483 895 484
rect 899 483 900 487
rect 894 482 900 483
rect 911 487 917 488
rect 911 483 912 487
rect 916 486 917 487
rect 962 487 968 488
rect 962 486 963 487
rect 916 484 963 486
rect 916 483 917 484
rect 911 482 917 483
rect 962 483 963 484
rect 967 483 968 487
rect 962 482 968 483
rect 1007 487 1013 488
rect 1007 483 1008 487
rect 1012 486 1013 487
rect 1058 487 1064 488
rect 1058 486 1059 487
rect 1012 484 1059 486
rect 1012 483 1013 484
rect 1007 482 1013 483
rect 1058 483 1059 484
rect 1063 483 1064 487
rect 1058 482 1064 483
rect 1103 487 1109 488
rect 1103 483 1104 487
rect 1108 486 1109 487
rect 1154 487 1160 488
rect 1154 486 1155 487
rect 1108 484 1155 486
rect 1108 483 1109 484
rect 1103 482 1109 483
rect 1154 483 1155 484
rect 1159 483 1160 487
rect 1154 482 1160 483
rect 1207 487 1213 488
rect 1207 483 1208 487
rect 1212 486 1213 487
rect 1266 487 1272 488
rect 1266 486 1267 487
rect 1212 484 1267 486
rect 1212 483 1213 484
rect 1207 482 1213 483
rect 1266 483 1267 484
rect 1271 483 1272 487
rect 1266 482 1272 483
rect 1278 487 1284 488
rect 1278 483 1279 487
rect 1283 486 1284 487
rect 1319 487 1325 488
rect 1319 486 1320 487
rect 1283 484 1320 486
rect 1283 483 1284 484
rect 1278 482 1284 483
rect 1319 483 1320 484
rect 1324 483 1325 487
rect 1319 482 1325 483
rect 1382 483 1389 484
rect 727 479 733 480
rect 688 476 698 478
rect 678 474 684 475
rect 696 472 698 476
rect 727 475 728 479
rect 732 478 733 479
rect 807 479 813 480
rect 732 476 750 478
rect 732 475 733 476
rect 727 474 733 475
rect 495 471 504 472
rect 599 471 608 472
rect 639 471 645 472
rect 695 471 701 472
rect 727 471 736 472
rect 332 468 358 470
rect 374 470 380 471
rect 332 467 333 468
rect 327 466 333 467
rect 374 466 375 470
rect 379 466 380 470
rect 430 470 436 471
rect 134 465 140 466
rect 158 465 164 466
rect 182 465 188 466
rect 222 465 228 466
rect 270 465 276 466
rect 318 465 324 466
rect 374 465 380 466
rect 383 467 389 468
rect 230 463 236 464
rect 230 459 231 463
rect 235 462 236 463
rect 383 463 384 467
rect 388 463 389 467
rect 430 466 431 470
rect 435 466 436 470
rect 486 470 492 471
rect 430 465 436 466
rect 439 467 448 468
rect 383 462 389 463
rect 439 463 440 467
rect 447 463 448 467
rect 486 466 487 470
rect 491 466 492 470
rect 495 467 496 471
rect 503 467 504 471
rect 495 466 504 467
rect 542 470 548 471
rect 542 466 543 470
rect 547 466 548 470
rect 590 470 596 471
rect 486 465 492 466
rect 542 465 548 466
rect 551 467 557 468
rect 439 462 448 463
rect 551 463 552 467
rect 556 466 557 467
rect 590 466 591 470
rect 595 466 596 470
rect 599 467 600 471
rect 607 467 608 471
rect 599 466 608 467
rect 630 470 636 471
rect 630 466 631 470
rect 635 466 636 470
rect 639 467 640 471
rect 644 467 645 471
rect 639 466 645 467
rect 662 470 668 471
rect 662 466 663 470
rect 667 466 668 470
rect 686 470 692 471
rect 556 464 586 466
rect 590 465 596 466
rect 630 465 636 466
rect 662 465 668 466
rect 671 467 677 468
rect 556 463 557 464
rect 551 462 557 463
rect 584 462 586 464
rect 654 463 660 464
rect 654 462 655 463
rect 235 460 386 462
rect 584 460 655 462
rect 235 459 236 460
rect 230 458 236 459
rect 654 459 655 460
rect 659 459 660 463
rect 671 463 672 467
rect 676 466 677 467
rect 686 466 687 470
rect 691 466 692 470
rect 695 467 696 471
rect 700 467 701 471
rect 695 466 701 467
rect 718 470 724 471
rect 718 466 719 470
rect 723 466 724 470
rect 727 467 728 471
rect 735 467 736 471
rect 727 466 736 467
rect 676 464 682 466
rect 686 465 692 466
rect 718 465 724 466
rect 676 463 677 464
rect 671 462 677 463
rect 680 462 682 464
rect 710 463 716 464
rect 710 462 711 463
rect 680 460 711 462
rect 654 458 660 459
rect 710 459 711 460
rect 715 459 716 463
rect 748 462 750 476
rect 807 475 808 479
rect 812 478 813 479
rect 855 479 861 480
rect 812 476 843 478
rect 812 475 813 476
rect 807 474 813 475
rect 807 471 816 472
rect 758 470 764 471
rect 758 466 759 470
rect 763 466 764 470
rect 798 470 804 471
rect 758 465 764 466
rect 767 467 773 468
rect 767 463 768 467
rect 772 463 773 467
rect 798 466 799 470
rect 803 466 804 470
rect 807 467 808 471
rect 815 467 816 471
rect 807 466 816 467
rect 798 465 804 466
rect 767 462 773 463
rect 841 462 843 476
rect 855 475 856 479
rect 860 478 861 479
rect 918 479 924 480
rect 860 476 915 478
rect 860 475 861 476
rect 855 474 861 475
rect 913 472 915 476
rect 918 475 919 479
rect 923 478 924 479
rect 959 479 965 480
rect 959 478 960 479
rect 923 476 960 478
rect 923 475 924 476
rect 918 474 924 475
rect 959 475 960 476
rect 964 475 965 479
rect 959 474 965 475
rect 1055 479 1061 480
rect 1055 475 1056 479
rect 1060 478 1061 479
rect 1151 479 1157 480
rect 1060 476 1082 478
rect 1060 475 1061 476
rect 1055 474 1061 475
rect 911 471 917 472
rect 959 471 968 472
rect 1055 471 1064 472
rect 846 470 852 471
rect 846 466 847 470
rect 851 466 852 470
rect 902 470 908 471
rect 846 465 852 466
rect 855 467 861 468
rect 855 463 856 467
rect 860 463 861 467
rect 902 466 903 470
rect 907 466 908 470
rect 911 467 912 471
rect 916 467 917 471
rect 911 466 917 467
rect 950 470 956 471
rect 950 466 951 470
rect 955 466 956 470
rect 959 467 960 471
rect 967 467 968 471
rect 959 466 968 467
rect 998 470 1004 471
rect 998 466 999 470
rect 1003 466 1004 470
rect 1046 470 1052 471
rect 902 465 908 466
rect 950 465 956 466
rect 998 465 1004 466
rect 1007 467 1013 468
rect 855 462 861 463
rect 922 463 928 464
rect 748 460 771 462
rect 841 460 858 462
rect 710 458 716 459
rect 922 459 923 463
rect 927 462 928 463
rect 1007 463 1008 467
rect 1012 466 1013 467
rect 1023 467 1029 468
rect 1023 466 1024 467
rect 1012 464 1024 466
rect 1012 463 1013 464
rect 1007 462 1013 463
rect 1023 463 1024 464
rect 1028 463 1029 467
rect 1046 466 1047 470
rect 1051 466 1052 470
rect 1055 467 1056 471
rect 1063 467 1064 471
rect 1055 466 1064 467
rect 1046 465 1052 466
rect 1023 462 1029 463
rect 1080 462 1082 476
rect 1151 475 1152 479
rect 1156 478 1157 479
rect 1263 479 1269 480
rect 1156 476 1195 478
rect 1156 475 1157 476
rect 1151 474 1157 475
rect 1151 471 1160 472
rect 1094 470 1100 471
rect 1094 466 1095 470
rect 1099 466 1100 470
rect 1142 470 1148 471
rect 1094 465 1100 466
rect 1103 467 1109 468
rect 1103 463 1104 467
rect 1108 463 1109 467
rect 1142 466 1143 470
rect 1147 466 1148 470
rect 1151 467 1152 471
rect 1159 467 1160 471
rect 1151 466 1160 467
rect 1142 465 1148 466
rect 1103 462 1109 463
rect 1193 462 1195 476
rect 1263 475 1264 479
rect 1268 478 1269 479
rect 1382 479 1383 483
rect 1388 479 1389 483
rect 1382 478 1389 479
rect 1423 479 1429 480
rect 1423 478 1424 479
rect 1268 476 1294 478
rect 1268 475 1269 476
rect 1263 474 1269 475
rect 1263 471 1272 472
rect 1198 470 1204 471
rect 1198 466 1199 470
rect 1203 466 1204 470
rect 1254 470 1260 471
rect 1198 465 1204 466
rect 1207 467 1213 468
rect 1207 463 1208 467
rect 1212 463 1213 467
rect 1254 466 1255 470
rect 1259 466 1260 470
rect 1263 467 1264 471
rect 1271 467 1272 471
rect 1263 466 1272 467
rect 1254 465 1260 466
rect 1207 462 1213 463
rect 1292 462 1294 476
rect 1404 476 1424 478
rect 1383 471 1389 472
rect 1310 470 1316 471
rect 1310 466 1311 470
rect 1315 466 1316 470
rect 1374 470 1380 471
rect 1310 465 1316 466
rect 1319 467 1325 468
rect 1319 463 1320 467
rect 1324 463 1325 467
rect 1374 466 1375 470
rect 1379 466 1380 470
rect 1383 467 1384 471
rect 1388 470 1389 471
rect 1404 470 1406 476
rect 1423 475 1424 476
rect 1428 475 1429 479
rect 1423 474 1429 475
rect 1446 475 1452 476
rect 1423 471 1432 472
rect 1388 468 1406 470
rect 1414 470 1420 471
rect 1388 467 1389 468
rect 1383 466 1389 467
rect 1414 466 1415 470
rect 1419 466 1420 470
rect 1423 467 1424 471
rect 1431 467 1432 471
rect 1446 471 1447 475
rect 1451 471 1452 475
rect 1446 470 1452 471
rect 1423 466 1432 467
rect 1374 465 1380 466
rect 1414 465 1420 466
rect 1319 462 1325 463
rect 927 460 954 462
rect 1080 460 1106 462
rect 1193 460 1211 462
rect 1292 460 1323 462
rect 927 459 928 460
rect 922 458 928 459
rect 952 456 954 460
rect 359 455 368 456
rect 799 455 805 456
rect 134 454 140 455
rect 134 450 135 454
rect 139 450 140 454
rect 158 454 164 455
rect 110 449 116 450
rect 134 449 140 450
rect 143 451 149 452
rect 110 445 111 449
rect 115 445 116 449
rect 143 447 144 451
rect 148 447 149 451
rect 158 450 159 454
rect 163 450 164 454
rect 190 454 196 455
rect 158 449 164 450
rect 167 451 173 452
rect 143 446 149 447
rect 167 447 168 451
rect 172 450 173 451
rect 190 450 191 454
rect 195 450 196 454
rect 238 454 244 455
rect 172 448 187 450
rect 190 449 196 450
rect 199 451 205 452
rect 172 447 173 448
rect 167 446 173 447
rect 110 444 116 445
rect 145 442 147 446
rect 167 443 173 444
rect 167 442 168 443
rect 145 440 168 442
rect 126 439 132 440
rect 126 435 127 439
rect 131 438 132 439
rect 167 439 168 440
rect 172 439 173 443
rect 185 442 187 448
rect 199 447 200 451
rect 204 450 205 451
rect 238 450 239 454
rect 243 450 244 454
rect 294 454 300 455
rect 204 448 235 450
rect 238 449 244 450
rect 247 451 253 452
rect 204 447 205 448
rect 199 446 205 447
rect 199 443 205 444
rect 199 442 200 443
rect 185 440 200 442
rect 167 438 173 439
rect 199 439 200 440
rect 204 439 205 443
rect 233 442 235 448
rect 247 447 248 451
rect 252 450 253 451
rect 294 450 295 454
rect 299 450 300 454
rect 350 454 356 455
rect 252 448 291 450
rect 294 449 300 450
rect 303 451 309 452
rect 252 447 253 448
rect 247 446 253 447
rect 247 443 253 444
rect 247 442 248 443
rect 233 440 248 442
rect 199 438 205 439
rect 247 439 248 440
rect 252 439 253 443
rect 289 442 291 448
rect 303 447 304 451
rect 308 450 309 451
rect 350 450 351 454
rect 355 450 356 454
rect 359 451 360 455
rect 367 451 368 455
rect 359 450 368 451
rect 414 454 420 455
rect 414 450 415 454
rect 419 450 420 454
rect 478 454 484 455
rect 308 448 347 450
rect 350 449 356 450
rect 414 449 420 450
rect 423 451 429 452
rect 308 447 309 448
rect 303 446 309 447
rect 303 443 309 444
rect 303 442 304 443
rect 289 440 304 442
rect 247 438 253 439
rect 303 439 304 440
rect 308 439 309 443
rect 345 442 347 448
rect 423 447 424 451
rect 428 450 429 451
rect 478 450 479 454
rect 483 450 484 454
rect 542 454 548 455
rect 428 448 458 450
rect 478 449 484 450
rect 487 451 493 452
rect 428 447 429 448
rect 423 446 429 447
rect 359 443 365 444
rect 359 442 360 443
rect 345 440 360 442
rect 303 438 309 439
rect 359 439 360 440
rect 364 439 365 443
rect 359 438 365 439
rect 423 443 429 444
rect 423 439 424 443
rect 428 442 429 443
rect 442 443 448 444
rect 442 442 443 443
rect 428 440 443 442
rect 428 439 429 440
rect 423 438 429 439
rect 442 439 443 440
rect 447 439 448 443
rect 456 442 458 448
rect 487 447 488 451
rect 492 450 493 451
rect 542 450 543 454
rect 547 450 548 454
rect 606 454 612 455
rect 492 448 522 450
rect 542 449 548 450
rect 551 451 557 452
rect 492 447 493 448
rect 487 446 493 447
rect 487 443 493 444
rect 487 442 488 443
rect 456 440 488 442
rect 442 438 448 439
rect 487 439 488 440
rect 492 439 493 443
rect 520 442 522 448
rect 551 447 552 451
rect 556 450 557 451
rect 606 450 607 454
rect 611 450 612 454
rect 670 454 676 455
rect 556 448 586 450
rect 606 449 612 450
rect 615 451 624 452
rect 556 447 557 448
rect 551 446 557 447
rect 551 443 557 444
rect 551 442 552 443
rect 520 440 552 442
rect 487 438 493 439
rect 551 439 552 440
rect 556 439 557 443
rect 584 442 586 448
rect 615 447 616 451
rect 623 447 624 451
rect 670 450 671 454
rect 675 450 676 454
rect 734 454 740 455
rect 670 449 676 450
rect 679 451 688 452
rect 615 446 624 447
rect 679 447 680 451
rect 687 447 688 451
rect 734 450 735 454
rect 739 450 740 454
rect 790 454 796 455
rect 734 449 740 450
rect 743 451 749 452
rect 679 446 688 447
rect 743 447 744 451
rect 748 447 749 451
rect 790 450 791 454
rect 795 450 796 454
rect 799 451 800 455
rect 804 454 805 455
rect 818 455 824 456
rect 951 455 957 456
rect 818 454 819 455
rect 804 452 819 454
rect 804 451 805 452
rect 799 450 805 451
rect 818 451 819 452
rect 823 451 824 455
rect 818 450 824 451
rect 838 454 844 455
rect 838 450 839 454
rect 843 450 844 454
rect 878 454 884 455
rect 790 449 796 450
rect 838 449 844 450
rect 847 451 856 452
rect 743 446 749 447
rect 847 447 848 451
rect 855 447 856 451
rect 878 450 879 454
rect 883 450 884 454
rect 910 454 916 455
rect 878 449 884 450
rect 887 451 896 452
rect 847 446 856 447
rect 887 447 888 451
rect 895 447 896 451
rect 910 450 911 454
rect 915 450 916 454
rect 942 454 948 455
rect 910 449 916 450
rect 919 451 925 452
rect 887 446 896 447
rect 919 447 920 451
rect 924 447 925 451
rect 942 450 943 454
rect 947 450 948 454
rect 951 451 952 455
rect 956 451 957 455
rect 951 450 957 451
rect 966 454 972 455
rect 966 450 967 454
rect 971 450 972 454
rect 998 454 1004 455
rect 942 449 948 450
rect 966 449 972 450
rect 975 451 981 452
rect 919 446 925 447
rect 975 447 976 451
rect 980 447 981 451
rect 998 450 999 454
rect 1003 450 1004 454
rect 1030 454 1036 455
rect 998 449 1004 450
rect 1007 451 1013 452
rect 975 446 981 447
rect 1007 447 1008 451
rect 1012 450 1013 451
rect 1022 451 1028 452
rect 1022 450 1023 451
rect 1012 448 1023 450
rect 1012 447 1013 448
rect 1007 446 1013 447
rect 1022 447 1023 448
rect 1027 447 1028 451
rect 1030 450 1031 454
rect 1035 450 1036 454
rect 1070 454 1076 455
rect 1030 449 1036 450
rect 1039 451 1045 452
rect 1022 446 1028 447
rect 1039 447 1040 451
rect 1044 447 1045 451
rect 1070 450 1071 454
rect 1075 450 1076 454
rect 1118 454 1124 455
rect 1070 449 1076 450
rect 1079 451 1085 452
rect 1039 446 1045 447
rect 1079 447 1080 451
rect 1084 447 1085 451
rect 1118 450 1119 454
rect 1123 450 1124 454
rect 1174 454 1180 455
rect 1118 449 1124 450
rect 1127 451 1133 452
rect 1079 446 1085 447
rect 1127 447 1128 451
rect 1132 447 1133 451
rect 1174 450 1175 454
rect 1179 450 1180 454
rect 1238 454 1244 455
rect 1174 449 1180 450
rect 1183 451 1189 452
rect 1127 446 1133 447
rect 1183 447 1184 451
rect 1188 447 1189 451
rect 1238 450 1239 454
rect 1243 450 1244 454
rect 1302 454 1308 455
rect 1238 449 1244 450
rect 1247 451 1253 452
rect 1183 446 1189 447
rect 1247 447 1248 451
rect 1252 447 1253 451
rect 1302 450 1303 454
rect 1307 450 1308 454
rect 1366 454 1372 455
rect 1302 449 1308 450
rect 1311 451 1317 452
rect 1247 446 1253 447
rect 1311 447 1312 451
rect 1316 450 1317 451
rect 1330 451 1336 452
rect 1330 450 1331 451
rect 1316 448 1331 450
rect 1316 447 1317 448
rect 1311 446 1317 447
rect 1330 447 1331 448
rect 1335 447 1336 451
rect 1366 450 1367 454
rect 1371 450 1372 454
rect 1414 454 1420 455
rect 1366 449 1372 450
rect 1375 451 1381 452
rect 1330 446 1336 447
rect 1375 447 1376 451
rect 1380 447 1381 451
rect 1414 450 1415 454
rect 1419 450 1420 454
rect 1414 449 1420 450
rect 1423 451 1429 452
rect 1375 446 1381 447
rect 1423 447 1424 451
rect 1428 447 1429 451
rect 1423 446 1429 447
rect 1446 449 1452 450
rect 615 443 621 444
rect 615 442 616 443
rect 584 440 616 442
rect 551 438 557 439
rect 615 439 616 440
rect 620 439 621 443
rect 615 438 621 439
rect 679 443 685 444
rect 679 439 680 443
rect 684 442 685 443
rect 744 442 746 446
rect 684 440 746 442
rect 799 443 805 444
rect 684 439 685 440
rect 679 438 685 439
rect 799 439 800 443
rect 804 442 805 443
rect 838 443 844 444
rect 838 442 839 443
rect 804 440 839 442
rect 804 439 805 440
rect 799 438 805 439
rect 838 439 839 440
rect 843 439 844 443
rect 838 438 844 439
rect 847 443 853 444
rect 847 439 848 443
rect 852 442 853 443
rect 878 443 884 444
rect 878 442 879 443
rect 852 440 879 442
rect 852 439 853 440
rect 847 438 853 439
rect 878 439 879 440
rect 883 439 884 443
rect 878 438 884 439
rect 887 443 893 444
rect 887 439 888 443
rect 892 442 893 443
rect 919 442 921 446
rect 892 440 921 442
rect 951 443 957 444
rect 892 439 893 440
rect 887 438 893 439
rect 951 439 952 443
rect 956 442 957 443
rect 977 442 979 446
rect 956 440 979 442
rect 1007 443 1013 444
rect 956 439 957 440
rect 951 438 957 439
rect 1007 439 1008 443
rect 1012 442 1013 443
rect 1041 442 1043 446
rect 1012 440 1043 442
rect 1012 439 1013 440
rect 1007 438 1013 439
rect 1080 438 1082 446
rect 1128 438 1130 446
rect 1184 438 1186 446
rect 1248 438 1250 446
rect 1375 443 1381 444
rect 1375 439 1376 443
rect 1380 442 1381 443
rect 1425 442 1427 446
rect 1446 445 1447 449
rect 1451 445 1452 449
rect 1446 444 1452 445
rect 1380 440 1427 442
rect 1380 439 1381 440
rect 1375 438 1381 439
rect 131 436 147 438
rect 712 436 746 438
rect 1041 436 1082 438
rect 1104 436 1130 438
rect 1156 436 1186 438
rect 1216 436 1250 438
rect 131 435 132 436
rect 126 434 132 435
rect 143 435 149 436
rect 110 431 116 432
rect 110 427 111 431
rect 115 427 116 431
rect 143 431 144 435
rect 148 431 149 435
rect 143 430 149 431
rect 710 435 716 436
rect 710 431 711 435
rect 715 431 716 435
rect 710 430 716 431
rect 743 435 749 436
rect 743 431 744 435
rect 748 431 749 435
rect 743 430 749 431
rect 919 435 928 436
rect 919 431 920 435
rect 927 431 928 435
rect 919 430 928 431
rect 1039 435 1045 436
rect 1039 431 1040 435
rect 1044 431 1045 435
rect 1039 430 1045 431
rect 1079 431 1085 432
rect 110 426 116 427
rect 134 428 140 429
rect 134 424 135 428
rect 139 424 140 428
rect 134 423 140 424
rect 158 428 164 429
rect 158 424 159 428
rect 163 424 164 428
rect 158 423 164 424
rect 190 428 196 429
rect 190 424 191 428
rect 195 424 196 428
rect 190 423 196 424
rect 238 428 244 429
rect 238 424 239 428
rect 243 424 244 428
rect 238 423 244 424
rect 294 428 300 429
rect 294 424 295 428
rect 299 424 300 428
rect 294 423 300 424
rect 350 428 356 429
rect 350 424 351 428
rect 355 424 356 428
rect 350 423 356 424
rect 414 428 420 429
rect 414 424 415 428
rect 419 424 420 428
rect 414 423 420 424
rect 478 428 484 429
rect 478 424 479 428
rect 483 424 484 428
rect 478 423 484 424
rect 542 428 548 429
rect 542 424 543 428
rect 547 424 548 428
rect 542 423 548 424
rect 606 428 612 429
rect 606 424 607 428
rect 611 424 612 428
rect 606 423 612 424
rect 670 428 676 429
rect 670 424 671 428
rect 675 424 676 428
rect 670 423 676 424
rect 734 428 740 429
rect 734 424 735 428
rect 739 424 740 428
rect 734 423 740 424
rect 790 428 796 429
rect 790 424 791 428
rect 795 424 796 428
rect 790 423 796 424
rect 838 428 844 429
rect 838 424 839 428
rect 843 424 844 428
rect 838 423 844 424
rect 878 428 884 429
rect 878 424 879 428
rect 883 424 884 428
rect 878 423 884 424
rect 910 428 916 429
rect 910 424 911 428
rect 915 424 916 428
rect 910 423 916 424
rect 942 428 948 429
rect 942 424 943 428
rect 947 424 948 428
rect 942 423 948 424
rect 966 428 972 429
rect 998 428 1004 429
rect 966 424 967 428
rect 971 424 972 428
rect 966 423 972 424
rect 975 427 981 428
rect 975 423 976 427
rect 980 426 981 427
rect 986 427 992 428
rect 986 426 987 427
rect 980 424 987 426
rect 980 423 981 424
rect 975 422 981 423
rect 986 423 987 424
rect 991 423 992 427
rect 998 424 999 428
rect 1003 424 1004 428
rect 998 423 1004 424
rect 1030 428 1036 429
rect 1030 424 1031 428
rect 1035 424 1036 428
rect 1030 423 1036 424
rect 1070 428 1076 429
rect 1070 424 1071 428
rect 1075 424 1076 428
rect 1079 427 1080 431
rect 1084 430 1085 431
rect 1104 430 1106 436
rect 1084 428 1106 430
rect 1127 431 1133 432
rect 1118 428 1124 429
rect 1084 427 1085 428
rect 1079 426 1085 427
rect 1070 423 1076 424
rect 1118 424 1119 428
rect 1123 424 1124 428
rect 1127 427 1128 431
rect 1132 430 1133 431
rect 1156 430 1158 436
rect 1132 428 1158 430
rect 1183 431 1189 432
rect 1174 428 1180 429
rect 1132 427 1133 428
rect 1127 426 1133 427
rect 1118 423 1124 424
rect 1174 424 1175 428
rect 1179 424 1180 428
rect 1183 427 1184 431
rect 1188 430 1189 431
rect 1216 430 1218 436
rect 1188 428 1218 430
rect 1446 431 1452 432
rect 1238 428 1244 429
rect 1302 428 1308 429
rect 1366 428 1372 429
rect 1188 427 1189 428
rect 1183 426 1189 427
rect 1174 423 1180 424
rect 1238 424 1239 428
rect 1243 424 1244 428
rect 1238 423 1244 424
rect 1247 427 1253 428
rect 1247 423 1248 427
rect 1252 426 1253 427
rect 1258 427 1264 428
rect 1258 426 1259 427
rect 1252 424 1259 426
rect 1252 423 1253 424
rect 986 422 992 423
rect 1247 422 1253 423
rect 1258 423 1259 424
rect 1263 423 1264 427
rect 1302 424 1303 428
rect 1307 424 1308 428
rect 1311 427 1317 428
rect 1311 424 1312 427
rect 1302 423 1308 424
rect 1310 423 1312 424
rect 1316 423 1317 427
rect 1366 424 1367 428
rect 1371 424 1372 428
rect 1366 423 1372 424
rect 1414 428 1420 429
rect 1414 424 1415 428
rect 1419 424 1420 428
rect 1414 423 1420 424
rect 1423 427 1432 428
rect 1423 423 1424 427
rect 1431 423 1432 427
rect 1446 427 1447 431
rect 1451 427 1452 431
rect 1446 426 1452 427
rect 1258 422 1264 423
rect 1310 419 1311 423
rect 1315 422 1317 423
rect 1423 422 1432 423
rect 1315 419 1316 422
rect 1310 418 1316 419
rect 134 416 140 417
rect 110 413 116 414
rect 110 409 111 413
rect 115 409 116 413
rect 134 412 135 416
rect 139 412 140 416
rect 134 411 140 412
rect 158 416 164 417
rect 158 412 159 416
rect 163 412 164 416
rect 158 411 164 412
rect 182 416 188 417
rect 182 412 183 416
rect 187 412 188 416
rect 182 411 188 412
rect 214 416 220 417
rect 214 412 215 416
rect 219 412 220 416
rect 214 411 220 412
rect 270 416 276 417
rect 270 412 271 416
rect 275 412 276 416
rect 270 411 276 412
rect 326 416 332 417
rect 326 412 327 416
rect 331 412 332 416
rect 326 411 332 412
rect 390 416 396 417
rect 390 412 391 416
rect 395 412 396 416
rect 390 411 396 412
rect 446 416 452 417
rect 446 412 447 416
rect 451 412 452 416
rect 446 411 452 412
rect 502 416 508 417
rect 502 412 503 416
rect 507 412 508 416
rect 502 411 508 412
rect 550 416 556 417
rect 550 412 551 416
rect 555 412 556 416
rect 550 411 556 412
rect 598 416 604 417
rect 598 412 599 416
rect 603 412 604 416
rect 598 411 604 412
rect 646 416 652 417
rect 646 412 647 416
rect 651 412 652 416
rect 646 411 652 412
rect 702 416 708 417
rect 702 412 703 416
rect 707 412 708 416
rect 702 411 708 412
rect 766 416 772 417
rect 766 412 767 416
rect 771 412 772 416
rect 766 411 772 412
rect 830 416 836 417
rect 830 412 831 416
rect 835 412 836 416
rect 830 411 836 412
rect 902 416 908 417
rect 902 412 903 416
rect 907 412 908 416
rect 902 411 908 412
rect 974 416 980 417
rect 974 412 975 416
rect 979 412 980 416
rect 974 411 980 412
rect 1038 416 1044 417
rect 1038 412 1039 416
rect 1043 412 1044 416
rect 1038 411 1044 412
rect 1102 416 1108 417
rect 1102 412 1103 416
rect 1107 412 1108 416
rect 1102 411 1108 412
rect 1158 416 1164 417
rect 1158 412 1159 416
rect 1163 412 1164 416
rect 1158 411 1164 412
rect 1206 416 1212 417
rect 1206 412 1207 416
rect 1211 412 1212 416
rect 1206 411 1212 412
rect 1246 416 1252 417
rect 1246 412 1247 416
rect 1251 412 1252 416
rect 1246 411 1252 412
rect 1278 416 1284 417
rect 1278 412 1279 416
rect 1283 412 1284 416
rect 1278 411 1284 412
rect 1318 416 1324 417
rect 1358 416 1364 417
rect 1318 412 1319 416
rect 1323 412 1324 416
rect 1318 411 1324 412
rect 1327 415 1336 416
rect 1327 411 1328 415
rect 1335 411 1336 415
rect 1358 412 1359 416
rect 1363 412 1364 416
rect 1358 411 1364 412
rect 1390 416 1396 417
rect 1390 412 1391 416
rect 1395 412 1396 416
rect 1390 411 1396 412
rect 1414 416 1420 417
rect 1414 412 1415 416
rect 1419 412 1420 416
rect 1414 411 1420 412
rect 1446 413 1452 414
rect 1327 410 1336 411
rect 110 408 116 409
rect 1446 409 1447 413
rect 1451 409 1452 413
rect 1446 408 1452 409
rect 143 407 149 408
rect 143 403 144 407
rect 148 406 149 407
rect 279 407 285 408
rect 148 404 267 406
rect 148 403 149 404
rect 143 402 149 403
rect 167 399 173 400
rect 167 398 168 399
rect 152 396 168 398
rect 110 395 116 396
rect 110 391 111 395
rect 115 391 116 395
rect 143 391 149 392
rect 110 390 116 391
rect 134 390 140 391
rect 134 386 135 390
rect 139 386 140 390
rect 143 387 144 391
rect 148 390 149 391
rect 152 390 154 396
rect 167 395 168 396
rect 172 395 173 399
rect 191 399 197 400
rect 191 398 192 399
rect 167 394 173 395
rect 176 396 192 398
rect 167 391 173 392
rect 148 388 154 390
rect 158 390 164 391
rect 148 387 149 388
rect 143 386 149 387
rect 158 386 159 390
rect 163 386 164 390
rect 167 387 168 391
rect 172 390 173 391
rect 176 390 178 396
rect 191 395 192 396
rect 196 395 197 399
rect 223 399 229 400
rect 223 398 224 399
rect 191 394 197 395
rect 209 396 224 398
rect 191 391 197 392
rect 172 388 178 390
rect 182 390 188 391
rect 172 387 173 388
rect 167 386 173 387
rect 182 386 183 390
rect 187 386 188 390
rect 191 387 192 391
rect 196 390 197 391
rect 209 390 211 396
rect 223 395 224 396
rect 228 395 229 399
rect 265 398 267 404
rect 279 403 280 407
rect 284 406 285 407
rect 338 407 344 408
rect 338 406 339 407
rect 284 404 339 406
rect 284 403 285 404
rect 279 402 285 403
rect 338 403 339 404
rect 343 403 344 407
rect 338 402 344 403
rect 346 407 352 408
rect 346 403 347 407
rect 351 406 352 407
rect 399 407 405 408
rect 399 406 400 407
rect 351 404 400 406
rect 351 403 352 404
rect 346 402 352 403
rect 399 403 400 404
rect 404 403 405 407
rect 399 402 405 403
rect 455 407 461 408
rect 455 403 456 407
rect 460 406 461 407
rect 618 407 624 408
rect 618 406 619 407
rect 460 404 619 406
rect 460 403 461 404
rect 455 402 461 403
rect 618 403 619 404
rect 623 403 624 407
rect 618 402 624 403
rect 983 407 989 408
rect 983 403 984 407
rect 988 406 989 407
rect 1050 407 1056 408
rect 1050 406 1051 407
rect 988 404 1051 406
rect 988 403 989 404
rect 983 402 989 403
rect 1050 403 1051 404
rect 1055 403 1056 407
rect 1050 402 1056 403
rect 1111 407 1117 408
rect 1111 403 1112 407
rect 1116 406 1117 407
rect 1238 407 1244 408
rect 1238 406 1239 407
rect 1116 404 1239 406
rect 1116 403 1117 404
rect 1111 402 1117 403
rect 1238 403 1239 404
rect 1243 403 1244 407
rect 1238 402 1244 403
rect 335 399 341 400
rect 265 396 283 398
rect 223 394 229 395
rect 281 392 283 396
rect 335 395 336 399
rect 340 398 341 399
rect 511 399 517 400
rect 511 398 512 399
rect 340 396 370 398
rect 340 395 341 396
rect 335 394 341 395
rect 279 391 285 392
rect 335 391 344 392
rect 196 388 211 390
rect 214 390 220 391
rect 196 387 197 388
rect 191 386 197 387
rect 214 386 215 390
rect 219 386 220 390
rect 270 390 276 391
rect 134 385 140 386
rect 158 385 164 386
rect 182 385 188 386
rect 214 385 220 386
rect 223 387 229 388
rect 126 383 132 384
rect 126 379 127 383
rect 131 382 132 383
rect 223 383 224 387
rect 228 383 229 387
rect 270 386 271 390
rect 275 386 276 390
rect 279 387 280 391
rect 284 387 285 391
rect 279 386 285 387
rect 326 390 332 391
rect 326 386 327 390
rect 331 386 332 390
rect 335 387 336 391
rect 343 387 344 391
rect 335 386 344 387
rect 270 385 276 386
rect 326 385 332 386
rect 223 382 229 383
rect 368 382 370 396
rect 484 396 512 398
rect 455 391 461 392
rect 390 390 396 391
rect 390 386 391 390
rect 395 386 396 390
rect 446 390 452 391
rect 390 385 396 386
rect 399 387 405 388
rect 399 383 400 387
rect 404 383 405 387
rect 446 386 447 390
rect 451 386 452 390
rect 455 387 456 391
rect 460 390 461 391
rect 484 390 486 396
rect 511 395 512 396
rect 516 395 517 399
rect 559 399 565 400
rect 559 398 560 399
rect 511 394 517 395
rect 536 396 560 398
rect 511 391 517 392
rect 460 388 486 390
rect 502 390 508 391
rect 460 387 461 388
rect 455 386 461 387
rect 502 386 503 390
rect 507 386 508 390
rect 511 387 512 391
rect 516 390 517 391
rect 536 390 538 396
rect 559 395 560 396
rect 564 395 565 399
rect 607 399 613 400
rect 607 398 608 399
rect 559 394 565 395
rect 584 396 608 398
rect 559 391 565 392
rect 516 388 538 390
rect 550 390 556 391
rect 516 387 517 388
rect 511 386 517 387
rect 550 386 551 390
rect 555 386 556 390
rect 559 387 560 391
rect 564 390 565 391
rect 584 390 586 396
rect 607 395 608 396
rect 612 395 613 399
rect 655 399 661 400
rect 655 398 656 399
rect 607 394 613 395
rect 632 396 656 398
rect 607 391 613 392
rect 564 388 586 390
rect 598 390 604 391
rect 564 387 565 388
rect 559 386 565 387
rect 598 386 599 390
rect 603 386 604 390
rect 607 387 608 391
rect 612 390 613 391
rect 632 390 634 396
rect 655 395 656 396
rect 660 395 661 399
rect 711 399 717 400
rect 711 398 712 399
rect 655 394 661 395
rect 679 396 712 398
rect 655 391 661 392
rect 612 388 634 390
rect 646 390 652 391
rect 612 387 613 388
rect 607 386 613 387
rect 646 386 647 390
rect 651 386 652 390
rect 655 387 656 391
rect 660 390 661 391
rect 679 390 681 396
rect 711 395 712 396
rect 716 395 717 399
rect 711 394 717 395
rect 738 399 744 400
rect 738 395 739 399
rect 743 398 744 399
rect 775 399 781 400
rect 775 398 776 399
rect 743 396 776 398
rect 743 395 744 396
rect 738 394 744 395
rect 775 395 776 396
rect 780 395 781 399
rect 839 399 845 400
rect 839 398 840 399
rect 775 394 781 395
rect 808 396 840 398
rect 775 391 781 392
rect 660 388 681 390
rect 702 390 708 391
rect 660 387 661 388
rect 655 386 661 387
rect 702 386 703 390
rect 707 386 708 390
rect 766 390 772 391
rect 446 385 452 386
rect 502 385 508 386
rect 550 385 556 386
rect 598 385 604 386
rect 646 385 652 386
rect 702 385 708 386
rect 711 387 720 388
rect 399 382 405 383
rect 711 383 712 387
rect 719 383 720 387
rect 766 386 767 390
rect 771 386 772 390
rect 775 387 776 391
rect 780 390 781 391
rect 808 390 810 396
rect 839 395 840 396
rect 844 395 845 399
rect 911 399 917 400
rect 911 398 912 399
rect 839 394 845 395
rect 876 396 912 398
rect 839 391 845 392
rect 780 388 810 390
rect 830 390 836 391
rect 780 387 781 388
rect 775 386 781 387
rect 830 386 831 390
rect 835 386 836 390
rect 839 387 840 391
rect 844 390 845 391
rect 876 390 878 396
rect 911 395 912 396
rect 916 395 917 399
rect 911 394 917 395
rect 1022 399 1028 400
rect 1022 395 1023 399
rect 1027 398 1028 399
rect 1047 399 1053 400
rect 1047 398 1048 399
rect 1027 396 1048 398
rect 1027 395 1028 396
rect 1022 394 1028 395
rect 1047 395 1048 396
rect 1052 395 1053 399
rect 1167 399 1173 400
rect 1167 398 1168 399
rect 1047 394 1053 395
rect 1140 396 1168 398
rect 983 391 992 392
rect 1047 391 1056 392
rect 1111 391 1117 392
rect 844 388 878 390
rect 902 390 908 391
rect 844 387 845 388
rect 839 386 845 387
rect 902 386 903 390
rect 907 386 908 390
rect 974 390 980 391
rect 766 385 772 386
rect 830 385 836 386
rect 902 385 908 386
rect 911 387 917 388
rect 711 382 720 383
rect 743 383 749 384
rect 131 380 227 382
rect 368 380 403 382
rect 131 379 132 380
rect 126 378 132 379
rect 346 379 352 380
rect 346 378 347 379
rect 145 376 347 378
rect 145 372 147 376
rect 346 375 347 376
rect 351 375 352 379
rect 346 374 352 375
rect 666 379 672 380
rect 666 375 667 379
rect 671 378 672 379
rect 727 379 733 380
rect 727 378 728 379
rect 671 376 728 378
rect 671 375 672 376
rect 666 374 672 375
rect 727 375 728 376
rect 732 375 733 379
rect 743 379 744 383
rect 748 382 749 383
rect 911 383 912 387
rect 916 383 917 387
rect 974 386 975 390
rect 979 386 980 390
rect 983 387 984 391
rect 991 387 992 391
rect 983 386 992 387
rect 1038 390 1044 391
rect 1038 386 1039 390
rect 1043 386 1044 390
rect 1047 387 1048 391
rect 1055 387 1056 391
rect 1047 386 1056 387
rect 1102 390 1108 391
rect 1102 386 1103 390
rect 1107 386 1108 390
rect 1111 387 1112 391
rect 1116 390 1117 391
rect 1140 390 1142 396
rect 1167 395 1168 396
rect 1172 395 1173 399
rect 1215 399 1221 400
rect 1215 398 1216 399
rect 1167 394 1173 395
rect 1176 396 1216 398
rect 1167 391 1173 392
rect 1116 388 1142 390
rect 1158 390 1164 391
rect 1116 387 1117 388
rect 1111 386 1117 387
rect 1158 386 1159 390
rect 1163 386 1164 390
rect 1167 387 1168 391
rect 1172 390 1173 391
rect 1176 390 1178 396
rect 1215 395 1216 396
rect 1220 395 1221 399
rect 1255 399 1261 400
rect 1255 398 1256 399
rect 1215 394 1221 395
rect 1236 396 1256 398
rect 1215 391 1221 392
rect 1172 388 1178 390
rect 1206 390 1212 391
rect 1172 387 1173 388
rect 1167 386 1173 387
rect 1206 386 1207 390
rect 1211 386 1212 390
rect 1215 387 1216 391
rect 1220 390 1221 391
rect 1236 390 1238 396
rect 1255 395 1256 396
rect 1260 395 1261 399
rect 1287 399 1293 400
rect 1287 398 1288 399
rect 1255 394 1261 395
rect 1272 396 1288 398
rect 1255 391 1261 392
rect 1220 388 1238 390
rect 1246 390 1252 391
rect 1220 387 1221 388
rect 1215 386 1221 387
rect 1246 386 1247 390
rect 1251 386 1252 390
rect 1255 387 1256 391
rect 1260 390 1261 391
rect 1272 390 1274 396
rect 1287 395 1288 396
rect 1292 395 1293 399
rect 1367 399 1373 400
rect 1367 398 1368 399
rect 1287 394 1293 395
rect 1348 396 1368 398
rect 1287 391 1293 392
rect 1260 388 1274 390
rect 1278 390 1284 391
rect 1260 387 1261 388
rect 1255 386 1261 387
rect 1278 386 1279 390
rect 1283 386 1284 390
rect 1287 387 1288 391
rect 1292 390 1293 391
rect 1310 391 1316 392
rect 1327 391 1333 392
rect 1310 390 1311 391
rect 1292 388 1311 390
rect 1292 387 1293 388
rect 1287 386 1293 387
rect 1310 387 1311 388
rect 1315 387 1316 391
rect 1310 386 1316 387
rect 1318 390 1324 391
rect 1318 386 1319 390
rect 1323 386 1324 390
rect 1327 387 1328 391
rect 1332 390 1333 391
rect 1348 390 1350 396
rect 1367 395 1368 396
rect 1372 395 1373 399
rect 1399 399 1405 400
rect 1399 398 1400 399
rect 1367 394 1373 395
rect 1384 396 1400 398
rect 1367 391 1373 392
rect 1332 388 1350 390
rect 1358 390 1364 391
rect 1332 387 1333 388
rect 1327 386 1333 387
rect 1358 386 1359 390
rect 1363 386 1364 390
rect 1367 387 1368 391
rect 1372 390 1373 391
rect 1384 390 1386 396
rect 1399 395 1400 396
rect 1404 395 1405 399
rect 1399 394 1405 395
rect 1423 399 1429 400
rect 1423 395 1424 399
rect 1428 398 1429 399
rect 1431 399 1437 400
rect 1431 398 1432 399
rect 1428 396 1432 398
rect 1428 395 1429 396
rect 1423 394 1429 395
rect 1431 395 1432 396
rect 1436 395 1437 399
rect 1431 394 1437 395
rect 1446 395 1452 396
rect 1423 391 1432 392
rect 1372 388 1386 390
rect 1390 390 1396 391
rect 1372 387 1373 388
rect 1367 386 1373 387
rect 1390 386 1391 390
rect 1395 386 1396 390
rect 1414 390 1420 391
rect 974 385 980 386
rect 1038 385 1044 386
rect 1102 385 1108 386
rect 1158 385 1164 386
rect 1206 385 1212 386
rect 1246 385 1252 386
rect 1278 385 1284 386
rect 1318 385 1324 386
rect 1358 385 1364 386
rect 1390 385 1396 386
rect 1399 387 1405 388
rect 911 382 917 383
rect 1023 383 1029 384
rect 748 380 915 382
rect 748 379 749 380
rect 743 378 749 379
rect 1023 379 1024 383
rect 1028 382 1029 383
rect 1258 383 1264 384
rect 1258 382 1259 383
rect 1028 380 1259 382
rect 1028 379 1029 380
rect 1023 378 1029 379
rect 1258 379 1259 380
rect 1263 379 1264 383
rect 1258 378 1264 379
rect 1382 383 1388 384
rect 1382 379 1383 383
rect 1387 382 1388 383
rect 1399 383 1400 387
rect 1404 383 1405 387
rect 1414 386 1415 390
rect 1419 386 1420 390
rect 1423 387 1424 391
rect 1431 387 1432 391
rect 1446 391 1447 395
rect 1451 391 1452 395
rect 1446 390 1452 391
rect 1423 386 1432 387
rect 1414 385 1420 386
rect 1399 382 1405 383
rect 1387 380 1403 382
rect 1387 379 1388 380
rect 1382 378 1388 379
rect 727 374 733 375
rect 1238 375 1244 376
rect 143 371 149 372
rect 735 371 744 372
rect 1238 371 1239 375
rect 1243 372 1244 375
rect 1243 371 1245 372
rect 1423 371 1429 372
rect 134 370 140 371
rect 134 366 135 370
rect 139 366 140 370
rect 143 367 144 371
rect 148 367 149 371
rect 143 366 149 367
rect 158 370 164 371
rect 158 366 159 370
rect 163 366 164 370
rect 182 370 188 371
rect 110 365 116 366
rect 134 365 140 366
rect 158 365 164 366
rect 167 367 173 368
rect 110 361 111 365
rect 115 361 116 365
rect 167 363 168 367
rect 172 363 173 367
rect 182 366 183 370
rect 187 366 188 370
rect 206 370 212 371
rect 182 365 188 366
rect 191 367 197 368
rect 167 362 173 363
rect 191 363 192 367
rect 196 363 197 367
rect 206 366 207 370
rect 211 366 212 370
rect 230 370 236 371
rect 206 365 212 366
rect 215 367 221 368
rect 191 362 197 363
rect 215 363 216 367
rect 220 363 221 367
rect 230 366 231 370
rect 235 366 236 370
rect 254 370 260 371
rect 230 365 236 366
rect 239 367 245 368
rect 215 362 221 363
rect 239 363 240 367
rect 244 363 245 367
rect 254 366 255 370
rect 259 366 260 370
rect 294 370 300 371
rect 254 365 260 366
rect 263 367 269 368
rect 239 362 245 363
rect 263 363 264 367
rect 268 363 269 367
rect 294 366 295 370
rect 299 366 300 370
rect 334 370 340 371
rect 294 365 300 366
rect 303 367 309 368
rect 263 362 269 363
rect 303 363 304 367
rect 308 363 309 367
rect 334 366 335 370
rect 339 366 340 370
rect 374 370 380 371
rect 334 365 340 366
rect 343 367 349 368
rect 303 362 309 363
rect 343 363 344 367
rect 348 363 349 367
rect 374 366 375 370
rect 379 366 380 370
rect 414 370 420 371
rect 374 365 380 366
rect 383 367 389 368
rect 343 362 349 363
rect 383 363 384 367
rect 388 366 389 367
rect 414 366 415 370
rect 419 366 420 370
rect 454 370 460 371
rect 388 364 406 366
rect 414 365 420 366
rect 423 367 429 368
rect 388 363 389 364
rect 383 362 389 363
rect 110 360 116 361
rect 143 359 149 360
rect 143 355 144 359
rect 148 358 149 359
rect 169 358 171 362
rect 148 356 171 358
rect 148 355 149 356
rect 143 354 149 355
rect 193 354 195 362
rect 217 354 219 362
rect 241 354 243 362
rect 265 354 267 362
rect 305 354 307 362
rect 345 354 347 362
rect 404 358 406 364
rect 423 363 424 367
rect 428 366 429 367
rect 454 366 455 370
rect 459 366 460 370
rect 494 370 500 371
rect 428 364 451 366
rect 454 365 460 366
rect 463 367 469 368
rect 428 363 429 364
rect 423 362 429 363
rect 423 359 429 360
rect 423 358 424 359
rect 404 356 424 358
rect 423 355 424 356
rect 428 355 429 359
rect 449 358 451 364
rect 463 363 464 367
rect 468 366 469 367
rect 494 366 495 370
rect 499 366 500 370
rect 534 370 540 371
rect 468 364 486 366
rect 494 365 500 366
rect 503 367 509 368
rect 468 363 469 364
rect 463 362 469 363
rect 463 359 469 360
rect 463 358 464 359
rect 449 356 464 358
rect 423 354 429 355
rect 463 355 464 356
rect 468 355 469 359
rect 484 358 486 364
rect 503 363 504 367
rect 508 366 509 367
rect 534 366 535 370
rect 539 366 540 370
rect 574 370 580 371
rect 508 364 526 366
rect 534 365 540 366
rect 543 367 549 368
rect 508 363 509 364
rect 503 362 509 363
rect 503 359 509 360
rect 503 358 504 359
rect 484 356 504 358
rect 463 354 469 355
rect 503 355 504 356
rect 508 355 509 359
rect 503 354 509 355
rect 524 354 526 364
rect 543 363 544 367
rect 548 363 549 367
rect 574 366 575 370
rect 579 366 580 370
rect 614 370 620 371
rect 574 365 580 366
rect 583 367 589 368
rect 543 362 549 363
rect 583 363 584 367
rect 588 366 589 367
rect 614 366 615 370
rect 619 366 620 370
rect 654 370 660 371
rect 588 364 606 366
rect 614 365 620 366
rect 623 367 632 368
rect 588 363 589 364
rect 583 362 589 363
rect 545 358 547 362
rect 583 359 589 360
rect 583 358 584 359
rect 545 356 584 358
rect 583 355 584 356
rect 588 355 589 359
rect 604 358 606 364
rect 623 363 624 367
rect 631 363 632 367
rect 654 366 655 370
rect 659 366 660 370
rect 686 370 692 371
rect 654 365 660 366
rect 663 367 669 368
rect 623 362 632 363
rect 663 363 664 367
rect 668 366 669 367
rect 686 366 687 370
rect 691 366 692 370
rect 726 370 732 371
rect 668 364 681 366
rect 686 365 692 366
rect 695 367 701 368
rect 668 363 669 364
rect 663 362 669 363
rect 623 359 629 360
rect 623 358 624 359
rect 604 356 624 358
rect 583 354 589 355
rect 623 355 624 356
rect 628 355 629 359
rect 623 354 629 355
rect 663 359 672 360
rect 663 355 664 359
rect 671 355 672 359
rect 679 358 681 364
rect 695 363 696 367
rect 700 366 701 367
rect 726 366 727 370
rect 731 366 732 370
rect 735 367 736 371
rect 743 367 744 371
rect 735 366 744 367
rect 774 370 780 371
rect 774 366 775 370
rect 779 366 780 370
rect 830 370 836 371
rect 700 364 722 366
rect 726 365 732 366
rect 774 365 780 366
rect 783 367 789 368
rect 700 363 701 364
rect 695 362 701 363
rect 695 359 701 360
rect 695 358 696 359
rect 679 356 696 358
rect 663 354 672 355
rect 695 355 696 356
rect 700 355 701 359
rect 720 358 722 364
rect 783 363 784 367
rect 788 366 789 367
rect 830 366 831 370
rect 835 366 836 370
rect 886 370 892 371
rect 788 364 814 366
rect 830 365 836 366
rect 839 367 845 368
rect 788 363 789 364
rect 783 362 789 363
rect 783 359 789 360
rect 783 358 784 359
rect 720 356 784 358
rect 695 354 701 355
rect 783 355 784 356
rect 788 355 789 359
rect 783 354 789 355
rect 812 354 814 364
rect 839 363 840 367
rect 844 363 845 367
rect 886 366 887 370
rect 891 366 892 370
rect 950 370 956 371
rect 886 365 892 366
rect 895 367 901 368
rect 839 362 845 363
rect 895 363 896 367
rect 900 366 901 367
rect 950 366 951 370
rect 955 366 956 370
rect 1014 370 1020 371
rect 900 364 930 366
rect 950 365 956 366
rect 959 367 965 368
rect 900 363 901 364
rect 895 362 901 363
rect 841 358 843 362
rect 895 359 901 360
rect 895 358 896 359
rect 841 356 896 358
rect 895 355 896 356
rect 900 355 901 359
rect 928 358 930 364
rect 959 363 960 367
rect 964 366 965 367
rect 1014 366 1015 370
rect 1019 366 1020 370
rect 1078 370 1084 371
rect 964 364 994 366
rect 1014 365 1020 366
rect 1023 367 1032 368
rect 964 363 965 364
rect 959 362 965 363
rect 959 359 965 360
rect 959 358 960 359
rect 928 356 960 358
rect 895 354 901 355
rect 959 355 960 356
rect 964 355 965 359
rect 992 358 994 364
rect 1023 363 1024 367
rect 1031 363 1032 367
rect 1078 366 1079 370
rect 1083 366 1084 370
rect 1134 370 1140 371
rect 1078 365 1084 366
rect 1087 367 1093 368
rect 1023 362 1032 363
rect 1087 363 1088 367
rect 1092 366 1093 367
rect 1134 366 1135 370
rect 1139 366 1140 370
rect 1182 370 1188 371
rect 1092 364 1118 366
rect 1134 365 1140 366
rect 1143 367 1149 368
rect 1092 363 1093 364
rect 1087 362 1093 363
rect 1023 359 1029 360
rect 1023 358 1024 359
rect 992 356 1024 358
rect 959 354 965 355
rect 1023 355 1024 356
rect 1028 355 1029 359
rect 1023 354 1029 355
rect 1116 354 1118 364
rect 1143 363 1144 367
rect 1148 363 1149 367
rect 1182 366 1183 370
rect 1187 366 1188 370
rect 1230 370 1236 371
rect 1238 370 1240 371
rect 1182 365 1188 366
rect 1191 367 1197 368
rect 1143 362 1149 363
rect 1191 363 1192 367
rect 1196 366 1197 367
rect 1230 366 1231 370
rect 1235 366 1236 370
rect 1239 367 1240 370
rect 1244 367 1245 371
rect 1239 366 1245 367
rect 1270 370 1276 371
rect 1270 366 1271 370
rect 1275 366 1276 370
rect 1310 370 1316 371
rect 1196 364 1218 366
rect 1230 365 1236 366
rect 1270 365 1276 366
rect 1279 367 1285 368
rect 1196 363 1197 364
rect 1191 362 1197 363
rect 1145 358 1147 362
rect 1191 359 1197 360
rect 1191 358 1192 359
rect 1145 356 1192 358
rect 1191 355 1192 356
rect 1196 355 1197 359
rect 1216 358 1218 364
rect 1279 363 1280 367
rect 1284 366 1285 367
rect 1290 367 1296 368
rect 1290 366 1291 367
rect 1284 364 1291 366
rect 1284 363 1285 364
rect 1279 362 1285 363
rect 1290 363 1291 364
rect 1295 363 1296 367
rect 1310 366 1311 370
rect 1315 366 1316 370
rect 1350 370 1356 371
rect 1310 365 1316 366
rect 1319 367 1325 368
rect 1290 362 1296 363
rect 1319 363 1320 367
rect 1324 363 1325 367
rect 1350 366 1351 370
rect 1355 366 1356 370
rect 1390 370 1396 371
rect 1350 365 1356 366
rect 1359 367 1365 368
rect 1319 362 1325 363
rect 1359 363 1360 367
rect 1364 363 1365 367
rect 1390 366 1391 370
rect 1395 366 1396 370
rect 1414 370 1420 371
rect 1390 365 1396 366
rect 1399 367 1405 368
rect 1359 362 1365 363
rect 1399 363 1400 367
rect 1404 363 1405 367
rect 1414 366 1415 370
rect 1419 366 1420 370
rect 1423 367 1424 371
rect 1428 370 1429 371
rect 1431 371 1437 372
rect 1431 370 1432 371
rect 1428 368 1432 370
rect 1428 367 1429 368
rect 1423 366 1429 367
rect 1431 367 1432 368
rect 1436 367 1437 371
rect 1431 366 1437 367
rect 1414 365 1420 366
rect 1446 365 1452 366
rect 1399 362 1405 363
rect 1239 359 1245 360
rect 1239 358 1240 359
rect 1216 356 1240 358
rect 1191 354 1197 355
rect 1239 355 1240 356
rect 1244 355 1245 359
rect 1239 354 1245 355
rect 1279 359 1285 360
rect 1279 355 1280 359
rect 1284 358 1285 359
rect 1321 358 1323 362
rect 1361 358 1363 362
rect 1284 356 1323 358
rect 1340 356 1363 358
rect 1401 358 1403 362
rect 1446 361 1447 365
rect 1451 361 1452 365
rect 1446 360 1452 361
rect 1423 359 1429 360
rect 1423 358 1424 359
rect 1401 356 1424 358
rect 1284 355 1285 356
rect 1279 354 1285 355
rect 169 352 195 354
rect 204 352 219 354
rect 228 352 243 354
rect 252 352 267 354
rect 284 352 307 354
rect 324 352 347 354
rect 524 352 547 354
rect 716 352 738 354
rect 812 352 843 354
rect 1116 352 1147 354
rect 167 351 173 352
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 167 347 168 351
rect 172 347 173 351
rect 204 350 206 352
rect 228 350 230 352
rect 252 350 254 352
rect 193 348 206 350
rect 217 348 230 350
rect 241 348 254 350
rect 167 346 173 347
rect 191 347 197 348
rect 110 342 116 343
rect 134 344 140 345
rect 134 340 135 344
rect 139 340 140 344
rect 134 339 140 340
rect 158 344 164 345
rect 158 340 159 344
rect 163 340 164 344
rect 158 339 164 340
rect 182 344 188 345
rect 182 340 183 344
rect 187 340 188 344
rect 191 343 192 347
rect 196 343 197 347
rect 215 347 221 348
rect 191 342 197 343
rect 206 344 212 345
rect 182 339 188 340
rect 206 340 207 344
rect 211 340 212 344
rect 215 343 216 347
rect 220 343 221 347
rect 239 347 245 348
rect 215 342 221 343
rect 230 344 236 345
rect 206 339 212 340
rect 230 340 231 344
rect 235 340 236 344
rect 239 343 240 347
rect 244 343 245 347
rect 263 347 269 348
rect 239 342 245 343
rect 254 344 260 345
rect 230 339 236 340
rect 254 340 255 344
rect 259 340 260 344
rect 263 343 264 347
rect 268 346 269 347
rect 284 346 286 352
rect 268 344 286 346
rect 303 347 309 348
rect 294 344 300 345
rect 268 343 269 344
rect 263 342 269 343
rect 254 339 260 340
rect 294 340 295 344
rect 299 340 300 344
rect 303 343 304 347
rect 308 346 309 347
rect 324 346 326 352
rect 543 351 549 352
rect 543 347 544 351
rect 548 347 549 351
rect 543 346 549 347
rect 714 351 720 352
rect 714 347 715 351
rect 719 347 720 351
rect 714 346 720 347
rect 735 351 741 352
rect 735 347 736 351
rect 740 347 741 351
rect 735 346 741 347
rect 839 351 845 352
rect 839 347 840 351
rect 844 347 845 351
rect 839 346 845 347
rect 1143 351 1149 352
rect 1143 347 1144 351
rect 1148 347 1149 351
rect 1143 346 1149 347
rect 1319 351 1325 352
rect 1319 347 1320 351
rect 1324 350 1325 351
rect 1340 350 1342 356
rect 1423 355 1424 356
rect 1428 355 1429 359
rect 1423 354 1429 355
rect 1324 348 1342 350
rect 1359 351 1365 352
rect 1324 347 1325 348
rect 1319 346 1325 347
rect 1359 347 1360 351
rect 1364 350 1365 351
rect 1382 351 1388 352
rect 1382 350 1383 351
rect 1364 348 1383 350
rect 1364 347 1365 348
rect 1359 346 1365 347
rect 1382 347 1383 348
rect 1387 347 1388 351
rect 1382 346 1388 347
rect 1446 347 1452 348
rect 308 344 326 346
rect 334 344 340 345
rect 374 344 380 345
rect 414 344 420 345
rect 308 343 309 344
rect 303 342 309 343
rect 294 339 300 340
rect 334 340 335 344
rect 339 340 340 344
rect 334 339 340 340
rect 343 343 352 344
rect 343 339 344 343
rect 351 339 352 343
rect 374 340 375 344
rect 379 340 380 344
rect 374 339 380 340
rect 383 343 389 344
rect 383 339 384 343
rect 388 342 389 343
rect 406 343 412 344
rect 406 342 407 343
rect 388 340 407 342
rect 388 339 389 340
rect 343 338 352 339
rect 383 338 389 339
rect 406 339 407 340
rect 411 339 412 343
rect 414 340 415 344
rect 419 340 420 344
rect 414 339 420 340
rect 454 344 460 345
rect 454 340 455 344
rect 459 340 460 344
rect 454 339 460 340
rect 494 344 500 345
rect 494 340 495 344
rect 499 340 500 344
rect 494 339 500 340
rect 534 344 540 345
rect 534 340 535 344
rect 539 340 540 344
rect 534 339 540 340
rect 574 344 580 345
rect 574 340 575 344
rect 579 340 580 344
rect 574 339 580 340
rect 614 344 620 345
rect 614 340 615 344
rect 619 340 620 344
rect 614 339 620 340
rect 654 344 660 345
rect 654 340 655 344
rect 659 340 660 344
rect 654 339 660 340
rect 686 344 692 345
rect 686 340 687 344
rect 691 340 692 344
rect 686 339 692 340
rect 726 344 732 345
rect 726 340 727 344
rect 731 340 732 344
rect 726 339 732 340
rect 774 344 780 345
rect 774 340 775 344
rect 779 340 780 344
rect 774 339 780 340
rect 830 344 836 345
rect 830 340 831 344
rect 835 340 836 344
rect 830 339 836 340
rect 886 344 892 345
rect 886 340 887 344
rect 891 340 892 344
rect 886 339 892 340
rect 950 344 956 345
rect 950 340 951 344
rect 955 340 956 344
rect 950 339 956 340
rect 1014 344 1020 345
rect 1014 340 1015 344
rect 1019 340 1020 344
rect 1014 339 1020 340
rect 1078 344 1084 345
rect 1134 344 1140 345
rect 1078 340 1079 344
rect 1083 340 1084 344
rect 1078 339 1084 340
rect 1087 343 1093 344
rect 1087 339 1088 343
rect 1092 342 1093 343
rect 1119 343 1125 344
rect 1119 342 1120 343
rect 1092 340 1120 342
rect 1092 339 1093 340
rect 406 338 412 339
rect 1087 338 1093 339
rect 1119 339 1120 340
rect 1124 339 1125 343
rect 1134 340 1135 344
rect 1139 340 1140 344
rect 1134 339 1140 340
rect 1182 344 1188 345
rect 1182 340 1183 344
rect 1187 340 1188 344
rect 1182 339 1188 340
rect 1230 344 1236 345
rect 1230 340 1231 344
rect 1235 340 1236 344
rect 1230 339 1236 340
rect 1270 344 1276 345
rect 1270 340 1271 344
rect 1275 340 1276 344
rect 1270 339 1276 340
rect 1310 344 1316 345
rect 1310 340 1311 344
rect 1315 340 1316 344
rect 1310 339 1316 340
rect 1350 344 1356 345
rect 1350 340 1351 344
rect 1355 340 1356 344
rect 1350 339 1356 340
rect 1390 344 1396 345
rect 1414 344 1420 345
rect 1390 340 1391 344
rect 1395 340 1396 344
rect 1390 339 1396 340
rect 1399 343 1408 344
rect 1399 339 1400 343
rect 1407 339 1408 343
rect 1414 340 1415 344
rect 1419 340 1420 344
rect 1446 343 1447 347
rect 1451 343 1452 347
rect 1446 342 1452 343
rect 1414 339 1420 340
rect 1119 338 1125 339
rect 1399 338 1408 339
rect 265 336 290 338
rect 263 335 269 336
rect 174 332 180 333
rect 110 329 116 330
rect 110 325 111 329
rect 115 325 116 329
rect 174 328 175 332
rect 179 328 180 332
rect 174 327 180 328
rect 198 332 204 333
rect 198 328 199 332
rect 203 328 204 332
rect 198 327 204 328
rect 222 332 228 333
rect 222 328 223 332
rect 227 328 228 332
rect 222 327 228 328
rect 246 332 252 333
rect 246 328 247 332
rect 251 328 252 332
rect 263 331 264 335
rect 268 331 269 335
rect 288 334 290 336
rect 304 336 330 338
rect 304 334 306 336
rect 263 330 269 331
rect 278 332 284 333
rect 288 332 306 334
rect 318 332 324 333
rect 246 327 252 328
rect 278 328 279 332
rect 283 328 284 332
rect 278 327 284 328
rect 318 328 319 332
rect 323 328 324 332
rect 328 330 330 336
rect 358 332 364 333
rect 328 328 342 330
rect 318 327 324 328
rect 110 324 116 325
rect 183 323 189 324
rect 183 319 184 323
rect 188 322 189 323
rect 210 323 216 324
rect 210 322 211 323
rect 188 320 211 322
rect 188 319 189 320
rect 183 318 189 319
rect 210 319 211 320
rect 215 319 216 323
rect 210 318 216 319
rect 231 323 237 324
rect 231 319 232 323
rect 236 322 237 323
rect 258 323 264 324
rect 258 322 259 323
rect 236 320 259 322
rect 236 319 237 320
rect 231 318 237 319
rect 258 319 259 320
rect 263 319 264 323
rect 258 318 264 319
rect 287 323 293 324
rect 287 319 288 323
rect 292 322 293 323
rect 330 323 336 324
rect 330 322 331 323
rect 292 320 331 322
rect 292 319 293 320
rect 287 318 293 319
rect 330 319 331 320
rect 335 319 336 323
rect 340 322 342 328
rect 358 328 359 332
rect 363 328 364 332
rect 358 327 364 328
rect 398 332 404 333
rect 398 328 399 332
rect 403 328 404 332
rect 398 327 404 328
rect 438 332 444 333
rect 438 328 439 332
rect 443 328 444 332
rect 438 327 444 328
rect 478 332 484 333
rect 478 328 479 332
rect 483 328 484 332
rect 478 327 484 328
rect 526 332 532 333
rect 526 328 527 332
rect 531 328 532 332
rect 526 327 532 328
rect 582 332 588 333
rect 582 328 583 332
rect 587 328 588 332
rect 582 327 588 328
rect 638 332 644 333
rect 638 328 639 332
rect 643 328 644 332
rect 638 327 644 328
rect 686 332 692 333
rect 686 328 687 332
rect 691 328 692 332
rect 686 327 692 328
rect 734 332 740 333
rect 734 328 735 332
rect 739 328 740 332
rect 734 327 740 328
rect 790 332 796 333
rect 790 328 791 332
rect 795 328 796 332
rect 790 327 796 328
rect 846 332 852 333
rect 846 328 847 332
rect 851 328 852 332
rect 846 327 852 328
rect 894 332 900 333
rect 894 328 895 332
rect 899 328 900 332
rect 894 327 900 328
rect 942 332 948 333
rect 942 328 943 332
rect 947 328 948 332
rect 942 327 948 328
rect 990 332 996 333
rect 990 328 991 332
rect 995 328 996 332
rect 990 327 996 328
rect 1038 332 1044 333
rect 1038 328 1039 332
rect 1043 328 1044 332
rect 1038 327 1044 328
rect 1086 332 1092 333
rect 1086 328 1087 332
rect 1091 328 1092 332
rect 1086 327 1092 328
rect 1134 332 1140 333
rect 1134 328 1135 332
rect 1139 328 1140 332
rect 1134 327 1140 328
rect 1182 332 1188 333
rect 1182 328 1183 332
rect 1187 328 1188 332
rect 1182 327 1188 328
rect 1230 332 1236 333
rect 1230 328 1231 332
rect 1235 328 1236 332
rect 1230 327 1236 328
rect 1278 332 1284 333
rect 1326 332 1332 333
rect 1278 328 1279 332
rect 1283 328 1284 332
rect 1278 327 1284 328
rect 1287 331 1296 332
rect 1287 327 1288 331
rect 1295 327 1296 331
rect 1326 328 1327 332
rect 1331 328 1332 332
rect 1326 327 1332 328
rect 1382 332 1388 333
rect 1382 328 1383 332
rect 1387 328 1388 332
rect 1382 327 1388 328
rect 1414 332 1420 333
rect 1414 328 1415 332
rect 1419 328 1420 332
rect 1414 327 1420 328
rect 1446 329 1452 330
rect 1287 326 1296 327
rect 1446 325 1447 329
rect 1451 325 1452 329
rect 1446 324 1452 325
rect 367 323 373 324
rect 367 322 368 323
rect 340 320 368 322
rect 330 318 336 319
rect 367 319 368 320
rect 372 319 373 323
rect 367 318 373 319
rect 407 323 413 324
rect 407 319 408 323
rect 412 322 413 323
rect 450 323 456 324
rect 450 322 451 323
rect 412 320 451 322
rect 412 319 413 320
rect 407 318 413 319
rect 450 319 451 320
rect 455 319 456 323
rect 450 318 456 319
rect 535 323 541 324
rect 535 319 536 323
rect 540 322 541 323
rect 626 323 632 324
rect 626 322 627 323
rect 540 320 627 322
rect 540 319 541 320
rect 535 318 541 319
rect 626 319 627 320
rect 631 319 632 323
rect 626 318 632 319
rect 743 323 749 324
rect 743 319 744 323
rect 748 322 749 323
rect 1026 323 1032 324
rect 1026 322 1027 323
rect 748 320 1027 322
rect 748 319 749 320
rect 743 318 749 319
rect 1026 319 1027 320
rect 1031 319 1032 323
rect 1026 318 1032 319
rect 1047 323 1053 324
rect 1047 319 1048 323
rect 1052 322 1053 323
rect 1258 323 1264 324
rect 1258 322 1259 323
rect 1052 320 1259 322
rect 1052 319 1053 320
rect 1047 318 1053 319
rect 1258 319 1259 320
rect 1263 319 1264 323
rect 1258 318 1264 319
rect 207 315 213 316
rect 110 311 116 312
rect 110 307 111 311
rect 115 307 116 311
rect 207 311 208 315
rect 212 314 213 315
rect 215 315 221 316
rect 215 314 216 315
rect 212 312 216 314
rect 212 311 213 312
rect 207 310 213 311
rect 215 311 216 312
rect 220 311 221 315
rect 215 310 221 311
rect 255 315 261 316
rect 255 311 256 315
rect 260 314 261 315
rect 327 315 333 316
rect 260 312 290 314
rect 260 311 261 312
rect 255 310 261 311
rect 288 308 290 312
rect 327 311 328 315
rect 332 314 333 315
rect 447 315 453 316
rect 332 312 350 314
rect 332 311 333 312
rect 327 310 333 311
rect 183 307 189 308
rect 207 307 216 308
rect 255 307 264 308
rect 287 307 293 308
rect 327 307 336 308
rect 110 306 116 307
rect 174 306 180 307
rect 174 302 175 306
rect 179 302 180 306
rect 183 303 184 307
rect 188 303 189 307
rect 183 302 189 303
rect 198 306 204 307
rect 198 302 199 306
rect 203 302 204 306
rect 207 303 208 307
rect 215 303 216 307
rect 207 302 216 303
rect 222 306 228 307
rect 222 302 223 306
rect 227 302 228 306
rect 246 306 252 307
rect 174 301 180 302
rect 198 301 204 302
rect 222 301 228 302
rect 231 303 237 304
rect 231 299 232 303
rect 236 299 237 303
rect 246 302 247 306
rect 251 302 252 306
rect 255 303 256 307
rect 263 303 264 307
rect 255 302 264 303
rect 278 306 284 307
rect 278 302 279 306
rect 283 302 284 306
rect 287 303 288 307
rect 292 303 293 307
rect 287 302 293 303
rect 318 306 324 307
rect 318 302 319 306
rect 323 302 324 306
rect 327 303 328 307
rect 335 303 336 307
rect 327 302 336 303
rect 246 301 252 302
rect 278 301 284 302
rect 318 301 324 302
rect 231 298 237 299
rect 263 299 269 300
rect 215 295 221 296
rect 215 291 216 295
rect 220 294 221 295
rect 233 294 235 298
rect 263 295 264 299
rect 268 295 269 299
rect 348 298 350 312
rect 447 311 448 315
rect 452 314 453 315
rect 487 315 493 316
rect 452 312 470 314
rect 452 311 453 312
rect 447 310 453 311
rect 407 307 416 308
rect 447 307 456 308
rect 358 306 364 307
rect 358 302 359 306
rect 363 302 364 306
rect 398 306 404 307
rect 358 301 364 302
rect 367 303 373 304
rect 367 299 368 303
rect 372 299 373 303
rect 398 302 399 306
rect 403 302 404 306
rect 407 303 408 307
rect 415 303 416 307
rect 407 302 416 303
rect 438 306 444 307
rect 438 302 439 306
rect 443 302 444 306
rect 447 303 448 307
rect 455 303 456 307
rect 447 302 456 303
rect 398 301 404 302
rect 438 301 444 302
rect 367 298 373 299
rect 468 298 470 312
rect 487 311 488 315
rect 492 314 493 315
rect 518 315 524 316
rect 518 314 519 315
rect 492 312 519 314
rect 492 311 493 312
rect 487 310 493 311
rect 518 311 519 312
rect 523 311 524 315
rect 591 315 597 316
rect 591 314 592 315
rect 518 310 524 311
rect 564 312 592 314
rect 535 307 541 308
rect 478 306 484 307
rect 478 302 479 306
rect 483 302 484 306
rect 526 306 532 307
rect 478 301 484 302
rect 487 303 493 304
rect 487 299 488 303
rect 492 299 493 303
rect 526 302 527 306
rect 531 302 532 306
rect 535 303 536 307
rect 540 306 541 307
rect 564 306 566 312
rect 591 311 592 312
rect 596 311 597 315
rect 647 315 653 316
rect 647 314 648 315
rect 591 310 597 311
rect 620 312 648 314
rect 591 307 597 308
rect 540 304 566 306
rect 582 306 588 307
rect 540 303 541 304
rect 535 302 541 303
rect 582 302 583 306
rect 587 302 588 306
rect 591 303 592 307
rect 596 306 597 307
rect 620 306 622 312
rect 647 311 648 312
rect 652 311 653 315
rect 695 315 701 316
rect 695 314 696 315
rect 647 310 653 311
rect 679 312 696 314
rect 647 307 653 308
rect 596 304 622 306
rect 638 306 644 307
rect 596 303 597 304
rect 591 302 597 303
rect 638 302 639 306
rect 643 302 644 306
rect 647 303 648 307
rect 652 306 653 307
rect 679 306 681 312
rect 695 311 696 312
rect 700 311 701 315
rect 799 315 805 316
rect 799 314 800 315
rect 695 310 701 311
rect 772 312 800 314
rect 743 307 749 308
rect 652 304 681 306
rect 686 306 692 307
rect 652 303 653 304
rect 647 302 653 303
rect 686 302 687 306
rect 691 302 692 306
rect 734 306 740 307
rect 526 301 532 302
rect 582 301 588 302
rect 638 301 644 302
rect 686 301 692 302
rect 695 303 701 304
rect 487 298 493 299
rect 570 299 576 300
rect 348 296 371 298
rect 468 296 491 298
rect 263 294 269 295
rect 518 295 524 296
rect 220 292 235 294
rect 220 291 221 292
rect 255 291 261 292
rect 215 290 221 291
rect 246 290 252 291
rect 246 286 247 290
rect 251 286 252 290
rect 255 287 256 291
rect 260 290 261 291
rect 265 290 267 294
rect 518 291 519 295
rect 523 292 524 295
rect 570 295 571 299
rect 575 298 576 299
rect 695 299 696 303
rect 700 299 701 303
rect 734 302 735 306
rect 739 302 740 306
rect 743 303 744 307
rect 748 306 749 307
rect 772 306 774 312
rect 799 311 800 312
rect 804 311 805 315
rect 855 315 861 316
rect 855 314 856 315
rect 799 310 805 311
rect 828 312 856 314
rect 799 307 805 308
rect 748 304 774 306
rect 790 306 796 307
rect 748 303 749 304
rect 743 302 749 303
rect 790 302 791 306
rect 795 302 796 306
rect 799 303 800 307
rect 804 306 805 307
rect 828 306 830 312
rect 855 311 856 312
rect 860 311 861 315
rect 903 315 909 316
rect 903 314 904 315
rect 855 310 861 311
rect 880 312 904 314
rect 855 307 861 308
rect 804 304 830 306
rect 846 306 852 307
rect 804 303 805 304
rect 799 302 805 303
rect 846 302 847 306
rect 851 302 852 306
rect 855 303 856 307
rect 860 306 861 307
rect 880 306 882 312
rect 903 311 904 312
rect 908 311 909 315
rect 951 315 957 316
rect 951 314 952 315
rect 903 310 909 311
rect 928 312 952 314
rect 903 307 909 308
rect 860 304 882 306
rect 894 306 900 307
rect 860 303 861 304
rect 855 302 861 303
rect 894 302 895 306
rect 899 302 900 306
rect 903 303 904 307
rect 908 306 909 307
rect 928 306 930 312
rect 951 311 952 312
rect 956 311 957 315
rect 999 315 1005 316
rect 999 314 1000 315
rect 951 310 957 311
rect 977 312 1000 314
rect 951 307 957 308
rect 908 304 930 306
rect 942 306 948 307
rect 908 303 909 304
rect 903 302 909 303
rect 942 302 943 306
rect 947 302 948 306
rect 951 303 952 307
rect 956 306 957 307
rect 977 306 979 312
rect 999 311 1000 312
rect 1004 311 1005 315
rect 1095 315 1101 316
rect 1095 314 1096 315
rect 999 310 1005 311
rect 1072 312 1096 314
rect 1047 307 1053 308
rect 956 304 979 306
rect 990 306 996 307
rect 956 303 957 304
rect 951 302 957 303
rect 990 302 991 306
rect 995 302 996 306
rect 1038 306 1044 307
rect 734 301 740 302
rect 790 301 796 302
rect 846 301 852 302
rect 894 301 900 302
rect 942 301 948 302
rect 990 301 996 302
rect 999 303 1005 304
rect 695 298 701 299
rect 770 299 776 300
rect 575 296 699 298
rect 575 295 576 296
rect 570 294 576 295
rect 770 295 771 299
rect 775 298 776 299
rect 999 299 1000 303
rect 1004 299 1005 303
rect 1038 302 1039 306
rect 1043 302 1044 306
rect 1047 303 1048 307
rect 1052 306 1053 307
rect 1072 306 1074 312
rect 1095 311 1096 312
rect 1100 311 1101 315
rect 1143 315 1149 316
rect 1143 314 1144 315
rect 1095 310 1101 311
rect 1120 312 1144 314
rect 1095 307 1101 308
rect 1052 304 1074 306
rect 1086 306 1092 307
rect 1052 303 1053 304
rect 1047 302 1053 303
rect 1086 302 1087 306
rect 1091 302 1092 306
rect 1095 303 1096 307
rect 1100 306 1101 307
rect 1120 306 1122 312
rect 1143 311 1144 312
rect 1148 311 1149 315
rect 1191 315 1197 316
rect 1191 314 1192 315
rect 1143 310 1149 311
rect 1168 312 1192 314
rect 1143 307 1149 308
rect 1100 304 1122 306
rect 1134 306 1140 307
rect 1100 303 1101 304
rect 1095 302 1101 303
rect 1134 302 1135 306
rect 1139 302 1140 306
rect 1143 303 1144 307
rect 1148 306 1149 307
rect 1168 306 1170 312
rect 1191 311 1192 312
rect 1196 311 1197 315
rect 1239 315 1245 316
rect 1239 314 1240 315
rect 1191 310 1197 311
rect 1216 312 1240 314
rect 1191 307 1197 308
rect 1148 304 1170 306
rect 1182 306 1188 307
rect 1148 303 1149 304
rect 1143 302 1149 303
rect 1182 302 1183 306
rect 1187 302 1188 306
rect 1191 303 1192 307
rect 1196 306 1197 307
rect 1216 306 1218 312
rect 1239 311 1240 312
rect 1244 311 1245 315
rect 1335 315 1341 316
rect 1335 314 1336 315
rect 1239 310 1245 311
rect 1289 312 1336 314
rect 1289 308 1291 312
rect 1335 311 1336 312
rect 1340 311 1341 315
rect 1335 310 1341 311
rect 1391 315 1397 316
rect 1391 311 1392 315
rect 1396 314 1397 315
rect 1399 315 1405 316
rect 1399 314 1400 315
rect 1396 312 1400 314
rect 1396 311 1397 312
rect 1391 310 1397 311
rect 1399 311 1400 312
rect 1404 311 1405 315
rect 1399 310 1405 311
rect 1423 315 1432 316
rect 1423 311 1424 315
rect 1431 311 1432 315
rect 1423 310 1432 311
rect 1446 311 1452 312
rect 1287 307 1293 308
rect 1391 307 1397 308
rect 1196 304 1218 306
rect 1230 306 1236 307
rect 1196 303 1197 304
rect 1191 302 1197 303
rect 1230 302 1231 306
rect 1235 302 1236 306
rect 1278 306 1284 307
rect 1038 301 1044 302
rect 1086 301 1092 302
rect 1134 301 1140 302
rect 1182 301 1188 302
rect 1230 301 1236 302
rect 1239 303 1245 304
rect 999 298 1005 299
rect 1119 299 1125 300
rect 775 296 1003 298
rect 775 295 776 296
rect 770 294 776 295
rect 1119 295 1120 299
rect 1124 298 1125 299
rect 1239 299 1240 303
rect 1244 299 1245 303
rect 1278 302 1279 306
rect 1283 302 1284 306
rect 1287 303 1288 307
rect 1292 303 1293 307
rect 1287 302 1293 303
rect 1326 306 1332 307
rect 1326 302 1327 306
rect 1331 302 1332 306
rect 1382 306 1388 307
rect 1278 301 1284 302
rect 1326 301 1332 302
rect 1335 303 1341 304
rect 1239 298 1245 299
rect 1335 299 1336 303
rect 1340 302 1341 303
rect 1374 303 1380 304
rect 1374 302 1375 303
rect 1340 300 1375 302
rect 1340 299 1341 300
rect 1335 298 1341 299
rect 1374 299 1375 300
rect 1379 299 1380 303
rect 1382 302 1383 306
rect 1387 302 1388 306
rect 1391 303 1392 307
rect 1396 306 1397 307
rect 1402 307 1408 308
rect 1446 307 1447 311
rect 1451 307 1452 311
rect 1402 306 1403 307
rect 1396 304 1403 306
rect 1396 303 1397 304
rect 1391 302 1397 303
rect 1402 303 1403 304
rect 1407 303 1408 307
rect 1402 302 1408 303
rect 1414 306 1420 307
rect 1446 306 1452 307
rect 1414 302 1415 306
rect 1419 302 1420 306
rect 1382 301 1388 302
rect 1414 301 1420 302
rect 1423 303 1429 304
rect 1374 298 1380 299
rect 1399 299 1405 300
rect 1124 296 1243 298
rect 1124 295 1125 296
rect 1119 294 1125 295
rect 1399 295 1400 299
rect 1404 298 1405 299
rect 1423 299 1424 303
rect 1428 299 1429 303
rect 1423 298 1429 299
rect 1404 296 1427 298
rect 1404 295 1405 296
rect 1399 294 1405 295
rect 523 291 525 292
rect 1255 291 1264 292
rect 1423 291 1432 292
rect 260 288 267 290
rect 270 290 276 291
rect 260 287 261 288
rect 255 286 261 287
rect 270 286 271 290
rect 275 286 276 290
rect 294 290 300 291
rect 110 285 116 286
rect 246 285 252 286
rect 270 285 276 286
rect 279 287 285 288
rect 110 281 111 285
rect 115 281 116 285
rect 279 283 280 287
rect 284 283 285 287
rect 294 286 295 290
rect 299 286 300 290
rect 318 290 324 291
rect 294 285 300 286
rect 303 287 312 288
rect 279 282 285 283
rect 303 283 304 287
rect 311 283 312 287
rect 318 286 319 290
rect 323 286 324 290
rect 342 290 348 291
rect 318 285 324 286
rect 327 287 333 288
rect 303 282 312 283
rect 327 283 328 287
rect 332 283 333 287
rect 342 286 343 290
rect 347 286 348 290
rect 366 290 372 291
rect 342 285 348 286
rect 351 287 357 288
rect 327 282 333 283
rect 351 283 352 287
rect 356 283 357 287
rect 366 286 367 290
rect 371 286 372 290
rect 398 290 404 291
rect 366 285 372 286
rect 375 287 381 288
rect 351 282 357 283
rect 375 283 376 287
rect 380 283 381 287
rect 398 286 399 290
rect 403 286 404 290
rect 430 290 436 291
rect 398 285 404 286
rect 407 287 413 288
rect 375 282 381 283
rect 407 283 408 287
rect 412 283 413 287
rect 430 286 431 290
rect 435 286 436 290
rect 470 290 476 291
rect 430 285 436 286
rect 439 287 445 288
rect 407 282 413 283
rect 439 283 440 287
rect 444 286 445 287
rect 470 286 471 290
rect 475 286 476 290
rect 510 290 516 291
rect 518 290 520 291
rect 444 284 462 286
rect 470 285 476 286
rect 479 287 485 288
rect 444 283 445 284
rect 439 282 445 283
rect 110 280 116 281
rect 255 279 261 280
rect 255 275 256 279
rect 260 278 261 279
rect 280 278 282 282
rect 260 276 282 278
rect 260 275 261 276
rect 255 274 261 275
rect 294 275 300 276
rect 294 274 295 275
rect 281 272 295 274
rect 279 271 285 272
rect 110 267 116 268
rect 110 263 111 267
rect 115 263 116 267
rect 279 267 280 271
rect 284 267 285 271
rect 294 271 295 272
rect 299 271 300 275
rect 294 270 300 271
rect 303 275 309 276
rect 303 271 304 275
rect 308 274 309 275
rect 329 274 331 282
rect 352 274 354 282
rect 376 274 378 282
rect 409 274 411 282
rect 460 278 462 284
rect 479 283 480 287
rect 484 286 485 287
rect 510 286 511 290
rect 515 286 516 290
rect 519 287 520 290
rect 524 287 525 291
rect 519 286 525 287
rect 558 290 564 291
rect 558 286 559 290
rect 563 286 564 290
rect 614 290 620 291
rect 484 284 502 286
rect 510 285 516 286
rect 558 285 564 286
rect 567 287 573 288
rect 484 283 485 284
rect 479 282 485 283
rect 479 279 485 280
rect 479 278 480 279
rect 460 276 480 278
rect 308 272 331 274
rect 340 272 354 274
rect 364 272 378 274
rect 392 272 411 274
rect 418 275 424 276
rect 308 271 309 272
rect 303 270 309 271
rect 340 270 342 272
rect 364 270 366 272
rect 329 268 342 270
rect 360 268 366 270
rect 279 266 285 267
rect 327 267 333 268
rect 110 262 116 263
rect 246 264 252 265
rect 246 260 247 264
rect 251 260 252 264
rect 246 259 252 260
rect 270 264 276 265
rect 270 260 271 264
rect 275 260 276 264
rect 270 259 276 260
rect 294 264 300 265
rect 294 260 295 264
rect 299 260 300 264
rect 294 259 300 260
rect 318 264 324 265
rect 318 260 319 264
rect 323 260 324 264
rect 327 263 328 267
rect 332 263 333 267
rect 351 267 357 268
rect 327 262 333 263
rect 342 264 348 265
rect 318 259 324 260
rect 342 260 343 264
rect 347 260 348 264
rect 351 263 352 267
rect 356 266 357 267
rect 360 266 362 268
rect 356 264 362 266
rect 375 267 381 268
rect 366 264 372 265
rect 356 263 357 264
rect 351 262 357 263
rect 342 259 348 260
rect 366 260 367 264
rect 371 260 372 264
rect 375 263 376 267
rect 380 266 381 267
rect 392 266 394 272
rect 418 271 419 275
rect 423 274 424 275
rect 439 275 445 276
rect 439 274 440 275
rect 423 272 440 274
rect 423 271 424 272
rect 418 270 424 271
rect 439 271 440 272
rect 444 271 445 275
rect 479 275 480 276
rect 484 275 485 279
rect 500 278 502 284
rect 567 283 568 287
rect 572 286 573 287
rect 614 286 615 290
rect 619 286 620 290
rect 662 290 668 291
rect 572 284 598 286
rect 614 285 620 286
rect 623 287 629 288
rect 572 283 573 284
rect 567 282 573 283
rect 519 279 525 280
rect 519 278 520 279
rect 500 276 520 278
rect 479 274 485 275
rect 519 275 520 276
rect 524 275 525 279
rect 519 274 525 275
rect 567 279 576 280
rect 567 275 568 279
rect 575 275 576 279
rect 596 278 598 284
rect 623 283 624 287
rect 628 286 629 287
rect 662 286 663 290
rect 667 286 668 290
rect 710 290 716 291
rect 628 284 650 286
rect 662 285 668 286
rect 671 287 677 288
rect 628 283 629 284
rect 623 282 629 283
rect 623 279 629 280
rect 623 278 624 279
rect 596 276 624 278
rect 567 274 576 275
rect 623 275 624 276
rect 628 275 629 279
rect 648 278 650 284
rect 671 283 672 287
rect 676 286 677 287
rect 710 286 711 290
rect 715 286 716 290
rect 758 290 764 291
rect 676 284 698 286
rect 710 285 716 286
rect 719 287 728 288
rect 676 283 677 284
rect 671 282 677 283
rect 671 279 677 280
rect 671 278 672 279
rect 648 276 672 278
rect 623 274 629 275
rect 671 275 672 276
rect 676 275 677 279
rect 696 278 698 284
rect 719 283 720 287
rect 727 283 728 287
rect 758 286 759 290
rect 763 286 764 290
rect 806 290 812 291
rect 758 285 764 286
rect 767 287 773 288
rect 719 282 728 283
rect 767 283 768 287
rect 772 286 773 287
rect 806 286 807 290
rect 811 286 812 290
rect 846 290 852 291
rect 772 284 794 286
rect 806 285 812 286
rect 815 287 821 288
rect 772 283 773 284
rect 767 282 773 283
rect 719 279 725 280
rect 719 278 720 279
rect 696 276 720 278
rect 671 274 677 275
rect 719 275 720 276
rect 724 275 725 279
rect 719 274 725 275
rect 767 279 776 280
rect 767 275 768 279
rect 775 275 776 279
rect 792 278 794 284
rect 815 283 816 287
rect 820 286 821 287
rect 846 286 847 290
rect 851 286 852 290
rect 878 290 884 291
rect 820 284 838 286
rect 846 285 852 286
rect 855 287 861 288
rect 820 283 821 284
rect 815 282 821 283
rect 815 279 821 280
rect 815 278 816 279
rect 792 276 816 278
rect 767 274 776 275
rect 815 275 816 276
rect 820 275 821 279
rect 815 274 821 275
rect 836 274 838 284
rect 855 283 856 287
rect 860 283 861 287
rect 878 286 879 290
rect 883 286 884 290
rect 902 290 908 291
rect 878 285 884 286
rect 887 287 893 288
rect 855 282 861 283
rect 887 283 888 287
rect 892 286 893 287
rect 902 286 903 290
rect 907 286 908 290
rect 926 290 932 291
rect 892 284 898 286
rect 902 285 908 286
rect 911 287 917 288
rect 892 283 893 284
rect 887 282 893 283
rect 857 278 859 282
rect 887 279 893 280
rect 887 278 888 279
rect 857 276 888 278
rect 887 275 888 276
rect 892 275 893 279
rect 896 278 898 284
rect 911 283 912 287
rect 916 286 917 287
rect 926 286 927 290
rect 931 286 932 290
rect 950 290 956 291
rect 916 284 922 286
rect 926 285 932 286
rect 935 287 941 288
rect 916 283 917 284
rect 911 282 917 283
rect 911 279 917 280
rect 911 278 912 279
rect 896 276 912 278
rect 887 274 893 275
rect 911 275 912 276
rect 916 275 917 279
rect 920 278 922 284
rect 935 283 936 287
rect 940 286 941 287
rect 950 286 951 290
rect 955 286 956 290
rect 974 290 980 291
rect 940 284 946 286
rect 950 285 956 286
rect 959 287 965 288
rect 940 283 941 284
rect 935 282 941 283
rect 935 279 941 280
rect 935 278 936 279
rect 920 276 936 278
rect 911 274 917 275
rect 935 275 936 276
rect 940 275 941 279
rect 944 278 946 284
rect 959 283 960 287
rect 964 286 965 287
rect 974 286 975 290
rect 979 286 980 290
rect 998 290 1004 291
rect 964 284 970 286
rect 974 285 980 286
rect 983 287 989 288
rect 964 283 965 284
rect 959 282 965 283
rect 959 279 965 280
rect 959 278 960 279
rect 944 276 960 278
rect 935 274 941 275
rect 959 275 960 276
rect 964 275 965 279
rect 968 278 970 284
rect 983 283 984 287
rect 988 286 989 287
rect 998 286 999 290
rect 1003 286 1004 290
rect 1022 290 1028 291
rect 988 284 994 286
rect 998 285 1004 286
rect 1007 287 1013 288
rect 988 283 989 284
rect 983 282 989 283
rect 983 279 989 280
rect 983 278 984 279
rect 968 276 984 278
rect 959 274 965 275
rect 983 275 984 276
rect 988 275 989 279
rect 992 278 994 284
rect 1007 283 1008 287
rect 1012 286 1013 287
rect 1022 286 1023 290
rect 1027 286 1028 290
rect 1046 290 1052 291
rect 1012 284 1018 286
rect 1022 285 1028 286
rect 1031 287 1037 288
rect 1012 283 1013 284
rect 1007 282 1013 283
rect 1007 279 1013 280
rect 1007 278 1008 279
rect 992 276 1008 278
rect 983 274 989 275
rect 1007 275 1008 276
rect 1012 275 1013 279
rect 1016 278 1018 284
rect 1031 283 1032 287
rect 1036 286 1037 287
rect 1046 286 1047 290
rect 1051 286 1052 290
rect 1070 290 1076 291
rect 1036 284 1042 286
rect 1046 285 1052 286
rect 1055 287 1061 288
rect 1036 283 1037 284
rect 1031 282 1037 283
rect 1031 279 1037 280
rect 1031 278 1032 279
rect 1016 276 1032 278
rect 1007 274 1013 275
rect 1031 275 1032 276
rect 1036 275 1037 279
rect 1040 278 1042 284
rect 1055 283 1056 287
rect 1060 286 1061 287
rect 1070 286 1071 290
rect 1075 286 1076 290
rect 1094 290 1100 291
rect 1060 284 1066 286
rect 1070 285 1076 286
rect 1079 287 1085 288
rect 1060 283 1061 284
rect 1055 282 1061 283
rect 1055 279 1061 280
rect 1055 278 1056 279
rect 1040 276 1056 278
rect 1031 274 1037 275
rect 1055 275 1056 276
rect 1060 275 1061 279
rect 1064 278 1066 284
rect 1079 283 1080 287
rect 1084 286 1085 287
rect 1094 286 1095 290
rect 1099 286 1100 290
rect 1126 290 1132 291
rect 1084 284 1090 286
rect 1094 285 1100 286
rect 1103 287 1109 288
rect 1084 283 1085 284
rect 1079 282 1085 283
rect 1079 279 1085 280
rect 1079 278 1080 279
rect 1064 276 1080 278
rect 1055 274 1061 275
rect 1079 275 1080 276
rect 1084 275 1085 279
rect 1088 278 1090 284
rect 1103 283 1104 287
rect 1108 286 1109 287
rect 1126 286 1127 290
rect 1131 286 1132 290
rect 1158 290 1164 291
rect 1108 284 1122 286
rect 1126 285 1132 286
rect 1135 287 1141 288
rect 1108 283 1109 284
rect 1103 282 1109 283
rect 1103 279 1109 280
rect 1103 278 1104 279
rect 1088 276 1104 278
rect 1079 274 1085 275
rect 1103 275 1104 276
rect 1108 275 1109 279
rect 1120 278 1122 284
rect 1135 283 1136 287
rect 1140 286 1141 287
rect 1158 286 1159 290
rect 1163 286 1164 290
rect 1198 290 1204 291
rect 1140 284 1150 286
rect 1158 285 1164 286
rect 1167 287 1173 288
rect 1140 283 1141 284
rect 1135 282 1141 283
rect 1135 279 1141 280
rect 1135 278 1136 279
rect 1120 276 1136 278
rect 1103 274 1109 275
rect 1135 275 1136 276
rect 1140 275 1141 279
rect 1148 278 1150 284
rect 1167 283 1168 287
rect 1172 286 1173 287
rect 1198 286 1199 290
rect 1203 286 1204 290
rect 1246 290 1252 291
rect 1172 284 1195 286
rect 1198 285 1204 286
rect 1207 287 1213 288
rect 1172 283 1173 284
rect 1167 282 1173 283
rect 1167 279 1173 280
rect 1167 278 1168 279
rect 1148 276 1168 278
rect 1135 274 1141 275
rect 1167 275 1168 276
rect 1172 275 1173 279
rect 1193 278 1195 284
rect 1207 283 1208 287
rect 1212 286 1213 287
rect 1246 286 1247 290
rect 1251 286 1252 290
rect 1255 287 1256 291
rect 1263 287 1264 291
rect 1255 286 1264 287
rect 1302 290 1308 291
rect 1302 286 1303 290
rect 1307 286 1308 290
rect 1366 290 1372 291
rect 1212 284 1234 286
rect 1246 285 1252 286
rect 1302 285 1308 286
rect 1311 287 1320 288
rect 1212 283 1213 284
rect 1207 282 1213 283
rect 1207 279 1213 280
rect 1207 278 1208 279
rect 1193 276 1208 278
rect 1167 274 1173 275
rect 1207 275 1208 276
rect 1212 275 1213 279
rect 1232 278 1234 284
rect 1311 283 1312 287
rect 1319 283 1320 287
rect 1366 286 1367 290
rect 1371 286 1372 290
rect 1414 290 1420 291
rect 1366 285 1372 286
rect 1375 287 1381 288
rect 1311 282 1320 283
rect 1375 283 1376 287
rect 1380 283 1381 287
rect 1414 286 1415 290
rect 1419 286 1420 290
rect 1423 287 1424 291
rect 1431 287 1432 291
rect 1423 286 1432 287
rect 1414 285 1420 286
rect 1446 285 1452 286
rect 1375 282 1381 283
rect 1255 279 1261 280
rect 1255 278 1256 279
rect 1232 276 1256 278
rect 1207 274 1213 275
rect 1255 275 1256 276
rect 1260 275 1261 279
rect 1255 274 1261 275
rect 1311 279 1317 280
rect 1311 275 1312 279
rect 1316 278 1317 279
rect 1376 278 1378 282
rect 1446 281 1447 285
rect 1451 281 1452 285
rect 1446 280 1452 281
rect 1316 276 1378 278
rect 1316 275 1317 276
rect 1311 274 1317 275
rect 1383 275 1389 276
rect 836 272 859 274
rect 439 270 445 271
rect 855 271 861 272
rect 380 264 394 266
rect 407 267 416 268
rect 398 264 404 265
rect 380 263 381 264
rect 375 262 381 263
rect 366 259 372 260
rect 398 260 399 264
rect 403 260 404 264
rect 407 263 408 267
rect 415 263 416 267
rect 855 267 856 271
rect 860 267 861 271
rect 1383 271 1384 275
rect 1388 274 1389 275
rect 1423 275 1429 276
rect 1423 274 1424 275
rect 1388 272 1424 274
rect 1388 271 1389 272
rect 1383 270 1389 271
rect 1423 271 1424 272
rect 1428 271 1429 275
rect 1423 270 1429 271
rect 855 266 861 267
rect 1375 267 1384 268
rect 407 262 416 263
rect 430 264 436 265
rect 398 259 404 260
rect 430 260 431 264
rect 435 260 436 264
rect 430 259 436 260
rect 470 264 476 265
rect 470 260 471 264
rect 475 260 476 264
rect 470 259 476 260
rect 510 264 516 265
rect 510 260 511 264
rect 515 260 516 264
rect 510 259 516 260
rect 558 264 564 265
rect 558 260 559 264
rect 563 260 564 264
rect 558 259 564 260
rect 614 264 620 265
rect 614 260 615 264
rect 619 260 620 264
rect 614 259 620 260
rect 662 264 668 265
rect 662 260 663 264
rect 667 260 668 264
rect 662 259 668 260
rect 710 264 716 265
rect 710 260 711 264
rect 715 260 716 264
rect 710 259 716 260
rect 758 264 764 265
rect 758 260 759 264
rect 763 260 764 264
rect 758 259 764 260
rect 806 264 812 265
rect 806 260 807 264
rect 811 260 812 264
rect 806 259 812 260
rect 846 264 852 265
rect 846 260 847 264
rect 851 260 852 264
rect 846 259 852 260
rect 878 264 884 265
rect 878 260 879 264
rect 883 260 884 264
rect 878 259 884 260
rect 902 264 908 265
rect 902 260 903 264
rect 907 260 908 264
rect 902 259 908 260
rect 926 264 932 265
rect 926 260 927 264
rect 931 260 932 264
rect 926 259 932 260
rect 950 264 956 265
rect 950 260 951 264
rect 955 260 956 264
rect 950 259 956 260
rect 974 264 980 265
rect 974 260 975 264
rect 979 260 980 264
rect 974 259 980 260
rect 998 264 1004 265
rect 998 260 999 264
rect 1003 260 1004 264
rect 998 259 1004 260
rect 1022 264 1028 265
rect 1022 260 1023 264
rect 1027 260 1028 264
rect 1022 259 1028 260
rect 1046 264 1052 265
rect 1046 260 1047 264
rect 1051 260 1052 264
rect 1046 259 1052 260
rect 1070 264 1076 265
rect 1070 260 1071 264
rect 1075 260 1076 264
rect 1070 259 1076 260
rect 1094 264 1100 265
rect 1094 260 1095 264
rect 1099 260 1100 264
rect 1094 259 1100 260
rect 1126 264 1132 265
rect 1126 260 1127 264
rect 1131 260 1132 264
rect 1126 259 1132 260
rect 1158 264 1164 265
rect 1158 260 1159 264
rect 1163 260 1164 264
rect 1158 259 1164 260
rect 1198 264 1204 265
rect 1198 260 1199 264
rect 1203 260 1204 264
rect 1198 259 1204 260
rect 1246 264 1252 265
rect 1246 260 1247 264
rect 1251 260 1252 264
rect 1246 259 1252 260
rect 1302 264 1308 265
rect 1302 260 1303 264
rect 1307 260 1308 264
rect 1302 259 1308 260
rect 1366 264 1372 265
rect 1366 260 1367 264
rect 1371 260 1372 264
rect 1375 263 1376 267
rect 1383 263 1384 267
rect 1446 267 1452 268
rect 1375 262 1384 263
rect 1414 264 1420 265
rect 1366 259 1372 260
rect 1414 260 1415 264
rect 1419 260 1420 264
rect 1446 263 1447 267
rect 1451 263 1452 267
rect 1446 262 1452 263
rect 1414 259 1420 260
rect 262 252 268 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 262 248 263 252
rect 267 248 268 252
rect 262 247 268 248
rect 286 252 292 253
rect 286 248 287 252
rect 291 248 292 252
rect 286 247 292 248
rect 310 252 316 253
rect 310 248 311 252
rect 315 248 316 252
rect 310 247 316 248
rect 334 252 340 253
rect 334 248 335 252
rect 339 248 340 252
rect 334 247 340 248
rect 358 252 364 253
rect 358 248 359 252
rect 363 248 364 252
rect 358 247 364 248
rect 382 252 388 253
rect 382 248 383 252
rect 387 248 388 252
rect 382 247 388 248
rect 406 252 412 253
rect 406 248 407 252
rect 411 248 412 252
rect 406 247 412 248
rect 430 252 436 253
rect 430 248 431 252
rect 435 248 436 252
rect 430 247 436 248
rect 462 252 468 253
rect 462 248 463 252
rect 467 248 468 252
rect 462 247 468 248
rect 502 252 508 253
rect 502 248 503 252
rect 507 248 508 252
rect 502 247 508 248
rect 542 252 548 253
rect 542 248 543 252
rect 547 248 548 252
rect 542 247 548 248
rect 582 252 588 253
rect 582 248 583 252
rect 587 248 588 252
rect 582 247 588 248
rect 622 252 628 253
rect 622 248 623 252
rect 627 248 628 252
rect 622 247 628 248
rect 678 252 684 253
rect 678 248 679 252
rect 683 248 684 252
rect 678 247 684 248
rect 742 252 748 253
rect 742 248 743 252
rect 747 248 748 252
rect 742 247 748 248
rect 806 252 812 253
rect 806 248 807 252
rect 811 248 812 252
rect 806 247 812 248
rect 878 252 884 253
rect 878 248 879 252
rect 883 248 884 252
rect 878 247 884 248
rect 958 252 964 253
rect 958 248 959 252
rect 963 248 964 252
rect 958 247 964 248
rect 1038 252 1044 253
rect 1038 248 1039 252
rect 1043 248 1044 252
rect 1038 247 1044 248
rect 1118 252 1124 253
rect 1118 248 1119 252
rect 1123 248 1124 252
rect 1118 247 1124 248
rect 1198 252 1204 253
rect 1198 248 1199 252
rect 1203 248 1204 252
rect 1198 247 1204 248
rect 1278 252 1284 253
rect 1358 252 1364 253
rect 1278 248 1279 252
rect 1283 248 1284 252
rect 1278 247 1284 248
rect 1287 251 1293 252
rect 1287 247 1288 251
rect 1292 250 1293 251
rect 1314 251 1320 252
rect 1314 250 1315 251
rect 1292 248 1315 250
rect 1292 247 1293 248
rect 1287 246 1293 247
rect 1314 247 1315 248
rect 1319 247 1320 251
rect 1358 248 1359 252
rect 1363 248 1364 252
rect 1358 247 1364 248
rect 1414 252 1420 253
rect 1414 248 1415 252
rect 1419 248 1420 252
rect 1414 247 1420 248
rect 1446 249 1452 250
rect 1314 246 1320 247
rect 110 244 116 245
rect 1446 245 1447 249
rect 1451 245 1452 249
rect 1446 244 1452 245
rect 295 243 301 244
rect 295 239 296 243
rect 300 242 301 243
rect 322 243 328 244
rect 322 242 323 243
rect 300 240 323 242
rect 300 239 301 240
rect 295 238 301 239
rect 322 239 323 240
rect 327 239 328 243
rect 346 243 352 244
rect 346 242 347 243
rect 322 238 328 239
rect 336 240 347 242
rect 271 235 277 236
rect 110 231 116 232
rect 110 227 111 231
rect 115 227 116 231
rect 271 231 272 235
rect 276 234 277 235
rect 319 235 325 236
rect 276 232 298 234
rect 276 231 277 232
rect 271 230 277 231
rect 296 228 298 232
rect 319 231 320 235
rect 324 234 325 235
rect 336 234 338 240
rect 346 239 347 240
rect 351 239 352 243
rect 367 243 373 244
rect 346 238 352 239
rect 358 239 364 240
rect 324 232 338 234
rect 343 235 349 236
rect 324 231 325 232
rect 319 230 325 231
rect 343 231 344 235
rect 348 234 349 235
rect 358 235 359 239
rect 363 235 364 239
rect 367 239 368 243
rect 372 242 373 243
rect 394 243 400 244
rect 394 242 395 243
rect 372 240 395 242
rect 372 239 373 240
rect 367 238 373 239
rect 394 239 395 240
rect 399 239 400 243
rect 394 238 400 239
rect 439 243 445 244
rect 439 239 440 243
rect 444 242 445 243
rect 474 243 480 244
rect 474 242 475 243
rect 444 240 475 242
rect 444 239 445 240
rect 439 238 445 239
rect 474 239 475 240
rect 479 239 480 243
rect 474 238 480 239
rect 511 243 517 244
rect 511 239 512 243
rect 516 242 517 243
rect 554 243 560 244
rect 554 242 555 243
rect 516 240 555 242
rect 516 239 517 240
rect 511 238 517 239
rect 554 239 555 240
rect 559 239 560 243
rect 631 243 637 244
rect 554 238 560 239
rect 590 239 597 240
rect 358 234 364 235
rect 391 235 397 236
rect 391 234 392 235
rect 348 232 362 234
rect 376 232 392 234
rect 348 231 349 232
rect 343 230 349 231
rect 271 227 280 228
rect 295 227 301 228
rect 319 227 328 228
rect 343 227 352 228
rect 367 227 373 228
rect 110 226 116 227
rect 262 226 268 227
rect 262 222 263 226
rect 267 222 268 226
rect 271 223 272 227
rect 279 223 280 227
rect 271 222 280 223
rect 286 226 292 227
rect 286 222 287 226
rect 291 222 292 226
rect 295 223 296 227
rect 300 223 301 227
rect 295 222 301 223
rect 310 226 316 227
rect 310 222 311 226
rect 315 222 316 226
rect 319 223 320 227
rect 327 223 328 227
rect 319 222 328 223
rect 334 226 340 227
rect 334 222 335 226
rect 339 222 340 226
rect 343 223 344 227
rect 351 223 352 227
rect 343 222 352 223
rect 358 226 364 227
rect 358 222 359 226
rect 363 222 364 226
rect 367 223 368 227
rect 372 226 373 227
rect 376 226 378 232
rect 391 231 392 232
rect 396 231 397 235
rect 415 235 421 236
rect 415 234 416 235
rect 391 230 397 231
rect 400 232 416 234
rect 391 227 397 228
rect 372 224 378 226
rect 382 226 388 227
rect 372 223 373 224
rect 367 222 373 223
rect 382 222 383 226
rect 387 222 388 226
rect 391 223 392 227
rect 396 226 397 227
rect 400 226 402 232
rect 415 231 416 232
rect 420 231 421 235
rect 415 230 421 231
rect 471 235 477 236
rect 471 231 472 235
rect 476 234 477 235
rect 551 235 557 236
rect 476 232 494 234
rect 476 231 477 232
rect 471 230 477 231
rect 415 227 424 228
rect 471 227 480 228
rect 396 224 402 226
rect 406 226 412 227
rect 396 223 397 224
rect 391 222 397 223
rect 406 222 407 226
rect 411 222 412 226
rect 415 223 416 227
rect 423 223 424 227
rect 415 222 424 223
rect 430 226 436 227
rect 430 222 431 226
rect 435 222 436 226
rect 462 226 468 227
rect 262 221 268 222
rect 286 221 292 222
rect 310 221 316 222
rect 334 221 340 222
rect 358 221 364 222
rect 382 221 388 222
rect 406 221 412 222
rect 430 221 436 222
rect 439 223 445 224
rect 366 219 372 220
rect 366 215 367 219
rect 371 218 372 219
rect 439 219 440 223
rect 444 219 445 223
rect 462 222 463 226
rect 467 222 468 226
rect 471 223 472 227
rect 479 223 480 227
rect 471 222 480 223
rect 462 221 468 222
rect 439 218 445 219
rect 492 218 494 232
rect 551 231 552 235
rect 556 234 557 235
rect 590 235 591 239
rect 596 235 597 239
rect 631 239 632 243
rect 636 242 637 243
rect 722 243 728 244
rect 722 242 723 243
rect 636 240 723 242
rect 636 239 637 240
rect 631 238 637 239
rect 722 239 723 240
rect 727 239 728 243
rect 722 238 728 239
rect 1047 243 1053 244
rect 1047 239 1048 243
rect 1052 242 1053 243
rect 1130 243 1136 244
rect 1130 242 1131 243
rect 1052 240 1131 242
rect 1052 239 1053 240
rect 1047 238 1053 239
rect 1130 239 1131 240
rect 1135 239 1136 243
rect 1130 238 1136 239
rect 590 234 597 235
rect 687 235 693 236
rect 687 234 688 235
rect 556 232 574 234
rect 556 231 557 232
rect 551 230 557 231
rect 551 227 560 228
rect 502 226 508 227
rect 502 222 503 226
rect 507 222 508 226
rect 542 226 548 227
rect 502 221 508 222
rect 511 223 517 224
rect 511 219 512 223
rect 516 219 517 223
rect 542 222 543 226
rect 547 222 548 226
rect 551 223 552 227
rect 559 223 560 227
rect 551 222 560 223
rect 542 221 548 222
rect 511 218 517 219
rect 572 218 574 232
rect 660 232 688 234
rect 631 227 637 228
rect 582 226 588 227
rect 582 222 583 226
rect 587 222 588 226
rect 622 226 628 227
rect 582 221 588 222
rect 591 223 597 224
rect 591 219 592 223
rect 596 219 597 223
rect 622 222 623 226
rect 627 222 628 226
rect 631 223 632 227
rect 636 226 637 227
rect 660 226 662 232
rect 687 231 688 232
rect 692 231 693 235
rect 751 235 757 236
rect 751 234 752 235
rect 687 230 693 231
rect 716 232 752 234
rect 687 227 693 228
rect 636 224 662 226
rect 678 226 684 227
rect 636 223 637 224
rect 631 222 637 223
rect 678 222 679 226
rect 683 222 684 226
rect 687 223 688 227
rect 692 226 693 227
rect 716 226 718 232
rect 751 231 752 232
rect 756 231 757 235
rect 815 235 821 236
rect 815 234 816 235
rect 751 230 757 231
rect 784 232 816 234
rect 751 227 757 228
rect 692 224 718 226
rect 742 226 748 227
rect 692 223 693 224
rect 687 222 693 223
rect 742 222 743 226
rect 747 222 748 226
rect 751 223 752 227
rect 756 226 757 227
rect 784 226 786 232
rect 815 231 816 232
rect 820 231 821 235
rect 887 235 893 236
rect 887 234 888 235
rect 815 230 821 231
rect 852 232 888 234
rect 815 227 821 228
rect 756 224 786 226
rect 806 226 812 227
rect 756 223 757 224
rect 751 222 757 223
rect 806 222 807 226
rect 811 222 812 226
rect 815 223 816 227
rect 820 226 821 227
rect 852 226 854 232
rect 887 231 888 232
rect 892 231 893 235
rect 967 235 973 236
rect 967 234 968 235
rect 887 230 893 231
rect 932 232 968 234
rect 887 227 893 228
rect 820 224 854 226
rect 878 226 884 227
rect 820 223 821 224
rect 815 222 821 223
rect 878 222 879 226
rect 883 222 884 226
rect 887 223 888 227
rect 892 226 893 227
rect 932 226 934 232
rect 967 231 968 232
rect 972 231 973 235
rect 967 230 973 231
rect 1127 235 1133 236
rect 1127 231 1128 235
rect 1132 234 1133 235
rect 1207 235 1213 236
rect 1132 232 1161 234
rect 1132 231 1133 232
rect 1127 230 1133 231
rect 1127 227 1136 228
rect 892 224 934 226
rect 958 226 964 227
rect 892 223 893 224
rect 887 222 893 223
rect 958 222 959 226
rect 963 222 964 226
rect 1038 226 1044 227
rect 622 221 628 222
rect 678 221 684 222
rect 742 221 748 222
rect 806 221 812 222
rect 878 221 884 222
rect 958 221 964 222
rect 967 223 973 224
rect 591 218 597 219
rect 730 219 736 220
rect 371 216 442 218
rect 492 216 514 218
rect 572 216 595 218
rect 371 215 372 216
rect 366 214 372 215
rect 730 215 731 219
rect 735 218 736 219
rect 967 219 968 223
rect 972 219 973 223
rect 1038 222 1039 226
rect 1043 222 1044 226
rect 1118 226 1124 227
rect 1038 221 1044 222
rect 1047 223 1053 224
rect 967 218 973 219
rect 1047 219 1048 223
rect 1052 222 1053 223
rect 1094 223 1100 224
rect 1094 222 1095 223
rect 1052 220 1095 222
rect 1052 219 1053 220
rect 1047 218 1053 219
rect 1094 219 1095 220
rect 1099 219 1100 223
rect 1118 222 1119 226
rect 1123 222 1124 226
rect 1127 223 1128 227
rect 1135 223 1136 227
rect 1127 222 1136 223
rect 1118 221 1124 222
rect 1094 218 1100 219
rect 1159 218 1161 232
rect 1207 231 1208 235
rect 1212 234 1213 235
rect 1367 235 1373 236
rect 1212 232 1291 234
rect 1212 231 1213 232
rect 1207 230 1213 231
rect 1289 228 1291 232
rect 1367 231 1368 235
rect 1372 234 1373 235
rect 1423 235 1432 236
rect 1372 232 1398 234
rect 1372 231 1373 232
rect 1367 230 1373 231
rect 1287 227 1293 228
rect 1367 227 1373 228
rect 1198 226 1204 227
rect 1198 222 1199 226
rect 1203 222 1204 226
rect 1278 226 1284 227
rect 1198 221 1204 222
rect 1207 223 1213 224
rect 1207 219 1208 223
rect 1212 219 1213 223
rect 1278 222 1279 226
rect 1283 222 1284 226
rect 1287 223 1288 227
rect 1292 223 1293 227
rect 1287 222 1293 223
rect 1358 226 1364 227
rect 1358 222 1359 226
rect 1363 222 1364 226
rect 1367 223 1368 227
rect 1372 226 1373 227
rect 1383 227 1389 228
rect 1383 226 1384 227
rect 1372 224 1384 226
rect 1372 223 1373 224
rect 1367 222 1373 223
rect 1383 223 1384 224
rect 1388 223 1389 227
rect 1383 222 1389 223
rect 1278 221 1284 222
rect 1358 221 1364 222
rect 1207 218 1213 219
rect 1396 218 1398 232
rect 1423 231 1424 235
rect 1431 231 1432 235
rect 1423 230 1432 231
rect 1446 231 1452 232
rect 1446 227 1447 231
rect 1451 227 1452 231
rect 1414 226 1420 227
rect 1446 226 1452 227
rect 1414 222 1415 226
rect 1419 222 1420 226
rect 1414 221 1420 222
rect 1423 223 1429 224
rect 1423 219 1424 223
rect 1428 219 1429 223
rect 1423 218 1429 219
rect 735 216 970 218
rect 1159 216 1210 218
rect 1396 216 1427 218
rect 735 215 736 216
rect 730 214 736 215
rect 391 211 400 212
rect 1423 211 1432 212
rect 238 210 244 211
rect 238 206 239 210
rect 243 206 244 210
rect 262 210 268 211
rect 110 205 116 206
rect 238 205 244 206
rect 247 207 253 208
rect 110 201 111 205
rect 115 201 116 205
rect 247 203 248 207
rect 252 206 253 207
rect 262 206 263 210
rect 267 206 268 210
rect 286 210 292 211
rect 252 204 259 206
rect 262 205 268 206
rect 271 207 277 208
rect 252 203 253 204
rect 247 202 253 203
rect 110 200 116 201
rect 257 198 259 204
rect 271 203 272 207
rect 276 206 277 207
rect 286 206 287 210
rect 291 206 292 210
rect 310 210 316 211
rect 276 204 282 206
rect 286 205 292 206
rect 295 207 301 208
rect 276 203 277 204
rect 271 202 277 203
rect 271 199 277 200
rect 271 198 272 199
rect 257 196 272 198
rect 271 195 272 196
rect 276 195 277 199
rect 280 198 282 204
rect 295 203 296 207
rect 300 206 301 207
rect 310 206 311 210
rect 315 206 316 210
rect 334 210 340 211
rect 300 204 306 206
rect 310 205 316 206
rect 319 207 325 208
rect 300 203 301 204
rect 295 202 301 203
rect 295 199 301 200
rect 295 198 296 199
rect 280 196 296 198
rect 271 194 277 195
rect 295 195 296 196
rect 300 195 301 199
rect 304 198 306 204
rect 319 203 320 207
rect 324 206 325 207
rect 334 206 335 210
rect 339 206 340 210
rect 358 210 364 211
rect 324 204 331 206
rect 334 205 340 206
rect 343 207 349 208
rect 324 203 325 204
rect 319 202 325 203
rect 319 199 325 200
rect 319 198 320 199
rect 304 196 320 198
rect 295 194 301 195
rect 319 195 320 196
rect 324 195 325 199
rect 329 198 331 204
rect 343 203 344 207
rect 348 206 349 207
rect 358 206 359 210
rect 363 206 364 210
rect 382 210 388 211
rect 348 204 354 206
rect 358 205 364 206
rect 367 207 373 208
rect 348 203 349 204
rect 343 202 349 203
rect 343 199 349 200
rect 343 198 344 199
rect 329 196 344 198
rect 319 194 325 195
rect 343 195 344 196
rect 348 195 349 199
rect 343 194 349 195
rect 352 194 354 204
rect 367 203 368 207
rect 372 203 373 207
rect 382 206 383 210
rect 387 206 388 210
rect 391 207 392 211
rect 399 207 400 211
rect 391 206 400 207
rect 406 210 412 211
rect 406 206 407 210
rect 411 206 412 210
rect 430 210 436 211
rect 382 205 388 206
rect 406 205 412 206
rect 415 207 424 208
rect 367 202 373 203
rect 415 203 416 207
rect 423 203 424 207
rect 430 206 431 210
rect 435 206 436 210
rect 462 210 468 211
rect 430 205 436 206
rect 439 207 445 208
rect 415 202 424 203
rect 439 203 440 207
rect 444 203 445 207
rect 462 206 463 210
rect 467 206 468 210
rect 510 210 516 211
rect 462 205 468 206
rect 471 207 477 208
rect 439 202 445 203
rect 471 203 472 207
rect 476 203 477 207
rect 510 206 511 210
rect 515 206 516 210
rect 558 210 564 211
rect 510 205 516 206
rect 519 207 525 208
rect 471 202 477 203
rect 519 203 520 207
rect 524 203 525 207
rect 558 206 559 210
rect 563 206 564 210
rect 614 210 620 211
rect 558 205 564 206
rect 567 207 573 208
rect 519 202 525 203
rect 567 203 568 207
rect 572 203 573 207
rect 614 206 615 210
rect 619 206 620 210
rect 670 210 676 211
rect 614 205 620 206
rect 623 207 629 208
rect 567 202 573 203
rect 623 203 624 207
rect 628 203 629 207
rect 670 206 671 210
rect 675 206 676 210
rect 718 210 724 211
rect 670 205 676 206
rect 679 207 685 208
rect 623 202 629 203
rect 679 203 680 207
rect 684 203 685 207
rect 718 206 719 210
rect 723 206 724 210
rect 766 210 772 211
rect 718 205 724 206
rect 727 207 733 208
rect 679 202 685 203
rect 727 203 728 207
rect 732 206 733 207
rect 766 206 767 210
rect 771 206 772 210
rect 814 210 820 211
rect 732 204 754 206
rect 766 205 772 206
rect 775 207 781 208
rect 732 203 733 204
rect 727 202 733 203
rect 369 198 371 202
rect 391 199 397 200
rect 391 198 392 199
rect 369 196 392 198
rect 391 195 392 196
rect 396 195 397 199
rect 391 194 397 195
rect 415 199 421 200
rect 415 195 416 199
rect 420 198 421 199
rect 440 198 442 202
rect 420 196 442 198
rect 420 195 421 196
rect 415 194 421 195
rect 472 194 474 202
rect 520 194 522 202
rect 568 194 570 202
rect 624 194 626 202
rect 679 194 681 202
rect 727 199 736 200
rect 727 195 728 199
rect 735 195 736 199
rect 752 198 754 204
rect 775 203 776 207
rect 780 206 781 207
rect 814 206 815 210
rect 819 206 820 210
rect 862 210 868 211
rect 780 204 802 206
rect 814 205 820 206
rect 823 207 829 208
rect 780 203 781 204
rect 775 202 781 203
rect 775 199 781 200
rect 775 198 776 199
rect 752 196 776 198
rect 727 194 736 195
rect 775 195 776 196
rect 780 195 781 199
rect 800 198 802 204
rect 823 203 824 207
rect 828 206 829 207
rect 862 206 863 210
rect 867 206 868 210
rect 918 210 924 211
rect 828 204 850 206
rect 862 205 868 206
rect 871 207 877 208
rect 828 203 829 204
rect 823 202 829 203
rect 823 199 829 200
rect 823 198 824 199
rect 800 196 824 198
rect 775 194 781 195
rect 823 195 824 196
rect 828 195 829 199
rect 848 198 850 204
rect 871 203 872 207
rect 876 206 877 207
rect 918 206 919 210
rect 923 206 924 210
rect 974 210 980 211
rect 876 204 902 206
rect 918 205 924 206
rect 927 207 933 208
rect 876 203 877 204
rect 871 202 877 203
rect 871 199 877 200
rect 871 198 872 199
rect 848 196 872 198
rect 823 194 829 195
rect 871 195 872 196
rect 876 195 877 199
rect 900 198 902 204
rect 927 203 928 207
rect 932 206 933 207
rect 974 206 975 210
rect 979 206 980 210
rect 1030 210 1036 211
rect 932 204 958 206
rect 974 205 980 206
rect 983 207 989 208
rect 932 203 933 204
rect 927 202 933 203
rect 927 199 933 200
rect 927 198 928 199
rect 900 196 928 198
rect 871 194 877 195
rect 927 195 928 196
rect 932 195 933 199
rect 956 198 958 204
rect 983 203 984 207
rect 988 206 989 207
rect 1030 206 1031 210
rect 1035 206 1036 210
rect 1086 210 1092 211
rect 988 204 1014 206
rect 1030 205 1036 206
rect 1039 207 1045 208
rect 988 203 989 204
rect 983 202 989 203
rect 983 199 989 200
rect 983 198 984 199
rect 956 196 984 198
rect 927 194 933 195
rect 983 195 984 196
rect 988 195 989 199
rect 1012 198 1014 204
rect 1039 203 1040 207
rect 1044 206 1045 207
rect 1071 207 1077 208
rect 1071 206 1072 207
rect 1044 204 1072 206
rect 1044 203 1045 204
rect 1039 202 1045 203
rect 1071 203 1072 204
rect 1076 203 1077 207
rect 1086 206 1087 210
rect 1091 206 1092 210
rect 1134 210 1140 211
rect 1086 205 1092 206
rect 1095 207 1101 208
rect 1071 202 1077 203
rect 1095 203 1096 207
rect 1100 206 1101 207
rect 1134 206 1135 210
rect 1139 206 1140 210
rect 1182 210 1188 211
rect 1100 204 1122 206
rect 1134 205 1140 206
rect 1143 207 1149 208
rect 1100 203 1101 204
rect 1095 202 1101 203
rect 1039 199 1045 200
rect 1039 198 1040 199
rect 1012 196 1040 198
rect 983 194 989 195
rect 1039 195 1040 196
rect 1044 195 1045 199
rect 1039 194 1045 195
rect 1094 199 1101 200
rect 1094 195 1095 199
rect 1100 195 1101 199
rect 1120 198 1122 204
rect 1143 203 1144 207
rect 1148 206 1149 207
rect 1182 206 1183 210
rect 1187 206 1188 210
rect 1230 210 1236 211
rect 1148 204 1161 206
rect 1182 205 1188 206
rect 1191 207 1200 208
rect 1148 203 1149 204
rect 1143 202 1149 203
rect 1143 199 1149 200
rect 1143 198 1144 199
rect 1120 196 1144 198
rect 1094 194 1101 195
rect 1143 195 1144 196
rect 1148 195 1149 199
rect 1159 198 1161 204
rect 1191 203 1192 207
rect 1199 203 1200 207
rect 1230 206 1231 210
rect 1235 206 1236 210
rect 1278 210 1284 211
rect 1230 205 1236 206
rect 1239 207 1245 208
rect 1191 202 1200 203
rect 1239 203 1240 207
rect 1244 203 1245 207
rect 1278 206 1279 210
rect 1283 206 1284 210
rect 1326 210 1332 211
rect 1278 205 1284 206
rect 1287 207 1293 208
rect 1239 202 1245 203
rect 1287 203 1288 207
rect 1292 203 1293 207
rect 1326 206 1327 210
rect 1331 206 1332 210
rect 1382 210 1388 211
rect 1326 205 1332 206
rect 1335 207 1341 208
rect 1287 202 1293 203
rect 1335 203 1336 207
rect 1340 206 1341 207
rect 1382 206 1383 210
rect 1387 206 1388 210
rect 1414 210 1420 211
rect 1340 204 1366 206
rect 1382 205 1388 206
rect 1391 207 1397 208
rect 1340 203 1341 204
rect 1335 202 1341 203
rect 1191 199 1197 200
rect 1191 198 1192 199
rect 1159 196 1192 198
rect 1143 194 1149 195
rect 1191 195 1192 196
rect 1196 195 1197 199
rect 1191 194 1197 195
rect 1241 194 1243 202
rect 1289 198 1291 202
rect 1335 199 1341 200
rect 1335 198 1336 199
rect 1289 196 1336 198
rect 1335 195 1336 196
rect 1340 195 1341 199
rect 1335 194 1341 195
rect 352 192 371 194
rect 456 192 474 194
rect 496 192 522 194
rect 544 192 570 194
rect 596 192 626 194
rect 652 192 681 194
rect 1241 192 1291 194
rect 367 191 373 192
rect 110 187 116 188
rect 110 183 111 187
rect 115 183 116 187
rect 367 187 368 191
rect 372 187 373 191
rect 367 186 373 187
rect 439 191 445 192
rect 439 187 440 191
rect 444 190 445 191
rect 456 190 458 192
rect 444 188 458 190
rect 444 187 445 188
rect 439 186 445 187
rect 471 187 477 188
rect 110 182 116 183
rect 238 184 244 185
rect 262 184 268 185
rect 238 180 239 184
rect 243 180 244 184
rect 238 179 244 180
rect 247 183 256 184
rect 247 179 248 183
rect 255 179 256 183
rect 262 180 263 184
rect 267 180 268 184
rect 262 179 268 180
rect 286 184 292 185
rect 286 180 287 184
rect 291 180 292 184
rect 286 179 292 180
rect 310 184 316 185
rect 310 180 311 184
rect 315 180 316 184
rect 310 179 316 180
rect 334 184 340 185
rect 334 180 335 184
rect 339 180 340 184
rect 334 179 340 180
rect 358 184 364 185
rect 358 180 359 184
rect 363 180 364 184
rect 358 179 364 180
rect 382 184 388 185
rect 382 180 383 184
rect 387 180 388 184
rect 382 179 388 180
rect 406 184 412 185
rect 406 180 407 184
rect 411 180 412 184
rect 406 179 412 180
rect 430 184 436 185
rect 430 180 431 184
rect 435 180 436 184
rect 430 179 436 180
rect 462 184 468 185
rect 462 180 463 184
rect 467 180 468 184
rect 471 183 472 187
rect 476 186 477 187
rect 496 186 498 192
rect 476 184 498 186
rect 519 187 525 188
rect 510 184 516 185
rect 476 183 477 184
rect 471 182 477 183
rect 462 179 468 180
rect 510 180 511 184
rect 515 180 516 184
rect 519 183 520 187
rect 524 186 525 187
rect 544 186 546 192
rect 524 184 546 186
rect 567 187 573 188
rect 558 184 564 185
rect 524 183 525 184
rect 519 182 525 183
rect 510 179 516 180
rect 558 180 559 184
rect 563 180 564 184
rect 567 183 568 187
rect 572 186 573 187
rect 596 186 598 192
rect 572 184 598 186
rect 623 187 629 188
rect 614 184 620 185
rect 572 183 573 184
rect 567 182 573 183
rect 558 179 564 180
rect 614 180 615 184
rect 619 180 620 184
rect 623 183 624 187
rect 628 186 629 187
rect 652 186 654 192
rect 1287 191 1293 192
rect 1287 187 1288 191
rect 1292 187 1293 191
rect 1364 190 1366 204
rect 1391 203 1392 207
rect 1396 203 1397 207
rect 1414 206 1415 210
rect 1419 206 1420 210
rect 1423 207 1424 211
rect 1431 207 1432 211
rect 1423 206 1432 207
rect 1414 205 1420 206
rect 1446 205 1452 206
rect 1391 202 1397 203
rect 1370 199 1376 200
rect 1370 195 1371 199
rect 1375 198 1376 199
rect 1393 198 1395 202
rect 1446 201 1447 205
rect 1451 201 1452 205
rect 1446 200 1452 201
rect 1375 196 1395 198
rect 1375 195 1376 196
rect 1370 194 1376 195
rect 1380 192 1395 194
rect 1380 190 1382 192
rect 1364 188 1382 190
rect 1391 191 1397 192
rect 1287 186 1293 187
rect 1391 187 1392 191
rect 1396 187 1397 191
rect 1391 186 1397 187
rect 1446 187 1452 188
rect 628 184 654 186
rect 670 184 676 185
rect 718 184 724 185
rect 628 183 629 184
rect 623 182 629 183
rect 614 179 620 180
rect 670 180 671 184
rect 675 180 676 184
rect 670 179 676 180
rect 679 183 688 184
rect 679 179 680 183
rect 687 179 688 183
rect 718 180 719 184
rect 723 180 724 184
rect 718 179 724 180
rect 766 184 772 185
rect 766 180 767 184
rect 771 180 772 184
rect 766 179 772 180
rect 814 184 820 185
rect 814 180 815 184
rect 819 180 820 184
rect 814 179 820 180
rect 862 184 868 185
rect 862 180 863 184
rect 867 180 868 184
rect 862 179 868 180
rect 918 184 924 185
rect 918 180 919 184
rect 923 180 924 184
rect 918 179 924 180
rect 974 184 980 185
rect 974 180 975 184
rect 979 180 980 184
rect 974 179 980 180
rect 1030 184 1036 185
rect 1030 180 1031 184
rect 1035 180 1036 184
rect 1030 179 1036 180
rect 1086 184 1092 185
rect 1086 180 1087 184
rect 1091 180 1092 184
rect 1086 179 1092 180
rect 1134 184 1140 185
rect 1134 180 1135 184
rect 1139 180 1140 184
rect 1134 179 1140 180
rect 1182 184 1188 185
rect 1182 180 1183 184
rect 1187 180 1188 184
rect 1182 179 1188 180
rect 1230 184 1236 185
rect 1278 184 1284 185
rect 1230 180 1231 184
rect 1235 180 1236 184
rect 1230 179 1236 180
rect 1239 183 1245 184
rect 1239 179 1240 183
rect 1244 182 1245 183
rect 1270 183 1276 184
rect 1270 182 1271 183
rect 1244 180 1271 182
rect 1244 179 1245 180
rect 247 178 256 179
rect 679 178 688 179
rect 1239 178 1245 179
rect 1270 179 1271 180
rect 1275 179 1276 183
rect 1278 180 1279 184
rect 1283 180 1284 184
rect 1278 179 1284 180
rect 1326 184 1332 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1382 184 1388 185
rect 1382 180 1383 184
rect 1387 180 1388 184
rect 1382 179 1388 180
rect 1414 184 1420 185
rect 1414 180 1415 184
rect 1419 180 1420 184
rect 1414 179 1420 180
rect 1423 183 1432 184
rect 1423 179 1424 183
rect 1431 179 1432 183
rect 1446 183 1447 187
rect 1451 183 1452 187
rect 1446 182 1452 183
rect 1270 178 1276 179
rect 1423 178 1432 179
rect 182 172 188 173
rect 110 169 116 170
rect 110 165 111 169
rect 115 165 116 169
rect 182 168 183 172
rect 187 168 188 172
rect 182 167 188 168
rect 206 172 212 173
rect 206 168 207 172
rect 211 168 212 172
rect 206 167 212 168
rect 238 172 244 173
rect 238 168 239 172
rect 243 168 244 172
rect 238 167 244 168
rect 278 172 284 173
rect 278 168 279 172
rect 283 168 284 172
rect 278 167 284 168
rect 326 172 332 173
rect 326 168 327 172
rect 331 168 332 172
rect 326 167 332 168
rect 374 172 380 173
rect 374 168 375 172
rect 379 168 380 172
rect 374 167 380 168
rect 422 172 428 173
rect 422 168 423 172
rect 427 168 428 172
rect 422 167 428 168
rect 470 172 476 173
rect 470 168 471 172
rect 475 168 476 172
rect 470 167 476 168
rect 526 172 532 173
rect 526 168 527 172
rect 531 168 532 172
rect 526 167 532 168
rect 590 172 596 173
rect 590 168 591 172
rect 595 168 596 172
rect 590 167 596 168
rect 654 172 660 173
rect 654 168 655 172
rect 659 168 660 172
rect 654 167 660 168
rect 710 172 716 173
rect 710 168 711 172
rect 715 168 716 172
rect 710 167 716 168
rect 766 172 772 173
rect 766 168 767 172
rect 771 168 772 172
rect 766 167 772 168
rect 822 172 828 173
rect 822 168 823 172
rect 827 168 828 172
rect 822 167 828 168
rect 870 172 876 173
rect 870 168 871 172
rect 875 168 876 172
rect 870 167 876 168
rect 918 172 924 173
rect 918 168 919 172
rect 923 168 924 172
rect 918 167 924 168
rect 974 172 980 173
rect 974 168 975 172
rect 979 168 980 172
rect 974 167 980 168
rect 1030 172 1036 173
rect 1030 168 1031 172
rect 1035 168 1036 172
rect 1030 167 1036 168
rect 1078 172 1084 173
rect 1078 168 1079 172
rect 1083 168 1084 172
rect 1078 167 1084 168
rect 1126 172 1132 173
rect 1126 168 1127 172
rect 1131 168 1132 172
rect 1126 167 1132 168
rect 1174 172 1180 173
rect 1174 168 1175 172
rect 1179 168 1180 172
rect 1174 167 1180 168
rect 1222 172 1228 173
rect 1222 168 1223 172
rect 1227 168 1228 172
rect 1222 167 1228 168
rect 1262 172 1268 173
rect 1262 168 1263 172
rect 1267 168 1268 172
rect 1262 167 1268 168
rect 1294 172 1300 173
rect 1294 168 1295 172
rect 1299 168 1300 172
rect 1294 167 1300 168
rect 1326 172 1332 173
rect 1326 168 1327 172
rect 1331 168 1332 172
rect 1326 167 1332 168
rect 1358 172 1364 173
rect 1390 172 1396 173
rect 1358 168 1359 172
rect 1363 168 1364 172
rect 1358 167 1364 168
rect 1367 171 1376 172
rect 1367 167 1368 171
rect 1375 167 1376 171
rect 1390 168 1391 172
rect 1395 168 1396 172
rect 1390 167 1396 168
rect 1414 172 1420 173
rect 1414 168 1415 172
rect 1419 168 1420 172
rect 1414 167 1420 168
rect 1446 169 1452 170
rect 1367 166 1376 167
rect 110 164 116 165
rect 1446 165 1447 169
rect 1451 165 1452 169
rect 1446 164 1452 165
rect 191 163 197 164
rect 191 159 192 163
rect 196 162 197 163
rect 410 163 416 164
rect 410 162 411 163
rect 196 160 411 162
rect 196 159 197 160
rect 191 158 197 159
rect 410 159 411 160
rect 415 159 416 163
rect 410 158 416 159
rect 431 163 437 164
rect 431 159 432 163
rect 436 162 437 163
rect 482 163 488 164
rect 482 162 483 163
rect 436 160 483 162
rect 436 159 437 160
rect 431 158 437 159
rect 482 159 483 160
rect 487 159 488 163
rect 482 158 488 159
rect 535 163 541 164
rect 535 159 536 163
rect 540 162 541 163
rect 602 163 608 164
rect 602 162 603 163
rect 540 160 603 162
rect 540 159 541 160
rect 535 158 541 159
rect 602 159 603 160
rect 607 159 608 163
rect 602 158 608 159
rect 663 163 669 164
rect 663 159 664 163
rect 668 162 669 163
rect 722 163 728 164
rect 722 162 723 163
rect 668 160 723 162
rect 668 159 669 160
rect 663 158 669 159
rect 722 159 723 160
rect 727 159 728 163
rect 722 158 728 159
rect 831 163 837 164
rect 831 159 832 163
rect 836 162 837 163
rect 882 163 888 164
rect 882 162 883 163
rect 836 160 883 162
rect 836 159 837 160
rect 831 158 837 159
rect 882 159 883 160
rect 887 159 888 163
rect 882 158 888 159
rect 927 163 933 164
rect 927 159 928 163
rect 932 162 933 163
rect 986 163 992 164
rect 986 162 987 163
rect 932 160 987 162
rect 932 159 933 160
rect 927 158 933 159
rect 986 159 987 160
rect 991 159 992 163
rect 986 158 992 159
rect 1039 163 1045 164
rect 1039 159 1040 163
rect 1044 162 1045 163
rect 1090 163 1096 164
rect 1090 162 1091 163
rect 1044 160 1091 162
rect 1044 159 1045 160
rect 1039 158 1045 159
rect 1090 159 1091 160
rect 1095 159 1096 163
rect 1090 158 1096 159
rect 1135 163 1141 164
rect 1135 159 1136 163
rect 1140 162 1141 163
rect 1194 163 1200 164
rect 1194 162 1195 163
rect 1140 160 1195 162
rect 1140 159 1141 160
rect 1135 158 1141 159
rect 1194 159 1195 160
rect 1199 159 1200 163
rect 1194 158 1200 159
rect 1398 159 1405 160
rect 215 155 221 156
rect 215 154 216 155
rect 200 152 216 154
rect 110 151 116 152
rect 110 147 111 151
rect 115 147 116 151
rect 191 147 197 148
rect 110 146 116 147
rect 182 146 188 147
rect 182 142 183 146
rect 187 142 188 146
rect 191 143 192 147
rect 196 146 197 147
rect 200 146 202 152
rect 215 151 216 152
rect 220 151 221 155
rect 247 155 253 156
rect 247 154 248 155
rect 215 150 221 151
rect 233 152 248 154
rect 215 147 221 148
rect 196 144 202 146
rect 206 146 212 147
rect 196 143 197 144
rect 191 142 197 143
rect 206 142 207 146
rect 211 142 212 146
rect 215 143 216 147
rect 220 146 221 147
rect 233 146 235 152
rect 247 151 248 152
rect 252 151 253 155
rect 287 155 293 156
rect 287 154 288 155
rect 247 150 253 151
rect 268 152 288 154
rect 247 147 253 148
rect 220 144 235 146
rect 238 146 244 147
rect 220 143 221 144
rect 215 142 221 143
rect 238 142 239 146
rect 243 142 244 146
rect 247 143 248 147
rect 252 146 253 147
rect 268 146 270 152
rect 287 151 288 152
rect 292 151 293 155
rect 335 155 341 156
rect 335 154 336 155
rect 287 150 293 151
rect 319 152 336 154
rect 287 147 293 148
rect 252 144 270 146
rect 278 146 284 147
rect 252 143 253 144
rect 247 142 253 143
rect 278 142 279 146
rect 283 142 284 146
rect 287 143 288 147
rect 292 146 293 147
rect 319 146 321 152
rect 335 151 336 152
rect 340 151 341 155
rect 383 155 389 156
rect 383 154 384 155
rect 335 150 341 151
rect 360 152 384 154
rect 335 147 341 148
rect 292 144 321 146
rect 326 146 332 147
rect 292 143 293 144
rect 287 142 293 143
rect 326 142 327 146
rect 331 142 332 146
rect 335 143 336 147
rect 340 146 341 147
rect 360 146 362 152
rect 383 151 384 152
rect 388 151 389 155
rect 383 150 389 151
rect 479 155 485 156
rect 479 151 480 155
rect 484 154 485 155
rect 599 155 605 156
rect 484 152 510 154
rect 484 151 485 152
rect 479 150 485 151
rect 479 147 488 148
rect 340 144 362 146
rect 374 146 380 147
rect 340 143 341 144
rect 335 142 341 143
rect 374 142 375 146
rect 379 142 380 146
rect 422 146 428 147
rect 182 141 188 142
rect 206 141 212 142
rect 238 141 244 142
rect 278 141 284 142
rect 326 141 332 142
rect 374 141 380 142
rect 383 143 389 144
rect 250 139 256 140
rect 250 135 251 139
rect 255 138 256 139
rect 383 139 384 143
rect 388 139 389 143
rect 422 142 423 146
rect 427 142 428 146
rect 470 146 476 147
rect 422 141 428 142
rect 431 143 437 144
rect 383 138 389 139
rect 431 139 432 143
rect 436 142 437 143
rect 470 142 471 146
rect 475 142 476 146
rect 479 143 480 147
rect 487 143 488 147
rect 479 142 488 143
rect 436 140 466 142
rect 470 141 476 142
rect 436 139 437 140
rect 431 138 437 139
rect 255 136 321 138
rect 255 135 256 136
rect 250 134 256 135
rect 319 134 321 136
rect 384 134 386 138
rect 319 132 386 134
rect 464 134 466 140
rect 508 138 510 152
rect 599 151 600 155
rect 604 154 605 155
rect 670 155 676 156
rect 604 152 666 154
rect 604 151 605 152
rect 599 150 605 151
rect 664 148 666 152
rect 670 151 671 155
rect 675 154 676 155
rect 719 155 725 156
rect 719 154 720 155
rect 675 152 720 154
rect 675 151 676 152
rect 670 150 676 151
rect 719 151 720 152
rect 724 151 725 155
rect 719 150 725 151
rect 775 155 781 156
rect 775 151 776 155
rect 780 154 781 155
rect 879 155 885 156
rect 780 152 834 154
rect 780 151 781 152
rect 775 150 781 151
rect 832 148 834 152
rect 879 151 880 155
rect 884 154 885 155
rect 983 155 989 156
rect 884 152 907 154
rect 884 151 885 152
rect 879 150 885 151
rect 599 147 608 148
rect 663 147 669 148
rect 719 147 728 148
rect 831 147 837 148
rect 879 147 888 148
rect 526 146 532 147
rect 526 142 527 146
rect 531 142 532 146
rect 590 146 596 147
rect 526 141 532 142
rect 535 143 541 144
rect 535 139 536 143
rect 540 139 541 143
rect 590 142 591 146
rect 595 142 596 146
rect 599 143 600 147
rect 607 143 608 147
rect 599 142 608 143
rect 654 146 660 147
rect 654 142 655 146
rect 659 142 660 146
rect 663 143 664 147
rect 668 143 669 147
rect 663 142 669 143
rect 710 146 716 147
rect 710 142 711 146
rect 715 142 716 146
rect 719 143 720 147
rect 727 143 728 147
rect 719 142 728 143
rect 766 146 772 147
rect 766 142 767 146
rect 771 142 772 146
rect 822 146 828 147
rect 590 141 596 142
rect 654 141 660 142
rect 710 141 716 142
rect 766 141 772 142
rect 775 143 781 144
rect 535 138 541 139
rect 775 139 776 143
rect 780 142 781 143
rect 822 142 823 146
rect 827 142 828 146
rect 831 143 832 147
rect 836 143 837 147
rect 831 142 837 143
rect 870 146 876 147
rect 870 142 871 146
rect 875 142 876 146
rect 879 143 880 147
rect 887 143 888 147
rect 879 142 888 143
rect 780 140 818 142
rect 822 141 828 142
rect 870 141 876 142
rect 780 139 781 140
rect 775 138 781 139
rect 508 136 539 138
rect 682 135 688 136
rect 682 134 683 135
rect 464 132 683 134
rect 682 131 683 132
rect 687 131 688 135
rect 816 134 818 140
rect 905 138 907 152
rect 983 151 984 155
rect 988 154 989 155
rect 1071 155 1077 156
rect 988 152 1042 154
rect 988 151 989 152
rect 983 150 989 151
rect 1040 148 1042 152
rect 1071 151 1072 155
rect 1076 154 1077 155
rect 1087 155 1093 156
rect 1087 154 1088 155
rect 1076 152 1088 154
rect 1076 151 1077 152
rect 1071 150 1077 151
rect 1087 151 1088 152
rect 1092 151 1093 155
rect 1087 150 1093 151
rect 1183 155 1189 156
rect 1183 151 1184 155
rect 1188 154 1189 155
rect 1199 155 1205 156
rect 1199 154 1200 155
rect 1188 152 1200 154
rect 1188 151 1189 152
rect 1183 150 1189 151
rect 1199 151 1200 152
rect 1204 151 1205 155
rect 1231 155 1237 156
rect 1231 154 1232 155
rect 1199 150 1205 151
rect 1208 152 1232 154
rect 983 147 992 148
rect 1039 147 1045 148
rect 1087 147 1096 148
rect 1183 147 1189 148
rect 918 146 924 147
rect 918 142 919 146
rect 923 142 924 146
rect 974 146 980 147
rect 918 141 924 142
rect 927 143 933 144
rect 927 139 928 143
rect 932 139 933 143
rect 974 142 975 146
rect 979 142 980 146
rect 983 143 984 147
rect 991 143 992 147
rect 983 142 992 143
rect 1030 146 1036 147
rect 1030 142 1031 146
rect 1035 142 1036 146
rect 1039 143 1040 147
rect 1044 143 1045 147
rect 1039 142 1045 143
rect 1078 146 1084 147
rect 1078 142 1079 146
rect 1083 142 1084 146
rect 1087 143 1088 147
rect 1095 143 1096 147
rect 1087 142 1096 143
rect 1126 146 1132 147
rect 1126 142 1127 146
rect 1131 142 1132 146
rect 1174 146 1180 147
rect 974 141 980 142
rect 1030 141 1036 142
rect 1078 141 1084 142
rect 1126 141 1132 142
rect 1135 143 1141 144
rect 927 138 933 139
rect 1054 139 1060 140
rect 905 136 930 138
rect 1022 135 1028 136
rect 1022 134 1023 135
rect 816 132 1023 134
rect 682 130 688 131
rect 1022 131 1023 132
rect 1027 131 1028 135
rect 1054 135 1055 139
rect 1059 138 1060 139
rect 1135 139 1136 143
rect 1140 139 1141 143
rect 1174 142 1175 146
rect 1179 142 1180 146
rect 1183 143 1184 147
rect 1188 146 1189 147
rect 1208 146 1210 152
rect 1231 151 1232 152
rect 1236 151 1237 155
rect 1271 155 1277 156
rect 1271 154 1272 155
rect 1231 150 1237 151
rect 1252 152 1272 154
rect 1231 147 1237 148
rect 1188 144 1210 146
rect 1222 146 1228 147
rect 1188 143 1189 144
rect 1183 142 1189 143
rect 1222 142 1223 146
rect 1227 142 1228 146
rect 1231 143 1232 147
rect 1236 146 1237 147
rect 1252 146 1254 152
rect 1271 151 1272 152
rect 1276 151 1277 155
rect 1303 155 1309 156
rect 1303 154 1304 155
rect 1271 150 1277 151
rect 1289 152 1304 154
rect 1271 147 1277 148
rect 1236 144 1254 146
rect 1262 146 1268 147
rect 1236 143 1237 144
rect 1231 142 1237 143
rect 1262 142 1263 146
rect 1267 142 1268 146
rect 1271 143 1272 147
rect 1276 146 1277 147
rect 1289 146 1291 152
rect 1303 151 1304 152
rect 1308 151 1309 155
rect 1303 150 1309 151
rect 1335 155 1341 156
rect 1335 151 1336 155
rect 1340 154 1341 155
rect 1398 155 1399 159
rect 1404 155 1405 159
rect 1398 154 1405 155
rect 1423 155 1429 156
rect 1423 154 1424 155
rect 1340 152 1370 154
rect 1340 151 1341 152
rect 1335 150 1341 151
rect 1368 148 1370 152
rect 1408 152 1424 154
rect 1367 147 1373 148
rect 1399 147 1405 148
rect 1276 144 1291 146
rect 1294 146 1300 147
rect 1276 143 1277 144
rect 1271 142 1277 143
rect 1294 142 1295 146
rect 1299 142 1300 146
rect 1326 146 1332 147
rect 1174 141 1180 142
rect 1222 141 1228 142
rect 1262 141 1268 142
rect 1294 141 1300 142
rect 1303 143 1309 144
rect 1135 138 1141 139
rect 1270 139 1276 140
rect 1059 136 1138 138
rect 1059 135 1060 136
rect 1054 134 1060 135
rect 1270 135 1271 139
rect 1275 138 1276 139
rect 1303 139 1304 143
rect 1308 139 1309 143
rect 1326 142 1327 146
rect 1331 142 1332 146
rect 1358 146 1364 147
rect 1326 141 1332 142
rect 1335 143 1341 144
rect 1303 138 1309 139
rect 1335 139 1336 143
rect 1340 139 1341 143
rect 1358 142 1359 146
rect 1363 142 1364 146
rect 1367 143 1368 147
rect 1372 143 1373 147
rect 1367 142 1373 143
rect 1390 146 1396 147
rect 1390 142 1391 146
rect 1395 142 1396 146
rect 1399 143 1400 147
rect 1404 146 1405 147
rect 1408 146 1410 152
rect 1423 151 1424 152
rect 1428 151 1429 155
rect 1423 150 1429 151
rect 1446 151 1452 152
rect 1423 147 1432 148
rect 1404 144 1410 146
rect 1414 146 1420 147
rect 1404 143 1405 144
rect 1399 142 1405 143
rect 1414 142 1415 146
rect 1419 142 1420 146
rect 1423 143 1424 147
rect 1431 143 1432 147
rect 1446 147 1447 151
rect 1451 147 1452 151
rect 1446 146 1452 147
rect 1423 142 1432 143
rect 1358 141 1364 142
rect 1390 141 1396 142
rect 1414 141 1420 142
rect 1335 138 1341 139
rect 1374 139 1380 140
rect 1374 138 1375 139
rect 1275 136 1306 138
rect 1337 136 1375 138
rect 1275 135 1276 136
rect 1270 134 1276 135
rect 1374 135 1375 136
rect 1379 135 1380 139
rect 1374 134 1380 135
rect 1022 130 1028 131
rect 670 127 676 128
rect 670 126 671 127
rect 456 124 671 126
rect 407 119 416 120
rect 439 119 445 120
rect 134 118 140 119
rect 134 114 135 118
rect 139 114 140 118
rect 158 118 164 119
rect 110 113 116 114
rect 134 113 140 114
rect 143 115 149 116
rect 110 109 111 113
rect 115 109 116 113
rect 143 111 144 115
rect 148 114 149 115
rect 158 114 159 118
rect 163 114 164 118
rect 182 118 188 119
rect 148 112 154 114
rect 158 113 164 114
rect 167 115 173 116
rect 148 111 149 112
rect 143 110 149 111
rect 110 108 116 109
rect 152 106 154 112
rect 167 111 168 115
rect 172 114 173 115
rect 182 114 183 118
rect 187 114 188 118
rect 206 118 212 119
rect 172 112 178 114
rect 182 113 188 114
rect 191 115 197 116
rect 172 111 173 112
rect 167 110 173 111
rect 167 107 173 108
rect 167 106 168 107
rect 152 104 168 106
rect 167 103 168 104
rect 172 103 173 107
rect 176 106 178 112
rect 191 111 192 115
rect 196 114 197 115
rect 206 114 207 118
rect 211 114 212 118
rect 230 118 236 119
rect 196 112 202 114
rect 206 113 212 114
rect 215 115 221 116
rect 196 111 197 112
rect 191 110 197 111
rect 191 107 197 108
rect 191 106 192 107
rect 176 104 192 106
rect 167 102 173 103
rect 191 103 192 104
rect 196 103 197 107
rect 191 102 197 103
rect 200 102 202 112
rect 215 111 216 115
rect 220 111 221 115
rect 230 114 231 118
rect 235 114 236 118
rect 254 118 260 119
rect 230 113 236 114
rect 239 115 248 116
rect 215 110 221 111
rect 239 111 240 115
rect 247 111 248 115
rect 254 114 255 118
rect 259 114 260 118
rect 278 118 284 119
rect 254 113 260 114
rect 263 115 269 116
rect 239 110 248 111
rect 263 111 264 115
rect 268 111 269 115
rect 278 114 279 118
rect 283 114 284 118
rect 302 118 308 119
rect 278 113 284 114
rect 287 115 293 116
rect 263 110 269 111
rect 287 111 288 115
rect 292 111 293 115
rect 302 114 303 118
rect 307 114 308 118
rect 326 118 332 119
rect 302 113 308 114
rect 311 115 317 116
rect 287 110 293 111
rect 311 111 312 115
rect 316 114 317 115
rect 326 114 327 118
rect 331 114 332 118
rect 350 118 356 119
rect 316 112 321 114
rect 326 113 332 114
rect 335 115 341 116
rect 316 111 317 112
rect 311 110 317 111
rect 217 106 219 110
rect 239 107 245 108
rect 239 106 240 107
rect 217 104 240 106
rect 239 103 240 104
rect 244 103 245 107
rect 239 102 245 103
rect 265 102 267 110
rect 289 106 291 110
rect 311 107 317 108
rect 311 106 312 107
rect 289 104 312 106
rect 311 103 312 104
rect 316 103 317 107
rect 319 106 321 112
rect 335 111 336 115
rect 340 114 341 115
rect 350 114 351 118
rect 355 114 356 118
rect 374 118 380 119
rect 340 112 346 114
rect 350 113 356 114
rect 359 115 365 116
rect 340 111 341 112
rect 335 110 341 111
rect 335 107 341 108
rect 335 106 336 107
rect 319 104 336 106
rect 311 102 317 103
rect 335 103 336 104
rect 340 103 341 107
rect 344 106 346 112
rect 359 111 360 115
rect 364 114 365 115
rect 374 114 375 118
rect 379 114 380 118
rect 398 118 404 119
rect 364 112 371 114
rect 374 113 380 114
rect 383 115 389 116
rect 364 111 365 112
rect 359 110 365 111
rect 359 107 365 108
rect 359 106 360 107
rect 344 104 360 106
rect 335 102 341 103
rect 359 103 360 104
rect 364 103 365 107
rect 369 106 371 112
rect 383 111 384 115
rect 388 114 389 115
rect 398 114 399 118
rect 403 114 404 118
rect 407 115 408 119
rect 415 115 416 119
rect 407 114 416 115
rect 430 118 436 119
rect 430 114 431 118
rect 435 114 436 118
rect 439 115 440 119
rect 444 118 445 119
rect 456 118 458 124
rect 670 123 671 124
rect 675 123 676 127
rect 670 122 676 123
rect 1199 127 1205 128
rect 1199 123 1200 127
rect 1204 126 1205 127
rect 1398 127 1404 128
rect 1204 124 1346 126
rect 1204 123 1205 124
rect 1199 122 1205 123
rect 1344 120 1346 124
rect 1398 123 1399 127
rect 1403 126 1404 127
rect 1403 124 1427 126
rect 1403 123 1404 124
rect 1398 122 1404 123
rect 1425 120 1427 124
rect 1343 119 1349 120
rect 1423 119 1429 120
rect 444 116 458 118
rect 462 118 468 119
rect 444 115 445 116
rect 439 114 445 115
rect 462 114 463 118
rect 467 114 468 118
rect 486 118 492 119
rect 388 112 394 114
rect 398 113 404 114
rect 430 113 436 114
rect 462 113 468 114
rect 471 115 480 116
rect 388 111 389 112
rect 383 110 389 111
rect 383 107 389 108
rect 383 106 384 107
rect 369 104 384 106
rect 359 102 365 103
rect 383 103 384 104
rect 388 103 389 107
rect 392 106 394 112
rect 471 111 472 115
rect 479 111 480 115
rect 486 114 487 118
rect 491 114 492 118
rect 510 118 516 119
rect 486 113 492 114
rect 495 115 501 116
rect 471 110 480 111
rect 495 111 496 115
rect 500 111 501 115
rect 510 114 511 118
rect 515 114 516 118
rect 534 118 540 119
rect 510 113 516 114
rect 519 115 525 116
rect 495 110 501 111
rect 519 111 520 115
rect 524 111 525 115
rect 534 114 535 118
rect 539 114 540 118
rect 558 118 564 119
rect 534 113 540 114
rect 543 115 549 116
rect 519 110 525 111
rect 543 111 544 115
rect 548 111 549 115
rect 558 114 559 118
rect 563 114 564 118
rect 582 118 588 119
rect 558 113 564 114
rect 567 115 573 116
rect 543 110 549 111
rect 567 111 568 115
rect 572 111 573 115
rect 582 114 583 118
rect 587 114 588 118
rect 606 118 612 119
rect 582 113 588 114
rect 591 115 597 116
rect 567 110 573 111
rect 591 111 592 115
rect 596 111 597 115
rect 606 114 607 118
rect 611 114 612 118
rect 630 118 636 119
rect 606 113 612 114
rect 615 115 621 116
rect 591 110 597 111
rect 615 111 616 115
rect 620 111 621 115
rect 630 114 631 118
rect 635 114 636 118
rect 654 118 660 119
rect 630 113 636 114
rect 639 115 645 116
rect 615 110 621 111
rect 639 111 640 115
rect 644 111 645 115
rect 654 114 655 118
rect 659 114 660 118
rect 678 118 684 119
rect 654 113 660 114
rect 663 115 669 116
rect 639 110 645 111
rect 663 111 664 115
rect 668 111 669 115
rect 678 114 679 118
rect 683 114 684 118
rect 702 118 708 119
rect 678 113 684 114
rect 687 115 693 116
rect 663 110 669 111
rect 687 111 688 115
rect 692 111 693 115
rect 702 114 703 118
rect 707 114 708 118
rect 726 118 732 119
rect 702 113 708 114
rect 711 115 717 116
rect 687 110 693 111
rect 711 111 712 115
rect 716 111 717 115
rect 726 114 727 118
rect 731 114 732 118
rect 750 118 756 119
rect 726 113 732 114
rect 735 115 741 116
rect 711 110 717 111
rect 735 111 736 115
rect 740 111 741 115
rect 750 114 751 118
rect 755 114 756 118
rect 774 118 780 119
rect 750 113 756 114
rect 759 115 765 116
rect 735 110 741 111
rect 759 111 760 115
rect 764 111 765 115
rect 774 114 775 118
rect 779 114 780 118
rect 798 118 804 119
rect 774 113 780 114
rect 783 115 789 116
rect 759 110 765 111
rect 783 111 784 115
rect 788 111 789 115
rect 798 114 799 118
rect 803 114 804 118
rect 822 118 828 119
rect 798 113 804 114
rect 807 115 813 116
rect 783 110 789 111
rect 807 111 808 115
rect 812 111 813 115
rect 822 114 823 118
rect 827 114 828 118
rect 854 118 860 119
rect 822 113 828 114
rect 831 115 837 116
rect 807 110 813 111
rect 831 111 832 115
rect 836 111 837 115
rect 854 114 855 118
rect 859 114 860 118
rect 886 118 892 119
rect 854 113 860 114
rect 863 115 869 116
rect 831 110 837 111
rect 863 111 864 115
rect 868 111 869 115
rect 886 114 887 118
rect 891 114 892 118
rect 918 118 924 119
rect 886 113 892 114
rect 895 115 901 116
rect 863 110 869 111
rect 895 111 896 115
rect 900 111 901 115
rect 918 114 919 118
rect 923 114 924 118
rect 950 118 956 119
rect 918 113 924 114
rect 927 115 933 116
rect 895 110 901 111
rect 927 111 928 115
rect 932 111 933 115
rect 950 114 951 118
rect 955 114 956 118
rect 982 118 988 119
rect 950 113 956 114
rect 959 115 965 116
rect 927 110 933 111
rect 959 111 960 115
rect 964 111 965 115
rect 982 114 983 118
rect 987 114 988 118
rect 1014 118 1020 119
rect 982 113 988 114
rect 991 115 997 116
rect 959 110 965 111
rect 991 111 992 115
rect 996 111 997 115
rect 1014 114 1015 118
rect 1019 114 1020 118
rect 1046 118 1052 119
rect 1014 113 1020 114
rect 1023 115 1029 116
rect 991 110 997 111
rect 1023 111 1024 115
rect 1028 111 1029 115
rect 1046 114 1047 118
rect 1051 114 1052 118
rect 1070 118 1076 119
rect 1046 113 1052 114
rect 1055 115 1061 116
rect 1023 110 1029 111
rect 1055 111 1056 115
rect 1060 114 1061 115
rect 1070 114 1071 118
rect 1075 114 1076 118
rect 1094 118 1100 119
rect 1060 112 1066 114
rect 1070 113 1076 114
rect 1079 115 1085 116
rect 1060 111 1061 112
rect 1055 110 1061 111
rect 407 107 413 108
rect 407 106 408 107
rect 392 104 408 106
rect 383 102 389 103
rect 407 103 408 104
rect 412 103 413 107
rect 407 102 413 103
rect 439 107 445 108
rect 439 103 440 107
rect 444 106 445 107
rect 462 107 468 108
rect 462 106 463 107
rect 444 104 463 106
rect 444 103 445 104
rect 439 102 445 103
rect 462 103 463 104
rect 467 103 468 107
rect 462 102 468 103
rect 471 107 477 108
rect 471 103 472 107
rect 476 106 477 107
rect 496 106 498 110
rect 476 104 498 106
rect 476 103 477 104
rect 471 102 477 103
rect 520 102 522 110
rect 544 102 546 110
rect 568 102 570 110
rect 593 102 595 110
rect 616 102 618 110
rect 640 102 642 110
rect 664 102 666 110
rect 688 102 690 110
rect 712 102 714 110
rect 736 102 738 110
rect 760 102 762 110
rect 784 102 786 110
rect 808 102 810 110
rect 832 102 834 110
rect 864 102 866 110
rect 896 102 898 110
rect 928 102 930 110
rect 960 102 962 110
rect 992 102 994 110
rect 1024 102 1026 110
rect 1054 107 1061 108
rect 1054 103 1055 107
rect 1060 103 1061 107
rect 1064 106 1066 112
rect 1079 111 1080 115
rect 1084 114 1085 115
rect 1094 114 1095 118
rect 1099 114 1100 118
rect 1118 118 1124 119
rect 1084 112 1090 114
rect 1094 113 1100 114
rect 1103 115 1109 116
rect 1084 111 1085 112
rect 1079 110 1085 111
rect 1079 107 1085 108
rect 1079 106 1080 107
rect 1064 104 1080 106
rect 1054 102 1061 103
rect 1079 103 1080 104
rect 1084 103 1085 107
rect 1088 106 1090 112
rect 1103 111 1104 115
rect 1108 114 1109 115
rect 1118 114 1119 118
rect 1123 114 1124 118
rect 1142 118 1148 119
rect 1108 112 1114 114
rect 1118 113 1124 114
rect 1127 115 1133 116
rect 1108 111 1109 112
rect 1103 110 1109 111
rect 1103 107 1109 108
rect 1103 106 1104 107
rect 1088 104 1104 106
rect 1079 102 1085 103
rect 1103 103 1104 104
rect 1108 103 1109 107
rect 1112 106 1114 112
rect 1127 111 1128 115
rect 1132 114 1133 115
rect 1142 114 1143 118
rect 1147 114 1148 118
rect 1174 118 1180 119
rect 1132 112 1138 114
rect 1142 113 1148 114
rect 1151 115 1157 116
rect 1132 111 1133 112
rect 1127 110 1133 111
rect 1127 107 1133 108
rect 1127 106 1128 107
rect 1112 104 1128 106
rect 1103 102 1109 103
rect 1127 103 1128 104
rect 1132 103 1133 107
rect 1136 106 1138 112
rect 1151 111 1152 115
rect 1156 114 1157 115
rect 1174 114 1175 118
rect 1179 114 1180 118
rect 1206 118 1212 119
rect 1156 112 1161 114
rect 1174 113 1180 114
rect 1183 115 1189 116
rect 1156 111 1157 112
rect 1151 110 1157 111
rect 1151 107 1157 108
rect 1151 106 1152 107
rect 1136 104 1152 106
rect 1127 102 1133 103
rect 1151 103 1152 104
rect 1156 103 1157 107
rect 1159 106 1161 112
rect 1183 111 1184 115
rect 1188 114 1189 115
rect 1206 114 1207 118
rect 1211 114 1212 118
rect 1238 118 1244 119
rect 1188 112 1202 114
rect 1206 113 1212 114
rect 1215 115 1221 116
rect 1188 111 1189 112
rect 1183 110 1189 111
rect 1183 107 1189 108
rect 1183 106 1184 107
rect 1159 104 1184 106
rect 1151 102 1157 103
rect 1183 103 1184 104
rect 1188 103 1189 107
rect 1200 106 1202 112
rect 1215 111 1216 115
rect 1220 114 1221 115
rect 1238 114 1239 118
rect 1243 114 1244 118
rect 1270 118 1276 119
rect 1220 112 1234 114
rect 1238 113 1244 114
rect 1247 115 1253 116
rect 1220 111 1221 112
rect 1215 110 1221 111
rect 1215 107 1221 108
rect 1215 106 1216 107
rect 1200 104 1216 106
rect 1183 102 1189 103
rect 1215 103 1216 104
rect 1220 103 1221 107
rect 1232 106 1234 112
rect 1247 111 1248 115
rect 1252 114 1253 115
rect 1270 114 1271 118
rect 1275 114 1276 118
rect 1302 118 1308 119
rect 1252 112 1266 114
rect 1270 113 1276 114
rect 1279 115 1285 116
rect 1252 111 1253 112
rect 1247 110 1253 111
rect 1247 107 1253 108
rect 1247 106 1248 107
rect 1232 104 1248 106
rect 1215 102 1221 103
rect 1247 103 1248 104
rect 1252 103 1253 107
rect 1264 106 1266 112
rect 1279 111 1280 115
rect 1284 114 1285 115
rect 1302 114 1303 118
rect 1307 114 1308 118
rect 1334 118 1340 119
rect 1284 112 1298 114
rect 1302 113 1308 114
rect 1311 115 1317 116
rect 1284 111 1285 112
rect 1279 110 1285 111
rect 1279 107 1285 108
rect 1279 106 1280 107
rect 1264 104 1280 106
rect 1247 102 1253 103
rect 1279 103 1280 104
rect 1284 103 1285 107
rect 1296 106 1298 112
rect 1311 111 1312 115
rect 1316 114 1317 115
rect 1334 114 1335 118
rect 1339 114 1340 118
rect 1343 115 1344 119
rect 1348 115 1349 119
rect 1343 114 1349 115
rect 1366 118 1372 119
rect 1366 114 1367 118
rect 1371 114 1372 118
rect 1390 118 1396 119
rect 1316 112 1330 114
rect 1334 113 1340 114
rect 1366 113 1372 114
rect 1375 115 1381 116
rect 1316 111 1317 112
rect 1311 110 1317 111
rect 1311 107 1317 108
rect 1311 106 1312 107
rect 1296 104 1312 106
rect 1279 102 1285 103
rect 1311 103 1312 104
rect 1316 103 1317 107
rect 1328 106 1330 112
rect 1375 111 1376 115
rect 1380 114 1381 115
rect 1390 114 1391 118
rect 1395 114 1396 118
rect 1414 118 1420 119
rect 1380 112 1386 114
rect 1390 113 1396 114
rect 1399 115 1405 116
rect 1380 111 1381 112
rect 1375 110 1381 111
rect 1343 107 1349 108
rect 1343 106 1344 107
rect 1328 104 1344 106
rect 1311 102 1317 103
rect 1343 103 1344 104
rect 1348 103 1349 107
rect 1343 102 1349 103
rect 1374 107 1381 108
rect 1374 103 1375 107
rect 1380 103 1381 107
rect 1374 102 1381 103
rect 1384 102 1386 112
rect 1399 111 1400 115
rect 1404 111 1405 115
rect 1414 114 1415 118
rect 1419 114 1420 118
rect 1423 115 1424 119
rect 1428 115 1429 119
rect 1423 114 1429 115
rect 1414 113 1420 114
rect 1446 113 1452 114
rect 1399 110 1405 111
rect 1401 106 1403 110
rect 1446 109 1447 113
rect 1451 109 1452 113
rect 1446 108 1452 109
rect 1423 107 1429 108
rect 1423 106 1424 107
rect 1401 104 1424 106
rect 1423 103 1424 104
rect 1428 103 1429 107
rect 1423 102 1429 103
rect 200 100 219 102
rect 265 100 291 102
rect 508 100 522 102
rect 532 100 546 102
rect 556 100 570 102
rect 580 100 595 102
rect 604 100 618 102
rect 628 100 642 102
rect 652 100 666 102
rect 676 100 690 102
rect 700 100 714 102
rect 724 100 738 102
rect 748 100 762 102
rect 772 100 786 102
rect 796 100 810 102
rect 820 100 834 102
rect 848 100 866 102
rect 880 100 898 102
rect 912 100 930 102
rect 944 100 962 102
rect 977 100 994 102
rect 1008 100 1026 102
rect 1384 100 1403 102
rect 215 99 221 100
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 215 95 216 99
rect 220 95 221 99
rect 215 94 221 95
rect 287 99 293 100
rect 287 95 288 99
rect 292 95 293 99
rect 287 94 293 95
rect 495 99 501 100
rect 495 95 496 99
rect 500 98 501 99
rect 508 98 510 100
rect 532 98 534 100
rect 556 98 558 100
rect 580 98 582 100
rect 604 98 606 100
rect 628 98 630 100
rect 652 98 654 100
rect 676 98 678 100
rect 700 98 702 100
rect 724 98 726 100
rect 748 98 750 100
rect 772 98 774 100
rect 796 98 798 100
rect 820 98 822 100
rect 500 96 510 98
rect 528 96 534 98
rect 552 96 558 98
rect 576 96 582 98
rect 593 96 606 98
rect 624 96 630 98
rect 649 96 654 98
rect 672 96 678 98
rect 697 96 702 98
rect 720 96 726 98
rect 745 96 750 98
rect 768 96 774 98
rect 792 96 798 98
rect 816 96 822 98
rect 500 95 501 96
rect 495 94 501 95
rect 519 95 525 96
rect 110 90 116 91
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 158 92 164 93
rect 158 88 159 92
rect 163 88 164 92
rect 158 87 164 88
rect 182 92 188 93
rect 182 88 183 92
rect 187 88 188 92
rect 182 87 188 88
rect 206 92 212 93
rect 206 88 207 92
rect 211 88 212 92
rect 206 87 212 88
rect 230 92 236 93
rect 230 88 231 92
rect 235 88 236 92
rect 230 87 236 88
rect 254 92 260 93
rect 278 92 284 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 263 91 269 92
rect 263 87 264 91
rect 268 87 269 91
rect 278 88 279 92
rect 283 88 284 92
rect 278 87 284 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 326 92 332 93
rect 326 88 327 92
rect 331 88 332 92
rect 326 87 332 88
rect 350 92 356 93
rect 350 88 351 92
rect 355 88 356 92
rect 350 87 356 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 398 92 404 93
rect 398 88 399 92
rect 403 88 404 92
rect 398 87 404 88
rect 430 92 436 93
rect 430 88 431 92
rect 435 88 436 92
rect 430 87 436 88
rect 462 92 468 93
rect 462 88 463 92
rect 467 88 468 92
rect 462 87 468 88
rect 486 92 492 93
rect 486 88 487 92
rect 491 88 492 92
rect 486 87 492 88
rect 510 92 516 93
rect 510 88 511 92
rect 515 88 516 92
rect 519 91 520 95
rect 524 94 525 95
rect 528 94 530 96
rect 524 92 530 94
rect 543 95 549 96
rect 534 92 540 93
rect 524 91 525 92
rect 519 90 525 91
rect 510 87 516 88
rect 534 88 535 92
rect 539 88 540 92
rect 543 91 544 95
rect 548 94 549 95
rect 552 94 554 96
rect 548 92 554 94
rect 567 95 573 96
rect 558 92 564 93
rect 548 91 549 92
rect 543 90 549 91
rect 534 87 540 88
rect 558 88 559 92
rect 563 88 564 92
rect 567 91 568 95
rect 572 94 573 95
rect 576 94 578 96
rect 572 92 578 94
rect 591 95 597 96
rect 582 92 588 93
rect 572 91 573 92
rect 567 90 573 91
rect 558 87 564 88
rect 582 88 583 92
rect 587 88 588 92
rect 591 91 592 95
rect 596 91 597 95
rect 615 95 621 96
rect 591 90 597 91
rect 606 92 612 93
rect 582 87 588 88
rect 606 88 607 92
rect 611 88 612 92
rect 615 91 616 95
rect 620 94 621 95
rect 624 94 626 96
rect 620 92 626 94
rect 639 95 645 96
rect 630 92 636 93
rect 620 91 621 92
rect 615 90 621 91
rect 606 87 612 88
rect 630 88 631 92
rect 635 88 636 92
rect 639 91 640 95
rect 644 94 645 95
rect 649 94 651 96
rect 644 92 651 94
rect 663 95 669 96
rect 654 92 660 93
rect 644 91 645 92
rect 639 90 645 91
rect 630 87 636 88
rect 654 88 655 92
rect 659 88 660 92
rect 663 91 664 95
rect 668 94 669 95
rect 672 94 674 96
rect 668 92 674 94
rect 687 95 693 96
rect 678 92 684 93
rect 668 91 669 92
rect 663 90 669 91
rect 654 87 660 88
rect 678 88 679 92
rect 683 88 684 92
rect 687 91 688 95
rect 692 94 693 95
rect 697 94 699 96
rect 692 92 699 94
rect 711 95 717 96
rect 702 92 708 93
rect 692 91 693 92
rect 687 90 693 91
rect 678 87 684 88
rect 702 88 703 92
rect 707 88 708 92
rect 711 91 712 95
rect 716 94 717 95
rect 720 94 722 96
rect 716 92 722 94
rect 735 95 741 96
rect 726 92 732 93
rect 716 91 717 92
rect 711 90 717 91
rect 702 87 708 88
rect 726 88 727 92
rect 731 88 732 92
rect 735 91 736 95
rect 740 94 741 95
rect 745 94 747 96
rect 740 92 747 94
rect 759 95 765 96
rect 750 92 756 93
rect 740 91 741 92
rect 735 90 741 91
rect 726 87 732 88
rect 750 88 751 92
rect 755 88 756 92
rect 759 91 760 95
rect 764 94 765 95
rect 768 94 770 96
rect 764 92 770 94
rect 783 95 789 96
rect 774 92 780 93
rect 764 91 765 92
rect 759 90 765 91
rect 750 87 756 88
rect 774 88 775 92
rect 779 88 780 92
rect 783 91 784 95
rect 788 94 789 95
rect 792 94 794 96
rect 788 92 794 94
rect 807 95 813 96
rect 798 92 804 93
rect 788 91 789 92
rect 783 90 789 91
rect 774 87 780 88
rect 798 88 799 92
rect 803 88 804 92
rect 807 91 808 95
rect 812 94 813 95
rect 816 94 818 96
rect 812 92 818 94
rect 831 95 837 96
rect 822 92 828 93
rect 812 91 813 92
rect 807 90 813 91
rect 798 87 804 88
rect 822 88 823 92
rect 827 88 828 92
rect 831 91 832 95
rect 836 94 837 95
rect 848 94 850 100
rect 836 92 850 94
rect 863 95 869 96
rect 854 92 860 93
rect 836 91 837 92
rect 831 90 837 91
rect 822 87 828 88
rect 854 88 855 92
rect 859 88 860 92
rect 863 91 864 95
rect 868 94 869 95
rect 880 94 882 100
rect 868 92 882 94
rect 895 95 901 96
rect 886 92 892 93
rect 868 91 869 92
rect 863 90 869 91
rect 854 87 860 88
rect 886 88 887 92
rect 891 88 892 92
rect 895 91 896 95
rect 900 94 901 95
rect 912 94 914 100
rect 900 92 914 94
rect 927 95 933 96
rect 918 92 924 93
rect 900 91 901 92
rect 895 90 901 91
rect 886 87 892 88
rect 918 88 919 92
rect 923 88 924 92
rect 927 91 928 95
rect 932 94 933 95
rect 944 94 946 100
rect 932 92 946 94
rect 959 95 965 96
rect 950 92 956 93
rect 932 91 933 92
rect 927 90 933 91
rect 918 87 924 88
rect 950 88 951 92
rect 955 88 956 92
rect 959 91 960 95
rect 964 94 965 95
rect 977 94 979 100
rect 964 92 979 94
rect 991 95 997 96
rect 982 92 988 93
rect 964 91 965 92
rect 959 90 965 91
rect 950 87 956 88
rect 982 88 983 92
rect 987 88 988 92
rect 991 91 992 95
rect 996 94 997 95
rect 1008 94 1010 100
rect 1399 99 1405 100
rect 996 92 1010 94
rect 1023 95 1032 96
rect 1014 92 1020 93
rect 996 91 997 92
rect 991 90 997 91
rect 982 87 988 88
rect 1014 88 1015 92
rect 1019 88 1020 92
rect 1023 91 1024 95
rect 1031 91 1032 95
rect 1399 95 1400 99
rect 1404 95 1405 99
rect 1399 94 1405 95
rect 1446 95 1452 96
rect 1023 90 1032 91
rect 1046 92 1052 93
rect 1014 87 1020 88
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1046 87 1052 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1094 92 1100 93
rect 1094 88 1095 92
rect 1099 88 1100 92
rect 1094 87 1100 88
rect 1118 92 1124 93
rect 1118 88 1119 92
rect 1123 88 1124 92
rect 1118 87 1124 88
rect 1142 92 1148 93
rect 1142 88 1143 92
rect 1147 88 1148 92
rect 1142 87 1148 88
rect 1174 92 1180 93
rect 1174 88 1175 92
rect 1179 88 1180 92
rect 1174 87 1180 88
rect 1206 92 1212 93
rect 1206 88 1207 92
rect 1211 88 1212 92
rect 1206 87 1212 88
rect 1238 92 1244 93
rect 1238 88 1239 92
rect 1243 88 1244 92
rect 1238 87 1244 88
rect 1270 92 1276 93
rect 1270 88 1271 92
rect 1275 88 1276 92
rect 1270 87 1276 88
rect 1302 92 1308 93
rect 1302 88 1303 92
rect 1307 88 1308 92
rect 1302 87 1308 88
rect 1334 92 1340 93
rect 1334 88 1335 92
rect 1339 88 1340 92
rect 1334 87 1340 88
rect 1366 92 1372 93
rect 1366 88 1367 92
rect 1371 88 1372 92
rect 1366 87 1372 88
rect 1390 92 1396 93
rect 1390 88 1391 92
rect 1395 88 1396 92
rect 1390 87 1396 88
rect 1414 92 1420 93
rect 1414 88 1415 92
rect 1419 88 1420 92
rect 1446 91 1447 95
rect 1451 91 1452 95
rect 1446 90 1452 91
rect 1414 87 1420 88
rect 263 86 269 87
rect 242 83 248 84
rect 242 79 243 83
rect 247 82 248 83
rect 265 82 267 86
rect 247 80 267 82
rect 247 79 248 80
rect 242 78 248 79
<< m3c >>
rect 819 1507 823 1511
rect 295 1498 299 1502
rect 111 1493 115 1497
rect 319 1498 323 1502
rect 343 1498 347 1502
rect 367 1498 371 1502
rect 407 1498 411 1502
rect 455 1498 459 1502
rect 511 1498 515 1502
rect 575 1498 579 1502
rect 647 1498 651 1502
rect 727 1498 731 1502
rect 807 1498 811 1502
rect 887 1498 891 1502
rect 959 1498 963 1502
rect 1031 1498 1035 1502
rect 1083 1495 1087 1499
rect 1103 1498 1107 1502
rect 1115 1495 1116 1499
rect 1116 1495 1119 1499
rect 1175 1498 1179 1502
rect 1247 1498 1251 1502
rect 1103 1487 1107 1491
rect 111 1475 115 1479
rect 819 1479 820 1483
rect 820 1479 823 1483
rect 1447 1493 1451 1497
rect 295 1472 299 1476
rect 307 1471 308 1475
rect 308 1471 311 1475
rect 319 1472 323 1476
rect 343 1472 347 1476
rect 367 1472 371 1476
rect 407 1472 411 1476
rect 455 1472 459 1476
rect 511 1472 515 1476
rect 575 1472 579 1476
rect 647 1472 651 1476
rect 727 1472 731 1476
rect 807 1472 811 1476
rect 887 1472 891 1476
rect 959 1472 963 1476
rect 1031 1472 1035 1476
rect 1103 1472 1107 1476
rect 1175 1472 1179 1476
rect 1247 1472 1251 1476
rect 1447 1475 1451 1479
rect 111 1457 115 1461
rect 151 1460 155 1464
rect 175 1460 179 1464
rect 199 1460 203 1464
rect 231 1460 235 1464
rect 271 1460 275 1464
rect 319 1460 323 1464
rect 367 1460 371 1464
rect 407 1460 411 1464
rect 455 1460 459 1464
rect 503 1460 507 1464
rect 551 1460 555 1464
rect 607 1460 611 1464
rect 663 1460 667 1464
rect 711 1460 715 1464
rect 759 1460 763 1464
rect 815 1460 819 1464
rect 871 1460 875 1464
rect 927 1460 931 1464
rect 975 1460 979 1464
rect 1023 1460 1027 1464
rect 1071 1460 1075 1464
rect 1083 1459 1084 1463
rect 1084 1459 1087 1463
rect 1119 1460 1123 1464
rect 1167 1460 1171 1464
rect 1215 1460 1219 1464
rect 1263 1460 1267 1464
rect 1311 1460 1315 1464
rect 1447 1457 1451 1461
rect 427 1451 431 1455
rect 827 1451 831 1455
rect 987 1451 991 1455
rect 1227 1451 1231 1455
rect 1323 1451 1327 1455
rect 111 1439 115 1443
rect 151 1434 155 1438
rect 175 1434 179 1438
rect 199 1434 203 1438
rect 231 1434 235 1438
rect 271 1434 275 1438
rect 319 1434 323 1438
rect 367 1434 371 1438
rect 207 1427 211 1431
rect 299 1427 303 1431
rect 307 1427 311 1431
rect 407 1434 411 1438
rect 455 1434 459 1438
rect 503 1434 507 1438
rect 551 1434 555 1438
rect 607 1434 611 1438
rect 663 1434 667 1438
rect 711 1434 715 1438
rect 559 1427 563 1431
rect 759 1434 763 1438
rect 815 1434 819 1438
rect 827 1435 828 1439
rect 828 1435 831 1439
rect 871 1434 875 1438
rect 927 1434 931 1438
rect 975 1434 979 1438
rect 987 1435 988 1439
rect 988 1435 991 1439
rect 1035 1443 1036 1447
rect 1036 1443 1039 1447
rect 1023 1434 1027 1438
rect 1071 1434 1075 1438
rect 1119 1434 1123 1438
rect 1131 1431 1132 1435
rect 1132 1431 1135 1435
rect 1167 1434 1171 1438
rect 1215 1434 1219 1438
rect 1227 1435 1228 1439
rect 1228 1435 1231 1439
rect 1275 1443 1279 1447
rect 1263 1434 1267 1438
rect 1311 1434 1315 1438
rect 1323 1435 1324 1439
rect 1324 1435 1327 1439
rect 1447 1439 1451 1443
rect 1355 1427 1359 1431
rect 135 1418 139 1422
rect 111 1413 115 1417
rect 159 1418 163 1422
rect 183 1418 187 1422
rect 223 1418 227 1422
rect 287 1418 291 1422
rect 351 1418 355 1422
rect 415 1418 419 1422
rect 427 1419 428 1423
rect 428 1419 431 1423
rect 479 1418 483 1422
rect 535 1418 539 1422
rect 583 1418 587 1422
rect 559 1407 563 1411
rect 631 1418 635 1422
rect 687 1418 691 1422
rect 743 1418 747 1422
rect 799 1418 803 1422
rect 855 1418 859 1422
rect 891 1415 895 1419
rect 911 1418 915 1422
rect 967 1418 971 1422
rect 1023 1418 1027 1422
rect 1035 1419 1036 1423
rect 1036 1419 1039 1423
rect 1071 1418 1075 1422
rect 1083 1415 1084 1419
rect 1084 1415 1087 1419
rect 1119 1418 1123 1422
rect 1139 1415 1143 1419
rect 1167 1418 1171 1422
rect 1215 1418 1219 1422
rect 111 1395 115 1399
rect 1119 1403 1123 1407
rect 1131 1407 1132 1411
rect 1132 1407 1135 1411
rect 1263 1418 1267 1422
rect 1275 1419 1276 1423
rect 1276 1419 1279 1423
rect 1303 1418 1307 1422
rect 1315 1415 1316 1419
rect 1316 1415 1319 1419
rect 1343 1418 1347 1422
rect 1391 1418 1395 1422
rect 1415 1418 1419 1422
rect 1447 1413 1451 1417
rect 1355 1399 1356 1403
rect 1356 1399 1359 1403
rect 135 1392 139 1396
rect 147 1391 148 1395
rect 148 1391 151 1395
rect 159 1392 163 1396
rect 183 1392 187 1396
rect 223 1392 227 1396
rect 287 1392 291 1396
rect 351 1392 355 1396
rect 415 1392 419 1396
rect 479 1392 483 1396
rect 535 1392 539 1396
rect 583 1392 587 1396
rect 631 1392 635 1396
rect 687 1392 691 1396
rect 743 1392 747 1396
rect 799 1392 803 1396
rect 855 1392 859 1396
rect 911 1392 915 1396
rect 947 1391 951 1395
rect 967 1392 971 1396
rect 1023 1392 1027 1396
rect 1071 1392 1075 1396
rect 1119 1392 1123 1396
rect 1167 1392 1171 1396
rect 1207 1391 1211 1395
rect 1215 1392 1219 1396
rect 1263 1392 1267 1396
rect 1303 1392 1307 1396
rect 1343 1392 1347 1396
rect 1391 1392 1395 1396
rect 1415 1392 1419 1396
rect 1427 1391 1428 1395
rect 1428 1391 1431 1395
rect 1447 1395 1451 1399
rect 111 1377 115 1381
rect 135 1380 139 1384
rect 159 1380 163 1384
rect 183 1380 187 1384
rect 231 1380 235 1384
rect 279 1380 283 1384
rect 335 1380 339 1384
rect 391 1380 395 1384
rect 439 1380 443 1384
rect 487 1380 491 1384
rect 527 1380 531 1384
rect 567 1380 571 1384
rect 615 1380 619 1384
rect 663 1380 667 1384
rect 711 1380 715 1384
rect 767 1380 771 1384
rect 823 1380 827 1384
rect 879 1380 883 1384
rect 891 1379 892 1383
rect 892 1379 895 1383
rect 935 1380 939 1384
rect 991 1380 995 1384
rect 1047 1380 1051 1384
rect 1083 1379 1087 1383
rect 1095 1380 1099 1384
rect 1143 1380 1147 1384
rect 1191 1380 1195 1384
rect 1239 1380 1243 1384
rect 1287 1380 1291 1384
rect 1315 1379 1319 1383
rect 1335 1380 1339 1384
rect 1383 1380 1387 1384
rect 1415 1380 1419 1384
rect 1447 1377 1451 1381
rect 171 1371 175 1375
rect 111 1359 115 1363
rect 195 1371 199 1375
rect 291 1371 295 1375
rect 299 1371 303 1375
rect 451 1371 455 1375
rect 539 1371 543 1375
rect 627 1371 631 1375
rect 135 1354 139 1358
rect 147 1355 148 1359
rect 148 1355 151 1359
rect 159 1354 163 1358
rect 171 1355 172 1359
rect 172 1355 175 1359
rect 183 1354 187 1358
rect 195 1355 196 1359
rect 196 1355 199 1359
rect 207 1347 211 1351
rect 723 1371 727 1375
rect 835 1371 839 1375
rect 1003 1371 1007 1375
rect 1395 1371 1399 1375
rect 1427 1371 1431 1375
rect 231 1354 235 1358
rect 279 1354 283 1358
rect 291 1355 292 1359
rect 292 1355 295 1359
rect 335 1354 339 1358
rect 391 1354 395 1358
rect 319 1347 323 1351
rect 439 1354 443 1358
rect 451 1355 452 1359
rect 452 1355 455 1359
rect 487 1354 491 1358
rect 527 1354 531 1358
rect 539 1355 540 1359
rect 540 1355 543 1359
rect 567 1354 571 1358
rect 495 1347 499 1351
rect 615 1354 619 1358
rect 627 1355 628 1359
rect 628 1355 631 1359
rect 167 1338 171 1342
rect 191 1338 195 1342
rect 111 1333 115 1337
rect 231 1338 235 1342
rect 279 1338 283 1342
rect 335 1338 339 1342
rect 391 1338 395 1342
rect 411 1335 415 1339
rect 455 1338 459 1342
rect 519 1338 523 1342
rect 575 1338 579 1342
rect 1019 1363 1023 1367
rect 663 1354 667 1358
rect 711 1354 715 1358
rect 723 1355 724 1359
rect 724 1355 727 1359
rect 767 1354 771 1358
rect 691 1347 695 1351
rect 823 1354 827 1358
rect 835 1355 836 1359
rect 836 1355 839 1359
rect 879 1354 883 1358
rect 935 1354 939 1358
rect 947 1355 948 1359
rect 948 1355 951 1359
rect 991 1354 995 1358
rect 1003 1355 1004 1359
rect 1004 1355 1007 1359
rect 1047 1354 1051 1358
rect 1171 1363 1175 1367
rect 1095 1354 1099 1358
rect 1115 1351 1119 1355
rect 1143 1354 1147 1358
rect 1191 1354 1195 1358
rect 1239 1354 1243 1358
rect 1207 1347 1211 1351
rect 1287 1354 1291 1358
rect 1335 1354 1339 1358
rect 1375 1351 1379 1355
rect 1383 1354 1387 1358
rect 1395 1355 1396 1359
rect 1396 1355 1399 1359
rect 1427 1363 1428 1367
rect 1428 1363 1431 1367
rect 1447 1359 1451 1363
rect 1415 1354 1419 1358
rect 631 1338 635 1342
rect 679 1338 683 1342
rect 727 1338 731 1342
rect 111 1315 115 1319
rect 319 1323 323 1327
rect 327 1323 331 1327
rect 691 1327 692 1331
rect 692 1327 695 1331
rect 767 1338 771 1342
rect 799 1338 803 1342
rect 831 1338 835 1342
rect 863 1338 867 1342
rect 895 1338 899 1342
rect 927 1338 931 1342
rect 967 1338 971 1342
rect 979 1335 980 1339
rect 980 1335 983 1339
rect 1007 1338 1011 1342
rect 1019 1339 1020 1343
rect 1020 1339 1023 1343
rect 1055 1338 1059 1342
rect 1103 1338 1107 1342
rect 1123 1335 1127 1339
rect 1159 1338 1163 1342
rect 1171 1339 1172 1343
rect 1172 1339 1175 1343
rect 1215 1338 1219 1342
rect 1271 1338 1275 1342
rect 1315 1335 1319 1339
rect 1327 1338 1331 1342
rect 1383 1338 1387 1342
rect 1415 1338 1419 1342
rect 1427 1339 1428 1343
rect 1428 1339 1431 1343
rect 1115 1327 1116 1331
rect 1116 1327 1119 1331
rect 1447 1333 1451 1337
rect 167 1312 171 1316
rect 191 1312 195 1316
rect 231 1312 235 1316
rect 279 1312 283 1316
rect 335 1312 339 1316
rect 391 1312 395 1316
rect 455 1312 459 1316
rect 519 1312 523 1316
rect 575 1312 579 1316
rect 631 1312 635 1316
rect 495 1307 499 1311
rect 671 1311 675 1315
rect 679 1312 683 1316
rect 727 1312 731 1316
rect 767 1312 771 1316
rect 799 1312 803 1316
rect 831 1312 835 1316
rect 863 1312 867 1316
rect 895 1312 899 1316
rect 927 1312 931 1316
rect 967 1312 971 1316
rect 1007 1312 1011 1316
rect 1055 1312 1059 1316
rect 1083 1311 1087 1315
rect 1103 1312 1107 1316
rect 1159 1312 1163 1316
rect 1215 1312 1219 1316
rect 1259 1311 1263 1315
rect 1271 1312 1275 1316
rect 1327 1312 1331 1316
rect 1383 1312 1387 1316
rect 1415 1312 1419 1316
rect 1427 1311 1428 1315
rect 1428 1311 1431 1315
rect 1447 1315 1451 1319
rect 1375 1307 1379 1311
rect 111 1297 115 1301
rect 231 1300 235 1304
rect 255 1300 259 1304
rect 279 1300 283 1304
rect 303 1300 307 1304
rect 327 1300 331 1304
rect 351 1300 355 1304
rect 375 1300 379 1304
rect 399 1300 403 1304
rect 423 1300 427 1304
rect 447 1300 451 1304
rect 471 1300 475 1304
rect 503 1300 507 1304
rect 543 1300 547 1304
rect 591 1300 595 1304
rect 647 1300 651 1304
rect 695 1300 699 1304
rect 743 1300 747 1304
rect 791 1300 795 1304
rect 839 1300 843 1304
rect 879 1300 883 1304
rect 911 1300 915 1304
rect 951 1300 955 1304
rect 991 1300 995 1304
rect 1031 1300 1035 1304
rect 1071 1300 1075 1304
rect 1111 1300 1115 1304
rect 1123 1299 1124 1303
rect 1124 1299 1127 1303
rect 1151 1300 1155 1304
rect 1199 1300 1203 1304
rect 1247 1300 1251 1304
rect 1303 1300 1307 1304
rect 1315 1299 1316 1303
rect 1316 1299 1319 1303
rect 1367 1300 1371 1304
rect 1415 1300 1419 1304
rect 1447 1297 1451 1301
rect 267 1291 271 1295
rect 339 1291 343 1295
rect 411 1291 415 1295
rect 755 1291 759 1295
rect 979 1291 983 1295
rect 111 1279 115 1283
rect 319 1283 323 1287
rect 231 1274 235 1278
rect 243 1275 244 1279
rect 244 1275 247 1279
rect 255 1274 259 1278
rect 267 1275 268 1279
rect 268 1275 271 1279
rect 279 1274 283 1278
rect 303 1274 307 1278
rect 327 1274 331 1278
rect 339 1275 340 1279
rect 340 1275 343 1279
rect 351 1274 355 1278
rect 363 1275 364 1279
rect 364 1275 367 1279
rect 375 1274 379 1278
rect 319 1263 323 1267
rect 343 1267 347 1271
rect 399 1274 403 1278
rect 423 1274 427 1278
rect 447 1274 451 1278
rect 471 1274 475 1278
rect 503 1274 507 1278
rect 543 1274 547 1278
rect 591 1274 595 1278
rect 671 1283 675 1287
rect 647 1274 651 1278
rect 531 1267 535 1271
rect 695 1274 699 1278
rect 743 1274 747 1278
rect 755 1275 756 1279
rect 756 1275 759 1279
rect 791 1274 795 1278
rect 839 1274 843 1278
rect 879 1274 883 1278
rect 911 1274 915 1278
rect 951 1274 955 1278
rect 991 1274 995 1278
rect 1031 1274 1035 1278
rect 1139 1283 1143 1287
rect 1071 1274 1075 1278
rect 1083 1275 1084 1279
rect 1084 1275 1087 1279
rect 1111 1274 1115 1278
rect 1151 1274 1155 1278
rect 1199 1274 1203 1278
rect 1247 1274 1251 1278
rect 1259 1275 1260 1279
rect 1260 1275 1263 1279
rect 1303 1274 1307 1278
rect 1387 1283 1391 1287
rect 1367 1274 1371 1278
rect 1003 1267 1007 1271
rect 1295 1267 1299 1271
rect 1323 1267 1327 1271
rect 1415 1274 1419 1278
rect 1427 1275 1428 1279
rect 1428 1275 1431 1279
rect 1447 1279 1451 1283
rect 311 1258 315 1262
rect 335 1258 339 1262
rect 111 1253 115 1257
rect 359 1258 363 1262
rect 383 1258 387 1262
rect 415 1258 419 1262
rect 367 1247 368 1251
rect 368 1247 371 1251
rect 447 1258 451 1262
rect 479 1258 483 1262
rect 519 1258 523 1262
rect 559 1258 563 1262
rect 615 1258 619 1262
rect 679 1258 683 1262
rect 691 1255 692 1259
rect 692 1255 695 1259
rect 751 1258 755 1262
rect 831 1258 835 1262
rect 911 1258 915 1262
rect 991 1258 995 1262
rect 1063 1258 1067 1262
rect 1127 1258 1131 1262
rect 1139 1259 1140 1263
rect 1140 1259 1143 1263
rect 1191 1258 1195 1262
rect 1003 1247 1004 1251
rect 1004 1247 1007 1251
rect 1247 1258 1251 1262
rect 1311 1258 1315 1262
rect 1375 1258 1379 1262
rect 1387 1259 1388 1263
rect 1388 1259 1391 1263
rect 1415 1258 1419 1262
rect 1323 1247 1324 1251
rect 1324 1247 1327 1251
rect 1447 1253 1451 1257
rect 111 1235 115 1239
rect 347 1239 348 1243
rect 348 1239 351 1243
rect 531 1239 532 1243
rect 532 1239 535 1243
rect 311 1232 315 1236
rect 335 1232 339 1236
rect 359 1232 363 1236
rect 383 1232 387 1236
rect 415 1232 419 1236
rect 447 1232 451 1236
rect 479 1232 483 1236
rect 519 1232 523 1236
rect 559 1232 563 1236
rect 615 1232 619 1236
rect 679 1232 683 1236
rect 751 1232 755 1236
rect 763 1231 764 1235
rect 764 1231 767 1235
rect 831 1232 835 1236
rect 911 1232 915 1236
rect 991 1232 995 1236
rect 1063 1232 1067 1236
rect 1127 1232 1131 1236
rect 1191 1232 1195 1236
rect 1247 1232 1251 1236
rect 1311 1232 1315 1236
rect 1375 1232 1379 1236
rect 1415 1232 1419 1236
rect 1427 1231 1428 1235
rect 1428 1231 1431 1235
rect 1447 1235 1451 1239
rect 111 1217 115 1221
rect 327 1220 331 1224
rect 367 1220 371 1224
rect 407 1220 411 1224
rect 447 1220 451 1224
rect 487 1220 491 1224
rect 527 1220 531 1224
rect 567 1220 571 1224
rect 607 1220 611 1224
rect 655 1220 659 1224
rect 703 1220 707 1224
rect 751 1220 755 1224
rect 799 1220 803 1224
rect 847 1220 851 1224
rect 895 1220 899 1224
rect 943 1220 947 1224
rect 991 1220 995 1224
rect 1039 1220 1043 1224
rect 1103 1220 1107 1224
rect 1175 1220 1179 1224
rect 1255 1220 1259 1224
rect 1343 1220 1347 1224
rect 1415 1220 1419 1224
rect 1447 1217 1451 1221
rect 459 1211 463 1215
rect 691 1211 695 1215
rect 811 1211 815 1215
rect 907 1211 911 1215
rect 1003 1211 1007 1215
rect 1115 1211 1119 1215
rect 1267 1211 1271 1215
rect 1295 1211 1299 1215
rect 111 1199 115 1203
rect 347 1203 351 1207
rect 327 1194 331 1198
rect 367 1194 371 1198
rect 407 1194 411 1198
rect 447 1194 451 1198
rect 459 1195 460 1199
rect 460 1195 463 1199
rect 487 1194 491 1198
rect 527 1194 531 1198
rect 567 1194 571 1198
rect 607 1194 611 1198
rect 655 1194 659 1198
rect 703 1194 707 1198
rect 171 1187 175 1191
rect 415 1187 419 1191
rect 695 1187 699 1191
rect 751 1194 755 1198
rect 763 1195 764 1199
rect 764 1195 767 1199
rect 799 1194 803 1198
rect 811 1195 812 1199
rect 812 1195 815 1199
rect 779 1187 783 1191
rect 923 1203 927 1207
rect 847 1194 851 1198
rect 895 1194 899 1198
rect 907 1195 908 1199
rect 908 1195 911 1199
rect 943 1194 947 1198
rect 991 1194 995 1198
rect 1003 1195 1004 1199
rect 1004 1195 1007 1199
rect 1039 1194 1043 1198
rect 1103 1194 1107 1198
rect 1115 1195 1116 1199
rect 1116 1195 1119 1199
rect 1115 1187 1119 1191
rect 1175 1194 1179 1198
rect 1255 1194 1259 1198
rect 1267 1195 1268 1199
rect 1268 1195 1271 1199
rect 1283 1187 1287 1191
rect 1343 1194 1347 1198
rect 1415 1194 1419 1198
rect 1427 1195 1428 1199
rect 1428 1195 1431 1199
rect 1447 1199 1451 1203
rect 135 1178 139 1182
rect 159 1178 163 1182
rect 111 1173 115 1177
rect 183 1178 187 1182
rect 207 1178 211 1182
rect 231 1178 235 1182
rect 255 1178 259 1182
rect 279 1178 283 1182
rect 303 1178 307 1182
rect 315 1175 316 1179
rect 316 1175 319 1179
rect 335 1178 339 1182
rect 347 1179 348 1183
rect 348 1179 351 1183
rect 383 1178 387 1182
rect 423 1178 427 1182
rect 463 1178 467 1182
rect 503 1178 507 1182
rect 543 1178 547 1182
rect 583 1178 587 1182
rect 623 1178 627 1182
rect 671 1178 675 1182
rect 719 1178 723 1182
rect 767 1178 771 1182
rect 815 1178 819 1182
rect 863 1178 867 1182
rect 111 1155 115 1159
rect 399 1163 403 1167
rect 911 1178 915 1182
rect 923 1179 924 1183
rect 924 1179 927 1183
rect 959 1178 963 1182
rect 999 1175 1003 1179
rect 1007 1178 1011 1182
rect 1055 1178 1059 1182
rect 1103 1178 1107 1182
rect 1151 1178 1155 1182
rect 1183 1175 1187 1179
rect 1191 1178 1195 1182
rect 1231 1178 1235 1182
rect 1271 1178 1275 1182
rect 1311 1178 1315 1182
rect 1351 1178 1355 1182
rect 1363 1175 1364 1179
rect 1364 1175 1367 1179
rect 1391 1178 1395 1182
rect 1415 1178 1419 1182
rect 1447 1173 1451 1177
rect 135 1152 139 1156
rect 147 1151 148 1155
rect 148 1151 151 1155
rect 159 1152 163 1156
rect 171 1151 172 1155
rect 172 1151 175 1155
rect 183 1152 187 1156
rect 207 1152 211 1156
rect 231 1152 235 1156
rect 255 1152 259 1156
rect 279 1152 283 1156
rect 303 1152 307 1156
rect 335 1152 339 1156
rect 383 1152 387 1156
rect 415 1155 419 1159
rect 423 1152 427 1156
rect 463 1152 467 1156
rect 503 1152 507 1156
rect 543 1152 547 1156
rect 583 1152 587 1156
rect 623 1152 627 1156
rect 671 1152 675 1156
rect 719 1152 723 1156
rect 767 1152 771 1156
rect 779 1155 780 1159
rect 780 1155 783 1159
rect 815 1152 819 1156
rect 863 1152 867 1156
rect 911 1152 915 1156
rect 959 1152 963 1156
rect 1007 1152 1011 1156
rect 1055 1152 1059 1156
rect 1103 1152 1107 1156
rect 1115 1155 1116 1159
rect 1116 1155 1119 1159
rect 1151 1152 1155 1156
rect 823 1147 827 1151
rect 1183 1151 1187 1155
rect 1191 1152 1195 1156
rect 1203 1155 1204 1159
rect 1204 1155 1207 1159
rect 1231 1152 1235 1156
rect 1271 1152 1275 1156
rect 1283 1151 1284 1155
rect 1284 1151 1287 1155
rect 1311 1152 1315 1156
rect 1351 1152 1355 1156
rect 1391 1152 1395 1156
rect 1403 1151 1404 1155
rect 1404 1151 1407 1155
rect 1415 1152 1419 1156
rect 1447 1155 1451 1159
rect 111 1137 115 1141
rect 135 1140 139 1144
rect 159 1140 163 1144
rect 183 1140 187 1144
rect 215 1140 219 1144
rect 255 1140 259 1144
rect 295 1140 299 1144
rect 335 1140 339 1144
rect 375 1140 379 1144
rect 415 1140 419 1144
rect 463 1140 467 1144
rect 519 1140 523 1144
rect 583 1140 587 1144
rect 647 1140 651 1144
rect 711 1140 715 1144
rect 767 1140 771 1144
rect 831 1140 835 1144
rect 887 1140 891 1144
rect 943 1140 947 1144
rect 999 1140 1003 1144
rect 1055 1140 1059 1144
rect 1103 1140 1107 1144
rect 1151 1140 1155 1144
rect 1191 1140 1195 1144
rect 1231 1140 1235 1144
rect 1271 1140 1275 1144
rect 1311 1140 1315 1144
rect 1351 1140 1355 1144
rect 1391 1140 1395 1144
rect 1415 1140 1419 1144
rect 1447 1137 1451 1141
rect 171 1131 175 1135
rect 315 1131 319 1135
rect 427 1131 431 1135
rect 531 1131 535 1135
rect 659 1131 663 1135
rect 695 1131 699 1135
rect 899 1131 903 1135
rect 1011 1131 1015 1135
rect 1019 1131 1023 1135
rect 1363 1131 1367 1135
rect 111 1119 115 1123
rect 195 1123 196 1127
rect 196 1123 199 1127
rect 135 1114 139 1118
rect 147 1115 148 1119
rect 148 1115 151 1119
rect 159 1114 163 1118
rect 171 1115 172 1119
rect 172 1115 175 1119
rect 183 1114 187 1118
rect 215 1114 219 1118
rect 255 1114 259 1118
rect 295 1114 299 1118
rect 335 1114 339 1118
rect 399 1123 403 1127
rect 375 1114 379 1118
rect 387 1111 388 1115
rect 388 1111 391 1115
rect 415 1114 419 1118
rect 427 1115 428 1119
rect 428 1115 431 1119
rect 463 1114 467 1118
rect 519 1114 523 1118
rect 531 1115 532 1119
rect 532 1115 535 1119
rect 583 1114 587 1118
rect 647 1114 651 1118
rect 659 1115 660 1119
rect 660 1115 663 1119
rect 711 1114 715 1118
rect 767 1114 771 1118
rect 823 1115 827 1119
rect 831 1114 835 1118
rect 887 1114 891 1118
rect 899 1115 900 1119
rect 900 1115 903 1119
rect 943 1114 947 1118
rect 999 1114 1003 1118
rect 1011 1115 1012 1119
rect 1012 1115 1015 1119
rect 1055 1114 1059 1118
rect 1103 1114 1107 1118
rect 1151 1114 1155 1118
rect 1191 1114 1195 1118
rect 1231 1114 1235 1118
rect 135 1094 139 1098
rect 111 1089 115 1093
rect 159 1094 163 1098
rect 183 1094 187 1098
rect 195 1095 196 1099
rect 196 1095 199 1099
rect 207 1094 211 1098
rect 219 1091 220 1095
rect 220 1091 223 1095
rect 247 1094 251 1098
rect 287 1094 291 1098
rect 327 1094 331 1098
rect 1123 1103 1127 1107
rect 1183 1107 1187 1111
rect 1271 1114 1275 1118
rect 1311 1114 1315 1118
rect 1427 1123 1428 1127
rect 1428 1123 1431 1127
rect 1351 1114 1355 1118
rect 1391 1114 1395 1118
rect 1403 1115 1404 1119
rect 1404 1115 1407 1119
rect 1415 1114 1419 1118
rect 1447 1119 1451 1123
rect 1339 1103 1343 1107
rect 367 1094 371 1098
rect 379 1091 380 1095
rect 380 1091 383 1095
rect 407 1094 411 1098
rect 455 1094 459 1098
rect 503 1094 507 1098
rect 111 1071 115 1075
rect 135 1068 139 1072
rect 144 1071 148 1075
rect 367 1079 371 1083
rect 387 1083 391 1087
rect 559 1094 563 1098
rect 607 1094 611 1098
rect 619 1091 620 1095
rect 620 1091 623 1095
rect 655 1094 659 1098
rect 703 1094 707 1098
rect 743 1094 747 1098
rect 791 1094 795 1098
rect 839 1094 843 1098
rect 887 1094 891 1098
rect 943 1094 947 1098
rect 999 1094 1003 1098
rect 1011 1091 1012 1095
rect 1012 1091 1015 1095
rect 1055 1094 1059 1098
rect 1111 1094 1115 1098
rect 1167 1094 1171 1098
rect 1215 1094 1219 1098
rect 1263 1091 1267 1095
rect 1271 1094 1275 1098
rect 1327 1094 1331 1098
rect 1383 1094 1387 1098
rect 1415 1094 1419 1098
rect 1427 1095 1428 1099
rect 1428 1095 1431 1099
rect 1123 1075 1124 1079
rect 1124 1075 1127 1079
rect 1139 1079 1143 1083
rect 1447 1089 1451 1093
rect 159 1068 163 1072
rect 183 1068 187 1072
rect 207 1068 211 1072
rect 247 1068 251 1072
rect 287 1068 291 1072
rect 299 1067 300 1071
rect 300 1067 303 1071
rect 327 1068 331 1072
rect 367 1068 371 1072
rect 407 1068 411 1072
rect 455 1068 459 1072
rect 503 1068 507 1072
rect 559 1068 563 1072
rect 607 1068 611 1072
rect 655 1068 659 1072
rect 695 1067 699 1071
rect 703 1068 707 1072
rect 743 1068 747 1072
rect 791 1068 795 1072
rect 839 1068 843 1072
rect 887 1068 891 1072
rect 943 1068 947 1072
rect 999 1068 1003 1072
rect 1055 1068 1059 1072
rect 1111 1068 1115 1072
rect 1167 1068 1171 1072
rect 1215 1068 1219 1072
rect 1271 1068 1275 1072
rect 1327 1068 1331 1072
rect 1339 1071 1340 1075
rect 1340 1071 1343 1075
rect 1383 1068 1387 1072
rect 1415 1068 1419 1072
rect 1427 1067 1428 1071
rect 1428 1067 1431 1071
rect 1447 1071 1451 1075
rect 111 1053 115 1057
rect 135 1056 139 1060
rect 159 1056 163 1060
rect 183 1056 187 1060
rect 207 1056 211 1060
rect 231 1056 235 1060
rect 271 1056 275 1060
rect 311 1056 315 1060
rect 351 1056 355 1060
rect 391 1056 395 1060
rect 431 1056 435 1060
rect 471 1056 475 1060
rect 511 1056 515 1060
rect 551 1056 555 1060
rect 591 1056 595 1060
rect 631 1056 635 1060
rect 671 1056 675 1060
rect 711 1056 715 1060
rect 743 1056 747 1060
rect 783 1056 787 1060
rect 823 1056 827 1060
rect 871 1056 875 1060
rect 919 1056 923 1060
rect 975 1056 979 1060
rect 1011 1055 1015 1059
rect 1031 1056 1035 1060
rect 1079 1056 1083 1060
rect 1127 1056 1131 1060
rect 1175 1056 1179 1060
rect 1223 1056 1227 1060
rect 1271 1056 1275 1060
rect 1327 1056 1331 1060
rect 1383 1056 1387 1060
rect 1415 1056 1419 1060
rect 1447 1053 1451 1057
rect 171 1047 175 1051
rect 111 1035 115 1039
rect 195 1047 199 1051
rect 219 1047 223 1051
rect 243 1047 247 1051
rect 323 1047 327 1051
rect 619 1047 623 1051
rect 775 1047 779 1051
rect 883 1047 887 1051
rect 1235 1047 1239 1051
rect 1339 1047 1343 1051
rect 135 1030 139 1034
rect 147 1031 148 1035
rect 148 1031 151 1035
rect 159 1030 163 1034
rect 171 1031 172 1035
rect 172 1031 175 1035
rect 183 1030 187 1034
rect 195 1031 196 1035
rect 196 1031 199 1035
rect 207 1030 211 1034
rect 219 1031 220 1035
rect 220 1031 223 1035
rect 231 1030 235 1034
rect 243 1031 244 1035
rect 244 1031 247 1035
rect 271 1030 275 1034
rect 311 1030 315 1034
rect 323 1031 324 1035
rect 324 1031 327 1035
rect 351 1030 355 1034
rect 391 1030 395 1034
rect 431 1030 435 1034
rect 471 1030 475 1034
rect 511 1030 515 1034
rect 551 1030 555 1034
rect 591 1030 595 1034
rect 539 1023 543 1027
rect 603 1027 604 1031
rect 604 1027 607 1031
rect 631 1030 635 1034
rect 671 1030 675 1034
rect 711 1030 715 1034
rect 743 1030 747 1034
rect 783 1030 787 1034
rect 795 1031 796 1035
rect 796 1031 799 1035
rect 823 1030 827 1034
rect 835 1027 836 1031
rect 836 1027 839 1031
rect 871 1030 875 1034
rect 883 1031 884 1035
rect 884 1031 887 1035
rect 1003 1039 1007 1043
rect 919 1030 923 1034
rect 975 1030 979 1034
rect 1031 1030 1035 1034
rect 1079 1030 1083 1034
rect 1127 1030 1131 1034
rect 1139 1031 1140 1035
rect 1140 1031 1143 1035
rect 1175 1030 1179 1034
rect 1187 1027 1188 1031
rect 1188 1027 1191 1031
rect 1223 1030 1227 1034
rect 1235 1031 1236 1035
rect 1236 1031 1239 1035
rect 1263 1039 1267 1043
rect 1395 1039 1396 1043
rect 1396 1039 1399 1043
rect 1271 1030 1275 1034
rect 1327 1030 1331 1034
rect 1339 1031 1340 1035
rect 1340 1031 1343 1035
rect 1383 1030 1387 1034
rect 1415 1030 1419 1034
rect 1427 1031 1428 1035
rect 1428 1031 1431 1035
rect 1447 1035 1451 1039
rect 775 1019 779 1023
rect 159 1014 163 1018
rect 183 1014 187 1018
rect 111 1009 115 1013
rect 207 1014 211 1018
rect 231 1014 235 1018
rect 263 1014 267 1018
rect 303 1014 307 1018
rect 343 1014 347 1018
rect 383 1014 387 1018
rect 411 1011 415 1015
rect 431 1014 435 1018
rect 479 1014 483 1018
rect 527 1014 531 1018
rect 575 1014 579 1018
rect 623 1014 627 1018
rect 671 1014 675 1018
rect 603 1003 607 1007
rect 719 1014 723 1018
rect 767 1014 771 1018
rect 823 1014 827 1018
rect 879 1014 883 1018
rect 835 1003 836 1007
rect 836 1003 839 1007
rect 935 1014 939 1018
rect 991 1014 995 1018
rect 1003 1015 1004 1019
rect 1004 1015 1007 1019
rect 1047 1014 1051 1018
rect 1103 1014 1107 1018
rect 1159 1014 1163 1018
rect 1215 1014 1219 1018
rect 111 991 115 995
rect 159 988 163 992
rect 183 988 187 992
rect 207 988 211 992
rect 231 988 235 992
rect 263 988 267 992
rect 303 988 307 992
rect 343 988 347 992
rect 355 991 356 995
rect 356 991 359 995
rect 383 988 387 992
rect 431 988 435 992
rect 479 988 483 992
rect 527 988 531 992
rect 539 991 540 995
rect 540 991 543 995
rect 575 988 579 992
rect 623 988 627 992
rect 663 987 667 991
rect 671 988 675 992
rect 719 988 723 992
rect 767 988 771 992
rect 823 988 827 992
rect 899 1003 903 1007
rect 1187 1003 1191 1007
rect 1271 1014 1275 1018
rect 1327 1014 1331 1018
rect 1347 1011 1351 1015
rect 1383 1014 1387 1018
rect 1395 1015 1396 1019
rect 1396 1015 1399 1019
rect 1415 1014 1419 1018
rect 1447 1009 1451 1013
rect 879 988 883 992
rect 935 988 939 992
rect 991 988 995 992
rect 1047 988 1051 992
rect 1103 988 1107 992
rect 1115 987 1116 991
rect 1116 987 1119 991
rect 1159 988 1163 992
rect 1215 988 1219 992
rect 1271 988 1275 992
rect 1327 988 1331 992
rect 1383 988 1387 992
rect 1415 988 1419 992
rect 1427 987 1428 991
rect 1428 987 1431 991
rect 1447 991 1451 995
rect 111 973 115 977
rect 207 976 211 980
rect 231 976 235 980
rect 255 976 259 980
rect 287 976 291 980
rect 327 976 331 980
rect 375 976 379 980
rect 423 976 427 980
rect 471 976 475 980
rect 519 976 523 980
rect 567 976 571 980
rect 623 976 627 980
rect 679 976 683 980
rect 727 976 731 980
rect 775 976 779 980
rect 831 976 835 980
rect 887 976 891 980
rect 899 975 900 979
rect 900 975 903 979
rect 943 976 947 980
rect 999 976 1003 980
rect 1047 976 1051 980
rect 1095 976 1099 980
rect 1143 976 1147 980
rect 1191 976 1195 980
rect 1239 976 1243 980
rect 1287 976 1291 980
rect 1335 976 1339 980
rect 1383 976 1387 980
rect 1415 976 1419 980
rect 1447 973 1451 977
rect 243 967 247 971
rect 111 955 115 959
rect 267 967 271 971
rect 339 967 343 971
rect 411 967 415 971
rect 739 967 743 971
rect 843 967 847 971
rect 1347 967 1351 971
rect 207 950 211 954
rect 219 951 220 955
rect 220 951 223 955
rect 231 950 235 954
rect 243 951 244 955
rect 244 951 247 955
rect 255 950 259 954
rect 267 951 268 955
rect 268 951 271 955
rect 287 950 291 954
rect 327 950 331 954
rect 339 951 340 955
rect 340 951 343 955
rect 275 943 279 947
rect 303 943 307 947
rect 375 950 379 954
rect 423 950 427 954
rect 471 950 475 954
rect 519 950 523 954
rect 531 947 532 951
rect 532 947 535 951
rect 567 950 571 954
rect 623 950 627 954
rect 679 950 683 954
rect 931 959 935 963
rect 727 950 731 954
rect 663 943 667 947
rect 775 950 779 954
rect 795 947 799 951
rect 831 950 835 954
rect 843 951 844 955
rect 844 951 847 955
rect 887 950 891 954
rect 943 950 947 954
rect 999 950 1003 954
rect 1047 950 1051 954
rect 1095 950 1099 954
rect 1115 951 1119 955
rect 1143 950 1147 954
rect 1191 950 1195 954
rect 1239 950 1243 954
rect 1287 950 1291 954
rect 1335 950 1339 954
rect 1383 950 1387 954
rect 1131 943 1135 947
rect 1415 950 1419 954
rect 1427 951 1428 955
rect 1428 951 1431 955
rect 1447 955 1451 959
rect 215 934 219 938
rect 111 929 115 933
rect 227 931 228 935
rect 228 931 231 935
rect 239 934 243 938
rect 263 934 267 938
rect 287 934 291 938
rect 319 934 323 938
rect 351 934 355 938
rect 391 934 395 938
rect 431 934 435 938
rect 471 934 475 938
rect 111 911 115 915
rect 443 923 444 927
rect 444 923 447 927
rect 507 931 511 935
rect 519 934 523 938
rect 539 931 543 935
rect 567 934 571 938
rect 615 934 619 938
rect 531 923 532 927
rect 532 923 535 927
rect 671 934 675 938
rect 727 934 731 938
rect 739 935 740 939
rect 740 935 743 939
rect 783 934 787 938
rect 847 934 851 938
rect 795 923 796 927
rect 796 923 799 927
rect 859 931 860 935
rect 860 931 863 935
rect 919 934 923 938
rect 931 935 932 939
rect 932 935 935 939
rect 991 934 995 938
rect 1003 931 1004 935
rect 1004 931 1007 935
rect 1055 934 1059 938
rect 1119 934 1123 938
rect 1175 934 1179 938
rect 215 908 219 912
rect 239 908 243 912
rect 263 908 267 912
rect 275 911 276 915
rect 276 911 279 915
rect 287 908 291 912
rect 319 908 323 912
rect 351 908 355 912
rect 991 919 995 923
rect 1131 923 1132 927
rect 1132 923 1135 927
rect 1223 934 1227 938
rect 1263 934 1267 938
rect 1295 934 1299 938
rect 1327 934 1331 938
rect 1359 934 1363 938
rect 1391 934 1395 938
rect 1415 934 1419 938
rect 1447 929 1451 933
rect 391 908 395 912
rect 403 907 404 911
rect 404 907 407 911
rect 431 908 435 912
rect 471 908 475 912
rect 519 908 523 912
rect 567 908 571 912
rect 607 907 611 911
rect 615 908 619 912
rect 671 908 675 912
rect 727 908 731 912
rect 783 908 787 912
rect 847 908 851 912
rect 919 908 923 912
rect 991 908 995 912
rect 1055 908 1059 912
rect 1067 907 1068 911
rect 1068 907 1071 911
rect 1119 908 1123 912
rect 1175 908 1179 912
rect 1223 908 1227 912
rect 1263 908 1267 912
rect 1295 908 1299 912
rect 1327 908 1331 912
rect 1359 908 1363 912
rect 1391 908 1395 912
rect 1403 907 1404 911
rect 1404 907 1407 911
rect 1415 908 1419 912
rect 1447 911 1451 915
rect 111 893 115 897
rect 231 896 235 900
rect 255 896 259 900
rect 279 896 283 900
rect 303 896 307 900
rect 327 896 331 900
rect 359 896 363 900
rect 391 896 395 900
rect 423 896 427 900
rect 455 896 459 900
rect 495 896 499 900
rect 507 895 508 899
rect 508 895 511 899
rect 535 896 539 900
rect 575 896 579 900
rect 623 896 627 900
rect 663 896 667 900
rect 703 896 707 900
rect 751 896 755 900
rect 807 896 811 900
rect 855 895 859 899
rect 863 896 867 900
rect 927 896 931 900
rect 991 896 995 900
rect 1055 896 1059 900
rect 1119 896 1123 900
rect 1175 896 1179 900
rect 1231 896 1235 900
rect 1279 896 1283 900
rect 1327 896 1331 900
rect 1383 896 1387 900
rect 1415 896 1419 900
rect 1447 893 1451 897
rect 239 883 240 887
rect 240 883 243 887
rect 467 887 471 891
rect 763 887 767 891
rect 1187 887 1191 891
rect 1291 887 1295 891
rect 111 875 115 879
rect 231 870 235 874
rect 255 870 259 874
rect 279 870 283 874
rect 303 870 307 874
rect 327 870 331 874
rect 359 870 363 874
rect 391 870 395 874
rect 403 871 404 875
rect 404 871 407 875
rect 423 870 427 874
rect 239 863 243 867
rect 399 863 403 867
rect 455 870 459 874
rect 467 871 468 875
rect 468 871 471 875
rect 495 870 499 874
rect 535 870 539 874
rect 575 870 579 874
rect 623 870 627 874
rect 663 870 667 874
rect 607 863 611 867
rect 703 870 707 874
rect 751 870 755 874
rect 763 871 764 875
rect 764 871 767 875
rect 807 870 811 874
rect 863 870 867 874
rect 927 870 931 874
rect 991 870 995 874
rect 1055 870 1059 874
rect 1067 871 1068 875
rect 1068 871 1071 875
rect 1119 870 1123 874
rect 779 863 783 867
rect 1175 870 1179 874
rect 1187 871 1188 875
rect 1188 871 1191 875
rect 1199 871 1203 875
rect 1231 870 1235 874
rect 1279 870 1283 874
rect 1291 871 1292 875
rect 1292 871 1295 875
rect 207 854 211 858
rect 111 849 115 853
rect 231 854 235 858
rect 255 854 259 858
rect 287 854 291 858
rect 319 854 323 858
rect 351 854 355 858
rect 383 854 387 858
rect 415 854 419 858
rect 392 843 396 847
rect 447 854 451 858
rect 479 854 483 858
rect 499 851 503 855
rect 511 854 515 858
rect 551 854 555 858
rect 599 854 603 858
rect 647 854 651 858
rect 703 854 707 858
rect 767 854 771 858
rect 839 854 843 858
rect 911 854 915 858
rect 667 843 671 847
rect 983 854 987 858
rect 1047 854 1051 858
rect 1103 854 1107 858
rect 1151 855 1155 859
rect 1159 854 1163 858
rect 1183 863 1187 867
rect 1303 863 1307 867
rect 1427 879 1428 883
rect 1428 879 1431 883
rect 1447 875 1451 879
rect 1327 870 1331 874
rect 1383 870 1387 874
rect 1415 870 1419 874
rect 1403 863 1407 867
rect 1199 855 1203 859
rect 1207 854 1211 858
rect 1247 854 1251 858
rect 1295 854 1299 858
rect 1343 854 1347 858
rect 1391 854 1395 858
rect 1415 854 1419 858
rect 1427 855 1428 859
rect 1428 855 1431 859
rect 1447 849 1451 853
rect 111 831 115 835
rect 207 828 211 832
rect 231 828 235 832
rect 255 828 259 832
rect 287 828 291 832
rect 319 828 323 832
rect 351 828 355 832
rect 383 828 387 832
rect 415 828 419 832
rect 447 828 451 832
rect 479 828 483 832
rect 511 828 515 832
rect 535 827 539 831
rect 551 828 555 832
rect 599 828 603 832
rect 647 828 651 832
rect 703 828 707 832
rect 767 828 771 832
rect 779 831 780 835
rect 780 831 783 835
rect 839 828 843 832
rect 851 827 852 831
rect 852 827 855 831
rect 911 828 915 832
rect 983 828 987 832
rect 1047 828 1051 832
rect 1103 828 1107 832
rect 1159 828 1163 832
rect 1183 831 1187 835
rect 1207 828 1211 832
rect 1247 828 1251 832
rect 1295 828 1299 832
rect 1343 828 1347 832
rect 1391 828 1395 832
rect 1403 827 1404 831
rect 1404 827 1407 831
rect 1415 828 1419 832
rect 1447 831 1451 835
rect 111 813 115 817
rect 135 816 139 820
rect 159 816 163 820
rect 183 816 187 820
rect 215 816 219 820
rect 1303 823 1307 827
rect 263 816 267 820
rect 311 816 315 820
rect 367 816 371 820
rect 431 816 435 820
rect 487 816 491 820
rect 543 816 547 820
rect 599 816 603 820
rect 655 816 659 820
rect 667 815 668 819
rect 668 815 671 819
rect 711 816 715 820
rect 767 816 771 820
rect 815 816 819 820
rect 863 816 867 820
rect 903 816 907 820
rect 935 816 939 820
rect 967 816 971 820
rect 991 816 995 820
rect 1015 816 1019 820
rect 1039 816 1043 820
rect 1063 816 1067 820
rect 1095 816 1099 820
rect 1127 816 1131 820
rect 1167 816 1171 820
rect 1207 816 1211 820
rect 1255 816 1259 820
rect 1311 816 1315 820
rect 1375 816 1379 820
rect 1415 816 1419 820
rect 1447 813 1451 817
rect 419 807 423 811
rect 499 807 503 811
rect 611 807 615 811
rect 779 807 783 811
rect 947 807 951 811
rect 1003 807 1007 811
rect 1051 807 1055 811
rect 111 795 115 799
rect 135 790 139 794
rect 159 790 163 794
rect 183 790 187 794
rect 215 790 219 794
rect 263 790 267 794
rect 311 790 315 794
rect 367 790 371 794
rect 431 790 435 794
rect 487 790 491 794
rect 807 799 811 803
rect 1075 807 1079 811
rect 1103 803 1104 807
rect 1104 803 1107 807
rect 1179 807 1183 811
rect 1267 807 1271 811
rect 1275 807 1279 811
rect 543 790 547 794
rect 535 783 539 787
rect 599 790 603 794
rect 611 791 612 795
rect 612 791 615 795
rect 655 790 659 794
rect 711 790 715 794
rect 731 787 735 791
rect 767 790 771 794
rect 779 791 780 795
rect 780 791 783 795
rect 815 790 819 794
rect 851 791 855 795
rect 863 790 867 794
rect 903 790 907 794
rect 935 790 939 794
rect 947 791 948 795
rect 948 791 951 795
rect 967 790 971 794
rect 991 790 995 794
rect 1003 791 1004 795
rect 1004 791 1007 795
rect 1015 790 1019 794
rect 807 779 811 783
rect 135 774 139 778
rect 111 769 115 773
rect 159 774 163 778
rect 183 774 187 778
rect 223 774 227 778
rect 279 774 283 778
rect 343 774 347 778
rect 407 774 411 778
rect 419 775 420 779
rect 420 775 423 779
rect 463 774 467 778
rect 511 771 515 775
rect 519 774 523 778
rect 575 774 579 778
rect 623 774 627 778
rect 635 771 636 775
rect 636 771 639 775
rect 671 774 675 778
rect 719 774 723 778
rect 759 774 763 778
rect 799 774 803 778
rect 839 774 843 778
rect 111 751 115 755
rect 623 759 627 763
rect 731 763 732 767
rect 732 763 735 767
rect 863 771 867 775
rect 879 774 883 778
rect 919 774 923 778
rect 951 783 955 787
rect 1039 790 1043 794
rect 1051 791 1052 795
rect 1052 791 1055 795
rect 1063 790 1067 794
rect 1075 791 1076 795
rect 1076 791 1079 795
rect 1095 790 1099 794
rect 1127 790 1131 794
rect 1159 791 1163 795
rect 1167 790 1171 794
rect 1179 791 1180 795
rect 1180 791 1183 795
rect 1207 790 1211 794
rect 1255 790 1259 794
rect 1267 791 1268 795
rect 1268 791 1271 795
rect 1151 779 1155 783
rect 1275 783 1279 787
rect 1427 799 1428 803
rect 1428 799 1431 803
rect 1311 790 1315 794
rect 1375 790 1379 794
rect 1447 795 1451 799
rect 1403 791 1407 795
rect 1415 790 1419 794
rect 959 774 963 778
rect 991 774 995 778
rect 1003 771 1004 775
rect 1004 771 1007 775
rect 1023 774 1027 778
rect 1055 774 1059 778
rect 1087 774 1091 778
rect 1127 774 1131 778
rect 1175 774 1179 778
rect 1231 774 1235 778
rect 1295 774 1299 778
rect 1367 774 1371 778
rect 1415 774 1419 778
rect 1427 775 1428 779
rect 1428 775 1431 779
rect 1447 769 1451 773
rect 135 748 139 752
rect 147 747 148 751
rect 148 747 151 751
rect 159 748 163 752
rect 183 748 187 752
rect 223 748 227 752
rect 279 748 283 752
rect 343 748 347 752
rect 407 748 411 752
rect 463 748 467 752
rect 519 748 523 752
rect 575 748 579 752
rect 623 748 627 752
rect 671 748 675 752
rect 127 739 131 743
rect 111 729 115 733
rect 135 732 139 736
rect 159 732 163 736
rect 183 732 187 736
rect 215 732 219 736
rect 263 732 267 736
rect 319 732 323 736
rect 511 739 515 743
rect 719 748 723 752
rect 759 748 763 752
rect 771 747 772 751
rect 772 747 775 751
rect 799 748 803 752
rect 839 748 843 752
rect 879 748 883 752
rect 919 748 923 752
rect 951 751 955 755
rect 959 748 963 752
rect 991 748 995 752
rect 1023 748 1027 752
rect 1055 748 1059 752
rect 1087 748 1091 752
rect 1127 748 1131 752
rect 1175 748 1179 752
rect 1231 748 1235 752
rect 1295 748 1299 752
rect 1367 748 1371 752
rect 1415 748 1419 752
rect 1447 751 1451 755
rect 375 732 379 736
rect 423 732 427 736
rect 471 732 475 736
rect 519 732 523 736
rect 567 732 571 736
rect 615 732 619 736
rect 863 739 867 743
rect 1003 739 1007 743
rect 1103 739 1107 743
rect 1159 739 1163 743
rect 1375 743 1379 747
rect 663 732 667 736
rect 703 732 707 736
rect 751 732 755 736
rect 807 732 811 736
rect 871 732 875 736
rect 943 732 947 736
rect 1015 732 1019 736
rect 1087 732 1091 736
rect 1151 732 1155 736
rect 1215 732 1219 736
rect 1271 732 1275 736
rect 1327 732 1331 736
rect 1383 732 1387 736
rect 1415 732 1419 736
rect 1447 729 1451 733
rect 171 723 175 727
rect 227 723 231 727
rect 331 723 335 727
rect 483 723 487 727
rect 579 723 583 727
rect 675 723 679 727
rect 883 723 887 727
rect 1027 723 1031 727
rect 1051 723 1055 727
rect 1291 723 1295 727
rect 111 711 115 715
rect 135 706 139 710
rect 147 707 148 711
rect 148 707 151 711
rect 159 706 163 710
rect 171 707 172 711
rect 172 707 175 711
rect 183 706 187 710
rect 127 699 131 703
rect 215 706 219 710
rect 227 707 228 711
rect 228 707 231 711
rect 263 706 267 710
rect 319 706 323 710
rect 331 707 332 711
rect 332 707 335 711
rect 375 706 379 710
rect 423 706 427 710
rect 471 706 475 710
rect 483 707 484 711
rect 484 707 487 711
rect 495 699 499 703
rect 519 706 523 710
rect 567 706 571 710
rect 579 707 580 711
rect 580 707 583 711
rect 615 706 619 710
rect 663 706 667 710
rect 675 707 676 711
rect 676 707 679 711
rect 703 706 707 710
rect 751 706 755 710
rect 771 707 775 711
rect 807 706 811 710
rect 839 703 843 707
rect 871 706 875 710
rect 883 707 884 711
rect 884 707 887 711
rect 847 699 851 703
rect 943 706 947 710
rect 1015 706 1019 710
rect 1027 707 1028 711
rect 1028 707 1031 711
rect 1051 699 1055 703
rect 1087 706 1091 710
rect 1151 706 1155 710
rect 1215 706 1219 710
rect 1427 715 1428 719
rect 1428 715 1431 719
rect 1271 706 1275 710
rect 1327 706 1331 710
rect 1375 707 1379 711
rect 1383 706 1387 710
rect 1447 711 1451 715
rect 1415 706 1419 710
rect 135 690 139 694
rect 159 690 163 694
rect 111 685 115 689
rect 199 690 203 694
rect 239 690 243 694
rect 287 690 291 694
rect 335 690 339 694
rect 391 690 395 694
rect 431 687 435 691
rect 439 690 443 694
rect 451 687 452 691
rect 452 687 455 691
rect 487 690 491 694
rect 535 690 539 694
rect 583 690 587 694
rect 639 690 643 694
rect 695 690 699 694
rect 111 667 115 671
rect 135 664 139 668
rect 159 664 163 668
rect 199 664 203 668
rect 239 664 243 668
rect 287 664 291 668
rect 439 679 443 683
rect 759 690 763 694
rect 831 690 835 694
rect 335 664 339 668
rect 347 663 348 667
rect 348 663 351 667
rect 391 664 395 668
rect 439 664 443 668
rect 487 664 491 668
rect 535 664 539 668
rect 903 690 907 694
rect 839 679 840 683
rect 840 679 843 683
rect 967 690 971 694
rect 1031 690 1035 694
rect 1087 690 1091 694
rect 1135 690 1139 694
rect 1175 690 1179 694
rect 1215 690 1219 694
rect 1247 690 1251 694
rect 1279 690 1283 694
rect 1291 691 1292 695
rect 1292 691 1295 695
rect 1311 690 1315 694
rect 1343 690 1347 694
rect 1355 687 1356 691
rect 1356 687 1359 691
rect 1367 690 1371 694
rect 1391 690 1395 694
rect 1415 690 1419 694
rect 1427 691 1428 695
rect 1428 691 1431 695
rect 1447 685 1451 689
rect 583 664 587 668
rect 639 664 643 668
rect 651 663 652 667
rect 652 663 655 667
rect 695 664 699 668
rect 759 664 763 668
rect 831 664 835 668
rect 903 664 907 668
rect 967 664 971 668
rect 1031 664 1035 668
rect 111 649 115 653
rect 191 652 195 656
rect 215 652 219 656
rect 239 652 243 656
rect 263 652 267 656
rect 295 652 299 656
rect 327 652 331 656
rect 367 652 371 656
rect 407 652 411 656
rect 431 655 435 659
rect 455 652 459 656
rect 227 643 231 647
rect 275 643 279 647
rect 339 643 343 647
rect 467 643 471 647
rect 495 659 499 663
rect 1079 663 1083 667
rect 1087 664 1091 668
rect 1135 664 1139 668
rect 1175 664 1179 668
rect 1215 664 1219 668
rect 1247 664 1251 668
rect 1279 664 1283 668
rect 1311 664 1315 668
rect 1343 664 1347 668
rect 1367 664 1371 668
rect 1391 664 1395 668
rect 1415 664 1419 668
rect 1447 667 1451 671
rect 503 652 507 656
rect 551 652 555 656
rect 607 652 611 656
rect 663 652 667 656
rect 719 652 723 656
rect 767 652 771 656
rect 815 652 819 656
rect 847 651 851 655
rect 863 652 867 656
rect 903 652 907 656
rect 935 652 939 656
rect 967 652 971 656
rect 1007 652 1011 656
rect 1047 652 1051 656
rect 1087 652 1091 656
rect 1127 652 1131 656
rect 1159 652 1163 656
rect 1191 652 1195 656
rect 1223 652 1227 656
rect 1263 652 1267 656
rect 1303 652 1307 656
rect 1343 652 1347 656
rect 1355 655 1359 659
rect 1447 649 1451 653
rect 563 643 567 647
rect 675 643 679 647
rect 987 643 991 647
rect 1079 643 1083 647
rect 1171 643 1175 647
rect 1235 643 1239 647
rect 1315 643 1319 647
rect 1323 643 1327 647
rect 111 631 115 635
rect 191 626 195 630
rect 203 627 204 631
rect 204 627 207 631
rect 215 626 219 630
rect 227 627 228 631
rect 228 627 231 631
rect 239 626 243 630
rect 263 626 267 630
rect 275 627 276 631
rect 276 627 279 631
rect 295 626 299 630
rect 327 626 331 630
rect 339 627 340 631
rect 340 627 343 631
rect 367 626 371 630
rect 407 626 411 630
rect 447 627 451 631
rect 455 626 459 630
rect 467 627 468 631
rect 468 627 471 631
rect 503 626 507 630
rect 551 626 555 630
rect 563 627 564 631
rect 564 627 567 631
rect 607 626 611 630
rect 651 627 655 631
rect 663 626 667 630
rect 675 627 676 631
rect 676 627 679 631
rect 711 635 715 639
rect 719 626 723 630
rect 767 626 771 630
rect 815 626 819 630
rect 863 626 867 630
rect 903 626 907 630
rect 935 626 939 630
rect 967 626 971 630
rect 1007 626 1011 630
rect 1047 626 1051 630
rect 1087 626 1091 630
rect 1127 626 1131 630
rect 423 615 427 619
rect 271 610 275 614
rect 295 610 299 614
rect 111 605 115 609
rect 307 607 308 611
rect 308 607 311 611
rect 319 610 323 614
rect 343 610 347 614
rect 367 610 371 614
rect 391 610 395 614
rect 403 607 404 611
rect 404 607 407 611
rect 415 610 419 614
rect 295 599 299 603
rect 391 595 395 599
rect 415 595 419 599
rect 111 587 115 591
rect 271 584 275 588
rect 295 584 299 588
rect 319 584 323 588
rect 343 584 347 588
rect 367 584 371 588
rect 391 584 395 588
rect 415 584 419 588
rect 775 619 779 623
rect 1035 619 1039 623
rect 1159 626 1163 630
rect 1171 627 1172 631
rect 1172 627 1175 631
rect 1191 626 1195 630
rect 1223 626 1227 630
rect 1235 627 1236 631
rect 1236 627 1239 631
rect 1263 626 1267 630
rect 1303 626 1307 630
rect 1315 627 1316 631
rect 1316 627 1319 631
rect 439 610 443 614
rect 479 610 483 614
rect 519 610 523 614
rect 567 610 571 614
rect 623 610 627 614
rect 679 610 683 614
rect 711 611 715 615
rect 735 610 739 614
rect 783 610 787 614
rect 795 607 796 611
rect 796 607 799 611
rect 831 610 835 614
rect 879 610 883 614
rect 927 610 931 614
rect 775 599 779 603
rect 439 584 443 588
rect 479 584 483 588
rect 975 610 979 614
rect 987 611 988 615
rect 988 611 991 615
rect 1023 610 1027 614
rect 1071 610 1075 614
rect 1035 599 1036 603
rect 1036 599 1039 603
rect 1111 610 1115 614
rect 1151 610 1155 614
rect 1191 610 1195 614
rect 1323 619 1327 623
rect 1447 631 1451 635
rect 1343 626 1347 630
rect 1239 610 1243 614
rect 1287 610 1291 614
rect 1335 610 1339 614
rect 1447 605 1451 609
rect 519 584 523 588
rect 531 587 532 591
rect 532 587 535 591
rect 567 584 571 588
rect 615 583 619 587
rect 623 584 627 588
rect 679 584 683 588
rect 735 584 739 588
rect 783 584 787 588
rect 831 584 835 588
rect 871 583 875 587
rect 879 584 883 588
rect 927 584 931 588
rect 975 584 979 588
rect 1023 584 1027 588
rect 1071 584 1075 588
rect 1111 584 1115 588
rect 1151 584 1155 588
rect 1191 584 1195 588
rect 1239 584 1243 588
rect 1287 584 1291 588
rect 1335 584 1339 588
rect 1387 583 1391 587
rect 1447 587 1451 591
rect 111 569 115 573
rect 263 572 267 576
rect 287 572 291 576
rect 311 572 315 576
rect 335 572 339 576
rect 359 572 363 576
rect 383 572 387 576
rect 407 572 411 576
rect 431 572 435 576
rect 463 572 467 576
rect 503 572 507 576
rect 551 572 555 576
rect 607 572 611 576
rect 663 572 667 576
rect 719 572 723 576
rect 775 572 779 576
rect 399 563 403 567
rect 440 567 444 571
rect 795 571 799 575
rect 831 572 835 576
rect 887 572 891 576
rect 943 572 947 576
rect 1007 572 1011 576
rect 1071 572 1075 576
rect 1127 572 1131 576
rect 1183 572 1187 576
rect 1247 572 1251 576
rect 1311 572 1315 576
rect 1375 572 1379 576
rect 1447 569 1451 573
rect 111 551 115 555
rect 263 546 267 550
rect 287 546 291 550
rect 311 546 315 550
rect 335 546 339 550
rect 359 546 363 550
rect 383 546 387 550
rect 407 546 411 550
rect 416 547 420 551
rect 431 546 435 550
rect 463 546 467 550
rect 675 563 679 567
rect 1035 563 1039 567
rect 1139 563 1143 567
rect 539 555 543 559
rect 503 546 507 550
rect 515 543 516 547
rect 516 543 519 547
rect 551 546 555 550
rect 607 546 611 550
rect 619 547 620 551
rect 620 547 623 551
rect 663 546 667 550
rect 675 547 676 551
rect 676 547 679 551
rect 719 546 723 550
rect 399 535 403 539
rect 587 539 591 543
rect 731 543 732 547
rect 732 543 735 547
rect 775 546 779 550
rect 831 546 835 550
rect 887 546 891 550
rect 943 546 947 550
rect 1007 546 1011 550
rect 871 539 875 543
rect 1071 546 1075 550
rect 1091 543 1095 547
rect 1127 546 1131 550
rect 1139 547 1140 551
rect 1140 547 1143 551
rect 1283 555 1287 559
rect 1183 546 1187 550
rect 1247 546 1251 550
rect 1311 546 1315 550
rect 1375 546 1379 550
rect 1387 547 1388 551
rect 1388 547 1391 551
rect 1447 551 1451 555
rect 1363 539 1367 543
rect 223 530 227 534
rect 111 525 115 529
rect 235 527 236 531
rect 236 527 239 531
rect 247 530 251 534
rect 271 530 275 534
rect 295 530 299 534
rect 327 530 331 534
rect 359 530 363 534
rect 391 530 395 534
rect 423 530 427 534
rect 447 527 451 531
rect 455 530 459 534
rect 467 527 468 531
rect 468 527 471 531
rect 487 530 491 534
rect 499 527 500 531
rect 500 527 503 531
rect 527 530 531 534
rect 539 531 540 535
rect 540 531 543 535
rect 575 530 579 534
rect 623 530 627 534
rect 671 530 675 534
rect 711 530 715 534
rect 759 530 763 534
rect 455 519 459 523
rect 487 519 491 523
rect 515 519 519 523
rect 111 507 115 511
rect 587 511 588 515
rect 588 511 591 515
rect 731 519 735 523
rect 807 530 811 534
rect 855 530 859 534
rect 911 530 915 534
rect 967 530 971 534
rect 1023 530 1027 534
rect 1035 531 1036 535
rect 1036 531 1039 535
rect 1079 530 1083 534
rect 1127 530 1131 534
rect 1091 519 1092 523
rect 1092 519 1095 523
rect 1175 530 1179 534
rect 1223 530 1227 534
rect 1263 527 1267 531
rect 1271 530 1275 534
rect 1283 531 1284 535
rect 1284 531 1287 535
rect 1311 530 1315 534
rect 1351 530 1355 534
rect 1391 530 1395 534
rect 1415 530 1419 534
rect 1447 525 1451 529
rect 223 504 227 508
rect 247 504 251 508
rect 271 504 275 508
rect 295 504 299 508
rect 327 504 331 508
rect 359 504 363 508
rect 391 504 395 508
rect 423 504 427 508
rect 455 504 459 508
rect 487 504 491 508
rect 527 504 531 508
rect 575 504 579 508
rect 623 504 627 508
rect 671 504 675 508
rect 711 504 715 508
rect 759 504 763 508
rect 807 504 811 508
rect 855 504 859 508
rect 911 504 915 508
rect 967 504 971 508
rect 1023 504 1027 508
rect 1079 504 1083 508
rect 1127 504 1131 508
rect 1175 504 1179 508
rect 1223 504 1227 508
rect 1271 504 1275 508
rect 1311 504 1315 508
rect 1351 504 1355 508
rect 1363 507 1364 511
rect 1364 507 1367 511
rect 1391 504 1395 508
rect 1415 504 1419 508
rect 1427 503 1428 507
rect 1428 503 1431 507
rect 1447 507 1451 511
rect 231 499 235 503
rect 111 489 115 493
rect 135 492 139 496
rect 159 492 163 496
rect 183 492 187 496
rect 223 492 227 496
rect 239 495 243 499
rect 679 499 683 503
rect 271 492 275 496
rect 319 492 323 496
rect 375 492 379 496
rect 431 492 435 496
rect 487 492 491 496
rect 543 492 547 496
rect 591 492 595 496
rect 631 492 635 496
rect 663 492 667 496
rect 687 492 691 496
rect 719 492 723 496
rect 759 492 763 496
rect 799 492 803 496
rect 847 492 851 496
rect 903 492 907 496
rect 951 492 955 496
rect 999 492 1003 496
rect 1047 492 1051 496
rect 1095 492 1099 496
rect 1143 492 1147 496
rect 1199 492 1203 496
rect 1255 492 1259 496
rect 1311 492 1315 496
rect 1375 492 1379 496
rect 1415 492 1419 496
rect 1447 489 1451 493
rect 363 483 367 487
rect 499 483 503 487
rect 603 483 607 487
rect 111 471 115 475
rect 135 466 139 470
rect 159 466 163 470
rect 183 466 187 470
rect 223 466 227 470
rect 271 466 275 470
rect 319 466 323 470
rect 447 475 451 479
rect 679 475 683 479
rect 731 483 735 487
rect 811 483 815 487
rect 819 483 823 487
rect 895 483 899 487
rect 963 483 967 487
rect 1059 483 1063 487
rect 1155 483 1159 487
rect 1267 483 1271 487
rect 1279 483 1283 487
rect 375 466 379 470
rect 231 459 235 463
rect 431 466 435 470
rect 443 463 444 467
rect 444 463 447 467
rect 487 466 491 470
rect 499 467 500 471
rect 500 467 503 471
rect 543 466 547 470
rect 591 466 595 470
rect 603 467 604 471
rect 604 467 607 471
rect 631 466 635 470
rect 663 466 667 470
rect 655 459 659 463
rect 687 466 691 470
rect 719 466 723 470
rect 731 467 732 471
rect 732 467 735 471
rect 711 459 715 463
rect 759 466 763 470
rect 799 466 803 470
rect 811 467 812 471
rect 812 467 815 471
rect 919 475 923 479
rect 847 466 851 470
rect 903 466 907 470
rect 951 466 955 470
rect 963 467 964 471
rect 964 467 967 471
rect 999 466 1003 470
rect 923 459 927 463
rect 1047 466 1051 470
rect 1059 467 1060 471
rect 1060 467 1063 471
rect 1095 466 1099 470
rect 1143 466 1147 470
rect 1155 467 1156 471
rect 1156 467 1159 471
rect 1383 479 1384 483
rect 1384 479 1387 483
rect 1199 466 1203 470
rect 1255 466 1259 470
rect 1267 467 1268 471
rect 1268 467 1271 471
rect 1311 466 1315 470
rect 1375 466 1379 470
rect 1415 466 1419 470
rect 1427 467 1428 471
rect 1428 467 1431 471
rect 1447 471 1451 475
rect 135 450 139 454
rect 111 445 115 449
rect 159 450 163 454
rect 191 450 195 454
rect 127 435 131 439
rect 239 450 243 454
rect 295 450 299 454
rect 351 450 355 454
rect 363 451 364 455
rect 364 451 367 455
rect 415 450 419 454
rect 479 450 483 454
rect 443 439 447 443
rect 543 450 547 454
rect 607 450 611 454
rect 619 447 620 451
rect 620 447 623 451
rect 671 450 675 454
rect 683 447 684 451
rect 684 447 687 451
rect 735 450 739 454
rect 791 450 795 454
rect 819 451 823 455
rect 839 450 843 454
rect 851 447 852 451
rect 852 447 855 451
rect 879 450 883 454
rect 891 447 892 451
rect 892 447 895 451
rect 911 450 915 454
rect 943 450 947 454
rect 967 450 971 454
rect 999 450 1003 454
rect 1023 447 1027 451
rect 1031 450 1035 454
rect 1071 450 1075 454
rect 1119 450 1123 454
rect 1175 450 1179 454
rect 1239 450 1243 454
rect 1303 450 1307 454
rect 1331 447 1335 451
rect 1367 450 1371 454
rect 1376 447 1380 451
rect 1415 450 1419 454
rect 839 439 843 443
rect 879 439 883 443
rect 1447 445 1451 449
rect 111 427 115 431
rect 711 431 715 435
rect 923 431 924 435
rect 924 431 927 435
rect 135 424 139 428
rect 159 424 163 428
rect 191 424 195 428
rect 239 424 243 428
rect 295 424 299 428
rect 351 424 355 428
rect 415 424 419 428
rect 479 424 483 428
rect 543 424 547 428
rect 607 424 611 428
rect 671 424 675 428
rect 735 424 739 428
rect 791 424 795 428
rect 839 424 843 428
rect 879 424 883 428
rect 911 424 915 428
rect 943 424 947 428
rect 967 424 971 428
rect 987 423 991 427
rect 999 424 1003 428
rect 1031 424 1035 428
rect 1071 424 1075 428
rect 1119 424 1123 428
rect 1175 424 1179 428
rect 1239 424 1243 428
rect 1259 423 1263 427
rect 1303 424 1307 428
rect 1367 424 1371 428
rect 1415 424 1419 428
rect 1427 423 1428 427
rect 1428 423 1431 427
rect 1447 427 1451 431
rect 1311 419 1315 423
rect 111 409 115 413
rect 135 412 139 416
rect 159 412 163 416
rect 183 412 187 416
rect 215 412 219 416
rect 271 412 275 416
rect 327 412 331 416
rect 391 412 395 416
rect 447 412 451 416
rect 503 412 507 416
rect 551 412 555 416
rect 599 412 603 416
rect 647 412 651 416
rect 703 412 707 416
rect 767 412 771 416
rect 831 412 835 416
rect 903 412 907 416
rect 975 412 979 416
rect 1039 412 1043 416
rect 1103 412 1107 416
rect 1159 412 1163 416
rect 1207 412 1211 416
rect 1247 412 1251 416
rect 1279 412 1283 416
rect 1319 412 1323 416
rect 1331 411 1332 415
rect 1332 411 1335 415
rect 1359 412 1363 416
rect 1391 412 1395 416
rect 1415 412 1419 416
rect 1447 409 1451 413
rect 111 391 115 395
rect 135 386 139 390
rect 159 386 163 390
rect 183 386 187 390
rect 339 403 343 407
rect 347 403 351 407
rect 619 403 623 407
rect 1051 403 1055 407
rect 1239 403 1243 407
rect 215 386 219 390
rect 127 379 131 383
rect 271 386 275 390
rect 327 386 331 390
rect 339 387 340 391
rect 340 387 343 391
rect 391 386 395 390
rect 447 386 451 390
rect 503 386 507 390
rect 551 386 555 390
rect 599 386 603 390
rect 647 386 651 390
rect 739 395 743 399
rect 703 386 707 390
rect 715 383 716 387
rect 716 383 719 387
rect 767 386 771 390
rect 831 386 835 390
rect 1023 395 1027 399
rect 903 386 907 390
rect 347 375 351 379
rect 667 375 671 379
rect 975 386 979 390
rect 987 387 988 391
rect 988 387 991 391
rect 1039 386 1043 390
rect 1051 387 1052 391
rect 1052 387 1055 391
rect 1103 386 1107 390
rect 1159 386 1163 390
rect 1207 386 1211 390
rect 1247 386 1251 390
rect 1279 386 1283 390
rect 1311 387 1315 391
rect 1319 386 1323 390
rect 1359 386 1363 390
rect 1391 386 1395 390
rect 1259 379 1263 383
rect 1383 379 1387 383
rect 1415 386 1419 390
rect 1427 387 1428 391
rect 1428 387 1431 391
rect 1447 391 1451 395
rect 1239 371 1243 375
rect 135 366 139 370
rect 159 366 163 370
rect 111 361 115 365
rect 183 366 187 370
rect 207 366 211 370
rect 231 366 235 370
rect 255 366 259 370
rect 295 366 299 370
rect 335 366 339 370
rect 375 366 379 370
rect 415 366 419 370
rect 455 366 459 370
rect 495 366 499 370
rect 535 366 539 370
rect 575 366 579 370
rect 615 366 619 370
rect 627 363 628 367
rect 628 363 631 367
rect 655 366 659 370
rect 687 366 691 370
rect 667 355 668 359
rect 668 355 671 359
rect 727 366 731 370
rect 739 367 740 371
rect 740 367 743 371
rect 775 366 779 370
rect 831 366 835 370
rect 887 366 891 370
rect 951 366 955 370
rect 1015 366 1019 370
rect 1027 363 1028 367
rect 1028 363 1031 367
rect 1079 366 1083 370
rect 1135 366 1139 370
rect 1183 366 1187 370
rect 1231 366 1235 370
rect 1271 366 1275 370
rect 1291 363 1295 367
rect 1311 366 1315 370
rect 1351 366 1355 370
rect 1391 366 1395 370
rect 1415 366 1419 370
rect 1447 361 1451 365
rect 111 343 115 347
rect 135 340 139 344
rect 159 340 163 344
rect 183 340 187 344
rect 207 340 211 344
rect 231 340 235 344
rect 255 340 259 344
rect 295 340 299 344
rect 715 347 719 351
rect 1383 347 1387 351
rect 335 340 339 344
rect 347 339 348 343
rect 348 339 351 343
rect 375 340 379 344
rect 407 339 411 343
rect 415 340 419 344
rect 455 340 459 344
rect 495 340 499 344
rect 535 340 539 344
rect 575 340 579 344
rect 615 340 619 344
rect 655 340 659 344
rect 687 340 691 344
rect 727 340 731 344
rect 775 340 779 344
rect 831 340 835 344
rect 887 340 891 344
rect 951 340 955 344
rect 1015 340 1019 344
rect 1079 340 1083 344
rect 1135 340 1139 344
rect 1183 340 1187 344
rect 1231 340 1235 344
rect 1271 340 1275 344
rect 1311 340 1315 344
rect 1351 340 1355 344
rect 1391 340 1395 344
rect 1403 339 1404 343
rect 1404 339 1407 343
rect 1415 340 1419 344
rect 1447 343 1451 347
rect 111 325 115 329
rect 175 328 179 332
rect 199 328 203 332
rect 223 328 227 332
rect 247 328 251 332
rect 279 328 283 332
rect 319 328 323 332
rect 211 319 215 323
rect 259 319 263 323
rect 331 319 335 323
rect 359 328 363 332
rect 399 328 403 332
rect 439 328 443 332
rect 479 328 483 332
rect 527 328 531 332
rect 583 328 587 332
rect 639 328 643 332
rect 687 328 691 332
rect 735 328 739 332
rect 791 328 795 332
rect 847 328 851 332
rect 895 328 899 332
rect 943 328 947 332
rect 991 328 995 332
rect 1039 328 1043 332
rect 1087 328 1091 332
rect 1135 328 1139 332
rect 1183 328 1187 332
rect 1231 328 1235 332
rect 1279 328 1283 332
rect 1291 327 1292 331
rect 1292 327 1295 331
rect 1327 328 1331 332
rect 1383 328 1387 332
rect 1415 328 1419 332
rect 1447 325 1451 329
rect 451 319 455 323
rect 627 319 631 323
rect 1027 319 1031 323
rect 1259 319 1263 323
rect 111 307 115 311
rect 175 302 179 306
rect 184 303 188 307
rect 199 302 203 306
rect 211 303 212 307
rect 212 303 215 307
rect 223 302 227 306
rect 247 302 251 306
rect 259 303 260 307
rect 260 303 263 307
rect 279 302 283 306
rect 319 302 323 306
rect 331 303 332 307
rect 332 303 335 307
rect 359 302 363 306
rect 399 302 403 306
rect 411 303 412 307
rect 412 303 415 307
rect 439 302 443 306
rect 451 303 452 307
rect 452 303 455 307
rect 519 311 523 315
rect 479 302 483 306
rect 527 302 531 306
rect 583 302 587 306
rect 639 302 643 306
rect 687 302 691 306
rect 247 286 251 290
rect 519 291 523 295
rect 571 295 575 299
rect 735 302 739 306
rect 791 302 795 306
rect 847 302 851 306
rect 895 302 899 306
rect 943 302 947 306
rect 991 302 995 306
rect 771 295 775 299
rect 1039 302 1043 306
rect 1087 302 1091 306
rect 1135 302 1139 306
rect 1183 302 1187 306
rect 1427 311 1428 315
rect 1428 311 1431 315
rect 1231 302 1235 306
rect 1279 302 1283 306
rect 1327 302 1331 306
rect 1375 299 1379 303
rect 1383 302 1387 306
rect 1447 307 1451 311
rect 1403 303 1407 307
rect 1415 302 1419 306
rect 271 286 275 290
rect 111 281 115 285
rect 295 286 299 290
rect 307 283 308 287
rect 308 283 311 287
rect 319 286 323 290
rect 343 286 347 290
rect 367 286 371 290
rect 399 286 403 290
rect 431 286 435 290
rect 471 286 475 290
rect 111 263 115 267
rect 295 271 299 275
rect 511 286 515 290
rect 559 286 563 290
rect 247 260 251 264
rect 271 260 275 264
rect 295 260 299 264
rect 319 260 323 264
rect 343 260 347 264
rect 367 260 371 264
rect 419 271 423 275
rect 615 286 619 290
rect 571 275 572 279
rect 572 275 575 279
rect 663 286 667 290
rect 711 286 715 290
rect 723 283 724 287
rect 724 283 727 287
rect 759 286 763 290
rect 807 286 811 290
rect 771 275 772 279
rect 772 275 775 279
rect 847 286 851 290
rect 879 286 883 290
rect 903 286 907 290
rect 927 286 931 290
rect 951 286 955 290
rect 975 286 979 290
rect 999 286 1003 290
rect 1023 286 1027 290
rect 1047 286 1051 290
rect 1071 286 1075 290
rect 1095 286 1099 290
rect 1127 286 1131 290
rect 1159 286 1163 290
rect 1199 286 1203 290
rect 1247 286 1251 290
rect 1259 287 1260 291
rect 1260 287 1263 291
rect 1303 286 1307 290
rect 1315 283 1316 287
rect 1316 283 1319 287
rect 1367 286 1371 290
rect 1415 286 1419 290
rect 1427 287 1428 291
rect 1428 287 1431 291
rect 1447 281 1451 285
rect 399 260 403 264
rect 411 263 412 267
rect 412 263 415 267
rect 431 260 435 264
rect 471 260 475 264
rect 511 260 515 264
rect 559 260 563 264
rect 615 260 619 264
rect 663 260 667 264
rect 711 260 715 264
rect 759 260 763 264
rect 807 260 811 264
rect 847 260 851 264
rect 879 260 883 264
rect 903 260 907 264
rect 927 260 931 264
rect 951 260 955 264
rect 975 260 979 264
rect 999 260 1003 264
rect 1023 260 1027 264
rect 1047 260 1051 264
rect 1071 260 1075 264
rect 1095 260 1099 264
rect 1127 260 1131 264
rect 1159 260 1163 264
rect 1199 260 1203 264
rect 1247 260 1251 264
rect 1303 260 1307 264
rect 1367 260 1371 264
rect 1379 263 1380 267
rect 1380 263 1383 267
rect 1415 260 1419 264
rect 1447 263 1451 267
rect 111 245 115 249
rect 263 248 267 252
rect 287 248 291 252
rect 311 248 315 252
rect 335 248 339 252
rect 359 248 363 252
rect 383 248 387 252
rect 407 248 411 252
rect 431 248 435 252
rect 463 248 467 252
rect 503 248 507 252
rect 543 248 547 252
rect 583 248 587 252
rect 623 248 627 252
rect 679 248 683 252
rect 743 248 747 252
rect 807 248 811 252
rect 879 248 883 252
rect 959 248 963 252
rect 1039 248 1043 252
rect 1119 248 1123 252
rect 1199 248 1203 252
rect 1279 248 1283 252
rect 1315 247 1319 251
rect 1359 248 1363 252
rect 1415 248 1419 252
rect 1447 245 1451 249
rect 323 239 327 243
rect 111 227 115 231
rect 347 239 351 243
rect 359 235 363 239
rect 395 239 399 243
rect 475 239 479 243
rect 555 239 559 243
rect 263 222 267 226
rect 275 223 276 227
rect 276 223 279 227
rect 287 222 291 226
rect 311 222 315 226
rect 323 223 324 227
rect 324 223 327 227
rect 335 222 339 226
rect 347 223 348 227
rect 348 223 351 227
rect 359 222 363 226
rect 383 222 387 226
rect 407 222 411 226
rect 419 223 420 227
rect 420 223 423 227
rect 431 222 435 226
rect 367 215 371 219
rect 463 222 467 226
rect 475 223 476 227
rect 476 223 479 227
rect 591 235 592 239
rect 592 235 595 239
rect 723 239 727 243
rect 1131 239 1135 243
rect 503 222 507 226
rect 543 222 547 226
rect 555 223 556 227
rect 556 223 559 227
rect 583 222 587 226
rect 623 222 627 226
rect 679 222 683 226
rect 743 222 747 226
rect 807 222 811 226
rect 879 222 883 226
rect 959 222 963 226
rect 731 215 735 219
rect 1039 222 1043 226
rect 1095 219 1099 223
rect 1119 222 1123 226
rect 1131 223 1132 227
rect 1132 223 1135 227
rect 1199 222 1203 226
rect 1279 222 1283 226
rect 1359 222 1363 226
rect 1427 231 1428 235
rect 1428 231 1431 235
rect 1447 227 1451 231
rect 1415 222 1419 226
rect 239 206 243 210
rect 111 201 115 205
rect 263 206 267 210
rect 287 206 291 210
rect 311 206 315 210
rect 335 206 339 210
rect 359 206 363 210
rect 383 206 387 210
rect 395 207 396 211
rect 396 207 399 211
rect 407 206 411 210
rect 419 203 420 207
rect 420 203 423 207
rect 431 206 435 210
rect 463 206 467 210
rect 511 206 515 210
rect 559 206 563 210
rect 615 206 619 210
rect 671 206 675 210
rect 719 206 723 210
rect 767 206 771 210
rect 731 195 732 199
rect 732 195 735 199
rect 815 206 819 210
rect 863 206 867 210
rect 919 206 923 210
rect 975 206 979 210
rect 1031 206 1035 210
rect 1087 206 1091 210
rect 1135 206 1139 210
rect 1095 195 1096 199
rect 1096 195 1099 199
rect 1183 206 1187 210
rect 1195 203 1196 207
rect 1196 203 1199 207
rect 1231 206 1235 210
rect 1279 206 1283 210
rect 1327 206 1331 210
rect 1383 206 1387 210
rect 111 183 115 187
rect 239 180 243 184
rect 251 179 252 183
rect 252 179 255 183
rect 263 180 267 184
rect 287 180 291 184
rect 311 180 315 184
rect 335 180 339 184
rect 359 180 363 184
rect 383 180 387 184
rect 407 180 411 184
rect 431 180 435 184
rect 463 180 467 184
rect 511 180 515 184
rect 559 180 563 184
rect 615 180 619 184
rect 1415 206 1419 210
rect 1427 207 1428 211
rect 1428 207 1431 211
rect 1371 195 1375 199
rect 1447 201 1451 205
rect 671 180 675 184
rect 683 179 684 183
rect 684 179 687 183
rect 719 180 723 184
rect 767 180 771 184
rect 815 180 819 184
rect 863 180 867 184
rect 919 180 923 184
rect 975 180 979 184
rect 1031 180 1035 184
rect 1087 180 1091 184
rect 1135 180 1139 184
rect 1183 180 1187 184
rect 1231 180 1235 184
rect 1271 179 1275 183
rect 1279 180 1283 184
rect 1327 180 1331 184
rect 1383 180 1387 184
rect 1415 180 1419 184
rect 1427 179 1428 183
rect 1428 179 1431 183
rect 1447 183 1451 187
rect 111 165 115 169
rect 183 168 187 172
rect 207 168 211 172
rect 239 168 243 172
rect 279 168 283 172
rect 327 168 331 172
rect 375 168 379 172
rect 423 168 427 172
rect 471 168 475 172
rect 527 168 531 172
rect 591 168 595 172
rect 655 168 659 172
rect 711 168 715 172
rect 767 168 771 172
rect 823 168 827 172
rect 871 168 875 172
rect 919 168 923 172
rect 975 168 979 172
rect 1031 168 1035 172
rect 1079 168 1083 172
rect 1127 168 1131 172
rect 1175 168 1179 172
rect 1223 168 1227 172
rect 1263 168 1267 172
rect 1295 168 1299 172
rect 1327 168 1331 172
rect 1359 168 1363 172
rect 1371 167 1372 171
rect 1372 167 1375 171
rect 1391 168 1395 172
rect 1415 168 1419 172
rect 1447 165 1451 169
rect 411 159 415 163
rect 483 159 487 163
rect 603 159 607 163
rect 723 159 727 163
rect 883 159 887 163
rect 987 159 991 163
rect 1091 159 1095 163
rect 1195 159 1199 163
rect 111 147 115 151
rect 183 142 187 146
rect 207 142 211 146
rect 239 142 243 146
rect 279 142 283 146
rect 327 142 331 146
rect 375 142 379 146
rect 251 135 255 139
rect 423 142 427 146
rect 471 142 475 146
rect 483 143 484 147
rect 484 143 487 147
rect 671 151 675 155
rect 527 142 531 146
rect 591 142 595 146
rect 603 143 604 147
rect 604 143 607 147
rect 655 142 659 146
rect 711 142 715 146
rect 723 143 724 147
rect 724 143 727 147
rect 767 142 771 146
rect 823 142 827 146
rect 871 142 875 146
rect 883 143 884 147
rect 884 143 887 147
rect 683 131 687 135
rect 919 142 923 146
rect 975 142 979 146
rect 987 143 988 147
rect 988 143 991 147
rect 1031 142 1035 146
rect 1079 142 1083 146
rect 1091 143 1092 147
rect 1092 143 1095 147
rect 1127 142 1131 146
rect 1023 131 1027 135
rect 1055 135 1059 139
rect 1175 142 1179 146
rect 1223 142 1227 146
rect 1263 142 1267 146
rect 1399 155 1400 159
rect 1400 155 1403 159
rect 1295 142 1299 146
rect 1271 135 1275 139
rect 1327 142 1331 146
rect 1359 142 1363 146
rect 1391 142 1395 146
rect 1415 142 1419 146
rect 1427 143 1428 147
rect 1428 143 1431 147
rect 1447 147 1451 151
rect 1375 135 1379 139
rect 135 114 139 118
rect 111 109 115 113
rect 159 114 163 118
rect 183 114 187 118
rect 207 114 211 118
rect 231 114 235 118
rect 243 111 244 115
rect 244 111 247 115
rect 255 114 259 118
rect 279 114 283 118
rect 303 114 307 118
rect 327 114 331 118
rect 351 114 355 118
rect 375 114 379 118
rect 399 114 403 118
rect 411 115 412 119
rect 412 115 415 119
rect 431 114 435 118
rect 671 123 675 127
rect 1399 123 1403 127
rect 463 114 467 118
rect 475 111 476 115
rect 476 111 479 115
rect 487 114 491 118
rect 511 114 515 118
rect 535 114 539 118
rect 559 114 563 118
rect 583 114 587 118
rect 607 114 611 118
rect 631 114 635 118
rect 655 114 659 118
rect 679 114 683 118
rect 703 114 707 118
rect 727 114 731 118
rect 751 114 755 118
rect 775 114 779 118
rect 799 114 803 118
rect 823 114 827 118
rect 855 114 859 118
rect 887 114 891 118
rect 919 114 923 118
rect 951 114 955 118
rect 983 114 987 118
rect 1015 114 1019 118
rect 1047 114 1051 118
rect 1071 114 1075 118
rect 463 103 467 107
rect 1055 103 1056 107
rect 1056 103 1059 107
rect 1095 114 1099 118
rect 1119 114 1123 118
rect 1143 114 1147 118
rect 1175 114 1179 118
rect 1207 114 1211 118
rect 1239 114 1243 118
rect 1271 114 1275 118
rect 1303 114 1307 118
rect 1335 114 1339 118
rect 1367 114 1371 118
rect 1391 114 1395 118
rect 1375 103 1376 107
rect 1376 103 1379 107
rect 1415 114 1419 118
rect 1447 109 1451 113
rect 111 91 115 95
rect 135 88 139 92
rect 159 88 163 92
rect 183 88 187 92
rect 207 88 211 92
rect 231 88 235 92
rect 255 88 259 92
rect 279 88 283 92
rect 303 88 307 92
rect 327 88 331 92
rect 351 88 355 92
rect 375 88 379 92
rect 399 88 403 92
rect 431 88 435 92
rect 463 88 467 92
rect 487 88 491 92
rect 511 88 515 92
rect 535 88 539 92
rect 559 88 563 92
rect 583 88 587 92
rect 607 88 611 92
rect 631 88 635 92
rect 655 88 659 92
rect 679 88 683 92
rect 703 88 707 92
rect 727 88 731 92
rect 751 88 755 92
rect 775 88 779 92
rect 799 88 803 92
rect 823 88 827 92
rect 855 88 859 92
rect 887 88 891 92
rect 919 88 923 92
rect 951 88 955 92
rect 983 88 987 92
rect 1015 88 1019 92
rect 1027 91 1028 95
rect 1028 91 1031 95
rect 1047 88 1051 92
rect 1071 88 1075 92
rect 1095 88 1099 92
rect 1119 88 1123 92
rect 1143 88 1147 92
rect 1175 88 1179 92
rect 1207 88 1211 92
rect 1239 88 1243 92
rect 1271 88 1275 92
rect 1303 88 1307 92
rect 1335 88 1339 92
rect 1367 88 1371 92
rect 1391 88 1395 92
rect 1415 88 1419 92
rect 1447 91 1451 95
rect 243 79 247 83
<< m3 >>
rect 818 1511 824 1512
rect 111 1510 115 1511
rect 111 1505 115 1506
rect 295 1510 299 1511
rect 295 1505 299 1506
rect 319 1510 323 1511
rect 319 1505 323 1506
rect 343 1510 347 1511
rect 343 1505 347 1506
rect 367 1510 371 1511
rect 367 1505 371 1506
rect 407 1510 411 1511
rect 407 1505 411 1506
rect 455 1510 459 1511
rect 455 1505 459 1506
rect 511 1510 515 1511
rect 511 1505 515 1506
rect 575 1510 579 1511
rect 575 1505 579 1506
rect 647 1510 651 1511
rect 647 1505 651 1506
rect 727 1510 731 1511
rect 727 1505 731 1506
rect 807 1510 811 1511
rect 818 1507 819 1511
rect 823 1507 824 1511
rect 818 1506 824 1507
rect 887 1510 891 1511
rect 807 1505 811 1506
rect 112 1498 114 1505
rect 296 1503 298 1505
rect 320 1503 322 1505
rect 344 1503 346 1505
rect 368 1503 370 1505
rect 408 1503 410 1505
rect 456 1503 458 1505
rect 512 1503 514 1505
rect 576 1503 578 1505
rect 648 1503 650 1505
rect 728 1503 730 1505
rect 808 1503 810 1505
rect 294 1502 300 1503
rect 294 1498 295 1502
rect 299 1498 300 1502
rect 110 1497 116 1498
rect 294 1497 300 1498
rect 318 1502 324 1503
rect 318 1498 319 1502
rect 323 1498 324 1502
rect 318 1497 324 1498
rect 342 1502 348 1503
rect 342 1498 343 1502
rect 347 1498 348 1502
rect 342 1497 348 1498
rect 366 1502 372 1503
rect 366 1498 367 1502
rect 371 1498 372 1502
rect 366 1497 372 1498
rect 406 1502 412 1503
rect 406 1498 407 1502
rect 411 1498 412 1502
rect 406 1497 412 1498
rect 454 1502 460 1503
rect 454 1498 455 1502
rect 459 1498 460 1502
rect 454 1497 460 1498
rect 510 1502 516 1503
rect 510 1498 511 1502
rect 515 1498 516 1502
rect 510 1497 516 1498
rect 574 1502 580 1503
rect 574 1498 575 1502
rect 579 1498 580 1502
rect 574 1497 580 1498
rect 646 1502 652 1503
rect 646 1498 647 1502
rect 651 1498 652 1502
rect 646 1497 652 1498
rect 726 1502 732 1503
rect 726 1498 727 1502
rect 731 1498 732 1502
rect 726 1497 732 1498
rect 806 1502 812 1503
rect 806 1498 807 1502
rect 811 1498 812 1502
rect 806 1497 812 1498
rect 110 1493 111 1497
rect 115 1493 116 1497
rect 110 1492 116 1493
rect 820 1484 822 1506
rect 887 1505 891 1506
rect 959 1510 963 1511
rect 959 1505 963 1506
rect 1031 1510 1035 1511
rect 1031 1505 1035 1506
rect 1103 1510 1107 1511
rect 1103 1505 1107 1506
rect 1175 1510 1179 1511
rect 1175 1505 1179 1506
rect 1247 1510 1251 1511
rect 1247 1505 1251 1506
rect 1447 1510 1451 1511
rect 1447 1505 1451 1506
rect 888 1503 890 1505
rect 960 1503 962 1505
rect 1032 1503 1034 1505
rect 1104 1503 1106 1505
rect 1176 1503 1178 1505
rect 1248 1503 1250 1505
rect 886 1502 892 1503
rect 886 1498 887 1502
rect 891 1498 892 1502
rect 886 1497 892 1498
rect 958 1502 964 1503
rect 958 1498 959 1502
rect 963 1498 964 1502
rect 958 1497 964 1498
rect 1030 1502 1036 1503
rect 1030 1498 1031 1502
rect 1035 1498 1036 1502
rect 1102 1502 1108 1503
rect 1030 1497 1036 1498
rect 1082 1499 1088 1500
rect 1082 1495 1083 1499
rect 1087 1495 1088 1499
rect 1102 1498 1103 1502
rect 1107 1498 1108 1502
rect 1174 1502 1180 1503
rect 1102 1497 1108 1498
rect 1114 1499 1120 1500
rect 1082 1494 1088 1495
rect 1114 1495 1115 1499
rect 1119 1495 1120 1499
rect 1174 1498 1175 1502
rect 1179 1498 1180 1502
rect 1174 1497 1180 1498
rect 1246 1502 1252 1503
rect 1246 1498 1247 1502
rect 1251 1498 1252 1502
rect 1448 1498 1450 1505
rect 1246 1497 1252 1498
rect 1446 1497 1452 1498
rect 1114 1494 1120 1495
rect 818 1483 824 1484
rect 110 1479 116 1480
rect 110 1475 111 1479
rect 115 1475 116 1479
rect 818 1479 819 1483
rect 823 1479 824 1483
rect 818 1478 824 1479
rect 110 1474 116 1475
rect 294 1476 300 1477
rect 318 1476 324 1477
rect 112 1471 114 1474
rect 294 1472 295 1476
rect 299 1472 300 1476
rect 294 1471 300 1472
rect 306 1475 312 1476
rect 306 1471 307 1475
rect 311 1471 312 1475
rect 318 1472 319 1476
rect 323 1472 324 1476
rect 318 1471 324 1472
rect 342 1476 348 1477
rect 342 1472 343 1476
rect 347 1472 348 1476
rect 342 1471 348 1472
rect 366 1476 372 1477
rect 366 1472 367 1476
rect 371 1472 372 1476
rect 366 1471 372 1472
rect 406 1476 412 1477
rect 406 1472 407 1476
rect 411 1472 412 1476
rect 406 1471 412 1472
rect 454 1476 460 1477
rect 454 1472 455 1476
rect 459 1472 460 1476
rect 454 1471 460 1472
rect 510 1476 516 1477
rect 510 1472 511 1476
rect 515 1472 516 1476
rect 510 1471 516 1472
rect 574 1476 580 1477
rect 574 1472 575 1476
rect 579 1472 580 1476
rect 574 1471 580 1472
rect 646 1476 652 1477
rect 646 1472 647 1476
rect 651 1472 652 1476
rect 646 1471 652 1472
rect 726 1476 732 1477
rect 726 1472 727 1476
rect 731 1472 732 1476
rect 726 1471 732 1472
rect 806 1476 812 1477
rect 806 1472 807 1476
rect 811 1472 812 1476
rect 806 1471 812 1472
rect 886 1476 892 1477
rect 886 1472 887 1476
rect 891 1472 892 1476
rect 886 1471 892 1472
rect 958 1476 964 1477
rect 958 1472 959 1476
rect 963 1472 964 1476
rect 958 1471 964 1472
rect 1030 1476 1036 1477
rect 1030 1472 1031 1476
rect 1035 1472 1036 1476
rect 1030 1471 1036 1472
rect 111 1470 115 1471
rect 111 1465 115 1466
rect 151 1470 155 1471
rect 151 1465 155 1466
rect 175 1470 179 1471
rect 175 1465 179 1466
rect 199 1470 203 1471
rect 199 1465 203 1466
rect 231 1470 235 1471
rect 231 1465 235 1466
rect 271 1470 275 1471
rect 271 1465 275 1466
rect 295 1470 299 1471
rect 306 1470 312 1471
rect 319 1470 323 1471
rect 295 1465 299 1466
rect 112 1462 114 1465
rect 150 1464 156 1465
rect 110 1461 116 1462
rect 110 1457 111 1461
rect 115 1457 116 1461
rect 150 1460 151 1464
rect 155 1460 156 1464
rect 150 1459 156 1460
rect 174 1464 180 1465
rect 174 1460 175 1464
rect 179 1460 180 1464
rect 174 1459 180 1460
rect 198 1464 204 1465
rect 198 1460 199 1464
rect 203 1460 204 1464
rect 198 1459 204 1460
rect 230 1464 236 1465
rect 230 1460 231 1464
rect 235 1460 236 1464
rect 230 1459 236 1460
rect 270 1464 276 1465
rect 270 1460 271 1464
rect 275 1460 276 1464
rect 270 1459 276 1460
rect 110 1456 116 1457
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 110 1438 116 1439
rect 150 1438 156 1439
rect 112 1431 114 1438
rect 150 1434 151 1438
rect 155 1434 156 1438
rect 150 1433 156 1434
rect 174 1438 180 1439
rect 174 1434 175 1438
rect 179 1434 180 1438
rect 174 1433 180 1434
rect 198 1438 204 1439
rect 198 1434 199 1438
rect 203 1434 204 1438
rect 198 1433 204 1434
rect 230 1438 236 1439
rect 230 1434 231 1438
rect 235 1434 236 1438
rect 230 1433 236 1434
rect 270 1438 276 1439
rect 270 1434 271 1438
rect 275 1434 276 1438
rect 270 1433 276 1434
rect 152 1431 154 1433
rect 176 1431 178 1433
rect 200 1431 202 1433
rect 206 1431 212 1432
rect 232 1431 234 1433
rect 272 1431 274 1433
rect 308 1432 310 1470
rect 319 1465 323 1466
rect 343 1470 347 1471
rect 343 1465 347 1466
rect 367 1470 371 1471
rect 367 1465 371 1466
rect 407 1470 411 1471
rect 407 1465 411 1466
rect 455 1470 459 1471
rect 455 1465 459 1466
rect 503 1470 507 1471
rect 503 1465 507 1466
rect 511 1470 515 1471
rect 511 1465 515 1466
rect 551 1470 555 1471
rect 551 1465 555 1466
rect 575 1470 579 1471
rect 575 1465 579 1466
rect 607 1470 611 1471
rect 607 1465 611 1466
rect 647 1470 651 1471
rect 647 1465 651 1466
rect 663 1470 667 1471
rect 663 1465 667 1466
rect 711 1470 715 1471
rect 711 1465 715 1466
rect 727 1470 731 1471
rect 727 1465 731 1466
rect 759 1470 763 1471
rect 759 1465 763 1466
rect 807 1470 811 1471
rect 807 1465 811 1466
rect 815 1470 819 1471
rect 815 1465 819 1466
rect 871 1470 875 1471
rect 871 1465 875 1466
rect 887 1470 891 1471
rect 887 1465 891 1466
rect 927 1470 931 1471
rect 927 1465 931 1466
rect 959 1470 963 1471
rect 959 1465 963 1466
rect 975 1470 979 1471
rect 975 1465 979 1466
rect 1023 1470 1027 1471
rect 1023 1465 1027 1466
rect 1031 1470 1035 1471
rect 1031 1465 1035 1466
rect 1071 1470 1075 1471
rect 1071 1465 1075 1466
rect 318 1464 324 1465
rect 318 1460 319 1464
rect 323 1460 324 1464
rect 318 1459 324 1460
rect 366 1464 372 1465
rect 366 1460 367 1464
rect 371 1460 372 1464
rect 366 1459 372 1460
rect 406 1464 412 1465
rect 406 1460 407 1464
rect 411 1460 412 1464
rect 406 1459 412 1460
rect 454 1464 460 1465
rect 454 1460 455 1464
rect 459 1460 460 1464
rect 454 1459 460 1460
rect 502 1464 508 1465
rect 502 1460 503 1464
rect 507 1460 508 1464
rect 502 1459 508 1460
rect 550 1464 556 1465
rect 550 1460 551 1464
rect 555 1460 556 1464
rect 550 1459 556 1460
rect 606 1464 612 1465
rect 606 1460 607 1464
rect 611 1460 612 1464
rect 606 1459 612 1460
rect 662 1464 668 1465
rect 662 1460 663 1464
rect 667 1460 668 1464
rect 662 1459 668 1460
rect 710 1464 716 1465
rect 710 1460 711 1464
rect 715 1460 716 1464
rect 710 1459 716 1460
rect 758 1464 764 1465
rect 758 1460 759 1464
rect 763 1460 764 1464
rect 758 1459 764 1460
rect 814 1464 820 1465
rect 814 1460 815 1464
rect 819 1460 820 1464
rect 814 1459 820 1460
rect 870 1464 876 1465
rect 870 1460 871 1464
rect 875 1460 876 1464
rect 870 1459 876 1460
rect 926 1464 932 1465
rect 926 1460 927 1464
rect 931 1460 932 1464
rect 926 1459 932 1460
rect 974 1464 980 1465
rect 974 1460 975 1464
rect 979 1460 980 1464
rect 974 1459 980 1460
rect 1022 1464 1028 1465
rect 1022 1460 1023 1464
rect 1027 1460 1028 1464
rect 1022 1459 1028 1460
rect 1070 1464 1076 1465
rect 1084 1464 1086 1494
rect 1102 1491 1108 1492
rect 1116 1491 1118 1494
rect 1446 1493 1447 1497
rect 1451 1493 1452 1497
rect 1446 1492 1452 1493
rect 1102 1487 1103 1491
rect 1107 1489 1118 1491
rect 1107 1487 1108 1489
rect 1102 1486 1108 1487
rect 1446 1479 1452 1480
rect 1102 1476 1108 1477
rect 1102 1472 1103 1476
rect 1107 1472 1108 1476
rect 1102 1471 1108 1472
rect 1174 1476 1180 1477
rect 1174 1472 1175 1476
rect 1179 1472 1180 1476
rect 1174 1471 1180 1472
rect 1246 1476 1252 1477
rect 1246 1472 1247 1476
rect 1251 1472 1252 1476
rect 1446 1475 1447 1479
rect 1451 1475 1452 1479
rect 1446 1474 1452 1475
rect 1246 1471 1252 1472
rect 1448 1471 1450 1474
rect 1103 1470 1107 1471
rect 1103 1465 1107 1466
rect 1119 1470 1123 1471
rect 1119 1465 1123 1466
rect 1167 1470 1171 1471
rect 1167 1465 1171 1466
rect 1175 1470 1179 1471
rect 1175 1465 1179 1466
rect 1215 1470 1219 1471
rect 1215 1465 1219 1466
rect 1247 1470 1251 1471
rect 1247 1465 1251 1466
rect 1263 1470 1267 1471
rect 1263 1465 1267 1466
rect 1311 1470 1315 1471
rect 1311 1465 1315 1466
rect 1447 1470 1451 1471
rect 1447 1465 1451 1466
rect 1118 1464 1124 1465
rect 1070 1460 1071 1464
rect 1075 1460 1076 1464
rect 1070 1459 1076 1460
rect 1082 1463 1088 1464
rect 1082 1459 1083 1463
rect 1087 1459 1088 1463
rect 1118 1460 1119 1464
rect 1123 1460 1124 1464
rect 1118 1459 1124 1460
rect 1166 1464 1172 1465
rect 1166 1460 1167 1464
rect 1171 1460 1172 1464
rect 1166 1459 1172 1460
rect 1214 1464 1220 1465
rect 1214 1460 1215 1464
rect 1219 1460 1220 1464
rect 1214 1459 1220 1460
rect 1262 1464 1268 1465
rect 1262 1460 1263 1464
rect 1267 1460 1268 1464
rect 1262 1459 1268 1460
rect 1310 1464 1316 1465
rect 1310 1460 1311 1464
rect 1315 1460 1316 1464
rect 1448 1462 1450 1465
rect 1310 1459 1316 1460
rect 1446 1461 1452 1462
rect 1082 1458 1088 1459
rect 1446 1457 1447 1461
rect 1451 1457 1452 1461
rect 1446 1456 1452 1457
rect 426 1455 432 1456
rect 426 1451 427 1455
rect 431 1451 432 1455
rect 426 1450 432 1451
rect 826 1455 832 1456
rect 826 1451 827 1455
rect 831 1451 832 1455
rect 826 1450 832 1451
rect 986 1455 992 1456
rect 986 1451 987 1455
rect 991 1451 992 1455
rect 986 1450 992 1451
rect 1226 1455 1232 1456
rect 1226 1451 1227 1455
rect 1231 1451 1232 1455
rect 1226 1450 1232 1451
rect 1322 1455 1328 1456
rect 1322 1451 1323 1455
rect 1327 1451 1328 1455
rect 1322 1450 1328 1451
rect 318 1438 324 1439
rect 318 1434 319 1438
rect 323 1434 324 1438
rect 318 1433 324 1434
rect 366 1438 372 1439
rect 366 1434 367 1438
rect 371 1434 372 1438
rect 366 1433 372 1434
rect 406 1438 412 1439
rect 406 1434 407 1438
rect 411 1434 412 1438
rect 406 1433 412 1434
rect 298 1431 304 1432
rect 111 1430 115 1431
rect 111 1425 115 1426
rect 135 1430 139 1431
rect 135 1425 139 1426
rect 151 1430 155 1431
rect 151 1425 155 1426
rect 159 1430 163 1431
rect 159 1425 163 1426
rect 175 1430 179 1431
rect 175 1425 179 1426
rect 183 1430 187 1431
rect 183 1425 187 1426
rect 199 1430 203 1431
rect 206 1427 207 1431
rect 211 1427 212 1431
rect 206 1426 212 1427
rect 223 1430 227 1431
rect 199 1425 203 1426
rect 112 1418 114 1425
rect 136 1423 138 1425
rect 160 1423 162 1425
rect 184 1423 186 1425
rect 134 1422 140 1423
rect 134 1418 135 1422
rect 139 1418 140 1422
rect 110 1417 116 1418
rect 134 1417 140 1418
rect 158 1422 164 1423
rect 158 1418 159 1422
rect 163 1418 164 1422
rect 158 1417 164 1418
rect 182 1422 188 1423
rect 182 1418 183 1422
rect 187 1418 188 1422
rect 182 1417 188 1418
rect 110 1413 111 1417
rect 115 1413 116 1417
rect 110 1412 116 1413
rect 110 1399 116 1400
rect 110 1395 111 1399
rect 115 1395 116 1399
rect 110 1394 116 1395
rect 134 1396 140 1397
rect 158 1396 164 1397
rect 112 1391 114 1394
rect 134 1392 135 1396
rect 139 1392 140 1396
rect 134 1391 140 1392
rect 146 1395 152 1396
rect 146 1391 147 1395
rect 151 1391 152 1395
rect 158 1392 159 1396
rect 163 1392 164 1396
rect 158 1391 164 1392
rect 182 1396 188 1397
rect 182 1392 183 1396
rect 187 1392 188 1396
rect 182 1391 188 1392
rect 111 1390 115 1391
rect 111 1385 115 1386
rect 135 1390 139 1391
rect 146 1390 152 1391
rect 159 1390 163 1391
rect 135 1385 139 1386
rect 112 1382 114 1385
rect 134 1384 140 1385
rect 110 1381 116 1382
rect 110 1377 111 1381
rect 115 1377 116 1381
rect 134 1380 135 1384
rect 139 1380 140 1384
rect 134 1379 140 1380
rect 110 1376 116 1377
rect 110 1363 116 1364
rect 110 1359 111 1363
rect 115 1359 116 1363
rect 148 1360 150 1390
rect 159 1385 163 1386
rect 183 1390 187 1391
rect 183 1385 187 1386
rect 158 1384 164 1385
rect 158 1380 159 1384
rect 163 1380 164 1384
rect 158 1379 164 1380
rect 182 1384 188 1385
rect 182 1380 183 1384
rect 187 1380 188 1384
rect 182 1379 188 1380
rect 170 1375 176 1376
rect 170 1371 171 1375
rect 175 1371 176 1375
rect 170 1370 176 1371
rect 194 1375 200 1376
rect 194 1371 195 1375
rect 199 1371 200 1375
rect 194 1370 200 1371
rect 172 1360 174 1370
rect 196 1360 198 1370
rect 146 1359 152 1360
rect 170 1359 176 1360
rect 194 1359 200 1360
rect 110 1358 116 1359
rect 134 1358 140 1359
rect 112 1351 114 1358
rect 134 1354 135 1358
rect 139 1354 140 1358
rect 146 1355 147 1359
rect 151 1355 152 1359
rect 146 1354 152 1355
rect 158 1358 164 1359
rect 158 1354 159 1358
rect 163 1354 164 1358
rect 170 1355 171 1359
rect 175 1355 176 1359
rect 170 1354 176 1355
rect 182 1358 188 1359
rect 182 1354 183 1358
rect 187 1354 188 1358
rect 194 1355 195 1359
rect 199 1355 200 1359
rect 194 1354 200 1355
rect 134 1353 140 1354
rect 158 1353 164 1354
rect 182 1353 188 1354
rect 136 1351 138 1353
rect 160 1351 162 1353
rect 184 1351 186 1353
rect 208 1352 210 1426
rect 223 1425 227 1426
rect 231 1430 235 1431
rect 231 1425 235 1426
rect 271 1430 275 1431
rect 271 1425 275 1426
rect 287 1430 291 1431
rect 298 1427 299 1431
rect 303 1427 304 1431
rect 298 1426 304 1427
rect 306 1431 312 1432
rect 320 1431 322 1433
rect 368 1431 370 1433
rect 408 1431 410 1433
rect 306 1427 307 1431
rect 311 1427 312 1431
rect 306 1426 312 1427
rect 319 1430 323 1431
rect 287 1425 291 1426
rect 224 1423 226 1425
rect 288 1423 290 1425
rect 222 1422 228 1423
rect 222 1418 223 1422
rect 227 1418 228 1422
rect 222 1417 228 1418
rect 286 1422 292 1423
rect 286 1418 287 1422
rect 291 1418 292 1422
rect 286 1417 292 1418
rect 222 1396 228 1397
rect 222 1392 223 1396
rect 227 1392 228 1396
rect 222 1391 228 1392
rect 286 1396 292 1397
rect 286 1392 287 1396
rect 291 1392 292 1396
rect 286 1391 292 1392
rect 223 1390 227 1391
rect 223 1385 227 1386
rect 231 1390 235 1391
rect 231 1385 235 1386
rect 279 1390 283 1391
rect 279 1385 283 1386
rect 287 1390 291 1391
rect 287 1385 291 1386
rect 230 1384 236 1385
rect 230 1380 231 1384
rect 235 1380 236 1384
rect 230 1379 236 1380
rect 278 1384 284 1385
rect 278 1380 279 1384
rect 283 1380 284 1384
rect 278 1379 284 1380
rect 300 1376 302 1426
rect 319 1425 323 1426
rect 351 1430 355 1431
rect 351 1425 355 1426
rect 367 1430 371 1431
rect 367 1425 371 1426
rect 407 1430 411 1431
rect 407 1425 411 1426
rect 415 1430 419 1431
rect 415 1425 419 1426
rect 352 1423 354 1425
rect 416 1423 418 1425
rect 428 1424 430 1450
rect 828 1440 830 1450
rect 988 1440 990 1450
rect 1034 1447 1040 1448
rect 1034 1443 1035 1447
rect 1039 1443 1040 1447
rect 1034 1442 1040 1443
rect 826 1439 832 1440
rect 986 1439 992 1440
rect 454 1438 460 1439
rect 454 1434 455 1438
rect 459 1434 460 1438
rect 454 1433 460 1434
rect 502 1438 508 1439
rect 502 1434 503 1438
rect 507 1434 508 1438
rect 502 1433 508 1434
rect 550 1438 556 1439
rect 550 1434 551 1438
rect 555 1434 556 1438
rect 550 1433 556 1434
rect 606 1438 612 1439
rect 606 1434 607 1438
rect 611 1434 612 1438
rect 606 1433 612 1434
rect 662 1438 668 1439
rect 662 1434 663 1438
rect 667 1434 668 1438
rect 662 1433 668 1434
rect 710 1438 716 1439
rect 710 1434 711 1438
rect 715 1434 716 1438
rect 710 1433 716 1434
rect 758 1438 764 1439
rect 758 1434 759 1438
rect 763 1434 764 1438
rect 758 1433 764 1434
rect 814 1438 820 1439
rect 814 1434 815 1438
rect 819 1434 820 1438
rect 826 1435 827 1439
rect 831 1435 832 1439
rect 826 1434 832 1435
rect 870 1438 876 1439
rect 870 1434 871 1438
rect 875 1434 876 1438
rect 814 1433 820 1434
rect 870 1433 876 1434
rect 926 1438 932 1439
rect 926 1434 927 1438
rect 931 1434 932 1438
rect 926 1433 932 1434
rect 974 1438 980 1439
rect 974 1434 975 1438
rect 979 1434 980 1438
rect 986 1435 987 1439
rect 991 1435 992 1439
rect 986 1434 992 1435
rect 1022 1438 1028 1439
rect 1022 1434 1023 1438
rect 1027 1434 1028 1438
rect 974 1433 980 1434
rect 1022 1433 1028 1434
rect 456 1431 458 1433
rect 504 1431 506 1433
rect 552 1431 554 1433
rect 558 1431 564 1432
rect 608 1431 610 1433
rect 664 1431 666 1433
rect 712 1431 714 1433
rect 760 1431 762 1433
rect 816 1431 818 1433
rect 872 1431 874 1433
rect 928 1431 930 1433
rect 976 1431 978 1433
rect 1024 1431 1026 1433
rect 455 1430 459 1431
rect 455 1425 459 1426
rect 479 1430 483 1431
rect 479 1425 483 1426
rect 503 1430 507 1431
rect 503 1425 507 1426
rect 535 1430 539 1431
rect 535 1425 539 1426
rect 551 1430 555 1431
rect 558 1427 559 1431
rect 563 1427 564 1431
rect 558 1426 564 1427
rect 583 1430 587 1431
rect 551 1425 555 1426
rect 426 1423 432 1424
rect 480 1423 482 1425
rect 536 1423 538 1425
rect 350 1422 356 1423
rect 350 1418 351 1422
rect 355 1418 356 1422
rect 350 1417 356 1418
rect 414 1422 420 1423
rect 414 1418 415 1422
rect 419 1418 420 1422
rect 426 1419 427 1423
rect 431 1419 432 1423
rect 426 1418 432 1419
rect 478 1422 484 1423
rect 478 1418 479 1422
rect 483 1418 484 1422
rect 414 1417 420 1418
rect 478 1417 484 1418
rect 534 1422 540 1423
rect 534 1418 535 1422
rect 539 1418 540 1422
rect 534 1417 540 1418
rect 560 1412 562 1426
rect 583 1425 587 1426
rect 607 1430 611 1431
rect 607 1425 611 1426
rect 631 1430 635 1431
rect 631 1425 635 1426
rect 663 1430 667 1431
rect 663 1425 667 1426
rect 687 1430 691 1431
rect 687 1425 691 1426
rect 711 1430 715 1431
rect 711 1425 715 1426
rect 743 1430 747 1431
rect 743 1425 747 1426
rect 759 1430 763 1431
rect 759 1425 763 1426
rect 799 1430 803 1431
rect 799 1425 803 1426
rect 815 1430 819 1431
rect 815 1425 819 1426
rect 855 1430 859 1431
rect 855 1425 859 1426
rect 871 1430 875 1431
rect 871 1425 875 1426
rect 911 1430 915 1431
rect 911 1425 915 1426
rect 927 1430 931 1431
rect 927 1425 931 1426
rect 967 1430 971 1431
rect 967 1425 971 1426
rect 975 1430 979 1431
rect 975 1425 979 1426
rect 1023 1430 1027 1431
rect 1023 1425 1027 1426
rect 584 1423 586 1425
rect 632 1423 634 1425
rect 688 1423 690 1425
rect 744 1423 746 1425
rect 800 1423 802 1425
rect 856 1423 858 1425
rect 912 1423 914 1425
rect 968 1423 970 1425
rect 1024 1423 1026 1425
rect 1036 1424 1038 1442
rect 1228 1440 1230 1450
rect 1274 1447 1280 1448
rect 1274 1443 1275 1447
rect 1279 1443 1280 1447
rect 1274 1442 1280 1443
rect 1226 1439 1232 1440
rect 1070 1438 1076 1439
rect 1070 1434 1071 1438
rect 1075 1434 1076 1438
rect 1070 1433 1076 1434
rect 1118 1438 1124 1439
rect 1118 1434 1119 1438
rect 1123 1434 1124 1438
rect 1166 1438 1172 1439
rect 1118 1433 1124 1434
rect 1130 1435 1136 1436
rect 1072 1431 1074 1433
rect 1120 1431 1122 1433
rect 1130 1431 1131 1435
rect 1135 1431 1136 1435
rect 1166 1434 1167 1438
rect 1171 1434 1172 1438
rect 1166 1433 1172 1434
rect 1214 1438 1220 1439
rect 1214 1434 1215 1438
rect 1219 1434 1220 1438
rect 1226 1435 1227 1439
rect 1231 1435 1232 1439
rect 1226 1434 1232 1435
rect 1262 1438 1268 1439
rect 1262 1434 1263 1438
rect 1267 1434 1268 1438
rect 1214 1433 1220 1434
rect 1262 1433 1268 1434
rect 1168 1431 1170 1433
rect 1216 1431 1218 1433
rect 1264 1431 1266 1433
rect 1071 1430 1075 1431
rect 1071 1425 1075 1426
rect 1119 1430 1123 1431
rect 1130 1430 1136 1431
rect 1167 1430 1171 1431
rect 1119 1425 1123 1426
rect 1034 1423 1040 1424
rect 1072 1423 1074 1425
rect 1120 1423 1122 1425
rect 582 1422 588 1423
rect 582 1418 583 1422
rect 587 1418 588 1422
rect 582 1417 588 1418
rect 630 1422 636 1423
rect 630 1418 631 1422
rect 635 1418 636 1422
rect 630 1417 636 1418
rect 686 1422 692 1423
rect 686 1418 687 1422
rect 691 1418 692 1422
rect 686 1417 692 1418
rect 742 1422 748 1423
rect 742 1418 743 1422
rect 747 1418 748 1422
rect 742 1417 748 1418
rect 798 1422 804 1423
rect 798 1418 799 1422
rect 803 1418 804 1422
rect 798 1417 804 1418
rect 854 1422 860 1423
rect 854 1418 855 1422
rect 859 1418 860 1422
rect 910 1422 916 1423
rect 854 1417 860 1418
rect 890 1419 896 1420
rect 890 1415 891 1419
rect 895 1415 896 1419
rect 910 1418 911 1422
rect 915 1418 916 1422
rect 910 1417 916 1418
rect 966 1422 972 1423
rect 966 1418 967 1422
rect 971 1418 972 1422
rect 966 1417 972 1418
rect 1022 1422 1028 1423
rect 1022 1418 1023 1422
rect 1027 1418 1028 1422
rect 1034 1419 1035 1423
rect 1039 1419 1040 1423
rect 1034 1418 1040 1419
rect 1070 1422 1076 1423
rect 1070 1418 1071 1422
rect 1075 1418 1076 1422
rect 1118 1422 1124 1423
rect 1022 1417 1028 1418
rect 1070 1417 1076 1418
rect 1082 1419 1088 1420
rect 890 1414 896 1415
rect 1082 1415 1083 1419
rect 1087 1415 1088 1419
rect 1118 1418 1119 1422
rect 1123 1418 1124 1422
rect 1118 1417 1124 1418
rect 1082 1414 1088 1415
rect 558 1411 564 1412
rect 558 1407 559 1411
rect 563 1407 564 1411
rect 558 1406 564 1407
rect 350 1396 356 1397
rect 350 1392 351 1396
rect 355 1392 356 1396
rect 350 1391 356 1392
rect 414 1396 420 1397
rect 414 1392 415 1396
rect 419 1392 420 1396
rect 414 1391 420 1392
rect 478 1396 484 1397
rect 478 1392 479 1396
rect 483 1392 484 1396
rect 478 1391 484 1392
rect 534 1396 540 1397
rect 534 1392 535 1396
rect 539 1392 540 1396
rect 534 1391 540 1392
rect 582 1396 588 1397
rect 582 1392 583 1396
rect 587 1392 588 1396
rect 582 1391 588 1392
rect 630 1396 636 1397
rect 630 1392 631 1396
rect 635 1392 636 1396
rect 630 1391 636 1392
rect 686 1396 692 1397
rect 686 1392 687 1396
rect 691 1392 692 1396
rect 686 1391 692 1392
rect 742 1396 748 1397
rect 742 1392 743 1396
rect 747 1392 748 1396
rect 742 1391 748 1392
rect 798 1396 804 1397
rect 798 1392 799 1396
rect 803 1392 804 1396
rect 798 1391 804 1392
rect 854 1396 860 1397
rect 854 1392 855 1396
rect 859 1392 860 1396
rect 854 1391 860 1392
rect 335 1390 339 1391
rect 335 1385 339 1386
rect 351 1390 355 1391
rect 351 1385 355 1386
rect 391 1390 395 1391
rect 391 1385 395 1386
rect 415 1390 419 1391
rect 415 1385 419 1386
rect 439 1390 443 1391
rect 439 1385 443 1386
rect 479 1390 483 1391
rect 479 1385 483 1386
rect 487 1390 491 1391
rect 487 1385 491 1386
rect 527 1390 531 1391
rect 527 1385 531 1386
rect 535 1390 539 1391
rect 535 1385 539 1386
rect 567 1390 571 1391
rect 567 1385 571 1386
rect 583 1390 587 1391
rect 583 1385 587 1386
rect 615 1390 619 1391
rect 615 1385 619 1386
rect 631 1390 635 1391
rect 631 1385 635 1386
rect 663 1390 667 1391
rect 663 1385 667 1386
rect 687 1390 691 1391
rect 687 1385 691 1386
rect 711 1390 715 1391
rect 711 1385 715 1386
rect 743 1390 747 1391
rect 743 1385 747 1386
rect 767 1390 771 1391
rect 767 1385 771 1386
rect 799 1390 803 1391
rect 799 1385 803 1386
rect 823 1390 827 1391
rect 823 1385 827 1386
rect 855 1390 859 1391
rect 855 1385 859 1386
rect 879 1390 883 1391
rect 879 1385 883 1386
rect 334 1384 340 1385
rect 334 1380 335 1384
rect 339 1380 340 1384
rect 334 1379 340 1380
rect 390 1384 396 1385
rect 390 1380 391 1384
rect 395 1380 396 1384
rect 390 1379 396 1380
rect 438 1384 444 1385
rect 438 1380 439 1384
rect 443 1380 444 1384
rect 438 1379 444 1380
rect 486 1384 492 1385
rect 486 1380 487 1384
rect 491 1380 492 1384
rect 486 1379 492 1380
rect 526 1384 532 1385
rect 526 1380 527 1384
rect 531 1380 532 1384
rect 526 1379 532 1380
rect 566 1384 572 1385
rect 566 1380 567 1384
rect 571 1380 572 1384
rect 566 1379 572 1380
rect 614 1384 620 1385
rect 614 1380 615 1384
rect 619 1380 620 1384
rect 614 1379 620 1380
rect 662 1384 668 1385
rect 662 1380 663 1384
rect 667 1380 668 1384
rect 662 1379 668 1380
rect 710 1384 716 1385
rect 710 1380 711 1384
rect 715 1380 716 1384
rect 710 1379 716 1380
rect 766 1384 772 1385
rect 766 1380 767 1384
rect 771 1380 772 1384
rect 766 1379 772 1380
rect 822 1384 828 1385
rect 822 1380 823 1384
rect 827 1380 828 1384
rect 822 1379 828 1380
rect 878 1384 884 1385
rect 892 1384 894 1414
rect 910 1396 916 1397
rect 966 1396 972 1397
rect 910 1392 911 1396
rect 915 1392 916 1396
rect 910 1391 916 1392
rect 946 1395 952 1396
rect 946 1391 947 1395
rect 951 1391 952 1395
rect 966 1392 967 1396
rect 971 1392 972 1396
rect 966 1391 972 1392
rect 1022 1396 1028 1397
rect 1022 1392 1023 1396
rect 1027 1392 1028 1396
rect 1022 1391 1028 1392
rect 1070 1396 1076 1397
rect 1070 1392 1071 1396
rect 1075 1392 1076 1396
rect 1070 1391 1076 1392
rect 911 1390 915 1391
rect 911 1385 915 1386
rect 935 1390 939 1391
rect 946 1390 952 1391
rect 967 1390 971 1391
rect 935 1385 939 1386
rect 934 1384 940 1385
rect 878 1380 879 1384
rect 883 1380 884 1384
rect 878 1379 884 1380
rect 890 1383 896 1384
rect 890 1379 891 1383
rect 895 1379 896 1383
rect 934 1380 935 1384
rect 939 1380 940 1384
rect 934 1379 940 1380
rect 890 1378 896 1379
rect 290 1375 296 1376
rect 290 1371 291 1375
rect 295 1371 296 1375
rect 290 1370 296 1371
rect 298 1375 304 1376
rect 298 1371 299 1375
rect 303 1371 304 1375
rect 298 1370 304 1371
rect 450 1375 456 1376
rect 450 1371 451 1375
rect 455 1371 456 1375
rect 450 1370 456 1371
rect 538 1375 544 1376
rect 538 1371 539 1375
rect 543 1371 544 1375
rect 538 1370 544 1371
rect 626 1375 632 1376
rect 626 1371 627 1375
rect 631 1371 632 1375
rect 626 1370 632 1371
rect 722 1375 728 1376
rect 722 1371 723 1375
rect 727 1371 728 1375
rect 722 1370 728 1371
rect 834 1375 840 1376
rect 834 1371 835 1375
rect 839 1371 840 1375
rect 834 1370 840 1371
rect 292 1360 294 1370
rect 452 1360 454 1370
rect 540 1360 542 1370
rect 628 1360 630 1370
rect 724 1360 726 1370
rect 836 1360 838 1370
rect 948 1360 950 1390
rect 967 1385 971 1386
rect 991 1390 995 1391
rect 991 1385 995 1386
rect 1023 1390 1027 1391
rect 1023 1385 1027 1386
rect 1047 1390 1051 1391
rect 1047 1385 1051 1386
rect 1071 1390 1075 1391
rect 1071 1385 1075 1386
rect 990 1384 996 1385
rect 990 1380 991 1384
rect 995 1380 996 1384
rect 990 1379 996 1380
rect 1046 1384 1052 1385
rect 1084 1384 1086 1414
rect 1132 1412 1134 1430
rect 1167 1425 1171 1426
rect 1215 1430 1219 1431
rect 1215 1425 1219 1426
rect 1263 1430 1267 1431
rect 1263 1425 1267 1426
rect 1168 1423 1170 1425
rect 1216 1423 1218 1425
rect 1264 1423 1266 1425
rect 1276 1424 1278 1442
rect 1324 1440 1326 1450
rect 1446 1443 1452 1444
rect 1322 1439 1328 1440
rect 1310 1438 1316 1439
rect 1310 1434 1311 1438
rect 1315 1434 1316 1438
rect 1322 1435 1323 1439
rect 1327 1435 1328 1439
rect 1446 1439 1447 1443
rect 1451 1439 1452 1443
rect 1446 1438 1452 1439
rect 1322 1434 1328 1435
rect 1310 1433 1316 1434
rect 1312 1431 1314 1433
rect 1354 1431 1360 1432
rect 1448 1431 1450 1438
rect 1303 1430 1307 1431
rect 1303 1425 1307 1426
rect 1311 1430 1315 1431
rect 1311 1425 1315 1426
rect 1343 1430 1347 1431
rect 1354 1427 1355 1431
rect 1359 1427 1360 1431
rect 1354 1426 1360 1427
rect 1391 1430 1395 1431
rect 1343 1425 1347 1426
rect 1274 1423 1280 1424
rect 1304 1423 1306 1425
rect 1344 1423 1346 1425
rect 1166 1422 1172 1423
rect 1138 1419 1144 1420
rect 1138 1415 1139 1419
rect 1143 1415 1144 1419
rect 1166 1418 1167 1422
rect 1171 1418 1172 1422
rect 1166 1417 1172 1418
rect 1214 1422 1220 1423
rect 1214 1418 1215 1422
rect 1219 1418 1220 1422
rect 1214 1417 1220 1418
rect 1262 1422 1268 1423
rect 1262 1418 1263 1422
rect 1267 1418 1268 1422
rect 1274 1419 1275 1423
rect 1279 1419 1280 1423
rect 1274 1418 1280 1419
rect 1302 1422 1308 1423
rect 1302 1418 1303 1422
rect 1307 1418 1308 1422
rect 1342 1422 1348 1423
rect 1262 1417 1268 1418
rect 1302 1417 1308 1418
rect 1314 1419 1320 1420
rect 1138 1414 1144 1415
rect 1314 1415 1315 1419
rect 1319 1415 1320 1419
rect 1342 1418 1343 1422
rect 1347 1418 1348 1422
rect 1342 1417 1348 1418
rect 1314 1414 1320 1415
rect 1130 1411 1136 1412
rect 1118 1407 1124 1408
rect 1118 1403 1119 1407
rect 1123 1403 1124 1407
rect 1130 1407 1131 1411
rect 1135 1407 1136 1411
rect 1130 1406 1136 1407
rect 1140 1403 1142 1414
rect 1118 1402 1142 1403
rect 1120 1401 1142 1402
rect 1118 1396 1124 1397
rect 1118 1392 1119 1396
rect 1123 1392 1124 1396
rect 1118 1391 1124 1392
rect 1166 1396 1172 1397
rect 1214 1396 1220 1397
rect 1166 1392 1167 1396
rect 1171 1392 1172 1396
rect 1166 1391 1172 1392
rect 1206 1395 1212 1396
rect 1206 1391 1207 1395
rect 1211 1391 1212 1395
rect 1214 1392 1215 1396
rect 1219 1392 1220 1396
rect 1214 1391 1220 1392
rect 1262 1396 1268 1397
rect 1262 1392 1263 1396
rect 1267 1392 1268 1396
rect 1262 1391 1268 1392
rect 1302 1396 1308 1397
rect 1302 1392 1303 1396
rect 1307 1392 1308 1396
rect 1302 1391 1308 1392
rect 1095 1390 1099 1391
rect 1095 1385 1099 1386
rect 1119 1390 1123 1391
rect 1119 1385 1123 1386
rect 1143 1390 1147 1391
rect 1143 1385 1147 1386
rect 1167 1390 1171 1391
rect 1167 1385 1171 1386
rect 1191 1390 1195 1391
rect 1206 1390 1212 1391
rect 1215 1390 1219 1391
rect 1191 1385 1195 1386
rect 1094 1384 1100 1385
rect 1046 1380 1047 1384
rect 1051 1380 1052 1384
rect 1046 1379 1052 1380
rect 1082 1383 1088 1384
rect 1082 1379 1083 1383
rect 1087 1379 1088 1383
rect 1094 1380 1095 1384
rect 1099 1380 1100 1384
rect 1094 1379 1100 1380
rect 1142 1384 1148 1385
rect 1142 1380 1143 1384
rect 1147 1380 1148 1384
rect 1142 1379 1148 1380
rect 1190 1384 1196 1385
rect 1190 1380 1191 1384
rect 1195 1380 1196 1384
rect 1190 1379 1196 1380
rect 1082 1378 1088 1379
rect 1002 1375 1008 1376
rect 1002 1371 1003 1375
rect 1007 1371 1008 1375
rect 1002 1370 1008 1371
rect 1004 1360 1006 1370
rect 1018 1367 1024 1368
rect 1018 1363 1019 1367
rect 1023 1363 1024 1367
rect 1018 1362 1024 1363
rect 1170 1367 1176 1368
rect 1170 1363 1171 1367
rect 1175 1363 1176 1367
rect 1170 1362 1176 1363
rect 290 1359 296 1360
rect 450 1359 456 1360
rect 538 1359 544 1360
rect 626 1359 632 1360
rect 722 1359 728 1360
rect 834 1359 840 1360
rect 946 1359 952 1360
rect 1002 1359 1008 1360
rect 230 1358 236 1359
rect 230 1354 231 1358
rect 235 1354 236 1358
rect 230 1353 236 1354
rect 278 1358 284 1359
rect 278 1354 279 1358
rect 283 1354 284 1358
rect 290 1355 291 1359
rect 295 1355 296 1359
rect 290 1354 296 1355
rect 334 1358 340 1359
rect 334 1354 335 1358
rect 339 1354 340 1358
rect 278 1353 284 1354
rect 334 1353 340 1354
rect 390 1358 396 1359
rect 390 1354 391 1358
rect 395 1354 396 1358
rect 390 1353 396 1354
rect 438 1358 444 1359
rect 438 1354 439 1358
rect 443 1354 444 1358
rect 450 1355 451 1359
rect 455 1355 456 1359
rect 450 1354 456 1355
rect 486 1358 492 1359
rect 486 1354 487 1358
rect 491 1354 492 1358
rect 438 1353 444 1354
rect 486 1353 492 1354
rect 526 1358 532 1359
rect 526 1354 527 1358
rect 531 1354 532 1358
rect 538 1355 539 1359
rect 543 1355 544 1359
rect 538 1354 544 1355
rect 566 1358 572 1359
rect 566 1354 567 1358
rect 571 1354 572 1358
rect 526 1353 532 1354
rect 566 1353 572 1354
rect 614 1358 620 1359
rect 614 1354 615 1358
rect 619 1354 620 1358
rect 626 1355 627 1359
rect 631 1355 632 1359
rect 626 1354 632 1355
rect 662 1358 668 1359
rect 662 1354 663 1358
rect 667 1354 668 1358
rect 614 1353 620 1354
rect 662 1353 668 1354
rect 710 1358 716 1359
rect 710 1354 711 1358
rect 715 1354 716 1358
rect 722 1355 723 1359
rect 727 1355 728 1359
rect 722 1354 728 1355
rect 766 1358 772 1359
rect 766 1354 767 1358
rect 771 1354 772 1358
rect 710 1353 716 1354
rect 766 1353 772 1354
rect 822 1358 828 1359
rect 822 1354 823 1358
rect 827 1354 828 1358
rect 834 1355 835 1359
rect 839 1355 840 1359
rect 834 1354 840 1355
rect 878 1358 884 1359
rect 878 1354 879 1358
rect 883 1354 884 1358
rect 822 1353 828 1354
rect 878 1353 884 1354
rect 934 1358 940 1359
rect 934 1354 935 1358
rect 939 1354 940 1358
rect 946 1355 947 1359
rect 951 1355 952 1359
rect 946 1354 952 1355
rect 990 1358 996 1359
rect 990 1354 991 1358
rect 995 1354 996 1358
rect 1002 1355 1003 1359
rect 1007 1355 1008 1359
rect 1002 1354 1008 1355
rect 934 1353 940 1354
rect 990 1353 996 1354
rect 206 1351 212 1352
rect 232 1351 234 1353
rect 280 1351 282 1353
rect 318 1351 324 1352
rect 336 1351 338 1353
rect 392 1351 394 1353
rect 440 1351 442 1353
rect 488 1351 490 1353
rect 494 1351 500 1352
rect 528 1351 530 1353
rect 568 1351 570 1353
rect 616 1351 618 1353
rect 664 1351 666 1353
rect 690 1351 696 1352
rect 712 1351 714 1353
rect 768 1351 770 1353
rect 824 1351 826 1353
rect 880 1351 882 1353
rect 936 1351 938 1353
rect 992 1351 994 1353
rect 111 1350 115 1351
rect 111 1345 115 1346
rect 135 1350 139 1351
rect 135 1345 139 1346
rect 159 1350 163 1351
rect 159 1345 163 1346
rect 167 1350 171 1351
rect 167 1345 171 1346
rect 183 1350 187 1351
rect 183 1345 187 1346
rect 191 1350 195 1351
rect 206 1347 207 1351
rect 211 1347 212 1351
rect 206 1346 212 1347
rect 231 1350 235 1351
rect 191 1345 195 1346
rect 231 1345 235 1346
rect 279 1350 283 1351
rect 318 1347 319 1351
rect 323 1347 324 1351
rect 318 1346 324 1347
rect 335 1350 339 1351
rect 279 1345 283 1346
rect 112 1338 114 1345
rect 168 1343 170 1345
rect 192 1343 194 1345
rect 232 1343 234 1345
rect 280 1343 282 1345
rect 166 1342 172 1343
rect 166 1338 167 1342
rect 171 1338 172 1342
rect 110 1337 116 1338
rect 166 1337 172 1338
rect 190 1342 196 1343
rect 190 1338 191 1342
rect 195 1338 196 1342
rect 190 1337 196 1338
rect 230 1342 236 1343
rect 230 1338 231 1342
rect 235 1338 236 1342
rect 230 1337 236 1338
rect 278 1342 284 1343
rect 278 1338 279 1342
rect 283 1338 284 1342
rect 278 1337 284 1338
rect 110 1333 111 1337
rect 115 1333 116 1337
rect 110 1332 116 1333
rect 320 1328 322 1346
rect 335 1345 339 1346
rect 391 1350 395 1351
rect 391 1345 395 1346
rect 439 1350 443 1351
rect 439 1345 443 1346
rect 455 1350 459 1351
rect 455 1345 459 1346
rect 487 1350 491 1351
rect 494 1347 495 1351
rect 499 1347 500 1351
rect 494 1346 500 1347
rect 519 1350 523 1351
rect 487 1345 491 1346
rect 336 1343 338 1345
rect 392 1343 394 1345
rect 456 1343 458 1345
rect 334 1342 340 1343
rect 334 1338 335 1342
rect 339 1338 340 1342
rect 334 1337 340 1338
rect 390 1342 396 1343
rect 390 1338 391 1342
rect 395 1338 396 1342
rect 454 1342 460 1343
rect 390 1337 396 1338
rect 410 1339 416 1340
rect 410 1335 411 1339
rect 415 1335 416 1339
rect 454 1338 455 1342
rect 459 1338 460 1342
rect 454 1337 460 1338
rect 410 1334 416 1335
rect 318 1327 324 1328
rect 243 1324 247 1325
rect 318 1323 319 1327
rect 323 1323 324 1327
rect 318 1322 324 1323
rect 326 1327 332 1328
rect 326 1322 327 1327
rect 110 1319 116 1320
rect 243 1319 247 1320
rect 331 1322 332 1327
rect 327 1319 331 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 110 1314 116 1315
rect 166 1316 172 1317
rect 112 1311 114 1314
rect 166 1312 167 1316
rect 171 1312 172 1316
rect 166 1311 172 1312
rect 190 1316 196 1317
rect 190 1312 191 1316
rect 195 1312 196 1316
rect 190 1311 196 1312
rect 230 1316 236 1317
rect 230 1312 231 1316
rect 235 1312 236 1316
rect 230 1311 236 1312
rect 111 1310 115 1311
rect 111 1305 115 1306
rect 167 1310 171 1311
rect 167 1305 171 1306
rect 191 1310 195 1311
rect 191 1305 195 1306
rect 231 1310 235 1311
rect 231 1305 235 1306
rect 112 1302 114 1305
rect 230 1304 236 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 230 1300 231 1304
rect 235 1300 236 1304
rect 230 1299 236 1300
rect 110 1296 116 1297
rect 110 1283 116 1284
rect 110 1279 111 1283
rect 115 1279 116 1283
rect 244 1280 246 1319
rect 278 1316 284 1317
rect 278 1312 279 1316
rect 283 1312 284 1316
rect 278 1311 284 1312
rect 334 1316 340 1317
rect 334 1312 335 1316
rect 339 1312 340 1316
rect 334 1311 340 1312
rect 390 1316 396 1317
rect 390 1312 391 1316
rect 395 1312 396 1316
rect 390 1311 396 1312
rect 255 1310 259 1311
rect 255 1305 259 1306
rect 279 1310 283 1311
rect 279 1305 283 1306
rect 303 1310 307 1311
rect 303 1305 307 1306
rect 327 1310 331 1311
rect 327 1305 331 1306
rect 335 1310 339 1311
rect 335 1305 339 1306
rect 351 1310 355 1311
rect 351 1305 355 1306
rect 375 1310 379 1311
rect 375 1305 379 1306
rect 391 1310 395 1311
rect 391 1305 395 1306
rect 399 1310 403 1311
rect 399 1305 403 1306
rect 254 1304 260 1305
rect 254 1300 255 1304
rect 259 1300 260 1304
rect 254 1299 260 1300
rect 278 1304 284 1305
rect 278 1300 279 1304
rect 283 1300 284 1304
rect 278 1299 284 1300
rect 302 1304 308 1305
rect 302 1300 303 1304
rect 307 1300 308 1304
rect 302 1299 308 1300
rect 326 1304 332 1305
rect 326 1300 327 1304
rect 331 1300 332 1304
rect 326 1299 332 1300
rect 350 1304 356 1305
rect 350 1300 351 1304
rect 355 1300 356 1304
rect 350 1299 356 1300
rect 374 1304 380 1305
rect 374 1300 375 1304
rect 379 1300 380 1304
rect 374 1299 380 1300
rect 398 1304 404 1305
rect 398 1300 399 1304
rect 403 1300 404 1304
rect 398 1299 404 1300
rect 412 1296 414 1334
rect 454 1316 460 1317
rect 454 1312 455 1316
rect 459 1312 460 1316
rect 496 1312 498 1346
rect 519 1345 523 1346
rect 527 1350 531 1351
rect 527 1345 531 1346
rect 567 1350 571 1351
rect 567 1345 571 1346
rect 575 1350 579 1351
rect 575 1345 579 1346
rect 615 1350 619 1351
rect 615 1345 619 1346
rect 631 1350 635 1351
rect 631 1345 635 1346
rect 663 1350 667 1351
rect 663 1345 667 1346
rect 679 1350 683 1351
rect 690 1347 691 1351
rect 695 1347 696 1351
rect 690 1346 696 1347
rect 711 1350 715 1351
rect 679 1345 683 1346
rect 520 1343 522 1345
rect 576 1343 578 1345
rect 632 1343 634 1345
rect 680 1343 682 1345
rect 518 1342 524 1343
rect 518 1338 519 1342
rect 523 1338 524 1342
rect 518 1337 524 1338
rect 574 1342 580 1343
rect 574 1338 575 1342
rect 579 1338 580 1342
rect 574 1337 580 1338
rect 630 1342 636 1343
rect 630 1338 631 1342
rect 635 1338 636 1342
rect 630 1337 636 1338
rect 678 1342 684 1343
rect 678 1338 679 1342
rect 683 1338 684 1342
rect 678 1337 684 1338
rect 692 1332 694 1346
rect 711 1345 715 1346
rect 727 1350 731 1351
rect 727 1345 731 1346
rect 767 1350 771 1351
rect 767 1345 771 1346
rect 799 1350 803 1351
rect 799 1345 803 1346
rect 823 1350 827 1351
rect 823 1345 827 1346
rect 831 1350 835 1351
rect 831 1345 835 1346
rect 863 1350 867 1351
rect 863 1345 867 1346
rect 879 1350 883 1351
rect 879 1345 883 1346
rect 895 1350 899 1351
rect 895 1345 899 1346
rect 927 1350 931 1351
rect 927 1345 931 1346
rect 935 1350 939 1351
rect 935 1345 939 1346
rect 967 1350 971 1351
rect 967 1345 971 1346
rect 991 1350 995 1351
rect 991 1345 995 1346
rect 1007 1350 1011 1351
rect 1007 1345 1011 1346
rect 728 1343 730 1345
rect 768 1343 770 1345
rect 800 1343 802 1345
rect 832 1343 834 1345
rect 864 1343 866 1345
rect 896 1343 898 1345
rect 928 1343 930 1345
rect 968 1343 970 1345
rect 1008 1343 1010 1345
rect 1020 1344 1022 1362
rect 1046 1358 1052 1359
rect 1046 1354 1047 1358
rect 1051 1354 1052 1358
rect 1046 1353 1052 1354
rect 1094 1358 1100 1359
rect 1094 1354 1095 1358
rect 1099 1354 1100 1358
rect 1142 1358 1148 1359
rect 1094 1353 1100 1354
rect 1114 1355 1120 1356
rect 1048 1351 1050 1353
rect 1096 1351 1098 1353
rect 1114 1351 1115 1355
rect 1119 1351 1120 1355
rect 1142 1354 1143 1358
rect 1147 1354 1148 1358
rect 1142 1353 1148 1354
rect 1144 1351 1146 1353
rect 1047 1350 1051 1351
rect 1047 1345 1051 1346
rect 1055 1350 1059 1351
rect 1055 1345 1059 1346
rect 1095 1350 1099 1351
rect 1095 1345 1099 1346
rect 1103 1350 1107 1351
rect 1114 1350 1120 1351
rect 1143 1350 1147 1351
rect 1103 1345 1107 1346
rect 1018 1343 1024 1344
rect 1056 1343 1058 1345
rect 1104 1343 1106 1345
rect 726 1342 732 1343
rect 726 1338 727 1342
rect 731 1338 732 1342
rect 726 1337 732 1338
rect 766 1342 772 1343
rect 766 1338 767 1342
rect 771 1338 772 1342
rect 766 1337 772 1338
rect 798 1342 804 1343
rect 798 1338 799 1342
rect 803 1338 804 1342
rect 798 1337 804 1338
rect 830 1342 836 1343
rect 830 1338 831 1342
rect 835 1338 836 1342
rect 830 1337 836 1338
rect 862 1342 868 1343
rect 862 1338 863 1342
rect 867 1338 868 1342
rect 862 1337 868 1338
rect 894 1342 900 1343
rect 894 1338 895 1342
rect 899 1338 900 1342
rect 894 1337 900 1338
rect 926 1342 932 1343
rect 926 1338 927 1342
rect 931 1338 932 1342
rect 926 1337 932 1338
rect 966 1342 972 1343
rect 966 1338 967 1342
rect 971 1338 972 1342
rect 1006 1342 1012 1343
rect 966 1337 972 1338
rect 978 1339 984 1340
rect 978 1335 979 1339
rect 983 1335 984 1339
rect 1006 1338 1007 1342
rect 1011 1338 1012 1342
rect 1018 1339 1019 1343
rect 1023 1339 1024 1343
rect 1018 1338 1024 1339
rect 1054 1342 1060 1343
rect 1054 1338 1055 1342
rect 1059 1338 1060 1342
rect 1006 1337 1012 1338
rect 1054 1337 1060 1338
rect 1102 1342 1108 1343
rect 1102 1338 1103 1342
rect 1107 1338 1108 1342
rect 1102 1337 1108 1338
rect 978 1334 984 1335
rect 690 1331 696 1332
rect 690 1327 691 1331
rect 695 1327 696 1331
rect 690 1326 696 1327
rect 518 1316 524 1317
rect 518 1312 519 1316
rect 523 1312 524 1316
rect 454 1311 460 1312
rect 494 1311 500 1312
rect 518 1311 524 1312
rect 574 1316 580 1317
rect 574 1312 575 1316
rect 579 1312 580 1316
rect 574 1311 580 1312
rect 630 1316 636 1317
rect 678 1316 684 1317
rect 630 1312 631 1316
rect 635 1312 636 1316
rect 630 1311 636 1312
rect 670 1315 676 1316
rect 670 1311 671 1315
rect 675 1311 676 1315
rect 678 1312 679 1316
rect 683 1312 684 1316
rect 678 1311 684 1312
rect 726 1316 732 1317
rect 726 1312 727 1316
rect 731 1312 732 1316
rect 726 1311 732 1312
rect 766 1316 772 1317
rect 766 1312 767 1316
rect 771 1312 772 1316
rect 766 1311 772 1312
rect 798 1316 804 1317
rect 798 1312 799 1316
rect 803 1312 804 1316
rect 798 1311 804 1312
rect 830 1316 836 1317
rect 830 1312 831 1316
rect 835 1312 836 1316
rect 830 1311 836 1312
rect 862 1316 868 1317
rect 862 1312 863 1316
rect 867 1312 868 1316
rect 862 1311 868 1312
rect 894 1316 900 1317
rect 894 1312 895 1316
rect 899 1312 900 1316
rect 894 1311 900 1312
rect 926 1316 932 1317
rect 926 1312 927 1316
rect 931 1312 932 1316
rect 926 1311 932 1312
rect 966 1316 972 1317
rect 966 1312 967 1316
rect 971 1312 972 1316
rect 966 1311 972 1312
rect 423 1310 427 1311
rect 423 1305 427 1306
rect 447 1310 451 1311
rect 447 1305 451 1306
rect 455 1310 459 1311
rect 455 1305 459 1306
rect 471 1310 475 1311
rect 494 1307 495 1311
rect 499 1307 500 1311
rect 494 1306 500 1307
rect 503 1310 507 1311
rect 471 1305 475 1306
rect 503 1305 507 1306
rect 519 1310 523 1311
rect 519 1305 523 1306
rect 543 1310 547 1311
rect 543 1305 547 1306
rect 575 1310 579 1311
rect 575 1305 579 1306
rect 591 1310 595 1311
rect 591 1305 595 1306
rect 631 1310 635 1311
rect 631 1305 635 1306
rect 647 1310 651 1311
rect 670 1310 676 1311
rect 679 1310 683 1311
rect 647 1305 651 1306
rect 422 1304 428 1305
rect 422 1300 423 1304
rect 427 1300 428 1304
rect 422 1299 428 1300
rect 446 1304 452 1305
rect 446 1300 447 1304
rect 451 1300 452 1304
rect 446 1299 452 1300
rect 470 1304 476 1305
rect 470 1300 471 1304
rect 475 1300 476 1304
rect 470 1299 476 1300
rect 502 1304 508 1305
rect 502 1300 503 1304
rect 507 1300 508 1304
rect 502 1299 508 1300
rect 542 1304 548 1305
rect 542 1300 543 1304
rect 547 1300 548 1304
rect 542 1299 548 1300
rect 590 1304 596 1305
rect 590 1300 591 1304
rect 595 1300 596 1304
rect 590 1299 596 1300
rect 646 1304 652 1305
rect 646 1300 647 1304
rect 651 1300 652 1304
rect 646 1299 652 1300
rect 266 1295 272 1296
rect 266 1291 267 1295
rect 271 1291 272 1295
rect 266 1290 272 1291
rect 338 1295 344 1296
rect 338 1291 339 1295
rect 343 1291 344 1295
rect 338 1290 344 1291
rect 410 1295 416 1296
rect 410 1291 411 1295
rect 415 1291 416 1295
rect 410 1290 416 1291
rect 268 1280 270 1290
rect 318 1287 324 1288
rect 318 1283 319 1287
rect 323 1283 324 1287
rect 318 1282 324 1283
rect 242 1279 248 1280
rect 266 1279 272 1280
rect 110 1278 116 1279
rect 230 1278 236 1279
rect 112 1271 114 1278
rect 230 1274 231 1278
rect 235 1274 236 1278
rect 242 1275 243 1279
rect 247 1275 248 1279
rect 242 1274 248 1275
rect 254 1278 260 1279
rect 254 1274 255 1278
rect 259 1274 260 1278
rect 266 1275 267 1279
rect 271 1275 272 1279
rect 266 1274 272 1275
rect 278 1278 284 1279
rect 278 1274 279 1278
rect 283 1274 284 1278
rect 230 1273 236 1274
rect 254 1273 260 1274
rect 278 1273 284 1274
rect 302 1278 308 1279
rect 302 1274 303 1278
rect 307 1274 308 1278
rect 302 1273 308 1274
rect 232 1271 234 1273
rect 256 1271 258 1273
rect 280 1271 282 1273
rect 304 1271 306 1273
rect 111 1270 115 1271
rect 111 1265 115 1266
rect 231 1270 235 1271
rect 231 1265 235 1266
rect 255 1270 259 1271
rect 255 1265 259 1266
rect 279 1270 283 1271
rect 279 1265 283 1266
rect 303 1270 307 1271
rect 303 1265 307 1266
rect 311 1270 315 1271
rect 320 1268 322 1282
rect 340 1280 342 1290
rect 672 1288 674 1310
rect 679 1305 683 1306
rect 695 1310 699 1311
rect 695 1305 699 1306
rect 727 1310 731 1311
rect 727 1305 731 1306
rect 743 1310 747 1311
rect 743 1305 747 1306
rect 767 1310 771 1311
rect 767 1305 771 1306
rect 791 1310 795 1311
rect 791 1305 795 1306
rect 799 1310 803 1311
rect 799 1305 803 1306
rect 831 1310 835 1311
rect 831 1305 835 1306
rect 839 1310 843 1311
rect 839 1305 843 1306
rect 863 1310 867 1311
rect 863 1305 867 1306
rect 879 1310 883 1311
rect 879 1305 883 1306
rect 895 1310 899 1311
rect 895 1305 899 1306
rect 911 1310 915 1311
rect 911 1305 915 1306
rect 927 1310 931 1311
rect 927 1305 931 1306
rect 951 1310 955 1311
rect 951 1305 955 1306
rect 967 1310 971 1311
rect 967 1305 971 1306
rect 694 1304 700 1305
rect 694 1300 695 1304
rect 699 1300 700 1304
rect 694 1299 700 1300
rect 742 1304 748 1305
rect 742 1300 743 1304
rect 747 1300 748 1304
rect 742 1299 748 1300
rect 790 1304 796 1305
rect 790 1300 791 1304
rect 795 1300 796 1304
rect 790 1299 796 1300
rect 838 1304 844 1305
rect 838 1300 839 1304
rect 843 1300 844 1304
rect 838 1299 844 1300
rect 878 1304 884 1305
rect 878 1300 879 1304
rect 883 1300 884 1304
rect 878 1299 884 1300
rect 910 1304 916 1305
rect 910 1300 911 1304
rect 915 1300 916 1304
rect 910 1299 916 1300
rect 950 1304 956 1305
rect 950 1300 951 1304
rect 955 1300 956 1304
rect 950 1299 956 1300
rect 980 1296 982 1334
rect 1116 1332 1118 1350
rect 1143 1345 1147 1346
rect 1159 1350 1163 1351
rect 1159 1345 1163 1346
rect 1160 1343 1162 1345
rect 1172 1344 1174 1362
rect 1190 1358 1196 1359
rect 1190 1354 1191 1358
rect 1195 1354 1196 1358
rect 1190 1353 1196 1354
rect 1192 1351 1194 1353
rect 1208 1352 1210 1390
rect 1215 1385 1219 1386
rect 1239 1390 1243 1391
rect 1239 1385 1243 1386
rect 1263 1390 1267 1391
rect 1263 1385 1267 1386
rect 1287 1390 1291 1391
rect 1287 1385 1291 1386
rect 1303 1390 1307 1391
rect 1303 1385 1307 1386
rect 1238 1384 1244 1385
rect 1238 1380 1239 1384
rect 1243 1380 1244 1384
rect 1238 1379 1244 1380
rect 1286 1384 1292 1385
rect 1316 1384 1318 1414
rect 1356 1404 1358 1426
rect 1391 1425 1395 1426
rect 1415 1430 1419 1431
rect 1415 1425 1419 1426
rect 1447 1430 1451 1431
rect 1447 1425 1451 1426
rect 1392 1423 1394 1425
rect 1416 1423 1418 1425
rect 1390 1422 1396 1423
rect 1390 1418 1391 1422
rect 1395 1418 1396 1422
rect 1390 1417 1396 1418
rect 1414 1422 1420 1423
rect 1414 1418 1415 1422
rect 1419 1418 1420 1422
rect 1448 1418 1450 1425
rect 1414 1417 1420 1418
rect 1446 1417 1452 1418
rect 1446 1413 1447 1417
rect 1451 1413 1452 1417
rect 1446 1412 1452 1413
rect 1354 1403 1360 1404
rect 1354 1399 1355 1403
rect 1359 1399 1360 1403
rect 1354 1398 1360 1399
rect 1446 1399 1452 1400
rect 1342 1396 1348 1397
rect 1342 1392 1343 1396
rect 1347 1392 1348 1396
rect 1342 1391 1348 1392
rect 1390 1396 1396 1397
rect 1390 1392 1391 1396
rect 1395 1392 1396 1396
rect 1390 1391 1396 1392
rect 1414 1396 1420 1397
rect 1414 1392 1415 1396
rect 1419 1392 1420 1396
rect 1414 1391 1420 1392
rect 1426 1395 1432 1396
rect 1426 1391 1427 1395
rect 1431 1391 1432 1395
rect 1446 1395 1447 1399
rect 1451 1395 1452 1399
rect 1446 1394 1452 1395
rect 1448 1391 1450 1394
rect 1335 1390 1339 1391
rect 1335 1385 1339 1386
rect 1343 1390 1347 1391
rect 1343 1385 1347 1386
rect 1383 1390 1387 1391
rect 1383 1385 1387 1386
rect 1391 1390 1395 1391
rect 1391 1385 1395 1386
rect 1415 1390 1419 1391
rect 1426 1390 1432 1391
rect 1447 1390 1451 1391
rect 1415 1385 1419 1386
rect 1334 1384 1340 1385
rect 1286 1380 1287 1384
rect 1291 1380 1292 1384
rect 1286 1379 1292 1380
rect 1314 1383 1320 1384
rect 1314 1379 1315 1383
rect 1319 1379 1320 1383
rect 1334 1380 1335 1384
rect 1339 1380 1340 1384
rect 1334 1379 1340 1380
rect 1382 1384 1388 1385
rect 1382 1380 1383 1384
rect 1387 1380 1388 1384
rect 1382 1379 1388 1380
rect 1414 1384 1420 1385
rect 1414 1380 1415 1384
rect 1419 1380 1420 1384
rect 1414 1379 1420 1380
rect 1314 1378 1320 1379
rect 1428 1376 1430 1390
rect 1447 1385 1451 1386
rect 1448 1382 1450 1385
rect 1446 1381 1452 1382
rect 1446 1377 1447 1381
rect 1451 1377 1452 1381
rect 1446 1376 1452 1377
rect 1394 1375 1400 1376
rect 1394 1371 1395 1375
rect 1399 1371 1400 1375
rect 1394 1370 1400 1371
rect 1426 1375 1432 1376
rect 1426 1371 1427 1375
rect 1431 1371 1432 1375
rect 1426 1370 1432 1371
rect 1396 1360 1398 1370
rect 1426 1367 1432 1368
rect 1426 1363 1427 1367
rect 1431 1363 1432 1367
rect 1426 1362 1432 1363
rect 1446 1363 1452 1364
rect 1394 1359 1400 1360
rect 1238 1358 1244 1359
rect 1238 1354 1239 1358
rect 1243 1354 1244 1358
rect 1238 1353 1244 1354
rect 1286 1358 1292 1359
rect 1286 1354 1287 1358
rect 1291 1354 1292 1358
rect 1286 1353 1292 1354
rect 1334 1358 1340 1359
rect 1334 1354 1335 1358
rect 1339 1354 1340 1358
rect 1382 1358 1388 1359
rect 1334 1353 1340 1354
rect 1374 1355 1380 1356
rect 1206 1351 1212 1352
rect 1240 1351 1242 1353
rect 1288 1351 1290 1353
rect 1336 1351 1338 1353
rect 1374 1351 1375 1355
rect 1379 1351 1380 1355
rect 1382 1354 1383 1358
rect 1387 1354 1388 1358
rect 1394 1355 1395 1359
rect 1399 1355 1400 1359
rect 1394 1354 1400 1355
rect 1414 1358 1420 1359
rect 1414 1354 1415 1358
rect 1419 1354 1420 1358
rect 1382 1353 1388 1354
rect 1414 1353 1420 1354
rect 1384 1351 1386 1353
rect 1416 1351 1418 1353
rect 1191 1350 1195 1351
rect 1206 1347 1207 1351
rect 1211 1347 1212 1351
rect 1206 1346 1212 1347
rect 1215 1350 1219 1351
rect 1191 1345 1195 1346
rect 1215 1345 1219 1346
rect 1239 1350 1243 1351
rect 1239 1345 1243 1346
rect 1271 1350 1275 1351
rect 1271 1345 1275 1346
rect 1287 1350 1291 1351
rect 1287 1345 1291 1346
rect 1327 1350 1331 1351
rect 1327 1345 1331 1346
rect 1335 1350 1339 1351
rect 1374 1350 1380 1351
rect 1383 1350 1387 1351
rect 1335 1345 1339 1346
rect 1170 1343 1176 1344
rect 1216 1343 1218 1345
rect 1272 1343 1274 1345
rect 1328 1343 1330 1345
rect 1158 1342 1164 1343
rect 1122 1339 1128 1340
rect 1122 1335 1123 1339
rect 1127 1335 1128 1339
rect 1158 1338 1159 1342
rect 1163 1338 1164 1342
rect 1170 1339 1171 1343
rect 1175 1339 1176 1343
rect 1170 1338 1176 1339
rect 1214 1342 1220 1343
rect 1214 1338 1215 1342
rect 1219 1338 1220 1342
rect 1158 1337 1164 1338
rect 1214 1337 1220 1338
rect 1270 1342 1276 1343
rect 1270 1338 1271 1342
rect 1275 1338 1276 1342
rect 1326 1342 1332 1343
rect 1270 1337 1276 1338
rect 1314 1339 1320 1340
rect 1122 1334 1128 1335
rect 1314 1335 1315 1339
rect 1319 1335 1320 1339
rect 1326 1338 1327 1342
rect 1331 1338 1332 1342
rect 1326 1337 1332 1338
rect 1314 1334 1320 1335
rect 1114 1331 1120 1332
rect 1114 1327 1115 1331
rect 1119 1327 1120 1331
rect 1114 1326 1120 1327
rect 1006 1316 1012 1317
rect 1006 1312 1007 1316
rect 1011 1312 1012 1316
rect 1006 1311 1012 1312
rect 1054 1316 1060 1317
rect 1102 1316 1108 1317
rect 1054 1312 1055 1316
rect 1059 1312 1060 1316
rect 1054 1311 1060 1312
rect 1082 1315 1088 1316
rect 1082 1311 1083 1315
rect 1087 1311 1088 1315
rect 1102 1312 1103 1316
rect 1107 1312 1108 1316
rect 1102 1311 1108 1312
rect 991 1310 995 1311
rect 991 1305 995 1306
rect 1007 1310 1011 1311
rect 1007 1305 1011 1306
rect 1031 1310 1035 1311
rect 1031 1305 1035 1306
rect 1055 1310 1059 1311
rect 1055 1305 1059 1306
rect 1071 1310 1075 1311
rect 1082 1310 1088 1311
rect 1103 1310 1107 1311
rect 1071 1305 1075 1306
rect 990 1304 996 1305
rect 990 1300 991 1304
rect 995 1300 996 1304
rect 990 1299 996 1300
rect 1030 1304 1036 1305
rect 1030 1300 1031 1304
rect 1035 1300 1036 1304
rect 1030 1299 1036 1300
rect 1070 1304 1076 1305
rect 1070 1300 1071 1304
rect 1075 1300 1076 1304
rect 1070 1299 1076 1300
rect 754 1295 760 1296
rect 754 1291 755 1295
rect 759 1291 760 1295
rect 754 1290 760 1291
rect 978 1295 984 1296
rect 978 1291 979 1295
rect 983 1291 984 1295
rect 978 1290 984 1291
rect 670 1287 676 1288
rect 670 1283 671 1287
rect 675 1283 676 1287
rect 670 1282 676 1283
rect 756 1280 758 1290
rect 1084 1280 1086 1310
rect 1103 1305 1107 1306
rect 1111 1310 1115 1311
rect 1111 1305 1115 1306
rect 1110 1304 1116 1305
rect 1124 1304 1126 1334
rect 1158 1316 1164 1317
rect 1158 1312 1159 1316
rect 1163 1312 1164 1316
rect 1158 1311 1164 1312
rect 1214 1316 1220 1317
rect 1270 1316 1276 1317
rect 1214 1312 1215 1316
rect 1219 1312 1220 1316
rect 1214 1311 1220 1312
rect 1258 1315 1264 1316
rect 1258 1311 1259 1315
rect 1263 1311 1264 1315
rect 1270 1312 1271 1316
rect 1275 1312 1276 1316
rect 1270 1311 1276 1312
rect 1151 1310 1155 1311
rect 1151 1305 1155 1306
rect 1159 1310 1163 1311
rect 1159 1305 1163 1306
rect 1199 1310 1203 1311
rect 1199 1305 1203 1306
rect 1215 1310 1219 1311
rect 1215 1305 1219 1306
rect 1247 1310 1251 1311
rect 1258 1310 1264 1311
rect 1271 1310 1275 1311
rect 1247 1305 1251 1306
rect 1150 1304 1156 1305
rect 1110 1300 1111 1304
rect 1115 1300 1116 1304
rect 1110 1299 1116 1300
rect 1122 1303 1128 1304
rect 1122 1299 1123 1303
rect 1127 1299 1128 1303
rect 1150 1300 1151 1304
rect 1155 1300 1156 1304
rect 1150 1299 1156 1300
rect 1198 1304 1204 1305
rect 1198 1300 1199 1304
rect 1203 1300 1204 1304
rect 1198 1299 1204 1300
rect 1246 1304 1252 1305
rect 1246 1300 1247 1304
rect 1251 1300 1252 1304
rect 1246 1299 1252 1300
rect 1122 1298 1128 1299
rect 1138 1287 1144 1288
rect 1138 1283 1139 1287
rect 1143 1283 1144 1287
rect 1138 1282 1144 1283
rect 338 1279 344 1280
rect 362 1279 368 1280
rect 754 1279 760 1280
rect 1082 1279 1088 1280
rect 326 1278 332 1279
rect 326 1274 327 1278
rect 331 1274 332 1278
rect 338 1275 339 1279
rect 343 1275 344 1279
rect 338 1274 344 1275
rect 350 1278 356 1279
rect 350 1274 351 1278
rect 355 1274 356 1278
rect 362 1275 363 1279
rect 367 1275 368 1279
rect 374 1278 380 1279
rect 362 1274 370 1275
rect 326 1273 332 1274
rect 350 1273 356 1274
rect 364 1273 370 1274
rect 374 1274 375 1278
rect 379 1274 380 1278
rect 374 1273 380 1274
rect 398 1278 404 1279
rect 398 1274 399 1278
rect 403 1274 404 1278
rect 398 1273 404 1274
rect 422 1278 428 1279
rect 422 1274 423 1278
rect 427 1274 428 1278
rect 422 1273 428 1274
rect 446 1278 452 1279
rect 446 1274 447 1278
rect 451 1274 452 1278
rect 446 1273 452 1274
rect 470 1278 476 1279
rect 470 1274 471 1278
rect 475 1274 476 1278
rect 470 1273 476 1274
rect 502 1278 508 1279
rect 502 1274 503 1278
rect 507 1274 508 1278
rect 502 1273 508 1274
rect 542 1278 548 1279
rect 542 1274 543 1278
rect 547 1274 548 1278
rect 542 1273 548 1274
rect 590 1278 596 1279
rect 590 1274 591 1278
rect 595 1274 596 1278
rect 590 1273 596 1274
rect 646 1278 652 1279
rect 646 1274 647 1278
rect 651 1274 652 1278
rect 646 1273 652 1274
rect 694 1278 700 1279
rect 694 1274 695 1278
rect 699 1274 700 1278
rect 694 1273 700 1274
rect 742 1278 748 1279
rect 742 1274 743 1278
rect 747 1274 748 1278
rect 754 1275 755 1279
rect 759 1275 760 1279
rect 754 1274 760 1275
rect 790 1278 796 1279
rect 790 1274 791 1278
rect 795 1274 796 1278
rect 742 1273 748 1274
rect 790 1273 796 1274
rect 838 1278 844 1279
rect 838 1274 839 1278
rect 843 1274 844 1278
rect 838 1273 844 1274
rect 878 1278 884 1279
rect 878 1274 879 1278
rect 883 1274 884 1278
rect 878 1273 884 1274
rect 910 1278 916 1279
rect 910 1274 911 1278
rect 915 1274 916 1278
rect 910 1273 916 1274
rect 950 1278 956 1279
rect 950 1274 951 1278
rect 955 1274 956 1278
rect 950 1273 956 1274
rect 990 1278 996 1279
rect 990 1274 991 1278
rect 995 1274 996 1278
rect 990 1273 996 1274
rect 1030 1278 1036 1279
rect 1030 1274 1031 1278
rect 1035 1274 1036 1278
rect 1030 1273 1036 1274
rect 1070 1278 1076 1279
rect 1070 1274 1071 1278
rect 1075 1274 1076 1278
rect 1082 1275 1083 1279
rect 1087 1275 1088 1279
rect 1082 1274 1088 1275
rect 1110 1278 1116 1279
rect 1110 1274 1111 1278
rect 1115 1274 1116 1278
rect 1070 1273 1076 1274
rect 1110 1273 1116 1274
rect 328 1271 330 1273
rect 342 1271 348 1272
rect 352 1271 354 1273
rect 327 1270 331 1271
rect 311 1265 315 1266
rect 318 1267 324 1268
rect 112 1258 114 1265
rect 312 1263 314 1265
rect 318 1263 319 1267
rect 323 1263 324 1267
rect 327 1265 331 1266
rect 335 1270 339 1271
rect 342 1267 343 1271
rect 347 1267 348 1271
rect 342 1266 348 1267
rect 351 1270 355 1271
rect 335 1265 339 1266
rect 336 1263 338 1265
rect 310 1262 316 1263
rect 318 1262 324 1263
rect 334 1262 340 1263
rect 310 1258 311 1262
rect 315 1258 316 1262
rect 110 1257 116 1258
rect 310 1257 316 1258
rect 334 1258 335 1262
rect 339 1258 340 1262
rect 334 1257 340 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 110 1252 116 1253
rect 344 1244 346 1266
rect 351 1265 355 1266
rect 359 1270 363 1271
rect 359 1265 363 1266
rect 360 1263 362 1265
rect 358 1262 364 1263
rect 358 1258 359 1262
rect 363 1258 364 1262
rect 358 1257 364 1258
rect 368 1252 370 1273
rect 376 1271 378 1273
rect 400 1271 402 1273
rect 424 1271 426 1273
rect 448 1271 450 1273
rect 472 1271 474 1273
rect 504 1271 506 1273
rect 530 1271 536 1272
rect 544 1271 546 1273
rect 592 1271 594 1273
rect 648 1271 650 1273
rect 696 1271 698 1273
rect 744 1271 746 1273
rect 792 1271 794 1273
rect 840 1271 842 1273
rect 880 1271 882 1273
rect 912 1271 914 1273
rect 952 1271 954 1273
rect 992 1271 994 1273
rect 1002 1271 1008 1272
rect 1032 1271 1034 1273
rect 1072 1271 1074 1273
rect 1112 1271 1114 1273
rect 375 1270 379 1271
rect 375 1265 379 1266
rect 383 1270 387 1271
rect 383 1265 387 1266
rect 399 1270 403 1271
rect 399 1265 403 1266
rect 415 1270 419 1271
rect 415 1265 419 1266
rect 423 1270 427 1271
rect 423 1265 427 1266
rect 447 1270 451 1271
rect 447 1265 451 1266
rect 471 1270 475 1271
rect 471 1265 475 1266
rect 479 1270 483 1271
rect 479 1265 483 1266
rect 503 1270 507 1271
rect 503 1265 507 1266
rect 519 1270 523 1271
rect 530 1267 531 1271
rect 535 1267 536 1271
rect 530 1266 536 1267
rect 543 1270 547 1271
rect 519 1265 523 1266
rect 384 1263 386 1265
rect 416 1263 418 1265
rect 448 1263 450 1265
rect 480 1263 482 1265
rect 520 1263 522 1265
rect 382 1262 388 1263
rect 382 1258 383 1262
rect 387 1258 388 1262
rect 382 1257 388 1258
rect 414 1262 420 1263
rect 414 1258 415 1262
rect 419 1258 420 1262
rect 414 1257 420 1258
rect 446 1262 452 1263
rect 446 1258 447 1262
rect 451 1258 452 1262
rect 446 1257 452 1258
rect 478 1262 484 1263
rect 478 1258 479 1262
rect 483 1258 484 1262
rect 478 1257 484 1258
rect 518 1262 524 1263
rect 518 1258 519 1262
rect 523 1258 524 1262
rect 518 1257 524 1258
rect 366 1251 372 1252
rect 366 1247 367 1251
rect 371 1247 372 1251
rect 366 1246 372 1247
rect 532 1244 534 1266
rect 543 1265 547 1266
rect 559 1270 563 1271
rect 559 1265 563 1266
rect 591 1270 595 1271
rect 591 1265 595 1266
rect 615 1270 619 1271
rect 615 1265 619 1266
rect 647 1270 651 1271
rect 647 1265 651 1266
rect 679 1270 683 1271
rect 679 1265 683 1266
rect 695 1270 699 1271
rect 695 1265 699 1266
rect 743 1270 747 1271
rect 743 1265 747 1266
rect 751 1270 755 1271
rect 751 1265 755 1266
rect 791 1270 795 1271
rect 791 1265 795 1266
rect 831 1270 835 1271
rect 831 1265 835 1266
rect 839 1270 843 1271
rect 839 1265 843 1266
rect 879 1270 883 1271
rect 879 1265 883 1266
rect 911 1270 915 1271
rect 911 1265 915 1266
rect 951 1270 955 1271
rect 951 1265 955 1266
rect 991 1270 995 1271
rect 1002 1267 1003 1271
rect 1007 1267 1008 1271
rect 1002 1266 1008 1267
rect 1031 1270 1035 1271
rect 991 1265 995 1266
rect 560 1263 562 1265
rect 616 1263 618 1265
rect 680 1263 682 1265
rect 752 1263 754 1265
rect 832 1263 834 1265
rect 912 1263 914 1265
rect 992 1263 994 1265
rect 558 1262 564 1263
rect 558 1258 559 1262
rect 563 1258 564 1262
rect 558 1257 564 1258
rect 614 1262 620 1263
rect 614 1258 615 1262
rect 619 1258 620 1262
rect 614 1257 620 1258
rect 678 1262 684 1263
rect 678 1258 679 1262
rect 683 1258 684 1262
rect 750 1262 756 1263
rect 678 1257 684 1258
rect 690 1259 696 1260
rect 690 1255 691 1259
rect 695 1255 696 1259
rect 750 1258 751 1262
rect 755 1258 756 1262
rect 750 1257 756 1258
rect 830 1262 836 1263
rect 830 1258 831 1262
rect 835 1258 836 1262
rect 830 1257 836 1258
rect 910 1262 916 1263
rect 910 1258 911 1262
rect 915 1258 916 1262
rect 910 1257 916 1258
rect 990 1262 996 1263
rect 990 1258 991 1262
rect 995 1258 996 1262
rect 990 1257 996 1258
rect 690 1254 696 1255
rect 344 1243 352 1244
rect 344 1241 347 1243
rect 110 1239 116 1240
rect 110 1235 111 1239
rect 115 1235 116 1239
rect 346 1239 347 1241
rect 351 1239 352 1243
rect 346 1238 352 1239
rect 530 1243 536 1244
rect 530 1239 531 1243
rect 535 1239 536 1243
rect 530 1238 536 1239
rect 110 1234 116 1235
rect 310 1236 316 1237
rect 112 1231 114 1234
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 334 1236 340 1237
rect 334 1232 335 1236
rect 339 1232 340 1236
rect 334 1231 340 1232
rect 358 1236 364 1237
rect 358 1232 359 1236
rect 363 1232 364 1236
rect 358 1231 364 1232
rect 382 1236 388 1237
rect 382 1232 383 1236
rect 387 1232 388 1236
rect 382 1231 388 1232
rect 414 1236 420 1237
rect 414 1232 415 1236
rect 419 1232 420 1236
rect 414 1231 420 1232
rect 446 1236 452 1237
rect 446 1232 447 1236
rect 451 1232 452 1236
rect 446 1231 452 1232
rect 478 1236 484 1237
rect 478 1232 479 1236
rect 483 1232 484 1236
rect 478 1231 484 1232
rect 518 1236 524 1237
rect 518 1232 519 1236
rect 523 1232 524 1236
rect 518 1231 524 1232
rect 558 1236 564 1237
rect 558 1232 559 1236
rect 563 1232 564 1236
rect 558 1231 564 1232
rect 614 1236 620 1237
rect 614 1232 615 1236
rect 619 1232 620 1236
rect 614 1231 620 1232
rect 678 1236 684 1237
rect 678 1232 679 1236
rect 683 1232 684 1236
rect 678 1231 684 1232
rect 111 1230 115 1231
rect 111 1225 115 1226
rect 311 1230 315 1231
rect 311 1225 315 1226
rect 327 1230 331 1231
rect 327 1225 331 1226
rect 335 1230 339 1231
rect 335 1225 339 1226
rect 359 1230 363 1231
rect 359 1225 363 1226
rect 367 1230 371 1231
rect 367 1225 371 1226
rect 383 1230 387 1231
rect 383 1225 387 1226
rect 407 1230 411 1231
rect 407 1225 411 1226
rect 415 1230 419 1231
rect 415 1225 419 1226
rect 447 1230 451 1231
rect 447 1225 451 1226
rect 479 1230 483 1231
rect 479 1225 483 1226
rect 487 1230 491 1231
rect 487 1225 491 1226
rect 519 1230 523 1231
rect 519 1225 523 1226
rect 527 1230 531 1231
rect 527 1225 531 1226
rect 559 1230 563 1231
rect 559 1225 563 1226
rect 567 1230 571 1231
rect 567 1225 571 1226
rect 607 1230 611 1231
rect 607 1225 611 1226
rect 615 1230 619 1231
rect 615 1225 619 1226
rect 655 1230 659 1231
rect 655 1225 659 1226
rect 679 1230 683 1231
rect 679 1225 683 1226
rect 112 1222 114 1225
rect 326 1224 332 1225
rect 110 1221 116 1222
rect 110 1217 111 1221
rect 115 1217 116 1221
rect 326 1220 327 1224
rect 331 1220 332 1224
rect 326 1219 332 1220
rect 366 1224 372 1225
rect 366 1220 367 1224
rect 371 1220 372 1224
rect 366 1219 372 1220
rect 406 1224 412 1225
rect 406 1220 407 1224
rect 411 1220 412 1224
rect 406 1219 412 1220
rect 446 1224 452 1225
rect 446 1220 447 1224
rect 451 1220 452 1224
rect 446 1219 452 1220
rect 486 1224 492 1225
rect 486 1220 487 1224
rect 491 1220 492 1224
rect 486 1219 492 1220
rect 526 1224 532 1225
rect 526 1220 527 1224
rect 531 1220 532 1224
rect 526 1219 532 1220
rect 566 1224 572 1225
rect 566 1220 567 1224
rect 571 1220 572 1224
rect 566 1219 572 1220
rect 606 1224 612 1225
rect 606 1220 607 1224
rect 611 1220 612 1224
rect 606 1219 612 1220
rect 654 1224 660 1225
rect 654 1220 655 1224
rect 659 1220 660 1224
rect 654 1219 660 1220
rect 110 1216 116 1217
rect 692 1216 694 1254
rect 1004 1252 1006 1266
rect 1031 1265 1035 1266
rect 1063 1270 1067 1271
rect 1063 1265 1067 1266
rect 1071 1270 1075 1271
rect 1071 1265 1075 1266
rect 1111 1270 1115 1271
rect 1111 1265 1115 1266
rect 1127 1270 1131 1271
rect 1127 1265 1131 1266
rect 1064 1263 1066 1265
rect 1128 1263 1130 1265
rect 1140 1264 1142 1282
rect 1260 1280 1262 1310
rect 1271 1305 1275 1306
rect 1303 1310 1307 1311
rect 1303 1305 1307 1306
rect 1302 1304 1308 1305
rect 1316 1304 1318 1334
rect 1326 1316 1332 1317
rect 1326 1312 1327 1316
rect 1331 1312 1332 1316
rect 1376 1312 1378 1350
rect 1383 1345 1387 1346
rect 1415 1350 1419 1351
rect 1415 1345 1419 1346
rect 1384 1343 1386 1345
rect 1416 1343 1418 1345
rect 1428 1344 1430 1362
rect 1446 1359 1447 1363
rect 1451 1359 1452 1363
rect 1446 1358 1452 1359
rect 1448 1351 1450 1358
rect 1447 1350 1451 1351
rect 1447 1345 1451 1346
rect 1426 1343 1432 1344
rect 1382 1342 1388 1343
rect 1382 1338 1383 1342
rect 1387 1338 1388 1342
rect 1382 1337 1388 1338
rect 1414 1342 1420 1343
rect 1414 1338 1415 1342
rect 1419 1338 1420 1342
rect 1426 1339 1427 1343
rect 1431 1339 1432 1343
rect 1426 1338 1432 1339
rect 1448 1338 1450 1345
rect 1414 1337 1420 1338
rect 1446 1337 1452 1338
rect 1446 1333 1447 1337
rect 1451 1333 1452 1337
rect 1446 1332 1452 1333
rect 1446 1319 1452 1320
rect 1382 1316 1388 1317
rect 1382 1312 1383 1316
rect 1387 1312 1388 1316
rect 1326 1311 1332 1312
rect 1374 1311 1380 1312
rect 1382 1311 1388 1312
rect 1414 1316 1420 1317
rect 1414 1312 1415 1316
rect 1419 1312 1420 1316
rect 1414 1311 1420 1312
rect 1426 1315 1432 1316
rect 1426 1311 1427 1315
rect 1431 1311 1432 1315
rect 1446 1315 1447 1319
rect 1451 1315 1452 1319
rect 1446 1314 1452 1315
rect 1448 1311 1450 1314
rect 1327 1310 1331 1311
rect 1327 1305 1331 1306
rect 1367 1310 1371 1311
rect 1374 1307 1375 1311
rect 1379 1307 1380 1311
rect 1374 1306 1380 1307
rect 1383 1310 1387 1311
rect 1367 1305 1371 1306
rect 1383 1305 1387 1306
rect 1415 1310 1419 1311
rect 1426 1310 1432 1311
rect 1447 1310 1451 1311
rect 1415 1305 1419 1306
rect 1366 1304 1372 1305
rect 1302 1300 1303 1304
rect 1307 1300 1308 1304
rect 1302 1299 1308 1300
rect 1314 1303 1320 1304
rect 1314 1299 1315 1303
rect 1319 1299 1320 1303
rect 1366 1300 1367 1304
rect 1371 1300 1372 1304
rect 1366 1299 1372 1300
rect 1414 1304 1420 1305
rect 1414 1300 1415 1304
rect 1419 1300 1420 1304
rect 1414 1299 1420 1300
rect 1314 1298 1320 1299
rect 1386 1287 1392 1288
rect 1386 1283 1387 1287
rect 1391 1283 1392 1287
rect 1386 1282 1392 1283
rect 1258 1279 1264 1280
rect 1150 1278 1156 1279
rect 1150 1274 1151 1278
rect 1155 1274 1156 1278
rect 1150 1273 1156 1274
rect 1198 1278 1204 1279
rect 1198 1274 1199 1278
rect 1203 1274 1204 1278
rect 1198 1273 1204 1274
rect 1246 1278 1252 1279
rect 1246 1274 1247 1278
rect 1251 1274 1252 1278
rect 1258 1275 1259 1279
rect 1263 1275 1264 1279
rect 1258 1274 1264 1275
rect 1302 1278 1308 1279
rect 1302 1274 1303 1278
rect 1307 1274 1308 1278
rect 1246 1273 1252 1274
rect 1302 1273 1308 1274
rect 1366 1278 1372 1279
rect 1366 1274 1367 1278
rect 1371 1274 1372 1278
rect 1366 1273 1372 1274
rect 1152 1271 1154 1273
rect 1200 1271 1202 1273
rect 1248 1271 1250 1273
rect 1294 1271 1300 1272
rect 1304 1271 1306 1273
rect 1322 1271 1328 1272
rect 1368 1271 1370 1273
rect 1151 1270 1155 1271
rect 1151 1265 1155 1266
rect 1191 1270 1195 1271
rect 1191 1265 1195 1266
rect 1199 1270 1203 1271
rect 1199 1265 1203 1266
rect 1247 1270 1251 1271
rect 1294 1267 1295 1271
rect 1299 1267 1300 1271
rect 1294 1266 1300 1267
rect 1303 1270 1307 1271
rect 1247 1265 1251 1266
rect 1138 1263 1144 1264
rect 1192 1263 1194 1265
rect 1248 1263 1250 1265
rect 1062 1262 1068 1263
rect 1062 1258 1063 1262
rect 1067 1258 1068 1262
rect 1062 1257 1068 1258
rect 1126 1262 1132 1263
rect 1126 1258 1127 1262
rect 1131 1258 1132 1262
rect 1138 1259 1139 1263
rect 1143 1259 1144 1263
rect 1138 1258 1144 1259
rect 1190 1262 1196 1263
rect 1190 1258 1191 1262
rect 1195 1258 1196 1262
rect 1126 1257 1132 1258
rect 1190 1257 1196 1258
rect 1246 1262 1252 1263
rect 1246 1258 1247 1262
rect 1251 1258 1252 1262
rect 1246 1257 1252 1258
rect 1002 1251 1008 1252
rect 1002 1247 1003 1251
rect 1007 1247 1008 1251
rect 1002 1246 1008 1247
rect 750 1236 756 1237
rect 830 1236 836 1237
rect 750 1232 751 1236
rect 755 1232 756 1236
rect 750 1231 756 1232
rect 762 1235 768 1236
rect 762 1231 763 1235
rect 767 1231 768 1235
rect 830 1232 831 1236
rect 835 1232 836 1236
rect 830 1231 836 1232
rect 910 1236 916 1237
rect 910 1232 911 1236
rect 915 1232 916 1236
rect 910 1231 916 1232
rect 990 1236 996 1237
rect 990 1232 991 1236
rect 995 1232 996 1236
rect 990 1231 996 1232
rect 1062 1236 1068 1237
rect 1062 1232 1063 1236
rect 1067 1232 1068 1236
rect 1062 1231 1068 1232
rect 1126 1236 1132 1237
rect 1126 1232 1127 1236
rect 1131 1232 1132 1236
rect 1126 1231 1132 1232
rect 1190 1236 1196 1237
rect 1190 1232 1191 1236
rect 1195 1232 1196 1236
rect 1190 1231 1196 1232
rect 1246 1236 1252 1237
rect 1246 1232 1247 1236
rect 1251 1232 1252 1236
rect 1246 1231 1252 1232
rect 703 1230 707 1231
rect 703 1225 707 1226
rect 751 1230 755 1231
rect 762 1230 768 1231
rect 799 1230 803 1231
rect 751 1225 755 1226
rect 702 1224 708 1225
rect 702 1220 703 1224
rect 707 1220 708 1224
rect 702 1219 708 1220
rect 750 1224 756 1225
rect 750 1220 751 1224
rect 755 1220 756 1224
rect 750 1219 756 1220
rect 458 1215 464 1216
rect 458 1211 459 1215
rect 463 1211 464 1215
rect 458 1210 464 1211
rect 690 1215 696 1216
rect 690 1211 691 1215
rect 695 1211 696 1215
rect 690 1210 696 1211
rect 346 1207 352 1208
rect 110 1203 116 1204
rect 110 1199 111 1203
rect 115 1199 116 1203
rect 346 1203 347 1207
rect 351 1203 352 1207
rect 346 1202 352 1203
rect 110 1198 116 1199
rect 326 1198 332 1199
rect 112 1191 114 1198
rect 326 1194 327 1198
rect 331 1194 332 1198
rect 326 1193 332 1194
rect 170 1191 176 1192
rect 328 1191 330 1193
rect 111 1190 115 1191
rect 111 1185 115 1186
rect 135 1190 139 1191
rect 135 1185 139 1186
rect 159 1190 163 1191
rect 170 1187 171 1191
rect 175 1187 176 1191
rect 170 1186 176 1187
rect 183 1190 187 1191
rect 159 1185 163 1186
rect 112 1178 114 1185
rect 136 1183 138 1185
rect 160 1183 162 1185
rect 134 1182 140 1183
rect 134 1178 135 1182
rect 139 1178 140 1182
rect 110 1177 116 1178
rect 134 1177 140 1178
rect 158 1182 164 1183
rect 158 1178 159 1182
rect 163 1178 164 1182
rect 158 1177 164 1178
rect 110 1173 111 1177
rect 115 1173 116 1177
rect 110 1172 116 1173
rect 110 1159 116 1160
rect 110 1155 111 1159
rect 115 1155 116 1159
rect 110 1154 116 1155
rect 134 1156 140 1157
rect 158 1156 164 1157
rect 172 1156 174 1186
rect 183 1185 187 1186
rect 207 1190 211 1191
rect 207 1185 211 1186
rect 231 1190 235 1191
rect 231 1185 235 1186
rect 255 1190 259 1191
rect 255 1185 259 1186
rect 279 1190 283 1191
rect 279 1185 283 1186
rect 303 1190 307 1191
rect 303 1185 307 1186
rect 327 1190 331 1191
rect 327 1185 331 1186
rect 335 1190 339 1191
rect 335 1185 339 1186
rect 184 1183 186 1185
rect 208 1183 210 1185
rect 232 1183 234 1185
rect 256 1183 258 1185
rect 280 1183 282 1185
rect 304 1183 306 1185
rect 336 1183 338 1185
rect 348 1184 350 1202
rect 460 1200 462 1210
rect 764 1200 766 1230
rect 799 1225 803 1226
rect 831 1230 835 1231
rect 831 1225 835 1226
rect 847 1230 851 1231
rect 847 1225 851 1226
rect 895 1230 899 1231
rect 895 1225 899 1226
rect 911 1230 915 1231
rect 911 1225 915 1226
rect 943 1230 947 1231
rect 943 1225 947 1226
rect 991 1230 995 1231
rect 991 1225 995 1226
rect 1039 1230 1043 1231
rect 1039 1225 1043 1226
rect 1063 1230 1067 1231
rect 1063 1225 1067 1226
rect 1103 1230 1107 1231
rect 1103 1225 1107 1226
rect 1127 1230 1131 1231
rect 1127 1225 1131 1226
rect 1175 1230 1179 1231
rect 1175 1225 1179 1226
rect 1191 1230 1195 1231
rect 1191 1225 1195 1226
rect 1247 1230 1251 1231
rect 1247 1225 1251 1226
rect 1255 1230 1259 1231
rect 1255 1225 1259 1226
rect 798 1224 804 1225
rect 798 1220 799 1224
rect 803 1220 804 1224
rect 798 1219 804 1220
rect 846 1224 852 1225
rect 846 1220 847 1224
rect 851 1220 852 1224
rect 846 1219 852 1220
rect 894 1224 900 1225
rect 894 1220 895 1224
rect 899 1220 900 1224
rect 894 1219 900 1220
rect 942 1224 948 1225
rect 942 1220 943 1224
rect 947 1220 948 1224
rect 942 1219 948 1220
rect 990 1224 996 1225
rect 990 1220 991 1224
rect 995 1220 996 1224
rect 990 1219 996 1220
rect 1038 1224 1044 1225
rect 1038 1220 1039 1224
rect 1043 1220 1044 1224
rect 1038 1219 1044 1220
rect 1102 1224 1108 1225
rect 1102 1220 1103 1224
rect 1107 1220 1108 1224
rect 1102 1219 1108 1220
rect 1174 1224 1180 1225
rect 1174 1220 1175 1224
rect 1179 1220 1180 1224
rect 1174 1219 1180 1220
rect 1254 1224 1260 1225
rect 1254 1220 1255 1224
rect 1259 1220 1260 1224
rect 1254 1219 1260 1220
rect 1296 1216 1298 1266
rect 1303 1265 1307 1266
rect 1311 1270 1315 1271
rect 1322 1267 1323 1271
rect 1327 1267 1328 1271
rect 1322 1266 1328 1267
rect 1367 1270 1371 1271
rect 1311 1265 1315 1266
rect 1312 1263 1314 1265
rect 1310 1262 1316 1263
rect 1310 1258 1311 1262
rect 1315 1258 1316 1262
rect 1310 1257 1316 1258
rect 1324 1252 1326 1266
rect 1367 1265 1371 1266
rect 1375 1270 1379 1271
rect 1375 1265 1379 1266
rect 1376 1263 1378 1265
rect 1388 1264 1390 1282
rect 1428 1280 1430 1310
rect 1447 1305 1451 1306
rect 1448 1302 1450 1305
rect 1446 1301 1452 1302
rect 1446 1297 1447 1301
rect 1451 1297 1452 1301
rect 1446 1296 1452 1297
rect 1446 1283 1452 1284
rect 1426 1279 1432 1280
rect 1414 1278 1420 1279
rect 1414 1274 1415 1278
rect 1419 1274 1420 1278
rect 1426 1275 1427 1279
rect 1431 1275 1432 1279
rect 1446 1279 1447 1283
rect 1451 1279 1452 1283
rect 1446 1278 1452 1279
rect 1426 1274 1432 1275
rect 1414 1273 1420 1274
rect 1416 1271 1418 1273
rect 1448 1271 1450 1278
rect 1415 1270 1419 1271
rect 1415 1265 1419 1266
rect 1447 1270 1451 1271
rect 1447 1265 1451 1266
rect 1386 1263 1392 1264
rect 1416 1263 1418 1265
rect 1374 1262 1380 1263
rect 1374 1258 1375 1262
rect 1379 1258 1380 1262
rect 1386 1259 1387 1263
rect 1391 1259 1392 1263
rect 1386 1258 1392 1259
rect 1414 1262 1420 1263
rect 1414 1258 1415 1262
rect 1419 1258 1420 1262
rect 1448 1258 1450 1265
rect 1374 1257 1380 1258
rect 1414 1257 1420 1258
rect 1446 1257 1452 1258
rect 1446 1253 1447 1257
rect 1451 1253 1452 1257
rect 1446 1252 1452 1253
rect 1322 1251 1328 1252
rect 1322 1247 1323 1251
rect 1327 1247 1328 1251
rect 1322 1246 1328 1247
rect 1446 1239 1452 1240
rect 1310 1236 1316 1237
rect 1310 1232 1311 1236
rect 1315 1232 1316 1236
rect 1310 1231 1316 1232
rect 1374 1236 1380 1237
rect 1374 1232 1375 1236
rect 1379 1232 1380 1236
rect 1374 1231 1380 1232
rect 1414 1236 1420 1237
rect 1414 1232 1415 1236
rect 1419 1232 1420 1236
rect 1414 1231 1420 1232
rect 1426 1235 1432 1236
rect 1426 1231 1427 1235
rect 1431 1231 1432 1235
rect 1446 1235 1447 1239
rect 1451 1235 1452 1239
rect 1446 1234 1452 1235
rect 1448 1231 1450 1234
rect 1311 1230 1315 1231
rect 1311 1225 1315 1226
rect 1343 1230 1347 1231
rect 1343 1225 1347 1226
rect 1375 1230 1379 1231
rect 1375 1225 1379 1226
rect 1415 1230 1419 1231
rect 1426 1230 1432 1231
rect 1447 1230 1451 1231
rect 1415 1225 1419 1226
rect 1342 1224 1348 1225
rect 1342 1220 1343 1224
rect 1347 1220 1348 1224
rect 1342 1219 1348 1220
rect 1414 1224 1420 1225
rect 1414 1220 1415 1224
rect 1419 1220 1420 1224
rect 1414 1219 1420 1220
rect 810 1215 816 1216
rect 810 1211 811 1215
rect 815 1211 816 1215
rect 810 1210 816 1211
rect 906 1215 912 1216
rect 906 1211 907 1215
rect 911 1211 912 1215
rect 906 1210 912 1211
rect 1002 1215 1008 1216
rect 1002 1211 1003 1215
rect 1007 1211 1008 1215
rect 1002 1210 1008 1211
rect 1114 1215 1120 1216
rect 1114 1211 1115 1215
rect 1119 1211 1120 1215
rect 1114 1210 1120 1211
rect 1266 1215 1272 1216
rect 1266 1211 1267 1215
rect 1271 1211 1272 1215
rect 1266 1210 1272 1211
rect 1294 1215 1300 1216
rect 1294 1211 1295 1215
rect 1299 1211 1300 1215
rect 1294 1210 1300 1211
rect 812 1200 814 1210
rect 908 1200 910 1210
rect 922 1207 928 1208
rect 922 1203 923 1207
rect 927 1203 928 1207
rect 922 1202 928 1203
rect 458 1199 464 1200
rect 762 1199 768 1200
rect 810 1199 816 1200
rect 906 1199 912 1200
rect 366 1198 372 1199
rect 366 1194 367 1198
rect 371 1194 372 1198
rect 366 1193 372 1194
rect 406 1198 412 1199
rect 406 1194 407 1198
rect 411 1194 412 1198
rect 406 1193 412 1194
rect 446 1198 452 1199
rect 446 1194 447 1198
rect 451 1194 452 1198
rect 458 1195 459 1199
rect 463 1195 464 1199
rect 458 1194 464 1195
rect 486 1198 492 1199
rect 486 1194 487 1198
rect 491 1194 492 1198
rect 446 1193 452 1194
rect 486 1193 492 1194
rect 526 1198 532 1199
rect 526 1194 527 1198
rect 531 1194 532 1198
rect 526 1193 532 1194
rect 566 1198 572 1199
rect 566 1194 567 1198
rect 571 1194 572 1198
rect 566 1193 572 1194
rect 606 1198 612 1199
rect 606 1194 607 1198
rect 611 1194 612 1198
rect 606 1193 612 1194
rect 654 1198 660 1199
rect 654 1194 655 1198
rect 659 1194 660 1198
rect 654 1193 660 1194
rect 702 1198 708 1199
rect 702 1194 703 1198
rect 707 1194 708 1198
rect 702 1193 708 1194
rect 750 1198 756 1199
rect 750 1194 751 1198
rect 755 1194 756 1198
rect 762 1195 763 1199
rect 767 1195 768 1199
rect 762 1194 768 1195
rect 798 1198 804 1199
rect 798 1194 799 1198
rect 803 1194 804 1198
rect 810 1195 811 1199
rect 815 1195 816 1199
rect 810 1194 816 1195
rect 846 1198 852 1199
rect 846 1194 847 1198
rect 851 1194 852 1198
rect 750 1193 756 1194
rect 798 1193 804 1194
rect 846 1193 852 1194
rect 894 1198 900 1199
rect 894 1194 895 1198
rect 899 1194 900 1198
rect 906 1195 907 1199
rect 911 1195 912 1199
rect 906 1194 912 1195
rect 894 1193 900 1194
rect 368 1191 370 1193
rect 408 1191 410 1193
rect 414 1191 420 1192
rect 448 1191 450 1193
rect 488 1191 490 1193
rect 528 1191 530 1193
rect 568 1191 570 1193
rect 608 1191 610 1193
rect 656 1191 658 1193
rect 694 1191 700 1192
rect 704 1191 706 1193
rect 752 1191 754 1193
rect 778 1191 784 1192
rect 800 1191 802 1193
rect 848 1191 850 1193
rect 896 1191 898 1193
rect 367 1190 371 1191
rect 367 1185 371 1186
rect 383 1190 387 1191
rect 383 1185 387 1186
rect 407 1190 411 1191
rect 414 1187 415 1191
rect 419 1187 420 1191
rect 414 1186 420 1187
rect 423 1190 427 1191
rect 407 1185 411 1186
rect 346 1183 352 1184
rect 384 1183 386 1185
rect 182 1182 188 1183
rect 182 1178 183 1182
rect 187 1178 188 1182
rect 182 1177 188 1178
rect 206 1182 212 1183
rect 206 1178 207 1182
rect 211 1178 212 1182
rect 206 1177 212 1178
rect 230 1182 236 1183
rect 230 1178 231 1182
rect 235 1178 236 1182
rect 230 1177 236 1178
rect 254 1182 260 1183
rect 254 1178 255 1182
rect 259 1178 260 1182
rect 254 1177 260 1178
rect 278 1182 284 1183
rect 278 1178 279 1182
rect 283 1178 284 1182
rect 278 1177 284 1178
rect 302 1182 308 1183
rect 302 1178 303 1182
rect 307 1178 308 1182
rect 334 1182 340 1183
rect 302 1177 308 1178
rect 314 1179 320 1180
rect 314 1175 315 1179
rect 319 1175 320 1179
rect 334 1178 335 1182
rect 339 1178 340 1182
rect 346 1179 347 1183
rect 351 1179 352 1183
rect 346 1178 352 1179
rect 382 1182 388 1183
rect 382 1178 383 1182
rect 387 1178 388 1182
rect 334 1177 340 1178
rect 382 1177 388 1178
rect 314 1174 320 1175
rect 182 1156 188 1157
rect 112 1151 114 1154
rect 134 1152 135 1156
rect 139 1152 140 1156
rect 134 1151 140 1152
rect 146 1155 152 1156
rect 146 1151 147 1155
rect 151 1151 152 1155
rect 158 1152 159 1156
rect 163 1152 164 1156
rect 158 1151 164 1152
rect 170 1155 176 1156
rect 170 1151 171 1155
rect 175 1151 176 1155
rect 182 1152 183 1156
rect 187 1152 188 1156
rect 182 1151 188 1152
rect 206 1156 212 1157
rect 206 1152 207 1156
rect 211 1152 212 1156
rect 206 1151 212 1152
rect 230 1156 236 1157
rect 230 1152 231 1156
rect 235 1152 236 1156
rect 230 1151 236 1152
rect 254 1156 260 1157
rect 254 1152 255 1156
rect 259 1152 260 1156
rect 254 1151 260 1152
rect 278 1156 284 1157
rect 278 1152 279 1156
rect 283 1152 284 1156
rect 278 1151 284 1152
rect 302 1156 308 1157
rect 302 1152 303 1156
rect 307 1152 308 1156
rect 302 1151 308 1152
rect 111 1150 115 1151
rect 111 1145 115 1146
rect 135 1150 139 1151
rect 146 1150 152 1151
rect 159 1150 163 1151
rect 170 1150 176 1151
rect 183 1150 187 1151
rect 135 1145 139 1146
rect 112 1142 114 1145
rect 134 1144 140 1145
rect 110 1141 116 1142
rect 110 1137 111 1141
rect 115 1137 116 1141
rect 134 1140 135 1144
rect 139 1140 140 1144
rect 134 1139 140 1140
rect 110 1136 116 1137
rect 110 1123 116 1124
rect 110 1119 111 1123
rect 115 1119 116 1123
rect 148 1120 150 1150
rect 159 1145 163 1146
rect 183 1145 187 1146
rect 207 1150 211 1151
rect 207 1145 211 1146
rect 215 1150 219 1151
rect 215 1145 219 1146
rect 231 1150 235 1151
rect 231 1145 235 1146
rect 255 1150 259 1151
rect 255 1145 259 1146
rect 279 1150 283 1151
rect 279 1145 283 1146
rect 295 1150 299 1151
rect 295 1145 299 1146
rect 303 1150 307 1151
rect 303 1145 307 1146
rect 158 1144 164 1145
rect 158 1140 159 1144
rect 163 1140 164 1144
rect 158 1139 164 1140
rect 182 1144 188 1145
rect 182 1140 183 1144
rect 187 1140 188 1144
rect 182 1139 188 1140
rect 214 1144 220 1145
rect 214 1140 215 1144
rect 219 1140 220 1144
rect 214 1139 220 1140
rect 254 1144 260 1145
rect 254 1140 255 1144
rect 259 1140 260 1144
rect 254 1139 260 1140
rect 294 1144 300 1145
rect 294 1140 295 1144
rect 299 1140 300 1144
rect 294 1139 300 1140
rect 316 1136 318 1174
rect 398 1167 404 1168
rect 398 1163 399 1167
rect 403 1163 404 1167
rect 398 1162 404 1163
rect 334 1156 340 1157
rect 334 1152 335 1156
rect 339 1152 340 1156
rect 334 1151 340 1152
rect 382 1156 388 1157
rect 382 1152 383 1156
rect 387 1152 388 1156
rect 382 1151 388 1152
rect 335 1150 339 1151
rect 335 1145 339 1146
rect 375 1150 379 1151
rect 375 1145 379 1146
rect 383 1150 387 1151
rect 383 1145 387 1146
rect 334 1144 340 1145
rect 334 1140 335 1144
rect 339 1140 340 1144
rect 334 1139 340 1140
rect 374 1144 380 1145
rect 374 1140 375 1144
rect 379 1140 380 1144
rect 374 1139 380 1140
rect 170 1135 176 1136
rect 170 1131 171 1135
rect 175 1131 176 1135
rect 170 1130 176 1131
rect 314 1135 320 1136
rect 314 1131 315 1135
rect 319 1131 320 1135
rect 314 1130 320 1131
rect 172 1120 174 1130
rect 400 1128 402 1162
rect 416 1160 418 1186
rect 423 1185 427 1186
rect 447 1190 451 1191
rect 447 1185 451 1186
rect 463 1190 467 1191
rect 463 1185 467 1186
rect 487 1190 491 1191
rect 487 1185 491 1186
rect 503 1190 507 1191
rect 503 1185 507 1186
rect 527 1190 531 1191
rect 527 1185 531 1186
rect 543 1190 547 1191
rect 543 1185 547 1186
rect 567 1190 571 1191
rect 567 1185 571 1186
rect 583 1190 587 1191
rect 583 1185 587 1186
rect 607 1190 611 1191
rect 607 1185 611 1186
rect 623 1190 627 1191
rect 623 1185 627 1186
rect 655 1190 659 1191
rect 655 1185 659 1186
rect 671 1190 675 1191
rect 694 1187 695 1191
rect 699 1187 700 1191
rect 694 1186 700 1187
rect 703 1190 707 1191
rect 671 1185 675 1186
rect 424 1183 426 1185
rect 464 1183 466 1185
rect 504 1183 506 1185
rect 544 1183 546 1185
rect 584 1183 586 1185
rect 624 1183 626 1185
rect 672 1183 674 1185
rect 422 1182 428 1183
rect 422 1178 423 1182
rect 427 1178 428 1182
rect 422 1177 428 1178
rect 462 1182 468 1183
rect 462 1178 463 1182
rect 467 1178 468 1182
rect 462 1177 468 1178
rect 502 1182 508 1183
rect 502 1178 503 1182
rect 507 1178 508 1182
rect 502 1177 508 1178
rect 542 1182 548 1183
rect 542 1178 543 1182
rect 547 1178 548 1182
rect 542 1177 548 1178
rect 582 1182 588 1183
rect 582 1178 583 1182
rect 587 1178 588 1182
rect 582 1177 588 1178
rect 622 1182 628 1183
rect 622 1178 623 1182
rect 627 1178 628 1182
rect 622 1177 628 1178
rect 670 1182 676 1183
rect 670 1178 671 1182
rect 675 1178 676 1182
rect 670 1177 676 1178
rect 414 1159 420 1160
rect 414 1155 415 1159
rect 419 1155 420 1159
rect 414 1154 420 1155
rect 422 1156 428 1157
rect 422 1152 423 1156
rect 427 1152 428 1156
rect 422 1151 428 1152
rect 462 1156 468 1157
rect 462 1152 463 1156
rect 467 1152 468 1156
rect 462 1151 468 1152
rect 502 1156 508 1157
rect 502 1152 503 1156
rect 507 1152 508 1156
rect 502 1151 508 1152
rect 542 1156 548 1157
rect 542 1152 543 1156
rect 547 1152 548 1156
rect 542 1151 548 1152
rect 582 1156 588 1157
rect 582 1152 583 1156
rect 587 1152 588 1156
rect 582 1151 588 1152
rect 622 1156 628 1157
rect 622 1152 623 1156
rect 627 1152 628 1156
rect 622 1151 628 1152
rect 670 1156 676 1157
rect 670 1152 671 1156
rect 675 1152 676 1156
rect 670 1151 676 1152
rect 415 1150 419 1151
rect 415 1145 419 1146
rect 423 1150 427 1151
rect 423 1145 427 1146
rect 463 1150 467 1151
rect 463 1145 467 1146
rect 503 1150 507 1151
rect 503 1145 507 1146
rect 519 1150 523 1151
rect 519 1145 523 1146
rect 543 1150 547 1151
rect 543 1145 547 1146
rect 583 1150 587 1151
rect 583 1145 587 1146
rect 623 1150 627 1151
rect 623 1145 627 1146
rect 647 1150 651 1151
rect 647 1145 651 1146
rect 671 1150 675 1151
rect 671 1145 675 1146
rect 414 1144 420 1145
rect 414 1140 415 1144
rect 419 1140 420 1144
rect 414 1139 420 1140
rect 462 1144 468 1145
rect 462 1140 463 1144
rect 467 1140 468 1144
rect 462 1139 468 1140
rect 518 1144 524 1145
rect 518 1140 519 1144
rect 523 1140 524 1144
rect 518 1139 524 1140
rect 582 1144 588 1145
rect 582 1140 583 1144
rect 587 1140 588 1144
rect 582 1139 588 1140
rect 646 1144 652 1145
rect 646 1140 647 1144
rect 651 1140 652 1144
rect 646 1139 652 1140
rect 696 1136 698 1186
rect 703 1185 707 1186
rect 719 1190 723 1191
rect 719 1185 723 1186
rect 751 1190 755 1191
rect 751 1185 755 1186
rect 767 1190 771 1191
rect 778 1187 779 1191
rect 783 1187 784 1191
rect 778 1186 784 1187
rect 799 1190 803 1191
rect 767 1185 771 1186
rect 720 1183 722 1185
rect 768 1183 770 1185
rect 718 1182 724 1183
rect 718 1178 719 1182
rect 723 1178 724 1182
rect 718 1177 724 1178
rect 766 1182 772 1183
rect 766 1178 767 1182
rect 771 1178 772 1182
rect 766 1177 772 1178
rect 780 1160 782 1186
rect 799 1185 803 1186
rect 815 1190 819 1191
rect 815 1185 819 1186
rect 847 1190 851 1191
rect 847 1185 851 1186
rect 863 1190 867 1191
rect 863 1185 867 1186
rect 895 1190 899 1191
rect 895 1185 899 1186
rect 911 1190 915 1191
rect 911 1185 915 1186
rect 816 1183 818 1185
rect 864 1183 866 1185
rect 912 1183 914 1185
rect 924 1184 926 1202
rect 1004 1200 1006 1210
rect 1116 1200 1118 1210
rect 1268 1200 1270 1210
rect 1428 1200 1430 1230
rect 1447 1225 1451 1226
rect 1448 1222 1450 1225
rect 1446 1221 1452 1222
rect 1446 1217 1447 1221
rect 1451 1217 1452 1221
rect 1446 1216 1452 1217
rect 1446 1203 1452 1204
rect 1002 1199 1008 1200
rect 1114 1199 1120 1200
rect 1266 1199 1272 1200
rect 1426 1199 1432 1200
rect 942 1198 948 1199
rect 942 1194 943 1198
rect 947 1194 948 1198
rect 942 1193 948 1194
rect 990 1198 996 1199
rect 990 1194 991 1198
rect 995 1194 996 1198
rect 1002 1195 1003 1199
rect 1007 1195 1008 1199
rect 1002 1194 1008 1195
rect 1038 1198 1044 1199
rect 1038 1194 1039 1198
rect 1043 1194 1044 1198
rect 990 1193 996 1194
rect 1038 1193 1044 1194
rect 1102 1198 1108 1199
rect 1102 1194 1103 1198
rect 1107 1194 1108 1198
rect 1114 1195 1115 1199
rect 1119 1195 1120 1199
rect 1114 1194 1120 1195
rect 1174 1198 1180 1199
rect 1174 1194 1175 1198
rect 1179 1194 1180 1198
rect 1102 1193 1108 1194
rect 1174 1193 1180 1194
rect 1254 1198 1260 1199
rect 1254 1194 1255 1198
rect 1259 1194 1260 1198
rect 1266 1195 1267 1199
rect 1271 1195 1272 1199
rect 1266 1194 1272 1195
rect 1342 1198 1348 1199
rect 1342 1194 1343 1198
rect 1347 1194 1348 1198
rect 1254 1193 1260 1194
rect 1342 1193 1348 1194
rect 1414 1198 1420 1199
rect 1414 1194 1415 1198
rect 1419 1194 1420 1198
rect 1426 1195 1427 1199
rect 1431 1195 1432 1199
rect 1446 1199 1447 1203
rect 1451 1199 1452 1203
rect 1446 1198 1452 1199
rect 1426 1194 1432 1195
rect 1414 1193 1420 1194
rect 944 1191 946 1193
rect 992 1191 994 1193
rect 1040 1191 1042 1193
rect 1104 1191 1106 1193
rect 1114 1191 1120 1192
rect 1176 1191 1178 1193
rect 1256 1191 1258 1193
rect 1282 1191 1288 1192
rect 1344 1191 1346 1193
rect 1416 1191 1418 1193
rect 1448 1191 1450 1198
rect 943 1190 947 1191
rect 943 1185 947 1186
rect 959 1190 963 1191
rect 959 1185 963 1186
rect 991 1190 995 1191
rect 991 1185 995 1186
rect 1007 1190 1011 1191
rect 1007 1185 1011 1186
rect 1039 1190 1043 1191
rect 1039 1185 1043 1186
rect 1055 1190 1059 1191
rect 1055 1185 1059 1186
rect 1103 1190 1107 1191
rect 1114 1187 1115 1191
rect 1119 1187 1120 1191
rect 1114 1186 1120 1187
rect 1151 1190 1155 1191
rect 1103 1185 1107 1186
rect 922 1183 928 1184
rect 960 1183 962 1185
rect 1008 1183 1010 1185
rect 1056 1183 1058 1185
rect 1104 1183 1106 1185
rect 814 1182 820 1183
rect 814 1178 815 1182
rect 819 1178 820 1182
rect 814 1177 820 1178
rect 862 1182 868 1183
rect 862 1178 863 1182
rect 867 1178 868 1182
rect 862 1177 868 1178
rect 910 1182 916 1183
rect 910 1178 911 1182
rect 915 1178 916 1182
rect 922 1179 923 1183
rect 927 1179 928 1183
rect 922 1178 928 1179
rect 958 1182 964 1183
rect 958 1178 959 1182
rect 963 1178 964 1182
rect 1006 1182 1012 1183
rect 910 1177 916 1178
rect 958 1177 964 1178
rect 998 1179 1004 1180
rect 998 1175 999 1179
rect 1003 1175 1004 1179
rect 1006 1178 1007 1182
rect 1011 1178 1012 1182
rect 1006 1177 1012 1178
rect 1054 1182 1060 1183
rect 1054 1178 1055 1182
rect 1059 1178 1060 1182
rect 1054 1177 1060 1178
rect 1102 1182 1108 1183
rect 1102 1178 1103 1182
rect 1107 1178 1108 1182
rect 1102 1177 1108 1178
rect 998 1174 1004 1175
rect 1000 1163 1002 1174
rect 1000 1161 1022 1163
rect 778 1159 784 1160
rect 718 1156 724 1157
rect 718 1152 719 1156
rect 723 1152 724 1156
rect 718 1151 724 1152
rect 766 1156 772 1157
rect 766 1152 767 1156
rect 771 1152 772 1156
rect 778 1155 779 1159
rect 783 1155 784 1159
rect 778 1154 784 1155
rect 814 1156 820 1157
rect 766 1151 772 1152
rect 814 1152 815 1156
rect 819 1152 820 1156
rect 862 1156 868 1157
rect 862 1152 863 1156
rect 867 1152 868 1156
rect 814 1151 820 1152
rect 822 1151 828 1152
rect 862 1151 868 1152
rect 910 1156 916 1157
rect 910 1152 911 1156
rect 915 1152 916 1156
rect 910 1151 916 1152
rect 958 1156 964 1157
rect 958 1152 959 1156
rect 963 1152 964 1156
rect 958 1151 964 1152
rect 1006 1156 1012 1157
rect 1006 1152 1007 1156
rect 1011 1152 1012 1156
rect 1006 1151 1012 1152
rect 711 1150 715 1151
rect 711 1145 715 1146
rect 719 1150 723 1151
rect 719 1145 723 1146
rect 767 1150 771 1151
rect 767 1145 771 1146
rect 815 1150 819 1151
rect 822 1147 823 1151
rect 827 1147 828 1151
rect 822 1146 828 1147
rect 831 1150 835 1151
rect 815 1145 819 1146
rect 710 1144 716 1145
rect 710 1140 711 1144
rect 715 1140 716 1144
rect 710 1139 716 1140
rect 766 1144 772 1145
rect 766 1140 767 1144
rect 771 1140 772 1144
rect 766 1139 772 1140
rect 426 1135 432 1136
rect 426 1131 427 1135
rect 431 1131 432 1135
rect 426 1130 432 1131
rect 530 1135 536 1136
rect 530 1131 531 1135
rect 535 1131 536 1135
rect 530 1130 536 1131
rect 658 1135 664 1136
rect 658 1131 659 1135
rect 663 1131 664 1135
rect 658 1130 664 1131
rect 694 1135 700 1136
rect 694 1131 695 1135
rect 699 1131 700 1135
rect 694 1130 700 1131
rect 194 1127 200 1128
rect 194 1123 195 1127
rect 199 1123 200 1127
rect 194 1122 200 1123
rect 398 1127 404 1128
rect 398 1123 399 1127
rect 403 1123 404 1127
rect 398 1122 404 1123
rect 146 1119 152 1120
rect 170 1119 176 1120
rect 110 1118 116 1119
rect 134 1118 140 1119
rect 112 1107 114 1118
rect 134 1114 135 1118
rect 139 1114 140 1118
rect 146 1115 147 1119
rect 151 1115 152 1119
rect 146 1114 152 1115
rect 158 1118 164 1119
rect 158 1114 159 1118
rect 163 1114 164 1118
rect 170 1115 171 1119
rect 175 1115 176 1119
rect 170 1114 176 1115
rect 182 1118 188 1119
rect 182 1114 183 1118
rect 187 1114 188 1118
rect 134 1113 140 1114
rect 158 1113 164 1114
rect 182 1113 188 1114
rect 136 1107 138 1113
rect 160 1107 162 1113
rect 184 1107 186 1113
rect 111 1106 115 1107
rect 111 1101 115 1102
rect 135 1106 139 1107
rect 135 1101 139 1102
rect 159 1106 163 1107
rect 159 1101 163 1102
rect 183 1106 187 1107
rect 183 1101 187 1102
rect 112 1094 114 1101
rect 136 1099 138 1101
rect 160 1099 162 1101
rect 184 1099 186 1101
rect 196 1100 198 1122
rect 428 1120 430 1130
rect 532 1120 534 1130
rect 660 1120 662 1130
rect 824 1120 826 1146
rect 831 1145 835 1146
rect 863 1150 867 1151
rect 863 1145 867 1146
rect 887 1150 891 1151
rect 887 1145 891 1146
rect 911 1150 915 1151
rect 911 1145 915 1146
rect 943 1150 947 1151
rect 943 1145 947 1146
rect 959 1150 963 1151
rect 959 1145 963 1146
rect 999 1150 1003 1151
rect 999 1145 1003 1146
rect 1007 1150 1011 1151
rect 1007 1145 1011 1146
rect 830 1144 836 1145
rect 830 1140 831 1144
rect 835 1140 836 1144
rect 830 1139 836 1140
rect 886 1144 892 1145
rect 886 1140 887 1144
rect 891 1140 892 1144
rect 886 1139 892 1140
rect 942 1144 948 1145
rect 942 1140 943 1144
rect 947 1140 948 1144
rect 942 1139 948 1140
rect 998 1144 1004 1145
rect 998 1140 999 1144
rect 1003 1140 1004 1144
rect 998 1139 1004 1140
rect 1020 1136 1022 1161
rect 1116 1160 1118 1186
rect 1151 1185 1155 1186
rect 1175 1190 1179 1191
rect 1175 1185 1179 1186
rect 1191 1190 1195 1191
rect 1191 1185 1195 1186
rect 1231 1190 1235 1191
rect 1231 1185 1235 1186
rect 1255 1190 1259 1191
rect 1255 1185 1259 1186
rect 1271 1190 1275 1191
rect 1282 1187 1283 1191
rect 1287 1187 1288 1191
rect 1282 1186 1288 1187
rect 1311 1190 1315 1191
rect 1271 1185 1275 1186
rect 1152 1183 1154 1185
rect 1192 1183 1194 1185
rect 1232 1183 1234 1185
rect 1272 1183 1274 1185
rect 1150 1182 1156 1183
rect 1150 1178 1151 1182
rect 1155 1178 1156 1182
rect 1190 1182 1196 1183
rect 1150 1177 1156 1178
rect 1182 1179 1188 1180
rect 1182 1175 1183 1179
rect 1187 1175 1188 1179
rect 1190 1178 1191 1182
rect 1195 1178 1196 1182
rect 1190 1177 1196 1178
rect 1230 1182 1236 1183
rect 1230 1178 1231 1182
rect 1235 1178 1236 1182
rect 1230 1177 1236 1178
rect 1270 1182 1276 1183
rect 1270 1178 1271 1182
rect 1275 1178 1276 1182
rect 1270 1177 1276 1178
rect 1182 1174 1188 1175
rect 1184 1171 1186 1174
rect 1184 1169 1206 1171
rect 1204 1160 1206 1169
rect 1114 1159 1120 1160
rect 1054 1156 1060 1157
rect 1054 1152 1055 1156
rect 1059 1152 1060 1156
rect 1054 1151 1060 1152
rect 1102 1156 1108 1157
rect 1102 1152 1103 1156
rect 1107 1152 1108 1156
rect 1114 1155 1115 1159
rect 1119 1155 1120 1159
rect 1202 1159 1208 1160
rect 1114 1154 1120 1155
rect 1150 1156 1156 1157
rect 1190 1156 1196 1157
rect 1102 1151 1108 1152
rect 1150 1152 1151 1156
rect 1155 1152 1156 1156
rect 1150 1151 1156 1152
rect 1182 1155 1188 1156
rect 1182 1151 1183 1155
rect 1187 1151 1188 1155
rect 1190 1152 1191 1156
rect 1195 1152 1196 1156
rect 1202 1155 1203 1159
rect 1207 1155 1208 1159
rect 1202 1154 1208 1155
rect 1230 1156 1236 1157
rect 1190 1151 1196 1152
rect 1230 1152 1231 1156
rect 1235 1152 1236 1156
rect 1230 1151 1236 1152
rect 1270 1156 1276 1157
rect 1284 1156 1286 1186
rect 1311 1185 1315 1186
rect 1343 1190 1347 1191
rect 1343 1185 1347 1186
rect 1351 1190 1355 1191
rect 1351 1185 1355 1186
rect 1391 1190 1395 1191
rect 1391 1185 1395 1186
rect 1415 1190 1419 1191
rect 1415 1185 1419 1186
rect 1447 1190 1451 1191
rect 1447 1185 1451 1186
rect 1312 1183 1314 1185
rect 1352 1183 1354 1185
rect 1392 1183 1394 1185
rect 1416 1183 1418 1185
rect 1310 1182 1316 1183
rect 1310 1178 1311 1182
rect 1315 1178 1316 1182
rect 1310 1177 1316 1178
rect 1350 1182 1356 1183
rect 1350 1178 1351 1182
rect 1355 1178 1356 1182
rect 1390 1182 1396 1183
rect 1350 1177 1356 1178
rect 1362 1179 1368 1180
rect 1362 1175 1363 1179
rect 1367 1175 1368 1179
rect 1390 1178 1391 1182
rect 1395 1178 1396 1182
rect 1390 1177 1396 1178
rect 1414 1182 1420 1183
rect 1414 1178 1415 1182
rect 1419 1178 1420 1182
rect 1448 1178 1450 1185
rect 1414 1177 1420 1178
rect 1446 1177 1452 1178
rect 1362 1174 1368 1175
rect 1310 1156 1316 1157
rect 1270 1152 1271 1156
rect 1275 1152 1276 1156
rect 1270 1151 1276 1152
rect 1282 1155 1288 1156
rect 1282 1151 1283 1155
rect 1287 1151 1288 1155
rect 1310 1152 1311 1156
rect 1315 1152 1316 1156
rect 1310 1151 1316 1152
rect 1350 1156 1356 1157
rect 1350 1152 1351 1156
rect 1355 1152 1356 1156
rect 1350 1151 1356 1152
rect 1055 1150 1059 1151
rect 1055 1145 1059 1146
rect 1103 1150 1107 1151
rect 1103 1145 1107 1146
rect 1151 1150 1155 1151
rect 1182 1150 1188 1151
rect 1191 1150 1195 1151
rect 1151 1145 1155 1146
rect 1054 1144 1060 1145
rect 1054 1140 1055 1144
rect 1059 1140 1060 1144
rect 1054 1139 1060 1140
rect 1102 1144 1108 1145
rect 1102 1140 1103 1144
rect 1107 1140 1108 1144
rect 1102 1139 1108 1140
rect 1150 1144 1156 1145
rect 1150 1140 1151 1144
rect 1155 1140 1156 1144
rect 1150 1139 1156 1140
rect 898 1135 904 1136
rect 898 1131 899 1135
rect 903 1131 904 1135
rect 898 1130 904 1131
rect 1010 1135 1016 1136
rect 1010 1131 1011 1135
rect 1015 1131 1016 1135
rect 1010 1130 1016 1131
rect 1018 1135 1024 1136
rect 1018 1131 1019 1135
rect 1023 1131 1024 1135
rect 1018 1130 1024 1131
rect 900 1120 902 1130
rect 1012 1120 1014 1130
rect 426 1119 432 1120
rect 530 1119 536 1120
rect 658 1119 664 1120
rect 822 1119 828 1120
rect 898 1119 904 1120
rect 1010 1119 1016 1120
rect 214 1118 220 1119
rect 214 1114 215 1118
rect 219 1114 220 1118
rect 214 1113 220 1114
rect 254 1118 260 1119
rect 254 1114 255 1118
rect 259 1114 260 1118
rect 254 1113 260 1114
rect 294 1118 300 1119
rect 294 1114 295 1118
rect 299 1114 300 1118
rect 294 1113 300 1114
rect 334 1118 340 1119
rect 334 1114 335 1118
rect 339 1114 340 1118
rect 334 1113 340 1114
rect 374 1118 380 1119
rect 374 1114 375 1118
rect 379 1114 380 1118
rect 414 1118 420 1119
rect 374 1113 380 1114
rect 386 1115 392 1116
rect 216 1107 218 1113
rect 256 1107 258 1113
rect 296 1107 298 1113
rect 336 1107 338 1113
rect 376 1107 378 1113
rect 386 1111 387 1115
rect 391 1111 392 1115
rect 414 1114 415 1118
rect 419 1114 420 1118
rect 426 1115 427 1119
rect 431 1115 432 1119
rect 426 1114 432 1115
rect 462 1118 468 1119
rect 462 1114 463 1118
rect 467 1114 468 1118
rect 414 1113 420 1114
rect 462 1113 468 1114
rect 518 1118 524 1119
rect 518 1114 519 1118
rect 523 1114 524 1118
rect 530 1115 531 1119
rect 535 1115 536 1119
rect 530 1114 536 1115
rect 582 1118 588 1119
rect 582 1114 583 1118
rect 587 1114 588 1118
rect 518 1113 524 1114
rect 582 1113 588 1114
rect 646 1118 652 1119
rect 646 1114 647 1118
rect 651 1114 652 1118
rect 658 1115 659 1119
rect 663 1115 664 1119
rect 658 1114 664 1115
rect 710 1118 716 1119
rect 710 1114 711 1118
rect 715 1114 716 1118
rect 646 1113 652 1114
rect 710 1113 716 1114
rect 766 1118 772 1119
rect 766 1114 767 1118
rect 771 1114 772 1118
rect 822 1115 823 1119
rect 827 1115 828 1119
rect 822 1114 828 1115
rect 830 1118 836 1119
rect 830 1114 831 1118
rect 835 1114 836 1118
rect 766 1113 772 1114
rect 830 1113 836 1114
rect 886 1118 892 1119
rect 886 1114 887 1118
rect 891 1114 892 1118
rect 898 1115 899 1119
rect 903 1115 904 1119
rect 898 1114 904 1115
rect 942 1118 948 1119
rect 942 1114 943 1118
rect 947 1114 948 1118
rect 886 1113 892 1114
rect 942 1113 948 1114
rect 998 1118 1004 1119
rect 998 1114 999 1118
rect 1003 1114 1004 1118
rect 1010 1115 1011 1119
rect 1015 1115 1016 1119
rect 1010 1114 1016 1115
rect 1054 1118 1060 1119
rect 1054 1114 1055 1118
rect 1059 1114 1060 1118
rect 998 1113 1004 1114
rect 1054 1113 1060 1114
rect 1102 1118 1108 1119
rect 1102 1114 1103 1118
rect 1107 1114 1108 1118
rect 1102 1113 1108 1114
rect 1150 1118 1156 1119
rect 1150 1114 1151 1118
rect 1155 1114 1156 1118
rect 1150 1113 1156 1114
rect 386 1110 392 1111
rect 207 1106 211 1107
rect 207 1101 211 1102
rect 215 1106 219 1107
rect 215 1101 219 1102
rect 247 1106 251 1107
rect 247 1101 251 1102
rect 255 1106 259 1107
rect 255 1101 259 1102
rect 287 1106 291 1107
rect 287 1101 291 1102
rect 295 1106 299 1107
rect 295 1101 299 1102
rect 327 1106 331 1107
rect 327 1101 331 1102
rect 335 1106 339 1107
rect 335 1101 339 1102
rect 367 1106 371 1107
rect 367 1101 371 1102
rect 375 1106 379 1107
rect 375 1101 379 1102
rect 194 1099 200 1100
rect 208 1099 210 1101
rect 248 1099 250 1101
rect 288 1099 290 1101
rect 328 1099 330 1101
rect 368 1099 370 1101
rect 134 1098 140 1099
rect 134 1094 135 1098
rect 139 1094 140 1098
rect 110 1093 116 1094
rect 134 1093 140 1094
rect 158 1098 164 1099
rect 158 1094 159 1098
rect 163 1094 164 1098
rect 158 1093 164 1094
rect 182 1098 188 1099
rect 182 1094 183 1098
rect 187 1094 188 1098
rect 194 1095 195 1099
rect 199 1095 200 1099
rect 194 1094 200 1095
rect 206 1098 212 1099
rect 206 1094 207 1098
rect 211 1094 212 1098
rect 246 1098 252 1099
rect 182 1093 188 1094
rect 206 1093 212 1094
rect 218 1095 224 1096
rect 110 1089 111 1093
rect 115 1089 116 1093
rect 218 1091 219 1095
rect 223 1091 224 1095
rect 246 1094 247 1098
rect 251 1094 252 1098
rect 246 1093 252 1094
rect 286 1098 292 1099
rect 286 1094 287 1098
rect 291 1094 292 1098
rect 286 1093 292 1094
rect 326 1098 332 1099
rect 326 1094 327 1098
rect 331 1094 332 1098
rect 326 1093 332 1094
rect 366 1098 372 1099
rect 366 1094 367 1098
rect 371 1094 372 1098
rect 366 1093 372 1094
rect 378 1095 384 1096
rect 378 1091 379 1095
rect 383 1091 384 1095
rect 218 1090 224 1091
rect 372 1090 384 1091
rect 110 1088 116 1089
rect 220 1077 222 1090
rect 372 1089 382 1090
rect 372 1084 374 1089
rect 388 1088 390 1110
rect 416 1107 418 1113
rect 464 1107 466 1113
rect 520 1107 522 1113
rect 584 1107 586 1113
rect 648 1107 650 1113
rect 712 1107 714 1113
rect 768 1107 770 1113
rect 832 1107 834 1113
rect 888 1107 890 1113
rect 944 1107 946 1113
rect 1000 1107 1002 1113
rect 1056 1107 1058 1113
rect 1104 1107 1106 1113
rect 1122 1107 1128 1108
rect 1152 1107 1154 1113
rect 1184 1112 1186 1150
rect 1191 1145 1195 1146
rect 1231 1150 1235 1151
rect 1231 1145 1235 1146
rect 1271 1150 1275 1151
rect 1282 1150 1288 1151
rect 1311 1150 1315 1151
rect 1271 1145 1275 1146
rect 1311 1145 1315 1146
rect 1351 1150 1355 1151
rect 1351 1145 1355 1146
rect 1190 1144 1196 1145
rect 1190 1140 1191 1144
rect 1195 1140 1196 1144
rect 1190 1139 1196 1140
rect 1230 1144 1236 1145
rect 1230 1140 1231 1144
rect 1235 1140 1236 1144
rect 1230 1139 1236 1140
rect 1270 1144 1276 1145
rect 1270 1140 1271 1144
rect 1275 1140 1276 1144
rect 1270 1139 1276 1140
rect 1310 1144 1316 1145
rect 1310 1140 1311 1144
rect 1315 1140 1316 1144
rect 1310 1139 1316 1140
rect 1350 1144 1356 1145
rect 1350 1140 1351 1144
rect 1355 1140 1356 1144
rect 1350 1139 1356 1140
rect 1364 1136 1366 1174
rect 1446 1173 1447 1177
rect 1451 1173 1452 1177
rect 1446 1172 1452 1173
rect 1446 1159 1452 1160
rect 1390 1156 1396 1157
rect 1414 1156 1420 1157
rect 1390 1152 1391 1156
rect 1395 1152 1396 1156
rect 1390 1151 1396 1152
rect 1402 1155 1408 1156
rect 1402 1151 1403 1155
rect 1407 1151 1408 1155
rect 1414 1152 1415 1156
rect 1419 1152 1420 1156
rect 1446 1155 1447 1159
rect 1451 1155 1452 1159
rect 1446 1154 1452 1155
rect 1414 1151 1420 1152
rect 1448 1151 1450 1154
rect 1391 1150 1395 1151
rect 1402 1150 1408 1151
rect 1415 1150 1419 1151
rect 1391 1145 1395 1146
rect 1390 1144 1396 1145
rect 1390 1140 1391 1144
rect 1395 1140 1396 1144
rect 1390 1139 1396 1140
rect 1362 1135 1368 1136
rect 1362 1131 1363 1135
rect 1367 1131 1368 1135
rect 1362 1130 1368 1131
rect 1404 1120 1406 1150
rect 1415 1145 1419 1146
rect 1447 1150 1451 1151
rect 1447 1145 1451 1146
rect 1414 1144 1420 1145
rect 1414 1140 1415 1144
rect 1419 1140 1420 1144
rect 1448 1142 1450 1145
rect 1414 1139 1420 1140
rect 1446 1141 1452 1142
rect 1446 1137 1447 1141
rect 1451 1137 1452 1141
rect 1446 1136 1452 1137
rect 1426 1127 1432 1128
rect 1426 1123 1427 1127
rect 1431 1123 1432 1127
rect 1426 1122 1432 1123
rect 1446 1123 1452 1124
rect 1402 1119 1408 1120
rect 1190 1118 1196 1119
rect 1190 1114 1191 1118
rect 1195 1114 1196 1118
rect 1190 1113 1196 1114
rect 1230 1118 1236 1119
rect 1230 1114 1231 1118
rect 1235 1114 1236 1118
rect 1230 1113 1236 1114
rect 1270 1118 1276 1119
rect 1270 1114 1271 1118
rect 1275 1114 1276 1118
rect 1270 1113 1276 1114
rect 1310 1118 1316 1119
rect 1310 1114 1311 1118
rect 1315 1114 1316 1118
rect 1310 1113 1316 1114
rect 1350 1118 1356 1119
rect 1350 1114 1351 1118
rect 1355 1114 1356 1118
rect 1350 1113 1356 1114
rect 1390 1118 1396 1119
rect 1390 1114 1391 1118
rect 1395 1114 1396 1118
rect 1402 1115 1403 1119
rect 1407 1115 1408 1119
rect 1402 1114 1408 1115
rect 1414 1118 1420 1119
rect 1414 1114 1415 1118
rect 1419 1114 1420 1118
rect 1390 1113 1396 1114
rect 1414 1113 1420 1114
rect 1182 1111 1188 1112
rect 1182 1107 1183 1111
rect 1187 1107 1188 1111
rect 1192 1107 1194 1113
rect 1232 1107 1234 1113
rect 1272 1107 1274 1113
rect 1312 1107 1314 1113
rect 1338 1107 1344 1108
rect 1352 1107 1354 1113
rect 1392 1107 1394 1113
rect 1416 1107 1418 1113
rect 407 1106 411 1107
rect 407 1101 411 1102
rect 415 1106 419 1107
rect 415 1101 419 1102
rect 455 1106 459 1107
rect 455 1101 459 1102
rect 463 1106 467 1107
rect 463 1101 467 1102
rect 503 1106 507 1107
rect 503 1101 507 1102
rect 519 1106 523 1107
rect 519 1101 523 1102
rect 559 1106 563 1107
rect 559 1101 563 1102
rect 583 1106 587 1107
rect 583 1101 587 1102
rect 607 1106 611 1107
rect 607 1101 611 1102
rect 647 1106 651 1107
rect 647 1101 651 1102
rect 655 1106 659 1107
rect 655 1101 659 1102
rect 703 1106 707 1107
rect 703 1101 707 1102
rect 711 1106 715 1107
rect 711 1101 715 1102
rect 743 1106 747 1107
rect 743 1101 747 1102
rect 767 1106 771 1107
rect 767 1101 771 1102
rect 791 1106 795 1107
rect 791 1101 795 1102
rect 831 1106 835 1107
rect 831 1101 835 1102
rect 839 1106 843 1107
rect 839 1101 843 1102
rect 887 1106 891 1107
rect 887 1101 891 1102
rect 943 1106 947 1107
rect 943 1101 947 1102
rect 999 1106 1003 1107
rect 999 1101 1003 1102
rect 1055 1106 1059 1107
rect 1055 1101 1059 1102
rect 1103 1106 1107 1107
rect 1103 1101 1107 1102
rect 1111 1106 1115 1107
rect 1122 1103 1123 1107
rect 1127 1103 1128 1107
rect 1122 1102 1128 1103
rect 1151 1106 1155 1107
rect 1111 1101 1115 1102
rect 408 1099 410 1101
rect 456 1099 458 1101
rect 504 1099 506 1101
rect 560 1099 562 1101
rect 608 1099 610 1101
rect 656 1099 658 1101
rect 704 1099 706 1101
rect 744 1099 746 1101
rect 792 1099 794 1101
rect 840 1099 842 1101
rect 888 1099 890 1101
rect 944 1099 946 1101
rect 1000 1099 1002 1101
rect 1056 1099 1058 1101
rect 1112 1099 1114 1101
rect 406 1098 412 1099
rect 406 1094 407 1098
rect 411 1094 412 1098
rect 406 1093 412 1094
rect 454 1098 460 1099
rect 454 1094 455 1098
rect 459 1094 460 1098
rect 454 1093 460 1094
rect 502 1098 508 1099
rect 502 1094 503 1098
rect 507 1094 508 1098
rect 502 1093 508 1094
rect 558 1098 564 1099
rect 558 1094 559 1098
rect 563 1094 564 1098
rect 558 1093 564 1094
rect 606 1098 612 1099
rect 606 1094 607 1098
rect 611 1094 612 1098
rect 654 1098 660 1099
rect 606 1093 612 1094
rect 618 1095 624 1096
rect 618 1091 619 1095
rect 623 1091 624 1095
rect 654 1094 655 1098
rect 659 1094 660 1098
rect 654 1093 660 1094
rect 702 1098 708 1099
rect 702 1094 703 1098
rect 707 1094 708 1098
rect 702 1093 708 1094
rect 742 1098 748 1099
rect 742 1094 743 1098
rect 747 1094 748 1098
rect 742 1093 748 1094
rect 790 1098 796 1099
rect 790 1094 791 1098
rect 795 1094 796 1098
rect 790 1093 796 1094
rect 838 1098 844 1099
rect 838 1094 839 1098
rect 843 1094 844 1098
rect 838 1093 844 1094
rect 886 1098 892 1099
rect 886 1094 887 1098
rect 891 1094 892 1098
rect 886 1093 892 1094
rect 942 1098 948 1099
rect 942 1094 943 1098
rect 947 1094 948 1098
rect 942 1093 948 1094
rect 998 1098 1004 1099
rect 998 1094 999 1098
rect 1003 1094 1004 1098
rect 1054 1098 1060 1099
rect 998 1093 1004 1094
rect 1010 1095 1016 1096
rect 618 1090 624 1091
rect 1010 1091 1011 1095
rect 1015 1091 1016 1095
rect 1054 1094 1055 1098
rect 1059 1094 1060 1098
rect 1054 1093 1060 1094
rect 1110 1098 1116 1099
rect 1110 1094 1111 1098
rect 1115 1094 1116 1098
rect 1110 1093 1116 1094
rect 1010 1090 1016 1091
rect 366 1083 374 1084
rect 366 1079 367 1083
rect 371 1081 374 1083
rect 386 1087 392 1088
rect 386 1083 387 1087
rect 391 1083 392 1087
rect 386 1082 392 1083
rect 371 1079 372 1081
rect 366 1078 372 1079
rect 147 1076 151 1077
rect 110 1075 116 1076
rect 110 1071 111 1075
rect 115 1071 116 1075
rect 143 1075 147 1076
rect 110 1070 116 1071
rect 134 1072 140 1073
rect 112 1067 114 1070
rect 134 1068 135 1072
rect 139 1068 140 1072
rect 143 1071 144 1075
rect 219 1076 223 1077
rect 148 1071 151 1072
rect 158 1072 164 1073
rect 143 1070 149 1071
rect 134 1067 140 1068
rect 158 1068 159 1072
rect 163 1068 164 1072
rect 158 1067 164 1068
rect 182 1072 188 1073
rect 182 1068 183 1072
rect 187 1068 188 1072
rect 182 1067 188 1068
rect 206 1072 212 1073
rect 206 1068 207 1072
rect 211 1068 212 1072
rect 219 1071 223 1072
rect 246 1072 252 1073
rect 206 1067 212 1068
rect 246 1068 247 1072
rect 251 1068 252 1072
rect 246 1067 252 1068
rect 286 1072 292 1073
rect 326 1072 332 1073
rect 286 1068 287 1072
rect 291 1068 292 1072
rect 286 1067 292 1068
rect 298 1071 304 1072
rect 298 1067 299 1071
rect 303 1067 304 1071
rect 326 1068 327 1072
rect 331 1068 332 1072
rect 326 1067 332 1068
rect 366 1072 372 1073
rect 366 1068 367 1072
rect 371 1068 372 1072
rect 366 1067 372 1068
rect 406 1072 412 1073
rect 406 1068 407 1072
rect 411 1068 412 1072
rect 406 1067 412 1068
rect 454 1072 460 1073
rect 454 1068 455 1072
rect 459 1068 460 1072
rect 454 1067 460 1068
rect 502 1072 508 1073
rect 502 1068 503 1072
rect 507 1068 508 1072
rect 502 1067 508 1068
rect 558 1072 564 1073
rect 558 1068 559 1072
rect 563 1068 564 1072
rect 558 1067 564 1068
rect 606 1072 612 1073
rect 606 1068 607 1072
rect 611 1068 612 1072
rect 606 1067 612 1068
rect 111 1066 115 1067
rect 111 1061 115 1062
rect 135 1066 139 1067
rect 135 1061 139 1062
rect 159 1066 163 1067
rect 159 1061 163 1062
rect 183 1066 187 1067
rect 183 1061 187 1062
rect 207 1066 211 1067
rect 207 1061 211 1062
rect 231 1066 235 1067
rect 231 1061 235 1062
rect 247 1066 251 1067
rect 247 1061 251 1062
rect 271 1066 275 1067
rect 271 1061 275 1062
rect 287 1066 291 1067
rect 298 1066 304 1067
rect 311 1066 315 1067
rect 287 1061 291 1062
rect 112 1058 114 1061
rect 134 1060 140 1061
rect 110 1057 116 1058
rect 110 1053 111 1057
rect 115 1053 116 1057
rect 134 1056 135 1060
rect 139 1056 140 1060
rect 134 1055 140 1056
rect 158 1060 164 1061
rect 158 1056 159 1060
rect 163 1056 164 1060
rect 158 1055 164 1056
rect 182 1060 188 1061
rect 182 1056 183 1060
rect 187 1056 188 1060
rect 182 1055 188 1056
rect 206 1060 212 1061
rect 206 1056 207 1060
rect 211 1056 212 1060
rect 206 1055 212 1056
rect 230 1060 236 1061
rect 230 1056 231 1060
rect 235 1056 236 1060
rect 230 1055 236 1056
rect 270 1060 276 1061
rect 270 1056 271 1060
rect 275 1056 276 1060
rect 270 1055 276 1056
rect 110 1052 116 1053
rect 170 1051 176 1052
rect 170 1047 171 1051
rect 175 1047 176 1051
rect 170 1046 176 1047
rect 194 1051 200 1052
rect 194 1047 195 1051
rect 199 1047 200 1051
rect 194 1046 200 1047
rect 218 1051 224 1052
rect 218 1047 219 1051
rect 223 1047 224 1051
rect 218 1046 224 1047
rect 242 1051 248 1052
rect 242 1047 243 1051
rect 247 1047 248 1051
rect 242 1046 248 1047
rect 147 1044 151 1045
rect 110 1039 116 1040
rect 147 1039 151 1040
rect 110 1035 111 1039
rect 115 1035 116 1039
rect 148 1036 150 1039
rect 172 1036 174 1046
rect 196 1036 198 1046
rect 220 1036 222 1046
rect 244 1036 246 1046
rect 300 1045 302 1066
rect 311 1061 315 1062
rect 327 1066 331 1067
rect 327 1061 331 1062
rect 351 1066 355 1067
rect 351 1061 355 1062
rect 367 1066 371 1067
rect 367 1061 371 1062
rect 391 1066 395 1067
rect 391 1061 395 1062
rect 407 1066 411 1067
rect 407 1061 411 1062
rect 431 1066 435 1067
rect 431 1061 435 1062
rect 455 1066 459 1067
rect 455 1061 459 1062
rect 471 1066 475 1067
rect 471 1061 475 1062
rect 503 1066 507 1067
rect 503 1061 507 1062
rect 511 1066 515 1067
rect 511 1061 515 1062
rect 551 1066 555 1067
rect 551 1061 555 1062
rect 559 1066 563 1067
rect 559 1061 563 1062
rect 591 1066 595 1067
rect 591 1061 595 1062
rect 607 1066 611 1067
rect 607 1061 611 1062
rect 310 1060 316 1061
rect 310 1056 311 1060
rect 315 1056 316 1060
rect 310 1055 316 1056
rect 350 1060 356 1061
rect 350 1056 351 1060
rect 355 1056 356 1060
rect 350 1055 356 1056
rect 390 1060 396 1061
rect 390 1056 391 1060
rect 395 1056 396 1060
rect 390 1055 396 1056
rect 430 1060 436 1061
rect 430 1056 431 1060
rect 435 1056 436 1060
rect 430 1055 436 1056
rect 470 1060 476 1061
rect 470 1056 471 1060
rect 475 1056 476 1060
rect 470 1055 476 1056
rect 510 1060 516 1061
rect 510 1056 511 1060
rect 515 1056 516 1060
rect 510 1055 516 1056
rect 550 1060 556 1061
rect 550 1056 551 1060
rect 555 1056 556 1060
rect 550 1055 556 1056
rect 590 1060 596 1061
rect 590 1056 591 1060
rect 595 1056 596 1060
rect 590 1055 596 1056
rect 620 1052 622 1090
rect 654 1072 660 1073
rect 702 1072 708 1073
rect 654 1068 655 1072
rect 659 1068 660 1072
rect 654 1067 660 1068
rect 694 1071 700 1072
rect 694 1067 695 1071
rect 699 1067 700 1071
rect 702 1068 703 1072
rect 707 1068 708 1072
rect 702 1067 708 1068
rect 742 1072 748 1073
rect 742 1068 743 1072
rect 747 1068 748 1072
rect 742 1067 748 1068
rect 790 1072 796 1073
rect 790 1068 791 1072
rect 795 1068 796 1072
rect 790 1067 796 1068
rect 838 1072 844 1073
rect 838 1068 839 1072
rect 843 1068 844 1072
rect 838 1067 844 1068
rect 886 1072 892 1073
rect 886 1068 887 1072
rect 891 1068 892 1072
rect 886 1067 892 1068
rect 942 1072 948 1073
rect 942 1068 943 1072
rect 947 1068 948 1072
rect 942 1067 948 1068
rect 998 1072 1004 1073
rect 998 1068 999 1072
rect 1003 1068 1004 1072
rect 998 1067 1004 1068
rect 631 1066 635 1067
rect 631 1061 635 1062
rect 655 1066 659 1067
rect 655 1061 659 1062
rect 671 1066 675 1067
rect 694 1066 700 1067
rect 703 1066 707 1067
rect 671 1061 675 1062
rect 630 1060 636 1061
rect 630 1056 631 1060
rect 635 1056 636 1060
rect 630 1055 636 1056
rect 670 1060 676 1061
rect 670 1056 671 1060
rect 675 1056 676 1060
rect 670 1055 676 1056
rect 322 1051 328 1052
rect 322 1047 323 1051
rect 327 1047 328 1051
rect 322 1046 328 1047
rect 618 1051 624 1052
rect 618 1047 619 1051
rect 623 1047 624 1051
rect 618 1046 624 1047
rect 299 1044 303 1045
rect 299 1039 303 1040
rect 324 1036 326 1046
rect 696 1037 698 1066
rect 703 1061 707 1062
rect 711 1066 715 1067
rect 711 1061 715 1062
rect 743 1066 747 1067
rect 743 1061 747 1062
rect 783 1066 787 1067
rect 783 1061 787 1062
rect 791 1066 795 1067
rect 791 1061 795 1062
rect 823 1066 827 1067
rect 823 1061 827 1062
rect 839 1066 843 1067
rect 839 1061 843 1062
rect 871 1066 875 1067
rect 871 1061 875 1062
rect 887 1066 891 1067
rect 887 1061 891 1062
rect 919 1066 923 1067
rect 919 1061 923 1062
rect 943 1066 947 1067
rect 943 1061 947 1062
rect 975 1066 979 1067
rect 975 1061 979 1062
rect 999 1066 1003 1067
rect 999 1061 1003 1062
rect 710 1060 716 1061
rect 710 1056 711 1060
rect 715 1056 716 1060
rect 710 1055 716 1056
rect 742 1060 748 1061
rect 742 1056 743 1060
rect 747 1056 748 1060
rect 742 1055 748 1056
rect 782 1060 788 1061
rect 782 1056 783 1060
rect 787 1056 788 1060
rect 782 1055 788 1056
rect 822 1060 828 1061
rect 822 1056 823 1060
rect 827 1056 828 1060
rect 822 1055 828 1056
rect 870 1060 876 1061
rect 870 1056 871 1060
rect 875 1056 876 1060
rect 870 1055 876 1056
rect 918 1060 924 1061
rect 918 1056 919 1060
rect 923 1056 924 1060
rect 918 1055 924 1056
rect 974 1060 980 1061
rect 1012 1060 1014 1090
rect 1124 1080 1126 1102
rect 1151 1101 1155 1102
rect 1167 1106 1171 1107
rect 1182 1106 1188 1107
rect 1191 1106 1195 1107
rect 1167 1101 1171 1102
rect 1191 1101 1195 1102
rect 1215 1106 1219 1107
rect 1215 1101 1219 1102
rect 1231 1106 1235 1107
rect 1231 1101 1235 1102
rect 1271 1106 1275 1107
rect 1271 1101 1275 1102
rect 1311 1106 1315 1107
rect 1311 1101 1315 1102
rect 1327 1106 1331 1107
rect 1338 1103 1339 1107
rect 1343 1103 1344 1107
rect 1338 1102 1344 1103
rect 1351 1106 1355 1107
rect 1327 1101 1331 1102
rect 1168 1099 1170 1101
rect 1216 1099 1218 1101
rect 1272 1099 1274 1101
rect 1328 1099 1330 1101
rect 1166 1098 1172 1099
rect 1166 1094 1167 1098
rect 1171 1094 1172 1098
rect 1166 1093 1172 1094
rect 1214 1098 1220 1099
rect 1214 1094 1215 1098
rect 1219 1094 1220 1098
rect 1270 1098 1276 1099
rect 1214 1093 1220 1094
rect 1262 1095 1268 1096
rect 1262 1091 1263 1095
rect 1267 1091 1268 1095
rect 1270 1094 1271 1098
rect 1275 1094 1276 1098
rect 1270 1093 1276 1094
rect 1326 1098 1332 1099
rect 1326 1094 1327 1098
rect 1331 1094 1332 1098
rect 1326 1093 1332 1094
rect 1262 1090 1268 1091
rect 1138 1083 1144 1084
rect 1122 1079 1128 1080
rect 1122 1075 1123 1079
rect 1127 1075 1128 1079
rect 1138 1079 1139 1083
rect 1143 1079 1144 1083
rect 1138 1078 1144 1079
rect 1122 1074 1128 1075
rect 1054 1072 1060 1073
rect 1054 1068 1055 1072
rect 1059 1068 1060 1072
rect 1054 1067 1060 1068
rect 1110 1072 1116 1073
rect 1110 1068 1111 1072
rect 1115 1068 1116 1072
rect 1110 1067 1116 1068
rect 1031 1066 1035 1067
rect 1031 1061 1035 1062
rect 1055 1066 1059 1067
rect 1055 1061 1059 1062
rect 1079 1066 1083 1067
rect 1079 1061 1083 1062
rect 1111 1066 1115 1067
rect 1111 1061 1115 1062
rect 1127 1066 1131 1067
rect 1127 1061 1131 1062
rect 1030 1060 1036 1061
rect 974 1056 975 1060
rect 979 1056 980 1060
rect 974 1055 980 1056
rect 1010 1059 1016 1060
rect 1010 1055 1011 1059
rect 1015 1055 1016 1059
rect 1030 1056 1031 1060
rect 1035 1056 1036 1060
rect 1030 1055 1036 1056
rect 1078 1060 1084 1061
rect 1078 1056 1079 1060
rect 1083 1056 1084 1060
rect 1078 1055 1084 1056
rect 1126 1060 1132 1061
rect 1126 1056 1127 1060
rect 1131 1056 1132 1060
rect 1126 1055 1132 1056
rect 1010 1054 1016 1055
rect 774 1051 780 1052
rect 774 1047 775 1051
rect 779 1047 780 1051
rect 774 1046 780 1047
rect 882 1051 888 1052
rect 882 1047 883 1051
rect 887 1047 888 1051
rect 882 1046 888 1047
rect 695 1036 699 1037
rect 146 1035 152 1036
rect 170 1035 176 1036
rect 194 1035 200 1036
rect 218 1035 224 1036
rect 242 1035 248 1036
rect 322 1035 328 1036
rect 110 1034 116 1035
rect 134 1034 140 1035
rect 112 1027 114 1034
rect 134 1030 135 1034
rect 139 1030 140 1034
rect 146 1031 147 1035
rect 151 1031 152 1035
rect 146 1030 152 1031
rect 158 1034 164 1035
rect 158 1030 159 1034
rect 163 1030 164 1034
rect 170 1031 171 1035
rect 175 1031 176 1035
rect 170 1030 176 1031
rect 182 1034 188 1035
rect 182 1030 183 1034
rect 187 1030 188 1034
rect 194 1031 195 1035
rect 199 1031 200 1035
rect 194 1030 200 1031
rect 206 1034 212 1035
rect 206 1030 207 1034
rect 211 1030 212 1034
rect 218 1031 219 1035
rect 223 1031 224 1035
rect 218 1030 224 1031
rect 230 1034 236 1035
rect 230 1030 231 1034
rect 235 1030 236 1034
rect 242 1031 243 1035
rect 247 1031 248 1035
rect 242 1030 248 1031
rect 270 1034 276 1035
rect 270 1030 271 1034
rect 275 1030 276 1034
rect 134 1029 140 1030
rect 158 1029 164 1030
rect 182 1029 188 1030
rect 206 1029 212 1030
rect 230 1029 236 1030
rect 270 1029 276 1030
rect 310 1034 316 1035
rect 310 1030 311 1034
rect 315 1030 316 1034
rect 322 1031 323 1035
rect 327 1031 328 1035
rect 322 1030 328 1031
rect 350 1034 356 1035
rect 350 1030 351 1034
rect 355 1030 356 1034
rect 310 1029 316 1030
rect 350 1029 356 1030
rect 390 1034 396 1035
rect 390 1030 391 1034
rect 395 1030 396 1034
rect 390 1029 396 1030
rect 430 1034 436 1035
rect 430 1030 431 1034
rect 435 1030 436 1034
rect 430 1029 436 1030
rect 470 1034 476 1035
rect 470 1030 471 1034
rect 475 1030 476 1034
rect 470 1029 476 1030
rect 510 1034 516 1035
rect 510 1030 511 1034
rect 515 1030 516 1034
rect 510 1029 516 1030
rect 550 1034 556 1035
rect 550 1030 551 1034
rect 555 1030 556 1034
rect 550 1029 556 1030
rect 590 1034 596 1035
rect 590 1030 591 1034
rect 595 1030 596 1034
rect 630 1034 636 1035
rect 590 1029 596 1030
rect 602 1031 608 1032
rect 136 1027 138 1029
rect 160 1027 162 1029
rect 184 1027 186 1029
rect 208 1027 210 1029
rect 232 1027 234 1029
rect 272 1027 274 1029
rect 312 1027 314 1029
rect 352 1027 354 1029
rect 392 1027 394 1029
rect 432 1027 434 1029
rect 472 1027 474 1029
rect 512 1027 514 1029
rect 538 1027 544 1028
rect 552 1027 554 1029
rect 592 1027 594 1029
rect 602 1027 603 1031
rect 607 1027 608 1031
rect 630 1030 631 1034
rect 635 1030 636 1034
rect 630 1029 636 1030
rect 670 1034 676 1035
rect 670 1030 671 1034
rect 675 1030 676 1034
rect 695 1031 699 1032
rect 710 1034 716 1035
rect 670 1029 676 1030
rect 710 1030 711 1034
rect 715 1030 716 1034
rect 710 1029 716 1030
rect 742 1034 748 1035
rect 742 1030 743 1034
rect 747 1030 748 1034
rect 742 1029 748 1030
rect 632 1027 634 1029
rect 672 1027 674 1029
rect 712 1027 714 1029
rect 744 1027 746 1029
rect 111 1026 115 1027
rect 111 1021 115 1022
rect 135 1026 139 1027
rect 135 1021 139 1022
rect 159 1026 163 1027
rect 159 1021 163 1022
rect 183 1026 187 1027
rect 183 1021 187 1022
rect 207 1026 211 1027
rect 207 1021 211 1022
rect 231 1026 235 1027
rect 231 1021 235 1022
rect 263 1026 267 1027
rect 263 1021 267 1022
rect 271 1026 275 1027
rect 271 1021 275 1022
rect 303 1026 307 1027
rect 303 1021 307 1022
rect 311 1026 315 1027
rect 311 1021 315 1022
rect 343 1026 347 1027
rect 343 1021 347 1022
rect 351 1026 355 1027
rect 351 1021 355 1022
rect 383 1026 387 1027
rect 383 1021 387 1022
rect 391 1026 395 1027
rect 391 1021 395 1022
rect 431 1026 435 1027
rect 431 1021 435 1022
rect 471 1026 475 1027
rect 471 1021 475 1022
rect 479 1026 483 1027
rect 479 1021 483 1022
rect 511 1026 515 1027
rect 511 1021 515 1022
rect 527 1026 531 1027
rect 538 1023 539 1027
rect 543 1023 544 1027
rect 538 1022 544 1023
rect 551 1026 555 1027
rect 527 1021 531 1022
rect 112 1014 114 1021
rect 160 1019 162 1021
rect 184 1019 186 1021
rect 208 1019 210 1021
rect 232 1019 234 1021
rect 264 1019 266 1021
rect 304 1019 306 1021
rect 344 1019 346 1021
rect 384 1019 386 1021
rect 432 1019 434 1021
rect 480 1019 482 1021
rect 528 1019 530 1021
rect 158 1018 164 1019
rect 158 1014 159 1018
rect 163 1014 164 1018
rect 110 1013 116 1014
rect 158 1013 164 1014
rect 182 1018 188 1019
rect 182 1014 183 1018
rect 187 1014 188 1018
rect 182 1013 188 1014
rect 206 1018 212 1019
rect 206 1014 207 1018
rect 211 1014 212 1018
rect 206 1013 212 1014
rect 230 1018 236 1019
rect 230 1014 231 1018
rect 235 1014 236 1018
rect 230 1013 236 1014
rect 262 1018 268 1019
rect 262 1014 263 1018
rect 267 1014 268 1018
rect 262 1013 268 1014
rect 302 1018 308 1019
rect 302 1014 303 1018
rect 307 1014 308 1018
rect 302 1013 308 1014
rect 342 1018 348 1019
rect 342 1014 343 1018
rect 347 1014 348 1018
rect 342 1013 348 1014
rect 382 1018 388 1019
rect 382 1014 383 1018
rect 387 1014 388 1018
rect 430 1018 436 1019
rect 382 1013 388 1014
rect 410 1015 416 1016
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 410 1011 411 1015
rect 415 1011 416 1015
rect 430 1014 431 1018
rect 435 1014 436 1018
rect 430 1013 436 1014
rect 478 1018 484 1019
rect 478 1014 479 1018
rect 483 1014 484 1018
rect 478 1013 484 1014
rect 526 1018 532 1019
rect 526 1014 527 1018
rect 531 1014 532 1018
rect 526 1013 532 1014
rect 410 1010 416 1011
rect 110 1008 116 1009
rect 219 996 223 997
rect 355 996 359 997
rect 110 995 116 996
rect 110 991 111 995
rect 115 991 116 995
rect 110 990 116 991
rect 158 992 164 993
rect 112 987 114 990
rect 158 988 159 992
rect 163 988 164 992
rect 158 987 164 988
rect 182 992 188 993
rect 182 988 183 992
rect 187 988 188 992
rect 182 987 188 988
rect 206 992 212 993
rect 206 988 207 992
rect 211 988 212 992
rect 219 991 223 992
rect 230 992 236 993
rect 206 987 212 988
rect 111 986 115 987
rect 111 981 115 982
rect 159 986 163 987
rect 159 981 163 982
rect 183 986 187 987
rect 183 981 187 982
rect 207 986 211 987
rect 207 981 211 982
rect 112 978 114 981
rect 206 980 212 981
rect 110 977 116 978
rect 110 973 111 977
rect 115 973 116 977
rect 206 976 207 980
rect 211 976 212 980
rect 206 975 212 976
rect 110 972 116 973
rect 110 959 116 960
rect 110 955 111 959
rect 115 955 116 959
rect 220 956 222 991
rect 230 988 231 992
rect 235 988 236 992
rect 230 987 236 988
rect 262 992 268 993
rect 262 988 263 992
rect 267 988 268 992
rect 262 987 268 988
rect 302 992 308 993
rect 302 988 303 992
rect 307 988 308 992
rect 302 987 308 988
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 354 991 355 996
rect 359 991 360 996
rect 354 990 360 991
rect 382 992 388 993
rect 342 987 348 988
rect 382 988 383 992
rect 387 988 388 992
rect 382 987 388 988
rect 231 986 235 987
rect 231 981 235 982
rect 255 986 259 987
rect 255 981 259 982
rect 263 986 267 987
rect 263 981 267 982
rect 287 986 291 987
rect 287 981 291 982
rect 303 986 307 987
rect 303 981 307 982
rect 327 986 331 987
rect 327 981 331 982
rect 343 986 347 987
rect 343 981 347 982
rect 375 986 379 987
rect 375 981 379 982
rect 383 986 387 987
rect 383 981 387 982
rect 230 980 236 981
rect 230 976 231 980
rect 235 976 236 980
rect 230 975 236 976
rect 254 980 260 981
rect 254 976 255 980
rect 259 976 260 980
rect 254 975 260 976
rect 286 980 292 981
rect 286 976 287 980
rect 291 976 292 980
rect 286 975 292 976
rect 326 980 332 981
rect 326 976 327 980
rect 331 976 332 980
rect 326 975 332 976
rect 374 980 380 981
rect 374 976 375 980
rect 379 976 380 980
rect 374 975 380 976
rect 412 972 414 1010
rect 540 996 542 1022
rect 551 1021 555 1022
rect 575 1026 579 1027
rect 575 1021 579 1022
rect 591 1026 595 1027
rect 602 1026 608 1027
rect 623 1026 627 1027
rect 591 1021 595 1022
rect 576 1019 578 1021
rect 574 1018 580 1019
rect 574 1014 575 1018
rect 579 1014 580 1018
rect 574 1013 580 1014
rect 604 1008 606 1026
rect 623 1021 627 1022
rect 631 1026 635 1027
rect 631 1021 635 1022
rect 671 1026 675 1027
rect 671 1021 675 1022
rect 711 1026 715 1027
rect 711 1021 715 1022
rect 719 1026 723 1027
rect 719 1021 723 1022
rect 743 1026 747 1027
rect 743 1021 747 1022
rect 767 1026 771 1027
rect 776 1024 778 1046
rect 795 1036 799 1037
rect 884 1036 886 1046
rect 1002 1043 1008 1044
rect 1002 1039 1003 1043
rect 1007 1039 1008 1043
rect 1002 1038 1008 1039
rect 782 1034 788 1035
rect 782 1030 783 1034
rect 787 1030 788 1034
rect 794 1031 795 1036
rect 799 1031 800 1036
rect 882 1035 888 1036
rect 794 1030 800 1031
rect 822 1034 828 1035
rect 822 1030 823 1034
rect 827 1030 828 1034
rect 870 1034 876 1035
rect 782 1029 788 1030
rect 822 1029 828 1030
rect 834 1031 840 1032
rect 784 1027 786 1029
rect 824 1027 826 1029
rect 834 1027 835 1031
rect 839 1027 840 1031
rect 870 1030 871 1034
rect 875 1030 876 1034
rect 882 1031 883 1035
rect 887 1031 888 1035
rect 882 1030 888 1031
rect 918 1034 924 1035
rect 918 1030 919 1034
rect 923 1030 924 1034
rect 870 1029 876 1030
rect 918 1029 924 1030
rect 974 1034 980 1035
rect 974 1030 975 1034
rect 979 1030 980 1034
rect 974 1029 980 1030
rect 872 1027 874 1029
rect 920 1027 922 1029
rect 976 1027 978 1029
rect 783 1026 787 1027
rect 767 1021 771 1022
rect 774 1023 780 1024
rect 624 1019 626 1021
rect 672 1019 674 1021
rect 720 1019 722 1021
rect 768 1019 770 1021
rect 774 1019 775 1023
rect 779 1019 780 1023
rect 783 1021 787 1022
rect 823 1026 827 1027
rect 834 1026 840 1027
rect 871 1026 875 1027
rect 823 1021 827 1022
rect 824 1019 826 1021
rect 622 1018 628 1019
rect 622 1014 623 1018
rect 627 1014 628 1018
rect 622 1013 628 1014
rect 670 1018 676 1019
rect 670 1014 671 1018
rect 675 1014 676 1018
rect 670 1013 676 1014
rect 718 1018 724 1019
rect 718 1014 719 1018
rect 723 1014 724 1018
rect 718 1013 724 1014
rect 766 1018 772 1019
rect 774 1018 780 1019
rect 822 1018 828 1019
rect 766 1014 767 1018
rect 771 1014 772 1018
rect 766 1013 772 1014
rect 822 1014 823 1018
rect 827 1014 828 1018
rect 822 1013 828 1014
rect 836 1008 838 1026
rect 871 1021 875 1022
rect 879 1026 883 1027
rect 879 1021 883 1022
rect 919 1026 923 1027
rect 919 1021 923 1022
rect 935 1026 939 1027
rect 935 1021 939 1022
rect 975 1026 979 1027
rect 975 1021 979 1022
rect 991 1026 995 1027
rect 991 1021 995 1022
rect 880 1019 882 1021
rect 936 1019 938 1021
rect 992 1019 994 1021
rect 1004 1020 1006 1038
rect 1140 1036 1142 1078
rect 1166 1072 1172 1073
rect 1166 1068 1167 1072
rect 1171 1068 1172 1072
rect 1166 1067 1172 1068
rect 1214 1072 1220 1073
rect 1214 1068 1215 1072
rect 1219 1068 1220 1072
rect 1214 1067 1220 1068
rect 1167 1066 1171 1067
rect 1167 1061 1171 1062
rect 1175 1066 1179 1067
rect 1175 1061 1179 1062
rect 1215 1066 1219 1067
rect 1215 1061 1219 1062
rect 1223 1066 1227 1067
rect 1223 1061 1227 1062
rect 1174 1060 1180 1061
rect 1174 1056 1175 1060
rect 1179 1056 1180 1060
rect 1174 1055 1180 1056
rect 1222 1060 1228 1061
rect 1222 1056 1223 1060
rect 1227 1056 1228 1060
rect 1222 1055 1228 1056
rect 1234 1051 1240 1052
rect 1234 1047 1235 1051
rect 1239 1047 1240 1051
rect 1234 1046 1240 1047
rect 1236 1036 1238 1046
rect 1264 1044 1266 1090
rect 1340 1076 1342 1102
rect 1351 1101 1355 1102
rect 1383 1106 1387 1107
rect 1383 1101 1387 1102
rect 1391 1106 1395 1107
rect 1391 1101 1395 1102
rect 1415 1106 1419 1107
rect 1415 1101 1419 1102
rect 1384 1099 1386 1101
rect 1416 1099 1418 1101
rect 1428 1100 1430 1122
rect 1446 1119 1447 1123
rect 1451 1119 1452 1123
rect 1446 1118 1452 1119
rect 1448 1107 1450 1118
rect 1447 1106 1451 1107
rect 1447 1101 1451 1102
rect 1426 1099 1432 1100
rect 1382 1098 1388 1099
rect 1382 1094 1383 1098
rect 1387 1094 1388 1098
rect 1382 1093 1388 1094
rect 1414 1098 1420 1099
rect 1414 1094 1415 1098
rect 1419 1094 1420 1098
rect 1426 1095 1427 1099
rect 1431 1095 1432 1099
rect 1426 1094 1432 1095
rect 1448 1094 1450 1101
rect 1414 1093 1420 1094
rect 1446 1093 1452 1094
rect 1446 1089 1447 1093
rect 1451 1089 1452 1093
rect 1446 1088 1452 1089
rect 1338 1075 1344 1076
rect 1270 1072 1276 1073
rect 1270 1068 1271 1072
rect 1275 1068 1276 1072
rect 1270 1067 1276 1068
rect 1326 1072 1332 1073
rect 1326 1068 1327 1072
rect 1331 1068 1332 1072
rect 1338 1071 1339 1075
rect 1343 1071 1344 1075
rect 1446 1075 1452 1076
rect 1338 1070 1344 1071
rect 1382 1072 1388 1073
rect 1326 1067 1332 1068
rect 1382 1068 1383 1072
rect 1387 1068 1388 1072
rect 1382 1067 1388 1068
rect 1414 1072 1420 1073
rect 1414 1068 1415 1072
rect 1419 1068 1420 1072
rect 1414 1067 1420 1068
rect 1426 1071 1432 1072
rect 1426 1067 1427 1071
rect 1431 1067 1432 1071
rect 1446 1071 1447 1075
rect 1451 1071 1452 1075
rect 1446 1070 1452 1071
rect 1448 1067 1450 1070
rect 1271 1066 1275 1067
rect 1271 1061 1275 1062
rect 1327 1066 1331 1067
rect 1327 1061 1331 1062
rect 1383 1066 1387 1067
rect 1383 1061 1387 1062
rect 1415 1066 1419 1067
rect 1426 1066 1432 1067
rect 1447 1066 1451 1067
rect 1415 1061 1419 1062
rect 1270 1060 1276 1061
rect 1270 1056 1271 1060
rect 1275 1056 1276 1060
rect 1270 1055 1276 1056
rect 1326 1060 1332 1061
rect 1326 1056 1327 1060
rect 1331 1056 1332 1060
rect 1326 1055 1332 1056
rect 1382 1060 1388 1061
rect 1382 1056 1383 1060
rect 1387 1056 1388 1060
rect 1382 1055 1388 1056
rect 1414 1060 1420 1061
rect 1414 1056 1415 1060
rect 1419 1056 1420 1060
rect 1414 1055 1420 1056
rect 1338 1051 1344 1052
rect 1338 1047 1339 1051
rect 1343 1047 1344 1051
rect 1338 1046 1344 1047
rect 1262 1043 1268 1044
rect 1262 1039 1263 1043
rect 1267 1039 1268 1043
rect 1262 1038 1268 1039
rect 1340 1036 1342 1046
rect 1394 1043 1400 1044
rect 1394 1039 1395 1043
rect 1399 1039 1400 1043
rect 1394 1038 1400 1039
rect 1138 1035 1144 1036
rect 1234 1035 1240 1036
rect 1338 1035 1344 1036
rect 1030 1034 1036 1035
rect 1030 1030 1031 1034
rect 1035 1030 1036 1034
rect 1030 1029 1036 1030
rect 1078 1034 1084 1035
rect 1078 1030 1079 1034
rect 1083 1030 1084 1034
rect 1078 1029 1084 1030
rect 1126 1034 1132 1035
rect 1126 1030 1127 1034
rect 1131 1030 1132 1034
rect 1138 1031 1139 1035
rect 1143 1031 1144 1035
rect 1138 1030 1144 1031
rect 1174 1034 1180 1035
rect 1174 1030 1175 1034
rect 1179 1030 1180 1034
rect 1222 1034 1228 1035
rect 1126 1029 1132 1030
rect 1174 1029 1180 1030
rect 1186 1031 1192 1032
rect 1032 1027 1034 1029
rect 1080 1027 1082 1029
rect 1128 1027 1130 1029
rect 1176 1027 1178 1029
rect 1186 1027 1187 1031
rect 1191 1027 1192 1031
rect 1222 1030 1223 1034
rect 1227 1030 1228 1034
rect 1234 1031 1235 1035
rect 1239 1031 1240 1035
rect 1234 1030 1240 1031
rect 1270 1034 1276 1035
rect 1270 1030 1271 1034
rect 1275 1030 1276 1034
rect 1222 1029 1228 1030
rect 1270 1029 1276 1030
rect 1326 1034 1332 1035
rect 1326 1030 1327 1034
rect 1331 1030 1332 1034
rect 1338 1031 1339 1035
rect 1343 1031 1344 1035
rect 1338 1030 1344 1031
rect 1382 1034 1388 1035
rect 1382 1030 1383 1034
rect 1387 1030 1388 1034
rect 1326 1029 1332 1030
rect 1382 1029 1388 1030
rect 1224 1027 1226 1029
rect 1272 1027 1274 1029
rect 1328 1027 1330 1029
rect 1384 1027 1386 1029
rect 1031 1026 1035 1027
rect 1031 1021 1035 1022
rect 1047 1026 1051 1027
rect 1047 1021 1051 1022
rect 1079 1026 1083 1027
rect 1079 1021 1083 1022
rect 1103 1026 1107 1027
rect 1103 1021 1107 1022
rect 1127 1026 1131 1027
rect 1127 1021 1131 1022
rect 1159 1026 1163 1027
rect 1159 1021 1163 1022
rect 1175 1026 1179 1027
rect 1186 1026 1192 1027
rect 1215 1026 1219 1027
rect 1175 1021 1179 1022
rect 1002 1019 1008 1020
rect 1048 1019 1050 1021
rect 1104 1019 1106 1021
rect 1160 1019 1162 1021
rect 878 1018 884 1019
rect 878 1014 879 1018
rect 883 1014 884 1018
rect 878 1013 884 1014
rect 934 1018 940 1019
rect 934 1014 935 1018
rect 939 1014 940 1018
rect 934 1013 940 1014
rect 990 1018 996 1019
rect 990 1014 991 1018
rect 995 1014 996 1018
rect 1002 1015 1003 1019
rect 1007 1015 1008 1019
rect 1002 1014 1008 1015
rect 1046 1018 1052 1019
rect 1046 1014 1047 1018
rect 1051 1014 1052 1018
rect 990 1013 996 1014
rect 1046 1013 1052 1014
rect 1102 1018 1108 1019
rect 1102 1014 1103 1018
rect 1107 1014 1108 1018
rect 1102 1013 1108 1014
rect 1158 1018 1164 1019
rect 1158 1014 1159 1018
rect 1163 1014 1164 1018
rect 1158 1013 1164 1014
rect 1188 1008 1190 1026
rect 1215 1021 1219 1022
rect 1223 1026 1227 1027
rect 1223 1021 1227 1022
rect 1271 1026 1275 1027
rect 1271 1021 1275 1022
rect 1327 1026 1331 1027
rect 1327 1021 1331 1022
rect 1383 1026 1387 1027
rect 1383 1021 1387 1022
rect 1216 1019 1218 1021
rect 1272 1019 1274 1021
rect 1328 1019 1330 1021
rect 1384 1019 1386 1021
rect 1396 1020 1398 1038
rect 1428 1036 1430 1066
rect 1447 1061 1451 1062
rect 1448 1058 1450 1061
rect 1446 1057 1452 1058
rect 1446 1053 1447 1057
rect 1451 1053 1452 1057
rect 1446 1052 1452 1053
rect 1446 1039 1452 1040
rect 1426 1035 1432 1036
rect 1414 1034 1420 1035
rect 1414 1030 1415 1034
rect 1419 1030 1420 1034
rect 1426 1031 1427 1035
rect 1431 1031 1432 1035
rect 1446 1035 1447 1039
rect 1451 1035 1452 1039
rect 1446 1034 1452 1035
rect 1426 1030 1432 1031
rect 1414 1029 1420 1030
rect 1416 1027 1418 1029
rect 1448 1027 1450 1034
rect 1415 1026 1419 1027
rect 1415 1021 1419 1022
rect 1447 1026 1451 1027
rect 1447 1021 1451 1022
rect 1394 1019 1400 1020
rect 1416 1019 1418 1021
rect 1214 1018 1220 1019
rect 1214 1014 1215 1018
rect 1219 1014 1220 1018
rect 1214 1013 1220 1014
rect 1270 1018 1276 1019
rect 1270 1014 1271 1018
rect 1275 1014 1276 1018
rect 1270 1013 1276 1014
rect 1326 1018 1332 1019
rect 1326 1014 1327 1018
rect 1331 1014 1332 1018
rect 1382 1018 1388 1019
rect 1326 1013 1332 1014
rect 1346 1015 1352 1016
rect 1346 1011 1347 1015
rect 1351 1011 1352 1015
rect 1382 1014 1383 1018
rect 1387 1014 1388 1018
rect 1394 1015 1395 1019
rect 1399 1015 1400 1019
rect 1394 1014 1400 1015
rect 1414 1018 1420 1019
rect 1414 1014 1415 1018
rect 1419 1014 1420 1018
rect 1448 1014 1450 1021
rect 1382 1013 1388 1014
rect 1414 1013 1420 1014
rect 1446 1013 1452 1014
rect 1346 1010 1352 1011
rect 602 1007 608 1008
rect 602 1003 603 1007
rect 607 1003 608 1007
rect 602 1002 608 1003
rect 834 1007 840 1008
rect 834 1003 835 1007
rect 839 1003 840 1007
rect 834 1002 840 1003
rect 898 1007 904 1008
rect 898 1003 899 1007
rect 903 1003 904 1007
rect 898 1002 904 1003
rect 1186 1007 1192 1008
rect 1186 1003 1187 1007
rect 1191 1003 1192 1007
rect 1186 1002 1192 1003
rect 538 995 544 996
rect 430 992 436 993
rect 430 988 431 992
rect 435 988 436 992
rect 430 987 436 988
rect 478 992 484 993
rect 478 988 479 992
rect 483 988 484 992
rect 478 987 484 988
rect 526 992 532 993
rect 526 988 527 992
rect 531 988 532 992
rect 538 991 539 995
rect 543 991 544 995
rect 538 990 544 991
rect 574 992 580 993
rect 526 987 532 988
rect 574 988 575 992
rect 579 988 580 992
rect 574 987 580 988
rect 622 992 628 993
rect 670 992 676 993
rect 622 988 623 992
rect 627 988 628 992
rect 622 987 628 988
rect 662 991 668 992
rect 662 987 663 991
rect 667 987 668 991
rect 670 988 671 992
rect 675 988 676 992
rect 670 987 676 988
rect 718 992 724 993
rect 718 988 719 992
rect 723 988 724 992
rect 718 987 724 988
rect 766 992 772 993
rect 766 988 767 992
rect 771 988 772 992
rect 766 987 772 988
rect 822 992 828 993
rect 822 988 823 992
rect 827 988 828 992
rect 822 987 828 988
rect 878 992 884 993
rect 878 988 879 992
rect 883 988 884 992
rect 878 987 884 988
rect 423 986 427 987
rect 423 981 427 982
rect 431 986 435 987
rect 431 981 435 982
rect 471 986 475 987
rect 471 981 475 982
rect 479 986 483 987
rect 479 981 483 982
rect 519 986 523 987
rect 519 981 523 982
rect 527 986 531 987
rect 527 981 531 982
rect 567 986 571 987
rect 567 981 571 982
rect 575 986 579 987
rect 575 981 579 982
rect 623 986 627 987
rect 662 986 668 987
rect 671 986 675 987
rect 623 981 627 982
rect 422 980 428 981
rect 422 976 423 980
rect 427 976 428 980
rect 422 975 428 976
rect 470 980 476 981
rect 470 976 471 980
rect 475 976 476 980
rect 470 975 476 976
rect 518 980 524 981
rect 518 976 519 980
rect 523 976 524 980
rect 518 975 524 976
rect 566 980 572 981
rect 566 976 567 980
rect 571 976 572 980
rect 566 975 572 976
rect 622 980 628 981
rect 622 976 623 980
rect 627 976 628 980
rect 622 975 628 976
rect 242 971 248 972
rect 242 967 243 971
rect 247 967 248 971
rect 242 966 248 967
rect 266 971 272 972
rect 266 967 267 971
rect 271 967 272 971
rect 266 966 272 967
rect 338 971 344 972
rect 338 967 339 971
rect 343 967 344 971
rect 338 966 344 967
rect 410 971 416 972
rect 410 967 411 971
rect 415 967 416 971
rect 410 966 416 967
rect 244 956 246 966
rect 268 956 270 966
rect 340 956 342 966
rect 218 955 224 956
rect 242 955 248 956
rect 266 955 272 956
rect 338 955 344 956
rect 110 954 116 955
rect 206 954 212 955
rect 112 947 114 954
rect 206 950 207 954
rect 211 950 212 954
rect 218 951 219 955
rect 223 951 224 955
rect 218 950 224 951
rect 230 954 236 955
rect 230 950 231 954
rect 235 950 236 954
rect 242 951 243 955
rect 247 951 248 955
rect 242 950 248 951
rect 254 954 260 955
rect 254 950 255 954
rect 259 950 260 954
rect 266 951 267 955
rect 271 951 272 955
rect 266 950 272 951
rect 286 954 292 955
rect 286 950 287 954
rect 291 950 292 954
rect 206 949 212 950
rect 230 949 236 950
rect 254 949 260 950
rect 286 949 292 950
rect 326 954 332 955
rect 326 950 327 954
rect 331 950 332 954
rect 338 951 339 955
rect 343 951 344 955
rect 338 950 344 951
rect 374 954 380 955
rect 374 950 375 954
rect 379 950 380 954
rect 326 949 332 950
rect 374 949 380 950
rect 422 954 428 955
rect 422 950 423 954
rect 427 950 428 954
rect 422 949 428 950
rect 470 954 476 955
rect 470 950 471 954
rect 475 950 476 954
rect 470 949 476 950
rect 518 954 524 955
rect 518 950 519 954
rect 523 950 524 954
rect 566 954 572 955
rect 518 949 524 950
rect 530 951 536 952
rect 208 947 210 949
rect 232 947 234 949
rect 256 947 258 949
rect 274 947 280 948
rect 288 947 290 949
rect 302 947 308 948
rect 328 947 330 949
rect 376 947 378 949
rect 424 947 426 949
rect 472 947 474 949
rect 520 947 522 949
rect 530 947 531 951
rect 535 947 536 951
rect 566 950 567 954
rect 571 950 572 954
rect 566 949 572 950
rect 622 954 628 955
rect 622 950 623 954
rect 627 950 628 954
rect 622 949 628 950
rect 568 947 570 949
rect 624 947 626 949
rect 664 948 666 986
rect 671 981 675 982
rect 679 986 683 987
rect 679 981 683 982
rect 719 986 723 987
rect 719 981 723 982
rect 727 986 731 987
rect 727 981 731 982
rect 767 986 771 987
rect 767 981 771 982
rect 775 986 779 987
rect 775 981 779 982
rect 823 986 827 987
rect 823 981 827 982
rect 831 986 835 987
rect 831 981 835 982
rect 879 986 883 987
rect 879 981 883 982
rect 887 986 891 987
rect 887 981 891 982
rect 678 980 684 981
rect 678 976 679 980
rect 683 976 684 980
rect 678 975 684 976
rect 726 980 732 981
rect 726 976 727 980
rect 731 976 732 980
rect 726 975 732 976
rect 774 980 780 981
rect 774 976 775 980
rect 779 976 780 980
rect 774 975 780 976
rect 830 980 836 981
rect 830 976 831 980
rect 835 976 836 980
rect 830 975 836 976
rect 886 980 892 981
rect 900 980 902 1002
rect 934 992 940 993
rect 934 988 935 992
rect 939 988 940 992
rect 934 987 940 988
rect 990 992 996 993
rect 990 988 991 992
rect 995 988 996 992
rect 990 987 996 988
rect 1046 992 1052 993
rect 1046 988 1047 992
rect 1051 988 1052 992
rect 1046 987 1052 988
rect 1102 992 1108 993
rect 1158 992 1164 993
rect 1102 988 1103 992
rect 1107 988 1108 992
rect 1102 987 1108 988
rect 1114 991 1120 992
rect 1114 987 1115 991
rect 1119 987 1120 991
rect 1158 988 1159 992
rect 1163 988 1164 992
rect 1158 987 1164 988
rect 1214 992 1220 993
rect 1214 988 1215 992
rect 1219 988 1220 992
rect 1214 987 1220 988
rect 1270 992 1276 993
rect 1270 988 1271 992
rect 1275 988 1276 992
rect 1270 987 1276 988
rect 1326 992 1332 993
rect 1326 988 1327 992
rect 1331 988 1332 992
rect 1326 987 1332 988
rect 935 986 939 987
rect 935 981 939 982
rect 943 986 947 987
rect 943 981 947 982
rect 991 986 995 987
rect 991 981 995 982
rect 999 986 1003 987
rect 999 981 1003 982
rect 1047 986 1051 987
rect 1047 981 1051 982
rect 1095 986 1099 987
rect 1095 981 1099 982
rect 1103 986 1107 987
rect 1114 986 1120 987
rect 1143 986 1147 987
rect 1103 981 1107 982
rect 942 980 948 981
rect 886 976 887 980
rect 891 976 892 980
rect 886 975 892 976
rect 898 979 904 980
rect 898 975 899 979
rect 903 975 904 979
rect 942 976 943 980
rect 947 976 948 980
rect 942 975 948 976
rect 998 980 1004 981
rect 998 976 999 980
rect 1003 976 1004 980
rect 998 975 1004 976
rect 1046 980 1052 981
rect 1046 976 1047 980
rect 1051 976 1052 980
rect 1046 975 1052 976
rect 1094 980 1100 981
rect 1094 976 1095 980
rect 1099 976 1100 980
rect 1094 975 1100 976
rect 898 974 904 975
rect 738 971 744 972
rect 738 967 739 971
rect 743 967 744 971
rect 738 966 744 967
rect 842 971 848 972
rect 842 967 843 971
rect 847 967 848 971
rect 842 966 848 967
rect 678 954 684 955
rect 678 950 679 954
rect 683 950 684 954
rect 678 949 684 950
rect 726 954 732 955
rect 726 950 727 954
rect 731 950 732 954
rect 726 949 732 950
rect 662 947 668 948
rect 680 947 682 949
rect 728 947 730 949
rect 111 946 115 947
rect 111 941 115 942
rect 207 946 211 947
rect 207 941 211 942
rect 215 946 219 947
rect 215 941 219 942
rect 231 946 235 947
rect 231 941 235 942
rect 239 946 243 947
rect 239 941 243 942
rect 255 946 259 947
rect 255 941 259 942
rect 263 946 267 947
rect 274 943 275 947
rect 279 943 280 947
rect 274 942 280 943
rect 287 946 291 947
rect 302 943 303 947
rect 307 943 308 947
rect 302 942 308 943
rect 319 946 323 947
rect 263 941 267 942
rect 112 934 114 941
rect 216 939 218 941
rect 240 939 242 941
rect 264 939 266 941
rect 214 938 220 939
rect 214 934 215 938
rect 219 934 220 938
rect 238 938 244 939
rect 110 933 116 934
rect 214 933 220 934
rect 226 935 232 936
rect 110 929 111 933
rect 115 929 116 933
rect 226 930 227 935
rect 110 928 116 929
rect 231 930 232 935
rect 238 934 239 938
rect 243 934 244 938
rect 238 933 244 934
rect 262 938 268 939
rect 262 934 263 938
rect 267 934 268 938
rect 262 933 268 934
rect 227 927 231 928
rect 276 916 278 942
rect 287 941 291 942
rect 288 939 290 941
rect 286 938 292 939
rect 286 934 287 938
rect 291 934 292 938
rect 286 933 292 934
rect 304 933 306 942
rect 319 941 323 942
rect 327 946 331 947
rect 327 941 331 942
rect 351 946 355 947
rect 351 941 355 942
rect 375 946 379 947
rect 375 941 379 942
rect 391 946 395 947
rect 391 941 395 942
rect 423 946 427 947
rect 423 941 427 942
rect 431 946 435 947
rect 431 941 435 942
rect 471 946 475 947
rect 471 941 475 942
rect 519 946 523 947
rect 530 946 536 947
rect 567 946 571 947
rect 519 941 523 942
rect 320 939 322 941
rect 352 939 354 941
rect 392 939 394 941
rect 432 939 434 941
rect 472 939 474 941
rect 520 939 522 941
rect 318 938 324 939
rect 318 934 319 938
rect 323 934 324 938
rect 318 933 324 934
rect 350 938 356 939
rect 350 934 351 938
rect 355 934 356 938
rect 350 933 356 934
rect 390 938 396 939
rect 390 934 391 938
rect 395 934 396 938
rect 390 933 396 934
rect 430 938 436 939
rect 430 934 431 938
rect 435 934 436 938
rect 430 933 436 934
rect 470 938 476 939
rect 470 934 471 938
rect 475 934 476 938
rect 518 938 524 939
rect 470 933 476 934
rect 506 935 512 936
rect 303 932 307 933
rect 443 932 447 933
rect 506 931 507 935
rect 511 931 512 935
rect 518 934 519 938
rect 523 934 524 938
rect 518 933 524 934
rect 506 930 512 931
rect 303 927 307 928
rect 442 927 448 928
rect 442 923 443 927
rect 447 923 448 927
rect 442 922 448 923
rect 110 915 116 916
rect 110 911 111 915
rect 115 911 116 915
rect 274 915 280 916
rect 110 910 116 911
rect 214 912 220 913
rect 112 907 114 910
rect 214 908 215 912
rect 219 908 220 912
rect 214 907 220 908
rect 238 912 244 913
rect 238 908 239 912
rect 243 908 244 912
rect 238 907 244 908
rect 262 912 268 913
rect 262 908 263 912
rect 267 908 268 912
rect 274 911 275 915
rect 279 911 280 915
rect 274 910 280 911
rect 286 912 292 913
rect 262 907 268 908
rect 286 908 287 912
rect 291 908 292 912
rect 286 907 292 908
rect 318 912 324 913
rect 318 908 319 912
rect 323 908 324 912
rect 318 907 324 908
rect 350 912 356 913
rect 350 908 351 912
rect 355 908 356 912
rect 350 907 356 908
rect 390 912 396 913
rect 430 912 436 913
rect 390 908 391 912
rect 395 908 396 912
rect 390 907 396 908
rect 402 911 408 912
rect 402 907 403 911
rect 407 907 408 911
rect 430 908 431 912
rect 435 908 436 912
rect 430 907 436 908
rect 470 912 476 913
rect 470 908 471 912
rect 475 908 476 912
rect 470 907 476 908
rect 111 906 115 907
rect 111 901 115 902
rect 215 906 219 907
rect 215 901 219 902
rect 231 906 235 907
rect 231 901 235 902
rect 239 906 243 907
rect 239 901 243 902
rect 255 906 259 907
rect 255 901 259 902
rect 263 906 267 907
rect 263 901 267 902
rect 279 906 283 907
rect 279 901 283 902
rect 287 906 291 907
rect 287 901 291 902
rect 303 906 307 907
rect 303 901 307 902
rect 319 906 323 907
rect 319 901 323 902
rect 327 906 331 907
rect 327 901 331 902
rect 351 906 355 907
rect 351 901 355 902
rect 359 906 363 907
rect 359 901 363 902
rect 391 906 395 907
rect 402 906 408 907
rect 423 906 427 907
rect 391 901 395 902
rect 112 898 114 901
rect 230 900 236 901
rect 110 897 116 898
rect 110 893 111 897
rect 115 893 116 897
rect 230 896 231 900
rect 235 896 236 900
rect 230 895 236 896
rect 254 900 260 901
rect 254 896 255 900
rect 259 896 260 900
rect 254 895 260 896
rect 278 900 284 901
rect 278 896 279 900
rect 283 896 284 900
rect 278 895 284 896
rect 302 900 308 901
rect 302 896 303 900
rect 307 896 308 900
rect 302 895 308 896
rect 326 900 332 901
rect 326 896 327 900
rect 331 896 332 900
rect 326 895 332 896
rect 358 900 364 901
rect 358 896 359 900
rect 363 896 364 900
rect 358 895 364 896
rect 390 900 396 901
rect 390 896 391 900
rect 395 896 396 900
rect 390 895 396 896
rect 110 892 116 893
rect 238 887 244 888
rect 238 883 239 887
rect 243 883 244 887
rect 238 882 244 883
rect 110 879 116 880
rect 110 875 111 879
rect 115 875 116 879
rect 110 874 116 875
rect 230 874 236 875
rect 112 867 114 874
rect 230 870 231 874
rect 235 870 236 874
rect 230 869 236 870
rect 232 867 234 869
rect 240 868 242 882
rect 404 876 406 906
rect 423 901 427 902
rect 431 906 435 907
rect 431 901 435 902
rect 455 906 459 907
rect 455 901 459 902
rect 471 906 475 907
rect 471 901 475 902
rect 495 906 499 907
rect 495 901 499 902
rect 422 900 428 901
rect 422 896 423 900
rect 427 896 428 900
rect 422 895 428 896
rect 454 900 460 901
rect 454 896 455 900
rect 459 896 460 900
rect 454 895 460 896
rect 494 900 500 901
rect 508 900 510 930
rect 532 928 534 946
rect 567 941 571 942
rect 615 946 619 947
rect 615 941 619 942
rect 623 946 627 947
rect 662 943 663 947
rect 667 943 668 947
rect 662 942 668 943
rect 671 946 675 947
rect 623 941 627 942
rect 671 941 675 942
rect 679 946 683 947
rect 679 941 683 942
rect 727 946 731 947
rect 727 941 731 942
rect 568 939 570 941
rect 616 939 618 941
rect 672 939 674 941
rect 728 939 730 941
rect 740 940 742 966
rect 844 956 846 966
rect 930 963 936 964
rect 930 959 931 963
rect 935 959 936 963
rect 930 958 936 959
rect 842 955 848 956
rect 774 954 780 955
rect 774 950 775 954
rect 779 950 780 954
rect 830 954 836 955
rect 774 949 780 950
rect 794 951 800 952
rect 776 947 778 949
rect 794 947 795 951
rect 799 947 800 951
rect 830 950 831 954
rect 835 950 836 954
rect 842 951 843 955
rect 847 951 848 955
rect 842 950 848 951
rect 886 954 892 955
rect 886 950 887 954
rect 891 950 892 954
rect 830 949 836 950
rect 886 949 892 950
rect 832 947 834 949
rect 888 947 890 949
rect 775 946 779 947
rect 775 941 779 942
rect 783 946 787 947
rect 794 946 800 947
rect 831 946 835 947
rect 783 941 787 942
rect 738 939 744 940
rect 784 939 786 941
rect 566 938 572 939
rect 538 935 544 936
rect 538 930 539 935
rect 543 930 544 935
rect 566 934 567 938
rect 571 934 572 938
rect 566 933 572 934
rect 614 938 620 939
rect 614 934 615 938
rect 619 934 620 938
rect 614 933 620 934
rect 670 938 676 939
rect 670 934 671 938
rect 675 934 676 938
rect 670 933 676 934
rect 726 938 732 939
rect 726 934 727 938
rect 731 934 732 938
rect 738 935 739 939
rect 743 935 744 939
rect 738 934 744 935
rect 782 938 788 939
rect 782 934 783 938
rect 787 934 788 938
rect 726 933 732 934
rect 782 933 788 934
rect 796 928 798 946
rect 831 941 835 942
rect 847 946 851 947
rect 847 941 851 942
rect 887 946 891 947
rect 887 941 891 942
rect 919 946 923 947
rect 919 941 923 942
rect 848 939 850 941
rect 920 939 922 941
rect 932 940 934 958
rect 1116 956 1118 986
rect 1143 981 1147 982
rect 1159 986 1163 987
rect 1159 981 1163 982
rect 1191 986 1195 987
rect 1191 981 1195 982
rect 1215 986 1219 987
rect 1215 981 1219 982
rect 1239 986 1243 987
rect 1239 981 1243 982
rect 1271 986 1275 987
rect 1271 981 1275 982
rect 1287 986 1291 987
rect 1287 981 1291 982
rect 1327 986 1331 987
rect 1327 981 1331 982
rect 1335 986 1339 987
rect 1335 981 1339 982
rect 1142 980 1148 981
rect 1142 976 1143 980
rect 1147 976 1148 980
rect 1142 975 1148 976
rect 1190 980 1196 981
rect 1190 976 1191 980
rect 1195 976 1196 980
rect 1190 975 1196 976
rect 1238 980 1244 981
rect 1238 976 1239 980
rect 1243 976 1244 980
rect 1238 975 1244 976
rect 1286 980 1292 981
rect 1286 976 1287 980
rect 1291 976 1292 980
rect 1286 975 1292 976
rect 1334 980 1340 981
rect 1334 976 1335 980
rect 1339 976 1340 980
rect 1334 975 1340 976
rect 1348 972 1350 1010
rect 1446 1009 1447 1013
rect 1451 1009 1452 1013
rect 1446 1008 1452 1009
rect 1446 995 1452 996
rect 1382 992 1388 993
rect 1382 988 1383 992
rect 1387 988 1388 992
rect 1382 987 1388 988
rect 1414 992 1420 993
rect 1414 988 1415 992
rect 1419 988 1420 992
rect 1414 987 1420 988
rect 1426 991 1432 992
rect 1426 987 1427 991
rect 1431 987 1432 991
rect 1446 991 1447 995
rect 1451 991 1452 995
rect 1446 990 1452 991
rect 1448 987 1450 990
rect 1383 986 1387 987
rect 1383 981 1387 982
rect 1415 986 1419 987
rect 1426 986 1432 987
rect 1447 986 1451 987
rect 1415 981 1419 982
rect 1382 980 1388 981
rect 1382 976 1383 980
rect 1387 976 1388 980
rect 1382 975 1388 976
rect 1414 980 1420 981
rect 1414 976 1415 980
rect 1419 976 1420 980
rect 1414 975 1420 976
rect 1346 971 1352 972
rect 1346 967 1347 971
rect 1351 967 1352 971
rect 1346 966 1352 967
rect 1428 956 1430 986
rect 1447 981 1451 982
rect 1448 978 1450 981
rect 1446 977 1452 978
rect 1446 973 1447 977
rect 1451 973 1452 977
rect 1446 972 1452 973
rect 1446 959 1452 960
rect 1114 955 1120 956
rect 1426 955 1432 956
rect 942 954 948 955
rect 942 950 943 954
rect 947 950 948 954
rect 942 949 948 950
rect 998 954 1004 955
rect 998 950 999 954
rect 1003 950 1004 954
rect 998 949 1004 950
rect 1046 954 1052 955
rect 1046 950 1047 954
rect 1051 950 1052 954
rect 1046 949 1052 950
rect 1094 954 1100 955
rect 1094 950 1095 954
rect 1099 950 1100 954
rect 1114 951 1115 955
rect 1119 951 1120 955
rect 1114 950 1120 951
rect 1142 954 1148 955
rect 1142 950 1143 954
rect 1147 950 1148 954
rect 1094 949 1100 950
rect 1142 949 1148 950
rect 1190 954 1196 955
rect 1190 950 1191 954
rect 1195 950 1196 954
rect 1190 949 1196 950
rect 1238 954 1244 955
rect 1238 950 1239 954
rect 1243 950 1244 954
rect 1238 949 1244 950
rect 1286 954 1292 955
rect 1286 950 1287 954
rect 1291 950 1292 954
rect 1286 949 1292 950
rect 1334 954 1340 955
rect 1334 950 1335 954
rect 1339 950 1340 954
rect 1334 949 1340 950
rect 1382 954 1388 955
rect 1382 950 1383 954
rect 1387 950 1388 954
rect 1382 949 1388 950
rect 1414 954 1420 955
rect 1414 950 1415 954
rect 1419 950 1420 954
rect 1426 951 1427 955
rect 1431 951 1432 955
rect 1446 955 1447 959
rect 1451 955 1452 959
rect 1446 954 1452 955
rect 1426 950 1432 951
rect 1414 949 1420 950
rect 944 947 946 949
rect 1000 947 1002 949
rect 1048 947 1050 949
rect 1096 947 1098 949
rect 1130 947 1136 948
rect 1144 947 1146 949
rect 1192 947 1194 949
rect 1240 947 1242 949
rect 1288 947 1290 949
rect 1336 947 1338 949
rect 1384 947 1386 949
rect 1416 947 1418 949
rect 1448 947 1450 954
rect 943 946 947 947
rect 943 941 947 942
rect 991 946 995 947
rect 991 941 995 942
rect 999 946 1003 947
rect 999 941 1003 942
rect 1047 946 1051 947
rect 1047 941 1051 942
rect 1055 946 1059 947
rect 1055 941 1059 942
rect 1095 946 1099 947
rect 1095 941 1099 942
rect 1119 946 1123 947
rect 1130 943 1131 947
rect 1135 943 1136 947
rect 1130 942 1136 943
rect 1143 946 1147 947
rect 1119 941 1123 942
rect 930 939 936 940
rect 992 939 994 941
rect 1056 939 1058 941
rect 1120 939 1122 941
rect 846 938 852 939
rect 846 934 847 938
rect 851 934 852 938
rect 918 938 924 939
rect 846 933 852 934
rect 858 935 864 936
rect 858 931 859 935
rect 863 931 864 935
rect 918 934 919 938
rect 923 934 924 938
rect 930 935 931 939
rect 935 935 936 939
rect 930 934 936 935
rect 990 938 996 939
rect 990 934 991 938
rect 995 934 996 938
rect 1054 938 1060 939
rect 918 933 924 934
rect 990 933 996 934
rect 1002 935 1008 936
rect 858 930 864 931
rect 1002 931 1003 935
rect 1007 931 1008 935
rect 1054 934 1055 938
rect 1059 934 1060 938
rect 1054 933 1060 934
rect 1118 938 1124 939
rect 1118 934 1119 938
rect 1123 934 1124 938
rect 1118 933 1124 934
rect 1002 930 1008 931
rect 530 927 536 928
rect 539 927 543 928
rect 794 927 800 928
rect 530 923 531 927
rect 535 923 536 927
rect 530 922 536 923
rect 794 923 795 927
rect 799 923 800 927
rect 794 922 800 923
rect 860 915 862 930
rect 990 923 996 924
rect 1004 923 1006 930
rect 1132 928 1134 942
rect 1143 941 1147 942
rect 1175 946 1179 947
rect 1175 941 1179 942
rect 1191 946 1195 947
rect 1191 941 1195 942
rect 1223 946 1227 947
rect 1223 941 1227 942
rect 1239 946 1243 947
rect 1239 941 1243 942
rect 1263 946 1267 947
rect 1263 941 1267 942
rect 1287 946 1291 947
rect 1287 941 1291 942
rect 1295 946 1299 947
rect 1295 941 1299 942
rect 1327 946 1331 947
rect 1327 941 1331 942
rect 1335 946 1339 947
rect 1335 941 1339 942
rect 1359 946 1363 947
rect 1359 941 1363 942
rect 1383 946 1387 947
rect 1383 941 1387 942
rect 1391 946 1395 947
rect 1391 941 1395 942
rect 1415 946 1419 947
rect 1415 941 1419 942
rect 1447 946 1451 947
rect 1447 941 1451 942
rect 1176 939 1178 941
rect 1224 939 1226 941
rect 1264 939 1266 941
rect 1296 939 1298 941
rect 1328 939 1330 941
rect 1360 939 1362 941
rect 1392 939 1394 941
rect 1416 939 1418 941
rect 1174 938 1180 939
rect 1174 934 1175 938
rect 1179 934 1180 938
rect 1174 933 1180 934
rect 1222 938 1228 939
rect 1222 934 1223 938
rect 1227 934 1228 938
rect 1222 933 1228 934
rect 1262 938 1268 939
rect 1262 934 1263 938
rect 1267 934 1268 938
rect 1262 933 1268 934
rect 1294 938 1300 939
rect 1294 934 1295 938
rect 1299 934 1300 938
rect 1294 933 1300 934
rect 1326 938 1332 939
rect 1326 934 1327 938
rect 1331 934 1332 938
rect 1326 933 1332 934
rect 1358 938 1364 939
rect 1358 934 1359 938
rect 1363 934 1364 938
rect 1358 933 1364 934
rect 1390 938 1396 939
rect 1390 934 1391 938
rect 1395 934 1396 938
rect 1390 933 1396 934
rect 1414 938 1420 939
rect 1414 934 1415 938
rect 1419 934 1420 938
rect 1448 934 1450 941
rect 1414 933 1420 934
rect 1446 933 1452 934
rect 1446 929 1447 933
rect 1451 929 1452 933
rect 1446 928 1452 929
rect 990 919 991 923
rect 995 921 1006 923
rect 1130 927 1136 928
rect 1130 923 1131 927
rect 1135 923 1136 927
rect 1130 922 1136 923
rect 995 919 996 921
rect 990 918 996 919
rect 856 913 862 915
rect 1446 915 1452 916
rect 518 912 524 913
rect 518 908 519 912
rect 523 908 524 912
rect 518 907 524 908
rect 566 912 572 913
rect 614 912 620 913
rect 566 908 567 912
rect 571 908 572 912
rect 566 907 572 908
rect 606 911 612 912
rect 606 907 607 911
rect 611 907 612 911
rect 614 908 615 912
rect 619 908 620 912
rect 614 907 620 908
rect 670 912 676 913
rect 670 908 671 912
rect 675 908 676 912
rect 670 907 676 908
rect 726 912 732 913
rect 726 908 727 912
rect 731 908 732 912
rect 726 907 732 908
rect 782 912 788 913
rect 782 908 783 912
rect 787 908 788 912
rect 782 907 788 908
rect 846 912 852 913
rect 846 908 847 912
rect 851 908 852 912
rect 846 907 852 908
rect 519 906 523 907
rect 519 901 523 902
rect 535 906 539 907
rect 535 901 539 902
rect 567 906 571 907
rect 567 901 571 902
rect 575 906 579 907
rect 606 906 612 907
rect 615 906 619 907
rect 575 901 579 902
rect 534 900 540 901
rect 494 896 495 900
rect 499 896 500 900
rect 494 895 500 896
rect 506 899 512 900
rect 506 895 507 899
rect 511 895 512 899
rect 534 896 535 900
rect 539 896 540 900
rect 534 895 540 896
rect 574 900 580 901
rect 574 896 575 900
rect 579 896 580 900
rect 574 895 580 896
rect 506 894 512 895
rect 466 891 472 892
rect 466 887 467 891
rect 471 887 472 891
rect 466 886 472 887
rect 468 876 470 886
rect 402 875 408 876
rect 466 875 472 876
rect 254 874 260 875
rect 254 870 255 874
rect 259 870 260 874
rect 254 869 260 870
rect 278 874 284 875
rect 278 870 279 874
rect 283 870 284 874
rect 278 869 284 870
rect 302 874 308 875
rect 302 870 303 874
rect 307 870 308 874
rect 302 869 308 870
rect 326 874 332 875
rect 326 870 327 874
rect 331 870 332 874
rect 326 869 332 870
rect 358 874 364 875
rect 358 870 359 874
rect 363 870 364 874
rect 358 869 364 870
rect 390 874 396 875
rect 390 870 391 874
rect 395 870 396 874
rect 402 871 403 875
rect 407 871 408 875
rect 402 870 408 871
rect 422 874 428 875
rect 422 870 423 874
rect 427 870 428 874
rect 390 869 396 870
rect 422 869 428 870
rect 454 874 460 875
rect 454 870 455 874
rect 459 870 460 874
rect 466 871 467 875
rect 471 871 472 875
rect 466 870 472 871
rect 494 874 500 875
rect 494 870 495 874
rect 499 870 500 874
rect 454 869 460 870
rect 494 869 500 870
rect 534 874 540 875
rect 534 870 535 874
rect 539 870 540 874
rect 534 869 540 870
rect 574 874 580 875
rect 574 870 575 874
rect 579 870 580 874
rect 574 869 580 870
rect 238 867 244 868
rect 256 867 258 869
rect 280 867 282 869
rect 304 867 306 869
rect 328 867 330 869
rect 360 867 362 869
rect 392 867 394 869
rect 398 867 404 868
rect 424 867 426 869
rect 456 867 458 869
rect 496 867 498 869
rect 536 867 538 869
rect 576 867 578 869
rect 608 868 610 906
rect 615 901 619 902
rect 623 906 627 907
rect 623 901 627 902
rect 663 906 667 907
rect 663 901 667 902
rect 671 906 675 907
rect 671 901 675 902
rect 703 906 707 907
rect 703 901 707 902
rect 727 906 731 907
rect 727 901 731 902
rect 751 906 755 907
rect 751 901 755 902
rect 783 906 787 907
rect 783 901 787 902
rect 807 906 811 907
rect 807 901 811 902
rect 847 906 851 907
rect 847 901 851 902
rect 622 900 628 901
rect 622 896 623 900
rect 627 896 628 900
rect 622 895 628 896
rect 662 900 668 901
rect 662 896 663 900
rect 667 896 668 900
rect 662 895 668 896
rect 702 900 708 901
rect 702 896 703 900
rect 707 896 708 900
rect 702 895 708 896
rect 750 900 756 901
rect 750 896 751 900
rect 755 896 756 900
rect 750 895 756 896
rect 806 900 812 901
rect 856 900 858 913
rect 918 912 924 913
rect 918 908 919 912
rect 923 908 924 912
rect 918 907 924 908
rect 990 912 996 913
rect 990 908 991 912
rect 995 908 996 912
rect 990 907 996 908
rect 1054 912 1060 913
rect 1118 912 1124 913
rect 1054 908 1055 912
rect 1059 908 1060 912
rect 1054 907 1060 908
rect 1066 911 1072 912
rect 1066 907 1067 911
rect 1071 907 1072 911
rect 1118 908 1119 912
rect 1123 908 1124 912
rect 1118 907 1124 908
rect 1174 912 1180 913
rect 1174 908 1175 912
rect 1179 908 1180 912
rect 1174 907 1180 908
rect 1222 912 1228 913
rect 1222 908 1223 912
rect 1227 908 1228 912
rect 1222 907 1228 908
rect 1262 912 1268 913
rect 1262 908 1263 912
rect 1267 908 1268 912
rect 1262 907 1268 908
rect 1294 912 1300 913
rect 1294 908 1295 912
rect 1299 908 1300 912
rect 1294 907 1300 908
rect 1326 912 1332 913
rect 1326 908 1327 912
rect 1331 908 1332 912
rect 1326 907 1332 908
rect 1358 912 1364 913
rect 1358 908 1359 912
rect 1363 908 1364 912
rect 1358 907 1364 908
rect 1390 912 1396 913
rect 1414 912 1420 913
rect 1390 908 1391 912
rect 1395 908 1396 912
rect 1390 907 1396 908
rect 1402 911 1408 912
rect 1402 907 1403 911
rect 1407 907 1408 911
rect 1414 908 1415 912
rect 1419 908 1420 912
rect 1446 911 1447 915
rect 1451 911 1452 915
rect 1446 910 1452 911
rect 1414 907 1420 908
rect 1448 907 1450 910
rect 863 906 867 907
rect 863 901 867 902
rect 919 906 923 907
rect 919 901 923 902
rect 927 906 931 907
rect 927 901 931 902
rect 991 906 995 907
rect 991 901 995 902
rect 1055 906 1059 907
rect 1066 906 1072 907
rect 1119 906 1123 907
rect 1055 901 1059 902
rect 862 900 868 901
rect 806 896 807 900
rect 811 896 812 900
rect 806 895 812 896
rect 854 899 860 900
rect 854 895 855 899
rect 859 895 860 899
rect 862 896 863 900
rect 867 896 868 900
rect 862 895 868 896
rect 926 900 932 901
rect 926 896 927 900
rect 931 896 932 900
rect 926 895 932 896
rect 990 900 996 901
rect 990 896 991 900
rect 995 896 996 900
rect 990 895 996 896
rect 1054 900 1060 901
rect 1054 896 1055 900
rect 1059 896 1060 900
rect 1054 895 1060 896
rect 854 894 860 895
rect 762 891 768 892
rect 762 887 763 891
rect 767 887 768 891
rect 762 886 768 887
rect 764 876 766 886
rect 1068 876 1070 906
rect 1119 901 1123 902
rect 1175 906 1179 907
rect 1175 901 1179 902
rect 1223 906 1227 907
rect 1223 901 1227 902
rect 1231 906 1235 907
rect 1231 901 1235 902
rect 1263 906 1267 907
rect 1263 901 1267 902
rect 1279 906 1283 907
rect 1279 901 1283 902
rect 1295 906 1299 907
rect 1295 901 1299 902
rect 1327 906 1331 907
rect 1327 901 1331 902
rect 1359 906 1363 907
rect 1359 901 1363 902
rect 1383 906 1387 907
rect 1383 901 1387 902
rect 1391 906 1395 907
rect 1402 906 1408 907
rect 1415 906 1419 907
rect 1391 901 1395 902
rect 1118 900 1124 901
rect 1118 896 1119 900
rect 1123 896 1124 900
rect 1118 895 1124 896
rect 1174 900 1180 901
rect 1174 896 1175 900
rect 1179 896 1180 900
rect 1174 895 1180 896
rect 1230 900 1236 901
rect 1230 896 1231 900
rect 1235 896 1236 900
rect 1230 895 1236 896
rect 1278 900 1284 901
rect 1278 896 1279 900
rect 1283 896 1284 900
rect 1278 895 1284 896
rect 1326 900 1332 901
rect 1326 896 1327 900
rect 1331 896 1332 900
rect 1326 895 1332 896
rect 1382 900 1388 901
rect 1382 896 1383 900
rect 1387 896 1388 900
rect 1382 895 1388 896
rect 1186 891 1192 892
rect 1186 887 1187 891
rect 1191 887 1192 891
rect 1186 886 1192 887
rect 1290 891 1296 892
rect 1290 887 1291 891
rect 1295 887 1296 891
rect 1290 886 1296 887
rect 1188 876 1190 886
rect 1292 876 1294 886
rect 762 875 768 876
rect 1066 875 1072 876
rect 1186 875 1192 876
rect 622 874 628 875
rect 622 870 623 874
rect 627 870 628 874
rect 622 869 628 870
rect 662 874 668 875
rect 662 870 663 874
rect 667 870 668 874
rect 662 869 668 870
rect 702 874 708 875
rect 702 870 703 874
rect 707 870 708 874
rect 702 869 708 870
rect 750 874 756 875
rect 750 870 751 874
rect 755 870 756 874
rect 762 871 763 875
rect 767 871 768 875
rect 762 870 768 871
rect 806 874 812 875
rect 806 870 807 874
rect 811 870 812 874
rect 750 869 756 870
rect 806 869 812 870
rect 862 874 868 875
rect 862 870 863 874
rect 867 870 868 874
rect 862 869 868 870
rect 926 874 932 875
rect 926 870 927 874
rect 931 870 932 874
rect 926 869 932 870
rect 990 874 996 875
rect 990 870 991 874
rect 995 870 996 874
rect 990 869 996 870
rect 1054 874 1060 875
rect 1054 870 1055 874
rect 1059 870 1060 874
rect 1066 871 1067 875
rect 1071 871 1072 875
rect 1066 870 1072 871
rect 1118 874 1124 875
rect 1118 870 1119 874
rect 1123 870 1124 874
rect 1054 869 1060 870
rect 1118 869 1124 870
rect 1174 874 1180 875
rect 1174 870 1175 874
rect 1179 870 1180 874
rect 1186 871 1187 875
rect 1191 871 1192 875
rect 1186 870 1192 871
rect 1198 875 1204 876
rect 1290 875 1296 876
rect 1198 871 1199 875
rect 1203 871 1204 875
rect 1198 870 1204 871
rect 1230 874 1236 875
rect 1230 870 1231 874
rect 1235 870 1236 874
rect 1174 869 1180 870
rect 606 867 612 868
rect 624 867 626 869
rect 664 867 666 869
rect 704 867 706 869
rect 752 867 754 869
rect 778 867 784 868
rect 808 867 810 869
rect 864 867 866 869
rect 928 867 930 869
rect 992 867 994 869
rect 1056 867 1058 869
rect 1120 867 1122 869
rect 1176 867 1178 869
rect 1182 867 1188 868
rect 111 866 115 867
rect 111 861 115 862
rect 207 866 211 867
rect 207 861 211 862
rect 231 866 235 867
rect 238 863 239 867
rect 243 863 244 867
rect 238 862 244 863
rect 255 866 259 867
rect 231 861 235 862
rect 255 861 259 862
rect 279 866 283 867
rect 279 861 283 862
rect 287 866 291 867
rect 287 861 291 862
rect 303 866 307 867
rect 303 861 307 862
rect 319 866 323 867
rect 319 861 323 862
rect 327 866 331 867
rect 327 861 331 862
rect 351 866 355 867
rect 351 861 355 862
rect 359 866 363 867
rect 359 861 363 862
rect 383 866 387 867
rect 383 861 387 862
rect 391 866 395 867
rect 398 863 399 867
rect 403 863 404 867
rect 398 862 404 863
rect 415 866 419 867
rect 391 861 395 862
rect 112 854 114 861
rect 208 859 210 861
rect 232 859 234 861
rect 256 859 258 861
rect 288 859 290 861
rect 320 859 322 861
rect 352 859 354 861
rect 384 859 386 861
rect 206 858 212 859
rect 206 854 207 858
rect 211 854 212 858
rect 110 853 116 854
rect 206 853 212 854
rect 230 858 236 859
rect 230 854 231 858
rect 235 854 236 858
rect 230 853 236 854
rect 254 858 260 859
rect 254 854 255 858
rect 259 854 260 858
rect 254 853 260 854
rect 286 858 292 859
rect 286 854 287 858
rect 291 854 292 858
rect 286 853 292 854
rect 318 858 324 859
rect 318 854 319 858
rect 323 854 324 858
rect 318 853 324 854
rect 350 858 356 859
rect 350 854 351 858
rect 355 854 356 858
rect 350 853 356 854
rect 382 858 388 859
rect 382 854 383 858
rect 387 854 388 858
rect 382 853 388 854
rect 110 849 111 853
rect 115 849 116 853
rect 110 848 116 849
rect 391 847 397 848
rect 391 843 392 847
rect 396 846 397 847
rect 400 846 402 862
rect 415 861 419 862
rect 423 866 427 867
rect 423 861 427 862
rect 447 866 451 867
rect 447 861 451 862
rect 455 866 459 867
rect 455 861 459 862
rect 479 866 483 867
rect 479 861 483 862
rect 495 866 499 867
rect 495 861 499 862
rect 511 866 515 867
rect 511 861 515 862
rect 535 866 539 867
rect 535 861 539 862
rect 551 866 555 867
rect 551 861 555 862
rect 575 866 579 867
rect 575 861 579 862
rect 599 866 603 867
rect 606 863 607 867
rect 611 863 612 867
rect 606 862 612 863
rect 623 866 627 867
rect 599 861 603 862
rect 623 861 627 862
rect 647 866 651 867
rect 647 861 651 862
rect 663 866 667 867
rect 663 861 667 862
rect 703 866 707 867
rect 703 861 707 862
rect 751 866 755 867
rect 751 861 755 862
rect 767 866 771 867
rect 778 863 779 867
rect 783 863 784 867
rect 778 862 784 863
rect 807 866 811 867
rect 767 861 771 862
rect 416 859 418 861
rect 448 859 450 861
rect 480 859 482 861
rect 512 859 514 861
rect 552 859 554 861
rect 600 859 602 861
rect 648 859 650 861
rect 704 859 706 861
rect 768 859 770 861
rect 414 858 420 859
rect 414 854 415 858
rect 419 854 420 858
rect 414 853 420 854
rect 446 858 452 859
rect 446 854 447 858
rect 451 854 452 858
rect 446 853 452 854
rect 478 858 484 859
rect 478 854 479 858
rect 483 854 484 858
rect 510 858 516 859
rect 478 853 484 854
rect 498 855 504 856
rect 498 851 499 855
rect 503 851 504 855
rect 510 854 511 858
rect 515 854 516 858
rect 510 853 516 854
rect 550 858 556 859
rect 550 854 551 858
rect 555 854 556 858
rect 550 853 556 854
rect 598 858 604 859
rect 598 854 599 858
rect 603 854 604 858
rect 598 853 604 854
rect 646 858 652 859
rect 646 854 647 858
rect 651 854 652 858
rect 646 853 652 854
rect 702 858 708 859
rect 702 854 703 858
rect 707 854 708 858
rect 702 853 708 854
rect 766 858 772 859
rect 766 854 767 858
rect 771 854 772 858
rect 766 853 772 854
rect 498 850 504 851
rect 396 844 402 846
rect 396 843 397 844
rect 391 842 397 843
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 206 832 212 833
rect 112 827 114 830
rect 206 828 207 832
rect 211 828 212 832
rect 206 827 212 828
rect 230 832 236 833
rect 230 828 231 832
rect 235 828 236 832
rect 230 827 236 828
rect 254 832 260 833
rect 254 828 255 832
rect 259 828 260 832
rect 254 827 260 828
rect 286 832 292 833
rect 286 828 287 832
rect 291 828 292 832
rect 286 827 292 828
rect 318 832 324 833
rect 318 828 319 832
rect 323 828 324 832
rect 318 827 324 828
rect 350 832 356 833
rect 350 828 351 832
rect 355 828 356 832
rect 350 827 356 828
rect 382 832 388 833
rect 382 828 383 832
rect 387 828 388 832
rect 382 827 388 828
rect 414 832 420 833
rect 414 828 415 832
rect 419 828 420 832
rect 414 827 420 828
rect 446 832 452 833
rect 446 828 447 832
rect 451 828 452 832
rect 446 827 452 828
rect 478 832 484 833
rect 478 828 479 832
rect 483 828 484 832
rect 478 827 484 828
rect 111 826 115 827
rect 111 821 115 822
rect 135 826 139 827
rect 135 821 139 822
rect 159 826 163 827
rect 159 821 163 822
rect 183 826 187 827
rect 183 821 187 822
rect 207 826 211 827
rect 207 821 211 822
rect 215 826 219 827
rect 215 821 219 822
rect 231 826 235 827
rect 231 821 235 822
rect 255 826 259 827
rect 255 821 259 822
rect 263 826 267 827
rect 263 821 267 822
rect 287 826 291 827
rect 287 821 291 822
rect 311 826 315 827
rect 311 821 315 822
rect 319 826 323 827
rect 319 821 323 822
rect 351 826 355 827
rect 351 821 355 822
rect 367 826 371 827
rect 367 821 371 822
rect 383 826 387 827
rect 383 821 387 822
rect 415 826 419 827
rect 415 821 419 822
rect 431 826 435 827
rect 431 821 435 822
rect 447 826 451 827
rect 447 821 451 822
rect 479 826 483 827
rect 479 821 483 822
rect 487 826 491 827
rect 487 821 491 822
rect 112 818 114 821
rect 134 820 140 821
rect 110 817 116 818
rect 110 813 111 817
rect 115 813 116 817
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 158 820 164 821
rect 158 816 159 820
rect 163 816 164 820
rect 158 815 164 816
rect 182 820 188 821
rect 182 816 183 820
rect 187 816 188 820
rect 182 815 188 816
rect 214 820 220 821
rect 214 816 215 820
rect 219 816 220 820
rect 214 815 220 816
rect 262 820 268 821
rect 262 816 263 820
rect 267 816 268 820
rect 262 815 268 816
rect 310 820 316 821
rect 310 816 311 820
rect 315 816 316 820
rect 310 815 316 816
rect 366 820 372 821
rect 366 816 367 820
rect 371 816 372 820
rect 366 815 372 816
rect 430 820 436 821
rect 430 816 431 820
rect 435 816 436 820
rect 430 815 436 816
rect 486 820 492 821
rect 486 816 487 820
rect 491 816 492 820
rect 486 815 492 816
rect 110 812 116 813
rect 500 812 502 850
rect 666 847 672 848
rect 666 843 667 847
rect 671 843 672 847
rect 666 842 672 843
rect 510 832 516 833
rect 550 832 556 833
rect 510 828 511 832
rect 515 828 516 832
rect 510 827 516 828
rect 534 831 540 832
rect 534 827 535 831
rect 539 827 540 831
rect 550 828 551 832
rect 555 828 556 832
rect 550 827 556 828
rect 598 832 604 833
rect 598 828 599 832
rect 603 828 604 832
rect 598 827 604 828
rect 646 832 652 833
rect 646 828 647 832
rect 651 828 652 832
rect 646 827 652 828
rect 511 826 515 827
rect 534 826 540 827
rect 543 826 547 827
rect 511 821 515 822
rect 418 811 424 812
rect 418 807 419 811
rect 423 807 424 811
rect 418 806 424 807
rect 498 811 504 812
rect 498 807 499 811
rect 503 807 504 811
rect 498 806 504 807
rect 110 799 116 800
rect 110 795 111 799
rect 115 795 116 799
rect 110 794 116 795
rect 134 794 140 795
rect 112 787 114 794
rect 134 790 135 794
rect 139 790 140 794
rect 134 789 140 790
rect 158 794 164 795
rect 158 790 159 794
rect 163 790 164 794
rect 158 789 164 790
rect 182 794 188 795
rect 182 790 183 794
rect 187 790 188 794
rect 182 789 188 790
rect 214 794 220 795
rect 214 790 215 794
rect 219 790 220 794
rect 214 789 220 790
rect 262 794 268 795
rect 262 790 263 794
rect 267 790 268 794
rect 262 789 268 790
rect 310 794 316 795
rect 310 790 311 794
rect 315 790 316 794
rect 310 789 316 790
rect 366 794 372 795
rect 366 790 367 794
rect 371 790 372 794
rect 366 789 372 790
rect 136 787 138 789
rect 160 787 162 789
rect 184 787 186 789
rect 216 787 218 789
rect 264 787 266 789
rect 312 787 314 789
rect 368 787 370 789
rect 111 786 115 787
rect 111 781 115 782
rect 135 786 139 787
rect 135 781 139 782
rect 159 786 163 787
rect 159 781 163 782
rect 183 786 187 787
rect 183 781 187 782
rect 215 786 219 787
rect 215 781 219 782
rect 223 786 227 787
rect 223 781 227 782
rect 263 786 267 787
rect 263 781 267 782
rect 279 786 283 787
rect 279 781 283 782
rect 311 786 315 787
rect 311 781 315 782
rect 343 786 347 787
rect 343 781 347 782
rect 367 786 371 787
rect 367 781 371 782
rect 407 786 411 787
rect 407 781 411 782
rect 112 774 114 781
rect 136 779 138 781
rect 160 779 162 781
rect 184 779 186 781
rect 224 779 226 781
rect 280 779 282 781
rect 344 779 346 781
rect 408 779 410 781
rect 420 780 422 806
rect 430 794 436 795
rect 430 790 431 794
rect 435 790 436 794
rect 430 789 436 790
rect 486 794 492 795
rect 486 790 487 794
rect 491 790 492 794
rect 486 789 492 790
rect 432 787 434 789
rect 488 787 490 789
rect 536 788 538 826
rect 543 821 547 822
rect 551 826 555 827
rect 551 821 555 822
rect 599 826 603 827
rect 599 821 603 822
rect 647 826 651 827
rect 647 821 651 822
rect 655 826 659 827
rect 655 821 659 822
rect 542 820 548 821
rect 542 816 543 820
rect 547 816 548 820
rect 542 815 548 816
rect 598 820 604 821
rect 598 816 599 820
rect 603 816 604 820
rect 598 815 604 816
rect 654 820 660 821
rect 668 820 670 842
rect 780 836 782 862
rect 807 861 811 862
rect 839 866 843 867
rect 839 861 843 862
rect 863 866 867 867
rect 863 861 867 862
rect 911 866 915 867
rect 911 861 915 862
rect 927 866 931 867
rect 927 861 931 862
rect 983 866 987 867
rect 983 861 987 862
rect 991 866 995 867
rect 991 861 995 862
rect 1047 866 1051 867
rect 1047 861 1051 862
rect 1055 866 1059 867
rect 1055 861 1059 862
rect 1103 866 1107 867
rect 1103 861 1107 862
rect 1119 866 1123 867
rect 1119 861 1123 862
rect 1159 866 1163 867
rect 1159 861 1163 862
rect 1175 866 1179 867
rect 1182 863 1183 867
rect 1187 863 1188 867
rect 1182 862 1188 863
rect 1175 861 1179 862
rect 840 859 842 861
rect 912 859 914 861
rect 984 859 986 861
rect 1048 859 1050 861
rect 1104 859 1106 861
rect 1150 859 1156 860
rect 1160 859 1162 861
rect 838 858 844 859
rect 838 854 839 858
rect 843 854 844 858
rect 838 853 844 854
rect 910 858 916 859
rect 910 854 911 858
rect 915 854 916 858
rect 910 853 916 854
rect 982 858 988 859
rect 982 854 983 858
rect 987 854 988 858
rect 982 853 988 854
rect 1046 858 1052 859
rect 1046 854 1047 858
rect 1051 854 1052 858
rect 1046 853 1052 854
rect 1102 858 1108 859
rect 1102 854 1103 858
rect 1107 854 1108 858
rect 1150 855 1151 859
rect 1155 855 1156 859
rect 1150 854 1156 855
rect 1158 858 1164 859
rect 1158 854 1159 858
rect 1163 854 1164 858
rect 1102 853 1108 854
rect 778 835 784 836
rect 702 832 708 833
rect 702 828 703 832
rect 707 828 708 832
rect 702 827 708 828
rect 766 832 772 833
rect 766 828 767 832
rect 771 828 772 832
rect 778 831 779 835
rect 783 831 784 835
rect 778 830 784 831
rect 838 832 844 833
rect 910 832 916 833
rect 766 827 772 828
rect 838 828 839 832
rect 843 828 844 832
rect 838 827 844 828
rect 850 831 856 832
rect 850 827 851 831
rect 855 827 856 831
rect 910 828 911 832
rect 915 828 916 832
rect 910 827 916 828
rect 982 832 988 833
rect 982 828 983 832
rect 987 828 988 832
rect 982 827 988 828
rect 1046 832 1052 833
rect 1046 828 1047 832
rect 1051 828 1052 832
rect 1046 827 1052 828
rect 1102 832 1108 833
rect 1102 828 1103 832
rect 1107 828 1108 832
rect 1102 827 1108 828
rect 703 826 707 827
rect 703 821 707 822
rect 711 826 715 827
rect 711 821 715 822
rect 767 826 771 827
rect 767 821 771 822
rect 815 826 819 827
rect 815 821 819 822
rect 839 826 843 827
rect 850 826 856 827
rect 863 826 867 827
rect 839 821 843 822
rect 710 820 716 821
rect 654 816 655 820
rect 659 816 660 820
rect 654 815 660 816
rect 666 819 672 820
rect 666 815 667 819
rect 671 815 672 819
rect 710 816 711 820
rect 715 816 716 820
rect 710 815 716 816
rect 766 820 772 821
rect 766 816 767 820
rect 771 816 772 820
rect 766 815 772 816
rect 814 820 820 821
rect 814 816 815 820
rect 819 816 820 820
rect 814 815 820 816
rect 666 814 672 815
rect 610 811 616 812
rect 610 807 611 811
rect 615 807 616 811
rect 610 806 616 807
rect 778 811 784 812
rect 778 807 779 811
rect 783 807 784 811
rect 778 806 784 807
rect 612 796 614 806
rect 780 796 782 806
rect 806 803 812 804
rect 806 799 807 803
rect 811 799 812 803
rect 806 798 812 799
rect 610 795 616 796
rect 778 795 784 796
rect 542 794 548 795
rect 542 790 543 794
rect 547 790 548 794
rect 542 789 548 790
rect 598 794 604 795
rect 598 790 599 794
rect 603 790 604 794
rect 610 791 611 795
rect 615 791 616 795
rect 610 790 616 791
rect 654 794 660 795
rect 654 790 655 794
rect 659 790 660 794
rect 598 789 604 790
rect 654 789 660 790
rect 710 794 716 795
rect 710 790 711 794
rect 715 790 716 794
rect 766 794 772 795
rect 710 789 716 790
rect 730 791 736 792
rect 534 787 540 788
rect 544 787 546 789
rect 600 787 602 789
rect 656 787 658 789
rect 712 787 714 789
rect 730 787 731 791
rect 735 787 736 791
rect 766 790 767 794
rect 771 790 772 794
rect 778 791 779 795
rect 783 791 784 795
rect 778 790 784 791
rect 766 789 772 790
rect 768 787 770 789
rect 431 786 435 787
rect 431 781 435 782
rect 463 786 467 787
rect 463 781 467 782
rect 487 786 491 787
rect 487 781 491 782
rect 519 786 523 787
rect 534 783 535 787
rect 539 783 540 787
rect 534 782 540 783
rect 543 786 547 787
rect 519 781 523 782
rect 543 781 547 782
rect 575 786 579 787
rect 575 781 579 782
rect 599 786 603 787
rect 599 781 603 782
rect 623 786 627 787
rect 623 781 627 782
rect 655 786 659 787
rect 655 781 659 782
rect 671 786 675 787
rect 671 781 675 782
rect 711 786 715 787
rect 711 781 715 782
rect 719 786 723 787
rect 730 786 736 787
rect 759 786 763 787
rect 719 781 723 782
rect 418 779 424 780
rect 464 779 466 781
rect 520 779 522 781
rect 576 779 578 781
rect 624 779 626 781
rect 672 779 674 781
rect 720 779 722 781
rect 134 778 140 779
rect 134 774 135 778
rect 139 774 140 778
rect 110 773 116 774
rect 134 773 140 774
rect 158 778 164 779
rect 158 774 159 778
rect 163 774 164 778
rect 158 773 164 774
rect 182 778 188 779
rect 182 774 183 778
rect 187 774 188 778
rect 182 773 188 774
rect 222 778 228 779
rect 222 774 223 778
rect 227 774 228 778
rect 222 773 228 774
rect 278 778 284 779
rect 278 774 279 778
rect 283 774 284 778
rect 278 773 284 774
rect 342 778 348 779
rect 342 774 343 778
rect 347 774 348 778
rect 342 773 348 774
rect 406 778 412 779
rect 406 774 407 778
rect 411 774 412 778
rect 418 775 419 779
rect 423 775 424 779
rect 418 774 424 775
rect 462 778 468 779
rect 462 774 463 778
rect 467 774 468 778
rect 518 778 524 779
rect 406 773 412 774
rect 462 773 468 774
rect 510 775 516 776
rect 110 769 111 773
rect 115 769 116 773
rect 510 771 511 775
rect 515 771 516 775
rect 518 774 519 778
rect 523 774 524 778
rect 518 773 524 774
rect 574 778 580 779
rect 574 774 575 778
rect 579 774 580 778
rect 574 773 580 774
rect 622 778 628 779
rect 622 774 623 778
rect 627 774 628 778
rect 670 778 676 779
rect 622 773 628 774
rect 634 775 640 776
rect 634 771 635 775
rect 639 771 640 775
rect 670 774 671 778
rect 675 774 676 778
rect 670 773 676 774
rect 718 778 724 779
rect 718 774 719 778
rect 723 774 724 778
rect 718 773 724 774
rect 510 770 516 771
rect 628 770 640 771
rect 110 768 116 769
rect 110 755 116 756
rect 110 751 111 755
rect 115 751 116 755
rect 110 750 116 751
rect 134 752 140 753
rect 158 752 164 753
rect 112 743 114 750
rect 134 748 135 752
rect 139 748 140 752
rect 134 747 140 748
rect 146 751 152 752
rect 146 747 147 751
rect 151 747 152 751
rect 158 748 159 752
rect 163 748 164 752
rect 158 747 164 748
rect 182 752 188 753
rect 182 748 183 752
rect 187 748 188 752
rect 182 747 188 748
rect 222 752 228 753
rect 222 748 223 752
rect 227 748 228 752
rect 222 747 228 748
rect 278 752 284 753
rect 278 748 279 752
rect 283 748 284 752
rect 278 747 284 748
rect 342 752 348 753
rect 342 748 343 752
rect 347 748 348 752
rect 342 747 348 748
rect 406 752 412 753
rect 406 748 407 752
rect 411 748 412 752
rect 406 747 412 748
rect 462 752 468 753
rect 462 748 463 752
rect 467 748 468 752
rect 462 747 468 748
rect 126 743 132 744
rect 136 743 138 747
rect 146 746 152 747
rect 111 742 115 743
rect 126 739 127 743
rect 131 739 132 743
rect 126 738 132 739
rect 135 742 139 743
rect 111 737 115 738
rect 112 734 114 737
rect 110 733 116 734
rect 110 729 111 733
rect 115 729 116 733
rect 110 728 116 729
rect 110 715 116 716
rect 110 711 111 715
rect 115 711 116 715
rect 110 710 116 711
rect 112 703 114 710
rect 128 704 130 738
rect 135 737 139 738
rect 134 736 140 737
rect 134 732 135 736
rect 139 732 140 736
rect 134 731 140 732
rect 148 712 150 746
rect 160 743 162 747
rect 184 743 186 747
rect 224 743 226 747
rect 280 743 282 747
rect 344 743 346 747
rect 408 743 410 747
rect 464 743 466 747
rect 512 744 514 770
rect 628 769 638 770
rect 628 764 630 769
rect 732 768 734 786
rect 759 781 763 782
rect 767 786 771 787
rect 767 781 771 782
rect 799 786 803 787
rect 808 784 810 798
rect 852 796 854 826
rect 863 821 867 822
rect 903 826 907 827
rect 903 821 907 822
rect 911 826 915 827
rect 911 821 915 822
rect 935 826 939 827
rect 935 821 939 822
rect 967 826 971 827
rect 967 821 971 822
rect 983 826 987 827
rect 983 821 987 822
rect 991 826 995 827
rect 991 821 995 822
rect 1015 826 1019 827
rect 1015 821 1019 822
rect 1039 826 1043 827
rect 1039 821 1043 822
rect 1047 826 1051 827
rect 1047 821 1051 822
rect 1063 826 1067 827
rect 1063 821 1067 822
rect 1095 826 1099 827
rect 1095 821 1099 822
rect 1103 826 1107 827
rect 1103 821 1107 822
rect 1127 826 1131 827
rect 1127 821 1131 822
rect 862 820 868 821
rect 862 816 863 820
rect 867 816 868 820
rect 862 815 868 816
rect 902 820 908 821
rect 902 816 903 820
rect 907 816 908 820
rect 902 815 908 816
rect 934 820 940 821
rect 934 816 935 820
rect 939 816 940 820
rect 934 815 940 816
rect 966 820 972 821
rect 966 816 967 820
rect 971 816 972 820
rect 966 815 972 816
rect 990 820 996 821
rect 990 816 991 820
rect 995 816 996 820
rect 990 815 996 816
rect 1014 820 1020 821
rect 1014 816 1015 820
rect 1019 816 1020 820
rect 1014 815 1020 816
rect 1038 820 1044 821
rect 1038 816 1039 820
rect 1043 816 1044 820
rect 1038 815 1044 816
rect 1062 820 1068 821
rect 1062 816 1063 820
rect 1067 816 1068 820
rect 1062 815 1068 816
rect 1094 820 1100 821
rect 1094 816 1095 820
rect 1099 816 1100 820
rect 1094 815 1100 816
rect 1126 820 1132 821
rect 1126 816 1127 820
rect 1131 816 1132 820
rect 1126 815 1132 816
rect 946 811 952 812
rect 946 807 947 811
rect 951 807 952 811
rect 946 806 952 807
rect 1002 811 1008 812
rect 1002 807 1003 811
rect 1007 807 1008 811
rect 1002 806 1008 807
rect 1050 811 1056 812
rect 1050 807 1051 811
rect 1055 807 1056 811
rect 1050 806 1056 807
rect 1074 811 1080 812
rect 1074 807 1075 811
rect 1079 807 1080 811
rect 1074 806 1080 807
rect 1102 807 1108 808
rect 948 796 950 806
rect 1004 796 1006 806
rect 1052 796 1054 806
rect 1076 796 1078 806
rect 1102 803 1103 807
rect 1107 803 1108 807
rect 1102 802 1108 803
rect 850 795 856 796
rect 946 795 952 796
rect 1002 795 1008 796
rect 1050 795 1056 796
rect 1074 795 1080 796
rect 814 794 820 795
rect 814 790 815 794
rect 819 790 820 794
rect 850 791 851 795
rect 855 791 856 795
rect 850 790 856 791
rect 862 794 868 795
rect 862 790 863 794
rect 867 790 868 794
rect 814 789 820 790
rect 862 789 868 790
rect 902 794 908 795
rect 902 790 903 794
rect 907 790 908 794
rect 902 789 908 790
rect 934 794 940 795
rect 934 790 935 794
rect 939 790 940 794
rect 946 791 947 795
rect 951 791 952 795
rect 946 790 952 791
rect 966 794 972 795
rect 966 790 967 794
rect 971 790 972 794
rect 934 789 940 790
rect 966 789 972 790
rect 990 794 996 795
rect 990 790 991 794
rect 995 790 996 794
rect 1002 791 1003 795
rect 1007 791 1008 795
rect 1002 790 1008 791
rect 1014 794 1020 795
rect 1014 790 1015 794
rect 1019 790 1020 794
rect 990 789 996 790
rect 1014 789 1020 790
rect 1038 794 1044 795
rect 1038 790 1039 794
rect 1043 790 1044 794
rect 1050 791 1051 795
rect 1055 791 1056 795
rect 1050 790 1056 791
rect 1062 794 1068 795
rect 1062 790 1063 794
rect 1067 790 1068 794
rect 1074 791 1075 795
rect 1079 791 1080 795
rect 1074 790 1080 791
rect 1094 794 1100 795
rect 1094 790 1095 794
rect 1099 790 1100 794
rect 1038 789 1044 790
rect 1062 789 1068 790
rect 1094 789 1100 790
rect 816 787 818 789
rect 864 787 866 789
rect 904 787 906 789
rect 936 787 938 789
rect 950 787 956 788
rect 968 787 970 789
rect 992 787 994 789
rect 1016 787 1018 789
rect 1040 787 1042 789
rect 1064 787 1066 789
rect 1096 787 1098 789
rect 815 786 819 787
rect 799 781 803 782
rect 806 783 812 784
rect 760 779 762 781
rect 800 779 802 781
rect 806 779 807 783
rect 811 779 812 783
rect 815 781 819 782
rect 839 786 843 787
rect 839 781 843 782
rect 863 786 867 787
rect 863 781 867 782
rect 879 786 883 787
rect 879 781 883 782
rect 903 786 907 787
rect 903 781 907 782
rect 919 786 923 787
rect 919 781 923 782
rect 935 786 939 787
rect 950 783 951 787
rect 955 783 956 787
rect 950 782 956 783
rect 959 786 963 787
rect 935 781 939 782
rect 840 779 842 781
rect 880 779 882 781
rect 920 779 922 781
rect 758 778 764 779
rect 758 774 759 778
rect 763 774 764 778
rect 758 773 764 774
rect 798 778 804 779
rect 806 778 812 779
rect 838 778 844 779
rect 798 774 799 778
rect 803 774 804 778
rect 798 773 804 774
rect 838 774 839 778
rect 843 774 844 778
rect 878 778 884 779
rect 838 773 844 774
rect 862 775 868 776
rect 862 771 863 775
rect 867 771 868 775
rect 878 774 879 778
rect 883 774 884 778
rect 878 773 884 774
rect 918 778 924 779
rect 918 774 919 778
rect 923 774 924 778
rect 918 773 924 774
rect 862 770 868 771
rect 622 763 630 764
rect 622 759 623 763
rect 627 761 630 763
rect 730 767 736 768
rect 730 763 731 767
rect 735 763 736 767
rect 730 762 736 763
rect 627 759 628 761
rect 622 758 628 759
rect 518 752 524 753
rect 518 748 519 752
rect 523 748 524 752
rect 518 747 524 748
rect 574 752 580 753
rect 574 748 575 752
rect 579 748 580 752
rect 574 747 580 748
rect 622 752 628 753
rect 622 748 623 752
rect 627 748 628 752
rect 622 747 628 748
rect 670 752 676 753
rect 670 748 671 752
rect 675 748 676 752
rect 670 747 676 748
rect 718 752 724 753
rect 718 748 719 752
rect 723 748 724 752
rect 718 747 724 748
rect 758 752 764 753
rect 798 752 804 753
rect 758 748 759 752
rect 763 748 764 752
rect 758 747 764 748
rect 770 751 776 752
rect 770 747 771 751
rect 775 747 776 751
rect 798 748 799 752
rect 803 748 804 752
rect 798 747 804 748
rect 838 752 844 753
rect 838 748 839 752
rect 843 748 844 752
rect 838 747 844 748
rect 510 743 516 744
rect 520 743 522 747
rect 576 743 578 747
rect 624 743 626 747
rect 672 743 674 747
rect 720 743 722 747
rect 760 743 762 747
rect 770 746 776 747
rect 159 742 163 743
rect 159 737 163 738
rect 183 742 187 743
rect 183 737 187 738
rect 215 742 219 743
rect 215 737 219 738
rect 223 742 227 743
rect 223 737 227 738
rect 263 742 267 743
rect 263 737 267 738
rect 279 742 283 743
rect 279 737 283 738
rect 319 742 323 743
rect 319 737 323 738
rect 343 742 347 743
rect 343 737 347 738
rect 375 742 379 743
rect 375 737 379 738
rect 407 742 411 743
rect 407 737 411 738
rect 423 742 427 743
rect 423 737 427 738
rect 463 742 467 743
rect 463 737 467 738
rect 471 742 475 743
rect 510 739 511 743
rect 515 739 516 743
rect 510 738 516 739
rect 519 742 523 743
rect 471 737 475 738
rect 519 737 523 738
rect 567 742 571 743
rect 567 737 571 738
rect 575 742 579 743
rect 575 737 579 738
rect 615 742 619 743
rect 615 737 619 738
rect 623 742 627 743
rect 623 737 627 738
rect 663 742 667 743
rect 663 737 667 738
rect 671 742 675 743
rect 671 737 675 738
rect 703 742 707 743
rect 703 737 707 738
rect 719 742 723 743
rect 719 737 723 738
rect 751 742 755 743
rect 751 737 755 738
rect 759 742 763 743
rect 759 737 763 738
rect 158 736 164 737
rect 158 732 159 736
rect 163 732 164 736
rect 158 731 164 732
rect 182 736 188 737
rect 182 732 183 736
rect 187 732 188 736
rect 182 731 188 732
rect 214 736 220 737
rect 214 732 215 736
rect 219 732 220 736
rect 214 731 220 732
rect 262 736 268 737
rect 262 732 263 736
rect 267 732 268 736
rect 262 731 268 732
rect 318 736 324 737
rect 318 732 319 736
rect 323 732 324 736
rect 318 731 324 732
rect 374 736 380 737
rect 374 732 375 736
rect 379 732 380 736
rect 374 731 380 732
rect 422 736 428 737
rect 422 732 423 736
rect 427 732 428 736
rect 422 731 428 732
rect 470 736 476 737
rect 470 732 471 736
rect 475 732 476 736
rect 470 731 476 732
rect 518 736 524 737
rect 518 732 519 736
rect 523 732 524 736
rect 518 731 524 732
rect 566 736 572 737
rect 566 732 567 736
rect 571 732 572 736
rect 566 731 572 732
rect 614 736 620 737
rect 614 732 615 736
rect 619 732 620 736
rect 614 731 620 732
rect 662 736 668 737
rect 662 732 663 736
rect 667 732 668 736
rect 662 731 668 732
rect 702 736 708 737
rect 702 732 703 736
rect 707 732 708 736
rect 702 731 708 732
rect 750 736 756 737
rect 750 732 751 736
rect 755 732 756 736
rect 750 731 756 732
rect 170 727 176 728
rect 170 723 171 727
rect 175 723 176 727
rect 170 722 176 723
rect 226 727 232 728
rect 226 723 227 727
rect 231 723 232 727
rect 226 722 232 723
rect 330 727 336 728
rect 330 723 331 727
rect 335 723 336 727
rect 330 722 336 723
rect 482 727 488 728
rect 482 723 483 727
rect 487 723 488 727
rect 482 722 488 723
rect 578 727 584 728
rect 578 723 579 727
rect 583 723 584 727
rect 578 722 584 723
rect 674 727 680 728
rect 674 723 675 727
rect 679 723 680 727
rect 674 722 680 723
rect 172 712 174 722
rect 228 712 230 722
rect 332 712 334 722
rect 484 712 486 722
rect 580 712 582 722
rect 676 712 678 722
rect 772 712 774 746
rect 800 743 802 747
rect 840 743 842 747
rect 864 744 866 770
rect 952 756 954 782
rect 959 781 963 782
rect 967 786 971 787
rect 967 781 971 782
rect 991 786 995 787
rect 991 781 995 782
rect 1015 786 1019 787
rect 1015 781 1019 782
rect 1023 786 1027 787
rect 1023 781 1027 782
rect 1039 786 1043 787
rect 1039 781 1043 782
rect 1055 786 1059 787
rect 1055 781 1059 782
rect 1063 786 1067 787
rect 1063 781 1067 782
rect 1087 786 1091 787
rect 1087 781 1091 782
rect 1095 786 1099 787
rect 1095 781 1099 782
rect 960 779 962 781
rect 992 779 994 781
rect 1024 779 1026 781
rect 1056 779 1058 781
rect 1088 779 1090 781
rect 958 778 964 779
rect 958 774 959 778
rect 963 774 964 778
rect 958 773 964 774
rect 990 778 996 779
rect 990 774 991 778
rect 995 774 996 778
rect 1022 778 1028 779
rect 990 773 996 774
rect 1002 775 1008 776
rect 1002 771 1003 775
rect 1007 771 1008 775
rect 1022 774 1023 778
rect 1027 774 1028 778
rect 1022 773 1028 774
rect 1054 778 1060 779
rect 1054 774 1055 778
rect 1059 774 1060 778
rect 1054 773 1060 774
rect 1086 778 1092 779
rect 1086 774 1087 778
rect 1091 774 1092 778
rect 1086 773 1092 774
rect 1002 770 1008 771
rect 950 755 956 756
rect 878 752 884 753
rect 878 748 879 752
rect 883 748 884 752
rect 878 747 884 748
rect 918 752 924 753
rect 918 748 919 752
rect 923 748 924 752
rect 950 751 951 755
rect 955 751 956 755
rect 950 750 956 751
rect 958 752 964 753
rect 918 747 924 748
rect 958 748 959 752
rect 963 748 964 752
rect 958 747 964 748
rect 990 752 996 753
rect 990 748 991 752
rect 995 748 996 752
rect 990 747 996 748
rect 862 743 868 744
rect 880 743 882 747
rect 920 743 922 747
rect 960 743 962 747
rect 992 743 994 747
rect 1004 744 1006 770
rect 1022 752 1028 753
rect 1022 748 1023 752
rect 1027 748 1028 752
rect 1022 747 1028 748
rect 1054 752 1060 753
rect 1054 748 1055 752
rect 1059 748 1060 752
rect 1054 747 1060 748
rect 1086 752 1092 753
rect 1086 748 1087 752
rect 1091 748 1092 752
rect 1086 747 1092 748
rect 1002 743 1008 744
rect 1024 743 1026 747
rect 1056 743 1058 747
rect 1088 743 1090 747
rect 1104 744 1106 802
rect 1126 794 1132 795
rect 1126 790 1127 794
rect 1131 790 1132 794
rect 1126 789 1132 790
rect 1128 787 1130 789
rect 1127 786 1131 787
rect 1152 784 1154 854
rect 1158 853 1164 854
rect 1184 836 1186 862
rect 1200 860 1202 870
rect 1230 869 1236 870
rect 1278 874 1284 875
rect 1278 870 1279 874
rect 1283 870 1284 874
rect 1290 871 1291 875
rect 1295 871 1296 875
rect 1290 870 1296 871
rect 1326 874 1332 875
rect 1326 870 1327 874
rect 1331 870 1332 874
rect 1278 869 1284 870
rect 1326 869 1332 870
rect 1382 874 1388 875
rect 1382 870 1383 874
rect 1387 870 1388 874
rect 1382 869 1388 870
rect 1232 867 1234 869
rect 1280 867 1282 869
rect 1302 867 1308 868
rect 1328 867 1330 869
rect 1384 867 1386 869
rect 1404 868 1406 906
rect 1415 901 1419 902
rect 1447 906 1451 907
rect 1447 901 1451 902
rect 1414 900 1420 901
rect 1414 896 1415 900
rect 1419 896 1420 900
rect 1448 898 1450 901
rect 1414 895 1420 896
rect 1446 897 1452 898
rect 1446 893 1447 897
rect 1451 893 1452 897
rect 1446 892 1452 893
rect 1426 883 1432 884
rect 1426 879 1427 883
rect 1431 879 1432 883
rect 1426 878 1432 879
rect 1446 879 1452 880
rect 1414 874 1420 875
rect 1414 870 1415 874
rect 1419 870 1420 874
rect 1414 869 1420 870
rect 1402 867 1408 868
rect 1416 867 1418 869
rect 1207 866 1211 867
rect 1207 861 1211 862
rect 1231 866 1235 867
rect 1231 861 1235 862
rect 1247 866 1251 867
rect 1247 861 1251 862
rect 1279 866 1283 867
rect 1279 861 1283 862
rect 1295 866 1299 867
rect 1302 863 1303 867
rect 1307 863 1308 867
rect 1302 862 1308 863
rect 1327 866 1331 867
rect 1295 861 1299 862
rect 1198 859 1204 860
rect 1208 859 1210 861
rect 1248 859 1250 861
rect 1296 859 1298 861
rect 1198 855 1199 859
rect 1203 855 1204 859
rect 1198 854 1204 855
rect 1206 858 1212 859
rect 1206 854 1207 858
rect 1211 854 1212 858
rect 1206 853 1212 854
rect 1246 858 1252 859
rect 1246 854 1247 858
rect 1251 854 1252 858
rect 1246 853 1252 854
rect 1294 858 1300 859
rect 1294 854 1295 858
rect 1299 854 1300 858
rect 1294 853 1300 854
rect 1182 835 1188 836
rect 1158 832 1164 833
rect 1158 828 1159 832
rect 1163 828 1164 832
rect 1182 831 1183 835
rect 1187 831 1188 835
rect 1182 830 1188 831
rect 1206 832 1212 833
rect 1158 827 1164 828
rect 1206 828 1207 832
rect 1211 828 1212 832
rect 1206 827 1212 828
rect 1246 832 1252 833
rect 1246 828 1247 832
rect 1251 828 1252 832
rect 1246 827 1252 828
rect 1294 832 1300 833
rect 1294 828 1295 832
rect 1299 828 1300 832
rect 1304 828 1306 862
rect 1327 861 1331 862
rect 1343 866 1347 867
rect 1343 861 1347 862
rect 1383 866 1387 867
rect 1383 861 1387 862
rect 1391 866 1395 867
rect 1402 863 1403 867
rect 1407 863 1408 867
rect 1402 862 1408 863
rect 1415 866 1419 867
rect 1391 861 1395 862
rect 1415 861 1419 862
rect 1344 859 1346 861
rect 1392 859 1394 861
rect 1416 859 1418 861
rect 1428 860 1430 878
rect 1446 875 1447 879
rect 1451 875 1452 879
rect 1446 874 1452 875
rect 1448 867 1450 874
rect 1447 866 1451 867
rect 1447 861 1451 862
rect 1426 859 1432 860
rect 1342 858 1348 859
rect 1342 854 1343 858
rect 1347 854 1348 858
rect 1342 853 1348 854
rect 1390 858 1396 859
rect 1390 854 1391 858
rect 1395 854 1396 858
rect 1390 853 1396 854
rect 1414 858 1420 859
rect 1414 854 1415 858
rect 1419 854 1420 858
rect 1426 855 1427 859
rect 1431 855 1432 859
rect 1426 854 1432 855
rect 1448 854 1450 861
rect 1414 853 1420 854
rect 1446 853 1452 854
rect 1446 849 1447 853
rect 1451 849 1452 853
rect 1446 848 1452 849
rect 1446 835 1452 836
rect 1342 832 1348 833
rect 1342 828 1343 832
rect 1347 828 1348 832
rect 1294 827 1300 828
rect 1302 827 1308 828
rect 1342 827 1348 828
rect 1390 832 1396 833
rect 1414 832 1420 833
rect 1390 828 1391 832
rect 1395 828 1396 832
rect 1390 827 1396 828
rect 1402 831 1408 832
rect 1402 827 1403 831
rect 1407 827 1408 831
rect 1414 828 1415 832
rect 1419 828 1420 832
rect 1446 831 1447 835
rect 1451 831 1452 835
rect 1446 830 1452 831
rect 1414 827 1420 828
rect 1448 827 1450 830
rect 1159 826 1163 827
rect 1159 821 1163 822
rect 1167 826 1171 827
rect 1167 821 1171 822
rect 1207 826 1211 827
rect 1207 821 1211 822
rect 1247 826 1251 827
rect 1247 821 1251 822
rect 1255 826 1259 827
rect 1255 821 1259 822
rect 1295 826 1299 827
rect 1302 823 1303 827
rect 1307 823 1308 827
rect 1302 822 1308 823
rect 1311 826 1315 827
rect 1295 821 1299 822
rect 1311 821 1315 822
rect 1343 826 1347 827
rect 1343 821 1347 822
rect 1375 826 1379 827
rect 1375 821 1379 822
rect 1391 826 1395 827
rect 1402 826 1408 827
rect 1415 826 1419 827
rect 1391 821 1395 822
rect 1166 820 1172 821
rect 1166 816 1167 820
rect 1171 816 1172 820
rect 1166 815 1172 816
rect 1206 820 1212 821
rect 1206 816 1207 820
rect 1211 816 1212 820
rect 1206 815 1212 816
rect 1254 820 1260 821
rect 1254 816 1255 820
rect 1259 816 1260 820
rect 1254 815 1260 816
rect 1310 820 1316 821
rect 1310 816 1311 820
rect 1315 816 1316 820
rect 1310 815 1316 816
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1178 811 1184 812
rect 1178 807 1179 811
rect 1183 807 1184 811
rect 1178 806 1184 807
rect 1266 811 1272 812
rect 1266 807 1267 811
rect 1271 807 1272 811
rect 1266 806 1272 807
rect 1274 811 1280 812
rect 1274 807 1275 811
rect 1279 807 1280 811
rect 1274 806 1280 807
rect 1180 796 1182 806
rect 1268 796 1270 806
rect 1158 795 1164 796
rect 1178 795 1184 796
rect 1266 795 1272 796
rect 1158 791 1159 795
rect 1163 791 1164 795
rect 1158 790 1164 791
rect 1166 794 1172 795
rect 1166 790 1167 794
rect 1171 790 1172 794
rect 1178 791 1179 795
rect 1183 791 1184 795
rect 1178 790 1184 791
rect 1206 794 1212 795
rect 1206 790 1207 794
rect 1211 790 1212 794
rect 1127 781 1131 782
rect 1150 783 1156 784
rect 1128 779 1130 781
rect 1150 779 1151 783
rect 1155 779 1156 783
rect 1126 778 1132 779
rect 1150 778 1156 779
rect 1126 774 1127 778
rect 1131 774 1132 778
rect 1126 773 1132 774
rect 1126 752 1132 753
rect 1126 748 1127 752
rect 1131 748 1132 752
rect 1126 747 1132 748
rect 1102 743 1108 744
rect 1128 743 1130 747
rect 1160 744 1162 790
rect 1166 789 1172 790
rect 1206 789 1212 790
rect 1254 794 1260 795
rect 1254 790 1255 794
rect 1259 790 1260 794
rect 1266 791 1267 795
rect 1271 791 1272 795
rect 1266 790 1272 791
rect 1254 789 1260 790
rect 1168 787 1170 789
rect 1208 787 1210 789
rect 1256 787 1258 789
rect 1276 788 1278 806
rect 1404 796 1406 826
rect 1415 821 1419 822
rect 1447 826 1451 827
rect 1447 821 1451 822
rect 1414 820 1420 821
rect 1414 816 1415 820
rect 1419 816 1420 820
rect 1448 818 1450 821
rect 1414 815 1420 816
rect 1446 817 1452 818
rect 1446 813 1447 817
rect 1451 813 1452 817
rect 1446 812 1452 813
rect 1426 803 1432 804
rect 1426 799 1427 803
rect 1431 799 1432 803
rect 1426 798 1432 799
rect 1446 799 1452 800
rect 1402 795 1408 796
rect 1310 794 1316 795
rect 1310 790 1311 794
rect 1315 790 1316 794
rect 1310 789 1316 790
rect 1374 794 1380 795
rect 1374 790 1375 794
rect 1379 790 1380 794
rect 1402 791 1403 795
rect 1407 791 1408 795
rect 1402 790 1408 791
rect 1414 794 1420 795
rect 1414 790 1415 794
rect 1419 790 1420 794
rect 1374 789 1380 790
rect 1414 789 1420 790
rect 1274 787 1280 788
rect 1312 787 1314 789
rect 1376 787 1378 789
rect 1416 787 1418 789
rect 1167 786 1171 787
rect 1167 781 1171 782
rect 1175 786 1179 787
rect 1175 781 1179 782
rect 1207 786 1211 787
rect 1207 781 1211 782
rect 1231 786 1235 787
rect 1231 781 1235 782
rect 1255 786 1259 787
rect 1274 783 1275 787
rect 1279 783 1280 787
rect 1274 782 1280 783
rect 1295 786 1299 787
rect 1255 781 1259 782
rect 1295 781 1299 782
rect 1311 786 1315 787
rect 1311 781 1315 782
rect 1367 786 1371 787
rect 1367 781 1371 782
rect 1375 786 1379 787
rect 1375 781 1379 782
rect 1415 786 1419 787
rect 1415 781 1419 782
rect 1176 779 1178 781
rect 1232 779 1234 781
rect 1296 779 1298 781
rect 1368 779 1370 781
rect 1416 779 1418 781
rect 1428 780 1430 798
rect 1446 795 1447 799
rect 1451 795 1452 799
rect 1446 794 1452 795
rect 1448 787 1450 794
rect 1447 786 1451 787
rect 1447 781 1451 782
rect 1426 779 1432 780
rect 1174 778 1180 779
rect 1174 774 1175 778
rect 1179 774 1180 778
rect 1174 773 1180 774
rect 1230 778 1236 779
rect 1230 774 1231 778
rect 1235 774 1236 778
rect 1230 773 1236 774
rect 1294 778 1300 779
rect 1294 774 1295 778
rect 1299 774 1300 778
rect 1294 773 1300 774
rect 1366 778 1372 779
rect 1366 774 1367 778
rect 1371 774 1372 778
rect 1366 773 1372 774
rect 1414 778 1420 779
rect 1414 774 1415 778
rect 1419 774 1420 778
rect 1426 775 1427 779
rect 1431 775 1432 779
rect 1426 774 1432 775
rect 1448 774 1450 781
rect 1414 773 1420 774
rect 1446 773 1452 774
rect 1446 769 1447 773
rect 1451 769 1452 773
rect 1446 768 1452 769
rect 1446 755 1452 756
rect 1174 752 1180 753
rect 1174 748 1175 752
rect 1179 748 1180 752
rect 1174 747 1180 748
rect 1230 752 1236 753
rect 1230 748 1231 752
rect 1235 748 1236 752
rect 1230 747 1236 748
rect 1294 752 1300 753
rect 1294 748 1295 752
rect 1299 748 1300 752
rect 1294 747 1300 748
rect 1366 752 1372 753
rect 1366 748 1367 752
rect 1371 748 1372 752
rect 1414 752 1420 753
rect 1414 748 1415 752
rect 1419 748 1420 752
rect 1446 751 1447 755
rect 1451 751 1452 755
rect 1446 750 1452 751
rect 1366 747 1372 748
rect 1374 747 1380 748
rect 1414 747 1420 748
rect 1158 743 1164 744
rect 1176 743 1178 747
rect 1232 743 1234 747
rect 1296 743 1298 747
rect 1368 743 1370 747
rect 1374 743 1375 747
rect 1379 743 1380 747
rect 1416 743 1418 747
rect 1448 743 1450 750
rect 799 742 803 743
rect 799 737 803 738
rect 807 742 811 743
rect 807 737 811 738
rect 839 742 843 743
rect 862 739 863 743
rect 867 739 868 743
rect 862 738 868 739
rect 871 742 875 743
rect 839 737 843 738
rect 871 737 875 738
rect 879 742 883 743
rect 879 737 883 738
rect 919 742 923 743
rect 919 737 923 738
rect 943 742 947 743
rect 943 737 947 738
rect 959 742 963 743
rect 959 737 963 738
rect 991 742 995 743
rect 1002 739 1003 743
rect 1007 739 1008 743
rect 1002 738 1008 739
rect 1015 742 1019 743
rect 991 737 995 738
rect 1015 737 1019 738
rect 1023 742 1027 743
rect 1023 737 1027 738
rect 1055 742 1059 743
rect 1055 737 1059 738
rect 1087 742 1091 743
rect 1102 739 1103 743
rect 1107 739 1108 743
rect 1102 738 1108 739
rect 1127 742 1131 743
rect 1087 737 1091 738
rect 1127 737 1131 738
rect 1151 742 1155 743
rect 1158 739 1159 743
rect 1163 739 1164 743
rect 1158 738 1164 739
rect 1175 742 1179 743
rect 1151 737 1155 738
rect 1175 737 1179 738
rect 1215 742 1219 743
rect 1215 737 1219 738
rect 1231 742 1235 743
rect 1231 737 1235 738
rect 1271 742 1275 743
rect 1271 737 1275 738
rect 1295 742 1299 743
rect 1295 737 1299 738
rect 1327 742 1331 743
rect 1327 737 1331 738
rect 1367 742 1371 743
rect 1374 742 1380 743
rect 1383 742 1387 743
rect 1367 737 1371 738
rect 806 736 812 737
rect 806 732 807 736
rect 811 732 812 736
rect 806 731 812 732
rect 870 736 876 737
rect 870 732 871 736
rect 875 732 876 736
rect 870 731 876 732
rect 942 736 948 737
rect 942 732 943 736
rect 947 732 948 736
rect 942 731 948 732
rect 1014 736 1020 737
rect 1014 732 1015 736
rect 1019 732 1020 736
rect 1014 731 1020 732
rect 1086 736 1092 737
rect 1086 732 1087 736
rect 1091 732 1092 736
rect 1086 731 1092 732
rect 1150 736 1156 737
rect 1150 732 1151 736
rect 1155 732 1156 736
rect 1150 731 1156 732
rect 1214 736 1220 737
rect 1214 732 1215 736
rect 1219 732 1220 736
rect 1214 731 1220 732
rect 1270 736 1276 737
rect 1270 732 1271 736
rect 1275 732 1276 736
rect 1270 731 1276 732
rect 1326 736 1332 737
rect 1326 732 1327 736
rect 1331 732 1332 736
rect 1326 731 1332 732
rect 882 727 888 728
rect 882 723 883 727
rect 887 723 888 727
rect 882 722 888 723
rect 1026 727 1032 728
rect 1026 723 1027 727
rect 1031 723 1032 727
rect 1026 722 1032 723
rect 1050 727 1056 728
rect 1050 723 1051 727
rect 1055 723 1056 727
rect 1050 722 1056 723
rect 1290 727 1296 728
rect 1290 723 1291 727
rect 1295 723 1296 727
rect 1290 722 1296 723
rect 884 712 886 722
rect 1028 712 1030 722
rect 146 711 152 712
rect 170 711 176 712
rect 226 711 232 712
rect 330 711 336 712
rect 482 711 488 712
rect 578 711 584 712
rect 674 711 680 712
rect 770 711 776 712
rect 882 711 888 712
rect 1026 711 1032 712
rect 134 710 140 711
rect 134 706 135 710
rect 139 706 140 710
rect 146 707 147 711
rect 151 707 152 711
rect 146 706 152 707
rect 158 710 164 711
rect 158 706 159 710
rect 163 706 164 710
rect 170 707 171 711
rect 175 707 176 711
rect 170 706 176 707
rect 182 710 188 711
rect 182 706 183 710
rect 187 706 188 710
rect 134 705 140 706
rect 158 705 164 706
rect 182 705 188 706
rect 214 710 220 711
rect 214 706 215 710
rect 219 706 220 710
rect 226 707 227 711
rect 231 707 232 711
rect 226 706 232 707
rect 262 710 268 711
rect 262 706 263 710
rect 267 706 268 710
rect 214 705 220 706
rect 262 705 268 706
rect 318 710 324 711
rect 318 706 319 710
rect 323 706 324 710
rect 330 707 331 711
rect 335 707 336 711
rect 330 706 336 707
rect 374 710 380 711
rect 374 706 375 710
rect 379 706 380 710
rect 318 705 324 706
rect 374 705 380 706
rect 422 710 428 711
rect 422 706 423 710
rect 427 706 428 710
rect 422 705 428 706
rect 470 710 476 711
rect 470 706 471 710
rect 475 706 476 710
rect 482 707 483 711
rect 487 707 488 711
rect 482 706 488 707
rect 518 710 524 711
rect 518 706 519 710
rect 523 706 524 710
rect 470 705 476 706
rect 518 705 524 706
rect 566 710 572 711
rect 566 706 567 710
rect 571 706 572 710
rect 578 707 579 711
rect 583 707 584 711
rect 578 706 584 707
rect 614 710 620 711
rect 614 706 615 710
rect 619 706 620 710
rect 566 705 572 706
rect 614 705 620 706
rect 662 710 668 711
rect 662 706 663 710
rect 667 706 668 710
rect 674 707 675 711
rect 679 707 680 711
rect 674 706 680 707
rect 702 710 708 711
rect 702 706 703 710
rect 707 706 708 710
rect 662 705 668 706
rect 702 705 708 706
rect 750 710 756 711
rect 750 706 751 710
rect 755 706 756 710
rect 770 707 771 711
rect 775 707 776 711
rect 770 706 776 707
rect 806 710 812 711
rect 806 706 807 710
rect 811 706 812 710
rect 870 710 876 711
rect 750 705 756 706
rect 806 705 812 706
rect 838 707 844 708
rect 126 703 132 704
rect 136 703 138 705
rect 160 703 162 705
rect 184 703 186 705
rect 216 703 218 705
rect 264 703 266 705
rect 320 703 322 705
rect 376 703 378 705
rect 424 703 426 705
rect 472 703 474 705
rect 494 703 500 704
rect 520 703 522 705
rect 568 703 570 705
rect 616 703 618 705
rect 664 703 666 705
rect 704 703 706 705
rect 752 703 754 705
rect 808 703 810 705
rect 838 703 839 707
rect 843 703 844 707
rect 870 706 871 710
rect 875 706 876 710
rect 882 707 883 711
rect 887 707 888 711
rect 882 706 888 707
rect 942 710 948 711
rect 942 706 943 710
rect 947 706 948 710
rect 870 705 876 706
rect 942 705 948 706
rect 1014 710 1020 711
rect 1014 706 1015 710
rect 1019 706 1020 710
rect 1026 707 1027 711
rect 1031 707 1032 711
rect 1026 706 1032 707
rect 1014 705 1020 706
rect 111 702 115 703
rect 126 699 127 703
rect 131 699 132 703
rect 126 698 132 699
rect 135 702 139 703
rect 111 697 115 698
rect 135 697 139 698
rect 159 702 163 703
rect 159 697 163 698
rect 183 702 187 703
rect 183 697 187 698
rect 199 702 203 703
rect 199 697 203 698
rect 215 702 219 703
rect 215 697 219 698
rect 239 702 243 703
rect 239 697 243 698
rect 263 702 267 703
rect 263 697 267 698
rect 287 702 291 703
rect 287 697 291 698
rect 319 702 323 703
rect 319 697 323 698
rect 335 702 339 703
rect 335 697 339 698
rect 375 702 379 703
rect 375 697 379 698
rect 391 702 395 703
rect 391 697 395 698
rect 423 702 427 703
rect 423 697 427 698
rect 439 702 443 703
rect 439 697 443 698
rect 471 702 475 703
rect 471 697 475 698
rect 487 702 491 703
rect 494 699 495 703
rect 499 699 500 703
rect 494 698 500 699
rect 519 702 523 703
rect 487 697 491 698
rect 112 690 114 697
rect 136 695 138 697
rect 160 695 162 697
rect 200 695 202 697
rect 240 695 242 697
rect 288 695 290 697
rect 336 695 338 697
rect 392 695 394 697
rect 440 695 442 697
rect 488 695 490 697
rect 134 694 140 695
rect 134 690 135 694
rect 139 690 140 694
rect 110 689 116 690
rect 134 689 140 690
rect 158 694 164 695
rect 158 690 159 694
rect 163 690 164 694
rect 158 689 164 690
rect 198 694 204 695
rect 198 690 199 694
rect 203 690 204 694
rect 198 689 204 690
rect 238 694 244 695
rect 238 690 239 694
rect 243 690 244 694
rect 238 689 244 690
rect 286 694 292 695
rect 286 690 287 694
rect 291 690 292 694
rect 286 689 292 690
rect 334 694 340 695
rect 334 690 335 694
rect 339 690 340 694
rect 334 689 340 690
rect 390 694 396 695
rect 390 690 391 694
rect 395 690 396 694
rect 438 694 444 695
rect 390 689 396 690
rect 430 691 436 692
rect 110 685 111 689
rect 115 685 116 689
rect 430 687 431 691
rect 435 687 436 691
rect 438 690 439 694
rect 443 690 444 694
rect 486 694 492 695
rect 438 689 444 690
rect 450 691 456 692
rect 430 686 436 687
rect 450 687 451 691
rect 455 687 456 691
rect 486 690 487 694
rect 491 690 492 694
rect 486 689 492 690
rect 450 686 456 687
rect 110 684 116 685
rect 110 671 116 672
rect 110 667 111 671
rect 115 667 116 671
rect 110 666 116 667
rect 134 668 140 669
rect 112 663 114 666
rect 134 664 135 668
rect 139 664 140 668
rect 134 663 140 664
rect 158 668 164 669
rect 158 664 159 668
rect 163 664 164 668
rect 158 663 164 664
rect 198 668 204 669
rect 198 664 199 668
rect 203 664 204 668
rect 198 663 204 664
rect 238 668 244 669
rect 238 664 239 668
rect 243 664 244 668
rect 238 663 244 664
rect 286 668 292 669
rect 286 664 287 668
rect 291 664 292 668
rect 286 663 292 664
rect 334 668 340 669
rect 390 668 396 669
rect 334 664 335 668
rect 339 664 340 668
rect 334 663 340 664
rect 346 667 352 668
rect 346 663 347 667
rect 351 663 352 667
rect 390 664 391 668
rect 395 664 396 668
rect 390 663 396 664
rect 111 662 115 663
rect 111 657 115 658
rect 135 662 139 663
rect 135 657 139 658
rect 159 662 163 663
rect 159 657 163 658
rect 191 662 195 663
rect 191 657 195 658
rect 199 662 203 663
rect 199 657 203 658
rect 215 662 219 663
rect 215 657 219 658
rect 239 662 243 663
rect 239 657 243 658
rect 263 662 267 663
rect 263 657 267 658
rect 287 662 291 663
rect 287 657 291 658
rect 295 662 299 663
rect 295 657 299 658
rect 327 662 331 663
rect 327 657 331 658
rect 335 662 339 663
rect 346 662 352 663
rect 367 662 371 663
rect 335 657 339 658
rect 112 654 114 657
rect 190 656 196 657
rect 110 653 116 654
rect 110 649 111 653
rect 115 649 116 653
rect 190 652 191 656
rect 195 652 196 656
rect 190 651 196 652
rect 214 656 220 657
rect 214 652 215 656
rect 219 652 220 656
rect 214 651 220 652
rect 238 656 244 657
rect 238 652 239 656
rect 243 652 244 656
rect 238 651 244 652
rect 262 656 268 657
rect 262 652 263 656
rect 267 652 268 656
rect 262 651 268 652
rect 294 656 300 657
rect 294 652 295 656
rect 299 652 300 656
rect 294 651 300 652
rect 326 656 332 657
rect 326 652 327 656
rect 331 652 332 656
rect 326 651 332 652
rect 110 648 116 649
rect 226 647 232 648
rect 226 643 227 647
rect 231 643 232 647
rect 226 642 232 643
rect 274 647 280 648
rect 274 643 275 647
rect 279 643 280 647
rect 274 642 280 643
rect 338 647 344 648
rect 338 643 339 647
rect 343 643 344 647
rect 338 642 344 643
rect 203 636 207 637
rect 110 635 116 636
rect 110 631 111 635
rect 115 631 116 635
rect 228 632 230 642
rect 276 632 278 642
rect 340 632 342 642
rect 348 637 350 662
rect 367 657 371 658
rect 391 662 395 663
rect 391 657 395 658
rect 407 662 411 663
rect 432 660 434 686
rect 438 683 444 684
rect 452 683 454 686
rect 438 679 439 683
rect 443 681 454 683
rect 443 679 444 681
rect 438 678 444 679
rect 438 668 444 669
rect 438 664 439 668
rect 443 664 444 668
rect 438 663 444 664
rect 486 668 492 669
rect 486 664 487 668
rect 491 664 492 668
rect 496 664 498 698
rect 519 697 523 698
rect 535 702 539 703
rect 535 697 539 698
rect 567 702 571 703
rect 567 697 571 698
rect 583 702 587 703
rect 583 697 587 698
rect 615 702 619 703
rect 615 697 619 698
rect 639 702 643 703
rect 639 697 643 698
rect 663 702 667 703
rect 663 697 667 698
rect 695 702 699 703
rect 695 697 699 698
rect 703 702 707 703
rect 703 697 707 698
rect 751 702 755 703
rect 751 697 755 698
rect 759 702 763 703
rect 759 697 763 698
rect 807 702 811 703
rect 807 697 811 698
rect 831 702 835 703
rect 838 702 844 703
rect 846 703 852 704
rect 872 703 874 705
rect 944 703 946 705
rect 1016 703 1018 705
rect 1052 704 1054 722
rect 1086 710 1092 711
rect 1086 706 1087 710
rect 1091 706 1092 710
rect 1086 705 1092 706
rect 1150 710 1156 711
rect 1150 706 1151 710
rect 1155 706 1156 710
rect 1150 705 1156 706
rect 1214 710 1220 711
rect 1214 706 1215 710
rect 1219 706 1220 710
rect 1214 705 1220 706
rect 1270 710 1276 711
rect 1270 706 1271 710
rect 1275 706 1276 710
rect 1270 705 1276 706
rect 1050 703 1056 704
rect 1088 703 1090 705
rect 1152 703 1154 705
rect 1216 703 1218 705
rect 1272 703 1274 705
rect 831 697 835 698
rect 536 695 538 697
rect 584 695 586 697
rect 640 695 642 697
rect 696 695 698 697
rect 760 695 762 697
rect 832 695 834 697
rect 534 694 540 695
rect 534 690 535 694
rect 539 690 540 694
rect 534 689 540 690
rect 582 694 588 695
rect 582 690 583 694
rect 587 690 588 694
rect 582 689 588 690
rect 638 694 644 695
rect 638 690 639 694
rect 643 690 644 694
rect 638 689 644 690
rect 694 694 700 695
rect 694 690 695 694
rect 699 690 700 694
rect 694 689 700 690
rect 758 694 764 695
rect 758 690 759 694
rect 763 690 764 694
rect 758 689 764 690
rect 830 694 836 695
rect 830 690 831 694
rect 835 690 836 694
rect 830 689 836 690
rect 840 684 842 702
rect 846 699 847 703
rect 851 699 852 703
rect 846 698 852 699
rect 871 702 875 703
rect 838 683 844 684
rect 838 679 839 683
rect 843 679 844 683
rect 838 678 844 679
rect 534 668 540 669
rect 534 664 535 668
rect 539 664 540 668
rect 486 663 492 664
rect 494 663 500 664
rect 534 663 540 664
rect 582 668 588 669
rect 582 664 583 668
rect 587 664 588 668
rect 582 663 588 664
rect 638 668 644 669
rect 694 668 700 669
rect 638 664 639 668
rect 643 664 644 668
rect 638 663 644 664
rect 650 667 656 668
rect 650 663 651 667
rect 655 663 656 667
rect 694 664 695 668
rect 699 664 700 668
rect 694 663 700 664
rect 758 668 764 669
rect 758 664 759 668
rect 763 664 764 668
rect 758 663 764 664
rect 830 668 836 669
rect 830 664 831 668
rect 835 664 836 668
rect 830 663 836 664
rect 439 662 443 663
rect 407 657 411 658
rect 430 659 436 660
rect 366 656 372 657
rect 366 652 367 656
rect 371 652 372 656
rect 366 651 372 652
rect 406 656 412 657
rect 406 652 407 656
rect 411 652 412 656
rect 430 655 431 659
rect 435 655 436 659
rect 439 657 443 658
rect 455 662 459 663
rect 455 657 459 658
rect 487 662 491 663
rect 494 659 495 663
rect 499 659 500 663
rect 494 658 500 659
rect 503 662 507 663
rect 487 657 491 658
rect 503 657 507 658
rect 535 662 539 663
rect 535 657 539 658
rect 551 662 555 663
rect 551 657 555 658
rect 583 662 587 663
rect 583 657 587 658
rect 607 662 611 663
rect 607 657 611 658
rect 639 662 643 663
rect 650 662 656 663
rect 663 662 667 663
rect 639 657 643 658
rect 430 654 436 655
rect 454 656 460 657
rect 406 651 412 652
rect 454 652 455 656
rect 459 652 460 656
rect 454 651 460 652
rect 502 656 508 657
rect 502 652 503 656
rect 507 652 508 656
rect 502 651 508 652
rect 550 656 556 657
rect 550 652 551 656
rect 555 652 556 656
rect 550 651 556 652
rect 606 656 612 657
rect 606 652 607 656
rect 611 652 612 656
rect 606 651 612 652
rect 466 647 472 648
rect 466 643 467 647
rect 471 643 472 647
rect 466 642 472 643
rect 562 647 568 648
rect 562 643 563 647
rect 567 643 568 647
rect 562 642 568 643
rect 347 636 351 637
rect 447 636 451 637
rect 468 632 470 642
rect 531 636 535 637
rect 564 632 566 642
rect 652 632 654 662
rect 663 657 667 658
rect 695 662 699 663
rect 695 657 699 658
rect 719 662 723 663
rect 719 657 723 658
rect 759 662 763 663
rect 759 657 763 658
rect 767 662 771 663
rect 767 657 771 658
rect 815 662 819 663
rect 815 657 819 658
rect 831 662 835 663
rect 831 657 835 658
rect 662 656 668 657
rect 662 652 663 656
rect 667 652 668 656
rect 662 651 668 652
rect 718 656 724 657
rect 718 652 719 656
rect 723 652 724 656
rect 718 651 724 652
rect 766 656 772 657
rect 766 652 767 656
rect 771 652 772 656
rect 766 651 772 652
rect 814 656 820 657
rect 848 656 850 698
rect 871 697 875 698
rect 903 702 907 703
rect 903 697 907 698
rect 943 702 947 703
rect 943 697 947 698
rect 967 702 971 703
rect 967 697 971 698
rect 1015 702 1019 703
rect 1015 697 1019 698
rect 1031 702 1035 703
rect 1050 699 1051 703
rect 1055 699 1056 703
rect 1050 698 1056 699
rect 1087 702 1091 703
rect 1031 697 1035 698
rect 1087 697 1091 698
rect 1135 702 1139 703
rect 1135 697 1139 698
rect 1151 702 1155 703
rect 1151 697 1155 698
rect 1175 702 1179 703
rect 1175 697 1179 698
rect 1215 702 1219 703
rect 1215 697 1219 698
rect 1247 702 1251 703
rect 1247 697 1251 698
rect 1271 702 1275 703
rect 1271 697 1275 698
rect 1279 702 1283 703
rect 1279 697 1283 698
rect 904 695 906 697
rect 968 695 970 697
rect 1032 695 1034 697
rect 1088 695 1090 697
rect 1136 695 1138 697
rect 1176 695 1178 697
rect 1216 695 1218 697
rect 1248 695 1250 697
rect 1280 695 1282 697
rect 1292 696 1294 722
rect 1376 712 1378 742
rect 1383 737 1387 738
rect 1415 742 1419 743
rect 1415 737 1419 738
rect 1447 742 1451 743
rect 1447 737 1451 738
rect 1382 736 1388 737
rect 1382 732 1383 736
rect 1387 732 1388 736
rect 1382 731 1388 732
rect 1414 736 1420 737
rect 1414 732 1415 736
rect 1419 732 1420 736
rect 1448 734 1450 737
rect 1414 731 1420 732
rect 1446 733 1452 734
rect 1446 729 1447 733
rect 1451 729 1452 733
rect 1446 728 1452 729
rect 1426 719 1432 720
rect 1426 715 1427 719
rect 1431 715 1432 719
rect 1426 714 1432 715
rect 1446 715 1452 716
rect 1374 711 1380 712
rect 1326 710 1332 711
rect 1326 706 1327 710
rect 1331 706 1332 710
rect 1374 707 1375 711
rect 1379 707 1380 711
rect 1374 706 1380 707
rect 1382 710 1388 711
rect 1382 706 1383 710
rect 1387 706 1388 710
rect 1326 705 1332 706
rect 1382 705 1388 706
rect 1414 710 1420 711
rect 1414 706 1415 710
rect 1419 706 1420 710
rect 1414 705 1420 706
rect 1328 703 1330 705
rect 1384 703 1386 705
rect 1416 703 1418 705
rect 1311 702 1315 703
rect 1311 697 1315 698
rect 1327 702 1331 703
rect 1327 697 1331 698
rect 1343 702 1347 703
rect 1343 697 1347 698
rect 1367 702 1371 703
rect 1367 697 1371 698
rect 1383 702 1387 703
rect 1383 697 1387 698
rect 1391 702 1395 703
rect 1391 697 1395 698
rect 1415 702 1419 703
rect 1415 697 1419 698
rect 1290 695 1296 696
rect 1312 695 1314 697
rect 1344 695 1346 697
rect 1368 695 1370 697
rect 1392 695 1394 697
rect 1416 695 1418 697
rect 1428 696 1430 714
rect 1446 711 1447 715
rect 1451 711 1452 715
rect 1446 710 1452 711
rect 1448 703 1450 710
rect 1447 702 1451 703
rect 1447 697 1451 698
rect 1426 695 1432 696
rect 902 694 908 695
rect 902 690 903 694
rect 907 690 908 694
rect 902 689 908 690
rect 966 694 972 695
rect 966 690 967 694
rect 971 690 972 694
rect 966 689 972 690
rect 1030 694 1036 695
rect 1030 690 1031 694
rect 1035 690 1036 694
rect 1030 689 1036 690
rect 1086 694 1092 695
rect 1086 690 1087 694
rect 1091 690 1092 694
rect 1086 689 1092 690
rect 1134 694 1140 695
rect 1134 690 1135 694
rect 1139 690 1140 694
rect 1134 689 1140 690
rect 1174 694 1180 695
rect 1174 690 1175 694
rect 1179 690 1180 694
rect 1174 689 1180 690
rect 1214 694 1220 695
rect 1214 690 1215 694
rect 1219 690 1220 694
rect 1214 689 1220 690
rect 1246 694 1252 695
rect 1246 690 1247 694
rect 1251 690 1252 694
rect 1246 689 1252 690
rect 1278 694 1284 695
rect 1278 690 1279 694
rect 1283 690 1284 694
rect 1290 691 1291 695
rect 1295 691 1296 695
rect 1290 690 1296 691
rect 1310 694 1316 695
rect 1310 690 1311 694
rect 1315 690 1316 694
rect 1278 689 1284 690
rect 1310 689 1316 690
rect 1342 694 1348 695
rect 1342 690 1343 694
rect 1347 690 1348 694
rect 1366 694 1372 695
rect 1342 689 1348 690
rect 1354 691 1360 692
rect 1354 687 1355 691
rect 1359 687 1360 691
rect 1366 690 1367 694
rect 1371 690 1372 694
rect 1366 689 1372 690
rect 1390 694 1396 695
rect 1390 690 1391 694
rect 1395 690 1396 694
rect 1390 689 1396 690
rect 1414 694 1420 695
rect 1414 690 1415 694
rect 1419 690 1420 694
rect 1426 691 1427 695
rect 1431 691 1432 695
rect 1426 690 1432 691
rect 1448 690 1450 697
rect 1414 689 1420 690
rect 1446 689 1452 690
rect 1354 686 1360 687
rect 902 668 908 669
rect 902 664 903 668
rect 907 664 908 668
rect 902 663 908 664
rect 966 668 972 669
rect 966 664 967 668
rect 971 664 972 668
rect 966 663 972 664
rect 1030 668 1036 669
rect 1086 668 1092 669
rect 1030 664 1031 668
rect 1035 664 1036 668
rect 1030 663 1036 664
rect 1078 667 1084 668
rect 1078 663 1079 667
rect 1083 663 1084 667
rect 1086 664 1087 668
rect 1091 664 1092 668
rect 1086 663 1092 664
rect 1134 668 1140 669
rect 1134 664 1135 668
rect 1139 664 1140 668
rect 1134 663 1140 664
rect 1174 668 1180 669
rect 1174 664 1175 668
rect 1179 664 1180 668
rect 1174 663 1180 664
rect 1214 668 1220 669
rect 1214 664 1215 668
rect 1219 664 1220 668
rect 1214 663 1220 664
rect 1246 668 1252 669
rect 1246 664 1247 668
rect 1251 664 1252 668
rect 1246 663 1252 664
rect 1278 668 1284 669
rect 1278 664 1279 668
rect 1283 664 1284 668
rect 1278 663 1284 664
rect 1310 668 1316 669
rect 1310 664 1311 668
rect 1315 664 1316 668
rect 1310 663 1316 664
rect 1342 668 1348 669
rect 1342 664 1343 668
rect 1347 664 1348 668
rect 1342 663 1348 664
rect 863 662 867 663
rect 863 657 867 658
rect 903 662 907 663
rect 903 657 907 658
rect 935 662 939 663
rect 935 657 939 658
rect 967 662 971 663
rect 967 657 971 658
rect 1007 662 1011 663
rect 1007 657 1011 658
rect 1031 662 1035 663
rect 1031 657 1035 658
rect 1047 662 1051 663
rect 1078 662 1084 663
rect 1087 662 1091 663
rect 1047 657 1051 658
rect 862 656 868 657
rect 814 652 815 656
rect 819 652 820 656
rect 814 651 820 652
rect 846 655 852 656
rect 846 651 847 655
rect 851 651 852 655
rect 862 652 863 656
rect 867 652 868 656
rect 862 651 868 652
rect 902 656 908 657
rect 902 652 903 656
rect 907 652 908 656
rect 902 651 908 652
rect 934 656 940 657
rect 934 652 935 656
rect 939 652 940 656
rect 934 651 940 652
rect 966 656 972 657
rect 966 652 967 656
rect 971 652 972 656
rect 966 651 972 652
rect 1006 656 1012 657
rect 1006 652 1007 656
rect 1011 652 1012 656
rect 1006 651 1012 652
rect 1046 656 1052 657
rect 1046 652 1047 656
rect 1051 652 1052 656
rect 1046 651 1052 652
rect 846 650 852 651
rect 1080 648 1082 662
rect 1087 657 1091 658
rect 1127 662 1131 663
rect 1127 657 1131 658
rect 1135 662 1139 663
rect 1135 657 1139 658
rect 1159 662 1163 663
rect 1159 657 1163 658
rect 1175 662 1179 663
rect 1175 657 1179 658
rect 1191 662 1195 663
rect 1191 657 1195 658
rect 1215 662 1219 663
rect 1215 657 1219 658
rect 1223 662 1227 663
rect 1223 657 1227 658
rect 1247 662 1251 663
rect 1247 657 1251 658
rect 1263 662 1267 663
rect 1263 657 1267 658
rect 1279 662 1283 663
rect 1279 657 1283 658
rect 1303 662 1307 663
rect 1303 657 1307 658
rect 1311 662 1315 663
rect 1311 657 1315 658
rect 1343 662 1347 663
rect 1356 660 1358 686
rect 1446 685 1447 689
rect 1451 685 1452 689
rect 1446 684 1452 685
rect 1446 671 1452 672
rect 1366 668 1372 669
rect 1366 664 1367 668
rect 1371 664 1372 668
rect 1366 663 1372 664
rect 1390 668 1396 669
rect 1390 664 1391 668
rect 1395 664 1396 668
rect 1390 663 1396 664
rect 1414 668 1420 669
rect 1414 664 1415 668
rect 1419 664 1420 668
rect 1446 667 1447 671
rect 1451 667 1452 671
rect 1446 666 1452 667
rect 1414 663 1420 664
rect 1448 663 1450 666
rect 1367 662 1371 663
rect 1343 657 1347 658
rect 1354 659 1360 660
rect 1086 656 1092 657
rect 1086 652 1087 656
rect 1091 652 1092 656
rect 1086 651 1092 652
rect 1126 656 1132 657
rect 1126 652 1127 656
rect 1131 652 1132 656
rect 1126 651 1132 652
rect 1158 656 1164 657
rect 1158 652 1159 656
rect 1163 652 1164 656
rect 1158 651 1164 652
rect 1190 656 1196 657
rect 1190 652 1191 656
rect 1195 652 1196 656
rect 1190 651 1196 652
rect 1222 656 1228 657
rect 1222 652 1223 656
rect 1227 652 1228 656
rect 1222 651 1228 652
rect 1262 656 1268 657
rect 1262 652 1263 656
rect 1267 652 1268 656
rect 1262 651 1268 652
rect 1302 656 1308 657
rect 1302 652 1303 656
rect 1307 652 1308 656
rect 1302 651 1308 652
rect 1342 656 1348 657
rect 1342 652 1343 656
rect 1347 652 1348 656
rect 1354 655 1355 659
rect 1359 655 1360 659
rect 1367 657 1371 658
rect 1391 662 1395 663
rect 1391 657 1395 658
rect 1415 662 1419 663
rect 1415 657 1419 658
rect 1447 662 1451 663
rect 1447 657 1451 658
rect 1354 654 1360 655
rect 1448 654 1450 657
rect 1342 651 1348 652
rect 1446 653 1452 654
rect 1446 649 1447 653
rect 1451 649 1452 653
rect 1446 648 1452 649
rect 674 647 680 648
rect 674 643 675 647
rect 679 643 680 647
rect 674 642 680 643
rect 986 647 992 648
rect 986 643 987 647
rect 991 643 992 647
rect 986 642 992 643
rect 1078 647 1084 648
rect 1078 643 1079 647
rect 1083 643 1084 647
rect 1078 642 1084 643
rect 1170 647 1176 648
rect 1170 643 1171 647
rect 1175 643 1176 647
rect 1170 642 1176 643
rect 1234 647 1240 648
rect 1234 643 1235 647
rect 1239 643 1240 647
rect 1234 642 1240 643
rect 1314 647 1320 648
rect 1314 643 1315 647
rect 1319 643 1320 647
rect 1314 642 1320 643
rect 1322 647 1328 648
rect 1322 643 1323 647
rect 1327 643 1328 647
rect 1322 642 1328 643
rect 676 632 678 642
rect 710 639 716 640
rect 710 635 711 639
rect 715 635 716 639
rect 710 634 716 635
rect 202 631 208 632
rect 226 631 232 632
rect 274 631 280 632
rect 338 631 344 632
rect 347 631 351 632
rect 446 631 452 632
rect 466 631 472 632
rect 531 631 535 632
rect 562 631 568 632
rect 650 631 656 632
rect 674 631 680 632
rect 110 630 116 631
rect 190 630 196 631
rect 112 623 114 630
rect 190 626 191 630
rect 195 626 196 630
rect 202 627 203 631
rect 207 627 208 631
rect 202 626 208 627
rect 214 630 220 631
rect 214 626 215 630
rect 219 626 220 630
rect 226 627 227 631
rect 231 627 232 631
rect 226 626 232 627
rect 238 630 244 631
rect 238 626 239 630
rect 243 626 244 630
rect 190 625 196 626
rect 214 625 220 626
rect 238 625 244 626
rect 262 630 268 631
rect 262 626 263 630
rect 267 626 268 630
rect 274 627 275 631
rect 279 627 280 631
rect 274 626 280 627
rect 294 630 300 631
rect 294 626 295 630
rect 299 626 300 630
rect 262 625 268 626
rect 294 625 300 626
rect 326 630 332 631
rect 326 626 327 630
rect 331 626 332 630
rect 338 627 339 631
rect 343 627 344 631
rect 338 626 344 627
rect 366 630 372 631
rect 366 626 367 630
rect 371 626 372 630
rect 326 625 332 626
rect 366 625 372 626
rect 406 630 412 631
rect 406 626 407 630
rect 411 626 412 630
rect 446 627 447 631
rect 451 627 452 631
rect 446 626 452 627
rect 454 630 460 631
rect 454 626 455 630
rect 459 626 460 630
rect 466 627 467 631
rect 471 627 472 631
rect 466 626 472 627
rect 502 630 508 631
rect 502 626 503 630
rect 507 626 508 630
rect 406 625 412 626
rect 454 625 460 626
rect 502 625 508 626
rect 192 623 194 625
rect 216 623 218 625
rect 240 623 242 625
rect 264 623 266 625
rect 296 623 298 625
rect 328 623 330 625
rect 368 623 370 625
rect 408 623 410 625
rect 456 623 458 625
rect 504 623 506 625
rect 111 622 115 623
rect 111 617 115 618
rect 191 622 195 623
rect 191 617 195 618
rect 215 622 219 623
rect 215 617 219 618
rect 239 622 243 623
rect 239 617 243 618
rect 263 622 267 623
rect 263 617 267 618
rect 271 622 275 623
rect 271 617 275 618
rect 295 622 299 623
rect 295 617 299 618
rect 319 622 323 623
rect 319 617 323 618
rect 327 622 331 623
rect 327 617 331 618
rect 343 622 347 623
rect 343 617 347 618
rect 367 622 371 623
rect 367 617 371 618
rect 391 622 395 623
rect 391 617 395 618
rect 407 622 411 623
rect 407 617 411 618
rect 415 622 419 623
rect 439 622 443 623
rect 415 617 419 618
rect 422 619 428 620
rect 112 610 114 617
rect 272 615 274 617
rect 296 615 298 617
rect 320 615 322 617
rect 344 615 346 617
rect 368 615 370 617
rect 392 615 394 617
rect 416 615 418 617
rect 422 615 423 619
rect 427 615 428 619
rect 439 617 443 618
rect 455 622 459 623
rect 455 617 459 618
rect 479 622 483 623
rect 479 617 483 618
rect 503 622 507 623
rect 503 617 507 618
rect 519 622 523 623
rect 519 617 523 618
rect 440 615 442 617
rect 480 615 482 617
rect 520 615 522 617
rect 270 614 276 615
rect 270 610 271 614
rect 275 610 276 614
rect 110 609 116 610
rect 270 609 276 610
rect 294 614 300 615
rect 294 610 295 614
rect 299 610 300 614
rect 318 614 324 615
rect 294 609 300 610
rect 306 611 312 612
rect 110 605 111 609
rect 115 605 116 609
rect 306 607 307 611
rect 311 607 312 611
rect 318 610 319 614
rect 323 610 324 614
rect 318 609 324 610
rect 342 614 348 615
rect 342 610 343 614
rect 347 610 348 614
rect 342 609 348 610
rect 366 614 372 615
rect 366 610 367 614
rect 371 610 372 614
rect 366 609 372 610
rect 390 614 396 615
rect 390 610 391 614
rect 395 610 396 614
rect 414 614 420 615
rect 422 614 428 615
rect 438 614 444 615
rect 402 611 408 612
rect 402 610 403 611
rect 390 609 396 610
rect 306 606 312 607
rect 400 607 403 610
rect 407 607 408 611
rect 414 610 415 614
rect 419 610 420 614
rect 414 609 420 610
rect 400 606 408 607
rect 110 604 116 605
rect 294 603 300 604
rect 308 603 310 606
rect 294 599 295 603
rect 299 601 310 603
rect 400 602 402 606
rect 299 599 300 601
rect 392 600 402 602
rect 424 602 426 614
rect 438 610 439 614
rect 443 610 444 614
rect 438 609 444 610
rect 478 614 484 615
rect 478 610 479 614
rect 483 610 484 614
rect 478 609 484 610
rect 518 614 524 615
rect 518 610 519 614
rect 523 610 524 614
rect 518 609 524 610
rect 424 600 450 602
rect 294 598 300 599
rect 390 599 396 600
rect 390 595 391 599
rect 395 595 396 599
rect 390 594 396 595
rect 414 599 420 600
rect 414 595 415 599
rect 419 598 420 599
rect 419 596 426 598
rect 419 595 420 596
rect 414 594 420 595
rect 110 591 116 592
rect 110 587 111 591
rect 115 587 116 591
rect 110 586 116 587
rect 270 588 276 589
rect 112 583 114 586
rect 270 584 271 588
rect 275 584 276 588
rect 270 583 276 584
rect 294 588 300 589
rect 294 584 295 588
rect 299 584 300 588
rect 294 583 300 584
rect 318 588 324 589
rect 318 584 319 588
rect 323 584 324 588
rect 318 583 324 584
rect 342 588 348 589
rect 342 584 343 588
rect 347 584 348 588
rect 342 583 348 584
rect 366 588 372 589
rect 366 584 367 588
rect 371 584 372 588
rect 366 583 372 584
rect 390 588 396 589
rect 390 584 391 588
rect 395 584 396 588
rect 390 583 396 584
rect 414 588 420 589
rect 414 584 415 588
rect 419 584 420 588
rect 414 583 420 584
rect 111 582 115 583
rect 111 577 115 578
rect 263 582 267 583
rect 263 577 267 578
rect 271 582 275 583
rect 271 577 275 578
rect 287 582 291 583
rect 287 577 291 578
rect 295 582 299 583
rect 295 577 299 578
rect 311 582 315 583
rect 311 577 315 578
rect 319 582 323 583
rect 319 577 323 578
rect 335 582 339 583
rect 335 577 339 578
rect 343 582 347 583
rect 343 577 347 578
rect 359 582 363 583
rect 359 577 363 578
rect 367 582 371 583
rect 367 577 371 578
rect 383 582 387 583
rect 383 577 387 578
rect 391 582 395 583
rect 391 577 395 578
rect 407 582 411 583
rect 407 577 411 578
rect 415 582 419 583
rect 415 577 419 578
rect 112 574 114 577
rect 262 576 268 577
rect 110 573 116 574
rect 110 569 111 573
rect 115 569 116 573
rect 262 572 263 576
rect 267 572 268 576
rect 262 571 268 572
rect 286 576 292 577
rect 286 572 287 576
rect 291 572 292 576
rect 286 571 292 572
rect 310 576 316 577
rect 310 572 311 576
rect 315 572 316 576
rect 310 571 316 572
rect 334 576 340 577
rect 334 572 335 576
rect 339 572 340 576
rect 334 571 340 572
rect 358 576 364 577
rect 358 572 359 576
rect 363 572 364 576
rect 358 571 364 572
rect 382 576 388 577
rect 382 572 383 576
rect 387 572 388 576
rect 382 571 388 572
rect 406 576 412 577
rect 406 572 407 576
rect 411 572 412 576
rect 406 571 412 572
rect 110 568 116 569
rect 398 567 404 568
rect 398 563 399 567
rect 403 563 404 567
rect 398 562 404 563
rect 110 555 116 556
rect 110 551 111 555
rect 115 551 116 555
rect 110 550 116 551
rect 262 550 268 551
rect 112 543 114 550
rect 262 546 263 550
rect 267 546 268 550
rect 262 545 268 546
rect 286 550 292 551
rect 286 546 287 550
rect 291 546 292 550
rect 286 545 292 546
rect 310 550 316 551
rect 310 546 311 550
rect 315 546 316 550
rect 310 545 316 546
rect 334 550 340 551
rect 334 546 335 550
rect 339 546 340 550
rect 334 545 340 546
rect 358 550 364 551
rect 358 546 359 550
rect 363 546 364 550
rect 358 545 364 546
rect 382 550 388 551
rect 382 546 383 550
rect 387 546 388 550
rect 382 545 388 546
rect 264 543 266 545
rect 288 543 290 545
rect 312 543 314 545
rect 336 543 338 545
rect 360 543 362 545
rect 384 543 386 545
rect 111 542 115 543
rect 111 537 115 538
rect 223 542 227 543
rect 223 537 227 538
rect 247 542 251 543
rect 247 537 251 538
rect 263 542 267 543
rect 263 537 267 538
rect 271 542 275 543
rect 271 537 275 538
rect 287 542 291 543
rect 287 537 291 538
rect 295 542 299 543
rect 295 537 299 538
rect 311 542 315 543
rect 311 537 315 538
rect 327 542 331 543
rect 327 537 331 538
rect 335 542 339 543
rect 335 537 339 538
rect 359 542 363 543
rect 359 537 363 538
rect 383 542 387 543
rect 383 537 387 538
rect 391 542 395 543
rect 400 540 402 562
rect 415 551 421 552
rect 406 550 412 551
rect 406 546 407 550
rect 411 546 412 550
rect 415 547 416 551
rect 420 550 421 551
rect 424 550 426 596
rect 438 588 444 589
rect 438 584 439 588
rect 443 584 444 588
rect 438 583 444 584
rect 431 582 435 583
rect 431 577 435 578
rect 439 582 443 583
rect 439 577 443 578
rect 430 576 436 577
rect 430 572 431 576
rect 435 572 436 576
rect 430 571 436 572
rect 439 571 445 572
rect 439 567 440 571
rect 444 570 445 571
rect 448 570 450 600
rect 532 592 534 631
rect 550 630 556 631
rect 550 626 551 630
rect 555 626 556 630
rect 562 627 563 631
rect 567 627 568 631
rect 562 626 568 627
rect 606 630 612 631
rect 606 626 607 630
rect 611 626 612 630
rect 650 627 651 631
rect 655 627 656 631
rect 650 626 656 627
rect 662 630 668 631
rect 662 626 663 630
rect 667 626 668 630
rect 674 627 675 631
rect 679 627 680 631
rect 674 626 680 627
rect 550 625 556 626
rect 606 625 612 626
rect 662 625 668 626
rect 552 623 554 625
rect 608 623 610 625
rect 664 623 666 625
rect 551 622 555 623
rect 551 617 555 618
rect 567 622 571 623
rect 567 617 571 618
rect 607 622 611 623
rect 607 617 611 618
rect 623 622 627 623
rect 623 617 627 618
rect 663 622 667 623
rect 663 617 667 618
rect 679 622 683 623
rect 679 617 683 618
rect 568 615 570 617
rect 624 615 626 617
rect 680 615 682 617
rect 712 616 714 634
rect 718 630 724 631
rect 718 626 719 630
rect 723 626 724 630
rect 718 625 724 626
rect 766 630 772 631
rect 766 626 767 630
rect 771 626 772 630
rect 766 625 772 626
rect 814 630 820 631
rect 814 626 815 630
rect 819 626 820 630
rect 814 625 820 626
rect 862 630 868 631
rect 862 626 863 630
rect 867 626 868 630
rect 862 625 868 626
rect 902 630 908 631
rect 902 626 903 630
rect 907 626 908 630
rect 902 625 908 626
rect 934 630 940 631
rect 934 626 935 630
rect 939 626 940 630
rect 934 625 940 626
rect 966 630 972 631
rect 966 626 967 630
rect 971 626 972 630
rect 966 625 972 626
rect 720 623 722 625
rect 768 623 770 625
rect 774 623 780 624
rect 816 623 818 625
rect 864 623 866 625
rect 904 623 906 625
rect 936 623 938 625
rect 968 623 970 625
rect 719 622 723 623
rect 719 617 723 618
rect 735 622 739 623
rect 735 617 739 618
rect 767 622 771 623
rect 774 619 775 623
rect 779 619 780 623
rect 774 618 780 619
rect 783 622 787 623
rect 767 617 771 618
rect 710 615 716 616
rect 736 615 738 617
rect 566 614 572 615
rect 566 610 567 614
rect 571 610 572 614
rect 566 609 572 610
rect 622 614 628 615
rect 622 610 623 614
rect 627 610 628 614
rect 622 609 628 610
rect 678 614 684 615
rect 678 610 679 614
rect 683 610 684 614
rect 710 611 711 615
rect 715 611 716 615
rect 710 610 716 611
rect 734 614 740 615
rect 734 610 735 614
rect 739 610 740 614
rect 678 609 684 610
rect 734 609 740 610
rect 776 604 778 618
rect 783 617 787 618
rect 815 622 819 623
rect 815 617 819 618
rect 831 622 835 623
rect 831 617 835 618
rect 863 622 867 623
rect 863 617 867 618
rect 879 622 883 623
rect 879 617 883 618
rect 903 622 907 623
rect 903 617 907 618
rect 927 622 931 623
rect 927 617 931 618
rect 935 622 939 623
rect 935 617 939 618
rect 967 622 971 623
rect 967 617 971 618
rect 975 622 979 623
rect 975 617 979 618
rect 784 615 786 617
rect 832 615 834 617
rect 880 615 882 617
rect 928 615 930 617
rect 976 615 978 617
rect 988 616 990 642
rect 1172 632 1174 642
rect 1236 632 1238 642
rect 1316 632 1318 642
rect 1170 631 1176 632
rect 1234 631 1240 632
rect 1314 631 1320 632
rect 1006 630 1012 631
rect 1006 626 1007 630
rect 1011 626 1012 630
rect 1006 625 1012 626
rect 1046 630 1052 631
rect 1046 626 1047 630
rect 1051 626 1052 630
rect 1046 625 1052 626
rect 1086 630 1092 631
rect 1086 626 1087 630
rect 1091 626 1092 630
rect 1086 625 1092 626
rect 1126 630 1132 631
rect 1126 626 1127 630
rect 1131 626 1132 630
rect 1126 625 1132 626
rect 1158 630 1164 631
rect 1158 626 1159 630
rect 1163 626 1164 630
rect 1170 627 1171 631
rect 1175 627 1176 631
rect 1170 626 1176 627
rect 1190 630 1196 631
rect 1190 626 1191 630
rect 1195 626 1196 630
rect 1158 625 1164 626
rect 1190 625 1196 626
rect 1222 630 1228 631
rect 1222 626 1223 630
rect 1227 626 1228 630
rect 1234 627 1235 631
rect 1239 627 1240 631
rect 1234 626 1240 627
rect 1262 630 1268 631
rect 1262 626 1263 630
rect 1267 626 1268 630
rect 1222 625 1228 626
rect 1262 625 1268 626
rect 1302 630 1308 631
rect 1302 626 1303 630
rect 1307 626 1308 630
rect 1314 627 1315 631
rect 1319 627 1320 631
rect 1314 626 1320 627
rect 1302 625 1308 626
rect 1008 623 1010 625
rect 1034 623 1040 624
rect 1048 623 1050 625
rect 1088 623 1090 625
rect 1128 623 1130 625
rect 1160 623 1162 625
rect 1192 623 1194 625
rect 1224 623 1226 625
rect 1264 623 1266 625
rect 1304 623 1306 625
rect 1324 624 1326 642
rect 1446 635 1452 636
rect 1446 631 1447 635
rect 1451 631 1452 635
rect 1342 630 1348 631
rect 1446 630 1452 631
rect 1342 626 1343 630
rect 1347 626 1348 630
rect 1342 625 1348 626
rect 1322 623 1328 624
rect 1344 623 1346 625
rect 1448 623 1450 630
rect 1007 622 1011 623
rect 1007 617 1011 618
rect 1023 622 1027 623
rect 1034 619 1035 623
rect 1039 619 1040 623
rect 1034 618 1040 619
rect 1047 622 1051 623
rect 1023 617 1027 618
rect 986 615 992 616
rect 1024 615 1026 617
rect 782 614 788 615
rect 782 610 783 614
rect 787 610 788 614
rect 830 614 836 615
rect 782 609 788 610
rect 794 611 800 612
rect 794 607 795 611
rect 799 607 800 611
rect 830 610 831 614
rect 835 610 836 614
rect 830 609 836 610
rect 878 614 884 615
rect 878 610 879 614
rect 883 610 884 614
rect 878 609 884 610
rect 926 614 932 615
rect 926 610 927 614
rect 931 610 932 614
rect 926 609 932 610
rect 974 614 980 615
rect 974 610 975 614
rect 979 610 980 614
rect 986 611 987 615
rect 991 611 992 615
rect 986 610 992 611
rect 1022 614 1028 615
rect 1022 610 1023 614
rect 1027 610 1028 614
rect 974 609 980 610
rect 1022 609 1028 610
rect 794 606 800 607
rect 774 603 780 604
rect 774 599 775 603
rect 779 599 780 603
rect 774 598 780 599
rect 530 591 536 592
rect 478 588 484 589
rect 478 584 479 588
rect 483 584 484 588
rect 478 583 484 584
rect 518 588 524 589
rect 518 584 519 588
rect 523 584 524 588
rect 530 587 531 591
rect 535 587 536 591
rect 530 586 536 587
rect 566 588 572 589
rect 622 588 628 589
rect 518 583 524 584
rect 566 584 567 588
rect 571 584 572 588
rect 566 583 572 584
rect 614 587 620 588
rect 614 583 615 587
rect 619 583 620 587
rect 622 584 623 588
rect 627 584 628 588
rect 622 583 628 584
rect 678 588 684 589
rect 678 584 679 588
rect 683 584 684 588
rect 678 583 684 584
rect 734 588 740 589
rect 734 584 735 588
rect 739 584 740 588
rect 734 583 740 584
rect 782 588 788 589
rect 782 584 783 588
rect 787 584 788 588
rect 782 583 788 584
rect 463 582 467 583
rect 463 577 467 578
rect 479 582 483 583
rect 479 577 483 578
rect 503 582 507 583
rect 503 577 507 578
rect 519 582 523 583
rect 519 577 523 578
rect 551 582 555 583
rect 551 577 555 578
rect 567 582 571 583
rect 567 577 571 578
rect 607 582 611 583
rect 614 582 620 583
rect 623 582 627 583
rect 607 577 611 578
rect 462 576 468 577
rect 462 572 463 576
rect 467 572 468 576
rect 462 571 468 572
rect 502 576 508 577
rect 502 572 503 576
rect 507 572 508 576
rect 502 571 508 572
rect 550 576 556 577
rect 550 572 551 576
rect 555 572 556 576
rect 550 571 556 572
rect 606 576 612 577
rect 606 572 607 576
rect 611 572 612 576
rect 606 571 612 572
rect 444 568 450 570
rect 444 567 445 568
rect 439 566 445 567
rect 616 563 618 582
rect 623 577 627 578
rect 663 582 667 583
rect 663 577 667 578
rect 679 582 683 583
rect 679 577 683 578
rect 719 582 723 583
rect 719 577 723 578
rect 735 582 739 583
rect 735 577 739 578
rect 775 582 779 583
rect 775 577 779 578
rect 783 582 787 583
rect 783 577 787 578
rect 662 576 668 577
rect 662 572 663 576
rect 667 572 668 576
rect 662 571 668 572
rect 718 576 724 577
rect 718 572 719 576
rect 723 572 724 576
rect 718 571 724 572
rect 774 576 780 577
rect 796 576 798 606
rect 1036 604 1038 618
rect 1047 617 1051 618
rect 1071 622 1075 623
rect 1071 617 1075 618
rect 1087 622 1091 623
rect 1087 617 1091 618
rect 1111 622 1115 623
rect 1111 617 1115 618
rect 1127 622 1131 623
rect 1127 617 1131 618
rect 1151 622 1155 623
rect 1151 617 1155 618
rect 1159 622 1163 623
rect 1159 617 1163 618
rect 1191 622 1195 623
rect 1191 617 1195 618
rect 1223 622 1227 623
rect 1223 617 1227 618
rect 1239 622 1243 623
rect 1239 617 1243 618
rect 1263 622 1267 623
rect 1263 617 1267 618
rect 1287 622 1291 623
rect 1287 617 1291 618
rect 1303 622 1307 623
rect 1322 619 1323 623
rect 1327 619 1328 623
rect 1322 618 1328 619
rect 1335 622 1339 623
rect 1303 617 1307 618
rect 1335 617 1339 618
rect 1343 622 1347 623
rect 1343 617 1347 618
rect 1447 622 1451 623
rect 1447 617 1451 618
rect 1072 615 1074 617
rect 1112 615 1114 617
rect 1152 615 1154 617
rect 1192 615 1194 617
rect 1240 615 1242 617
rect 1288 615 1290 617
rect 1336 615 1338 617
rect 1070 614 1076 615
rect 1070 610 1071 614
rect 1075 610 1076 614
rect 1070 609 1076 610
rect 1110 614 1116 615
rect 1110 610 1111 614
rect 1115 610 1116 614
rect 1110 609 1116 610
rect 1150 614 1156 615
rect 1150 610 1151 614
rect 1155 610 1156 614
rect 1150 609 1156 610
rect 1190 614 1196 615
rect 1190 610 1191 614
rect 1195 610 1196 614
rect 1190 609 1196 610
rect 1238 614 1244 615
rect 1238 610 1239 614
rect 1243 610 1244 614
rect 1238 609 1244 610
rect 1286 614 1292 615
rect 1286 610 1287 614
rect 1291 610 1292 614
rect 1286 609 1292 610
rect 1334 614 1340 615
rect 1334 610 1335 614
rect 1339 610 1340 614
rect 1448 610 1450 617
rect 1334 609 1340 610
rect 1446 609 1452 610
rect 1446 605 1447 609
rect 1451 605 1452 609
rect 1446 604 1452 605
rect 1034 603 1040 604
rect 1034 599 1035 603
rect 1039 599 1040 603
rect 1034 598 1040 599
rect 1446 591 1452 592
rect 830 588 836 589
rect 878 588 884 589
rect 830 584 831 588
rect 835 584 836 588
rect 830 583 836 584
rect 870 587 876 588
rect 870 583 871 587
rect 875 583 876 587
rect 878 584 879 588
rect 883 584 884 588
rect 878 583 884 584
rect 926 588 932 589
rect 926 584 927 588
rect 931 584 932 588
rect 926 583 932 584
rect 974 588 980 589
rect 974 584 975 588
rect 979 584 980 588
rect 974 583 980 584
rect 1022 588 1028 589
rect 1022 584 1023 588
rect 1027 584 1028 588
rect 1022 583 1028 584
rect 1070 588 1076 589
rect 1070 584 1071 588
rect 1075 584 1076 588
rect 1070 583 1076 584
rect 1110 588 1116 589
rect 1110 584 1111 588
rect 1115 584 1116 588
rect 1110 583 1116 584
rect 1150 588 1156 589
rect 1150 584 1151 588
rect 1155 584 1156 588
rect 1150 583 1156 584
rect 1190 588 1196 589
rect 1190 584 1191 588
rect 1195 584 1196 588
rect 1190 583 1196 584
rect 1238 588 1244 589
rect 1238 584 1239 588
rect 1243 584 1244 588
rect 1238 583 1244 584
rect 1286 588 1292 589
rect 1286 584 1287 588
rect 1291 584 1292 588
rect 1286 583 1292 584
rect 1334 588 1340 589
rect 1334 584 1335 588
rect 1339 584 1340 588
rect 1334 583 1340 584
rect 1386 587 1392 588
rect 1386 583 1387 587
rect 1391 583 1392 587
rect 1446 587 1447 591
rect 1451 587 1452 591
rect 1446 586 1452 587
rect 1448 583 1450 586
rect 831 582 835 583
rect 870 582 876 583
rect 879 582 883 583
rect 831 577 835 578
rect 830 576 836 577
rect 774 572 775 576
rect 779 572 780 576
rect 774 571 780 572
rect 794 575 800 576
rect 794 571 795 575
rect 799 571 800 575
rect 830 572 831 576
rect 835 572 836 576
rect 830 571 836 572
rect 794 570 800 571
rect 674 567 680 568
rect 674 563 675 567
rect 679 563 680 567
rect 616 561 622 563
rect 674 562 680 563
rect 538 559 544 560
rect 538 555 539 559
rect 543 555 544 559
rect 538 554 544 555
rect 420 548 426 550
rect 430 550 436 551
rect 420 547 421 548
rect 415 546 421 547
rect 430 546 431 550
rect 435 546 436 550
rect 406 545 412 546
rect 430 545 436 546
rect 462 550 468 551
rect 462 546 463 550
rect 467 546 468 550
rect 462 545 468 546
rect 502 550 508 551
rect 502 546 503 550
rect 507 546 508 550
rect 502 545 508 546
rect 514 547 520 548
rect 408 543 410 545
rect 432 543 434 545
rect 464 543 466 545
rect 504 543 506 545
rect 514 543 515 547
rect 519 543 520 547
rect 407 542 411 543
rect 391 537 395 538
rect 398 539 404 540
rect 112 530 114 537
rect 224 535 226 537
rect 248 535 250 537
rect 272 535 274 537
rect 296 535 298 537
rect 328 535 330 537
rect 360 535 362 537
rect 392 535 394 537
rect 398 535 399 539
rect 403 535 404 539
rect 407 537 411 538
rect 423 542 427 543
rect 423 537 427 538
rect 431 542 435 543
rect 431 537 435 538
rect 455 542 459 543
rect 455 537 459 538
rect 463 542 467 543
rect 463 537 467 538
rect 487 542 491 543
rect 487 537 491 538
rect 503 542 507 543
rect 514 542 520 543
rect 527 542 531 543
rect 503 537 507 538
rect 424 535 426 537
rect 456 535 458 537
rect 488 535 490 537
rect 222 534 228 535
rect 222 530 223 534
rect 227 530 228 534
rect 246 534 252 535
rect 110 529 116 530
rect 222 529 228 530
rect 234 531 240 532
rect 110 525 111 529
rect 115 525 116 529
rect 234 527 235 531
rect 239 527 240 531
rect 246 530 247 534
rect 251 530 252 534
rect 246 529 252 530
rect 270 534 276 535
rect 270 530 271 534
rect 275 530 276 534
rect 270 529 276 530
rect 294 534 300 535
rect 294 530 295 534
rect 299 530 300 534
rect 294 529 300 530
rect 326 534 332 535
rect 326 530 327 534
rect 331 530 332 534
rect 326 529 332 530
rect 358 534 364 535
rect 358 530 359 534
rect 363 530 364 534
rect 358 529 364 530
rect 390 534 396 535
rect 398 534 404 535
rect 422 534 428 535
rect 390 530 391 534
rect 395 530 396 534
rect 390 529 396 530
rect 422 530 423 534
rect 427 530 428 534
rect 454 534 460 535
rect 422 529 428 530
rect 446 531 452 532
rect 234 526 240 527
rect 446 527 447 531
rect 451 527 452 531
rect 454 530 455 534
rect 459 530 460 534
rect 486 534 492 535
rect 454 529 460 530
rect 466 531 472 532
rect 446 526 452 527
rect 466 527 467 531
rect 471 527 472 531
rect 486 530 487 534
rect 491 530 492 534
rect 486 529 492 530
rect 498 531 504 532
rect 466 526 472 527
rect 498 527 499 531
rect 503 527 504 531
rect 498 526 504 527
rect 110 524 116 525
rect 236 514 238 526
rect 236 512 242 514
rect 110 511 116 512
rect 110 507 111 511
rect 115 507 116 511
rect 110 506 116 507
rect 222 508 228 509
rect 112 503 114 506
rect 222 504 223 508
rect 227 504 228 508
rect 222 503 228 504
rect 230 503 236 504
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 135 497 139 498
rect 159 502 163 503
rect 159 497 163 498
rect 183 502 187 503
rect 183 497 187 498
rect 223 502 227 503
rect 230 499 231 503
rect 235 499 236 503
rect 240 500 242 512
rect 246 508 252 509
rect 246 504 247 508
rect 251 504 252 508
rect 246 503 252 504
rect 270 508 276 509
rect 270 504 271 508
rect 275 504 276 508
rect 270 503 276 504
rect 294 508 300 509
rect 294 504 295 508
rect 299 504 300 508
rect 294 503 300 504
rect 326 508 332 509
rect 326 504 327 508
rect 331 504 332 508
rect 326 503 332 504
rect 358 508 364 509
rect 358 504 359 508
rect 363 504 364 508
rect 358 503 364 504
rect 390 508 396 509
rect 390 504 391 508
rect 395 504 396 508
rect 390 503 396 504
rect 422 508 428 509
rect 422 504 423 508
rect 427 504 428 508
rect 422 503 428 504
rect 247 502 251 503
rect 230 498 236 499
rect 238 499 244 500
rect 223 497 227 498
rect 112 494 114 497
rect 134 496 140 497
rect 110 493 116 494
rect 110 489 111 493
rect 115 489 116 493
rect 134 492 135 496
rect 139 492 140 496
rect 134 491 140 492
rect 158 496 164 497
rect 158 492 159 496
rect 163 492 164 496
rect 158 491 164 492
rect 182 496 188 497
rect 182 492 183 496
rect 187 492 188 496
rect 182 491 188 492
rect 222 496 228 497
rect 222 492 223 496
rect 227 492 228 496
rect 222 491 228 492
rect 110 488 116 489
rect 110 475 116 476
rect 110 471 111 475
rect 115 471 116 475
rect 110 470 116 471
rect 134 470 140 471
rect 112 463 114 470
rect 134 466 135 470
rect 139 466 140 470
rect 134 465 140 466
rect 158 470 164 471
rect 158 466 159 470
rect 163 466 164 470
rect 158 465 164 466
rect 182 470 188 471
rect 182 466 183 470
rect 187 466 188 470
rect 182 465 188 466
rect 222 470 228 471
rect 222 466 223 470
rect 227 466 228 470
rect 222 465 228 466
rect 136 463 138 465
rect 160 463 162 465
rect 184 463 186 465
rect 224 463 226 465
rect 232 464 234 498
rect 238 495 239 499
rect 243 495 244 499
rect 247 497 251 498
rect 271 502 275 503
rect 271 497 275 498
rect 295 502 299 503
rect 295 497 299 498
rect 319 502 323 503
rect 319 497 323 498
rect 327 502 331 503
rect 327 497 331 498
rect 359 502 363 503
rect 359 497 363 498
rect 375 502 379 503
rect 375 497 379 498
rect 391 502 395 503
rect 391 497 395 498
rect 423 502 427 503
rect 423 497 427 498
rect 431 502 435 503
rect 431 497 435 498
rect 238 494 244 495
rect 270 496 276 497
rect 270 492 271 496
rect 275 492 276 496
rect 270 491 276 492
rect 318 496 324 497
rect 318 492 319 496
rect 323 492 324 496
rect 318 491 324 492
rect 374 496 380 497
rect 374 492 375 496
rect 379 492 380 496
rect 374 491 380 492
rect 430 496 436 497
rect 430 492 431 496
rect 435 492 436 496
rect 430 491 436 492
rect 362 487 368 488
rect 362 483 363 487
rect 367 483 368 487
rect 362 482 368 483
rect 270 470 276 471
rect 270 466 271 470
rect 275 466 276 470
rect 270 465 276 466
rect 318 470 324 471
rect 318 466 319 470
rect 323 466 324 470
rect 318 465 324 466
rect 230 463 236 464
rect 272 463 274 465
rect 320 463 322 465
rect 111 462 115 463
rect 111 457 115 458
rect 135 462 139 463
rect 135 457 139 458
rect 159 462 163 463
rect 159 457 163 458
rect 183 462 187 463
rect 183 457 187 458
rect 191 462 195 463
rect 191 457 195 458
rect 223 462 227 463
rect 230 459 231 463
rect 235 459 236 463
rect 230 458 236 459
rect 239 462 243 463
rect 223 457 227 458
rect 239 457 243 458
rect 271 462 275 463
rect 271 457 275 458
rect 295 462 299 463
rect 295 457 299 458
rect 319 462 323 463
rect 319 457 323 458
rect 351 462 355 463
rect 351 457 355 458
rect 112 450 114 457
rect 136 455 138 457
rect 160 455 162 457
rect 192 455 194 457
rect 240 455 242 457
rect 296 455 298 457
rect 352 455 354 457
rect 364 456 366 482
rect 448 480 450 526
rect 454 523 460 524
rect 468 523 470 526
rect 454 519 455 523
rect 459 521 470 523
rect 486 523 492 524
rect 500 523 502 526
rect 516 524 518 542
rect 527 537 531 538
rect 528 535 530 537
rect 540 536 542 554
rect 620 552 622 561
rect 676 552 678 562
rect 618 551 624 552
rect 674 551 680 552
rect 550 550 556 551
rect 550 546 551 550
rect 555 546 556 550
rect 550 545 556 546
rect 606 550 612 551
rect 606 546 607 550
rect 611 546 612 550
rect 618 547 619 551
rect 623 547 624 551
rect 618 546 624 547
rect 662 550 668 551
rect 662 546 663 550
rect 667 546 668 550
rect 674 547 675 551
rect 679 547 680 551
rect 674 546 680 547
rect 718 550 724 551
rect 718 546 719 550
rect 723 546 724 550
rect 774 550 780 551
rect 606 545 612 546
rect 662 545 668 546
rect 718 545 724 546
rect 730 547 736 548
rect 552 543 554 545
rect 586 543 592 544
rect 608 543 610 545
rect 664 543 666 545
rect 720 543 722 545
rect 730 543 731 547
rect 735 543 736 547
rect 774 546 775 550
rect 779 546 780 550
rect 774 545 780 546
rect 830 550 836 551
rect 830 546 831 550
rect 835 546 836 550
rect 830 545 836 546
rect 776 543 778 545
rect 832 543 834 545
rect 872 544 874 582
rect 879 577 883 578
rect 887 582 891 583
rect 887 577 891 578
rect 927 582 931 583
rect 927 577 931 578
rect 943 582 947 583
rect 943 577 947 578
rect 975 582 979 583
rect 975 577 979 578
rect 1007 582 1011 583
rect 1007 577 1011 578
rect 1023 582 1027 583
rect 1023 577 1027 578
rect 1071 582 1075 583
rect 1071 577 1075 578
rect 1111 582 1115 583
rect 1111 577 1115 578
rect 1127 582 1131 583
rect 1127 577 1131 578
rect 1151 582 1155 583
rect 1151 577 1155 578
rect 1183 582 1187 583
rect 1183 577 1187 578
rect 1191 582 1195 583
rect 1191 577 1195 578
rect 1239 582 1243 583
rect 1239 577 1243 578
rect 1247 582 1251 583
rect 1247 577 1251 578
rect 1287 582 1291 583
rect 1287 577 1291 578
rect 1311 582 1315 583
rect 1311 577 1315 578
rect 1335 582 1339 583
rect 1335 577 1339 578
rect 1375 582 1379 583
rect 1386 582 1392 583
rect 1447 582 1451 583
rect 1375 577 1379 578
rect 886 576 892 577
rect 886 572 887 576
rect 891 572 892 576
rect 886 571 892 572
rect 942 576 948 577
rect 942 572 943 576
rect 947 572 948 576
rect 942 571 948 572
rect 1006 576 1012 577
rect 1006 572 1007 576
rect 1011 572 1012 576
rect 1006 571 1012 572
rect 1070 576 1076 577
rect 1070 572 1071 576
rect 1075 572 1076 576
rect 1070 571 1076 572
rect 1126 576 1132 577
rect 1126 572 1127 576
rect 1131 572 1132 576
rect 1126 571 1132 572
rect 1182 576 1188 577
rect 1182 572 1183 576
rect 1187 572 1188 576
rect 1182 571 1188 572
rect 1246 576 1252 577
rect 1246 572 1247 576
rect 1251 572 1252 576
rect 1246 571 1252 572
rect 1310 576 1316 577
rect 1310 572 1311 576
rect 1315 572 1316 576
rect 1310 571 1316 572
rect 1374 576 1380 577
rect 1374 572 1375 576
rect 1379 572 1380 576
rect 1374 571 1380 572
rect 1034 567 1040 568
rect 1034 563 1035 567
rect 1039 563 1040 567
rect 1034 562 1040 563
rect 1138 567 1144 568
rect 1138 563 1139 567
rect 1143 563 1144 567
rect 1138 562 1144 563
rect 886 550 892 551
rect 886 546 887 550
rect 891 546 892 550
rect 886 545 892 546
rect 942 550 948 551
rect 942 546 943 550
rect 947 546 948 550
rect 942 545 948 546
rect 1006 550 1012 551
rect 1006 546 1007 550
rect 1011 546 1012 550
rect 1006 545 1012 546
rect 870 543 876 544
rect 888 543 890 545
rect 944 543 946 545
rect 1008 543 1010 545
rect 551 542 555 543
rect 551 537 555 538
rect 575 542 579 543
rect 586 539 587 543
rect 591 539 592 543
rect 586 538 592 539
rect 607 542 611 543
rect 575 537 579 538
rect 538 535 544 536
rect 576 535 578 537
rect 526 534 532 535
rect 526 530 527 534
rect 531 530 532 534
rect 538 531 539 535
rect 543 531 544 535
rect 538 530 544 531
rect 574 534 580 535
rect 574 530 575 534
rect 579 530 580 534
rect 526 529 532 530
rect 574 529 580 530
rect 459 519 460 521
rect 454 518 460 519
rect 486 519 487 523
rect 491 521 502 523
rect 514 523 520 524
rect 491 519 492 521
rect 486 518 492 519
rect 514 519 515 523
rect 519 519 520 523
rect 514 518 520 519
rect 588 516 590 538
rect 607 537 611 538
rect 623 542 627 543
rect 623 537 627 538
rect 663 542 667 543
rect 663 537 667 538
rect 671 542 675 543
rect 671 537 675 538
rect 711 542 715 543
rect 711 537 715 538
rect 719 542 723 543
rect 730 542 736 543
rect 759 542 763 543
rect 719 537 723 538
rect 624 535 626 537
rect 672 535 674 537
rect 712 535 714 537
rect 622 534 628 535
rect 622 530 623 534
rect 627 530 628 534
rect 622 529 628 530
rect 670 534 676 535
rect 670 530 671 534
rect 675 530 676 534
rect 670 529 676 530
rect 710 534 716 535
rect 710 530 711 534
rect 715 530 716 534
rect 710 529 716 530
rect 732 524 734 542
rect 759 537 763 538
rect 775 542 779 543
rect 775 537 779 538
rect 807 542 811 543
rect 807 537 811 538
rect 831 542 835 543
rect 831 537 835 538
rect 855 542 859 543
rect 870 539 871 543
rect 875 539 876 543
rect 870 538 876 539
rect 887 542 891 543
rect 855 537 859 538
rect 887 537 891 538
rect 911 542 915 543
rect 911 537 915 538
rect 943 542 947 543
rect 943 537 947 538
rect 967 542 971 543
rect 967 537 971 538
rect 1007 542 1011 543
rect 1007 537 1011 538
rect 1023 542 1027 543
rect 1023 537 1027 538
rect 760 535 762 537
rect 808 535 810 537
rect 856 535 858 537
rect 912 535 914 537
rect 968 535 970 537
rect 1024 535 1026 537
rect 1036 536 1038 562
rect 1140 552 1142 562
rect 1282 559 1288 560
rect 1282 555 1283 559
rect 1287 555 1288 559
rect 1282 554 1288 555
rect 1138 551 1144 552
rect 1070 550 1076 551
rect 1070 546 1071 550
rect 1075 546 1076 550
rect 1126 550 1132 551
rect 1070 545 1076 546
rect 1090 547 1096 548
rect 1072 543 1074 545
rect 1090 543 1091 547
rect 1095 543 1096 547
rect 1126 546 1127 550
rect 1131 546 1132 550
rect 1138 547 1139 551
rect 1143 547 1144 551
rect 1138 546 1144 547
rect 1182 550 1188 551
rect 1182 546 1183 550
rect 1187 546 1188 550
rect 1126 545 1132 546
rect 1182 545 1188 546
rect 1246 550 1252 551
rect 1246 546 1247 550
rect 1251 546 1252 550
rect 1246 545 1252 546
rect 1128 543 1130 545
rect 1184 543 1186 545
rect 1248 543 1250 545
rect 1071 542 1075 543
rect 1071 537 1075 538
rect 1079 542 1083 543
rect 1090 542 1096 543
rect 1127 542 1131 543
rect 1079 537 1083 538
rect 1034 535 1040 536
rect 1080 535 1082 537
rect 758 534 764 535
rect 758 530 759 534
rect 763 530 764 534
rect 758 529 764 530
rect 806 534 812 535
rect 806 530 807 534
rect 811 530 812 534
rect 806 529 812 530
rect 854 534 860 535
rect 854 530 855 534
rect 859 530 860 534
rect 854 529 860 530
rect 910 534 916 535
rect 910 530 911 534
rect 915 530 916 534
rect 910 529 916 530
rect 966 534 972 535
rect 966 530 967 534
rect 971 530 972 534
rect 966 529 972 530
rect 1022 534 1028 535
rect 1022 530 1023 534
rect 1027 530 1028 534
rect 1034 531 1035 535
rect 1039 531 1040 535
rect 1034 530 1040 531
rect 1078 534 1084 535
rect 1078 530 1079 534
rect 1083 530 1084 534
rect 1022 529 1028 530
rect 1078 529 1084 530
rect 1092 524 1094 542
rect 1127 537 1131 538
rect 1175 542 1179 543
rect 1175 537 1179 538
rect 1183 542 1187 543
rect 1183 537 1187 538
rect 1223 542 1227 543
rect 1223 537 1227 538
rect 1247 542 1251 543
rect 1247 537 1251 538
rect 1271 542 1275 543
rect 1271 537 1275 538
rect 1128 535 1130 537
rect 1176 535 1178 537
rect 1224 535 1226 537
rect 1272 535 1274 537
rect 1284 536 1286 554
rect 1388 552 1390 582
rect 1447 577 1451 578
rect 1448 574 1450 577
rect 1446 573 1452 574
rect 1446 569 1447 573
rect 1451 569 1452 573
rect 1446 568 1452 569
rect 1446 555 1452 556
rect 1386 551 1392 552
rect 1310 550 1316 551
rect 1310 546 1311 550
rect 1315 546 1316 550
rect 1310 545 1316 546
rect 1374 550 1380 551
rect 1374 546 1375 550
rect 1379 546 1380 550
rect 1386 547 1387 551
rect 1391 547 1392 551
rect 1446 551 1447 555
rect 1451 551 1452 555
rect 1446 550 1452 551
rect 1386 546 1392 547
rect 1374 545 1380 546
rect 1312 543 1314 545
rect 1362 543 1368 544
rect 1376 543 1378 545
rect 1448 543 1450 550
rect 1311 542 1315 543
rect 1311 537 1315 538
rect 1351 542 1355 543
rect 1362 539 1363 543
rect 1367 539 1368 543
rect 1362 538 1368 539
rect 1375 542 1379 543
rect 1351 537 1355 538
rect 1282 535 1288 536
rect 1312 535 1314 537
rect 1352 535 1354 537
rect 1126 534 1132 535
rect 1126 530 1127 534
rect 1131 530 1132 534
rect 1126 529 1132 530
rect 1174 534 1180 535
rect 1174 530 1175 534
rect 1179 530 1180 534
rect 1174 529 1180 530
rect 1222 534 1228 535
rect 1222 530 1223 534
rect 1227 530 1228 534
rect 1270 534 1276 535
rect 1222 529 1228 530
rect 1262 531 1268 532
rect 1262 527 1263 531
rect 1267 527 1268 531
rect 1270 530 1271 534
rect 1275 530 1276 534
rect 1282 531 1283 535
rect 1287 531 1288 535
rect 1282 530 1288 531
rect 1310 534 1316 535
rect 1310 530 1311 534
rect 1315 530 1316 534
rect 1270 529 1276 530
rect 1310 529 1316 530
rect 1350 534 1356 535
rect 1350 530 1351 534
rect 1355 530 1356 534
rect 1350 529 1356 530
rect 1262 526 1268 527
rect 730 523 736 524
rect 730 519 731 523
rect 735 519 736 523
rect 730 518 736 519
rect 1090 523 1096 524
rect 1090 519 1091 523
rect 1095 519 1096 523
rect 1090 518 1096 519
rect 586 515 592 516
rect 586 511 587 515
rect 591 511 592 515
rect 1264 515 1266 526
rect 1264 513 1282 515
rect 586 510 592 511
rect 454 508 460 509
rect 454 504 455 508
rect 459 504 460 508
rect 454 503 460 504
rect 486 508 492 509
rect 486 504 487 508
rect 491 504 492 508
rect 486 503 492 504
rect 526 508 532 509
rect 526 504 527 508
rect 531 504 532 508
rect 526 503 532 504
rect 574 508 580 509
rect 574 504 575 508
rect 579 504 580 508
rect 574 503 580 504
rect 622 508 628 509
rect 622 504 623 508
rect 627 504 628 508
rect 622 503 628 504
rect 670 508 676 509
rect 670 504 671 508
rect 675 504 676 508
rect 710 508 716 509
rect 710 504 711 508
rect 715 504 716 508
rect 670 503 676 504
rect 678 503 684 504
rect 710 503 716 504
rect 758 508 764 509
rect 758 504 759 508
rect 763 504 764 508
rect 758 503 764 504
rect 806 508 812 509
rect 806 504 807 508
rect 811 504 812 508
rect 806 503 812 504
rect 854 508 860 509
rect 854 504 855 508
rect 859 504 860 508
rect 854 503 860 504
rect 910 508 916 509
rect 910 504 911 508
rect 915 504 916 508
rect 910 503 916 504
rect 966 508 972 509
rect 966 504 967 508
rect 971 504 972 508
rect 966 503 972 504
rect 1022 508 1028 509
rect 1022 504 1023 508
rect 1027 504 1028 508
rect 1022 503 1028 504
rect 1078 508 1084 509
rect 1078 504 1079 508
rect 1083 504 1084 508
rect 1078 503 1084 504
rect 1126 508 1132 509
rect 1126 504 1127 508
rect 1131 504 1132 508
rect 1126 503 1132 504
rect 1174 508 1180 509
rect 1174 504 1175 508
rect 1179 504 1180 508
rect 1174 503 1180 504
rect 1222 508 1228 509
rect 1222 504 1223 508
rect 1227 504 1228 508
rect 1222 503 1228 504
rect 1270 508 1276 509
rect 1270 504 1271 508
rect 1275 504 1276 508
rect 1270 503 1276 504
rect 455 502 459 503
rect 455 497 459 498
rect 487 502 491 503
rect 487 497 491 498
rect 527 502 531 503
rect 527 497 531 498
rect 543 502 547 503
rect 543 497 547 498
rect 575 502 579 503
rect 575 497 579 498
rect 591 502 595 503
rect 591 497 595 498
rect 623 502 627 503
rect 623 497 627 498
rect 631 502 635 503
rect 631 497 635 498
rect 663 502 667 503
rect 663 497 667 498
rect 671 502 675 503
rect 678 499 679 503
rect 683 499 684 503
rect 678 498 684 499
rect 687 502 691 503
rect 671 497 675 498
rect 486 496 492 497
rect 486 492 487 496
rect 491 492 492 496
rect 486 491 492 492
rect 542 496 548 497
rect 542 492 543 496
rect 547 492 548 496
rect 542 491 548 492
rect 590 496 596 497
rect 590 492 591 496
rect 595 492 596 496
rect 590 491 596 492
rect 630 496 636 497
rect 630 492 631 496
rect 635 492 636 496
rect 630 491 636 492
rect 662 496 668 497
rect 662 492 663 496
rect 667 492 668 496
rect 662 491 668 492
rect 680 491 682 498
rect 687 497 691 498
rect 711 502 715 503
rect 711 497 715 498
rect 719 502 723 503
rect 719 497 723 498
rect 759 502 763 503
rect 759 497 763 498
rect 799 502 803 503
rect 799 497 803 498
rect 807 502 811 503
rect 807 497 811 498
rect 847 502 851 503
rect 847 497 851 498
rect 855 502 859 503
rect 855 497 859 498
rect 903 502 907 503
rect 903 497 907 498
rect 911 502 915 503
rect 911 497 915 498
rect 951 502 955 503
rect 951 497 955 498
rect 967 502 971 503
rect 967 497 971 498
rect 999 502 1003 503
rect 999 497 1003 498
rect 1023 502 1027 503
rect 1023 497 1027 498
rect 1047 502 1051 503
rect 1047 497 1051 498
rect 1079 502 1083 503
rect 1079 497 1083 498
rect 1095 502 1099 503
rect 1095 497 1099 498
rect 1127 502 1131 503
rect 1127 497 1131 498
rect 1143 502 1147 503
rect 1143 497 1147 498
rect 1175 502 1179 503
rect 1175 497 1179 498
rect 1199 502 1203 503
rect 1199 497 1203 498
rect 1223 502 1227 503
rect 1223 497 1227 498
rect 1255 502 1259 503
rect 1255 497 1259 498
rect 1271 502 1275 503
rect 1271 497 1275 498
rect 686 496 692 497
rect 686 492 687 496
rect 691 492 692 496
rect 686 491 692 492
rect 718 496 724 497
rect 718 492 719 496
rect 723 492 724 496
rect 718 491 724 492
rect 758 496 764 497
rect 758 492 759 496
rect 763 492 764 496
rect 758 491 764 492
rect 798 496 804 497
rect 798 492 799 496
rect 803 492 804 496
rect 798 491 804 492
rect 846 496 852 497
rect 846 492 847 496
rect 851 492 852 496
rect 846 491 852 492
rect 902 496 908 497
rect 902 492 903 496
rect 907 492 908 496
rect 902 491 908 492
rect 950 496 956 497
rect 950 492 951 496
rect 955 492 956 496
rect 950 491 956 492
rect 998 496 1004 497
rect 998 492 999 496
rect 1003 492 1004 496
rect 998 491 1004 492
rect 1046 496 1052 497
rect 1046 492 1047 496
rect 1051 492 1052 496
rect 1046 491 1052 492
rect 1094 496 1100 497
rect 1094 492 1095 496
rect 1099 492 1100 496
rect 1094 491 1100 492
rect 1142 496 1148 497
rect 1142 492 1143 496
rect 1147 492 1148 496
rect 1142 491 1148 492
rect 1198 496 1204 497
rect 1198 492 1199 496
rect 1203 492 1204 496
rect 1198 491 1204 492
rect 1254 496 1260 497
rect 1254 492 1255 496
rect 1259 492 1260 496
rect 1254 491 1260 492
rect 672 489 682 491
rect 498 487 504 488
rect 498 483 499 487
rect 503 483 504 487
rect 498 482 504 483
rect 602 487 608 488
rect 602 483 603 487
rect 607 483 608 487
rect 602 482 608 483
rect 446 479 452 480
rect 446 475 447 479
rect 451 475 452 479
rect 446 474 452 475
rect 500 472 502 482
rect 604 472 606 482
rect 672 475 674 489
rect 1280 488 1282 513
rect 1364 512 1366 538
rect 1375 537 1379 538
rect 1391 542 1395 543
rect 1391 537 1395 538
rect 1415 542 1419 543
rect 1415 537 1419 538
rect 1447 542 1451 543
rect 1447 537 1451 538
rect 1392 535 1394 537
rect 1416 535 1418 537
rect 1390 534 1396 535
rect 1390 530 1391 534
rect 1395 530 1396 534
rect 1390 529 1396 530
rect 1414 534 1420 535
rect 1414 530 1415 534
rect 1419 530 1420 534
rect 1448 530 1450 537
rect 1414 529 1420 530
rect 1446 529 1452 530
rect 1446 525 1447 529
rect 1451 525 1452 529
rect 1446 524 1452 525
rect 1362 511 1368 512
rect 1310 508 1316 509
rect 1310 504 1311 508
rect 1315 504 1316 508
rect 1310 503 1316 504
rect 1350 508 1356 509
rect 1350 504 1351 508
rect 1355 504 1356 508
rect 1362 507 1363 511
rect 1367 507 1368 511
rect 1446 511 1452 512
rect 1362 506 1368 507
rect 1390 508 1396 509
rect 1350 503 1356 504
rect 1390 504 1391 508
rect 1395 504 1396 508
rect 1390 503 1396 504
rect 1414 508 1420 509
rect 1414 504 1415 508
rect 1419 504 1420 508
rect 1414 503 1420 504
rect 1426 507 1432 508
rect 1426 503 1427 507
rect 1431 503 1432 507
rect 1446 507 1447 511
rect 1451 507 1452 511
rect 1446 506 1452 507
rect 1448 503 1450 506
rect 1311 502 1315 503
rect 1311 497 1315 498
rect 1351 502 1355 503
rect 1351 497 1355 498
rect 1375 502 1379 503
rect 1375 497 1379 498
rect 1391 502 1395 503
rect 1391 497 1395 498
rect 1415 502 1419 503
rect 1426 502 1432 503
rect 1447 502 1451 503
rect 1415 497 1419 498
rect 1310 496 1316 497
rect 1310 492 1311 496
rect 1315 492 1316 496
rect 1310 491 1316 492
rect 1374 496 1380 497
rect 1374 492 1375 496
rect 1379 492 1380 496
rect 1374 491 1380 492
rect 1414 496 1420 497
rect 1414 492 1415 496
rect 1419 492 1420 496
rect 1414 491 1420 492
rect 730 487 736 488
rect 730 483 731 487
rect 735 483 736 487
rect 730 482 736 483
rect 810 487 816 488
rect 810 483 811 487
rect 815 483 816 487
rect 810 482 816 483
rect 818 487 824 488
rect 818 483 819 487
rect 823 483 824 487
rect 818 482 824 483
rect 894 487 900 488
rect 894 483 895 487
rect 899 483 900 487
rect 894 482 900 483
rect 962 487 968 488
rect 962 483 963 487
rect 967 483 968 487
rect 962 482 968 483
rect 1058 487 1064 488
rect 1058 483 1059 487
rect 1063 483 1064 487
rect 1058 482 1064 483
rect 1154 487 1160 488
rect 1154 483 1155 487
rect 1159 483 1160 487
rect 1154 482 1160 483
rect 1266 487 1272 488
rect 1266 483 1267 487
rect 1271 483 1272 487
rect 1266 482 1272 483
rect 1278 487 1284 488
rect 1278 483 1279 487
rect 1283 483 1284 487
rect 1278 482 1284 483
rect 1382 483 1388 484
rect 656 473 674 475
rect 678 479 684 480
rect 678 475 679 479
rect 683 475 684 479
rect 678 474 684 475
rect 498 471 504 472
rect 602 471 608 472
rect 374 470 380 471
rect 374 466 375 470
rect 379 466 380 470
rect 374 465 380 466
rect 430 470 436 471
rect 430 466 431 470
rect 435 466 436 470
rect 486 470 492 471
rect 430 465 436 466
rect 442 467 448 468
rect 376 463 378 465
rect 432 463 434 465
rect 442 463 443 467
rect 447 463 448 467
rect 486 466 487 470
rect 491 466 492 470
rect 498 467 499 471
rect 503 467 504 471
rect 498 466 504 467
rect 542 470 548 471
rect 542 466 543 470
rect 547 466 548 470
rect 486 465 492 466
rect 542 465 548 466
rect 590 470 596 471
rect 590 466 591 470
rect 595 466 596 470
rect 602 467 603 471
rect 607 467 608 471
rect 602 466 608 467
rect 630 470 636 471
rect 630 466 631 470
rect 635 466 636 470
rect 590 465 596 466
rect 630 465 636 466
rect 488 463 490 465
rect 544 463 546 465
rect 592 463 594 465
rect 632 463 634 465
rect 656 464 658 473
rect 662 470 668 471
rect 662 466 663 470
rect 667 466 668 470
rect 662 465 668 466
rect 654 463 660 464
rect 664 463 666 465
rect 375 462 379 463
rect 375 457 379 458
rect 415 462 419 463
rect 415 457 419 458
rect 431 462 435 463
rect 442 462 448 463
rect 479 462 483 463
rect 431 457 435 458
rect 362 455 368 456
rect 416 455 418 457
rect 134 454 140 455
rect 134 450 135 454
rect 139 450 140 454
rect 110 449 116 450
rect 134 449 140 450
rect 158 454 164 455
rect 158 450 159 454
rect 163 450 164 454
rect 158 449 164 450
rect 190 454 196 455
rect 190 450 191 454
rect 195 450 196 454
rect 190 449 196 450
rect 238 454 244 455
rect 238 450 239 454
rect 243 450 244 454
rect 238 449 244 450
rect 294 454 300 455
rect 294 450 295 454
rect 299 450 300 454
rect 294 449 300 450
rect 350 454 356 455
rect 350 450 351 454
rect 355 450 356 454
rect 362 451 363 455
rect 367 451 368 455
rect 362 450 368 451
rect 414 454 420 455
rect 414 450 415 454
rect 419 450 420 454
rect 350 449 356 450
rect 414 449 420 450
rect 110 445 111 449
rect 115 445 116 449
rect 110 444 116 445
rect 444 444 446 462
rect 479 457 483 458
rect 487 462 491 463
rect 487 457 491 458
rect 543 462 547 463
rect 543 457 547 458
rect 591 462 595 463
rect 591 457 595 458
rect 607 462 611 463
rect 607 457 611 458
rect 631 462 635 463
rect 654 459 655 463
rect 659 459 660 463
rect 654 458 660 459
rect 663 462 667 463
rect 631 457 635 458
rect 663 457 667 458
rect 671 462 675 463
rect 671 457 675 458
rect 480 455 482 457
rect 544 455 546 457
rect 608 455 610 457
rect 672 455 674 457
rect 478 454 484 455
rect 478 450 479 454
rect 483 450 484 454
rect 478 449 484 450
rect 542 454 548 455
rect 542 450 543 454
rect 547 450 548 454
rect 542 449 548 450
rect 606 454 612 455
rect 606 450 607 454
rect 611 450 612 454
rect 670 454 676 455
rect 606 449 612 450
rect 618 451 624 452
rect 618 447 619 451
rect 623 447 624 451
rect 670 450 671 454
rect 675 450 676 454
rect 670 449 676 450
rect 680 452 682 474
rect 732 472 734 482
rect 812 472 814 482
rect 730 471 736 472
rect 810 471 816 472
rect 686 470 692 471
rect 686 466 687 470
rect 691 466 692 470
rect 686 465 692 466
rect 718 470 724 471
rect 718 466 719 470
rect 723 466 724 470
rect 730 467 731 471
rect 735 467 736 471
rect 730 466 736 467
rect 758 470 764 471
rect 758 466 759 470
rect 763 466 764 470
rect 718 465 724 466
rect 758 465 764 466
rect 798 470 804 471
rect 798 466 799 470
rect 803 466 804 470
rect 810 467 811 471
rect 815 467 816 471
rect 810 466 816 467
rect 798 465 804 466
rect 688 463 690 465
rect 710 463 716 464
rect 720 463 722 465
rect 760 463 762 465
rect 800 463 802 465
rect 687 462 691 463
rect 710 459 711 463
rect 715 459 716 463
rect 710 458 716 459
rect 719 462 723 463
rect 687 457 691 458
rect 680 451 688 452
rect 680 449 683 451
rect 618 446 624 447
rect 682 447 683 449
rect 687 447 688 451
rect 682 446 688 447
rect 442 443 448 444
rect 126 439 132 440
rect 126 435 127 439
rect 131 435 132 439
rect 442 439 443 443
rect 447 439 448 443
rect 442 438 448 439
rect 126 434 132 435
rect 110 431 116 432
rect 110 427 111 431
rect 115 427 116 431
rect 110 426 116 427
rect 112 423 114 426
rect 111 422 115 423
rect 111 417 115 418
rect 112 414 114 417
rect 110 413 116 414
rect 110 409 111 413
rect 115 409 116 413
rect 110 408 116 409
rect 110 395 116 396
rect 110 391 111 395
rect 115 391 116 395
rect 110 390 116 391
rect 112 379 114 390
rect 128 384 130 434
rect 134 428 140 429
rect 134 424 135 428
rect 139 424 140 428
rect 134 423 140 424
rect 158 428 164 429
rect 158 424 159 428
rect 163 424 164 428
rect 158 423 164 424
rect 190 428 196 429
rect 190 424 191 428
rect 195 424 196 428
rect 190 423 196 424
rect 238 428 244 429
rect 238 424 239 428
rect 243 424 244 428
rect 238 423 244 424
rect 294 428 300 429
rect 294 424 295 428
rect 299 424 300 428
rect 294 423 300 424
rect 350 428 356 429
rect 350 424 351 428
rect 355 424 356 428
rect 350 423 356 424
rect 414 428 420 429
rect 414 424 415 428
rect 419 424 420 428
rect 414 423 420 424
rect 478 428 484 429
rect 478 424 479 428
rect 483 424 484 428
rect 478 423 484 424
rect 542 428 548 429
rect 542 424 543 428
rect 547 424 548 428
rect 542 423 548 424
rect 606 428 612 429
rect 606 424 607 428
rect 611 424 612 428
rect 606 423 612 424
rect 135 422 139 423
rect 135 417 139 418
rect 159 422 163 423
rect 159 417 163 418
rect 183 422 187 423
rect 183 417 187 418
rect 191 422 195 423
rect 191 417 195 418
rect 215 422 219 423
rect 215 417 219 418
rect 239 422 243 423
rect 239 417 243 418
rect 271 422 275 423
rect 271 417 275 418
rect 295 422 299 423
rect 295 417 299 418
rect 327 422 331 423
rect 327 417 331 418
rect 351 422 355 423
rect 351 417 355 418
rect 391 422 395 423
rect 391 417 395 418
rect 415 422 419 423
rect 415 417 419 418
rect 447 422 451 423
rect 447 417 451 418
rect 479 422 483 423
rect 479 417 483 418
rect 503 422 507 423
rect 503 417 507 418
rect 543 422 547 423
rect 543 417 547 418
rect 551 422 555 423
rect 551 417 555 418
rect 599 422 603 423
rect 599 417 603 418
rect 607 422 611 423
rect 607 417 611 418
rect 134 416 140 417
rect 134 412 135 416
rect 139 412 140 416
rect 134 411 140 412
rect 158 416 164 417
rect 158 412 159 416
rect 163 412 164 416
rect 158 411 164 412
rect 182 416 188 417
rect 182 412 183 416
rect 187 412 188 416
rect 182 411 188 412
rect 214 416 220 417
rect 214 412 215 416
rect 219 412 220 416
rect 214 411 220 412
rect 270 416 276 417
rect 270 412 271 416
rect 275 412 276 416
rect 270 411 276 412
rect 326 416 332 417
rect 326 412 327 416
rect 331 412 332 416
rect 326 411 332 412
rect 390 416 396 417
rect 390 412 391 416
rect 395 412 396 416
rect 390 411 396 412
rect 446 416 452 417
rect 446 412 447 416
rect 451 412 452 416
rect 446 411 452 412
rect 502 416 508 417
rect 502 412 503 416
rect 507 412 508 416
rect 502 411 508 412
rect 550 416 556 417
rect 550 412 551 416
rect 555 412 556 416
rect 550 411 556 412
rect 598 416 604 417
rect 598 412 599 416
rect 603 412 604 416
rect 598 411 604 412
rect 620 408 622 446
rect 712 436 714 458
rect 719 457 723 458
rect 735 462 739 463
rect 735 457 739 458
rect 759 462 763 463
rect 759 457 763 458
rect 791 462 795 463
rect 791 457 795 458
rect 799 462 803 463
rect 799 457 803 458
rect 736 455 738 457
rect 792 455 794 457
rect 820 456 822 482
rect 896 475 898 482
rect 918 479 924 480
rect 918 475 919 479
rect 923 475 924 479
rect 896 474 924 475
rect 896 473 922 474
rect 964 472 966 482
rect 1060 472 1062 482
rect 1156 472 1158 482
rect 1268 472 1270 482
rect 1382 479 1383 483
rect 1387 479 1388 483
rect 1382 478 1388 479
rect 962 471 968 472
rect 1058 471 1064 472
rect 1154 471 1160 472
rect 1266 471 1272 472
rect 846 470 852 471
rect 846 466 847 470
rect 851 466 852 470
rect 846 465 852 466
rect 902 470 908 471
rect 902 466 903 470
rect 907 466 908 470
rect 902 465 908 466
rect 950 470 956 471
rect 950 466 951 470
rect 955 466 956 470
rect 962 467 963 471
rect 967 467 968 471
rect 962 466 968 467
rect 998 470 1004 471
rect 998 466 999 470
rect 1003 466 1004 470
rect 950 465 956 466
rect 998 465 1004 466
rect 1046 470 1052 471
rect 1046 466 1047 470
rect 1051 466 1052 470
rect 1058 467 1059 471
rect 1063 467 1064 471
rect 1058 466 1064 467
rect 1094 470 1100 471
rect 1094 466 1095 470
rect 1099 466 1100 470
rect 1046 465 1052 466
rect 1094 465 1100 466
rect 1142 470 1148 471
rect 1142 466 1143 470
rect 1147 466 1148 470
rect 1154 467 1155 471
rect 1159 467 1160 471
rect 1154 466 1160 467
rect 1198 470 1204 471
rect 1198 466 1199 470
rect 1203 466 1204 470
rect 1142 465 1148 466
rect 1198 465 1204 466
rect 1254 470 1260 471
rect 1254 466 1255 470
rect 1259 466 1260 470
rect 1266 467 1267 471
rect 1271 467 1272 471
rect 1266 466 1272 467
rect 1310 470 1316 471
rect 1310 466 1311 470
rect 1315 466 1316 470
rect 1254 465 1260 466
rect 1310 465 1316 466
rect 1374 470 1380 471
rect 1374 466 1375 470
rect 1379 466 1380 470
rect 1374 465 1380 466
rect 848 463 850 465
rect 904 463 906 465
rect 922 463 928 464
rect 952 463 954 465
rect 1000 463 1002 465
rect 1048 463 1050 465
rect 1096 463 1098 465
rect 1144 463 1146 465
rect 1200 463 1202 465
rect 1256 463 1258 465
rect 1312 463 1314 465
rect 1376 463 1378 465
rect 839 462 843 463
rect 839 457 843 458
rect 847 462 851 463
rect 847 457 851 458
rect 879 462 883 463
rect 879 457 883 458
rect 903 462 907 463
rect 903 457 907 458
rect 911 462 915 463
rect 922 459 923 463
rect 927 459 928 463
rect 922 458 928 459
rect 943 462 947 463
rect 911 457 915 458
rect 818 455 824 456
rect 840 455 842 457
rect 880 455 882 457
rect 912 455 914 457
rect 734 454 740 455
rect 734 450 735 454
rect 739 450 740 454
rect 734 449 740 450
rect 790 454 796 455
rect 790 450 791 454
rect 795 450 796 454
rect 818 451 819 455
rect 823 451 824 455
rect 818 450 824 451
rect 838 454 844 455
rect 838 450 839 454
rect 843 450 844 454
rect 878 454 884 455
rect 790 449 796 450
rect 838 449 844 450
rect 850 451 856 452
rect 850 447 851 451
rect 855 447 856 451
rect 878 450 879 454
rect 883 450 884 454
rect 910 454 916 455
rect 878 449 884 450
rect 890 451 896 452
rect 850 446 856 447
rect 890 447 891 451
rect 895 447 896 451
rect 910 450 911 454
rect 915 450 916 454
rect 910 449 916 450
rect 890 446 896 447
rect 838 443 844 444
rect 852 443 854 446
rect 838 439 839 443
rect 843 441 854 443
rect 878 443 884 444
rect 892 443 894 446
rect 843 439 844 441
rect 838 438 844 439
rect 878 439 879 443
rect 883 441 894 443
rect 883 439 884 441
rect 878 438 884 439
rect 924 436 926 458
rect 943 457 947 458
rect 951 462 955 463
rect 951 457 955 458
rect 967 462 971 463
rect 967 457 971 458
rect 999 462 1003 463
rect 999 457 1003 458
rect 1031 462 1035 463
rect 1031 457 1035 458
rect 1047 462 1051 463
rect 1047 457 1051 458
rect 1071 462 1075 463
rect 1071 457 1075 458
rect 1095 462 1099 463
rect 1095 457 1099 458
rect 1119 462 1123 463
rect 1119 457 1123 458
rect 1143 462 1147 463
rect 1143 457 1147 458
rect 1175 462 1179 463
rect 1175 457 1179 458
rect 1199 462 1203 463
rect 1199 457 1203 458
rect 1239 462 1243 463
rect 1239 457 1243 458
rect 1255 462 1259 463
rect 1255 457 1259 458
rect 1303 462 1307 463
rect 1303 457 1307 458
rect 1311 462 1315 463
rect 1311 457 1315 458
rect 1367 462 1371 463
rect 1367 457 1371 458
rect 1375 462 1379 463
rect 1375 457 1379 458
rect 944 455 946 457
rect 968 455 970 457
rect 1000 455 1002 457
rect 1032 455 1034 457
rect 1072 455 1074 457
rect 1120 455 1122 457
rect 1176 455 1178 457
rect 1240 455 1242 457
rect 1304 455 1306 457
rect 1368 455 1370 457
rect 942 454 948 455
rect 942 450 943 454
rect 947 450 948 454
rect 942 449 948 450
rect 966 454 972 455
rect 966 450 967 454
rect 971 450 972 454
rect 966 449 972 450
rect 998 454 1004 455
rect 998 450 999 454
rect 1003 450 1004 454
rect 1030 454 1036 455
rect 998 449 1004 450
rect 1022 451 1028 452
rect 1022 447 1023 451
rect 1027 447 1028 451
rect 1030 450 1031 454
rect 1035 450 1036 454
rect 1030 449 1036 450
rect 1070 454 1076 455
rect 1070 450 1071 454
rect 1075 450 1076 454
rect 1070 449 1076 450
rect 1118 454 1124 455
rect 1118 450 1119 454
rect 1123 450 1124 454
rect 1118 449 1124 450
rect 1174 454 1180 455
rect 1174 450 1175 454
rect 1179 450 1180 454
rect 1174 449 1180 450
rect 1238 454 1244 455
rect 1238 450 1239 454
rect 1243 450 1244 454
rect 1238 449 1244 450
rect 1302 454 1308 455
rect 1302 450 1303 454
rect 1307 450 1308 454
rect 1366 454 1372 455
rect 1302 449 1308 450
rect 1330 451 1336 452
rect 1022 446 1028 447
rect 1330 447 1331 451
rect 1335 447 1336 451
rect 1366 450 1367 454
rect 1371 450 1372 454
rect 1366 449 1372 450
rect 1375 451 1381 452
rect 1330 446 1336 447
rect 1375 447 1376 451
rect 1380 450 1381 451
rect 1384 450 1386 478
rect 1428 472 1430 502
rect 1447 497 1451 498
rect 1448 494 1450 497
rect 1446 493 1452 494
rect 1446 489 1447 493
rect 1451 489 1452 493
rect 1446 488 1452 489
rect 1446 475 1452 476
rect 1426 471 1432 472
rect 1414 470 1420 471
rect 1414 466 1415 470
rect 1419 466 1420 470
rect 1426 467 1427 471
rect 1431 467 1432 471
rect 1446 471 1447 475
rect 1451 471 1452 475
rect 1446 470 1452 471
rect 1426 466 1432 467
rect 1414 465 1420 466
rect 1416 463 1418 465
rect 1448 463 1450 470
rect 1415 462 1419 463
rect 1415 457 1419 458
rect 1447 462 1451 463
rect 1447 457 1451 458
rect 1416 455 1418 457
rect 1380 448 1386 450
rect 1414 454 1420 455
rect 1414 450 1415 454
rect 1419 450 1420 454
rect 1448 450 1450 457
rect 1414 449 1420 450
rect 1446 449 1452 450
rect 1380 447 1381 448
rect 1375 446 1381 447
rect 710 435 716 436
rect 710 431 711 435
rect 715 431 716 435
rect 710 430 716 431
rect 922 435 928 436
rect 922 431 923 435
rect 927 431 928 435
rect 922 430 928 431
rect 670 428 676 429
rect 670 424 671 428
rect 675 424 676 428
rect 670 423 676 424
rect 734 428 740 429
rect 734 424 735 428
rect 739 424 740 428
rect 734 423 740 424
rect 790 428 796 429
rect 790 424 791 428
rect 795 424 796 428
rect 790 423 796 424
rect 838 428 844 429
rect 838 424 839 428
rect 843 424 844 428
rect 838 423 844 424
rect 878 428 884 429
rect 878 424 879 428
rect 883 424 884 428
rect 878 423 884 424
rect 910 428 916 429
rect 910 424 911 428
rect 915 424 916 428
rect 910 423 916 424
rect 942 428 948 429
rect 942 424 943 428
rect 947 424 948 428
rect 942 423 948 424
rect 966 428 972 429
rect 998 428 1004 429
rect 966 424 967 428
rect 971 424 972 428
rect 966 423 972 424
rect 986 427 992 428
rect 986 423 987 427
rect 991 423 992 427
rect 998 424 999 428
rect 1003 424 1004 428
rect 998 423 1004 424
rect 647 422 651 423
rect 647 417 651 418
rect 671 422 675 423
rect 671 417 675 418
rect 703 422 707 423
rect 703 417 707 418
rect 735 422 739 423
rect 735 417 739 418
rect 767 422 771 423
rect 767 417 771 418
rect 791 422 795 423
rect 791 417 795 418
rect 831 422 835 423
rect 831 417 835 418
rect 839 422 843 423
rect 839 417 843 418
rect 879 422 883 423
rect 879 417 883 418
rect 903 422 907 423
rect 903 417 907 418
rect 911 422 915 423
rect 911 417 915 418
rect 943 422 947 423
rect 943 417 947 418
rect 967 422 971 423
rect 967 417 971 418
rect 975 422 979 423
rect 986 422 992 423
rect 999 422 1003 423
rect 975 417 979 418
rect 646 416 652 417
rect 646 412 647 416
rect 651 412 652 416
rect 646 411 652 412
rect 702 416 708 417
rect 702 412 703 416
rect 707 412 708 416
rect 702 411 708 412
rect 766 416 772 417
rect 766 412 767 416
rect 771 412 772 416
rect 766 411 772 412
rect 830 416 836 417
rect 830 412 831 416
rect 835 412 836 416
rect 830 411 836 412
rect 902 416 908 417
rect 902 412 903 416
rect 907 412 908 416
rect 902 411 908 412
rect 974 416 980 417
rect 974 412 975 416
rect 979 412 980 416
rect 974 411 980 412
rect 338 407 344 408
rect 338 403 339 407
rect 343 403 344 407
rect 338 402 344 403
rect 346 407 352 408
rect 346 403 347 407
rect 351 403 352 407
rect 346 402 352 403
rect 618 407 624 408
rect 618 403 619 407
rect 623 403 624 407
rect 618 402 624 403
rect 340 392 342 402
rect 338 391 344 392
rect 134 390 140 391
rect 134 386 135 390
rect 139 386 140 390
rect 134 385 140 386
rect 158 390 164 391
rect 158 386 159 390
rect 163 386 164 390
rect 158 385 164 386
rect 182 390 188 391
rect 182 386 183 390
rect 187 386 188 390
rect 182 385 188 386
rect 214 390 220 391
rect 214 386 215 390
rect 219 386 220 390
rect 214 385 220 386
rect 270 390 276 391
rect 270 386 271 390
rect 275 386 276 390
rect 270 385 276 386
rect 326 390 332 391
rect 326 386 327 390
rect 331 386 332 390
rect 338 387 339 391
rect 343 387 344 391
rect 338 386 344 387
rect 326 385 332 386
rect 126 383 132 384
rect 126 379 127 383
rect 131 379 132 383
rect 136 379 138 385
rect 160 379 162 385
rect 184 379 186 385
rect 216 379 218 385
rect 272 379 274 385
rect 328 379 330 385
rect 348 380 350 402
rect 738 399 744 400
rect 738 395 739 399
rect 743 395 744 399
rect 738 394 744 395
rect 390 390 396 391
rect 390 386 391 390
rect 395 386 396 390
rect 390 385 396 386
rect 446 390 452 391
rect 446 386 447 390
rect 451 386 452 390
rect 446 385 452 386
rect 502 390 508 391
rect 502 386 503 390
rect 507 386 508 390
rect 502 385 508 386
rect 550 390 556 391
rect 550 386 551 390
rect 555 386 556 390
rect 550 385 556 386
rect 598 390 604 391
rect 598 386 599 390
rect 603 386 604 390
rect 598 385 604 386
rect 646 390 652 391
rect 646 386 647 390
rect 651 386 652 390
rect 646 385 652 386
rect 702 390 708 391
rect 702 386 703 390
rect 707 386 708 390
rect 702 385 708 386
rect 714 387 720 388
rect 346 379 352 380
rect 392 379 394 385
rect 448 379 450 385
rect 504 379 506 385
rect 552 379 554 385
rect 600 379 602 385
rect 648 379 650 385
rect 666 379 672 380
rect 704 379 706 385
rect 714 383 715 387
rect 719 383 720 387
rect 714 382 720 383
rect 111 378 115 379
rect 126 378 132 379
rect 135 378 139 379
rect 111 373 115 374
rect 135 373 139 374
rect 159 378 163 379
rect 159 373 163 374
rect 183 378 187 379
rect 183 373 187 374
rect 207 378 211 379
rect 207 373 211 374
rect 215 378 219 379
rect 215 373 219 374
rect 231 378 235 379
rect 231 373 235 374
rect 255 378 259 379
rect 255 373 259 374
rect 271 378 275 379
rect 271 373 275 374
rect 295 378 299 379
rect 295 373 299 374
rect 327 378 331 379
rect 327 373 331 374
rect 335 378 339 379
rect 346 375 347 379
rect 351 375 352 379
rect 346 374 352 375
rect 375 378 379 379
rect 335 373 339 374
rect 375 373 379 374
rect 391 378 395 379
rect 391 373 395 374
rect 415 378 419 379
rect 415 373 419 374
rect 447 378 451 379
rect 447 373 451 374
rect 455 378 459 379
rect 455 373 459 374
rect 495 378 499 379
rect 495 373 499 374
rect 503 378 507 379
rect 503 373 507 374
rect 535 378 539 379
rect 535 373 539 374
rect 551 378 555 379
rect 551 373 555 374
rect 575 378 579 379
rect 575 373 579 374
rect 599 378 603 379
rect 599 373 603 374
rect 615 378 619 379
rect 615 373 619 374
rect 647 378 651 379
rect 647 373 651 374
rect 655 378 659 379
rect 666 375 667 379
rect 671 375 672 379
rect 666 374 672 375
rect 687 378 691 379
rect 655 373 659 374
rect 112 366 114 373
rect 136 371 138 373
rect 160 371 162 373
rect 184 371 186 373
rect 208 371 210 373
rect 232 371 234 373
rect 256 371 258 373
rect 296 371 298 373
rect 336 371 338 373
rect 376 371 378 373
rect 416 371 418 373
rect 456 371 458 373
rect 496 371 498 373
rect 536 371 538 373
rect 576 371 578 373
rect 616 371 618 373
rect 656 371 658 373
rect 134 370 140 371
rect 134 366 135 370
rect 139 366 140 370
rect 110 365 116 366
rect 134 365 140 366
rect 158 370 164 371
rect 158 366 159 370
rect 163 366 164 370
rect 158 365 164 366
rect 182 370 188 371
rect 182 366 183 370
rect 187 366 188 370
rect 182 365 188 366
rect 206 370 212 371
rect 206 366 207 370
rect 211 366 212 370
rect 206 365 212 366
rect 230 370 236 371
rect 230 366 231 370
rect 235 366 236 370
rect 230 365 236 366
rect 254 370 260 371
rect 254 366 255 370
rect 259 366 260 370
rect 254 365 260 366
rect 294 370 300 371
rect 294 366 295 370
rect 299 366 300 370
rect 294 365 300 366
rect 334 370 340 371
rect 334 366 335 370
rect 339 366 340 370
rect 334 365 340 366
rect 374 370 380 371
rect 374 366 375 370
rect 379 366 380 370
rect 374 365 380 366
rect 414 370 420 371
rect 414 366 415 370
rect 419 366 420 370
rect 414 365 420 366
rect 454 370 460 371
rect 454 366 455 370
rect 459 366 460 370
rect 454 365 460 366
rect 494 370 500 371
rect 494 366 495 370
rect 499 366 500 370
rect 494 365 500 366
rect 534 370 540 371
rect 534 366 535 370
rect 539 366 540 370
rect 534 365 540 366
rect 574 370 580 371
rect 574 366 575 370
rect 579 366 580 370
rect 574 365 580 366
rect 614 370 620 371
rect 614 366 615 370
rect 619 366 620 370
rect 654 370 660 371
rect 614 365 620 366
rect 626 367 632 368
rect 110 361 111 365
rect 115 361 116 365
rect 626 363 627 367
rect 631 363 632 367
rect 654 366 655 370
rect 659 366 660 370
rect 654 365 660 366
rect 626 362 632 363
rect 110 360 116 361
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 110 342 116 343
rect 134 344 140 345
rect 112 339 114 342
rect 134 340 135 344
rect 139 340 140 344
rect 134 339 140 340
rect 158 344 164 345
rect 158 340 159 344
rect 163 340 164 344
rect 158 339 164 340
rect 182 344 188 345
rect 182 340 183 344
rect 187 340 188 344
rect 182 339 188 340
rect 206 344 212 345
rect 206 340 207 344
rect 211 340 212 344
rect 206 339 212 340
rect 230 344 236 345
rect 230 340 231 344
rect 235 340 236 344
rect 230 339 236 340
rect 254 344 260 345
rect 254 340 255 344
rect 259 340 260 344
rect 254 339 260 340
rect 294 344 300 345
rect 294 340 295 344
rect 299 340 300 344
rect 294 339 300 340
rect 334 344 340 345
rect 374 344 380 345
rect 414 344 420 345
rect 334 340 335 344
rect 339 340 340 344
rect 334 339 340 340
rect 346 343 352 344
rect 346 339 347 343
rect 351 339 352 343
rect 374 340 375 344
rect 379 340 380 344
rect 374 339 380 340
rect 406 343 412 344
rect 406 339 407 343
rect 411 339 412 343
rect 414 340 415 344
rect 419 340 420 344
rect 414 339 420 340
rect 454 344 460 345
rect 454 340 455 344
rect 459 340 460 344
rect 454 339 460 340
rect 494 344 500 345
rect 494 340 495 344
rect 499 340 500 344
rect 494 339 500 340
rect 534 344 540 345
rect 534 340 535 344
rect 539 340 540 344
rect 534 339 540 340
rect 574 344 580 345
rect 574 340 575 344
rect 579 340 580 344
rect 574 339 580 340
rect 614 344 620 345
rect 614 340 615 344
rect 619 340 620 344
rect 614 339 620 340
rect 111 338 115 339
rect 111 333 115 334
rect 135 338 139 339
rect 135 333 139 334
rect 159 338 163 339
rect 159 333 163 334
rect 175 338 179 339
rect 175 333 179 334
rect 183 338 187 339
rect 183 333 187 334
rect 199 338 203 339
rect 199 333 203 334
rect 207 338 211 339
rect 207 333 211 334
rect 223 338 227 339
rect 223 333 227 334
rect 231 338 235 339
rect 231 333 235 334
rect 247 338 251 339
rect 247 333 251 334
rect 255 338 259 339
rect 255 333 259 334
rect 279 338 283 339
rect 279 333 283 334
rect 295 338 299 339
rect 295 333 299 334
rect 319 338 323 339
rect 319 333 323 334
rect 335 338 339 339
rect 346 338 352 339
rect 359 338 363 339
rect 335 333 339 334
rect 112 330 114 333
rect 174 332 180 333
rect 110 329 116 330
rect 110 325 111 329
rect 115 325 116 329
rect 174 328 175 332
rect 179 328 180 332
rect 174 327 180 328
rect 198 332 204 333
rect 198 328 199 332
rect 203 328 204 332
rect 198 327 204 328
rect 222 332 228 333
rect 222 328 223 332
rect 227 328 228 332
rect 222 327 228 328
rect 246 332 252 333
rect 246 328 247 332
rect 251 328 252 332
rect 246 327 252 328
rect 278 332 284 333
rect 278 328 279 332
rect 283 328 284 332
rect 278 327 284 328
rect 318 332 324 333
rect 318 328 319 332
rect 323 328 324 332
rect 318 327 324 328
rect 110 324 116 325
rect 210 323 216 324
rect 210 319 211 323
rect 215 319 216 323
rect 210 318 216 319
rect 258 323 264 324
rect 258 319 259 323
rect 263 319 264 323
rect 258 318 264 319
rect 330 323 336 324
rect 330 319 331 323
rect 335 319 336 323
rect 330 318 336 319
rect 187 316 191 317
rect 110 311 116 312
rect 187 311 191 312
rect 110 307 111 311
rect 115 307 116 311
rect 188 308 190 311
rect 212 308 214 318
rect 260 308 262 318
rect 332 308 334 318
rect 348 317 350 338
rect 359 333 363 334
rect 375 338 379 339
rect 375 333 379 334
rect 399 338 403 339
rect 406 338 412 339
rect 415 338 419 339
rect 399 333 403 334
rect 358 332 364 333
rect 358 328 359 332
rect 363 328 364 332
rect 358 327 364 328
rect 398 332 404 333
rect 398 328 399 332
rect 403 328 404 332
rect 398 327 404 328
rect 347 316 351 317
rect 408 315 410 338
rect 415 333 419 334
rect 439 338 443 339
rect 439 333 443 334
rect 455 338 459 339
rect 455 333 459 334
rect 479 338 483 339
rect 479 333 483 334
rect 495 338 499 339
rect 495 333 499 334
rect 527 338 531 339
rect 527 333 531 334
rect 535 338 539 339
rect 535 333 539 334
rect 575 338 579 339
rect 575 333 579 334
rect 583 338 587 339
rect 583 333 587 334
rect 615 338 619 339
rect 615 333 619 334
rect 438 332 444 333
rect 438 328 439 332
rect 443 328 444 332
rect 438 327 444 328
rect 478 332 484 333
rect 478 328 479 332
rect 483 328 484 332
rect 478 327 484 328
rect 526 332 532 333
rect 526 328 527 332
rect 531 328 532 332
rect 526 327 532 328
rect 582 332 588 333
rect 582 328 583 332
rect 587 328 588 332
rect 582 327 588 328
rect 628 324 630 362
rect 668 360 670 374
rect 687 373 691 374
rect 703 378 707 379
rect 703 373 707 374
rect 688 371 690 373
rect 686 370 692 371
rect 686 366 687 370
rect 691 366 692 370
rect 686 365 692 366
rect 666 359 672 360
rect 666 355 667 359
rect 671 355 672 359
rect 666 354 672 355
rect 716 352 718 382
rect 727 378 731 379
rect 727 373 731 374
rect 728 371 730 373
rect 740 372 742 394
rect 988 392 990 422
rect 999 417 1003 418
rect 1024 400 1026 446
rect 1030 428 1036 429
rect 1030 424 1031 428
rect 1035 424 1036 428
rect 1030 423 1036 424
rect 1070 428 1076 429
rect 1070 424 1071 428
rect 1075 424 1076 428
rect 1070 423 1076 424
rect 1118 428 1124 429
rect 1118 424 1119 428
rect 1123 424 1124 428
rect 1118 423 1124 424
rect 1174 428 1180 429
rect 1174 424 1175 428
rect 1179 424 1180 428
rect 1174 423 1180 424
rect 1238 428 1244 429
rect 1302 428 1308 429
rect 1238 424 1239 428
rect 1243 424 1244 428
rect 1238 423 1244 424
rect 1258 427 1264 428
rect 1258 423 1259 427
rect 1263 423 1264 427
rect 1302 424 1303 428
rect 1307 424 1308 428
rect 1302 423 1308 424
rect 1310 423 1316 424
rect 1031 422 1035 423
rect 1031 417 1035 418
rect 1039 422 1043 423
rect 1039 417 1043 418
rect 1071 422 1075 423
rect 1071 417 1075 418
rect 1103 422 1107 423
rect 1103 417 1107 418
rect 1119 422 1123 423
rect 1119 417 1123 418
rect 1159 422 1163 423
rect 1159 417 1163 418
rect 1175 422 1179 423
rect 1175 417 1179 418
rect 1207 422 1211 423
rect 1207 417 1211 418
rect 1239 422 1243 423
rect 1239 417 1243 418
rect 1247 422 1251 423
rect 1258 422 1264 423
rect 1279 422 1283 423
rect 1247 417 1251 418
rect 1038 416 1044 417
rect 1038 412 1039 416
rect 1043 412 1044 416
rect 1038 411 1044 412
rect 1102 416 1108 417
rect 1102 412 1103 416
rect 1107 412 1108 416
rect 1102 411 1108 412
rect 1158 416 1164 417
rect 1158 412 1159 416
rect 1163 412 1164 416
rect 1158 411 1164 412
rect 1206 416 1212 417
rect 1206 412 1207 416
rect 1211 412 1212 416
rect 1206 411 1212 412
rect 1246 416 1252 417
rect 1246 412 1247 416
rect 1251 412 1252 416
rect 1246 411 1252 412
rect 1050 407 1056 408
rect 1050 403 1051 407
rect 1055 403 1056 407
rect 1050 402 1056 403
rect 1238 407 1244 408
rect 1238 403 1239 407
rect 1243 403 1244 407
rect 1238 402 1244 403
rect 1022 399 1028 400
rect 1022 395 1023 399
rect 1027 395 1028 399
rect 1022 394 1028 395
rect 1052 392 1054 402
rect 986 391 992 392
rect 1050 391 1056 392
rect 766 390 772 391
rect 766 386 767 390
rect 771 386 772 390
rect 766 385 772 386
rect 830 390 836 391
rect 830 386 831 390
rect 835 386 836 390
rect 830 385 836 386
rect 902 390 908 391
rect 902 386 903 390
rect 907 386 908 390
rect 902 385 908 386
rect 974 390 980 391
rect 974 386 975 390
rect 979 386 980 390
rect 986 387 987 391
rect 991 387 992 391
rect 986 386 992 387
rect 1038 390 1044 391
rect 1038 386 1039 390
rect 1043 386 1044 390
rect 1050 387 1051 391
rect 1055 387 1056 391
rect 1050 386 1056 387
rect 1102 390 1108 391
rect 1102 386 1103 390
rect 1107 386 1108 390
rect 974 385 980 386
rect 1038 385 1044 386
rect 1102 385 1108 386
rect 1158 390 1164 391
rect 1158 386 1159 390
rect 1163 386 1164 390
rect 1158 385 1164 386
rect 1206 390 1212 391
rect 1206 386 1207 390
rect 1211 386 1212 390
rect 1206 385 1212 386
rect 768 379 770 385
rect 832 379 834 385
rect 904 379 906 385
rect 976 379 978 385
rect 1040 379 1042 385
rect 1104 379 1106 385
rect 1160 379 1162 385
rect 1208 379 1210 385
rect 767 378 771 379
rect 767 373 771 374
rect 775 378 779 379
rect 775 373 779 374
rect 831 378 835 379
rect 831 373 835 374
rect 887 378 891 379
rect 887 373 891 374
rect 903 378 907 379
rect 903 373 907 374
rect 951 378 955 379
rect 951 373 955 374
rect 975 378 979 379
rect 975 373 979 374
rect 1015 378 1019 379
rect 1015 373 1019 374
rect 1039 378 1043 379
rect 1039 373 1043 374
rect 1079 378 1083 379
rect 1079 373 1083 374
rect 1103 378 1107 379
rect 1103 373 1107 374
rect 1135 378 1139 379
rect 1135 373 1139 374
rect 1159 378 1163 379
rect 1159 373 1163 374
rect 1183 378 1187 379
rect 1183 373 1187 374
rect 1207 378 1211 379
rect 1207 373 1211 374
rect 1231 378 1235 379
rect 1240 376 1242 402
rect 1246 390 1252 391
rect 1246 386 1247 390
rect 1251 386 1252 390
rect 1246 385 1252 386
rect 1248 379 1250 385
rect 1260 384 1262 422
rect 1279 417 1283 418
rect 1303 422 1307 423
rect 1310 419 1311 423
rect 1315 419 1316 423
rect 1310 418 1316 419
rect 1319 422 1323 423
rect 1303 417 1307 418
rect 1278 416 1284 417
rect 1278 412 1279 416
rect 1283 412 1284 416
rect 1278 411 1284 412
rect 1312 392 1314 418
rect 1319 417 1323 418
rect 1318 416 1324 417
rect 1332 416 1334 446
rect 1446 445 1447 449
rect 1451 445 1452 449
rect 1446 444 1452 445
rect 1446 431 1452 432
rect 1366 428 1372 429
rect 1366 424 1367 428
rect 1371 424 1372 428
rect 1366 423 1372 424
rect 1414 428 1420 429
rect 1414 424 1415 428
rect 1419 424 1420 428
rect 1414 423 1420 424
rect 1426 427 1432 428
rect 1426 423 1427 427
rect 1431 423 1432 427
rect 1446 427 1447 431
rect 1451 427 1452 431
rect 1446 426 1452 427
rect 1448 423 1450 426
rect 1359 422 1363 423
rect 1359 417 1363 418
rect 1367 422 1371 423
rect 1367 417 1371 418
rect 1391 422 1395 423
rect 1391 417 1395 418
rect 1415 422 1419 423
rect 1426 422 1432 423
rect 1447 422 1451 423
rect 1415 417 1419 418
rect 1358 416 1364 417
rect 1318 412 1319 416
rect 1323 412 1324 416
rect 1318 411 1324 412
rect 1330 415 1336 416
rect 1330 411 1331 415
rect 1335 411 1336 415
rect 1358 412 1359 416
rect 1363 412 1364 416
rect 1358 411 1364 412
rect 1390 416 1396 417
rect 1390 412 1391 416
rect 1395 412 1396 416
rect 1390 411 1396 412
rect 1414 416 1420 417
rect 1414 412 1415 416
rect 1419 412 1420 416
rect 1414 411 1420 412
rect 1330 410 1336 411
rect 1428 392 1430 422
rect 1447 417 1451 418
rect 1448 414 1450 417
rect 1446 413 1452 414
rect 1446 409 1447 413
rect 1451 409 1452 413
rect 1446 408 1452 409
rect 1446 395 1452 396
rect 1310 391 1316 392
rect 1426 391 1432 392
rect 1278 390 1284 391
rect 1278 386 1279 390
rect 1283 386 1284 390
rect 1310 387 1311 391
rect 1315 387 1316 391
rect 1310 386 1316 387
rect 1318 390 1324 391
rect 1318 386 1319 390
rect 1323 386 1324 390
rect 1278 385 1284 386
rect 1318 385 1324 386
rect 1358 390 1364 391
rect 1358 386 1359 390
rect 1363 386 1364 390
rect 1358 385 1364 386
rect 1390 390 1396 391
rect 1390 386 1391 390
rect 1395 386 1396 390
rect 1390 385 1396 386
rect 1414 390 1420 391
rect 1414 386 1415 390
rect 1419 386 1420 390
rect 1426 387 1427 391
rect 1431 387 1432 391
rect 1446 391 1447 395
rect 1451 391 1452 395
rect 1446 390 1452 391
rect 1426 386 1432 387
rect 1414 385 1420 386
rect 1258 383 1264 384
rect 1258 379 1259 383
rect 1263 379 1264 383
rect 1280 379 1282 385
rect 1320 379 1322 385
rect 1360 379 1362 385
rect 1382 383 1388 384
rect 1382 379 1383 383
rect 1387 379 1388 383
rect 1392 379 1394 385
rect 1416 379 1418 385
rect 1448 379 1450 390
rect 1247 378 1251 379
rect 1258 378 1264 379
rect 1271 378 1275 379
rect 1231 373 1235 374
rect 1238 375 1244 376
rect 738 371 744 372
rect 776 371 778 373
rect 832 371 834 373
rect 888 371 890 373
rect 952 371 954 373
rect 1016 371 1018 373
rect 1080 371 1082 373
rect 1136 371 1138 373
rect 1184 371 1186 373
rect 1232 371 1234 373
rect 1238 371 1239 375
rect 1243 371 1244 375
rect 1247 373 1251 374
rect 1271 373 1275 374
rect 1279 378 1283 379
rect 1279 373 1283 374
rect 1311 378 1315 379
rect 1311 373 1315 374
rect 1319 378 1323 379
rect 1319 373 1323 374
rect 1351 378 1355 379
rect 1351 373 1355 374
rect 1359 378 1363 379
rect 1382 378 1388 379
rect 1391 378 1395 379
rect 1359 373 1363 374
rect 1272 371 1274 373
rect 1312 371 1314 373
rect 1352 371 1354 373
rect 726 370 732 371
rect 726 366 727 370
rect 731 366 732 370
rect 738 367 739 371
rect 743 367 744 371
rect 738 366 744 367
rect 774 370 780 371
rect 774 366 775 370
rect 779 366 780 370
rect 726 365 732 366
rect 774 365 780 366
rect 830 370 836 371
rect 830 366 831 370
rect 835 366 836 370
rect 830 365 836 366
rect 886 370 892 371
rect 886 366 887 370
rect 891 366 892 370
rect 886 365 892 366
rect 950 370 956 371
rect 950 366 951 370
rect 955 366 956 370
rect 950 365 956 366
rect 1014 370 1020 371
rect 1014 366 1015 370
rect 1019 366 1020 370
rect 1078 370 1084 371
rect 1014 365 1020 366
rect 1026 367 1032 368
rect 1026 363 1027 367
rect 1031 363 1032 367
rect 1078 366 1079 370
rect 1083 366 1084 370
rect 1078 365 1084 366
rect 1134 370 1140 371
rect 1134 366 1135 370
rect 1139 366 1140 370
rect 1134 365 1140 366
rect 1182 370 1188 371
rect 1182 366 1183 370
rect 1187 366 1188 370
rect 1182 365 1188 366
rect 1230 370 1236 371
rect 1238 370 1244 371
rect 1270 370 1276 371
rect 1230 366 1231 370
rect 1235 366 1236 370
rect 1230 365 1236 366
rect 1270 366 1271 370
rect 1275 366 1276 370
rect 1310 370 1316 371
rect 1270 365 1276 366
rect 1290 367 1296 368
rect 1026 362 1032 363
rect 1290 363 1291 367
rect 1295 363 1296 367
rect 1310 366 1311 370
rect 1315 366 1316 370
rect 1310 365 1316 366
rect 1350 370 1356 371
rect 1350 366 1351 370
rect 1355 366 1356 370
rect 1350 365 1356 366
rect 1290 362 1296 363
rect 714 351 720 352
rect 714 347 715 351
rect 719 347 720 351
rect 714 346 720 347
rect 654 344 660 345
rect 654 340 655 344
rect 659 340 660 344
rect 654 339 660 340
rect 686 344 692 345
rect 686 340 687 344
rect 691 340 692 344
rect 686 339 692 340
rect 726 344 732 345
rect 726 340 727 344
rect 731 340 732 344
rect 726 339 732 340
rect 774 344 780 345
rect 774 340 775 344
rect 779 340 780 344
rect 774 339 780 340
rect 830 344 836 345
rect 830 340 831 344
rect 835 340 836 344
rect 830 339 836 340
rect 886 344 892 345
rect 886 340 887 344
rect 891 340 892 344
rect 886 339 892 340
rect 950 344 956 345
rect 950 340 951 344
rect 955 340 956 344
rect 950 339 956 340
rect 1014 344 1020 345
rect 1014 340 1015 344
rect 1019 340 1020 344
rect 1014 339 1020 340
rect 639 338 643 339
rect 639 333 643 334
rect 655 338 659 339
rect 655 333 659 334
rect 687 338 691 339
rect 687 333 691 334
rect 727 338 731 339
rect 727 333 731 334
rect 735 338 739 339
rect 735 333 739 334
rect 775 338 779 339
rect 775 333 779 334
rect 791 338 795 339
rect 791 333 795 334
rect 831 338 835 339
rect 831 333 835 334
rect 847 338 851 339
rect 847 333 851 334
rect 887 338 891 339
rect 887 333 891 334
rect 895 338 899 339
rect 895 333 899 334
rect 943 338 947 339
rect 943 333 947 334
rect 951 338 955 339
rect 951 333 955 334
rect 991 338 995 339
rect 991 333 995 334
rect 1015 338 1019 339
rect 1015 333 1019 334
rect 638 332 644 333
rect 638 328 639 332
rect 643 328 644 332
rect 638 327 644 328
rect 686 332 692 333
rect 686 328 687 332
rect 691 328 692 332
rect 686 327 692 328
rect 734 332 740 333
rect 734 328 735 332
rect 739 328 740 332
rect 734 327 740 328
rect 790 332 796 333
rect 790 328 791 332
rect 795 328 796 332
rect 790 327 796 328
rect 846 332 852 333
rect 846 328 847 332
rect 851 328 852 332
rect 846 327 852 328
rect 894 332 900 333
rect 894 328 895 332
rect 899 328 900 332
rect 894 327 900 328
rect 942 332 948 333
rect 942 328 943 332
rect 947 328 948 332
rect 942 327 948 328
rect 990 332 996 333
rect 990 328 991 332
rect 995 328 996 332
rect 990 327 996 328
rect 1028 324 1030 362
rect 1078 344 1084 345
rect 1078 340 1079 344
rect 1083 340 1084 344
rect 1078 339 1084 340
rect 1134 344 1140 345
rect 1134 340 1135 344
rect 1139 340 1140 344
rect 1134 339 1140 340
rect 1182 344 1188 345
rect 1182 340 1183 344
rect 1187 340 1188 344
rect 1182 339 1188 340
rect 1230 344 1236 345
rect 1230 340 1231 344
rect 1235 340 1236 344
rect 1230 339 1236 340
rect 1270 344 1276 345
rect 1270 340 1271 344
rect 1275 340 1276 344
rect 1270 339 1276 340
rect 1039 338 1043 339
rect 1039 333 1043 334
rect 1079 338 1083 339
rect 1079 333 1083 334
rect 1087 338 1091 339
rect 1087 333 1091 334
rect 1135 338 1139 339
rect 1135 333 1139 334
rect 1183 338 1187 339
rect 1183 333 1187 334
rect 1231 338 1235 339
rect 1231 333 1235 334
rect 1271 338 1275 339
rect 1271 333 1275 334
rect 1279 338 1283 339
rect 1279 333 1283 334
rect 1038 332 1044 333
rect 1038 328 1039 332
rect 1043 328 1044 332
rect 1038 327 1044 328
rect 1086 332 1092 333
rect 1086 328 1087 332
rect 1091 328 1092 332
rect 1086 327 1092 328
rect 1134 332 1140 333
rect 1134 328 1135 332
rect 1139 328 1140 332
rect 1134 327 1140 328
rect 1182 332 1188 333
rect 1182 328 1183 332
rect 1187 328 1188 332
rect 1182 327 1188 328
rect 1230 332 1236 333
rect 1230 328 1231 332
rect 1235 328 1236 332
rect 1230 327 1236 328
rect 1278 332 1284 333
rect 1292 332 1294 362
rect 1384 352 1386 378
rect 1391 373 1395 374
rect 1415 378 1419 379
rect 1415 373 1419 374
rect 1447 378 1451 379
rect 1447 373 1451 374
rect 1392 371 1394 373
rect 1416 371 1418 373
rect 1390 370 1396 371
rect 1390 366 1391 370
rect 1395 366 1396 370
rect 1390 365 1396 366
rect 1414 370 1420 371
rect 1414 366 1415 370
rect 1419 366 1420 370
rect 1448 366 1450 373
rect 1414 365 1420 366
rect 1446 365 1452 366
rect 1446 361 1447 365
rect 1451 361 1452 365
rect 1446 360 1452 361
rect 1382 351 1388 352
rect 1382 347 1383 351
rect 1387 347 1388 351
rect 1382 346 1388 347
rect 1446 347 1452 348
rect 1310 344 1316 345
rect 1310 340 1311 344
rect 1315 340 1316 344
rect 1310 339 1316 340
rect 1350 344 1356 345
rect 1350 340 1351 344
rect 1355 340 1356 344
rect 1350 339 1356 340
rect 1390 344 1396 345
rect 1414 344 1420 345
rect 1390 340 1391 344
rect 1395 340 1396 344
rect 1390 339 1396 340
rect 1402 343 1408 344
rect 1402 339 1403 343
rect 1407 339 1408 343
rect 1414 340 1415 344
rect 1419 340 1420 344
rect 1446 343 1447 347
rect 1451 343 1452 347
rect 1446 342 1452 343
rect 1414 339 1420 340
rect 1448 339 1450 342
rect 1311 338 1315 339
rect 1311 333 1315 334
rect 1327 338 1331 339
rect 1327 333 1331 334
rect 1351 338 1355 339
rect 1351 333 1355 334
rect 1383 338 1387 339
rect 1383 333 1387 334
rect 1391 338 1395 339
rect 1402 338 1408 339
rect 1415 338 1419 339
rect 1391 333 1395 334
rect 1326 332 1332 333
rect 1278 328 1279 332
rect 1283 328 1284 332
rect 1278 327 1284 328
rect 1290 331 1296 332
rect 1290 327 1291 331
rect 1295 327 1296 331
rect 1326 328 1327 332
rect 1331 328 1332 332
rect 1326 327 1332 328
rect 1382 332 1388 333
rect 1382 328 1383 332
rect 1387 328 1388 332
rect 1382 327 1388 328
rect 1290 326 1296 327
rect 450 323 456 324
rect 450 319 451 323
rect 455 319 456 323
rect 450 318 456 319
rect 626 323 632 324
rect 626 319 627 323
rect 631 319 632 323
rect 626 318 632 319
rect 1026 323 1032 324
rect 1026 319 1027 323
rect 1031 319 1032 323
rect 1026 318 1032 319
rect 1258 323 1264 324
rect 1258 319 1259 323
rect 1263 319 1264 323
rect 1258 318 1264 319
rect 408 313 414 315
rect 347 311 351 312
rect 412 308 414 313
rect 452 308 454 318
rect 518 315 524 316
rect 518 311 519 315
rect 523 311 524 315
rect 518 310 524 311
rect 183 307 190 308
rect 210 307 216 308
rect 258 307 264 308
rect 330 307 336 308
rect 410 307 416 308
rect 450 307 456 308
rect 110 306 116 307
rect 174 306 180 307
rect 112 299 114 306
rect 174 302 175 306
rect 179 302 180 306
rect 183 303 184 307
rect 188 304 190 307
rect 198 306 204 307
rect 188 303 189 304
rect 183 302 189 303
rect 198 302 199 306
rect 203 302 204 306
rect 210 303 211 307
rect 215 303 216 307
rect 210 302 216 303
rect 222 306 228 307
rect 222 302 223 306
rect 227 302 228 306
rect 174 301 180 302
rect 198 301 204 302
rect 222 301 228 302
rect 246 306 252 307
rect 246 302 247 306
rect 251 302 252 306
rect 258 303 259 307
rect 263 303 264 307
rect 258 302 264 303
rect 278 306 284 307
rect 278 302 279 306
rect 283 302 284 306
rect 246 301 252 302
rect 278 301 284 302
rect 318 306 324 307
rect 318 302 319 306
rect 323 302 324 306
rect 330 303 331 307
rect 335 303 336 307
rect 330 302 336 303
rect 358 306 364 307
rect 358 302 359 306
rect 363 302 364 306
rect 318 301 324 302
rect 358 301 364 302
rect 398 306 404 307
rect 398 302 399 306
rect 403 302 404 306
rect 410 303 411 307
rect 415 303 416 307
rect 410 302 416 303
rect 438 306 444 307
rect 438 302 439 306
rect 443 302 444 306
rect 450 303 451 307
rect 455 303 456 307
rect 450 302 456 303
rect 478 306 484 307
rect 478 302 479 306
rect 483 302 484 306
rect 398 301 404 302
rect 438 301 444 302
rect 478 301 484 302
rect 176 299 178 301
rect 200 299 202 301
rect 224 299 226 301
rect 248 299 250 301
rect 280 299 282 301
rect 320 299 322 301
rect 360 299 362 301
rect 400 299 402 301
rect 440 299 442 301
rect 480 299 482 301
rect 111 298 115 299
rect 111 293 115 294
rect 175 298 179 299
rect 175 293 179 294
rect 199 298 203 299
rect 199 293 203 294
rect 223 298 227 299
rect 223 293 227 294
rect 247 298 251 299
rect 247 293 251 294
rect 271 298 275 299
rect 271 293 275 294
rect 279 298 283 299
rect 279 293 283 294
rect 295 298 299 299
rect 295 293 299 294
rect 319 298 323 299
rect 319 293 323 294
rect 343 298 347 299
rect 343 293 347 294
rect 359 298 363 299
rect 359 293 363 294
rect 367 298 371 299
rect 367 293 371 294
rect 399 298 403 299
rect 399 293 403 294
rect 431 298 435 299
rect 431 293 435 294
rect 439 298 443 299
rect 439 293 443 294
rect 471 298 475 299
rect 471 293 475 294
rect 479 298 483 299
rect 479 293 483 294
rect 511 298 515 299
rect 520 296 522 310
rect 526 306 532 307
rect 526 302 527 306
rect 531 302 532 306
rect 526 301 532 302
rect 582 306 588 307
rect 582 302 583 306
rect 587 302 588 306
rect 582 301 588 302
rect 638 306 644 307
rect 638 302 639 306
rect 643 302 644 306
rect 638 301 644 302
rect 686 306 692 307
rect 686 302 687 306
rect 691 302 692 306
rect 686 301 692 302
rect 734 306 740 307
rect 734 302 735 306
rect 739 302 740 306
rect 734 301 740 302
rect 790 306 796 307
rect 790 302 791 306
rect 795 302 796 306
rect 790 301 796 302
rect 846 306 852 307
rect 846 302 847 306
rect 851 302 852 306
rect 846 301 852 302
rect 894 306 900 307
rect 894 302 895 306
rect 899 302 900 306
rect 894 301 900 302
rect 942 306 948 307
rect 942 302 943 306
rect 947 302 948 306
rect 942 301 948 302
rect 990 306 996 307
rect 990 302 991 306
rect 995 302 996 306
rect 990 301 996 302
rect 1038 306 1044 307
rect 1038 302 1039 306
rect 1043 302 1044 306
rect 1038 301 1044 302
rect 1086 306 1092 307
rect 1086 302 1087 306
rect 1091 302 1092 306
rect 1086 301 1092 302
rect 1134 306 1140 307
rect 1134 302 1135 306
rect 1139 302 1140 306
rect 1134 301 1140 302
rect 1182 306 1188 307
rect 1182 302 1183 306
rect 1187 302 1188 306
rect 1182 301 1188 302
rect 1230 306 1236 307
rect 1230 302 1231 306
rect 1235 302 1236 306
rect 1230 301 1236 302
rect 528 299 530 301
rect 570 299 576 300
rect 584 299 586 301
rect 640 299 642 301
rect 688 299 690 301
rect 736 299 738 301
rect 770 299 776 300
rect 792 299 794 301
rect 848 299 850 301
rect 896 299 898 301
rect 944 299 946 301
rect 992 299 994 301
rect 1040 299 1042 301
rect 1088 299 1090 301
rect 1136 299 1138 301
rect 1184 299 1186 301
rect 1232 299 1234 301
rect 527 298 531 299
rect 511 293 515 294
rect 518 295 524 296
rect 112 286 114 293
rect 248 291 250 293
rect 272 291 274 293
rect 296 291 298 293
rect 320 291 322 293
rect 344 291 346 293
rect 368 291 370 293
rect 400 291 402 293
rect 432 291 434 293
rect 472 291 474 293
rect 512 291 514 293
rect 518 291 519 295
rect 523 291 524 295
rect 527 293 531 294
rect 559 298 563 299
rect 570 295 571 299
rect 575 295 576 299
rect 570 294 576 295
rect 583 298 587 299
rect 559 293 563 294
rect 560 291 562 293
rect 246 290 252 291
rect 246 286 247 290
rect 251 286 252 290
rect 110 285 116 286
rect 246 285 252 286
rect 270 290 276 291
rect 270 286 271 290
rect 275 286 276 290
rect 270 285 276 286
rect 294 290 300 291
rect 294 286 295 290
rect 299 286 300 290
rect 318 290 324 291
rect 306 287 312 288
rect 306 286 307 287
rect 294 285 300 286
rect 110 281 111 285
rect 115 281 116 285
rect 304 283 307 286
rect 311 283 312 287
rect 318 286 319 290
rect 323 286 324 290
rect 318 285 324 286
rect 342 290 348 291
rect 342 286 343 290
rect 347 286 348 290
rect 342 285 348 286
rect 366 290 372 291
rect 366 286 367 290
rect 371 286 372 290
rect 366 285 372 286
rect 398 290 404 291
rect 398 286 399 290
rect 403 286 404 290
rect 398 285 404 286
rect 430 290 436 291
rect 430 286 431 290
rect 435 286 436 290
rect 430 285 436 286
rect 470 290 476 291
rect 470 286 471 290
rect 475 286 476 290
rect 470 285 476 286
rect 510 290 516 291
rect 518 290 524 291
rect 558 290 564 291
rect 510 286 511 290
rect 515 286 516 290
rect 510 285 516 286
rect 558 286 559 290
rect 563 286 564 290
rect 558 285 564 286
rect 110 280 116 281
rect 296 282 312 283
rect 296 281 306 282
rect 296 276 298 281
rect 572 280 574 294
rect 583 293 587 294
rect 615 298 619 299
rect 615 293 619 294
rect 639 298 643 299
rect 639 293 643 294
rect 663 298 667 299
rect 663 293 667 294
rect 687 298 691 299
rect 687 293 691 294
rect 711 298 715 299
rect 711 293 715 294
rect 735 298 739 299
rect 735 293 739 294
rect 759 298 763 299
rect 770 295 771 299
rect 775 295 776 299
rect 770 294 776 295
rect 791 298 795 299
rect 759 293 763 294
rect 616 291 618 293
rect 664 291 666 293
rect 712 291 714 293
rect 760 291 762 293
rect 614 290 620 291
rect 614 286 615 290
rect 619 286 620 290
rect 614 285 620 286
rect 662 290 668 291
rect 662 286 663 290
rect 667 286 668 290
rect 662 285 668 286
rect 710 290 716 291
rect 710 286 711 290
rect 715 286 716 290
rect 758 290 764 291
rect 710 285 716 286
rect 722 287 728 288
rect 722 283 723 287
rect 727 283 728 287
rect 758 286 759 290
rect 763 286 764 290
rect 758 285 764 286
rect 722 282 728 283
rect 570 279 576 280
rect 294 275 300 276
rect 294 271 295 275
rect 299 271 300 275
rect 294 270 300 271
rect 418 275 424 276
rect 418 271 419 275
rect 423 271 424 275
rect 570 275 571 279
rect 575 275 576 279
rect 570 274 576 275
rect 418 270 424 271
rect 279 268 283 269
rect 411 268 415 269
rect 110 267 116 268
rect 110 263 111 267
rect 115 263 116 267
rect 110 262 116 263
rect 246 264 252 265
rect 112 259 114 262
rect 246 260 247 264
rect 251 260 252 264
rect 246 259 252 260
rect 270 264 276 265
rect 270 260 271 264
rect 275 260 276 264
rect 279 263 283 264
rect 294 264 300 265
rect 270 259 276 260
rect 111 258 115 259
rect 111 253 115 254
rect 247 258 251 259
rect 247 253 251 254
rect 263 258 267 259
rect 263 253 267 254
rect 271 258 275 259
rect 271 253 275 254
rect 112 250 114 253
rect 262 252 268 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 262 248 263 252
rect 267 248 268 252
rect 262 247 268 248
rect 110 244 116 245
rect 110 231 116 232
rect 110 227 111 231
rect 115 227 116 231
rect 280 228 282 263
rect 294 260 295 264
rect 299 260 300 264
rect 294 259 300 260
rect 318 264 324 265
rect 318 260 319 264
rect 323 260 324 264
rect 318 259 324 260
rect 342 264 348 265
rect 342 260 343 264
rect 347 260 348 264
rect 342 259 348 260
rect 366 264 372 265
rect 366 260 367 264
rect 371 260 372 264
rect 366 259 372 260
rect 398 264 404 265
rect 398 260 399 264
rect 403 260 404 264
rect 410 263 411 268
rect 415 263 416 268
rect 410 262 416 263
rect 398 259 404 260
rect 287 258 291 259
rect 287 253 291 254
rect 295 258 299 259
rect 295 253 299 254
rect 311 258 315 259
rect 311 253 315 254
rect 319 258 323 259
rect 319 253 323 254
rect 335 258 339 259
rect 335 253 339 254
rect 343 258 347 259
rect 343 253 347 254
rect 359 258 363 259
rect 359 253 363 254
rect 367 258 371 259
rect 367 253 371 254
rect 383 258 387 259
rect 383 253 387 254
rect 399 258 403 259
rect 399 253 403 254
rect 407 258 411 259
rect 407 253 411 254
rect 286 252 292 253
rect 286 248 287 252
rect 291 248 292 252
rect 286 247 292 248
rect 310 252 316 253
rect 310 248 311 252
rect 315 248 316 252
rect 310 247 316 248
rect 334 252 340 253
rect 334 248 335 252
rect 339 248 340 252
rect 334 247 340 248
rect 358 252 364 253
rect 358 248 359 252
rect 363 248 364 252
rect 358 247 364 248
rect 382 252 388 253
rect 382 248 383 252
rect 387 248 388 252
rect 382 247 388 248
rect 406 252 412 253
rect 406 248 407 252
rect 411 248 412 252
rect 406 247 412 248
rect 322 243 328 244
rect 322 239 323 243
rect 327 239 328 243
rect 322 238 328 239
rect 346 243 352 244
rect 346 239 347 243
rect 351 239 352 243
rect 394 243 400 244
rect 346 238 352 239
rect 358 239 364 240
rect 324 228 326 238
rect 348 228 350 238
rect 358 235 359 239
rect 363 235 364 239
rect 394 239 395 243
rect 399 239 400 243
rect 394 238 400 239
rect 358 234 370 235
rect 360 233 370 234
rect 274 227 282 228
rect 322 227 328 228
rect 346 227 352 228
rect 110 226 116 227
rect 262 226 268 227
rect 112 219 114 226
rect 262 222 263 226
rect 267 222 268 226
rect 274 223 275 227
rect 279 224 282 227
rect 286 226 292 227
rect 279 223 280 224
rect 274 222 280 223
rect 286 222 287 226
rect 291 222 292 226
rect 262 221 268 222
rect 286 221 292 222
rect 310 226 316 227
rect 310 222 311 226
rect 315 222 316 226
rect 322 223 323 227
rect 327 223 328 227
rect 322 222 328 223
rect 334 226 340 227
rect 334 222 335 226
rect 339 222 340 226
rect 346 223 347 227
rect 351 223 352 227
rect 346 222 352 223
rect 358 226 364 227
rect 358 222 359 226
rect 363 222 364 226
rect 310 221 316 222
rect 334 221 340 222
rect 358 221 364 222
rect 264 219 266 221
rect 288 219 290 221
rect 312 219 314 221
rect 336 219 338 221
rect 360 219 362 221
rect 368 220 370 233
rect 382 226 388 227
rect 382 222 383 226
rect 387 222 388 226
rect 382 221 388 222
rect 366 219 372 220
rect 384 219 386 221
rect 111 218 115 219
rect 111 213 115 214
rect 239 218 243 219
rect 239 213 243 214
rect 263 218 267 219
rect 263 213 267 214
rect 287 218 291 219
rect 287 213 291 214
rect 311 218 315 219
rect 311 213 315 214
rect 335 218 339 219
rect 335 213 339 214
rect 359 218 363 219
rect 366 215 367 219
rect 371 215 372 219
rect 366 214 372 215
rect 383 218 387 219
rect 359 213 363 214
rect 383 213 387 214
rect 112 206 114 213
rect 240 211 242 213
rect 264 211 266 213
rect 288 211 290 213
rect 312 211 314 213
rect 336 211 338 213
rect 360 211 362 213
rect 384 211 386 213
rect 396 212 398 238
rect 420 228 422 270
rect 430 264 436 265
rect 430 260 431 264
rect 435 260 436 264
rect 430 259 436 260
rect 470 264 476 265
rect 470 260 471 264
rect 475 260 476 264
rect 470 259 476 260
rect 510 264 516 265
rect 510 260 511 264
rect 515 260 516 264
rect 510 259 516 260
rect 558 264 564 265
rect 558 260 559 264
rect 563 260 564 264
rect 558 259 564 260
rect 614 264 620 265
rect 614 260 615 264
rect 619 260 620 264
rect 614 259 620 260
rect 662 264 668 265
rect 662 260 663 264
rect 667 260 668 264
rect 662 259 668 260
rect 710 264 716 265
rect 710 260 711 264
rect 715 260 716 264
rect 710 259 716 260
rect 431 258 435 259
rect 431 253 435 254
rect 463 258 467 259
rect 463 253 467 254
rect 471 258 475 259
rect 471 253 475 254
rect 503 258 507 259
rect 503 253 507 254
rect 511 258 515 259
rect 511 253 515 254
rect 543 258 547 259
rect 543 253 547 254
rect 559 258 563 259
rect 559 253 563 254
rect 583 258 587 259
rect 583 253 587 254
rect 615 258 619 259
rect 615 253 619 254
rect 623 258 627 259
rect 623 253 627 254
rect 663 258 667 259
rect 663 253 667 254
rect 679 258 683 259
rect 679 253 683 254
rect 711 258 715 259
rect 711 253 715 254
rect 430 252 436 253
rect 430 248 431 252
rect 435 248 436 252
rect 430 247 436 248
rect 462 252 468 253
rect 462 248 463 252
rect 467 248 468 252
rect 462 247 468 248
rect 502 252 508 253
rect 502 248 503 252
rect 507 248 508 252
rect 502 247 508 248
rect 542 252 548 253
rect 542 248 543 252
rect 547 248 548 252
rect 542 247 548 248
rect 582 252 588 253
rect 582 248 583 252
rect 587 248 588 252
rect 582 247 588 248
rect 622 252 628 253
rect 622 248 623 252
rect 627 248 628 252
rect 622 247 628 248
rect 678 252 684 253
rect 678 248 679 252
rect 683 248 684 252
rect 678 247 684 248
rect 724 244 726 282
rect 772 280 774 294
rect 791 293 795 294
rect 807 298 811 299
rect 807 293 811 294
rect 847 298 851 299
rect 847 293 851 294
rect 879 298 883 299
rect 879 293 883 294
rect 895 298 899 299
rect 895 293 899 294
rect 903 298 907 299
rect 903 293 907 294
rect 927 298 931 299
rect 927 293 931 294
rect 943 298 947 299
rect 943 293 947 294
rect 951 298 955 299
rect 951 293 955 294
rect 975 298 979 299
rect 975 293 979 294
rect 991 298 995 299
rect 991 293 995 294
rect 999 298 1003 299
rect 999 293 1003 294
rect 1023 298 1027 299
rect 1023 293 1027 294
rect 1039 298 1043 299
rect 1039 293 1043 294
rect 1047 298 1051 299
rect 1047 293 1051 294
rect 1071 298 1075 299
rect 1071 293 1075 294
rect 1087 298 1091 299
rect 1087 293 1091 294
rect 1095 298 1099 299
rect 1095 293 1099 294
rect 1127 298 1131 299
rect 1127 293 1131 294
rect 1135 298 1139 299
rect 1135 293 1139 294
rect 1159 298 1163 299
rect 1159 293 1163 294
rect 1183 298 1187 299
rect 1183 293 1187 294
rect 1199 298 1203 299
rect 1199 293 1203 294
rect 1231 298 1235 299
rect 1231 293 1235 294
rect 1247 298 1251 299
rect 1247 293 1251 294
rect 808 291 810 293
rect 848 291 850 293
rect 880 291 882 293
rect 904 291 906 293
rect 928 291 930 293
rect 952 291 954 293
rect 976 291 978 293
rect 1000 291 1002 293
rect 1024 291 1026 293
rect 1048 291 1050 293
rect 1072 291 1074 293
rect 1096 291 1098 293
rect 1128 291 1130 293
rect 1160 291 1162 293
rect 1200 291 1202 293
rect 1248 291 1250 293
rect 1260 292 1262 318
rect 1404 308 1406 338
rect 1415 333 1419 334
rect 1447 338 1451 339
rect 1447 333 1451 334
rect 1414 332 1420 333
rect 1414 328 1415 332
rect 1419 328 1420 332
rect 1448 330 1450 333
rect 1414 327 1420 328
rect 1446 329 1452 330
rect 1446 325 1447 329
rect 1451 325 1452 329
rect 1446 324 1452 325
rect 1426 315 1432 316
rect 1426 311 1427 315
rect 1431 311 1432 315
rect 1426 310 1432 311
rect 1446 311 1452 312
rect 1402 307 1408 308
rect 1278 306 1284 307
rect 1278 302 1279 306
rect 1283 302 1284 306
rect 1278 301 1284 302
rect 1326 306 1332 307
rect 1326 302 1327 306
rect 1331 302 1332 306
rect 1382 306 1388 307
rect 1326 301 1332 302
rect 1374 303 1380 304
rect 1280 299 1282 301
rect 1328 299 1330 301
rect 1374 299 1375 303
rect 1379 299 1380 303
rect 1382 302 1383 306
rect 1387 302 1388 306
rect 1402 303 1403 307
rect 1407 303 1408 307
rect 1402 302 1408 303
rect 1414 306 1420 307
rect 1414 302 1415 306
rect 1419 302 1420 306
rect 1382 301 1388 302
rect 1414 301 1420 302
rect 1384 299 1386 301
rect 1416 299 1418 301
rect 1279 298 1283 299
rect 1279 293 1283 294
rect 1303 298 1307 299
rect 1303 293 1307 294
rect 1327 298 1331 299
rect 1327 293 1331 294
rect 1367 298 1371 299
rect 1374 298 1380 299
rect 1383 298 1387 299
rect 1367 293 1371 294
rect 1258 291 1264 292
rect 1304 291 1306 293
rect 1368 291 1370 293
rect 806 290 812 291
rect 806 286 807 290
rect 811 286 812 290
rect 806 285 812 286
rect 846 290 852 291
rect 846 286 847 290
rect 851 286 852 290
rect 846 285 852 286
rect 878 290 884 291
rect 878 286 879 290
rect 883 286 884 290
rect 878 285 884 286
rect 902 290 908 291
rect 902 286 903 290
rect 907 286 908 290
rect 902 285 908 286
rect 926 290 932 291
rect 926 286 927 290
rect 931 286 932 290
rect 926 285 932 286
rect 950 290 956 291
rect 950 286 951 290
rect 955 286 956 290
rect 950 285 956 286
rect 974 290 980 291
rect 974 286 975 290
rect 979 286 980 290
rect 974 285 980 286
rect 998 290 1004 291
rect 998 286 999 290
rect 1003 286 1004 290
rect 998 285 1004 286
rect 1022 290 1028 291
rect 1022 286 1023 290
rect 1027 286 1028 290
rect 1022 285 1028 286
rect 1046 290 1052 291
rect 1046 286 1047 290
rect 1051 286 1052 290
rect 1046 285 1052 286
rect 1070 290 1076 291
rect 1070 286 1071 290
rect 1075 286 1076 290
rect 1070 285 1076 286
rect 1094 290 1100 291
rect 1094 286 1095 290
rect 1099 286 1100 290
rect 1094 285 1100 286
rect 1126 290 1132 291
rect 1126 286 1127 290
rect 1131 286 1132 290
rect 1126 285 1132 286
rect 1158 290 1164 291
rect 1158 286 1159 290
rect 1163 286 1164 290
rect 1158 285 1164 286
rect 1198 290 1204 291
rect 1198 286 1199 290
rect 1203 286 1204 290
rect 1198 285 1204 286
rect 1246 290 1252 291
rect 1246 286 1247 290
rect 1251 286 1252 290
rect 1258 287 1259 291
rect 1263 287 1264 291
rect 1258 286 1264 287
rect 1302 290 1308 291
rect 1302 286 1303 290
rect 1307 286 1308 290
rect 1366 290 1372 291
rect 1246 285 1252 286
rect 1302 285 1308 286
rect 1314 287 1320 288
rect 1314 283 1315 287
rect 1319 283 1320 287
rect 1366 286 1367 290
rect 1371 286 1372 290
rect 1366 285 1372 286
rect 1314 282 1320 283
rect 770 279 776 280
rect 770 275 771 279
rect 775 275 776 279
rect 770 274 776 275
rect 758 264 764 265
rect 758 260 759 264
rect 763 260 764 264
rect 758 259 764 260
rect 806 264 812 265
rect 806 260 807 264
rect 811 260 812 264
rect 806 259 812 260
rect 846 264 852 265
rect 846 260 847 264
rect 851 260 852 264
rect 846 259 852 260
rect 878 264 884 265
rect 878 260 879 264
rect 883 260 884 264
rect 878 259 884 260
rect 902 264 908 265
rect 902 260 903 264
rect 907 260 908 264
rect 902 259 908 260
rect 926 264 932 265
rect 926 260 927 264
rect 931 260 932 264
rect 926 259 932 260
rect 950 264 956 265
rect 950 260 951 264
rect 955 260 956 264
rect 950 259 956 260
rect 974 264 980 265
rect 974 260 975 264
rect 979 260 980 264
rect 974 259 980 260
rect 998 264 1004 265
rect 998 260 999 264
rect 1003 260 1004 264
rect 998 259 1004 260
rect 1022 264 1028 265
rect 1022 260 1023 264
rect 1027 260 1028 264
rect 1022 259 1028 260
rect 1046 264 1052 265
rect 1046 260 1047 264
rect 1051 260 1052 264
rect 1046 259 1052 260
rect 1070 264 1076 265
rect 1070 260 1071 264
rect 1075 260 1076 264
rect 1070 259 1076 260
rect 1094 264 1100 265
rect 1094 260 1095 264
rect 1099 260 1100 264
rect 1094 259 1100 260
rect 1126 264 1132 265
rect 1126 260 1127 264
rect 1131 260 1132 264
rect 1126 259 1132 260
rect 1158 264 1164 265
rect 1158 260 1159 264
rect 1163 260 1164 264
rect 1158 259 1164 260
rect 1198 264 1204 265
rect 1198 260 1199 264
rect 1203 260 1204 264
rect 1198 259 1204 260
rect 1246 264 1252 265
rect 1246 260 1247 264
rect 1251 260 1252 264
rect 1246 259 1252 260
rect 1302 264 1308 265
rect 1302 260 1303 264
rect 1307 260 1308 264
rect 1302 259 1308 260
rect 743 258 747 259
rect 743 253 747 254
rect 759 258 763 259
rect 759 253 763 254
rect 807 258 811 259
rect 807 253 811 254
rect 847 258 851 259
rect 847 253 851 254
rect 879 258 883 259
rect 879 253 883 254
rect 903 258 907 259
rect 903 253 907 254
rect 927 258 931 259
rect 927 253 931 254
rect 951 258 955 259
rect 951 253 955 254
rect 959 258 963 259
rect 959 253 963 254
rect 975 258 979 259
rect 975 253 979 254
rect 999 258 1003 259
rect 999 253 1003 254
rect 1023 258 1027 259
rect 1023 253 1027 254
rect 1039 258 1043 259
rect 1039 253 1043 254
rect 1047 258 1051 259
rect 1047 253 1051 254
rect 1071 258 1075 259
rect 1071 253 1075 254
rect 1095 258 1099 259
rect 1095 253 1099 254
rect 1119 258 1123 259
rect 1119 253 1123 254
rect 1127 258 1131 259
rect 1127 253 1131 254
rect 1159 258 1163 259
rect 1159 253 1163 254
rect 1199 258 1203 259
rect 1199 253 1203 254
rect 1247 258 1251 259
rect 1247 253 1251 254
rect 1279 258 1283 259
rect 1279 253 1283 254
rect 1303 258 1307 259
rect 1303 253 1307 254
rect 742 252 748 253
rect 742 248 743 252
rect 747 248 748 252
rect 742 247 748 248
rect 806 252 812 253
rect 806 248 807 252
rect 811 248 812 252
rect 806 247 812 248
rect 878 252 884 253
rect 878 248 879 252
rect 883 248 884 252
rect 878 247 884 248
rect 958 252 964 253
rect 958 248 959 252
rect 963 248 964 252
rect 958 247 964 248
rect 1038 252 1044 253
rect 1038 248 1039 252
rect 1043 248 1044 252
rect 1038 247 1044 248
rect 1118 252 1124 253
rect 1118 248 1119 252
rect 1123 248 1124 252
rect 1118 247 1124 248
rect 1198 252 1204 253
rect 1198 248 1199 252
rect 1203 248 1204 252
rect 1198 247 1204 248
rect 1278 252 1284 253
rect 1316 252 1318 282
rect 1376 268 1378 298
rect 1383 293 1387 294
rect 1415 298 1419 299
rect 1415 293 1419 294
rect 1416 291 1418 293
rect 1428 292 1430 310
rect 1446 307 1447 311
rect 1451 307 1452 311
rect 1446 306 1452 307
rect 1448 299 1450 306
rect 1447 298 1451 299
rect 1447 293 1451 294
rect 1426 291 1432 292
rect 1414 290 1420 291
rect 1414 286 1415 290
rect 1419 286 1420 290
rect 1426 287 1427 291
rect 1431 287 1432 291
rect 1426 286 1432 287
rect 1448 286 1450 293
rect 1414 285 1420 286
rect 1446 285 1452 286
rect 1446 281 1447 285
rect 1451 281 1452 285
rect 1446 280 1452 281
rect 1376 267 1384 268
rect 1376 265 1379 267
rect 1366 264 1372 265
rect 1366 260 1367 264
rect 1371 260 1372 264
rect 1378 263 1379 265
rect 1383 263 1384 267
rect 1446 267 1452 268
rect 1378 262 1384 263
rect 1414 264 1420 265
rect 1366 259 1372 260
rect 1414 260 1415 264
rect 1419 260 1420 264
rect 1446 263 1447 267
rect 1451 263 1452 267
rect 1446 262 1452 263
rect 1414 259 1420 260
rect 1448 259 1450 262
rect 1359 258 1363 259
rect 1359 253 1363 254
rect 1367 258 1371 259
rect 1367 253 1371 254
rect 1415 258 1419 259
rect 1415 253 1419 254
rect 1447 258 1451 259
rect 1447 253 1451 254
rect 1358 252 1364 253
rect 1278 248 1279 252
rect 1283 248 1284 252
rect 1278 247 1284 248
rect 1314 251 1320 252
rect 1314 247 1315 251
rect 1319 247 1320 251
rect 1358 248 1359 252
rect 1363 248 1364 252
rect 1358 247 1364 248
rect 1414 252 1420 253
rect 1414 248 1415 252
rect 1419 248 1420 252
rect 1448 250 1450 253
rect 1414 247 1420 248
rect 1446 249 1452 250
rect 1314 246 1320 247
rect 1446 245 1447 249
rect 1451 245 1452 249
rect 1446 244 1452 245
rect 474 243 480 244
rect 474 239 475 243
rect 479 239 480 243
rect 474 238 480 239
rect 554 243 560 244
rect 554 239 555 243
rect 559 239 560 243
rect 722 243 728 244
rect 554 238 560 239
rect 590 239 596 240
rect 476 228 478 238
rect 556 228 558 238
rect 590 235 591 239
rect 595 235 596 239
rect 722 239 723 243
rect 727 239 728 243
rect 722 238 728 239
rect 1130 243 1136 244
rect 1130 239 1131 243
rect 1135 239 1136 243
rect 1130 238 1136 239
rect 590 234 596 235
rect 418 227 424 228
rect 474 227 480 228
rect 554 227 560 228
rect 406 226 412 227
rect 406 222 407 226
rect 411 222 412 226
rect 418 223 419 227
rect 423 223 424 227
rect 418 222 424 223
rect 430 226 436 227
rect 430 222 431 226
rect 435 222 436 226
rect 406 221 412 222
rect 430 221 436 222
rect 462 226 468 227
rect 462 222 463 226
rect 467 222 468 226
rect 474 223 475 227
rect 479 223 480 227
rect 474 222 480 223
rect 502 226 508 227
rect 502 222 503 226
rect 507 222 508 226
rect 462 221 468 222
rect 502 221 508 222
rect 542 226 548 227
rect 542 222 543 226
rect 547 222 548 226
rect 554 223 555 227
rect 559 223 560 227
rect 554 222 560 223
rect 582 226 588 227
rect 582 222 583 226
rect 587 222 588 226
rect 542 221 548 222
rect 582 221 588 222
rect 408 219 410 221
rect 432 219 434 221
rect 464 219 466 221
rect 504 219 506 221
rect 544 219 546 221
rect 584 219 586 221
rect 407 218 411 219
rect 407 213 411 214
rect 431 218 435 219
rect 431 213 435 214
rect 463 218 467 219
rect 463 213 467 214
rect 503 218 507 219
rect 503 213 507 214
rect 511 218 515 219
rect 511 213 515 214
rect 543 218 547 219
rect 543 213 547 214
rect 559 218 563 219
rect 559 213 563 214
rect 583 218 587 219
rect 583 213 587 214
rect 394 211 400 212
rect 408 211 410 213
rect 432 211 434 213
rect 464 211 466 213
rect 512 211 514 213
rect 560 211 562 213
rect 238 210 244 211
rect 238 206 239 210
rect 243 206 244 210
rect 110 205 116 206
rect 238 205 244 206
rect 262 210 268 211
rect 262 206 263 210
rect 267 206 268 210
rect 262 205 268 206
rect 286 210 292 211
rect 286 206 287 210
rect 291 206 292 210
rect 286 205 292 206
rect 310 210 316 211
rect 310 206 311 210
rect 315 206 316 210
rect 310 205 316 206
rect 334 210 340 211
rect 334 206 335 210
rect 339 206 340 210
rect 334 205 340 206
rect 358 210 364 211
rect 358 206 359 210
rect 363 206 364 210
rect 358 205 364 206
rect 382 210 388 211
rect 382 206 383 210
rect 387 206 388 210
rect 394 207 395 211
rect 399 207 400 211
rect 394 206 400 207
rect 406 210 412 211
rect 406 206 407 210
rect 411 206 412 210
rect 430 210 436 211
rect 382 205 388 206
rect 406 205 412 206
rect 418 207 424 208
rect 110 201 111 205
rect 115 201 116 205
rect 418 202 419 207
rect 110 200 116 201
rect 423 202 424 207
rect 430 206 431 210
rect 435 206 436 210
rect 430 205 436 206
rect 462 210 468 211
rect 462 206 463 210
rect 467 206 468 210
rect 462 205 468 206
rect 510 210 516 211
rect 510 206 511 210
rect 515 206 516 210
rect 510 205 516 206
rect 558 210 564 211
rect 558 206 559 210
rect 563 206 564 210
rect 558 205 564 206
rect 592 205 594 234
rect 1132 228 1134 238
rect 1426 235 1432 236
rect 1426 231 1427 235
rect 1431 231 1432 235
rect 1426 230 1432 231
rect 1446 231 1452 232
rect 1130 227 1136 228
rect 622 226 628 227
rect 622 222 623 226
rect 627 222 628 226
rect 622 221 628 222
rect 678 226 684 227
rect 678 222 679 226
rect 683 222 684 226
rect 678 221 684 222
rect 742 226 748 227
rect 742 222 743 226
rect 747 222 748 226
rect 742 221 748 222
rect 806 226 812 227
rect 806 222 807 226
rect 811 222 812 226
rect 806 221 812 222
rect 878 226 884 227
rect 878 222 879 226
rect 883 222 884 226
rect 878 221 884 222
rect 958 226 964 227
rect 958 222 959 226
rect 963 222 964 226
rect 958 221 964 222
rect 1038 226 1044 227
rect 1038 222 1039 226
rect 1043 222 1044 226
rect 1118 226 1124 227
rect 1038 221 1044 222
rect 1094 223 1100 224
rect 624 219 626 221
rect 680 219 682 221
rect 730 219 736 220
rect 744 219 746 221
rect 808 219 810 221
rect 880 219 882 221
rect 960 219 962 221
rect 1040 219 1042 221
rect 1094 219 1095 223
rect 1099 219 1100 223
rect 1118 222 1119 226
rect 1123 222 1124 226
rect 1130 223 1131 227
rect 1135 223 1136 227
rect 1130 222 1136 223
rect 1198 226 1204 227
rect 1198 222 1199 226
rect 1203 222 1204 226
rect 1118 221 1124 222
rect 1198 221 1204 222
rect 1278 226 1284 227
rect 1278 222 1279 226
rect 1283 222 1284 226
rect 1278 221 1284 222
rect 1358 226 1364 227
rect 1358 222 1359 226
rect 1363 222 1364 226
rect 1358 221 1364 222
rect 1414 226 1420 227
rect 1414 222 1415 226
rect 1419 222 1420 226
rect 1414 221 1420 222
rect 1120 219 1122 221
rect 1200 219 1202 221
rect 1280 219 1282 221
rect 1360 219 1362 221
rect 1416 219 1418 221
rect 615 218 619 219
rect 615 213 619 214
rect 623 218 627 219
rect 623 213 627 214
rect 671 218 675 219
rect 671 213 675 214
rect 679 218 683 219
rect 679 213 683 214
rect 719 218 723 219
rect 730 215 731 219
rect 735 215 736 219
rect 730 214 736 215
rect 743 218 747 219
rect 719 213 723 214
rect 616 211 618 213
rect 672 211 674 213
rect 720 211 722 213
rect 614 210 620 211
rect 614 206 615 210
rect 619 206 620 210
rect 614 205 620 206
rect 670 210 676 211
rect 670 206 671 210
rect 675 206 676 210
rect 670 205 676 206
rect 718 210 724 211
rect 718 206 719 210
rect 723 206 724 210
rect 718 205 724 206
rect 591 204 595 205
rect 419 199 423 200
rect 732 200 734 214
rect 743 213 747 214
rect 767 218 771 219
rect 767 213 771 214
rect 807 218 811 219
rect 807 213 811 214
rect 815 218 819 219
rect 815 213 819 214
rect 863 218 867 219
rect 863 213 867 214
rect 879 218 883 219
rect 879 213 883 214
rect 919 218 923 219
rect 919 213 923 214
rect 959 218 963 219
rect 959 213 963 214
rect 975 218 979 219
rect 975 213 979 214
rect 1031 218 1035 219
rect 1031 213 1035 214
rect 1039 218 1043 219
rect 1039 213 1043 214
rect 1087 218 1091 219
rect 1094 218 1100 219
rect 1119 218 1123 219
rect 1087 213 1091 214
rect 768 211 770 213
rect 816 211 818 213
rect 864 211 866 213
rect 920 211 922 213
rect 976 211 978 213
rect 1032 211 1034 213
rect 1088 211 1090 213
rect 766 210 772 211
rect 766 206 767 210
rect 771 206 772 210
rect 766 205 772 206
rect 814 210 820 211
rect 814 206 815 210
rect 819 206 820 210
rect 814 205 820 206
rect 862 210 868 211
rect 862 206 863 210
rect 867 206 868 210
rect 862 205 868 206
rect 918 210 924 211
rect 918 206 919 210
rect 923 206 924 210
rect 918 205 924 206
rect 974 210 980 211
rect 974 206 975 210
rect 979 206 980 210
rect 974 205 980 206
rect 1030 210 1036 211
rect 1030 206 1031 210
rect 1035 206 1036 210
rect 1030 205 1036 206
rect 1086 210 1092 211
rect 1086 206 1087 210
rect 1091 206 1092 210
rect 1086 205 1092 206
rect 1096 200 1098 218
rect 1119 213 1123 214
rect 1135 218 1139 219
rect 1135 213 1139 214
rect 1183 218 1187 219
rect 1183 213 1187 214
rect 1199 218 1203 219
rect 1199 213 1203 214
rect 1231 218 1235 219
rect 1231 213 1235 214
rect 1279 218 1283 219
rect 1279 213 1283 214
rect 1327 218 1331 219
rect 1327 213 1331 214
rect 1359 218 1363 219
rect 1359 213 1363 214
rect 1383 218 1387 219
rect 1383 213 1387 214
rect 1415 218 1419 219
rect 1415 213 1419 214
rect 1136 211 1138 213
rect 1184 211 1186 213
rect 1232 211 1234 213
rect 1280 211 1282 213
rect 1328 211 1330 213
rect 1384 211 1386 213
rect 1416 211 1418 213
rect 1428 212 1430 230
rect 1446 227 1447 231
rect 1451 227 1452 231
rect 1446 226 1452 227
rect 1448 219 1450 226
rect 1447 218 1451 219
rect 1447 213 1451 214
rect 1426 211 1432 212
rect 1134 210 1140 211
rect 1134 206 1135 210
rect 1139 206 1140 210
rect 1134 205 1140 206
rect 1182 210 1188 211
rect 1182 206 1183 210
rect 1187 206 1188 210
rect 1230 210 1236 211
rect 1182 205 1188 206
rect 1194 207 1200 208
rect 1194 203 1195 207
rect 1199 203 1200 207
rect 1230 206 1231 210
rect 1235 206 1236 210
rect 1230 205 1236 206
rect 1278 210 1284 211
rect 1278 206 1279 210
rect 1283 206 1284 210
rect 1278 205 1284 206
rect 1326 210 1332 211
rect 1326 206 1327 210
rect 1331 206 1332 210
rect 1326 205 1332 206
rect 1382 210 1388 211
rect 1382 206 1383 210
rect 1387 206 1388 210
rect 1382 205 1388 206
rect 1414 210 1420 211
rect 1414 206 1415 210
rect 1419 206 1420 210
rect 1426 207 1427 211
rect 1431 207 1432 211
rect 1426 206 1432 207
rect 1448 206 1450 213
rect 1414 205 1420 206
rect 1446 205 1452 206
rect 1194 202 1200 203
rect 591 199 595 200
rect 730 199 736 200
rect 730 195 731 199
rect 735 195 736 199
rect 730 194 736 195
rect 1094 199 1100 200
rect 1094 195 1095 199
rect 1099 195 1100 199
rect 1094 194 1100 195
rect 110 187 116 188
rect 110 183 111 187
rect 115 183 116 187
rect 110 182 116 183
rect 238 184 244 185
rect 262 184 268 185
rect 112 179 114 182
rect 238 180 239 184
rect 243 180 244 184
rect 238 179 244 180
rect 250 183 256 184
rect 250 179 251 183
rect 255 179 256 183
rect 262 180 263 184
rect 267 180 268 184
rect 262 179 268 180
rect 286 184 292 185
rect 286 180 287 184
rect 291 180 292 184
rect 286 179 292 180
rect 310 184 316 185
rect 310 180 311 184
rect 315 180 316 184
rect 310 179 316 180
rect 334 184 340 185
rect 334 180 335 184
rect 339 180 340 184
rect 334 179 340 180
rect 358 184 364 185
rect 358 180 359 184
rect 363 180 364 184
rect 358 179 364 180
rect 382 184 388 185
rect 382 180 383 184
rect 387 180 388 184
rect 382 179 388 180
rect 406 184 412 185
rect 406 180 407 184
rect 411 180 412 184
rect 406 179 412 180
rect 430 184 436 185
rect 430 180 431 184
rect 435 180 436 184
rect 430 179 436 180
rect 462 184 468 185
rect 462 180 463 184
rect 467 180 468 184
rect 462 179 468 180
rect 510 184 516 185
rect 510 180 511 184
rect 515 180 516 184
rect 510 179 516 180
rect 558 184 564 185
rect 558 180 559 184
rect 563 180 564 184
rect 558 179 564 180
rect 614 184 620 185
rect 614 180 615 184
rect 619 180 620 184
rect 614 179 620 180
rect 670 184 676 185
rect 718 184 724 185
rect 670 180 671 184
rect 675 180 676 184
rect 670 179 676 180
rect 682 183 688 184
rect 682 179 683 183
rect 687 179 688 183
rect 718 180 719 184
rect 723 180 724 184
rect 718 179 724 180
rect 766 184 772 185
rect 766 180 767 184
rect 771 180 772 184
rect 766 179 772 180
rect 814 184 820 185
rect 814 180 815 184
rect 819 180 820 184
rect 814 179 820 180
rect 862 184 868 185
rect 862 180 863 184
rect 867 180 868 184
rect 862 179 868 180
rect 918 184 924 185
rect 918 180 919 184
rect 923 180 924 184
rect 918 179 924 180
rect 974 184 980 185
rect 974 180 975 184
rect 979 180 980 184
rect 974 179 980 180
rect 1030 184 1036 185
rect 1030 180 1031 184
rect 1035 180 1036 184
rect 1030 179 1036 180
rect 1086 184 1092 185
rect 1086 180 1087 184
rect 1091 180 1092 184
rect 1086 179 1092 180
rect 1134 184 1140 185
rect 1134 180 1135 184
rect 1139 180 1140 184
rect 1134 179 1140 180
rect 1182 184 1188 185
rect 1182 180 1183 184
rect 1187 180 1188 184
rect 1182 179 1188 180
rect 111 178 115 179
rect 111 173 115 174
rect 183 178 187 179
rect 183 173 187 174
rect 207 178 211 179
rect 207 173 211 174
rect 239 178 243 179
rect 250 178 256 179
rect 263 178 267 179
rect 239 173 243 174
rect 112 170 114 173
rect 182 172 188 173
rect 110 169 116 170
rect 110 165 111 169
rect 115 165 116 169
rect 182 168 183 172
rect 187 168 188 172
rect 182 167 188 168
rect 206 172 212 173
rect 206 168 207 172
rect 211 168 212 172
rect 206 167 212 168
rect 238 172 244 173
rect 238 168 239 172
rect 243 168 244 172
rect 238 167 244 168
rect 110 164 116 165
rect 110 151 116 152
rect 110 147 111 151
rect 115 147 116 151
rect 110 146 116 147
rect 182 146 188 147
rect 112 127 114 146
rect 182 142 183 146
rect 187 142 188 146
rect 182 141 188 142
rect 206 146 212 147
rect 206 142 207 146
rect 211 142 212 146
rect 206 141 212 142
rect 238 146 244 147
rect 238 142 239 146
rect 243 142 244 146
rect 238 141 244 142
rect 184 127 186 141
rect 208 127 210 141
rect 240 127 242 141
rect 252 140 254 178
rect 263 173 267 174
rect 279 178 283 179
rect 279 173 283 174
rect 287 178 291 179
rect 287 173 291 174
rect 311 178 315 179
rect 311 173 315 174
rect 327 178 331 179
rect 327 173 331 174
rect 335 178 339 179
rect 335 173 339 174
rect 359 178 363 179
rect 359 173 363 174
rect 375 178 379 179
rect 375 173 379 174
rect 383 178 387 179
rect 383 173 387 174
rect 407 178 411 179
rect 407 173 411 174
rect 423 178 427 179
rect 423 173 427 174
rect 431 178 435 179
rect 431 173 435 174
rect 463 178 467 179
rect 463 173 467 174
rect 471 178 475 179
rect 471 173 475 174
rect 511 178 515 179
rect 511 173 515 174
rect 527 178 531 179
rect 527 173 531 174
rect 559 178 563 179
rect 559 173 563 174
rect 591 178 595 179
rect 591 173 595 174
rect 615 178 619 179
rect 615 173 619 174
rect 655 178 659 179
rect 655 173 659 174
rect 671 178 675 179
rect 682 178 688 179
rect 711 178 715 179
rect 671 173 675 174
rect 278 172 284 173
rect 278 168 279 172
rect 283 168 284 172
rect 278 167 284 168
rect 326 172 332 173
rect 326 168 327 172
rect 331 168 332 172
rect 326 167 332 168
rect 374 172 380 173
rect 374 168 375 172
rect 379 168 380 172
rect 374 167 380 168
rect 422 172 428 173
rect 422 168 423 172
rect 427 168 428 172
rect 422 167 428 168
rect 470 172 476 173
rect 470 168 471 172
rect 475 168 476 172
rect 470 167 476 168
rect 526 172 532 173
rect 526 168 527 172
rect 531 168 532 172
rect 526 167 532 168
rect 590 172 596 173
rect 590 168 591 172
rect 595 168 596 172
rect 590 167 596 168
rect 654 172 660 173
rect 654 168 655 172
rect 659 168 660 172
rect 654 167 660 168
rect 410 163 416 164
rect 410 159 411 163
rect 415 159 416 163
rect 410 158 416 159
rect 482 163 488 164
rect 482 159 483 163
rect 487 159 488 163
rect 482 158 488 159
rect 602 163 608 164
rect 602 159 603 163
rect 607 159 608 163
rect 602 158 608 159
rect 278 146 284 147
rect 278 142 279 146
rect 283 142 284 146
rect 278 141 284 142
rect 326 146 332 147
rect 326 142 327 146
rect 331 142 332 146
rect 326 141 332 142
rect 374 146 380 147
rect 374 142 375 146
rect 379 142 380 146
rect 374 141 380 142
rect 250 139 256 140
rect 250 135 251 139
rect 255 135 256 139
rect 250 134 256 135
rect 280 127 282 141
rect 328 127 330 141
rect 376 127 378 141
rect 111 126 115 127
rect 111 121 115 122
rect 135 126 139 127
rect 135 121 139 122
rect 159 126 163 127
rect 159 121 163 122
rect 183 126 187 127
rect 183 121 187 122
rect 207 126 211 127
rect 207 121 211 122
rect 231 126 235 127
rect 231 121 235 122
rect 239 126 243 127
rect 239 121 243 122
rect 255 126 259 127
rect 255 121 259 122
rect 279 126 283 127
rect 279 121 283 122
rect 303 126 307 127
rect 303 121 307 122
rect 327 126 331 127
rect 327 121 331 122
rect 351 126 355 127
rect 351 121 355 122
rect 375 126 379 127
rect 375 121 379 122
rect 399 126 403 127
rect 399 121 403 122
rect 112 114 114 121
rect 136 119 138 121
rect 160 119 162 121
rect 184 119 186 121
rect 208 119 210 121
rect 232 119 234 121
rect 256 119 258 121
rect 280 119 282 121
rect 304 119 306 121
rect 328 119 330 121
rect 352 119 354 121
rect 376 119 378 121
rect 400 119 402 121
rect 412 120 414 158
rect 484 148 486 158
rect 604 148 606 158
rect 670 155 676 156
rect 670 151 671 155
rect 675 151 676 155
rect 670 150 676 151
rect 482 147 488 148
rect 602 147 608 148
rect 422 146 428 147
rect 422 142 423 146
rect 427 142 428 146
rect 422 141 428 142
rect 470 146 476 147
rect 470 142 471 146
rect 475 142 476 146
rect 482 143 483 147
rect 487 143 488 147
rect 482 142 488 143
rect 526 146 532 147
rect 526 142 527 146
rect 531 142 532 146
rect 470 141 476 142
rect 526 141 532 142
rect 590 146 596 147
rect 590 142 591 146
rect 595 142 596 146
rect 602 143 603 147
rect 607 143 608 147
rect 602 142 608 143
rect 654 146 660 147
rect 654 142 655 146
rect 659 142 660 146
rect 590 141 596 142
rect 654 141 660 142
rect 424 127 426 141
rect 472 127 474 141
rect 528 127 530 141
rect 592 127 594 141
rect 656 127 658 141
rect 672 128 674 150
rect 684 136 686 178
rect 711 173 715 174
rect 719 178 723 179
rect 719 173 723 174
rect 767 178 771 179
rect 767 173 771 174
rect 815 178 819 179
rect 815 173 819 174
rect 823 178 827 179
rect 823 173 827 174
rect 863 178 867 179
rect 863 173 867 174
rect 871 178 875 179
rect 871 173 875 174
rect 919 178 923 179
rect 919 173 923 174
rect 975 178 979 179
rect 975 173 979 174
rect 1031 178 1035 179
rect 1031 173 1035 174
rect 1079 178 1083 179
rect 1079 173 1083 174
rect 1087 178 1091 179
rect 1087 173 1091 174
rect 1127 178 1131 179
rect 1127 173 1131 174
rect 1135 178 1139 179
rect 1135 173 1139 174
rect 1175 178 1179 179
rect 1175 173 1179 174
rect 1183 178 1187 179
rect 1183 173 1187 174
rect 710 172 716 173
rect 710 168 711 172
rect 715 168 716 172
rect 710 167 716 168
rect 766 172 772 173
rect 766 168 767 172
rect 771 168 772 172
rect 766 167 772 168
rect 822 172 828 173
rect 822 168 823 172
rect 827 168 828 172
rect 822 167 828 168
rect 870 172 876 173
rect 870 168 871 172
rect 875 168 876 172
rect 870 167 876 168
rect 918 172 924 173
rect 918 168 919 172
rect 923 168 924 172
rect 918 167 924 168
rect 974 172 980 173
rect 974 168 975 172
rect 979 168 980 172
rect 974 167 980 168
rect 1030 172 1036 173
rect 1030 168 1031 172
rect 1035 168 1036 172
rect 1030 167 1036 168
rect 1078 172 1084 173
rect 1078 168 1079 172
rect 1083 168 1084 172
rect 1078 167 1084 168
rect 1126 172 1132 173
rect 1126 168 1127 172
rect 1131 168 1132 172
rect 1126 167 1132 168
rect 1174 172 1180 173
rect 1174 168 1175 172
rect 1179 168 1180 172
rect 1174 167 1180 168
rect 1196 164 1198 202
rect 1446 201 1447 205
rect 1451 201 1452 205
rect 1446 200 1452 201
rect 1370 199 1376 200
rect 1370 195 1371 199
rect 1375 195 1376 199
rect 1370 194 1376 195
rect 1230 184 1236 185
rect 1278 184 1284 185
rect 1230 180 1231 184
rect 1235 180 1236 184
rect 1230 179 1236 180
rect 1270 183 1276 184
rect 1270 179 1271 183
rect 1275 179 1276 183
rect 1278 180 1279 184
rect 1283 180 1284 184
rect 1278 179 1284 180
rect 1326 184 1332 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1223 178 1227 179
rect 1223 173 1227 174
rect 1231 178 1235 179
rect 1231 173 1235 174
rect 1263 178 1267 179
rect 1270 178 1276 179
rect 1279 178 1283 179
rect 1263 173 1267 174
rect 1222 172 1228 173
rect 1222 168 1223 172
rect 1227 168 1228 172
rect 1222 167 1228 168
rect 1262 172 1268 173
rect 1262 168 1263 172
rect 1267 168 1268 172
rect 1262 167 1268 168
rect 722 163 728 164
rect 722 159 723 163
rect 727 159 728 163
rect 722 158 728 159
rect 882 163 888 164
rect 882 159 883 163
rect 887 159 888 163
rect 882 158 888 159
rect 986 163 992 164
rect 986 159 987 163
rect 991 159 992 163
rect 986 158 992 159
rect 1090 163 1096 164
rect 1090 159 1091 163
rect 1095 159 1096 163
rect 1090 158 1096 159
rect 1194 163 1200 164
rect 1194 159 1195 163
rect 1199 159 1200 163
rect 1194 158 1200 159
rect 724 148 726 158
rect 884 148 886 158
rect 988 148 990 158
rect 1092 148 1094 158
rect 722 147 728 148
rect 882 147 888 148
rect 986 147 992 148
rect 1090 147 1096 148
rect 710 146 716 147
rect 710 142 711 146
rect 715 142 716 146
rect 722 143 723 147
rect 727 143 728 147
rect 722 142 728 143
rect 766 146 772 147
rect 766 142 767 146
rect 771 142 772 146
rect 710 141 716 142
rect 766 141 772 142
rect 822 146 828 147
rect 822 142 823 146
rect 827 142 828 146
rect 822 141 828 142
rect 870 146 876 147
rect 870 142 871 146
rect 875 142 876 146
rect 882 143 883 147
rect 887 143 888 147
rect 882 142 888 143
rect 918 146 924 147
rect 918 142 919 146
rect 923 142 924 146
rect 870 141 876 142
rect 918 141 924 142
rect 974 146 980 147
rect 974 142 975 146
rect 979 142 980 146
rect 986 143 987 147
rect 991 143 992 147
rect 986 142 992 143
rect 1030 146 1036 147
rect 1030 142 1031 146
rect 1035 142 1036 146
rect 974 141 980 142
rect 1030 141 1036 142
rect 1078 146 1084 147
rect 1078 142 1079 146
rect 1083 142 1084 146
rect 1090 143 1091 147
rect 1095 143 1096 147
rect 1090 142 1096 143
rect 1126 146 1132 147
rect 1126 142 1127 146
rect 1131 142 1132 146
rect 1078 141 1084 142
rect 1126 141 1132 142
rect 1174 146 1180 147
rect 1174 142 1175 146
rect 1179 142 1180 146
rect 1174 141 1180 142
rect 1222 146 1228 147
rect 1222 142 1223 146
rect 1227 142 1228 146
rect 1222 141 1228 142
rect 1262 146 1268 147
rect 1262 142 1263 146
rect 1267 142 1268 146
rect 1262 141 1268 142
rect 682 135 688 136
rect 682 131 683 135
rect 687 131 688 135
rect 682 130 688 131
rect 670 127 676 128
rect 712 127 714 141
rect 768 127 770 141
rect 824 127 826 141
rect 872 127 874 141
rect 920 127 922 141
rect 976 127 978 141
rect 1022 135 1028 136
rect 1022 131 1023 135
rect 1027 131 1028 135
rect 1022 130 1028 131
rect 423 126 427 127
rect 423 121 427 122
rect 431 126 435 127
rect 431 121 435 122
rect 463 126 467 127
rect 463 121 467 122
rect 471 126 475 127
rect 471 121 475 122
rect 487 126 491 127
rect 487 121 491 122
rect 511 126 515 127
rect 511 121 515 122
rect 527 126 531 127
rect 527 121 531 122
rect 535 126 539 127
rect 535 121 539 122
rect 559 126 563 127
rect 559 121 563 122
rect 583 126 587 127
rect 583 121 587 122
rect 591 126 595 127
rect 591 121 595 122
rect 607 126 611 127
rect 607 121 611 122
rect 631 126 635 127
rect 631 121 635 122
rect 655 126 659 127
rect 670 123 671 127
rect 675 123 676 127
rect 670 122 676 123
rect 679 126 683 127
rect 655 121 659 122
rect 679 121 683 122
rect 703 126 707 127
rect 703 121 707 122
rect 711 126 715 127
rect 711 121 715 122
rect 727 126 731 127
rect 727 121 731 122
rect 751 126 755 127
rect 751 121 755 122
rect 767 126 771 127
rect 767 121 771 122
rect 775 126 779 127
rect 775 121 779 122
rect 799 126 803 127
rect 799 121 803 122
rect 823 126 827 127
rect 823 121 827 122
rect 855 126 859 127
rect 855 121 859 122
rect 871 126 875 127
rect 871 121 875 122
rect 887 126 891 127
rect 887 121 891 122
rect 919 126 923 127
rect 919 121 923 122
rect 951 126 955 127
rect 951 121 955 122
rect 975 126 979 127
rect 975 121 979 122
rect 983 126 987 127
rect 983 121 987 122
rect 1015 126 1019 127
rect 1015 121 1019 122
rect 410 119 416 120
rect 432 119 434 121
rect 464 119 466 121
rect 488 119 490 121
rect 512 119 514 121
rect 536 119 538 121
rect 560 119 562 121
rect 584 119 586 121
rect 608 119 610 121
rect 632 119 634 121
rect 656 119 658 121
rect 680 119 682 121
rect 704 119 706 121
rect 728 119 730 121
rect 752 119 754 121
rect 776 119 778 121
rect 800 119 802 121
rect 824 119 826 121
rect 856 119 858 121
rect 888 119 890 121
rect 920 119 922 121
rect 952 119 954 121
rect 984 119 986 121
rect 1016 119 1018 121
rect 134 118 140 119
rect 134 114 135 118
rect 139 114 140 118
rect 110 113 116 114
rect 134 113 140 114
rect 158 118 164 119
rect 158 114 159 118
rect 163 114 164 118
rect 158 113 164 114
rect 182 118 188 119
rect 182 114 183 118
rect 187 114 188 118
rect 182 113 188 114
rect 206 118 212 119
rect 206 114 207 118
rect 211 114 212 118
rect 206 113 212 114
rect 230 118 236 119
rect 230 114 231 118
rect 235 114 236 118
rect 254 118 260 119
rect 230 113 236 114
rect 242 115 248 116
rect 110 109 111 113
rect 115 109 116 113
rect 242 111 243 115
rect 247 111 248 115
rect 254 114 255 118
rect 259 114 260 118
rect 254 113 260 114
rect 278 118 284 119
rect 278 114 279 118
rect 283 114 284 118
rect 278 113 284 114
rect 302 118 308 119
rect 302 114 303 118
rect 307 114 308 118
rect 302 113 308 114
rect 326 118 332 119
rect 326 114 327 118
rect 331 114 332 118
rect 326 113 332 114
rect 350 118 356 119
rect 350 114 351 118
rect 355 114 356 118
rect 350 113 356 114
rect 374 118 380 119
rect 374 114 375 118
rect 379 114 380 118
rect 374 113 380 114
rect 398 118 404 119
rect 398 114 399 118
rect 403 114 404 118
rect 410 115 411 119
rect 415 115 416 119
rect 410 114 416 115
rect 430 118 436 119
rect 430 114 431 118
rect 435 114 436 118
rect 398 113 404 114
rect 430 113 436 114
rect 462 118 468 119
rect 462 114 463 118
rect 467 114 468 118
rect 486 118 492 119
rect 462 113 468 114
rect 474 115 480 116
rect 242 110 248 111
rect 474 111 475 115
rect 479 111 480 115
rect 486 114 487 118
rect 491 114 492 118
rect 486 113 492 114
rect 510 118 516 119
rect 510 114 511 118
rect 515 114 516 118
rect 510 113 516 114
rect 534 118 540 119
rect 534 114 535 118
rect 539 114 540 118
rect 534 113 540 114
rect 558 118 564 119
rect 558 114 559 118
rect 563 114 564 118
rect 558 113 564 114
rect 582 118 588 119
rect 582 114 583 118
rect 587 114 588 118
rect 582 113 588 114
rect 606 118 612 119
rect 606 114 607 118
rect 611 114 612 118
rect 606 113 612 114
rect 630 118 636 119
rect 630 114 631 118
rect 635 114 636 118
rect 630 113 636 114
rect 654 118 660 119
rect 654 114 655 118
rect 659 114 660 118
rect 654 113 660 114
rect 678 118 684 119
rect 678 114 679 118
rect 683 114 684 118
rect 678 113 684 114
rect 702 118 708 119
rect 702 114 703 118
rect 707 114 708 118
rect 702 113 708 114
rect 726 118 732 119
rect 726 114 727 118
rect 731 114 732 118
rect 726 113 732 114
rect 750 118 756 119
rect 750 114 751 118
rect 755 114 756 118
rect 750 113 756 114
rect 774 118 780 119
rect 774 114 775 118
rect 779 114 780 118
rect 774 113 780 114
rect 798 118 804 119
rect 798 114 799 118
rect 803 114 804 118
rect 798 113 804 114
rect 822 118 828 119
rect 822 114 823 118
rect 827 114 828 118
rect 822 113 828 114
rect 854 118 860 119
rect 854 114 855 118
rect 859 114 860 118
rect 854 113 860 114
rect 886 118 892 119
rect 886 114 887 118
rect 891 114 892 118
rect 886 113 892 114
rect 918 118 924 119
rect 918 114 919 118
rect 923 114 924 118
rect 918 113 924 114
rect 950 118 956 119
rect 950 114 951 118
rect 955 114 956 118
rect 950 113 956 114
rect 982 118 988 119
rect 982 114 983 118
rect 987 114 988 118
rect 982 113 988 114
rect 1014 118 1020 119
rect 1014 114 1015 118
rect 1019 114 1020 118
rect 1014 113 1020 114
rect 474 110 480 111
rect 110 108 116 109
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 110 90 116 91
rect 134 92 140 93
rect 112 87 114 90
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 158 92 164 93
rect 158 88 159 92
rect 163 88 164 92
rect 158 87 164 88
rect 182 92 188 93
rect 182 88 183 92
rect 187 88 188 92
rect 182 87 188 88
rect 206 92 212 93
rect 206 88 207 92
rect 211 88 212 92
rect 206 87 212 88
rect 230 92 236 93
rect 230 88 231 92
rect 235 88 236 92
rect 230 87 236 88
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 159 86 163 87
rect 159 81 163 82
rect 183 86 187 87
rect 183 81 187 82
rect 207 86 211 87
rect 207 81 211 82
rect 231 86 235 87
rect 244 84 246 110
rect 462 107 468 108
rect 476 107 478 110
rect 462 103 463 107
rect 467 105 478 107
rect 1024 107 1026 130
rect 1032 127 1034 141
rect 1054 139 1060 140
rect 1054 135 1055 139
rect 1059 135 1060 139
rect 1054 134 1060 135
rect 1031 126 1035 127
rect 1031 121 1035 122
rect 1047 126 1051 127
rect 1047 121 1051 122
rect 1048 119 1050 121
rect 1046 118 1052 119
rect 1046 114 1047 118
rect 1051 114 1052 118
rect 1046 113 1052 114
rect 1056 108 1058 134
rect 1080 127 1082 141
rect 1128 127 1130 141
rect 1176 127 1178 141
rect 1224 127 1226 141
rect 1264 127 1266 141
rect 1272 140 1274 178
rect 1279 173 1283 174
rect 1295 178 1299 179
rect 1295 173 1299 174
rect 1327 178 1331 179
rect 1327 173 1331 174
rect 1359 178 1363 179
rect 1359 173 1363 174
rect 1294 172 1300 173
rect 1294 168 1295 172
rect 1299 168 1300 172
rect 1294 167 1300 168
rect 1326 172 1332 173
rect 1326 168 1327 172
rect 1331 168 1332 172
rect 1326 167 1332 168
rect 1358 172 1364 173
rect 1372 172 1374 194
rect 1446 187 1452 188
rect 1382 184 1388 185
rect 1382 180 1383 184
rect 1387 180 1388 184
rect 1382 179 1388 180
rect 1414 184 1420 185
rect 1414 180 1415 184
rect 1419 180 1420 184
rect 1414 179 1420 180
rect 1426 183 1432 184
rect 1426 179 1427 183
rect 1431 179 1432 183
rect 1446 183 1447 187
rect 1451 183 1452 187
rect 1446 182 1452 183
rect 1448 179 1450 182
rect 1383 178 1387 179
rect 1383 173 1387 174
rect 1391 178 1395 179
rect 1391 173 1395 174
rect 1415 178 1419 179
rect 1426 178 1432 179
rect 1447 178 1451 179
rect 1415 173 1419 174
rect 1390 172 1396 173
rect 1358 168 1359 172
rect 1363 168 1364 172
rect 1358 167 1364 168
rect 1370 171 1376 172
rect 1370 167 1371 171
rect 1375 167 1376 171
rect 1390 168 1391 172
rect 1395 168 1396 172
rect 1390 167 1396 168
rect 1414 172 1420 173
rect 1414 168 1415 172
rect 1419 168 1420 172
rect 1414 167 1420 168
rect 1370 166 1376 167
rect 1398 159 1404 160
rect 1398 155 1399 159
rect 1403 155 1404 159
rect 1398 154 1404 155
rect 1294 146 1300 147
rect 1294 142 1295 146
rect 1299 142 1300 146
rect 1294 141 1300 142
rect 1326 146 1332 147
rect 1326 142 1327 146
rect 1331 142 1332 146
rect 1326 141 1332 142
rect 1358 146 1364 147
rect 1358 142 1359 146
rect 1363 142 1364 146
rect 1358 141 1364 142
rect 1390 146 1396 147
rect 1390 142 1391 146
rect 1395 142 1396 146
rect 1390 141 1396 142
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1296 127 1298 141
rect 1328 127 1330 141
rect 1360 127 1362 141
rect 1374 139 1380 140
rect 1374 135 1375 139
rect 1379 135 1380 139
rect 1374 134 1380 135
rect 1071 126 1075 127
rect 1071 121 1075 122
rect 1079 126 1083 127
rect 1079 121 1083 122
rect 1095 126 1099 127
rect 1095 121 1099 122
rect 1119 126 1123 127
rect 1119 121 1123 122
rect 1127 126 1131 127
rect 1127 121 1131 122
rect 1143 126 1147 127
rect 1143 121 1147 122
rect 1175 126 1179 127
rect 1175 121 1179 122
rect 1207 126 1211 127
rect 1207 121 1211 122
rect 1223 126 1227 127
rect 1223 121 1227 122
rect 1239 126 1243 127
rect 1239 121 1243 122
rect 1263 126 1267 127
rect 1263 121 1267 122
rect 1271 126 1275 127
rect 1271 121 1275 122
rect 1295 126 1299 127
rect 1295 121 1299 122
rect 1303 126 1307 127
rect 1303 121 1307 122
rect 1327 126 1331 127
rect 1327 121 1331 122
rect 1335 126 1339 127
rect 1335 121 1339 122
rect 1359 126 1363 127
rect 1359 121 1363 122
rect 1367 126 1371 127
rect 1367 121 1371 122
rect 1072 119 1074 121
rect 1096 119 1098 121
rect 1120 119 1122 121
rect 1144 119 1146 121
rect 1176 119 1178 121
rect 1208 119 1210 121
rect 1240 119 1242 121
rect 1272 119 1274 121
rect 1304 119 1306 121
rect 1336 119 1338 121
rect 1368 119 1370 121
rect 1070 118 1076 119
rect 1070 114 1071 118
rect 1075 114 1076 118
rect 1070 113 1076 114
rect 1094 118 1100 119
rect 1094 114 1095 118
rect 1099 114 1100 118
rect 1094 113 1100 114
rect 1118 118 1124 119
rect 1118 114 1119 118
rect 1123 114 1124 118
rect 1118 113 1124 114
rect 1142 118 1148 119
rect 1142 114 1143 118
rect 1147 114 1148 118
rect 1142 113 1148 114
rect 1174 118 1180 119
rect 1174 114 1175 118
rect 1179 114 1180 118
rect 1174 113 1180 114
rect 1206 118 1212 119
rect 1206 114 1207 118
rect 1211 114 1212 118
rect 1206 113 1212 114
rect 1238 118 1244 119
rect 1238 114 1239 118
rect 1243 114 1244 118
rect 1238 113 1244 114
rect 1270 118 1276 119
rect 1270 114 1271 118
rect 1275 114 1276 118
rect 1270 113 1276 114
rect 1302 118 1308 119
rect 1302 114 1303 118
rect 1307 114 1308 118
rect 1302 113 1308 114
rect 1334 118 1340 119
rect 1334 114 1335 118
rect 1339 114 1340 118
rect 1334 113 1340 114
rect 1366 118 1372 119
rect 1366 114 1367 118
rect 1371 114 1372 118
rect 1366 113 1372 114
rect 1376 108 1378 134
rect 1392 127 1394 141
rect 1400 128 1402 154
rect 1428 148 1430 178
rect 1447 173 1451 174
rect 1448 170 1450 173
rect 1446 169 1452 170
rect 1446 165 1447 169
rect 1451 165 1452 169
rect 1446 164 1452 165
rect 1446 151 1452 152
rect 1426 147 1432 148
rect 1414 146 1420 147
rect 1414 142 1415 146
rect 1419 142 1420 146
rect 1426 143 1427 147
rect 1431 143 1432 147
rect 1446 147 1447 151
rect 1451 147 1452 151
rect 1446 146 1452 147
rect 1426 142 1432 143
rect 1414 141 1420 142
rect 1398 127 1404 128
rect 1416 127 1418 141
rect 1448 127 1450 146
rect 1391 126 1395 127
rect 1398 123 1399 127
rect 1403 123 1404 127
rect 1398 122 1404 123
rect 1415 126 1419 127
rect 1391 121 1395 122
rect 1415 121 1419 122
rect 1447 126 1451 127
rect 1447 121 1451 122
rect 1392 119 1394 121
rect 1416 119 1418 121
rect 1390 118 1396 119
rect 1390 114 1391 118
rect 1395 114 1396 118
rect 1390 113 1396 114
rect 1414 118 1420 119
rect 1414 114 1415 118
rect 1419 114 1420 118
rect 1448 114 1450 121
rect 1414 113 1420 114
rect 1446 113 1452 114
rect 1446 109 1447 113
rect 1451 109 1452 113
rect 1446 108 1452 109
rect 1054 107 1060 108
rect 1024 105 1030 107
rect 467 103 468 105
rect 462 102 468 103
rect 1028 96 1030 105
rect 1054 103 1055 107
rect 1059 103 1060 107
rect 1054 102 1060 103
rect 1374 107 1380 108
rect 1374 103 1375 107
rect 1379 103 1380 107
rect 1374 102 1380 103
rect 1026 95 1032 96
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 278 92 284 93
rect 278 88 279 92
rect 283 88 284 92
rect 278 87 284 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 326 92 332 93
rect 326 88 327 92
rect 331 88 332 92
rect 326 87 332 88
rect 350 92 356 93
rect 350 88 351 92
rect 355 88 356 92
rect 350 87 356 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 398 92 404 93
rect 398 88 399 92
rect 403 88 404 92
rect 398 87 404 88
rect 430 92 436 93
rect 430 88 431 92
rect 435 88 436 92
rect 430 87 436 88
rect 462 92 468 93
rect 462 88 463 92
rect 467 88 468 92
rect 462 87 468 88
rect 486 92 492 93
rect 486 88 487 92
rect 491 88 492 92
rect 486 87 492 88
rect 510 92 516 93
rect 510 88 511 92
rect 515 88 516 92
rect 510 87 516 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 558 92 564 93
rect 558 88 559 92
rect 563 88 564 92
rect 558 87 564 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 606 92 612 93
rect 606 88 607 92
rect 611 88 612 92
rect 606 87 612 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 654 92 660 93
rect 654 88 655 92
rect 659 88 660 92
rect 654 87 660 88
rect 678 92 684 93
rect 678 88 679 92
rect 683 88 684 92
rect 678 87 684 88
rect 702 92 708 93
rect 702 88 703 92
rect 707 88 708 92
rect 702 87 708 88
rect 726 92 732 93
rect 726 88 727 92
rect 731 88 732 92
rect 726 87 732 88
rect 750 92 756 93
rect 750 88 751 92
rect 755 88 756 92
rect 750 87 756 88
rect 774 92 780 93
rect 774 88 775 92
rect 779 88 780 92
rect 774 87 780 88
rect 798 92 804 93
rect 798 88 799 92
rect 803 88 804 92
rect 798 87 804 88
rect 822 92 828 93
rect 822 88 823 92
rect 827 88 828 92
rect 822 87 828 88
rect 854 92 860 93
rect 854 88 855 92
rect 859 88 860 92
rect 854 87 860 88
rect 886 92 892 93
rect 886 88 887 92
rect 891 88 892 92
rect 886 87 892 88
rect 918 92 924 93
rect 918 88 919 92
rect 923 88 924 92
rect 918 87 924 88
rect 950 92 956 93
rect 950 88 951 92
rect 955 88 956 92
rect 950 87 956 88
rect 982 92 988 93
rect 982 88 983 92
rect 987 88 988 92
rect 982 87 988 88
rect 1014 92 1020 93
rect 1014 88 1015 92
rect 1019 88 1020 92
rect 1026 91 1027 95
rect 1031 91 1032 95
rect 1446 95 1452 96
rect 1026 90 1032 91
rect 1046 92 1052 93
rect 1014 87 1020 88
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1046 87 1052 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1094 92 1100 93
rect 1094 88 1095 92
rect 1099 88 1100 92
rect 1094 87 1100 88
rect 1118 92 1124 93
rect 1118 88 1119 92
rect 1123 88 1124 92
rect 1118 87 1124 88
rect 1142 92 1148 93
rect 1142 88 1143 92
rect 1147 88 1148 92
rect 1142 87 1148 88
rect 1174 92 1180 93
rect 1174 88 1175 92
rect 1179 88 1180 92
rect 1174 87 1180 88
rect 1206 92 1212 93
rect 1206 88 1207 92
rect 1211 88 1212 92
rect 1206 87 1212 88
rect 1238 92 1244 93
rect 1238 88 1239 92
rect 1243 88 1244 92
rect 1238 87 1244 88
rect 1270 92 1276 93
rect 1270 88 1271 92
rect 1275 88 1276 92
rect 1270 87 1276 88
rect 1302 92 1308 93
rect 1302 88 1303 92
rect 1307 88 1308 92
rect 1302 87 1308 88
rect 1334 92 1340 93
rect 1334 88 1335 92
rect 1339 88 1340 92
rect 1334 87 1340 88
rect 1366 92 1372 93
rect 1366 88 1367 92
rect 1371 88 1372 92
rect 1366 87 1372 88
rect 1390 92 1396 93
rect 1390 88 1391 92
rect 1395 88 1396 92
rect 1390 87 1396 88
rect 1414 92 1420 93
rect 1414 88 1415 92
rect 1419 88 1420 92
rect 1446 91 1447 95
rect 1451 91 1452 95
rect 1446 90 1452 91
rect 1414 87 1420 88
rect 1448 87 1450 90
rect 255 86 259 87
rect 231 81 235 82
rect 242 83 248 84
rect 242 79 243 83
rect 247 79 248 83
rect 255 81 259 82
rect 279 86 283 87
rect 279 81 283 82
rect 303 86 307 87
rect 303 81 307 82
rect 327 86 331 87
rect 327 81 331 82
rect 351 86 355 87
rect 351 81 355 82
rect 375 86 379 87
rect 375 81 379 82
rect 399 86 403 87
rect 399 81 403 82
rect 431 86 435 87
rect 431 81 435 82
rect 463 86 467 87
rect 463 81 467 82
rect 487 86 491 87
rect 487 81 491 82
rect 511 86 515 87
rect 511 81 515 82
rect 535 86 539 87
rect 535 81 539 82
rect 559 86 563 87
rect 559 81 563 82
rect 583 86 587 87
rect 583 81 587 82
rect 607 86 611 87
rect 607 81 611 82
rect 631 86 635 87
rect 631 81 635 82
rect 655 86 659 87
rect 655 81 659 82
rect 679 86 683 87
rect 679 81 683 82
rect 703 86 707 87
rect 703 81 707 82
rect 727 86 731 87
rect 727 81 731 82
rect 751 86 755 87
rect 751 81 755 82
rect 775 86 779 87
rect 775 81 779 82
rect 799 86 803 87
rect 799 81 803 82
rect 823 86 827 87
rect 823 81 827 82
rect 855 86 859 87
rect 855 81 859 82
rect 887 86 891 87
rect 887 81 891 82
rect 919 86 923 87
rect 919 81 923 82
rect 951 86 955 87
rect 951 81 955 82
rect 983 86 987 87
rect 983 81 987 82
rect 1015 86 1019 87
rect 1015 81 1019 82
rect 1047 86 1051 87
rect 1047 81 1051 82
rect 1071 86 1075 87
rect 1071 81 1075 82
rect 1095 86 1099 87
rect 1095 81 1099 82
rect 1119 86 1123 87
rect 1119 81 1123 82
rect 1143 86 1147 87
rect 1143 81 1147 82
rect 1175 86 1179 87
rect 1175 81 1179 82
rect 1207 86 1211 87
rect 1207 81 1211 82
rect 1239 86 1243 87
rect 1239 81 1243 82
rect 1271 86 1275 87
rect 1271 81 1275 82
rect 1303 86 1307 87
rect 1303 81 1307 82
rect 1335 86 1339 87
rect 1335 81 1339 82
rect 1367 86 1371 87
rect 1367 81 1371 82
rect 1391 86 1395 87
rect 1391 81 1395 82
rect 1415 86 1419 87
rect 1415 81 1419 82
rect 1447 86 1451 87
rect 1447 81 1451 82
rect 242 78 248 79
<< m4c >>
rect 111 1506 115 1510
rect 295 1506 299 1510
rect 319 1506 323 1510
rect 343 1506 347 1510
rect 367 1506 371 1510
rect 407 1506 411 1510
rect 455 1506 459 1510
rect 511 1506 515 1510
rect 575 1506 579 1510
rect 647 1506 651 1510
rect 727 1506 731 1510
rect 807 1506 811 1510
rect 887 1506 891 1510
rect 959 1506 963 1510
rect 1031 1506 1035 1510
rect 1103 1506 1107 1510
rect 1175 1506 1179 1510
rect 1247 1506 1251 1510
rect 1447 1506 1451 1510
rect 111 1466 115 1470
rect 151 1466 155 1470
rect 175 1466 179 1470
rect 199 1466 203 1470
rect 231 1466 235 1470
rect 271 1466 275 1470
rect 295 1466 299 1470
rect 319 1466 323 1470
rect 343 1466 347 1470
rect 367 1466 371 1470
rect 407 1466 411 1470
rect 455 1466 459 1470
rect 503 1466 507 1470
rect 511 1466 515 1470
rect 551 1466 555 1470
rect 575 1466 579 1470
rect 607 1466 611 1470
rect 647 1466 651 1470
rect 663 1466 667 1470
rect 711 1466 715 1470
rect 727 1466 731 1470
rect 759 1466 763 1470
rect 807 1466 811 1470
rect 815 1466 819 1470
rect 871 1466 875 1470
rect 887 1466 891 1470
rect 927 1466 931 1470
rect 959 1466 963 1470
rect 975 1466 979 1470
rect 1023 1466 1027 1470
rect 1031 1466 1035 1470
rect 1071 1466 1075 1470
rect 1103 1466 1107 1470
rect 1119 1466 1123 1470
rect 1167 1466 1171 1470
rect 1175 1466 1179 1470
rect 1215 1466 1219 1470
rect 1247 1466 1251 1470
rect 1263 1466 1267 1470
rect 1311 1466 1315 1470
rect 1447 1466 1451 1470
rect 111 1426 115 1430
rect 135 1426 139 1430
rect 151 1426 155 1430
rect 159 1426 163 1430
rect 175 1426 179 1430
rect 183 1426 187 1430
rect 199 1426 203 1430
rect 223 1426 227 1430
rect 111 1386 115 1390
rect 135 1386 139 1390
rect 159 1386 163 1390
rect 183 1386 187 1390
rect 231 1426 235 1430
rect 271 1426 275 1430
rect 287 1426 291 1430
rect 319 1426 323 1430
rect 223 1386 227 1390
rect 231 1386 235 1390
rect 279 1386 283 1390
rect 287 1386 291 1390
rect 351 1426 355 1430
rect 367 1426 371 1430
rect 407 1426 411 1430
rect 415 1426 419 1430
rect 455 1426 459 1430
rect 479 1426 483 1430
rect 503 1426 507 1430
rect 535 1426 539 1430
rect 551 1426 555 1430
rect 583 1426 587 1430
rect 607 1426 611 1430
rect 631 1426 635 1430
rect 663 1426 667 1430
rect 687 1426 691 1430
rect 711 1426 715 1430
rect 743 1426 747 1430
rect 759 1426 763 1430
rect 799 1426 803 1430
rect 815 1426 819 1430
rect 855 1426 859 1430
rect 871 1426 875 1430
rect 911 1426 915 1430
rect 927 1426 931 1430
rect 967 1426 971 1430
rect 975 1426 979 1430
rect 1023 1426 1027 1430
rect 1071 1426 1075 1430
rect 1119 1426 1123 1430
rect 335 1386 339 1390
rect 351 1386 355 1390
rect 391 1386 395 1390
rect 415 1386 419 1390
rect 439 1386 443 1390
rect 479 1386 483 1390
rect 487 1386 491 1390
rect 527 1386 531 1390
rect 535 1386 539 1390
rect 567 1386 571 1390
rect 583 1386 587 1390
rect 615 1386 619 1390
rect 631 1386 635 1390
rect 663 1386 667 1390
rect 687 1386 691 1390
rect 711 1386 715 1390
rect 743 1386 747 1390
rect 767 1386 771 1390
rect 799 1386 803 1390
rect 823 1386 827 1390
rect 855 1386 859 1390
rect 879 1386 883 1390
rect 911 1386 915 1390
rect 935 1386 939 1390
rect 967 1386 971 1390
rect 991 1386 995 1390
rect 1023 1386 1027 1390
rect 1047 1386 1051 1390
rect 1071 1386 1075 1390
rect 1167 1426 1171 1430
rect 1215 1426 1219 1430
rect 1263 1426 1267 1430
rect 1303 1426 1307 1430
rect 1311 1426 1315 1430
rect 1343 1426 1347 1430
rect 1391 1426 1395 1430
rect 1095 1386 1099 1390
rect 1119 1386 1123 1390
rect 1143 1386 1147 1390
rect 1167 1386 1171 1390
rect 1191 1386 1195 1390
rect 111 1346 115 1350
rect 135 1346 139 1350
rect 159 1346 163 1350
rect 167 1346 171 1350
rect 183 1346 187 1350
rect 191 1346 195 1350
rect 231 1346 235 1350
rect 279 1346 283 1350
rect 335 1346 339 1350
rect 391 1346 395 1350
rect 439 1346 443 1350
rect 455 1346 459 1350
rect 487 1346 491 1350
rect 519 1346 523 1350
rect 243 1320 247 1324
rect 327 1323 331 1324
rect 327 1320 331 1323
rect 111 1306 115 1310
rect 167 1306 171 1310
rect 191 1306 195 1310
rect 231 1306 235 1310
rect 255 1306 259 1310
rect 279 1306 283 1310
rect 303 1306 307 1310
rect 327 1306 331 1310
rect 335 1306 339 1310
rect 351 1306 355 1310
rect 375 1306 379 1310
rect 391 1306 395 1310
rect 399 1306 403 1310
rect 527 1346 531 1350
rect 567 1346 571 1350
rect 575 1346 579 1350
rect 615 1346 619 1350
rect 631 1346 635 1350
rect 663 1346 667 1350
rect 679 1346 683 1350
rect 711 1346 715 1350
rect 727 1346 731 1350
rect 767 1346 771 1350
rect 799 1346 803 1350
rect 823 1346 827 1350
rect 831 1346 835 1350
rect 863 1346 867 1350
rect 879 1346 883 1350
rect 895 1346 899 1350
rect 927 1346 931 1350
rect 935 1346 939 1350
rect 967 1346 971 1350
rect 991 1346 995 1350
rect 1007 1346 1011 1350
rect 1047 1346 1051 1350
rect 1055 1346 1059 1350
rect 1095 1346 1099 1350
rect 1103 1346 1107 1350
rect 423 1306 427 1310
rect 447 1306 451 1310
rect 455 1306 459 1310
rect 471 1306 475 1310
rect 503 1306 507 1310
rect 519 1306 523 1310
rect 543 1306 547 1310
rect 575 1306 579 1310
rect 591 1306 595 1310
rect 631 1306 635 1310
rect 647 1306 651 1310
rect 111 1266 115 1270
rect 231 1266 235 1270
rect 255 1266 259 1270
rect 279 1266 283 1270
rect 303 1266 307 1270
rect 311 1266 315 1270
rect 679 1306 683 1310
rect 695 1306 699 1310
rect 727 1306 731 1310
rect 743 1306 747 1310
rect 767 1306 771 1310
rect 791 1306 795 1310
rect 799 1306 803 1310
rect 831 1306 835 1310
rect 839 1306 843 1310
rect 863 1306 867 1310
rect 879 1306 883 1310
rect 895 1306 899 1310
rect 911 1306 915 1310
rect 927 1306 931 1310
rect 951 1306 955 1310
rect 967 1306 971 1310
rect 1143 1346 1147 1350
rect 1159 1346 1163 1350
rect 1215 1386 1219 1390
rect 1239 1386 1243 1390
rect 1263 1386 1267 1390
rect 1287 1386 1291 1390
rect 1303 1386 1307 1390
rect 1415 1426 1419 1430
rect 1447 1426 1451 1430
rect 1335 1386 1339 1390
rect 1343 1386 1347 1390
rect 1383 1386 1387 1390
rect 1391 1386 1395 1390
rect 1415 1386 1419 1390
rect 1447 1386 1451 1390
rect 1191 1346 1195 1350
rect 1215 1346 1219 1350
rect 1239 1346 1243 1350
rect 1271 1346 1275 1350
rect 1287 1346 1291 1350
rect 1327 1346 1331 1350
rect 1335 1346 1339 1350
rect 991 1306 995 1310
rect 1007 1306 1011 1310
rect 1031 1306 1035 1310
rect 1055 1306 1059 1310
rect 1071 1306 1075 1310
rect 1103 1306 1107 1310
rect 1111 1306 1115 1310
rect 1151 1306 1155 1310
rect 1159 1306 1163 1310
rect 1199 1306 1203 1310
rect 1215 1306 1219 1310
rect 1247 1306 1251 1310
rect 327 1266 331 1270
rect 335 1266 339 1270
rect 351 1266 355 1270
rect 359 1266 363 1270
rect 375 1266 379 1270
rect 383 1266 387 1270
rect 399 1266 403 1270
rect 415 1266 419 1270
rect 423 1266 427 1270
rect 447 1266 451 1270
rect 471 1266 475 1270
rect 479 1266 483 1270
rect 503 1266 507 1270
rect 519 1266 523 1270
rect 543 1266 547 1270
rect 559 1266 563 1270
rect 591 1266 595 1270
rect 615 1266 619 1270
rect 647 1266 651 1270
rect 679 1266 683 1270
rect 695 1266 699 1270
rect 743 1266 747 1270
rect 751 1266 755 1270
rect 791 1266 795 1270
rect 831 1266 835 1270
rect 839 1266 843 1270
rect 879 1266 883 1270
rect 911 1266 915 1270
rect 951 1266 955 1270
rect 991 1266 995 1270
rect 1031 1266 1035 1270
rect 111 1226 115 1230
rect 311 1226 315 1230
rect 327 1226 331 1230
rect 335 1226 339 1230
rect 359 1226 363 1230
rect 367 1226 371 1230
rect 383 1226 387 1230
rect 407 1226 411 1230
rect 415 1226 419 1230
rect 447 1226 451 1230
rect 479 1226 483 1230
rect 487 1226 491 1230
rect 519 1226 523 1230
rect 527 1226 531 1230
rect 559 1226 563 1230
rect 567 1226 571 1230
rect 607 1226 611 1230
rect 615 1226 619 1230
rect 655 1226 659 1230
rect 679 1226 683 1230
rect 1063 1266 1067 1270
rect 1071 1266 1075 1270
rect 1111 1266 1115 1270
rect 1127 1266 1131 1270
rect 1271 1306 1275 1310
rect 1303 1306 1307 1310
rect 1383 1346 1387 1350
rect 1415 1346 1419 1350
rect 1447 1346 1451 1350
rect 1327 1306 1331 1310
rect 1367 1306 1371 1310
rect 1383 1306 1387 1310
rect 1415 1306 1419 1310
rect 1151 1266 1155 1270
rect 1191 1266 1195 1270
rect 1199 1266 1203 1270
rect 1247 1266 1251 1270
rect 1303 1266 1307 1270
rect 703 1226 707 1230
rect 751 1226 755 1230
rect 111 1186 115 1190
rect 135 1186 139 1190
rect 159 1186 163 1190
rect 183 1186 187 1190
rect 207 1186 211 1190
rect 231 1186 235 1190
rect 255 1186 259 1190
rect 279 1186 283 1190
rect 303 1186 307 1190
rect 327 1186 331 1190
rect 335 1186 339 1190
rect 799 1226 803 1230
rect 831 1226 835 1230
rect 847 1226 851 1230
rect 895 1226 899 1230
rect 911 1226 915 1230
rect 943 1226 947 1230
rect 991 1226 995 1230
rect 1039 1226 1043 1230
rect 1063 1226 1067 1230
rect 1103 1226 1107 1230
rect 1127 1226 1131 1230
rect 1175 1226 1179 1230
rect 1191 1226 1195 1230
rect 1247 1226 1251 1230
rect 1255 1226 1259 1230
rect 1311 1266 1315 1270
rect 1367 1266 1371 1270
rect 1375 1266 1379 1270
rect 1447 1306 1451 1310
rect 1415 1266 1419 1270
rect 1447 1266 1451 1270
rect 1311 1226 1315 1230
rect 1343 1226 1347 1230
rect 1375 1226 1379 1230
rect 1415 1226 1419 1230
rect 367 1186 371 1190
rect 383 1186 387 1190
rect 407 1186 411 1190
rect 423 1186 427 1190
rect 111 1146 115 1150
rect 135 1146 139 1150
rect 159 1146 163 1150
rect 183 1146 187 1150
rect 207 1146 211 1150
rect 215 1146 219 1150
rect 231 1146 235 1150
rect 255 1146 259 1150
rect 279 1146 283 1150
rect 295 1146 299 1150
rect 303 1146 307 1150
rect 335 1146 339 1150
rect 375 1146 379 1150
rect 383 1146 387 1150
rect 447 1186 451 1190
rect 463 1186 467 1190
rect 487 1186 491 1190
rect 503 1186 507 1190
rect 527 1186 531 1190
rect 543 1186 547 1190
rect 567 1186 571 1190
rect 583 1186 587 1190
rect 607 1186 611 1190
rect 623 1186 627 1190
rect 655 1186 659 1190
rect 671 1186 675 1190
rect 703 1186 707 1190
rect 415 1146 419 1150
rect 423 1146 427 1150
rect 463 1146 467 1150
rect 503 1146 507 1150
rect 519 1146 523 1150
rect 543 1146 547 1150
rect 583 1146 587 1150
rect 623 1146 627 1150
rect 647 1146 651 1150
rect 671 1146 675 1150
rect 719 1186 723 1190
rect 751 1186 755 1190
rect 767 1186 771 1190
rect 799 1186 803 1190
rect 815 1186 819 1190
rect 847 1186 851 1190
rect 863 1186 867 1190
rect 895 1186 899 1190
rect 911 1186 915 1190
rect 1447 1226 1451 1230
rect 943 1186 947 1190
rect 959 1186 963 1190
rect 991 1186 995 1190
rect 1007 1186 1011 1190
rect 1039 1186 1043 1190
rect 1055 1186 1059 1190
rect 1103 1186 1107 1190
rect 1151 1186 1155 1190
rect 711 1146 715 1150
rect 719 1146 723 1150
rect 767 1146 771 1150
rect 815 1146 819 1150
rect 831 1146 835 1150
rect 111 1102 115 1106
rect 135 1102 139 1106
rect 159 1102 163 1106
rect 183 1102 187 1106
rect 863 1146 867 1150
rect 887 1146 891 1150
rect 911 1146 915 1150
rect 943 1146 947 1150
rect 959 1146 963 1150
rect 999 1146 1003 1150
rect 1007 1146 1011 1150
rect 1175 1186 1179 1190
rect 1191 1186 1195 1190
rect 1231 1186 1235 1190
rect 1255 1186 1259 1190
rect 1271 1186 1275 1190
rect 1311 1186 1315 1190
rect 1343 1186 1347 1190
rect 1351 1186 1355 1190
rect 1391 1186 1395 1190
rect 1415 1186 1419 1190
rect 1447 1186 1451 1190
rect 1055 1146 1059 1150
rect 1103 1146 1107 1150
rect 1151 1146 1155 1150
rect 207 1102 211 1106
rect 215 1102 219 1106
rect 247 1102 251 1106
rect 255 1102 259 1106
rect 287 1102 291 1106
rect 295 1102 299 1106
rect 327 1102 331 1106
rect 335 1102 339 1106
rect 367 1102 371 1106
rect 375 1102 379 1106
rect 1191 1146 1195 1150
rect 1231 1146 1235 1150
rect 1271 1146 1275 1150
rect 1311 1146 1315 1150
rect 1351 1146 1355 1150
rect 1391 1146 1395 1150
rect 1415 1146 1419 1150
rect 1447 1146 1451 1150
rect 407 1102 411 1106
rect 415 1102 419 1106
rect 455 1102 459 1106
rect 463 1102 467 1106
rect 503 1102 507 1106
rect 519 1102 523 1106
rect 559 1102 563 1106
rect 583 1102 587 1106
rect 607 1102 611 1106
rect 647 1102 651 1106
rect 655 1102 659 1106
rect 703 1102 707 1106
rect 711 1102 715 1106
rect 743 1102 747 1106
rect 767 1102 771 1106
rect 791 1102 795 1106
rect 831 1102 835 1106
rect 839 1102 843 1106
rect 887 1102 891 1106
rect 943 1102 947 1106
rect 999 1102 1003 1106
rect 1055 1102 1059 1106
rect 1103 1102 1107 1106
rect 1111 1102 1115 1106
rect 1151 1102 1155 1106
rect 147 1075 151 1076
rect 147 1072 148 1075
rect 148 1072 151 1075
rect 219 1072 223 1076
rect 111 1062 115 1066
rect 135 1062 139 1066
rect 159 1062 163 1066
rect 183 1062 187 1066
rect 207 1062 211 1066
rect 231 1062 235 1066
rect 247 1062 251 1066
rect 271 1062 275 1066
rect 287 1062 291 1066
rect 147 1040 151 1044
rect 311 1062 315 1066
rect 327 1062 331 1066
rect 351 1062 355 1066
rect 367 1062 371 1066
rect 391 1062 395 1066
rect 407 1062 411 1066
rect 431 1062 435 1066
rect 455 1062 459 1066
rect 471 1062 475 1066
rect 503 1062 507 1066
rect 511 1062 515 1066
rect 551 1062 555 1066
rect 559 1062 563 1066
rect 591 1062 595 1066
rect 607 1062 611 1066
rect 631 1062 635 1066
rect 655 1062 659 1066
rect 671 1062 675 1066
rect 299 1040 303 1044
rect 703 1062 707 1066
rect 711 1062 715 1066
rect 743 1062 747 1066
rect 783 1062 787 1066
rect 791 1062 795 1066
rect 823 1062 827 1066
rect 839 1062 843 1066
rect 871 1062 875 1066
rect 887 1062 891 1066
rect 919 1062 923 1066
rect 943 1062 947 1066
rect 975 1062 979 1066
rect 999 1062 1003 1066
rect 1167 1102 1171 1106
rect 1191 1102 1195 1106
rect 1215 1102 1219 1106
rect 1231 1102 1235 1106
rect 1271 1102 1275 1106
rect 1311 1102 1315 1106
rect 1327 1102 1331 1106
rect 1351 1102 1355 1106
rect 1031 1062 1035 1066
rect 1055 1062 1059 1066
rect 1079 1062 1083 1066
rect 1111 1062 1115 1066
rect 1127 1062 1131 1066
rect 695 1032 699 1036
rect 111 1022 115 1026
rect 135 1022 139 1026
rect 159 1022 163 1026
rect 183 1022 187 1026
rect 207 1022 211 1026
rect 231 1022 235 1026
rect 263 1022 267 1026
rect 271 1022 275 1026
rect 303 1022 307 1026
rect 311 1022 315 1026
rect 343 1022 347 1026
rect 351 1022 355 1026
rect 383 1022 387 1026
rect 391 1022 395 1026
rect 431 1022 435 1026
rect 471 1022 475 1026
rect 479 1022 483 1026
rect 511 1022 515 1026
rect 527 1022 531 1026
rect 551 1022 555 1026
rect 219 992 223 996
rect 111 982 115 986
rect 159 982 163 986
rect 183 982 187 986
rect 207 982 211 986
rect 355 995 359 996
rect 355 992 359 995
rect 231 982 235 986
rect 255 982 259 986
rect 263 982 267 986
rect 287 982 291 986
rect 303 982 307 986
rect 327 982 331 986
rect 343 982 347 986
rect 375 982 379 986
rect 383 982 387 986
rect 575 1022 579 1026
rect 591 1022 595 1026
rect 623 1022 627 1026
rect 631 1022 635 1026
rect 671 1022 675 1026
rect 711 1022 715 1026
rect 719 1022 723 1026
rect 743 1022 747 1026
rect 767 1022 771 1026
rect 795 1035 799 1036
rect 795 1032 799 1035
rect 783 1022 787 1026
rect 823 1022 827 1026
rect 871 1022 875 1026
rect 879 1022 883 1026
rect 919 1022 923 1026
rect 935 1022 939 1026
rect 975 1022 979 1026
rect 991 1022 995 1026
rect 1167 1062 1171 1066
rect 1175 1062 1179 1066
rect 1215 1062 1219 1066
rect 1223 1062 1227 1066
rect 1383 1102 1387 1106
rect 1391 1102 1395 1106
rect 1415 1102 1419 1106
rect 1447 1102 1451 1106
rect 1271 1062 1275 1066
rect 1327 1062 1331 1066
rect 1383 1062 1387 1066
rect 1415 1062 1419 1066
rect 1031 1022 1035 1026
rect 1047 1022 1051 1026
rect 1079 1022 1083 1026
rect 1103 1022 1107 1026
rect 1127 1022 1131 1026
rect 1159 1022 1163 1026
rect 1175 1022 1179 1026
rect 1215 1022 1219 1026
rect 1223 1022 1227 1026
rect 1271 1022 1275 1026
rect 1327 1022 1331 1026
rect 1383 1022 1387 1026
rect 1447 1062 1451 1066
rect 1415 1022 1419 1026
rect 1447 1022 1451 1026
rect 423 982 427 986
rect 431 982 435 986
rect 471 982 475 986
rect 479 982 483 986
rect 519 982 523 986
rect 527 982 531 986
rect 567 982 571 986
rect 575 982 579 986
rect 623 982 627 986
rect 671 982 675 986
rect 679 982 683 986
rect 719 982 723 986
rect 727 982 731 986
rect 767 982 771 986
rect 775 982 779 986
rect 823 982 827 986
rect 831 982 835 986
rect 879 982 883 986
rect 887 982 891 986
rect 935 982 939 986
rect 943 982 947 986
rect 991 982 995 986
rect 999 982 1003 986
rect 1047 982 1051 986
rect 1095 982 1099 986
rect 1103 982 1107 986
rect 111 942 115 946
rect 207 942 211 946
rect 215 942 219 946
rect 231 942 235 946
rect 239 942 243 946
rect 255 942 259 946
rect 263 942 267 946
rect 287 942 291 946
rect 319 942 323 946
rect 227 931 231 932
rect 227 928 231 931
rect 327 942 331 946
rect 351 942 355 946
rect 375 942 379 946
rect 391 942 395 946
rect 423 942 427 946
rect 431 942 435 946
rect 471 942 475 946
rect 519 942 523 946
rect 303 928 307 932
rect 443 928 447 932
rect 111 902 115 906
rect 215 902 219 906
rect 231 902 235 906
rect 239 902 243 906
rect 255 902 259 906
rect 263 902 267 906
rect 279 902 283 906
rect 287 902 291 906
rect 303 902 307 906
rect 319 902 323 906
rect 327 902 331 906
rect 351 902 355 906
rect 359 902 363 906
rect 391 902 395 906
rect 423 902 427 906
rect 431 902 435 906
rect 455 902 459 906
rect 471 902 475 906
rect 495 902 499 906
rect 567 942 571 946
rect 615 942 619 946
rect 623 942 627 946
rect 671 942 675 946
rect 679 942 683 946
rect 727 942 731 946
rect 775 942 779 946
rect 783 942 787 946
rect 539 931 543 932
rect 539 928 543 931
rect 831 942 835 946
rect 847 942 851 946
rect 887 942 891 946
rect 919 942 923 946
rect 1143 982 1147 986
rect 1159 982 1163 986
rect 1191 982 1195 986
rect 1215 982 1219 986
rect 1239 982 1243 986
rect 1271 982 1275 986
rect 1287 982 1291 986
rect 1327 982 1331 986
rect 1335 982 1339 986
rect 1383 982 1387 986
rect 1415 982 1419 986
rect 1447 982 1451 986
rect 943 942 947 946
rect 991 942 995 946
rect 999 942 1003 946
rect 1047 942 1051 946
rect 1055 942 1059 946
rect 1095 942 1099 946
rect 1119 942 1123 946
rect 1143 942 1147 946
rect 1175 942 1179 946
rect 1191 942 1195 946
rect 1223 942 1227 946
rect 1239 942 1243 946
rect 1263 942 1267 946
rect 1287 942 1291 946
rect 1295 942 1299 946
rect 1327 942 1331 946
rect 1335 942 1339 946
rect 1359 942 1363 946
rect 1383 942 1387 946
rect 1391 942 1395 946
rect 1415 942 1419 946
rect 1447 942 1451 946
rect 519 902 523 906
rect 535 902 539 906
rect 567 902 571 906
rect 575 902 579 906
rect 615 902 619 906
rect 623 902 627 906
rect 663 902 667 906
rect 671 902 675 906
rect 703 902 707 906
rect 727 902 731 906
rect 751 902 755 906
rect 783 902 787 906
rect 807 902 811 906
rect 847 902 851 906
rect 863 902 867 906
rect 919 902 923 906
rect 927 902 931 906
rect 991 902 995 906
rect 1055 902 1059 906
rect 1119 902 1123 906
rect 1175 902 1179 906
rect 1223 902 1227 906
rect 1231 902 1235 906
rect 1263 902 1267 906
rect 1279 902 1283 906
rect 1295 902 1299 906
rect 1327 902 1331 906
rect 1359 902 1363 906
rect 1383 902 1387 906
rect 1391 902 1395 906
rect 111 862 115 866
rect 207 862 211 866
rect 231 862 235 866
rect 255 862 259 866
rect 279 862 283 866
rect 287 862 291 866
rect 303 862 307 866
rect 319 862 323 866
rect 327 862 331 866
rect 351 862 355 866
rect 359 862 363 866
rect 383 862 387 866
rect 391 862 395 866
rect 415 862 419 866
rect 423 862 427 866
rect 447 862 451 866
rect 455 862 459 866
rect 479 862 483 866
rect 495 862 499 866
rect 511 862 515 866
rect 535 862 539 866
rect 551 862 555 866
rect 575 862 579 866
rect 599 862 603 866
rect 623 862 627 866
rect 647 862 651 866
rect 663 862 667 866
rect 703 862 707 866
rect 751 862 755 866
rect 767 862 771 866
rect 807 862 811 866
rect 111 822 115 826
rect 135 822 139 826
rect 159 822 163 826
rect 183 822 187 826
rect 207 822 211 826
rect 215 822 219 826
rect 231 822 235 826
rect 255 822 259 826
rect 263 822 267 826
rect 287 822 291 826
rect 311 822 315 826
rect 319 822 323 826
rect 351 822 355 826
rect 367 822 371 826
rect 383 822 387 826
rect 415 822 419 826
rect 431 822 435 826
rect 447 822 451 826
rect 479 822 483 826
rect 487 822 491 826
rect 511 822 515 826
rect 111 782 115 786
rect 135 782 139 786
rect 159 782 163 786
rect 183 782 187 786
rect 215 782 219 786
rect 223 782 227 786
rect 263 782 267 786
rect 279 782 283 786
rect 311 782 315 786
rect 343 782 347 786
rect 367 782 371 786
rect 407 782 411 786
rect 543 822 547 826
rect 551 822 555 826
rect 599 822 603 826
rect 647 822 651 826
rect 655 822 659 826
rect 839 862 843 866
rect 863 862 867 866
rect 911 862 915 866
rect 927 862 931 866
rect 983 862 987 866
rect 991 862 995 866
rect 1047 862 1051 866
rect 1055 862 1059 866
rect 1103 862 1107 866
rect 1119 862 1123 866
rect 1159 862 1163 866
rect 1175 862 1179 866
rect 703 822 707 826
rect 711 822 715 826
rect 767 822 771 826
rect 815 822 819 826
rect 839 822 843 826
rect 431 782 435 786
rect 463 782 467 786
rect 487 782 491 786
rect 519 782 523 786
rect 543 782 547 786
rect 575 782 579 786
rect 599 782 603 786
rect 623 782 627 786
rect 655 782 659 786
rect 671 782 675 786
rect 711 782 715 786
rect 719 782 723 786
rect 111 738 115 742
rect 135 738 139 742
rect 759 782 763 786
rect 767 782 771 786
rect 799 782 803 786
rect 863 822 867 826
rect 903 822 907 826
rect 911 822 915 826
rect 935 822 939 826
rect 967 822 971 826
rect 983 822 987 826
rect 991 822 995 826
rect 1015 822 1019 826
rect 1039 822 1043 826
rect 1047 822 1051 826
rect 1063 822 1067 826
rect 1095 822 1099 826
rect 1103 822 1107 826
rect 1127 822 1131 826
rect 815 782 819 786
rect 839 782 843 786
rect 863 782 867 786
rect 879 782 883 786
rect 903 782 907 786
rect 919 782 923 786
rect 935 782 939 786
rect 959 782 963 786
rect 159 738 163 742
rect 183 738 187 742
rect 215 738 219 742
rect 223 738 227 742
rect 263 738 267 742
rect 279 738 283 742
rect 319 738 323 742
rect 343 738 347 742
rect 375 738 379 742
rect 407 738 411 742
rect 423 738 427 742
rect 463 738 467 742
rect 471 738 475 742
rect 519 738 523 742
rect 567 738 571 742
rect 575 738 579 742
rect 615 738 619 742
rect 623 738 627 742
rect 663 738 667 742
rect 671 738 675 742
rect 703 738 707 742
rect 719 738 723 742
rect 751 738 755 742
rect 759 738 763 742
rect 967 782 971 786
rect 991 782 995 786
rect 1015 782 1019 786
rect 1023 782 1027 786
rect 1039 782 1043 786
rect 1055 782 1059 786
rect 1063 782 1067 786
rect 1087 782 1091 786
rect 1095 782 1099 786
rect 1127 782 1131 786
rect 1415 902 1419 906
rect 1447 902 1451 906
rect 1207 862 1211 866
rect 1231 862 1235 866
rect 1247 862 1251 866
rect 1279 862 1283 866
rect 1295 862 1299 866
rect 1327 862 1331 866
rect 1343 862 1347 866
rect 1383 862 1387 866
rect 1391 862 1395 866
rect 1415 862 1419 866
rect 1447 862 1451 866
rect 1159 822 1163 826
rect 1167 822 1171 826
rect 1207 822 1211 826
rect 1247 822 1251 826
rect 1255 822 1259 826
rect 1295 822 1299 826
rect 1311 822 1315 826
rect 1343 822 1347 826
rect 1375 822 1379 826
rect 1391 822 1395 826
rect 1415 822 1419 826
rect 1447 822 1451 826
rect 1167 782 1171 786
rect 1175 782 1179 786
rect 1207 782 1211 786
rect 1231 782 1235 786
rect 1255 782 1259 786
rect 1295 782 1299 786
rect 1311 782 1315 786
rect 1367 782 1371 786
rect 1375 782 1379 786
rect 1415 782 1419 786
rect 1447 782 1451 786
rect 799 738 803 742
rect 807 738 811 742
rect 839 738 843 742
rect 871 738 875 742
rect 879 738 883 742
rect 919 738 923 742
rect 943 738 947 742
rect 959 738 963 742
rect 991 738 995 742
rect 1015 738 1019 742
rect 1023 738 1027 742
rect 1055 738 1059 742
rect 1087 738 1091 742
rect 1127 738 1131 742
rect 1151 738 1155 742
rect 1175 738 1179 742
rect 1215 738 1219 742
rect 1231 738 1235 742
rect 1271 738 1275 742
rect 1295 738 1299 742
rect 1327 738 1331 742
rect 1367 738 1371 742
rect 111 698 115 702
rect 135 698 139 702
rect 159 698 163 702
rect 183 698 187 702
rect 199 698 203 702
rect 215 698 219 702
rect 239 698 243 702
rect 263 698 267 702
rect 287 698 291 702
rect 319 698 323 702
rect 335 698 339 702
rect 375 698 379 702
rect 391 698 395 702
rect 423 698 427 702
rect 439 698 443 702
rect 471 698 475 702
rect 487 698 491 702
rect 519 698 523 702
rect 111 658 115 662
rect 135 658 139 662
rect 159 658 163 662
rect 191 658 195 662
rect 199 658 203 662
rect 215 658 219 662
rect 239 658 243 662
rect 263 658 267 662
rect 287 658 291 662
rect 295 658 299 662
rect 327 658 331 662
rect 335 658 339 662
rect 203 632 207 636
rect 367 658 371 662
rect 391 658 395 662
rect 407 658 411 662
rect 535 698 539 702
rect 567 698 571 702
rect 583 698 587 702
rect 615 698 619 702
rect 639 698 643 702
rect 663 698 667 702
rect 695 698 699 702
rect 703 698 707 702
rect 751 698 755 702
rect 759 698 763 702
rect 807 698 811 702
rect 831 698 835 702
rect 871 698 875 702
rect 439 658 443 662
rect 455 658 459 662
rect 487 658 491 662
rect 503 658 507 662
rect 535 658 539 662
rect 551 658 555 662
rect 583 658 587 662
rect 607 658 611 662
rect 639 658 643 662
rect 347 632 351 636
rect 447 632 451 636
rect 531 632 535 636
rect 663 658 667 662
rect 695 658 699 662
rect 719 658 723 662
rect 759 658 763 662
rect 767 658 771 662
rect 815 658 819 662
rect 831 658 835 662
rect 903 698 907 702
rect 943 698 947 702
rect 967 698 971 702
rect 1015 698 1019 702
rect 1031 698 1035 702
rect 1087 698 1091 702
rect 1135 698 1139 702
rect 1151 698 1155 702
rect 1175 698 1179 702
rect 1215 698 1219 702
rect 1247 698 1251 702
rect 1271 698 1275 702
rect 1279 698 1283 702
rect 1383 738 1387 742
rect 1415 738 1419 742
rect 1447 738 1451 742
rect 1311 698 1315 702
rect 1327 698 1331 702
rect 1343 698 1347 702
rect 1367 698 1371 702
rect 1383 698 1387 702
rect 1391 698 1395 702
rect 1415 698 1419 702
rect 1447 698 1451 702
rect 863 658 867 662
rect 903 658 907 662
rect 935 658 939 662
rect 967 658 971 662
rect 1007 658 1011 662
rect 1031 658 1035 662
rect 1047 658 1051 662
rect 1087 658 1091 662
rect 1127 658 1131 662
rect 1135 658 1139 662
rect 1159 658 1163 662
rect 1175 658 1179 662
rect 1191 658 1195 662
rect 1215 658 1219 662
rect 1223 658 1227 662
rect 1247 658 1251 662
rect 1263 658 1267 662
rect 1279 658 1283 662
rect 1303 658 1307 662
rect 1311 658 1315 662
rect 1343 658 1347 662
rect 1367 658 1371 662
rect 1391 658 1395 662
rect 1415 658 1419 662
rect 1447 658 1451 662
rect 111 618 115 622
rect 191 618 195 622
rect 215 618 219 622
rect 239 618 243 622
rect 263 618 267 622
rect 271 618 275 622
rect 295 618 299 622
rect 319 618 323 622
rect 327 618 331 622
rect 343 618 347 622
rect 367 618 371 622
rect 391 618 395 622
rect 407 618 411 622
rect 415 618 419 622
rect 439 618 443 622
rect 455 618 459 622
rect 479 618 483 622
rect 503 618 507 622
rect 519 618 523 622
rect 111 578 115 582
rect 263 578 267 582
rect 271 578 275 582
rect 287 578 291 582
rect 295 578 299 582
rect 311 578 315 582
rect 319 578 323 582
rect 335 578 339 582
rect 343 578 347 582
rect 359 578 363 582
rect 367 578 371 582
rect 383 578 387 582
rect 391 578 395 582
rect 407 578 411 582
rect 415 578 419 582
rect 111 538 115 542
rect 223 538 227 542
rect 247 538 251 542
rect 263 538 267 542
rect 271 538 275 542
rect 287 538 291 542
rect 295 538 299 542
rect 311 538 315 542
rect 327 538 331 542
rect 335 538 339 542
rect 359 538 363 542
rect 383 538 387 542
rect 391 538 395 542
rect 431 578 435 582
rect 439 578 443 582
rect 551 618 555 622
rect 567 618 571 622
rect 607 618 611 622
rect 623 618 627 622
rect 663 618 667 622
rect 679 618 683 622
rect 719 618 723 622
rect 735 618 739 622
rect 767 618 771 622
rect 783 618 787 622
rect 815 618 819 622
rect 831 618 835 622
rect 863 618 867 622
rect 879 618 883 622
rect 903 618 907 622
rect 927 618 931 622
rect 935 618 939 622
rect 967 618 971 622
rect 975 618 979 622
rect 1007 618 1011 622
rect 1023 618 1027 622
rect 1047 618 1051 622
rect 463 578 467 582
rect 479 578 483 582
rect 503 578 507 582
rect 519 578 523 582
rect 551 578 555 582
rect 567 578 571 582
rect 607 578 611 582
rect 623 578 627 582
rect 663 578 667 582
rect 679 578 683 582
rect 719 578 723 582
rect 735 578 739 582
rect 775 578 779 582
rect 783 578 787 582
rect 1071 618 1075 622
rect 1087 618 1091 622
rect 1111 618 1115 622
rect 1127 618 1131 622
rect 1151 618 1155 622
rect 1159 618 1163 622
rect 1191 618 1195 622
rect 1223 618 1227 622
rect 1239 618 1243 622
rect 1263 618 1267 622
rect 1287 618 1291 622
rect 1303 618 1307 622
rect 1335 618 1339 622
rect 1343 618 1347 622
rect 1447 618 1451 622
rect 831 578 835 582
rect 407 538 411 542
rect 423 538 427 542
rect 431 538 435 542
rect 455 538 459 542
rect 463 538 467 542
rect 487 538 491 542
rect 503 538 507 542
rect 111 498 115 502
rect 135 498 139 502
rect 159 498 163 502
rect 183 498 187 502
rect 223 498 227 502
rect 247 498 251 502
rect 271 498 275 502
rect 295 498 299 502
rect 319 498 323 502
rect 327 498 331 502
rect 359 498 363 502
rect 375 498 379 502
rect 391 498 395 502
rect 423 498 427 502
rect 431 498 435 502
rect 111 458 115 462
rect 135 458 139 462
rect 159 458 163 462
rect 183 458 187 462
rect 191 458 195 462
rect 223 458 227 462
rect 239 458 243 462
rect 271 458 275 462
rect 295 458 299 462
rect 319 458 323 462
rect 351 458 355 462
rect 527 538 531 542
rect 879 578 883 582
rect 887 578 891 582
rect 927 578 931 582
rect 943 578 947 582
rect 975 578 979 582
rect 1007 578 1011 582
rect 1023 578 1027 582
rect 1071 578 1075 582
rect 1111 578 1115 582
rect 1127 578 1131 582
rect 1151 578 1155 582
rect 1183 578 1187 582
rect 1191 578 1195 582
rect 1239 578 1243 582
rect 1247 578 1251 582
rect 1287 578 1291 582
rect 1311 578 1315 582
rect 1335 578 1339 582
rect 1375 578 1379 582
rect 551 538 555 542
rect 575 538 579 542
rect 607 538 611 542
rect 623 538 627 542
rect 663 538 667 542
rect 671 538 675 542
rect 711 538 715 542
rect 719 538 723 542
rect 759 538 763 542
rect 775 538 779 542
rect 807 538 811 542
rect 831 538 835 542
rect 855 538 859 542
rect 887 538 891 542
rect 911 538 915 542
rect 943 538 947 542
rect 967 538 971 542
rect 1007 538 1011 542
rect 1023 538 1027 542
rect 1071 538 1075 542
rect 1079 538 1083 542
rect 1127 538 1131 542
rect 1175 538 1179 542
rect 1183 538 1187 542
rect 1223 538 1227 542
rect 1247 538 1251 542
rect 1271 538 1275 542
rect 1447 578 1451 582
rect 1311 538 1315 542
rect 1351 538 1355 542
rect 1375 538 1379 542
rect 455 498 459 502
rect 487 498 491 502
rect 527 498 531 502
rect 543 498 547 502
rect 575 498 579 502
rect 591 498 595 502
rect 623 498 627 502
rect 631 498 635 502
rect 663 498 667 502
rect 671 498 675 502
rect 687 498 691 502
rect 711 498 715 502
rect 719 498 723 502
rect 759 498 763 502
rect 799 498 803 502
rect 807 498 811 502
rect 847 498 851 502
rect 855 498 859 502
rect 903 498 907 502
rect 911 498 915 502
rect 951 498 955 502
rect 967 498 971 502
rect 999 498 1003 502
rect 1023 498 1027 502
rect 1047 498 1051 502
rect 1079 498 1083 502
rect 1095 498 1099 502
rect 1127 498 1131 502
rect 1143 498 1147 502
rect 1175 498 1179 502
rect 1199 498 1203 502
rect 1223 498 1227 502
rect 1255 498 1259 502
rect 1271 498 1275 502
rect 1391 538 1395 542
rect 1415 538 1419 542
rect 1447 538 1451 542
rect 1311 498 1315 502
rect 1351 498 1355 502
rect 1375 498 1379 502
rect 1391 498 1395 502
rect 1415 498 1419 502
rect 375 458 379 462
rect 415 458 419 462
rect 431 458 435 462
rect 479 458 483 462
rect 487 458 491 462
rect 543 458 547 462
rect 591 458 595 462
rect 607 458 611 462
rect 631 458 635 462
rect 663 458 667 462
rect 671 458 675 462
rect 687 458 691 462
rect 719 458 723 462
rect 111 418 115 422
rect 135 418 139 422
rect 159 418 163 422
rect 183 418 187 422
rect 191 418 195 422
rect 215 418 219 422
rect 239 418 243 422
rect 271 418 275 422
rect 295 418 299 422
rect 327 418 331 422
rect 351 418 355 422
rect 391 418 395 422
rect 415 418 419 422
rect 447 418 451 422
rect 479 418 483 422
rect 503 418 507 422
rect 543 418 547 422
rect 551 418 555 422
rect 599 418 603 422
rect 607 418 611 422
rect 735 458 739 462
rect 759 458 763 462
rect 791 458 795 462
rect 799 458 803 462
rect 839 458 843 462
rect 847 458 851 462
rect 879 458 883 462
rect 903 458 907 462
rect 911 458 915 462
rect 943 458 947 462
rect 951 458 955 462
rect 967 458 971 462
rect 999 458 1003 462
rect 1031 458 1035 462
rect 1047 458 1051 462
rect 1071 458 1075 462
rect 1095 458 1099 462
rect 1119 458 1123 462
rect 1143 458 1147 462
rect 1175 458 1179 462
rect 1199 458 1203 462
rect 1239 458 1243 462
rect 1255 458 1259 462
rect 1303 458 1307 462
rect 1311 458 1315 462
rect 1367 458 1371 462
rect 1375 458 1379 462
rect 1447 498 1451 502
rect 1415 458 1419 462
rect 1447 458 1451 462
rect 647 418 651 422
rect 671 418 675 422
rect 703 418 707 422
rect 735 418 739 422
rect 767 418 771 422
rect 791 418 795 422
rect 831 418 835 422
rect 839 418 843 422
rect 879 418 883 422
rect 903 418 907 422
rect 911 418 915 422
rect 943 418 947 422
rect 967 418 971 422
rect 975 418 979 422
rect 111 374 115 378
rect 135 374 139 378
rect 159 374 163 378
rect 183 374 187 378
rect 207 374 211 378
rect 215 374 219 378
rect 231 374 235 378
rect 255 374 259 378
rect 271 374 275 378
rect 295 374 299 378
rect 327 374 331 378
rect 335 374 339 378
rect 375 374 379 378
rect 391 374 395 378
rect 415 374 419 378
rect 447 374 451 378
rect 455 374 459 378
rect 495 374 499 378
rect 503 374 507 378
rect 535 374 539 378
rect 551 374 555 378
rect 575 374 579 378
rect 599 374 603 378
rect 615 374 619 378
rect 647 374 651 378
rect 655 374 659 378
rect 687 374 691 378
rect 111 334 115 338
rect 135 334 139 338
rect 159 334 163 338
rect 175 334 179 338
rect 183 334 187 338
rect 199 334 203 338
rect 207 334 211 338
rect 223 334 227 338
rect 231 334 235 338
rect 247 334 251 338
rect 255 334 259 338
rect 279 334 283 338
rect 295 334 299 338
rect 319 334 323 338
rect 335 334 339 338
rect 187 312 191 316
rect 359 334 363 338
rect 375 334 379 338
rect 399 334 403 338
rect 347 312 351 316
rect 415 334 419 338
rect 439 334 443 338
rect 455 334 459 338
rect 479 334 483 338
rect 495 334 499 338
rect 527 334 531 338
rect 535 334 539 338
rect 575 334 579 338
rect 583 334 587 338
rect 615 334 619 338
rect 703 374 707 378
rect 727 374 731 378
rect 999 418 1003 422
rect 1031 418 1035 422
rect 1039 418 1043 422
rect 1071 418 1075 422
rect 1103 418 1107 422
rect 1119 418 1123 422
rect 1159 418 1163 422
rect 1175 418 1179 422
rect 1207 418 1211 422
rect 1239 418 1243 422
rect 1247 418 1251 422
rect 767 374 771 378
rect 775 374 779 378
rect 831 374 835 378
rect 887 374 891 378
rect 903 374 907 378
rect 951 374 955 378
rect 975 374 979 378
rect 1015 374 1019 378
rect 1039 374 1043 378
rect 1079 374 1083 378
rect 1103 374 1107 378
rect 1135 374 1139 378
rect 1159 374 1163 378
rect 1183 374 1187 378
rect 1207 374 1211 378
rect 1231 374 1235 378
rect 1279 418 1283 422
rect 1303 418 1307 422
rect 1319 418 1323 422
rect 1359 418 1363 422
rect 1367 418 1371 422
rect 1391 418 1395 422
rect 1415 418 1419 422
rect 1447 418 1451 422
rect 1247 374 1251 378
rect 1271 374 1275 378
rect 1279 374 1283 378
rect 1311 374 1315 378
rect 1319 374 1323 378
rect 1351 374 1355 378
rect 1359 374 1363 378
rect 639 334 643 338
rect 655 334 659 338
rect 687 334 691 338
rect 727 334 731 338
rect 735 334 739 338
rect 775 334 779 338
rect 791 334 795 338
rect 831 334 835 338
rect 847 334 851 338
rect 887 334 891 338
rect 895 334 899 338
rect 943 334 947 338
rect 951 334 955 338
rect 991 334 995 338
rect 1015 334 1019 338
rect 1039 334 1043 338
rect 1079 334 1083 338
rect 1087 334 1091 338
rect 1135 334 1139 338
rect 1183 334 1187 338
rect 1231 334 1235 338
rect 1271 334 1275 338
rect 1279 334 1283 338
rect 1391 374 1395 378
rect 1415 374 1419 378
rect 1447 374 1451 378
rect 1311 334 1315 338
rect 1327 334 1331 338
rect 1351 334 1355 338
rect 1383 334 1387 338
rect 1391 334 1395 338
rect 111 294 115 298
rect 175 294 179 298
rect 199 294 203 298
rect 223 294 227 298
rect 247 294 251 298
rect 271 294 275 298
rect 279 294 283 298
rect 295 294 299 298
rect 319 294 323 298
rect 343 294 347 298
rect 359 294 363 298
rect 367 294 371 298
rect 399 294 403 298
rect 431 294 435 298
rect 439 294 443 298
rect 471 294 475 298
rect 479 294 483 298
rect 511 294 515 298
rect 527 294 531 298
rect 559 294 563 298
rect 583 294 587 298
rect 615 294 619 298
rect 639 294 643 298
rect 663 294 667 298
rect 687 294 691 298
rect 711 294 715 298
rect 735 294 739 298
rect 759 294 763 298
rect 791 294 795 298
rect 279 264 283 268
rect 111 254 115 258
rect 247 254 251 258
rect 263 254 267 258
rect 271 254 275 258
rect 411 267 415 268
rect 411 264 415 267
rect 287 254 291 258
rect 295 254 299 258
rect 311 254 315 258
rect 319 254 323 258
rect 335 254 339 258
rect 343 254 347 258
rect 359 254 363 258
rect 367 254 371 258
rect 383 254 387 258
rect 399 254 403 258
rect 407 254 411 258
rect 111 214 115 218
rect 239 214 243 218
rect 263 214 267 218
rect 287 214 291 218
rect 311 214 315 218
rect 335 214 339 218
rect 359 214 363 218
rect 383 214 387 218
rect 431 254 435 258
rect 463 254 467 258
rect 471 254 475 258
rect 503 254 507 258
rect 511 254 515 258
rect 543 254 547 258
rect 559 254 563 258
rect 583 254 587 258
rect 615 254 619 258
rect 623 254 627 258
rect 663 254 667 258
rect 679 254 683 258
rect 711 254 715 258
rect 807 294 811 298
rect 847 294 851 298
rect 879 294 883 298
rect 895 294 899 298
rect 903 294 907 298
rect 927 294 931 298
rect 943 294 947 298
rect 951 294 955 298
rect 975 294 979 298
rect 991 294 995 298
rect 999 294 1003 298
rect 1023 294 1027 298
rect 1039 294 1043 298
rect 1047 294 1051 298
rect 1071 294 1075 298
rect 1087 294 1091 298
rect 1095 294 1099 298
rect 1127 294 1131 298
rect 1135 294 1139 298
rect 1159 294 1163 298
rect 1183 294 1187 298
rect 1199 294 1203 298
rect 1231 294 1235 298
rect 1247 294 1251 298
rect 1415 334 1419 338
rect 1447 334 1451 338
rect 1279 294 1283 298
rect 1303 294 1307 298
rect 1327 294 1331 298
rect 1367 294 1371 298
rect 743 254 747 258
rect 759 254 763 258
rect 807 254 811 258
rect 847 254 851 258
rect 879 254 883 258
rect 903 254 907 258
rect 927 254 931 258
rect 951 254 955 258
rect 959 254 963 258
rect 975 254 979 258
rect 999 254 1003 258
rect 1023 254 1027 258
rect 1039 254 1043 258
rect 1047 254 1051 258
rect 1071 254 1075 258
rect 1095 254 1099 258
rect 1119 254 1123 258
rect 1127 254 1131 258
rect 1159 254 1163 258
rect 1199 254 1203 258
rect 1247 254 1251 258
rect 1279 254 1283 258
rect 1303 254 1307 258
rect 1383 294 1387 298
rect 1415 294 1419 298
rect 1447 294 1451 298
rect 1359 254 1363 258
rect 1367 254 1371 258
rect 1415 254 1419 258
rect 1447 254 1451 258
rect 407 214 411 218
rect 431 214 435 218
rect 463 214 467 218
rect 503 214 507 218
rect 511 214 515 218
rect 543 214 547 218
rect 559 214 563 218
rect 583 214 587 218
rect 419 203 423 204
rect 419 200 423 203
rect 615 214 619 218
rect 623 214 627 218
rect 671 214 675 218
rect 679 214 683 218
rect 719 214 723 218
rect 743 214 747 218
rect 591 200 595 204
rect 767 214 771 218
rect 807 214 811 218
rect 815 214 819 218
rect 863 214 867 218
rect 879 214 883 218
rect 919 214 923 218
rect 959 214 963 218
rect 975 214 979 218
rect 1031 214 1035 218
rect 1039 214 1043 218
rect 1087 214 1091 218
rect 1119 214 1123 218
rect 1135 214 1139 218
rect 1183 214 1187 218
rect 1199 214 1203 218
rect 1231 214 1235 218
rect 1279 214 1283 218
rect 1327 214 1331 218
rect 1359 214 1363 218
rect 1383 214 1387 218
rect 1415 214 1419 218
rect 1447 214 1451 218
rect 111 174 115 178
rect 183 174 187 178
rect 207 174 211 178
rect 239 174 243 178
rect 263 174 267 178
rect 279 174 283 178
rect 287 174 291 178
rect 311 174 315 178
rect 327 174 331 178
rect 335 174 339 178
rect 359 174 363 178
rect 375 174 379 178
rect 383 174 387 178
rect 407 174 411 178
rect 423 174 427 178
rect 431 174 435 178
rect 463 174 467 178
rect 471 174 475 178
rect 511 174 515 178
rect 527 174 531 178
rect 559 174 563 178
rect 591 174 595 178
rect 615 174 619 178
rect 655 174 659 178
rect 671 174 675 178
rect 111 122 115 126
rect 135 122 139 126
rect 159 122 163 126
rect 183 122 187 126
rect 207 122 211 126
rect 231 122 235 126
rect 239 122 243 126
rect 255 122 259 126
rect 279 122 283 126
rect 303 122 307 126
rect 327 122 331 126
rect 351 122 355 126
rect 375 122 379 126
rect 399 122 403 126
rect 711 174 715 178
rect 719 174 723 178
rect 767 174 771 178
rect 815 174 819 178
rect 823 174 827 178
rect 863 174 867 178
rect 871 174 875 178
rect 919 174 923 178
rect 975 174 979 178
rect 1031 174 1035 178
rect 1079 174 1083 178
rect 1087 174 1091 178
rect 1127 174 1131 178
rect 1135 174 1139 178
rect 1175 174 1179 178
rect 1183 174 1187 178
rect 1223 174 1227 178
rect 1231 174 1235 178
rect 1263 174 1267 178
rect 423 122 427 126
rect 431 122 435 126
rect 463 122 467 126
rect 471 122 475 126
rect 487 122 491 126
rect 511 122 515 126
rect 527 122 531 126
rect 535 122 539 126
rect 559 122 563 126
rect 583 122 587 126
rect 591 122 595 126
rect 607 122 611 126
rect 631 122 635 126
rect 655 122 659 126
rect 679 122 683 126
rect 703 122 707 126
rect 711 122 715 126
rect 727 122 731 126
rect 751 122 755 126
rect 767 122 771 126
rect 775 122 779 126
rect 799 122 803 126
rect 823 122 827 126
rect 855 122 859 126
rect 871 122 875 126
rect 887 122 891 126
rect 919 122 923 126
rect 951 122 955 126
rect 975 122 979 126
rect 983 122 987 126
rect 1015 122 1019 126
rect 111 82 115 86
rect 135 82 139 86
rect 159 82 163 86
rect 183 82 187 86
rect 207 82 211 86
rect 231 82 235 86
rect 1031 122 1035 126
rect 1047 122 1051 126
rect 1279 174 1283 178
rect 1295 174 1299 178
rect 1327 174 1331 178
rect 1359 174 1363 178
rect 1383 174 1387 178
rect 1391 174 1395 178
rect 1415 174 1419 178
rect 1071 122 1075 126
rect 1079 122 1083 126
rect 1095 122 1099 126
rect 1119 122 1123 126
rect 1127 122 1131 126
rect 1143 122 1147 126
rect 1175 122 1179 126
rect 1207 122 1211 126
rect 1223 122 1227 126
rect 1239 122 1243 126
rect 1263 122 1267 126
rect 1271 122 1275 126
rect 1295 122 1299 126
rect 1303 122 1307 126
rect 1327 122 1331 126
rect 1335 122 1339 126
rect 1359 122 1363 126
rect 1367 122 1371 126
rect 1447 174 1451 178
rect 1391 122 1395 126
rect 1415 122 1419 126
rect 1447 122 1451 126
rect 255 82 259 86
rect 279 82 283 86
rect 303 82 307 86
rect 327 82 331 86
rect 351 82 355 86
rect 375 82 379 86
rect 399 82 403 86
rect 431 82 435 86
rect 463 82 467 86
rect 487 82 491 86
rect 511 82 515 86
rect 535 82 539 86
rect 559 82 563 86
rect 583 82 587 86
rect 607 82 611 86
rect 631 82 635 86
rect 655 82 659 86
rect 679 82 683 86
rect 703 82 707 86
rect 727 82 731 86
rect 751 82 755 86
rect 775 82 779 86
rect 799 82 803 86
rect 823 82 827 86
rect 855 82 859 86
rect 887 82 891 86
rect 919 82 923 86
rect 951 82 955 86
rect 983 82 987 86
rect 1015 82 1019 86
rect 1047 82 1051 86
rect 1071 82 1075 86
rect 1095 82 1099 86
rect 1119 82 1123 86
rect 1143 82 1147 86
rect 1175 82 1179 86
rect 1207 82 1211 86
rect 1239 82 1243 86
rect 1271 82 1275 86
rect 1303 82 1307 86
rect 1335 82 1339 86
rect 1367 82 1371 86
rect 1391 82 1395 86
rect 1415 82 1419 86
rect 1447 82 1451 86
<< m4 >>
rect 96 1505 97 1511
rect 103 1510 1483 1511
rect 103 1506 111 1510
rect 115 1506 295 1510
rect 299 1506 319 1510
rect 323 1506 343 1510
rect 347 1506 367 1510
rect 371 1506 407 1510
rect 411 1506 455 1510
rect 459 1506 511 1510
rect 515 1506 575 1510
rect 579 1506 647 1510
rect 651 1506 727 1510
rect 731 1506 807 1510
rect 811 1506 887 1510
rect 891 1506 959 1510
rect 963 1506 1031 1510
rect 1035 1506 1103 1510
rect 1107 1506 1175 1510
rect 1179 1506 1247 1510
rect 1251 1506 1447 1510
rect 1451 1506 1483 1510
rect 103 1505 1483 1506
rect 1489 1505 1490 1511
rect 84 1465 85 1471
rect 91 1470 1471 1471
rect 91 1466 111 1470
rect 115 1466 151 1470
rect 155 1466 175 1470
rect 179 1466 199 1470
rect 203 1466 231 1470
rect 235 1466 271 1470
rect 275 1466 295 1470
rect 299 1466 319 1470
rect 323 1466 343 1470
rect 347 1466 367 1470
rect 371 1466 407 1470
rect 411 1466 455 1470
rect 459 1466 503 1470
rect 507 1466 511 1470
rect 515 1466 551 1470
rect 555 1466 575 1470
rect 579 1466 607 1470
rect 611 1466 647 1470
rect 651 1466 663 1470
rect 667 1466 711 1470
rect 715 1466 727 1470
rect 731 1466 759 1470
rect 763 1466 807 1470
rect 811 1466 815 1470
rect 819 1466 871 1470
rect 875 1466 887 1470
rect 891 1466 927 1470
rect 931 1466 959 1470
rect 963 1466 975 1470
rect 979 1466 1023 1470
rect 1027 1466 1031 1470
rect 1035 1466 1071 1470
rect 1075 1466 1103 1470
rect 1107 1466 1119 1470
rect 1123 1466 1167 1470
rect 1171 1466 1175 1470
rect 1179 1466 1215 1470
rect 1219 1466 1247 1470
rect 1251 1466 1263 1470
rect 1267 1466 1311 1470
rect 1315 1466 1447 1470
rect 1451 1466 1471 1470
rect 91 1465 1471 1466
rect 1477 1465 1478 1471
rect 96 1425 97 1431
rect 103 1430 1483 1431
rect 103 1426 111 1430
rect 115 1426 135 1430
rect 139 1426 151 1430
rect 155 1426 159 1430
rect 163 1426 175 1430
rect 179 1426 183 1430
rect 187 1426 199 1430
rect 203 1426 223 1430
rect 227 1426 231 1430
rect 235 1426 271 1430
rect 275 1426 287 1430
rect 291 1426 319 1430
rect 323 1426 351 1430
rect 355 1426 367 1430
rect 371 1426 407 1430
rect 411 1426 415 1430
rect 419 1426 455 1430
rect 459 1426 479 1430
rect 483 1426 503 1430
rect 507 1426 535 1430
rect 539 1426 551 1430
rect 555 1426 583 1430
rect 587 1426 607 1430
rect 611 1426 631 1430
rect 635 1426 663 1430
rect 667 1426 687 1430
rect 691 1426 711 1430
rect 715 1426 743 1430
rect 747 1426 759 1430
rect 763 1426 799 1430
rect 803 1426 815 1430
rect 819 1426 855 1430
rect 859 1426 871 1430
rect 875 1426 911 1430
rect 915 1426 927 1430
rect 931 1426 967 1430
rect 971 1426 975 1430
rect 979 1426 1023 1430
rect 1027 1426 1071 1430
rect 1075 1426 1119 1430
rect 1123 1426 1167 1430
rect 1171 1426 1215 1430
rect 1219 1426 1263 1430
rect 1267 1426 1303 1430
rect 1307 1426 1311 1430
rect 1315 1426 1343 1430
rect 1347 1426 1391 1430
rect 1395 1426 1415 1430
rect 1419 1426 1447 1430
rect 1451 1426 1483 1430
rect 103 1425 1483 1426
rect 1489 1425 1490 1431
rect 84 1385 85 1391
rect 91 1390 1471 1391
rect 91 1386 111 1390
rect 115 1386 135 1390
rect 139 1386 159 1390
rect 163 1386 183 1390
rect 187 1386 223 1390
rect 227 1386 231 1390
rect 235 1386 279 1390
rect 283 1386 287 1390
rect 291 1386 335 1390
rect 339 1386 351 1390
rect 355 1386 391 1390
rect 395 1386 415 1390
rect 419 1386 439 1390
rect 443 1386 479 1390
rect 483 1386 487 1390
rect 491 1386 527 1390
rect 531 1386 535 1390
rect 539 1386 567 1390
rect 571 1386 583 1390
rect 587 1386 615 1390
rect 619 1386 631 1390
rect 635 1386 663 1390
rect 667 1386 687 1390
rect 691 1386 711 1390
rect 715 1386 743 1390
rect 747 1386 767 1390
rect 771 1386 799 1390
rect 803 1386 823 1390
rect 827 1386 855 1390
rect 859 1386 879 1390
rect 883 1386 911 1390
rect 915 1386 935 1390
rect 939 1386 967 1390
rect 971 1386 991 1390
rect 995 1386 1023 1390
rect 1027 1386 1047 1390
rect 1051 1386 1071 1390
rect 1075 1386 1095 1390
rect 1099 1386 1119 1390
rect 1123 1386 1143 1390
rect 1147 1386 1167 1390
rect 1171 1386 1191 1390
rect 1195 1386 1215 1390
rect 1219 1386 1239 1390
rect 1243 1386 1263 1390
rect 1267 1386 1287 1390
rect 1291 1386 1303 1390
rect 1307 1386 1335 1390
rect 1339 1386 1343 1390
rect 1347 1386 1383 1390
rect 1387 1386 1391 1390
rect 1395 1386 1415 1390
rect 1419 1386 1447 1390
rect 1451 1386 1471 1390
rect 91 1385 1471 1386
rect 1477 1385 1478 1391
rect 96 1345 97 1351
rect 103 1350 1483 1351
rect 103 1346 111 1350
rect 115 1346 135 1350
rect 139 1346 159 1350
rect 163 1346 167 1350
rect 171 1346 183 1350
rect 187 1346 191 1350
rect 195 1346 231 1350
rect 235 1346 279 1350
rect 283 1346 335 1350
rect 339 1346 391 1350
rect 395 1346 439 1350
rect 443 1346 455 1350
rect 459 1346 487 1350
rect 491 1346 519 1350
rect 523 1346 527 1350
rect 531 1346 567 1350
rect 571 1346 575 1350
rect 579 1346 615 1350
rect 619 1346 631 1350
rect 635 1346 663 1350
rect 667 1346 679 1350
rect 683 1346 711 1350
rect 715 1346 727 1350
rect 731 1346 767 1350
rect 771 1346 799 1350
rect 803 1346 823 1350
rect 827 1346 831 1350
rect 835 1346 863 1350
rect 867 1346 879 1350
rect 883 1346 895 1350
rect 899 1346 927 1350
rect 931 1346 935 1350
rect 939 1346 967 1350
rect 971 1346 991 1350
rect 995 1346 1007 1350
rect 1011 1346 1047 1350
rect 1051 1346 1055 1350
rect 1059 1346 1095 1350
rect 1099 1346 1103 1350
rect 1107 1346 1143 1350
rect 1147 1346 1159 1350
rect 1163 1346 1191 1350
rect 1195 1346 1215 1350
rect 1219 1346 1239 1350
rect 1243 1346 1271 1350
rect 1275 1346 1287 1350
rect 1291 1346 1327 1350
rect 1331 1346 1335 1350
rect 1339 1346 1383 1350
rect 1387 1346 1415 1350
rect 1419 1346 1447 1350
rect 1451 1346 1483 1350
rect 103 1345 1483 1346
rect 1489 1345 1490 1351
rect 242 1324 248 1325
rect 326 1324 332 1325
rect 242 1320 243 1324
rect 247 1320 327 1324
rect 331 1320 332 1324
rect 242 1319 248 1320
rect 326 1319 332 1320
rect 84 1305 85 1311
rect 91 1310 1471 1311
rect 91 1306 111 1310
rect 115 1306 167 1310
rect 171 1306 191 1310
rect 195 1306 231 1310
rect 235 1306 255 1310
rect 259 1306 279 1310
rect 283 1306 303 1310
rect 307 1306 327 1310
rect 331 1306 335 1310
rect 339 1306 351 1310
rect 355 1306 375 1310
rect 379 1306 391 1310
rect 395 1306 399 1310
rect 403 1306 423 1310
rect 427 1306 447 1310
rect 451 1306 455 1310
rect 459 1306 471 1310
rect 475 1306 503 1310
rect 507 1306 519 1310
rect 523 1306 543 1310
rect 547 1306 575 1310
rect 579 1306 591 1310
rect 595 1306 631 1310
rect 635 1306 647 1310
rect 651 1306 679 1310
rect 683 1306 695 1310
rect 699 1306 727 1310
rect 731 1306 743 1310
rect 747 1306 767 1310
rect 771 1306 791 1310
rect 795 1306 799 1310
rect 803 1306 831 1310
rect 835 1306 839 1310
rect 843 1306 863 1310
rect 867 1306 879 1310
rect 883 1306 895 1310
rect 899 1306 911 1310
rect 915 1306 927 1310
rect 931 1306 951 1310
rect 955 1306 967 1310
rect 971 1306 991 1310
rect 995 1306 1007 1310
rect 1011 1306 1031 1310
rect 1035 1306 1055 1310
rect 1059 1306 1071 1310
rect 1075 1306 1103 1310
rect 1107 1306 1111 1310
rect 1115 1306 1151 1310
rect 1155 1306 1159 1310
rect 1163 1306 1199 1310
rect 1203 1306 1215 1310
rect 1219 1306 1247 1310
rect 1251 1306 1271 1310
rect 1275 1306 1303 1310
rect 1307 1306 1327 1310
rect 1331 1306 1367 1310
rect 1371 1306 1383 1310
rect 1387 1306 1415 1310
rect 1419 1306 1447 1310
rect 1451 1306 1471 1310
rect 91 1305 1471 1306
rect 1477 1305 1478 1311
rect 96 1265 97 1271
rect 103 1270 1483 1271
rect 103 1266 111 1270
rect 115 1266 231 1270
rect 235 1266 255 1270
rect 259 1266 279 1270
rect 283 1266 303 1270
rect 307 1266 311 1270
rect 315 1266 327 1270
rect 331 1266 335 1270
rect 339 1266 351 1270
rect 355 1266 359 1270
rect 363 1266 375 1270
rect 379 1266 383 1270
rect 387 1266 399 1270
rect 403 1266 415 1270
rect 419 1266 423 1270
rect 427 1266 447 1270
rect 451 1266 471 1270
rect 475 1266 479 1270
rect 483 1266 503 1270
rect 507 1266 519 1270
rect 523 1266 543 1270
rect 547 1266 559 1270
rect 563 1266 591 1270
rect 595 1266 615 1270
rect 619 1266 647 1270
rect 651 1266 679 1270
rect 683 1266 695 1270
rect 699 1266 743 1270
rect 747 1266 751 1270
rect 755 1266 791 1270
rect 795 1266 831 1270
rect 835 1266 839 1270
rect 843 1266 879 1270
rect 883 1266 911 1270
rect 915 1266 951 1270
rect 955 1266 991 1270
rect 995 1266 1031 1270
rect 1035 1266 1063 1270
rect 1067 1266 1071 1270
rect 1075 1266 1111 1270
rect 1115 1266 1127 1270
rect 1131 1266 1151 1270
rect 1155 1266 1191 1270
rect 1195 1266 1199 1270
rect 1203 1266 1247 1270
rect 1251 1266 1303 1270
rect 1307 1266 1311 1270
rect 1315 1266 1367 1270
rect 1371 1266 1375 1270
rect 1379 1266 1415 1270
rect 1419 1266 1447 1270
rect 1451 1266 1483 1270
rect 103 1265 1483 1266
rect 1489 1265 1490 1271
rect 84 1225 85 1231
rect 91 1230 1471 1231
rect 91 1226 111 1230
rect 115 1226 311 1230
rect 315 1226 327 1230
rect 331 1226 335 1230
rect 339 1226 359 1230
rect 363 1226 367 1230
rect 371 1226 383 1230
rect 387 1226 407 1230
rect 411 1226 415 1230
rect 419 1226 447 1230
rect 451 1226 479 1230
rect 483 1226 487 1230
rect 491 1226 519 1230
rect 523 1226 527 1230
rect 531 1226 559 1230
rect 563 1226 567 1230
rect 571 1226 607 1230
rect 611 1226 615 1230
rect 619 1226 655 1230
rect 659 1226 679 1230
rect 683 1226 703 1230
rect 707 1226 751 1230
rect 755 1226 799 1230
rect 803 1226 831 1230
rect 835 1226 847 1230
rect 851 1226 895 1230
rect 899 1226 911 1230
rect 915 1226 943 1230
rect 947 1226 991 1230
rect 995 1226 1039 1230
rect 1043 1226 1063 1230
rect 1067 1226 1103 1230
rect 1107 1226 1127 1230
rect 1131 1226 1175 1230
rect 1179 1226 1191 1230
rect 1195 1226 1247 1230
rect 1251 1226 1255 1230
rect 1259 1226 1311 1230
rect 1315 1226 1343 1230
rect 1347 1226 1375 1230
rect 1379 1226 1415 1230
rect 1419 1226 1447 1230
rect 1451 1226 1471 1230
rect 91 1225 1471 1226
rect 1477 1225 1478 1231
rect 96 1185 97 1191
rect 103 1190 1483 1191
rect 103 1186 111 1190
rect 115 1186 135 1190
rect 139 1186 159 1190
rect 163 1186 183 1190
rect 187 1186 207 1190
rect 211 1186 231 1190
rect 235 1186 255 1190
rect 259 1186 279 1190
rect 283 1186 303 1190
rect 307 1186 327 1190
rect 331 1186 335 1190
rect 339 1186 367 1190
rect 371 1186 383 1190
rect 387 1186 407 1190
rect 411 1186 423 1190
rect 427 1186 447 1190
rect 451 1186 463 1190
rect 467 1186 487 1190
rect 491 1186 503 1190
rect 507 1186 527 1190
rect 531 1186 543 1190
rect 547 1186 567 1190
rect 571 1186 583 1190
rect 587 1186 607 1190
rect 611 1186 623 1190
rect 627 1186 655 1190
rect 659 1186 671 1190
rect 675 1186 703 1190
rect 707 1186 719 1190
rect 723 1186 751 1190
rect 755 1186 767 1190
rect 771 1186 799 1190
rect 803 1186 815 1190
rect 819 1186 847 1190
rect 851 1186 863 1190
rect 867 1186 895 1190
rect 899 1186 911 1190
rect 915 1186 943 1190
rect 947 1186 959 1190
rect 963 1186 991 1190
rect 995 1186 1007 1190
rect 1011 1186 1039 1190
rect 1043 1186 1055 1190
rect 1059 1186 1103 1190
rect 1107 1186 1151 1190
rect 1155 1186 1175 1190
rect 1179 1186 1191 1190
rect 1195 1186 1231 1190
rect 1235 1186 1255 1190
rect 1259 1186 1271 1190
rect 1275 1186 1311 1190
rect 1315 1186 1343 1190
rect 1347 1186 1351 1190
rect 1355 1186 1391 1190
rect 1395 1186 1415 1190
rect 1419 1186 1447 1190
rect 1451 1186 1483 1190
rect 103 1185 1483 1186
rect 1489 1185 1490 1191
rect 84 1145 85 1151
rect 91 1150 1471 1151
rect 91 1146 111 1150
rect 115 1146 135 1150
rect 139 1146 159 1150
rect 163 1146 183 1150
rect 187 1146 207 1150
rect 211 1146 215 1150
rect 219 1146 231 1150
rect 235 1146 255 1150
rect 259 1146 279 1150
rect 283 1146 295 1150
rect 299 1146 303 1150
rect 307 1146 335 1150
rect 339 1146 375 1150
rect 379 1146 383 1150
rect 387 1146 415 1150
rect 419 1146 423 1150
rect 427 1146 463 1150
rect 467 1146 503 1150
rect 507 1146 519 1150
rect 523 1146 543 1150
rect 547 1146 583 1150
rect 587 1146 623 1150
rect 627 1146 647 1150
rect 651 1146 671 1150
rect 675 1146 711 1150
rect 715 1146 719 1150
rect 723 1146 767 1150
rect 771 1146 815 1150
rect 819 1146 831 1150
rect 835 1146 863 1150
rect 867 1146 887 1150
rect 891 1146 911 1150
rect 915 1146 943 1150
rect 947 1146 959 1150
rect 963 1146 999 1150
rect 1003 1146 1007 1150
rect 1011 1146 1055 1150
rect 1059 1146 1103 1150
rect 1107 1146 1151 1150
rect 1155 1146 1191 1150
rect 1195 1146 1231 1150
rect 1235 1146 1271 1150
rect 1275 1146 1311 1150
rect 1315 1146 1351 1150
rect 1355 1146 1391 1150
rect 1395 1146 1415 1150
rect 1419 1146 1447 1150
rect 1451 1146 1471 1150
rect 91 1145 1471 1146
rect 1477 1145 1478 1151
rect 96 1101 97 1107
rect 103 1106 1483 1107
rect 103 1102 111 1106
rect 115 1102 135 1106
rect 139 1102 159 1106
rect 163 1102 183 1106
rect 187 1102 207 1106
rect 211 1102 215 1106
rect 219 1102 247 1106
rect 251 1102 255 1106
rect 259 1102 287 1106
rect 291 1102 295 1106
rect 299 1102 327 1106
rect 331 1102 335 1106
rect 339 1102 367 1106
rect 371 1102 375 1106
rect 379 1102 407 1106
rect 411 1102 415 1106
rect 419 1102 455 1106
rect 459 1102 463 1106
rect 467 1102 503 1106
rect 507 1102 519 1106
rect 523 1102 559 1106
rect 563 1102 583 1106
rect 587 1102 607 1106
rect 611 1102 647 1106
rect 651 1102 655 1106
rect 659 1102 703 1106
rect 707 1102 711 1106
rect 715 1102 743 1106
rect 747 1102 767 1106
rect 771 1102 791 1106
rect 795 1102 831 1106
rect 835 1102 839 1106
rect 843 1102 887 1106
rect 891 1102 943 1106
rect 947 1102 999 1106
rect 1003 1102 1055 1106
rect 1059 1102 1103 1106
rect 1107 1102 1111 1106
rect 1115 1102 1151 1106
rect 1155 1102 1167 1106
rect 1171 1102 1191 1106
rect 1195 1102 1215 1106
rect 1219 1102 1231 1106
rect 1235 1102 1271 1106
rect 1275 1102 1311 1106
rect 1315 1102 1327 1106
rect 1331 1102 1351 1106
rect 1355 1102 1383 1106
rect 1387 1102 1391 1106
rect 1395 1102 1415 1106
rect 1419 1102 1447 1106
rect 1451 1102 1483 1106
rect 103 1101 1483 1102
rect 1489 1101 1490 1107
rect 146 1076 152 1077
rect 218 1076 224 1077
rect 146 1072 147 1076
rect 151 1072 219 1076
rect 223 1072 224 1076
rect 146 1071 152 1072
rect 218 1071 224 1072
rect 84 1061 85 1067
rect 91 1066 1471 1067
rect 91 1062 111 1066
rect 115 1062 135 1066
rect 139 1062 159 1066
rect 163 1062 183 1066
rect 187 1062 207 1066
rect 211 1062 231 1066
rect 235 1062 247 1066
rect 251 1062 271 1066
rect 275 1062 287 1066
rect 291 1062 311 1066
rect 315 1062 327 1066
rect 331 1062 351 1066
rect 355 1062 367 1066
rect 371 1062 391 1066
rect 395 1062 407 1066
rect 411 1062 431 1066
rect 435 1062 455 1066
rect 459 1062 471 1066
rect 475 1062 503 1066
rect 507 1062 511 1066
rect 515 1062 551 1066
rect 555 1062 559 1066
rect 563 1062 591 1066
rect 595 1062 607 1066
rect 611 1062 631 1066
rect 635 1062 655 1066
rect 659 1062 671 1066
rect 675 1062 703 1066
rect 707 1062 711 1066
rect 715 1062 743 1066
rect 747 1062 783 1066
rect 787 1062 791 1066
rect 795 1062 823 1066
rect 827 1062 839 1066
rect 843 1062 871 1066
rect 875 1062 887 1066
rect 891 1062 919 1066
rect 923 1062 943 1066
rect 947 1062 975 1066
rect 979 1062 999 1066
rect 1003 1062 1031 1066
rect 1035 1062 1055 1066
rect 1059 1062 1079 1066
rect 1083 1062 1111 1066
rect 1115 1062 1127 1066
rect 1131 1062 1167 1066
rect 1171 1062 1175 1066
rect 1179 1062 1215 1066
rect 1219 1062 1223 1066
rect 1227 1062 1271 1066
rect 1275 1062 1327 1066
rect 1331 1062 1383 1066
rect 1387 1062 1415 1066
rect 1419 1062 1447 1066
rect 1451 1062 1471 1066
rect 91 1061 1471 1062
rect 1477 1061 1478 1067
rect 146 1044 152 1045
rect 298 1044 304 1045
rect 146 1040 147 1044
rect 151 1040 299 1044
rect 303 1040 304 1044
rect 146 1039 152 1040
rect 298 1039 304 1040
rect 694 1036 700 1037
rect 794 1036 800 1037
rect 694 1032 695 1036
rect 699 1032 795 1036
rect 799 1032 800 1036
rect 694 1031 700 1032
rect 794 1031 800 1032
rect 96 1021 97 1027
rect 103 1026 1483 1027
rect 103 1022 111 1026
rect 115 1022 135 1026
rect 139 1022 159 1026
rect 163 1022 183 1026
rect 187 1022 207 1026
rect 211 1022 231 1026
rect 235 1022 263 1026
rect 267 1022 271 1026
rect 275 1022 303 1026
rect 307 1022 311 1026
rect 315 1022 343 1026
rect 347 1022 351 1026
rect 355 1022 383 1026
rect 387 1022 391 1026
rect 395 1022 431 1026
rect 435 1022 471 1026
rect 475 1022 479 1026
rect 483 1022 511 1026
rect 515 1022 527 1026
rect 531 1022 551 1026
rect 555 1022 575 1026
rect 579 1022 591 1026
rect 595 1022 623 1026
rect 627 1022 631 1026
rect 635 1022 671 1026
rect 675 1022 711 1026
rect 715 1022 719 1026
rect 723 1022 743 1026
rect 747 1022 767 1026
rect 771 1022 783 1026
rect 787 1022 823 1026
rect 827 1022 871 1026
rect 875 1022 879 1026
rect 883 1022 919 1026
rect 923 1022 935 1026
rect 939 1022 975 1026
rect 979 1022 991 1026
rect 995 1022 1031 1026
rect 1035 1022 1047 1026
rect 1051 1022 1079 1026
rect 1083 1022 1103 1026
rect 1107 1022 1127 1026
rect 1131 1022 1159 1026
rect 1163 1022 1175 1026
rect 1179 1022 1215 1026
rect 1219 1022 1223 1026
rect 1227 1022 1271 1026
rect 1275 1022 1327 1026
rect 1331 1022 1383 1026
rect 1387 1022 1415 1026
rect 1419 1022 1447 1026
rect 1451 1022 1483 1026
rect 103 1021 1483 1022
rect 1489 1021 1490 1027
rect 218 996 224 997
rect 354 996 360 997
rect 218 992 219 996
rect 223 992 355 996
rect 359 992 360 996
rect 218 991 224 992
rect 354 991 360 992
rect 84 981 85 987
rect 91 986 1471 987
rect 91 982 111 986
rect 115 982 159 986
rect 163 982 183 986
rect 187 982 207 986
rect 211 982 231 986
rect 235 982 255 986
rect 259 982 263 986
rect 267 982 287 986
rect 291 982 303 986
rect 307 982 327 986
rect 331 982 343 986
rect 347 982 375 986
rect 379 982 383 986
rect 387 982 423 986
rect 427 982 431 986
rect 435 982 471 986
rect 475 982 479 986
rect 483 982 519 986
rect 523 982 527 986
rect 531 982 567 986
rect 571 982 575 986
rect 579 982 623 986
rect 627 982 671 986
rect 675 982 679 986
rect 683 982 719 986
rect 723 982 727 986
rect 731 982 767 986
rect 771 982 775 986
rect 779 982 823 986
rect 827 982 831 986
rect 835 982 879 986
rect 883 982 887 986
rect 891 982 935 986
rect 939 982 943 986
rect 947 982 991 986
rect 995 982 999 986
rect 1003 982 1047 986
rect 1051 982 1095 986
rect 1099 982 1103 986
rect 1107 982 1143 986
rect 1147 982 1159 986
rect 1163 982 1191 986
rect 1195 982 1215 986
rect 1219 982 1239 986
rect 1243 982 1271 986
rect 1275 982 1287 986
rect 1291 982 1327 986
rect 1331 982 1335 986
rect 1339 982 1383 986
rect 1387 982 1415 986
rect 1419 982 1447 986
rect 1451 982 1471 986
rect 91 981 1471 982
rect 1477 981 1478 987
rect 96 941 97 947
rect 103 946 1483 947
rect 103 942 111 946
rect 115 942 207 946
rect 211 942 215 946
rect 219 942 231 946
rect 235 942 239 946
rect 243 942 255 946
rect 259 942 263 946
rect 267 942 287 946
rect 291 942 319 946
rect 323 942 327 946
rect 331 942 351 946
rect 355 942 375 946
rect 379 942 391 946
rect 395 942 423 946
rect 427 942 431 946
rect 435 942 471 946
rect 475 942 519 946
rect 523 942 567 946
rect 571 942 615 946
rect 619 942 623 946
rect 627 942 671 946
rect 675 942 679 946
rect 683 942 727 946
rect 731 942 775 946
rect 779 942 783 946
rect 787 942 831 946
rect 835 942 847 946
rect 851 942 887 946
rect 891 942 919 946
rect 923 942 943 946
rect 947 942 991 946
rect 995 942 999 946
rect 1003 942 1047 946
rect 1051 942 1055 946
rect 1059 942 1095 946
rect 1099 942 1119 946
rect 1123 942 1143 946
rect 1147 942 1175 946
rect 1179 942 1191 946
rect 1195 942 1223 946
rect 1227 942 1239 946
rect 1243 942 1263 946
rect 1267 942 1287 946
rect 1291 942 1295 946
rect 1299 942 1327 946
rect 1331 942 1335 946
rect 1339 942 1359 946
rect 1363 942 1383 946
rect 1387 942 1391 946
rect 1395 942 1415 946
rect 1419 942 1447 946
rect 1451 942 1483 946
rect 103 941 1483 942
rect 1489 941 1490 947
rect 226 932 232 933
rect 302 932 308 933
rect 226 928 227 932
rect 231 928 303 932
rect 307 928 308 932
rect 226 927 232 928
rect 302 927 308 928
rect 442 932 448 933
rect 538 932 544 933
rect 442 928 443 932
rect 447 928 539 932
rect 543 928 544 932
rect 442 927 448 928
rect 538 927 544 928
rect 84 901 85 907
rect 91 906 1471 907
rect 91 902 111 906
rect 115 902 215 906
rect 219 902 231 906
rect 235 902 239 906
rect 243 902 255 906
rect 259 902 263 906
rect 267 902 279 906
rect 283 902 287 906
rect 291 902 303 906
rect 307 902 319 906
rect 323 902 327 906
rect 331 902 351 906
rect 355 902 359 906
rect 363 902 391 906
rect 395 902 423 906
rect 427 902 431 906
rect 435 902 455 906
rect 459 902 471 906
rect 475 902 495 906
rect 499 902 519 906
rect 523 902 535 906
rect 539 902 567 906
rect 571 902 575 906
rect 579 902 615 906
rect 619 902 623 906
rect 627 902 663 906
rect 667 902 671 906
rect 675 902 703 906
rect 707 902 727 906
rect 731 902 751 906
rect 755 902 783 906
rect 787 902 807 906
rect 811 902 847 906
rect 851 902 863 906
rect 867 902 919 906
rect 923 902 927 906
rect 931 902 991 906
rect 995 902 1055 906
rect 1059 902 1119 906
rect 1123 902 1175 906
rect 1179 902 1223 906
rect 1227 902 1231 906
rect 1235 902 1263 906
rect 1267 902 1279 906
rect 1283 902 1295 906
rect 1299 902 1327 906
rect 1331 902 1359 906
rect 1363 902 1383 906
rect 1387 902 1391 906
rect 1395 902 1415 906
rect 1419 902 1447 906
rect 1451 902 1471 906
rect 91 901 1471 902
rect 1477 901 1478 907
rect 96 861 97 867
rect 103 866 1483 867
rect 103 862 111 866
rect 115 862 207 866
rect 211 862 231 866
rect 235 862 255 866
rect 259 862 279 866
rect 283 862 287 866
rect 291 862 303 866
rect 307 862 319 866
rect 323 862 327 866
rect 331 862 351 866
rect 355 862 359 866
rect 363 862 383 866
rect 387 862 391 866
rect 395 862 415 866
rect 419 862 423 866
rect 427 862 447 866
rect 451 862 455 866
rect 459 862 479 866
rect 483 862 495 866
rect 499 862 511 866
rect 515 862 535 866
rect 539 862 551 866
rect 555 862 575 866
rect 579 862 599 866
rect 603 862 623 866
rect 627 862 647 866
rect 651 862 663 866
rect 667 862 703 866
rect 707 862 751 866
rect 755 862 767 866
rect 771 862 807 866
rect 811 862 839 866
rect 843 862 863 866
rect 867 862 911 866
rect 915 862 927 866
rect 931 862 983 866
rect 987 862 991 866
rect 995 862 1047 866
rect 1051 862 1055 866
rect 1059 862 1103 866
rect 1107 862 1119 866
rect 1123 862 1159 866
rect 1163 862 1175 866
rect 1179 862 1207 866
rect 1211 862 1231 866
rect 1235 862 1247 866
rect 1251 862 1279 866
rect 1283 862 1295 866
rect 1299 862 1327 866
rect 1331 862 1343 866
rect 1347 862 1383 866
rect 1387 862 1391 866
rect 1395 862 1415 866
rect 1419 862 1447 866
rect 1451 862 1483 866
rect 103 861 1483 862
rect 1489 861 1490 867
rect 84 821 85 827
rect 91 826 1471 827
rect 91 822 111 826
rect 115 822 135 826
rect 139 822 159 826
rect 163 822 183 826
rect 187 822 207 826
rect 211 822 215 826
rect 219 822 231 826
rect 235 822 255 826
rect 259 822 263 826
rect 267 822 287 826
rect 291 822 311 826
rect 315 822 319 826
rect 323 822 351 826
rect 355 822 367 826
rect 371 822 383 826
rect 387 822 415 826
rect 419 822 431 826
rect 435 822 447 826
rect 451 822 479 826
rect 483 822 487 826
rect 491 822 511 826
rect 515 822 543 826
rect 547 822 551 826
rect 555 822 599 826
rect 603 822 647 826
rect 651 822 655 826
rect 659 822 703 826
rect 707 822 711 826
rect 715 822 767 826
rect 771 822 815 826
rect 819 822 839 826
rect 843 822 863 826
rect 867 822 903 826
rect 907 822 911 826
rect 915 822 935 826
rect 939 822 967 826
rect 971 822 983 826
rect 987 822 991 826
rect 995 822 1015 826
rect 1019 822 1039 826
rect 1043 822 1047 826
rect 1051 822 1063 826
rect 1067 822 1095 826
rect 1099 822 1103 826
rect 1107 822 1127 826
rect 1131 822 1159 826
rect 1163 822 1167 826
rect 1171 822 1207 826
rect 1211 822 1247 826
rect 1251 822 1255 826
rect 1259 822 1295 826
rect 1299 822 1311 826
rect 1315 822 1343 826
rect 1347 822 1375 826
rect 1379 822 1391 826
rect 1395 822 1415 826
rect 1419 822 1447 826
rect 1451 822 1471 826
rect 91 821 1471 822
rect 1477 821 1478 827
rect 96 781 97 787
rect 103 786 1483 787
rect 103 782 111 786
rect 115 782 135 786
rect 139 782 159 786
rect 163 782 183 786
rect 187 782 215 786
rect 219 782 223 786
rect 227 782 263 786
rect 267 782 279 786
rect 283 782 311 786
rect 315 782 343 786
rect 347 782 367 786
rect 371 782 407 786
rect 411 782 431 786
rect 435 782 463 786
rect 467 782 487 786
rect 491 782 519 786
rect 523 782 543 786
rect 547 782 575 786
rect 579 782 599 786
rect 603 782 623 786
rect 627 782 655 786
rect 659 782 671 786
rect 675 782 711 786
rect 715 782 719 786
rect 723 782 759 786
rect 763 782 767 786
rect 771 782 799 786
rect 803 782 815 786
rect 819 782 839 786
rect 843 782 863 786
rect 867 782 879 786
rect 883 782 903 786
rect 907 782 919 786
rect 923 782 935 786
rect 939 782 959 786
rect 963 782 967 786
rect 971 782 991 786
rect 995 782 1015 786
rect 1019 782 1023 786
rect 1027 782 1039 786
rect 1043 782 1055 786
rect 1059 782 1063 786
rect 1067 782 1087 786
rect 1091 782 1095 786
rect 1099 782 1127 786
rect 1131 782 1167 786
rect 1171 782 1175 786
rect 1179 782 1207 786
rect 1211 782 1231 786
rect 1235 782 1255 786
rect 1259 782 1295 786
rect 1299 782 1311 786
rect 1315 782 1367 786
rect 1371 782 1375 786
rect 1379 782 1415 786
rect 1419 782 1447 786
rect 1451 782 1483 786
rect 103 781 1483 782
rect 1489 781 1490 787
rect 84 737 85 743
rect 91 742 1471 743
rect 91 738 111 742
rect 115 738 135 742
rect 139 738 159 742
rect 163 738 183 742
rect 187 738 215 742
rect 219 738 223 742
rect 227 738 263 742
rect 267 738 279 742
rect 283 738 319 742
rect 323 738 343 742
rect 347 738 375 742
rect 379 738 407 742
rect 411 738 423 742
rect 427 738 463 742
rect 467 738 471 742
rect 475 738 519 742
rect 523 738 567 742
rect 571 738 575 742
rect 579 738 615 742
rect 619 738 623 742
rect 627 738 663 742
rect 667 738 671 742
rect 675 738 703 742
rect 707 738 719 742
rect 723 738 751 742
rect 755 738 759 742
rect 763 738 799 742
rect 803 738 807 742
rect 811 738 839 742
rect 843 738 871 742
rect 875 738 879 742
rect 883 738 919 742
rect 923 738 943 742
rect 947 738 959 742
rect 963 738 991 742
rect 995 738 1015 742
rect 1019 738 1023 742
rect 1027 738 1055 742
rect 1059 738 1087 742
rect 1091 738 1127 742
rect 1131 738 1151 742
rect 1155 738 1175 742
rect 1179 738 1215 742
rect 1219 738 1231 742
rect 1235 738 1271 742
rect 1275 738 1295 742
rect 1299 738 1327 742
rect 1331 738 1367 742
rect 1371 738 1383 742
rect 1387 738 1415 742
rect 1419 738 1447 742
rect 1451 738 1471 742
rect 91 737 1471 738
rect 1477 737 1478 743
rect 96 697 97 703
rect 103 702 1483 703
rect 103 698 111 702
rect 115 698 135 702
rect 139 698 159 702
rect 163 698 183 702
rect 187 698 199 702
rect 203 698 215 702
rect 219 698 239 702
rect 243 698 263 702
rect 267 698 287 702
rect 291 698 319 702
rect 323 698 335 702
rect 339 698 375 702
rect 379 698 391 702
rect 395 698 423 702
rect 427 698 439 702
rect 443 698 471 702
rect 475 698 487 702
rect 491 698 519 702
rect 523 698 535 702
rect 539 698 567 702
rect 571 698 583 702
rect 587 698 615 702
rect 619 698 639 702
rect 643 698 663 702
rect 667 698 695 702
rect 699 698 703 702
rect 707 698 751 702
rect 755 698 759 702
rect 763 698 807 702
rect 811 698 831 702
rect 835 698 871 702
rect 875 698 903 702
rect 907 698 943 702
rect 947 698 967 702
rect 971 698 1015 702
rect 1019 698 1031 702
rect 1035 698 1087 702
rect 1091 698 1135 702
rect 1139 698 1151 702
rect 1155 698 1175 702
rect 1179 698 1215 702
rect 1219 698 1247 702
rect 1251 698 1271 702
rect 1275 698 1279 702
rect 1283 698 1311 702
rect 1315 698 1327 702
rect 1331 698 1343 702
rect 1347 698 1367 702
rect 1371 698 1383 702
rect 1387 698 1391 702
rect 1395 698 1415 702
rect 1419 698 1447 702
rect 1451 698 1483 702
rect 103 697 1483 698
rect 1489 697 1490 703
rect 84 657 85 663
rect 91 662 1471 663
rect 91 658 111 662
rect 115 658 135 662
rect 139 658 159 662
rect 163 658 191 662
rect 195 658 199 662
rect 203 658 215 662
rect 219 658 239 662
rect 243 658 263 662
rect 267 658 287 662
rect 291 658 295 662
rect 299 658 327 662
rect 331 658 335 662
rect 339 658 367 662
rect 371 658 391 662
rect 395 658 407 662
rect 411 658 439 662
rect 443 658 455 662
rect 459 658 487 662
rect 491 658 503 662
rect 507 658 535 662
rect 539 658 551 662
rect 555 658 583 662
rect 587 658 607 662
rect 611 658 639 662
rect 643 658 663 662
rect 667 658 695 662
rect 699 658 719 662
rect 723 658 759 662
rect 763 658 767 662
rect 771 658 815 662
rect 819 658 831 662
rect 835 658 863 662
rect 867 658 903 662
rect 907 658 935 662
rect 939 658 967 662
rect 971 658 1007 662
rect 1011 658 1031 662
rect 1035 658 1047 662
rect 1051 658 1087 662
rect 1091 658 1127 662
rect 1131 658 1135 662
rect 1139 658 1159 662
rect 1163 658 1175 662
rect 1179 658 1191 662
rect 1195 658 1215 662
rect 1219 658 1223 662
rect 1227 658 1247 662
rect 1251 658 1263 662
rect 1267 658 1279 662
rect 1283 658 1303 662
rect 1307 658 1311 662
rect 1315 658 1343 662
rect 1347 658 1367 662
rect 1371 658 1391 662
rect 1395 658 1415 662
rect 1419 658 1447 662
rect 1451 658 1471 662
rect 91 657 1471 658
rect 1477 657 1478 663
rect 202 636 208 637
rect 346 636 352 637
rect 202 632 203 636
rect 207 632 347 636
rect 351 632 352 636
rect 202 631 208 632
rect 346 631 352 632
rect 446 636 452 637
rect 530 636 536 637
rect 446 632 447 636
rect 451 632 531 636
rect 535 632 536 636
rect 446 631 452 632
rect 530 631 536 632
rect 96 617 97 623
rect 103 622 1483 623
rect 103 618 111 622
rect 115 618 191 622
rect 195 618 215 622
rect 219 618 239 622
rect 243 618 263 622
rect 267 618 271 622
rect 275 618 295 622
rect 299 618 319 622
rect 323 618 327 622
rect 331 618 343 622
rect 347 618 367 622
rect 371 618 391 622
rect 395 618 407 622
rect 411 618 415 622
rect 419 618 439 622
rect 443 618 455 622
rect 459 618 479 622
rect 483 618 503 622
rect 507 618 519 622
rect 523 618 551 622
rect 555 618 567 622
rect 571 618 607 622
rect 611 618 623 622
rect 627 618 663 622
rect 667 618 679 622
rect 683 618 719 622
rect 723 618 735 622
rect 739 618 767 622
rect 771 618 783 622
rect 787 618 815 622
rect 819 618 831 622
rect 835 618 863 622
rect 867 618 879 622
rect 883 618 903 622
rect 907 618 927 622
rect 931 618 935 622
rect 939 618 967 622
rect 971 618 975 622
rect 979 618 1007 622
rect 1011 618 1023 622
rect 1027 618 1047 622
rect 1051 618 1071 622
rect 1075 618 1087 622
rect 1091 618 1111 622
rect 1115 618 1127 622
rect 1131 618 1151 622
rect 1155 618 1159 622
rect 1163 618 1191 622
rect 1195 618 1223 622
rect 1227 618 1239 622
rect 1243 618 1263 622
rect 1267 618 1287 622
rect 1291 618 1303 622
rect 1307 618 1335 622
rect 1339 618 1343 622
rect 1347 618 1447 622
rect 1451 618 1483 622
rect 103 617 1483 618
rect 1489 617 1490 623
rect 84 577 85 583
rect 91 582 1471 583
rect 91 578 111 582
rect 115 578 263 582
rect 267 578 271 582
rect 275 578 287 582
rect 291 578 295 582
rect 299 578 311 582
rect 315 578 319 582
rect 323 578 335 582
rect 339 578 343 582
rect 347 578 359 582
rect 363 578 367 582
rect 371 578 383 582
rect 387 578 391 582
rect 395 578 407 582
rect 411 578 415 582
rect 419 578 431 582
rect 435 578 439 582
rect 443 578 463 582
rect 467 578 479 582
rect 483 578 503 582
rect 507 578 519 582
rect 523 578 551 582
rect 555 578 567 582
rect 571 578 607 582
rect 611 578 623 582
rect 627 578 663 582
rect 667 578 679 582
rect 683 578 719 582
rect 723 578 735 582
rect 739 578 775 582
rect 779 578 783 582
rect 787 578 831 582
rect 835 578 879 582
rect 883 578 887 582
rect 891 578 927 582
rect 931 578 943 582
rect 947 578 975 582
rect 979 578 1007 582
rect 1011 578 1023 582
rect 1027 578 1071 582
rect 1075 578 1111 582
rect 1115 578 1127 582
rect 1131 578 1151 582
rect 1155 578 1183 582
rect 1187 578 1191 582
rect 1195 578 1239 582
rect 1243 578 1247 582
rect 1251 578 1287 582
rect 1291 578 1311 582
rect 1315 578 1335 582
rect 1339 578 1375 582
rect 1379 578 1447 582
rect 1451 578 1471 582
rect 91 577 1471 578
rect 1477 577 1478 583
rect 96 537 97 543
rect 103 542 1483 543
rect 103 538 111 542
rect 115 538 223 542
rect 227 538 247 542
rect 251 538 263 542
rect 267 538 271 542
rect 275 538 287 542
rect 291 538 295 542
rect 299 538 311 542
rect 315 538 327 542
rect 331 538 335 542
rect 339 538 359 542
rect 363 538 383 542
rect 387 538 391 542
rect 395 538 407 542
rect 411 538 423 542
rect 427 538 431 542
rect 435 538 455 542
rect 459 538 463 542
rect 467 538 487 542
rect 491 538 503 542
rect 507 538 527 542
rect 531 538 551 542
rect 555 538 575 542
rect 579 538 607 542
rect 611 538 623 542
rect 627 538 663 542
rect 667 538 671 542
rect 675 538 711 542
rect 715 538 719 542
rect 723 538 759 542
rect 763 538 775 542
rect 779 538 807 542
rect 811 538 831 542
rect 835 538 855 542
rect 859 538 887 542
rect 891 538 911 542
rect 915 538 943 542
rect 947 538 967 542
rect 971 538 1007 542
rect 1011 538 1023 542
rect 1027 538 1071 542
rect 1075 538 1079 542
rect 1083 538 1127 542
rect 1131 538 1175 542
rect 1179 538 1183 542
rect 1187 538 1223 542
rect 1227 538 1247 542
rect 1251 538 1271 542
rect 1275 538 1311 542
rect 1315 538 1351 542
rect 1355 538 1375 542
rect 1379 538 1391 542
rect 1395 538 1415 542
rect 1419 538 1447 542
rect 1451 538 1483 542
rect 103 537 1483 538
rect 1489 537 1490 543
rect 84 497 85 503
rect 91 502 1471 503
rect 91 498 111 502
rect 115 498 135 502
rect 139 498 159 502
rect 163 498 183 502
rect 187 498 223 502
rect 227 498 247 502
rect 251 498 271 502
rect 275 498 295 502
rect 299 498 319 502
rect 323 498 327 502
rect 331 498 359 502
rect 363 498 375 502
rect 379 498 391 502
rect 395 498 423 502
rect 427 498 431 502
rect 435 498 455 502
rect 459 498 487 502
rect 491 498 527 502
rect 531 498 543 502
rect 547 498 575 502
rect 579 498 591 502
rect 595 498 623 502
rect 627 498 631 502
rect 635 498 663 502
rect 667 498 671 502
rect 675 498 687 502
rect 691 498 711 502
rect 715 498 719 502
rect 723 498 759 502
rect 763 498 799 502
rect 803 498 807 502
rect 811 498 847 502
rect 851 498 855 502
rect 859 498 903 502
rect 907 498 911 502
rect 915 498 951 502
rect 955 498 967 502
rect 971 498 999 502
rect 1003 498 1023 502
rect 1027 498 1047 502
rect 1051 498 1079 502
rect 1083 498 1095 502
rect 1099 498 1127 502
rect 1131 498 1143 502
rect 1147 498 1175 502
rect 1179 498 1199 502
rect 1203 498 1223 502
rect 1227 498 1255 502
rect 1259 498 1271 502
rect 1275 498 1311 502
rect 1315 498 1351 502
rect 1355 498 1375 502
rect 1379 498 1391 502
rect 1395 498 1415 502
rect 1419 498 1447 502
rect 1451 498 1471 502
rect 91 497 1471 498
rect 1477 497 1478 503
rect 96 457 97 463
rect 103 462 1483 463
rect 103 458 111 462
rect 115 458 135 462
rect 139 458 159 462
rect 163 458 183 462
rect 187 458 191 462
rect 195 458 223 462
rect 227 458 239 462
rect 243 458 271 462
rect 275 458 295 462
rect 299 458 319 462
rect 323 458 351 462
rect 355 458 375 462
rect 379 458 415 462
rect 419 458 431 462
rect 435 458 479 462
rect 483 458 487 462
rect 491 458 543 462
rect 547 458 591 462
rect 595 458 607 462
rect 611 458 631 462
rect 635 458 663 462
rect 667 458 671 462
rect 675 458 687 462
rect 691 458 719 462
rect 723 458 735 462
rect 739 458 759 462
rect 763 458 791 462
rect 795 458 799 462
rect 803 458 839 462
rect 843 458 847 462
rect 851 458 879 462
rect 883 458 903 462
rect 907 458 911 462
rect 915 458 943 462
rect 947 458 951 462
rect 955 458 967 462
rect 971 458 999 462
rect 1003 458 1031 462
rect 1035 458 1047 462
rect 1051 458 1071 462
rect 1075 458 1095 462
rect 1099 458 1119 462
rect 1123 458 1143 462
rect 1147 458 1175 462
rect 1179 458 1199 462
rect 1203 458 1239 462
rect 1243 458 1255 462
rect 1259 458 1303 462
rect 1307 458 1311 462
rect 1315 458 1367 462
rect 1371 458 1375 462
rect 1379 458 1415 462
rect 1419 458 1447 462
rect 1451 458 1483 462
rect 103 457 1483 458
rect 1489 457 1490 463
rect 84 417 85 423
rect 91 422 1471 423
rect 91 418 111 422
rect 115 418 135 422
rect 139 418 159 422
rect 163 418 183 422
rect 187 418 191 422
rect 195 418 215 422
rect 219 418 239 422
rect 243 418 271 422
rect 275 418 295 422
rect 299 418 327 422
rect 331 418 351 422
rect 355 418 391 422
rect 395 418 415 422
rect 419 418 447 422
rect 451 418 479 422
rect 483 418 503 422
rect 507 418 543 422
rect 547 418 551 422
rect 555 418 599 422
rect 603 418 607 422
rect 611 418 647 422
rect 651 418 671 422
rect 675 418 703 422
rect 707 418 735 422
rect 739 418 767 422
rect 771 418 791 422
rect 795 418 831 422
rect 835 418 839 422
rect 843 418 879 422
rect 883 418 903 422
rect 907 418 911 422
rect 915 418 943 422
rect 947 418 967 422
rect 971 418 975 422
rect 979 418 999 422
rect 1003 418 1031 422
rect 1035 418 1039 422
rect 1043 418 1071 422
rect 1075 418 1103 422
rect 1107 418 1119 422
rect 1123 418 1159 422
rect 1163 418 1175 422
rect 1179 418 1207 422
rect 1211 418 1239 422
rect 1243 418 1247 422
rect 1251 418 1279 422
rect 1283 418 1303 422
rect 1307 418 1319 422
rect 1323 418 1359 422
rect 1363 418 1367 422
rect 1371 418 1391 422
rect 1395 418 1415 422
rect 1419 418 1447 422
rect 1451 418 1471 422
rect 91 417 1471 418
rect 1477 417 1478 423
rect 96 373 97 379
rect 103 378 1483 379
rect 103 374 111 378
rect 115 374 135 378
rect 139 374 159 378
rect 163 374 183 378
rect 187 374 207 378
rect 211 374 215 378
rect 219 374 231 378
rect 235 374 255 378
rect 259 374 271 378
rect 275 374 295 378
rect 299 374 327 378
rect 331 374 335 378
rect 339 374 375 378
rect 379 374 391 378
rect 395 374 415 378
rect 419 374 447 378
rect 451 374 455 378
rect 459 374 495 378
rect 499 374 503 378
rect 507 374 535 378
rect 539 374 551 378
rect 555 374 575 378
rect 579 374 599 378
rect 603 374 615 378
rect 619 374 647 378
rect 651 374 655 378
rect 659 374 687 378
rect 691 374 703 378
rect 707 374 727 378
rect 731 374 767 378
rect 771 374 775 378
rect 779 374 831 378
rect 835 374 887 378
rect 891 374 903 378
rect 907 374 951 378
rect 955 374 975 378
rect 979 374 1015 378
rect 1019 374 1039 378
rect 1043 374 1079 378
rect 1083 374 1103 378
rect 1107 374 1135 378
rect 1139 374 1159 378
rect 1163 374 1183 378
rect 1187 374 1207 378
rect 1211 374 1231 378
rect 1235 374 1247 378
rect 1251 374 1271 378
rect 1275 374 1279 378
rect 1283 374 1311 378
rect 1315 374 1319 378
rect 1323 374 1351 378
rect 1355 374 1359 378
rect 1363 374 1391 378
rect 1395 374 1415 378
rect 1419 374 1447 378
rect 1451 374 1483 378
rect 103 373 1483 374
rect 1489 373 1490 379
rect 84 333 85 339
rect 91 338 1471 339
rect 91 334 111 338
rect 115 334 135 338
rect 139 334 159 338
rect 163 334 175 338
rect 179 334 183 338
rect 187 334 199 338
rect 203 334 207 338
rect 211 334 223 338
rect 227 334 231 338
rect 235 334 247 338
rect 251 334 255 338
rect 259 334 279 338
rect 283 334 295 338
rect 299 334 319 338
rect 323 334 335 338
rect 339 334 359 338
rect 363 334 375 338
rect 379 334 399 338
rect 403 334 415 338
rect 419 334 439 338
rect 443 334 455 338
rect 459 334 479 338
rect 483 334 495 338
rect 499 334 527 338
rect 531 334 535 338
rect 539 334 575 338
rect 579 334 583 338
rect 587 334 615 338
rect 619 334 639 338
rect 643 334 655 338
rect 659 334 687 338
rect 691 334 727 338
rect 731 334 735 338
rect 739 334 775 338
rect 779 334 791 338
rect 795 334 831 338
rect 835 334 847 338
rect 851 334 887 338
rect 891 334 895 338
rect 899 334 943 338
rect 947 334 951 338
rect 955 334 991 338
rect 995 334 1015 338
rect 1019 334 1039 338
rect 1043 334 1079 338
rect 1083 334 1087 338
rect 1091 334 1135 338
rect 1139 334 1183 338
rect 1187 334 1231 338
rect 1235 334 1271 338
rect 1275 334 1279 338
rect 1283 334 1311 338
rect 1315 334 1327 338
rect 1331 334 1351 338
rect 1355 334 1383 338
rect 1387 334 1391 338
rect 1395 334 1415 338
rect 1419 334 1447 338
rect 1451 334 1471 338
rect 91 333 1471 334
rect 1477 333 1478 339
rect 186 316 192 317
rect 346 316 352 317
rect 186 312 187 316
rect 191 312 347 316
rect 351 312 352 316
rect 186 311 192 312
rect 346 311 352 312
rect 96 293 97 299
rect 103 298 1483 299
rect 103 294 111 298
rect 115 294 175 298
rect 179 294 199 298
rect 203 294 223 298
rect 227 294 247 298
rect 251 294 271 298
rect 275 294 279 298
rect 283 294 295 298
rect 299 294 319 298
rect 323 294 343 298
rect 347 294 359 298
rect 363 294 367 298
rect 371 294 399 298
rect 403 294 431 298
rect 435 294 439 298
rect 443 294 471 298
rect 475 294 479 298
rect 483 294 511 298
rect 515 294 527 298
rect 531 294 559 298
rect 563 294 583 298
rect 587 294 615 298
rect 619 294 639 298
rect 643 294 663 298
rect 667 294 687 298
rect 691 294 711 298
rect 715 294 735 298
rect 739 294 759 298
rect 763 294 791 298
rect 795 294 807 298
rect 811 294 847 298
rect 851 294 879 298
rect 883 294 895 298
rect 899 294 903 298
rect 907 294 927 298
rect 931 294 943 298
rect 947 294 951 298
rect 955 294 975 298
rect 979 294 991 298
rect 995 294 999 298
rect 1003 294 1023 298
rect 1027 294 1039 298
rect 1043 294 1047 298
rect 1051 294 1071 298
rect 1075 294 1087 298
rect 1091 294 1095 298
rect 1099 294 1127 298
rect 1131 294 1135 298
rect 1139 294 1159 298
rect 1163 294 1183 298
rect 1187 294 1199 298
rect 1203 294 1231 298
rect 1235 294 1247 298
rect 1251 294 1279 298
rect 1283 294 1303 298
rect 1307 294 1327 298
rect 1331 294 1367 298
rect 1371 294 1383 298
rect 1387 294 1415 298
rect 1419 294 1447 298
rect 1451 294 1483 298
rect 103 293 1483 294
rect 1489 293 1490 299
rect 278 268 284 269
rect 410 268 416 269
rect 278 264 279 268
rect 283 264 411 268
rect 415 264 416 268
rect 278 263 284 264
rect 410 263 416 264
rect 84 253 85 259
rect 91 258 1471 259
rect 91 254 111 258
rect 115 254 247 258
rect 251 254 263 258
rect 267 254 271 258
rect 275 254 287 258
rect 291 254 295 258
rect 299 254 311 258
rect 315 254 319 258
rect 323 254 335 258
rect 339 254 343 258
rect 347 254 359 258
rect 363 254 367 258
rect 371 254 383 258
rect 387 254 399 258
rect 403 254 407 258
rect 411 254 431 258
rect 435 254 463 258
rect 467 254 471 258
rect 475 254 503 258
rect 507 254 511 258
rect 515 254 543 258
rect 547 254 559 258
rect 563 254 583 258
rect 587 254 615 258
rect 619 254 623 258
rect 627 254 663 258
rect 667 254 679 258
rect 683 254 711 258
rect 715 254 743 258
rect 747 254 759 258
rect 763 254 807 258
rect 811 254 847 258
rect 851 254 879 258
rect 883 254 903 258
rect 907 254 927 258
rect 931 254 951 258
rect 955 254 959 258
rect 963 254 975 258
rect 979 254 999 258
rect 1003 254 1023 258
rect 1027 254 1039 258
rect 1043 254 1047 258
rect 1051 254 1071 258
rect 1075 254 1095 258
rect 1099 254 1119 258
rect 1123 254 1127 258
rect 1131 254 1159 258
rect 1163 254 1199 258
rect 1203 254 1247 258
rect 1251 254 1279 258
rect 1283 254 1303 258
rect 1307 254 1359 258
rect 1363 254 1367 258
rect 1371 254 1415 258
rect 1419 254 1447 258
rect 1451 254 1471 258
rect 91 253 1471 254
rect 1477 253 1478 259
rect 96 213 97 219
rect 103 218 1483 219
rect 103 214 111 218
rect 115 214 239 218
rect 243 214 263 218
rect 267 214 287 218
rect 291 214 311 218
rect 315 214 335 218
rect 339 214 359 218
rect 363 214 383 218
rect 387 214 407 218
rect 411 214 431 218
rect 435 214 463 218
rect 467 214 503 218
rect 507 214 511 218
rect 515 214 543 218
rect 547 214 559 218
rect 563 214 583 218
rect 587 214 615 218
rect 619 214 623 218
rect 627 214 671 218
rect 675 214 679 218
rect 683 214 719 218
rect 723 214 743 218
rect 747 214 767 218
rect 771 214 807 218
rect 811 214 815 218
rect 819 214 863 218
rect 867 214 879 218
rect 883 214 919 218
rect 923 214 959 218
rect 963 214 975 218
rect 979 214 1031 218
rect 1035 214 1039 218
rect 1043 214 1087 218
rect 1091 214 1119 218
rect 1123 214 1135 218
rect 1139 214 1183 218
rect 1187 214 1199 218
rect 1203 214 1231 218
rect 1235 214 1279 218
rect 1283 214 1327 218
rect 1331 214 1359 218
rect 1363 214 1383 218
rect 1387 214 1415 218
rect 1419 214 1447 218
rect 1451 214 1483 218
rect 103 213 1483 214
rect 1489 213 1490 219
rect 418 204 424 205
rect 590 204 596 205
rect 418 200 419 204
rect 423 200 591 204
rect 595 200 596 204
rect 418 199 424 200
rect 590 199 596 200
rect 84 173 85 179
rect 91 178 1471 179
rect 91 174 111 178
rect 115 174 183 178
rect 187 174 207 178
rect 211 174 239 178
rect 243 174 263 178
rect 267 174 279 178
rect 283 174 287 178
rect 291 174 311 178
rect 315 174 327 178
rect 331 174 335 178
rect 339 174 359 178
rect 363 174 375 178
rect 379 174 383 178
rect 387 174 407 178
rect 411 174 423 178
rect 427 174 431 178
rect 435 174 463 178
rect 467 174 471 178
rect 475 174 511 178
rect 515 174 527 178
rect 531 174 559 178
rect 563 174 591 178
rect 595 174 615 178
rect 619 174 655 178
rect 659 174 671 178
rect 675 174 711 178
rect 715 174 719 178
rect 723 174 767 178
rect 771 174 815 178
rect 819 174 823 178
rect 827 174 863 178
rect 867 174 871 178
rect 875 174 919 178
rect 923 174 975 178
rect 979 174 1031 178
rect 1035 174 1079 178
rect 1083 174 1087 178
rect 1091 174 1127 178
rect 1131 174 1135 178
rect 1139 174 1175 178
rect 1179 174 1183 178
rect 1187 174 1223 178
rect 1227 174 1231 178
rect 1235 174 1263 178
rect 1267 174 1279 178
rect 1283 174 1295 178
rect 1299 174 1327 178
rect 1331 174 1359 178
rect 1363 174 1383 178
rect 1387 174 1391 178
rect 1395 174 1415 178
rect 1419 174 1447 178
rect 1451 174 1471 178
rect 91 173 1471 174
rect 1477 173 1478 179
rect 96 121 97 127
rect 103 126 1483 127
rect 103 122 111 126
rect 115 122 135 126
rect 139 122 159 126
rect 163 122 183 126
rect 187 122 207 126
rect 211 122 231 126
rect 235 122 239 126
rect 243 122 255 126
rect 259 122 279 126
rect 283 122 303 126
rect 307 122 327 126
rect 331 122 351 126
rect 355 122 375 126
rect 379 122 399 126
rect 403 122 423 126
rect 427 122 431 126
rect 435 122 463 126
rect 467 122 471 126
rect 475 122 487 126
rect 491 122 511 126
rect 515 122 527 126
rect 531 122 535 126
rect 539 122 559 126
rect 563 122 583 126
rect 587 122 591 126
rect 595 122 607 126
rect 611 122 631 126
rect 635 122 655 126
rect 659 122 679 126
rect 683 122 703 126
rect 707 122 711 126
rect 715 122 727 126
rect 731 122 751 126
rect 755 122 767 126
rect 771 122 775 126
rect 779 122 799 126
rect 803 122 823 126
rect 827 122 855 126
rect 859 122 871 126
rect 875 122 887 126
rect 891 122 919 126
rect 923 122 951 126
rect 955 122 975 126
rect 979 122 983 126
rect 987 122 1015 126
rect 1019 122 1031 126
rect 1035 122 1047 126
rect 1051 122 1071 126
rect 1075 122 1079 126
rect 1083 122 1095 126
rect 1099 122 1119 126
rect 1123 122 1127 126
rect 1131 122 1143 126
rect 1147 122 1175 126
rect 1179 122 1207 126
rect 1211 122 1223 126
rect 1227 122 1239 126
rect 1243 122 1263 126
rect 1267 122 1271 126
rect 1275 122 1295 126
rect 1299 122 1303 126
rect 1307 122 1327 126
rect 1331 122 1335 126
rect 1339 122 1359 126
rect 1363 122 1367 126
rect 1371 122 1391 126
rect 1395 122 1415 126
rect 1419 122 1447 126
rect 1451 122 1483 126
rect 103 121 1483 122
rect 1489 121 1490 127
rect 84 81 85 87
rect 91 86 1471 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 159 86
rect 163 82 183 86
rect 187 82 207 86
rect 211 82 231 86
rect 235 82 255 86
rect 259 82 279 86
rect 283 82 303 86
rect 307 82 327 86
rect 331 82 351 86
rect 355 82 375 86
rect 379 82 399 86
rect 403 82 431 86
rect 435 82 463 86
rect 467 82 487 86
rect 491 82 511 86
rect 515 82 535 86
rect 539 82 559 86
rect 563 82 583 86
rect 587 82 607 86
rect 611 82 631 86
rect 635 82 655 86
rect 659 82 679 86
rect 683 82 703 86
rect 707 82 727 86
rect 731 82 751 86
rect 755 82 775 86
rect 779 82 799 86
rect 803 82 823 86
rect 827 82 855 86
rect 859 82 887 86
rect 891 82 919 86
rect 923 82 951 86
rect 955 82 983 86
rect 987 82 1015 86
rect 1019 82 1047 86
rect 1051 82 1071 86
rect 1075 82 1095 86
rect 1099 82 1119 86
rect 1123 82 1143 86
rect 1147 82 1175 86
rect 1179 82 1207 86
rect 1211 82 1239 86
rect 1243 82 1271 86
rect 1275 82 1303 86
rect 1307 82 1335 86
rect 1339 82 1367 86
rect 1371 82 1391 86
rect 1395 82 1415 86
rect 1419 82 1447 86
rect 1451 82 1471 86
rect 91 81 1471 82
rect 1477 81 1478 87
<< m5c >>
rect 97 1505 103 1511
rect 1483 1505 1489 1511
rect 85 1465 91 1471
rect 1471 1465 1477 1471
rect 97 1425 103 1431
rect 1483 1425 1489 1431
rect 85 1385 91 1391
rect 1471 1385 1477 1391
rect 97 1345 103 1351
rect 1483 1345 1489 1351
rect 85 1305 91 1311
rect 1471 1305 1477 1311
rect 97 1265 103 1271
rect 1483 1265 1489 1271
rect 85 1225 91 1231
rect 1471 1225 1477 1231
rect 97 1185 103 1191
rect 1483 1185 1489 1191
rect 85 1145 91 1151
rect 1471 1145 1477 1151
rect 97 1101 103 1107
rect 1483 1101 1489 1107
rect 85 1061 91 1067
rect 1471 1061 1477 1067
rect 97 1021 103 1027
rect 1483 1021 1489 1027
rect 85 981 91 987
rect 1471 981 1477 987
rect 97 941 103 947
rect 1483 941 1489 947
rect 85 901 91 907
rect 1471 901 1477 907
rect 97 861 103 867
rect 1483 861 1489 867
rect 85 821 91 827
rect 1471 821 1477 827
rect 97 781 103 787
rect 1483 781 1489 787
rect 85 737 91 743
rect 1471 737 1477 743
rect 97 697 103 703
rect 1483 697 1489 703
rect 85 657 91 663
rect 1471 657 1477 663
rect 97 617 103 623
rect 1483 617 1489 623
rect 85 577 91 583
rect 1471 577 1477 583
rect 97 537 103 543
rect 1483 537 1489 543
rect 85 497 91 503
rect 1471 497 1477 503
rect 97 457 103 463
rect 1483 457 1489 463
rect 85 417 91 423
rect 1471 417 1477 423
rect 97 373 103 379
rect 1483 373 1489 379
rect 85 333 91 339
rect 1471 333 1477 339
rect 97 293 103 299
rect 1483 293 1489 299
rect 85 253 91 259
rect 1471 253 1477 259
rect 97 213 103 219
rect 1483 213 1489 219
rect 85 173 91 179
rect 1471 173 1477 179
rect 97 121 103 127
rect 1483 121 1489 127
rect 85 81 91 87
rect 1471 81 1477 87
<< m5 >>
rect 84 1471 92 1512
rect 84 1465 85 1471
rect 91 1465 92 1471
rect 84 1391 92 1465
rect 84 1385 85 1391
rect 91 1385 92 1391
rect 84 1311 92 1385
rect 84 1305 85 1311
rect 91 1305 92 1311
rect 84 1231 92 1305
rect 84 1225 85 1231
rect 91 1225 92 1231
rect 84 1151 92 1225
rect 84 1145 85 1151
rect 91 1145 92 1151
rect 84 1067 92 1145
rect 84 1061 85 1067
rect 91 1061 92 1067
rect 84 987 92 1061
rect 84 981 85 987
rect 91 981 92 987
rect 84 907 92 981
rect 84 901 85 907
rect 91 901 92 907
rect 84 827 92 901
rect 84 821 85 827
rect 91 821 92 827
rect 84 743 92 821
rect 84 737 85 743
rect 91 737 92 743
rect 84 663 92 737
rect 84 657 85 663
rect 91 657 92 663
rect 84 583 92 657
rect 84 577 85 583
rect 91 577 92 583
rect 84 503 92 577
rect 84 497 85 503
rect 91 497 92 503
rect 84 423 92 497
rect 84 417 85 423
rect 91 417 92 423
rect 84 339 92 417
rect 84 333 85 339
rect 91 333 92 339
rect 84 259 92 333
rect 84 253 85 259
rect 91 253 92 259
rect 84 179 92 253
rect 84 173 85 179
rect 91 173 92 179
rect 84 87 92 173
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 1511 104 1512
rect 96 1505 97 1511
rect 103 1505 104 1511
rect 96 1431 104 1505
rect 96 1425 97 1431
rect 103 1425 104 1431
rect 96 1351 104 1425
rect 96 1345 97 1351
rect 103 1345 104 1351
rect 96 1271 104 1345
rect 96 1265 97 1271
rect 103 1265 104 1271
rect 96 1191 104 1265
rect 96 1185 97 1191
rect 103 1185 104 1191
rect 96 1107 104 1185
rect 96 1101 97 1107
rect 103 1101 104 1107
rect 96 1027 104 1101
rect 96 1021 97 1027
rect 103 1021 104 1027
rect 96 947 104 1021
rect 96 941 97 947
rect 103 941 104 947
rect 96 867 104 941
rect 96 861 97 867
rect 103 861 104 867
rect 96 787 104 861
rect 96 781 97 787
rect 103 781 104 787
rect 96 703 104 781
rect 96 697 97 703
rect 103 697 104 703
rect 96 623 104 697
rect 96 617 97 623
rect 103 617 104 623
rect 96 543 104 617
rect 96 537 97 543
rect 103 537 104 543
rect 96 463 104 537
rect 96 457 97 463
rect 103 457 104 463
rect 96 379 104 457
rect 96 373 97 379
rect 103 373 104 379
rect 96 299 104 373
rect 96 293 97 299
rect 103 293 104 299
rect 96 219 104 293
rect 96 213 97 219
rect 103 213 104 219
rect 96 127 104 213
rect 96 121 97 127
rect 103 121 104 127
rect 96 72 104 121
rect 1470 1471 1478 1512
rect 1470 1465 1471 1471
rect 1477 1465 1478 1471
rect 1470 1391 1478 1465
rect 1470 1385 1471 1391
rect 1477 1385 1478 1391
rect 1470 1311 1478 1385
rect 1470 1305 1471 1311
rect 1477 1305 1478 1311
rect 1470 1231 1478 1305
rect 1470 1225 1471 1231
rect 1477 1225 1478 1231
rect 1470 1151 1478 1225
rect 1470 1145 1471 1151
rect 1477 1145 1478 1151
rect 1470 1067 1478 1145
rect 1470 1061 1471 1067
rect 1477 1061 1478 1067
rect 1470 987 1478 1061
rect 1470 981 1471 987
rect 1477 981 1478 987
rect 1470 907 1478 981
rect 1470 901 1471 907
rect 1477 901 1478 907
rect 1470 827 1478 901
rect 1470 821 1471 827
rect 1477 821 1478 827
rect 1470 743 1478 821
rect 1470 737 1471 743
rect 1477 737 1478 743
rect 1470 663 1478 737
rect 1470 657 1471 663
rect 1477 657 1478 663
rect 1470 583 1478 657
rect 1470 577 1471 583
rect 1477 577 1478 583
rect 1470 503 1478 577
rect 1470 497 1471 503
rect 1477 497 1478 503
rect 1470 423 1478 497
rect 1470 417 1471 423
rect 1477 417 1478 423
rect 1470 339 1478 417
rect 1470 333 1471 339
rect 1477 333 1478 339
rect 1470 259 1478 333
rect 1470 253 1471 259
rect 1477 253 1478 259
rect 1470 179 1478 253
rect 1470 173 1471 179
rect 1477 173 1478 179
rect 1470 87 1478 173
rect 1470 81 1471 87
rect 1477 81 1478 87
rect 1470 72 1478 81
rect 1482 1511 1490 1512
rect 1482 1505 1483 1511
rect 1489 1505 1490 1511
rect 1482 1431 1490 1505
rect 1482 1425 1483 1431
rect 1489 1425 1490 1431
rect 1482 1351 1490 1425
rect 1482 1345 1483 1351
rect 1489 1345 1490 1351
rect 1482 1271 1490 1345
rect 1482 1265 1483 1271
rect 1489 1265 1490 1271
rect 1482 1191 1490 1265
rect 1482 1185 1483 1191
rect 1489 1185 1490 1191
rect 1482 1107 1490 1185
rect 1482 1101 1483 1107
rect 1489 1101 1490 1107
rect 1482 1027 1490 1101
rect 1482 1021 1483 1027
rect 1489 1021 1490 1027
rect 1482 947 1490 1021
rect 1482 941 1483 947
rect 1489 941 1490 947
rect 1482 867 1490 941
rect 1482 861 1483 867
rect 1489 861 1490 867
rect 1482 787 1490 861
rect 1482 781 1483 787
rect 1489 781 1490 787
rect 1482 703 1490 781
rect 1482 697 1483 703
rect 1489 697 1490 703
rect 1482 623 1490 697
rect 1482 617 1483 623
rect 1489 617 1490 623
rect 1482 543 1490 617
rect 1482 537 1483 543
rect 1489 537 1490 543
rect 1482 463 1490 537
rect 1482 457 1483 463
rect 1489 457 1490 463
rect 1482 379 1490 457
rect 1482 373 1483 379
rect 1489 373 1490 379
rect 1482 299 1490 373
rect 1482 293 1483 299
rect 1489 293 1490 299
rect 1482 219 1490 293
rect 1482 213 1483 219
rect 1489 213 1490 219
rect 1482 127 1490 213
rect 1482 121 1483 127
rect 1489 121 1490 127
rect 1482 72 1490 121
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730589202
transform 1 0 104 0 1 88
box 8 4 12 24
use welltap_svt  __well_tap__0
timestamp 1730589202
transform 1 0 104 0 1 88
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0INVX1  inv_5999_6
timestamp 1730589202
transform 1 0 128 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5998_6
timestamp 1730589202
transform 1 0 152 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5998_6
timestamp 1730589202
transform 1 0 152 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5999_6
timestamp 1730589202
transform 1 0 128 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5997_6
timestamp 1730589202
transform 1 0 176 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5997_6
timestamp 1730589202
transform 1 0 176 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5996_6
timestamp 1730589202
transform 1 0 200 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5995_6
timestamp 1730589202
transform 1 0 224 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5995_6
timestamp 1730589202
transform 1 0 224 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5996_6
timestamp 1730589202
transform 1 0 200 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5994_6
timestamp 1730589202
transform 1 0 248 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5993_6
timestamp 1730589202
transform 1 0 272 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5993_6
timestamp 1730589202
transform 1 0 272 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5994_6
timestamp 1730589202
transform 1 0 248 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5992_6
timestamp 1730589202
transform 1 0 296 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5991_6
timestamp 1730589202
transform 1 0 320 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5991_6
timestamp 1730589202
transform 1 0 320 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5992_6
timestamp 1730589202
transform 1 0 296 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5990_6
timestamp 1730589202
transform 1 0 344 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5990_6
timestamp 1730589202
transform 1 0 344 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5989_6
timestamp 1730589202
transform 1 0 368 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5988_6
timestamp 1730589202
transform 1 0 392 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5988_6
timestamp 1730589202
transform 1 0 392 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5989_6
timestamp 1730589202
transform 1 0 368 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5908_6
timestamp 1730589202
transform 1 0 424 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5908_6
timestamp 1730589202
transform 1 0 424 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5910_6
timestamp 1730589202
transform 1 0 480 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5909_6
timestamp 1730589202
transform 1 0 456 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5909_6
timestamp 1730589202
transform 1 0 456 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5910_6
timestamp 1730589202
transform 1 0 480 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5912_6
timestamp 1730589202
transform 1 0 528 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5911_6
timestamp 1730589202
transform 1 0 504 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5911_6
timestamp 1730589202
transform 1 0 504 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5912_6
timestamp 1730589202
transform 1 0 528 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5913_6
timestamp 1730589202
transform 1 0 552 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5913_6
timestamp 1730589202
transform 1 0 552 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5915_6
timestamp 1730589202
transform 1 0 600 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5914_6
timestamp 1730589202
transform 1 0 576 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5914_6
timestamp 1730589202
transform 1 0 576 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5915_6
timestamp 1730589202
transform 1 0 600 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5917_6
timestamp 1730589202
transform 1 0 648 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5916_6
timestamp 1730589202
transform 1 0 624 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5916_6
timestamp 1730589202
transform 1 0 624 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5917_6
timestamp 1730589202
transform 1 0 648 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5919_6
timestamp 1730589202
transform 1 0 696 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5918_6
timestamp 1730589202
transform 1 0 672 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5918_6
timestamp 1730589202
transform 1 0 672 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5919_6
timestamp 1730589202
transform 1 0 696 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5920_6
timestamp 1730589202
transform 1 0 720 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5920_6
timestamp 1730589202
transform 1 0 720 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5922_6
timestamp 1730589202
transform 1 0 768 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5921_6
timestamp 1730589202
transform 1 0 744 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5921_6
timestamp 1730589202
transform 1 0 744 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5922_6
timestamp 1730589202
transform 1 0 768 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5924_6
timestamp 1730589202
transform 1 0 816 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5923_6
timestamp 1730589202
transform 1 0 792 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5923_6
timestamp 1730589202
transform 1 0 792 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5924_6
timestamp 1730589202
transform 1 0 816 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5925_6
timestamp 1730589202
transform 1 0 848 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5925_6
timestamp 1730589202
transform 1 0 848 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5926_6
timestamp 1730589202
transform 1 0 880 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5926_6
timestamp 1730589202
transform 1 0 880 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5928_6
timestamp 1730589202
transform 1 0 944 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5927_6
timestamp 1730589202
transform 1 0 912 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5927_6
timestamp 1730589202
transform 1 0 912 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5928_6
timestamp 1730589202
transform 1 0 944 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5929_6
timestamp 1730589202
transform 1 0 976 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5929_6
timestamp 1730589202
transform 1 0 976 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5930_6
timestamp 1730589202
transform 1 0 1008 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5930_6
timestamp 1730589202
transform 1 0 1008 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5282_6
timestamp 1730589202
transform 1 0 1040 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5281_6
timestamp 1730589202
transform 1 0 1064 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5281_6
timestamp 1730589202
transform 1 0 1064 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5282_6
timestamp 1730589202
transform 1 0 1040 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5280_6
timestamp 1730589202
transform 1 0 1088 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5279_6
timestamp 1730589202
transform 1 0 1112 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5279_6
timestamp 1730589202
transform 1 0 1112 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5280_6
timestamp 1730589202
transform 1 0 1088 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5278_6
timestamp 1730589202
transform 1 0 1136 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5278_6
timestamp 1730589202
transform 1 0 1136 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5277_6
timestamp 1730589202
transform 1 0 1168 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5276_6
timestamp 1730589202
transform 1 0 1200 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5276_6
timestamp 1730589202
transform 1 0 1200 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5277_6
timestamp 1730589202
transform 1 0 1168 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5275_6
timestamp 1730589202
transform 1 0 1232 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5275_6
timestamp 1730589202
transform 1 0 1232 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5274_6
timestamp 1730589202
transform 1 0 1264 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5274_6
timestamp 1730589202
transform 1 0 1264 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5273_6
timestamp 1730589202
transform 1 0 1296 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5272_6
timestamp 1730589202
transform 1 0 1328 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5272_6
timestamp 1730589202
transform 1 0 1328 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5273_6
timestamp 1730589202
transform 1 0 1296 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5261_6
timestamp 1730589202
transform 1 0 1360 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5261_6
timestamp 1730589202
transform 1 0 1360 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5260_6
timestamp 1730589202
transform 1 0 1384 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5259_6
timestamp 1730589202
transform 1 0 1408 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5259_6
timestamp 1730589202
transform 1 0 1408 0 1 84
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5260_6
timestamp 1730589202
transform 1 0 1384 0 1 84
box 8 4 20 35
use welltap_svt  __well_tap__1
timestamp 1730589202
transform 1 0 1440 0 1 88
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730589202
transform 1 0 1440 0 1 88
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730589202
transform 1 0 104 0 -1 172
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730589202
transform 1 0 104 0 -1 172
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5987_6
timestamp 1730589202
transform 1 0 176 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5987_6
timestamp 1730589202
transform 1 0 176 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5986_6
timestamp 1730589202
transform 1 0 200 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5985_6
timestamp 1730589202
transform 1 0 232 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5985_6
timestamp 1730589202
transform 1 0 232 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5986_6
timestamp 1730589202
transform 1 0 200 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5984_6
timestamp 1730589202
transform 1 0 272 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5984_6
timestamp 1730589202
transform 1 0 272 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5983_6
timestamp 1730589202
transform 1 0 320 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5983_6
timestamp 1730589202
transform 1 0 320 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5982_6
timestamp 1730589202
transform 1 0 368 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5982_6
timestamp 1730589202
transform 1 0 368 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5902_6
timestamp 1730589202
transform 1 0 416 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5902_6
timestamp 1730589202
transform 1 0 416 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5903_6
timestamp 1730589202
transform 1 0 464 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5903_6
timestamp 1730589202
transform 1 0 464 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5904_6
timestamp 1730589202
transform 1 0 520 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5904_6
timestamp 1730589202
transform 1 0 520 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5905_6
timestamp 1730589202
transform 1 0 584 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5905_6
timestamp 1730589202
transform 1 0 584 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5906_6
timestamp 1730589202
transform 1 0 648 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5906_6
timestamp 1730589202
transform 1 0 648 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5907_6
timestamp 1730589202
transform 1 0 704 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5907_6
timestamp 1730589202
transform 1 0 704 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5931_6
timestamp 1730589202
transform 1 0 760 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5931_6
timestamp 1730589202
transform 1 0 760 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5932_6
timestamp 1730589202
transform 1 0 816 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5932_6
timestamp 1730589202
transform 1 0 816 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5933_6
timestamp 1730589202
transform 1 0 864 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5933_6
timestamp 1730589202
transform 1 0 864 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5934_6
timestamp 1730589202
transform 1 0 912 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5934_6
timestamp 1730589202
transform 1 0 912 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5935_6
timestamp 1730589202
transform 1 0 968 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5935_6
timestamp 1730589202
transform 1 0 968 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5936_6
timestamp 1730589202
transform 1 0 1024 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5936_6
timestamp 1730589202
transform 1 0 1024 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5937_6
timestamp 1730589202
transform 1 0 1072 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5937_6
timestamp 1730589202
transform 1 0 1072 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5283_6
timestamp 1730589202
transform 1 0 1120 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5283_6
timestamp 1730589202
transform 1 0 1120 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5271_6
timestamp 1730589202
transform 1 0 1168 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5271_6
timestamp 1730589202
transform 1 0 1168 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5270_6
timestamp 1730589202
transform 1 0 1216 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5270_6
timestamp 1730589202
transform 1 0 1216 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5269_6
timestamp 1730589202
transform 1 0 1256 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5268_6
timestamp 1730589202
transform 1 0 1288 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5268_6
timestamp 1730589202
transform 1 0 1288 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5269_6
timestamp 1730589202
transform 1 0 1256 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5262_6
timestamp 1730589202
transform 1 0 1320 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5262_6
timestamp 1730589202
transform 1 0 1320 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5263_6
timestamp 1730589202
transform 1 0 1352 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5263_6
timestamp 1730589202
transform 1 0 1352 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5258_6
timestamp 1730589202
transform 1 0 1384 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5257_6
timestamp 1730589202
transform 1 0 1408 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5257_6
timestamp 1730589202
transform 1 0 1408 0 -1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5258_6
timestamp 1730589202
transform 1 0 1384 0 -1 176
box 8 4 20 35
use welltap_svt  __well_tap__3
timestamp 1730589202
transform 1 0 1440 0 -1 172
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730589202
transform 1 0 1440 0 -1 172
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730589202
transform 1 0 104 0 1 180
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730589202
transform 1 0 104 0 1 180
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5981_6
timestamp 1730589202
transform 1 0 232 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5981_6
timestamp 1730589202
transform 1 0 232 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5980_6
timestamp 1730589202
transform 1 0 256 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5979_6
timestamp 1730589202
transform 1 0 280 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5979_6
timestamp 1730589202
transform 1 0 280 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5980_6
timestamp 1730589202
transform 1 0 256 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5978_6
timestamp 1730589202
transform 1 0 304 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5978_6
timestamp 1730589202
transform 1 0 304 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5977_6
timestamp 1730589202
transform 1 0 328 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5976_6
timestamp 1730589202
transform 1 0 352 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5976_6
timestamp 1730589202
transform 1 0 352 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5977_6
timestamp 1730589202
transform 1 0 328 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5975_6
timestamp 1730589202
transform 1 0 376 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5895_6
timestamp 1730589202
transform 1 0 400 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5895_6
timestamp 1730589202
transform 1 0 400 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5975_6
timestamp 1730589202
transform 1 0 376 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5896_6
timestamp 1730589202
transform 1 0 424 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5896_6
timestamp 1730589202
transform 1 0 424 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5897_6
timestamp 1730589202
transform 1 0 456 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5897_6
timestamp 1730589202
transform 1 0 456 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5898_6
timestamp 1730589202
transform 1 0 504 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5898_6
timestamp 1730589202
transform 1 0 504 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5899_6
timestamp 1730589202
transform 1 0 552 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5899_6
timestamp 1730589202
transform 1 0 552 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5900_6
timestamp 1730589202
transform 1 0 608 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5900_6
timestamp 1730589202
transform 1 0 608 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5901_6
timestamp 1730589202
transform 1 0 664 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5901_6
timestamp 1730589202
transform 1 0 664 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5944_6
timestamp 1730589202
transform 1 0 712 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5944_6
timestamp 1730589202
transform 1 0 712 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5943_6
timestamp 1730589202
transform 1 0 760 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5943_6
timestamp 1730589202
transform 1 0 760 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5942_6
timestamp 1730589202
transform 1 0 808 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5942_6
timestamp 1730589202
transform 1 0 808 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5941_6
timestamp 1730589202
transform 1 0 856 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5941_6
timestamp 1730589202
transform 1 0 856 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5940_6
timestamp 1730589202
transform 1 0 912 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5940_6
timestamp 1730589202
transform 1 0 912 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5939_6
timestamp 1730589202
transform 1 0 968 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5939_6
timestamp 1730589202
transform 1 0 968 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5938_6
timestamp 1730589202
transform 1 0 1024 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5938_6
timestamp 1730589202
transform 1 0 1024 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5286_6
timestamp 1730589202
transform 1 0 1080 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5286_6
timestamp 1730589202
transform 1 0 1080 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5285_6
timestamp 1730589202
transform 1 0 1128 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5285_6
timestamp 1730589202
transform 1 0 1128 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5284_6
timestamp 1730589202
transform 1 0 1176 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5284_6
timestamp 1730589202
transform 1 0 1176 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5267_6
timestamp 1730589202
transform 1 0 1224 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5267_6
timestamp 1730589202
transform 1 0 1224 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5266_6
timestamp 1730589202
transform 1 0 1272 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5266_6
timestamp 1730589202
transform 1 0 1272 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5265_6
timestamp 1730589202
transform 1 0 1320 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5265_6
timestamp 1730589202
transform 1 0 1320 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5264_6
timestamp 1730589202
transform 1 0 1376 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5256_6
timestamp 1730589202
transform 1 0 1408 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5256_6
timestamp 1730589202
transform 1 0 1408 0 1 176
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5264_6
timestamp 1730589202
transform 1 0 1376 0 1 176
box 8 4 20 35
use welltap_svt  __well_tap__5
timestamp 1730589202
transform 1 0 1440 0 1 180
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730589202
transform 1 0 1440 0 1 180
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730589202
transform 1 0 104 0 -1 252
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730589202
transform 1 0 104 0 -1 252
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5887_6
timestamp 1730589202
transform 1 0 280 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5886_6
timestamp 1730589202
transform 1 0 256 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5886_6
timestamp 1730589202
transform 1 0 256 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5887_6
timestamp 1730589202
transform 1 0 280 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5888_6
timestamp 1730589202
transform 1 0 304 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5888_6
timestamp 1730589202
transform 1 0 304 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5974_6
timestamp 1730589202
transform 1 0 352 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5889_6
timestamp 1730589202
transform 1 0 328 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5889_6
timestamp 1730589202
transform 1 0 328 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5974_6
timestamp 1730589202
transform 1 0 352 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5973_6
timestamp 1730589202
transform 1 0 376 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5972_6
timestamp 1730589202
transform 1 0 400 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5972_6
timestamp 1730589202
transform 1 0 400 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5973_6
timestamp 1730589202
transform 1 0 376 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5890_6
timestamp 1730589202
transform 1 0 424 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5890_6
timestamp 1730589202
transform 1 0 424 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5891_6
timestamp 1730589202
transform 1 0 456 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5891_6
timestamp 1730589202
transform 1 0 456 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5892_6
timestamp 1730589202
transform 1 0 496 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5892_6
timestamp 1730589202
transform 1 0 496 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5893_6
timestamp 1730589202
transform 1 0 536 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5893_6
timestamp 1730589202
transform 1 0 536 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5950_6
timestamp 1730589202
transform 1 0 616 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5894_6
timestamp 1730589202
transform 1 0 576 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5894_6
timestamp 1730589202
transform 1 0 576 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5950_6
timestamp 1730589202
transform 1 0 616 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5949_6
timestamp 1730589202
transform 1 0 672 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5949_6
timestamp 1730589202
transform 1 0 672 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5948_6
timestamp 1730589202
transform 1 0 736 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5948_6
timestamp 1730589202
transform 1 0 736 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5947_6
timestamp 1730589202
transform 1 0 800 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5947_6
timestamp 1730589202
transform 1 0 800 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5946_6
timestamp 1730589202
transform 1 0 872 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5946_6
timestamp 1730589202
transform 1 0 872 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5945_6
timestamp 1730589202
transform 1 0 952 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5945_6
timestamp 1730589202
transform 1 0 952 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5287_6
timestamp 1730589202
transform 1 0 1032 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5287_6
timestamp 1730589202
transform 1 0 1032 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5288_6
timestamp 1730589202
transform 1 0 1112 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5288_6
timestamp 1730589202
transform 1 0 1112 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5289_6
timestamp 1730589202
transform 1 0 1192 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5289_6
timestamp 1730589202
transform 1 0 1192 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5290_6
timestamp 1730589202
transform 1 0 1272 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5290_6
timestamp 1730589202
transform 1 0 1272 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5254_6
timestamp 1730589202
transform 1 0 1352 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5254_6
timestamp 1730589202
transform 1 0 1352 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5255_6
timestamp 1730589202
transform 1 0 1408 0 -1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5255_6
timestamp 1730589202
transform 1 0 1408 0 -1 256
box 8 4 20 35
use welltap_svt  __well_tap__7
timestamp 1730589202
transform 1 0 1440 0 -1 252
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730589202
transform 1 0 1440 0 -1 252
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730589202
transform 1 0 104 0 1 260
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730589202
transform 1 0 104 0 1 260
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5880_6
timestamp 1730589202
transform 1 0 264 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5879_6
timestamp 1730589202
transform 1 0 240 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5879_6
timestamp 1730589202
transform 1 0 240 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5880_6
timestamp 1730589202
transform 1 0 264 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5882_6
timestamp 1730589202
transform 1 0 312 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5881_6
timestamp 1730589202
transform 1 0 288 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5881_6
timestamp 1730589202
transform 1 0 288 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5882_6
timestamp 1730589202
transform 1 0 312 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5884_6
timestamp 1730589202
transform 1 0 360 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5883_6
timestamp 1730589202
transform 1 0 336 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5883_6
timestamp 1730589202
transform 1 0 336 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5884_6
timestamp 1730589202
transform 1 0 360 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5885_6
timestamp 1730589202
transform 1 0 392 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5885_6
timestamp 1730589202
transform 1 0 392 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5971_6
timestamp 1730589202
transform 1 0 424 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5971_6
timestamp 1730589202
transform 1 0 424 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5970_6
timestamp 1730589202
transform 1 0 464 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5970_6
timestamp 1730589202
transform 1 0 464 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5969_6
timestamp 1730589202
transform 1 0 504 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5969_6
timestamp 1730589202
transform 1 0 504 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5954_6
timestamp 1730589202
transform 1 0 552 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5954_6
timestamp 1730589202
transform 1 0 552 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5953_6
timestamp 1730589202
transform 1 0 608 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5953_6
timestamp 1730589202
transform 1 0 608 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5952_6
timestamp 1730589202
transform 1 0 656 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5952_6
timestamp 1730589202
transform 1 0 656 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5951_6
timestamp 1730589202
transform 1 0 704 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5951_6
timestamp 1730589202
transform 1 0 704 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5332_6
timestamp 1730589202
transform 1 0 752 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5332_6
timestamp 1730589202
transform 1 0 752 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5331_6
timestamp 1730589202
transform 1 0 800 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5331_6
timestamp 1730589202
transform 1 0 800 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5330_6
timestamp 1730589202
transform 1 0 840 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5330_6
timestamp 1730589202
transform 1 0 840 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5329_6
timestamp 1730589202
transform 1 0 872 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5328_6
timestamp 1730589202
transform 1 0 896 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5328_6
timestamp 1730589202
transform 1 0 896 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5329_6
timestamp 1730589202
transform 1 0 872 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5327_6
timestamp 1730589202
transform 1 0 920 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5326_6
timestamp 1730589202
transform 1 0 944 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5326_6
timestamp 1730589202
transform 1 0 944 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5327_6
timestamp 1730589202
transform 1 0 920 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5325_6
timestamp 1730589202
transform 1 0 968 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5324_6
timestamp 1730589202
transform 1 0 992 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5324_6
timestamp 1730589202
transform 1 0 992 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5325_6
timestamp 1730589202
transform 1 0 968 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5323_6
timestamp 1730589202
transform 1 0 1016 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5323_6
timestamp 1730589202
transform 1 0 1016 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5322_6
timestamp 1730589202
transform 1 0 1040 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5321_6
timestamp 1730589202
transform 1 0 1064 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5321_6
timestamp 1730589202
transform 1 0 1064 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5322_6
timestamp 1730589202
transform 1 0 1040 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5320_6
timestamp 1730589202
transform 1 0 1088 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5319_6
timestamp 1730589202
transform 1 0 1120 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5319_6
timestamp 1730589202
transform 1 0 1120 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5320_6
timestamp 1730589202
transform 1 0 1088 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5318_6
timestamp 1730589202
transform 1 0 1152 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5318_6
timestamp 1730589202
transform 1 0 1152 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5317_6
timestamp 1730589202
transform 1 0 1192 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5317_6
timestamp 1730589202
transform 1 0 1192 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5316_6
timestamp 1730589202
transform 1 0 1240 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5316_6
timestamp 1730589202
transform 1 0 1240 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5291_6
timestamp 1730589202
transform 1 0 1296 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5291_6
timestamp 1730589202
transform 1 0 1296 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5292_6
timestamp 1730589202
transform 1 0 1360 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5292_6
timestamp 1730589202
transform 1 0 1360 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5253_6
timestamp 1730589202
transform 1 0 1408 0 1 256
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5253_6
timestamp 1730589202
transform 1 0 1408 0 1 256
box 8 4 20 35
use welltap_svt  __well_tap__9
timestamp 1730589202
transform 1 0 1440 0 1 260
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730589202
transform 1 0 1440 0 1 260
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730589202
transform 1 0 104 0 -1 332
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730589202
transform 1 0 104 0 -1 332
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5873_6
timestamp 1730589202
transform 1 0 192 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5872_6
timestamp 1730589202
transform 1 0 168 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5872_6
timestamp 1730589202
transform 1 0 168 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5873_6
timestamp 1730589202
transform 1 0 192 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5874_6
timestamp 1730589202
transform 1 0 216 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5874_6
timestamp 1730589202
transform 1 0 216 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5876_6
timestamp 1730589202
transform 1 0 272 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5875_6
timestamp 1730589202
transform 1 0 240 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5875_6
timestamp 1730589202
transform 1 0 240 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5876_6
timestamp 1730589202
transform 1 0 272 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5877_6
timestamp 1730589202
transform 1 0 312 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5877_6
timestamp 1730589202
transform 1 0 312 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5878_6
timestamp 1730589202
transform 1 0 352 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5878_6
timestamp 1730589202
transform 1 0 352 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5966_6
timestamp 1730589202
transform 1 0 392 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5966_6
timestamp 1730589202
transform 1 0 392 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5967_6
timestamp 1730589202
transform 1 0 432 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5967_6
timestamp 1730589202
transform 1 0 432 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5968_6
timestamp 1730589202
transform 1 0 472 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5968_6
timestamp 1730589202
transform 1 0 472 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5958_6
timestamp 1730589202
transform 1 0 520 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5958_6
timestamp 1730589202
transform 1 0 520 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5957_6
timestamp 1730589202
transform 1 0 576 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5957_6
timestamp 1730589202
transform 1 0 576 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5956_6
timestamp 1730589202
transform 1 0 632 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5956_6
timestamp 1730589202
transform 1 0 632 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5955_6
timestamp 1730589202
transform 1 0 680 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5955_6
timestamp 1730589202
transform 1 0 680 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5338_6
timestamp 1730589202
transform 1 0 728 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5338_6
timestamp 1730589202
transform 1 0 728 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5337_6
timestamp 1730589202
transform 1 0 784 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5337_6
timestamp 1730589202
transform 1 0 784 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5336_6
timestamp 1730589202
transform 1 0 840 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5336_6
timestamp 1730589202
transform 1 0 840 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5335_6
timestamp 1730589202
transform 1 0 888 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5335_6
timestamp 1730589202
transform 1 0 888 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5334_6
timestamp 1730589202
transform 1 0 936 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5334_6
timestamp 1730589202
transform 1 0 936 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5333_6
timestamp 1730589202
transform 1 0 984 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5333_6
timestamp 1730589202
transform 1 0 984 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5315_6
timestamp 1730589202
transform 1 0 1032 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5315_6
timestamp 1730589202
transform 1 0 1032 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5314_6
timestamp 1730589202
transform 1 0 1080 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5314_6
timestamp 1730589202
transform 1 0 1080 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5313_6
timestamp 1730589202
transform 1 0 1128 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5313_6
timestamp 1730589202
transform 1 0 1128 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5312_6
timestamp 1730589202
transform 1 0 1176 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5312_6
timestamp 1730589202
transform 1 0 1176 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5311_6
timestamp 1730589202
transform 1 0 1224 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5311_6
timestamp 1730589202
transform 1 0 1224 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5294_6
timestamp 1730589202
transform 1 0 1272 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5294_6
timestamp 1730589202
transform 1 0 1272 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5293_6
timestamp 1730589202
transform 1 0 1320 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5293_6
timestamp 1730589202
transform 1 0 1320 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5252_6
timestamp 1730589202
transform 1 0 1408 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5251_6
timestamp 1730589202
transform 1 0 1376 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5251_6
timestamp 1730589202
transform 1 0 1376 0 -1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5252_6
timestamp 1730589202
transform 1 0 1408 0 -1 336
box 8 4 20 35
use welltap_svt  __well_tap__11
timestamp 1730589202
transform 1 0 1440 0 -1 332
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730589202
transform 1 0 1440 0 -1 332
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730589202
transform 1 0 104 0 1 340
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730589202
transform 1 0 104 0 1 340
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5865_6
timestamp 1730589202
transform 1 0 152 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5864_6
timestamp 1730589202
transform 1 0 128 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5864_6
timestamp 1730589202
transform 1 0 128 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5865_6
timestamp 1730589202
transform 1 0 152 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5866_6
timestamp 1730589202
transform 1 0 176 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5866_6
timestamp 1730589202
transform 1 0 176 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5868_6
timestamp 1730589202
transform 1 0 224 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5867_6
timestamp 1730589202
transform 1 0 200 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5867_6
timestamp 1730589202
transform 1 0 200 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5868_6
timestamp 1730589202
transform 1 0 224 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5869_6
timestamp 1730589202
transform 1 0 248 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5869_6
timestamp 1730589202
transform 1 0 248 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5870_6
timestamp 1730589202
transform 1 0 288 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5870_6
timestamp 1730589202
transform 1 0 288 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5871_6
timestamp 1730589202
transform 1 0 328 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5871_6
timestamp 1730589202
transform 1 0 328 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5965_6
timestamp 1730589202
transform 1 0 368 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5965_6
timestamp 1730589202
transform 1 0 368 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5964_6
timestamp 1730589202
transform 1 0 408 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5963_6
timestamp 1730589202
transform 1 0 448 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5963_6
timestamp 1730589202
transform 1 0 448 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5964_6
timestamp 1730589202
transform 1 0 408 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5962_6
timestamp 1730589202
transform 1 0 488 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5962_6
timestamp 1730589202
transform 1 0 488 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5961_6
timestamp 1730589202
transform 1 0 528 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5961_6
timestamp 1730589202
transform 1 0 528 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5960_6
timestamp 1730589202
transform 1 0 568 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5960_6
timestamp 1730589202
transform 1 0 568 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5959_6
timestamp 1730589202
transform 1 0 608 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5959_6
timestamp 1730589202
transform 1 0 608 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5345_6
timestamp 1730589202
transform 1 0 648 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5345_6
timestamp 1730589202
transform 1 0 648 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5344_6
timestamp 1730589202
transform 1 0 680 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5344_6
timestamp 1730589202
transform 1 0 680 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5349_6
timestamp 1730589202
transform 1 0 720 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5349_6
timestamp 1730589202
transform 1 0 720 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5343_6
timestamp 1730589202
transform 1 0 768 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5343_6
timestamp 1730589202
transform 1 0 768 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5342_6
timestamp 1730589202
transform 1 0 824 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5342_6
timestamp 1730589202
transform 1 0 824 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5341_6
timestamp 1730589202
transform 1 0 880 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5341_6
timestamp 1730589202
transform 1 0 880 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5340_6
timestamp 1730589202
transform 1 0 944 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5340_6
timestamp 1730589202
transform 1 0 944 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5339_6
timestamp 1730589202
transform 1 0 1008 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5339_6
timestamp 1730589202
transform 1 0 1008 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5310_6
timestamp 1730589202
transform 1 0 1072 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5310_6
timestamp 1730589202
transform 1 0 1072 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5309_6
timestamp 1730589202
transform 1 0 1128 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5309_6
timestamp 1730589202
transform 1 0 1128 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5308_6
timestamp 1730589202
transform 1 0 1176 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5308_6
timestamp 1730589202
transform 1 0 1176 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5307_6
timestamp 1730589202
transform 1 0 1224 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5307_6
timestamp 1730589202
transform 1 0 1224 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5295_6
timestamp 1730589202
transform 1 0 1264 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5295_6
timestamp 1730589202
transform 1 0 1264 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5296_6
timestamp 1730589202
transform 1 0 1304 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5296_6
timestamp 1730589202
transform 1 0 1304 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5297_6
timestamp 1730589202
transform 1 0 1344 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5297_6
timestamp 1730589202
transform 1 0 1344 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5250_6
timestamp 1730589202
transform 1 0 1384 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5249_6
timestamp 1730589202
transform 1 0 1408 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5249_6
timestamp 1730589202
transform 1 0 1408 0 1 336
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5250_6
timestamp 1730589202
transform 1 0 1384 0 1 336
box 8 4 20 35
use welltap_svt  __well_tap__13
timestamp 1730589202
transform 1 0 1440 0 1 340
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730589202
transform 1 0 1440 0 1 340
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730589202
transform 1 0 104 0 -1 416
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730589202
transform 1 0 104 0 -1 416
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5860_6
timestamp 1730589202
transform 1 0 128 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5859_6
timestamp 1730589202
transform 1 0 152 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5859_6
timestamp 1730589202
transform 1 0 152 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5860_6
timestamp 1730589202
transform 1 0 128 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5858_6
timestamp 1730589202
transform 1 0 176 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5858_6
timestamp 1730589202
transform 1 0 176 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5857_6
timestamp 1730589202
transform 1 0 208 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5857_6
timestamp 1730589202
transform 1 0 208 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5861_6
timestamp 1730589202
transform 1 0 264 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5861_6
timestamp 1730589202
transform 1 0 264 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5862_6
timestamp 1730589202
transform 1 0 320 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5862_6
timestamp 1730589202
transform 1 0 320 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5863_6
timestamp 1730589202
transform 1 0 384 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5863_6
timestamp 1730589202
transform 1 0 384 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5355_6
timestamp 1730589202
transform 1 0 440 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5355_6
timestamp 1730589202
transform 1 0 440 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5354_6
timestamp 1730589202
transform 1 0 496 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5354_6
timestamp 1730589202
transform 1 0 496 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5353_6
timestamp 1730589202
transform 1 0 544 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5353_6
timestamp 1730589202
transform 1 0 544 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5352_6
timestamp 1730589202
transform 1 0 592 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5352_6
timestamp 1730589202
transform 1 0 592 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5351_6
timestamp 1730589202
transform 1 0 640 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5351_6
timestamp 1730589202
transform 1 0 640 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5350_6
timestamp 1730589202
transform 1 0 696 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5350_6
timestamp 1730589202
transform 1 0 696 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5348_6
timestamp 1730589202
transform 1 0 760 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5348_6
timestamp 1730589202
transform 1 0 760 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5347_6
timestamp 1730589202
transform 1 0 824 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5347_6
timestamp 1730589202
transform 1 0 824 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5346_6
timestamp 1730589202
transform 1 0 896 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5346_6
timestamp 1730589202
transform 1 0 896 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5389_6
timestamp 1730589202
transform 1 0 968 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5389_6
timestamp 1730589202
transform 1 0 968 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5390_6
timestamp 1730589202
transform 1 0 1032 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5390_6
timestamp 1730589202
transform 1 0 1032 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5306_6
timestamp 1730589202
transform 1 0 1096 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5306_6
timestamp 1730589202
transform 1 0 1096 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5305_6
timestamp 1730589202
transform 1 0 1152 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5305_6
timestamp 1730589202
transform 1 0 1152 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5304_6
timestamp 1730589202
transform 1 0 1200 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5304_6
timestamp 1730589202
transform 1 0 1200 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5303_6
timestamp 1730589202
transform 1 0 1240 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5303_6
timestamp 1730589202
transform 1 0 1240 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5302_6
timestamp 1730589202
transform 1 0 1272 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5302_6
timestamp 1730589202
transform 1 0 1272 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5300_6
timestamp 1730589202
transform 1 0 1312 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5300_6
timestamp 1730589202
transform 1 0 1312 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5299_6
timestamp 1730589202
transform 1 0 1352 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5299_6
timestamp 1730589202
transform 1 0 1352 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5298_6
timestamp 1730589202
transform 1 0 1384 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5248_6
timestamp 1730589202
transform 1 0 1408 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5248_6
timestamp 1730589202
transform 1 0 1408 0 -1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5298_6
timestamp 1730589202
transform 1 0 1384 0 -1 420
box 8 4 20 35
use welltap_svt  __well_tap__15
timestamp 1730589202
transform 1 0 1440 0 -1 416
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730589202
transform 1 0 1440 0 -1 416
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730589202
transform 1 0 104 0 1 424
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730589202
transform 1 0 104 0 1 424
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5856_6
timestamp 1730589202
transform 1 0 128 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5855_6
timestamp 1730589202
transform 1 0 152 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5855_6
timestamp 1730589202
transform 1 0 152 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5856_6
timestamp 1730589202
transform 1 0 128 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5854_6
timestamp 1730589202
transform 1 0 184 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5854_6
timestamp 1730589202
transform 1 0 184 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5853_6
timestamp 1730589202
transform 1 0 232 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5853_6
timestamp 1730589202
transform 1 0 232 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5852_6
timestamp 1730589202
transform 1 0 288 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5852_6
timestamp 1730589202
transform 1 0 288 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5851_6
timestamp 1730589202
transform 1 0 344 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5851_6
timestamp 1730589202
transform 1 0 344 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5359_6
timestamp 1730589202
transform 1 0 408 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5359_6
timestamp 1730589202
transform 1 0 408 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5358_6
timestamp 1730589202
transform 1 0 472 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5358_6
timestamp 1730589202
transform 1 0 472 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5357_6
timestamp 1730589202
transform 1 0 536 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5357_6
timestamp 1730589202
transform 1 0 536 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5356_6
timestamp 1730589202
transform 1 0 600 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5356_6
timestamp 1730589202
transform 1 0 600 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5373_6
timestamp 1730589202
transform 1 0 664 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5373_6
timestamp 1730589202
transform 1 0 664 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5374_6
timestamp 1730589202
transform 1 0 728 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5374_6
timestamp 1730589202
transform 1 0 728 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5383_6
timestamp 1730589202
transform 1 0 784 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5383_6
timestamp 1730589202
transform 1 0 784 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5384_6
timestamp 1730589202
transform 1 0 832 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5384_6
timestamp 1730589202
transform 1 0 832 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5386_6
timestamp 1730589202
transform 1 0 904 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5385_6
timestamp 1730589202
transform 1 0 872 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5385_6
timestamp 1730589202
transform 1 0 872 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5386_6
timestamp 1730589202
transform 1 0 904 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5387_6
timestamp 1730589202
transform 1 0 936 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5387_6
timestamp 1730589202
transform 1 0 936 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5391_6
timestamp 1730589202
transform 1 0 992 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5388_6
timestamp 1730589202
transform 1 0 960 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5388_6
timestamp 1730589202
transform 1 0 960 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5391_6
timestamp 1730589202
transform 1 0 992 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5392_6
timestamp 1730589202
transform 1 0 1024 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5392_6
timestamp 1730589202
transform 1 0 1024 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5393_6
timestamp 1730589202
transform 1 0 1064 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5393_6
timestamp 1730589202
transform 1 0 1064 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5394_6
timestamp 1730589202
transform 1 0 1112 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5394_6
timestamp 1730589202
transform 1 0 1112 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5395_6
timestamp 1730589202
transform 1 0 1168 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5395_6
timestamp 1730589202
transform 1 0 1168 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5396_6
timestamp 1730589202
transform 1 0 1232 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5396_6
timestamp 1730589202
transform 1 0 1232 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5301_6
timestamp 1730589202
transform 1 0 1296 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5301_6
timestamp 1730589202
transform 1 0 1296 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5246_6
timestamp 1730589202
transform 1 0 1360 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5246_6
timestamp 1730589202
transform 1 0 1360 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5247_6
timestamp 1730589202
transform 1 0 1408 0 1 420
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5247_6
timestamp 1730589202
transform 1 0 1408 0 1 420
box 8 4 20 35
use welltap_svt  __well_tap__17
timestamp 1730589202
transform 1 0 1440 0 1 424
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730589202
transform 1 0 1440 0 1 424
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730589202
transform 1 0 104 0 -1 496
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730589202
transform 1 0 104 0 -1 496
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5850_6
timestamp 1730589202
transform 1 0 128 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5849_6
timestamp 1730589202
transform 1 0 152 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5849_6
timestamp 1730589202
transform 1 0 152 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5850_6
timestamp 1730589202
transform 1 0 128 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5848_6
timestamp 1730589202
transform 1 0 176 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5848_6
timestamp 1730589202
transform 1 0 176 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5847_6
timestamp 1730589202
transform 1 0 216 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5847_6
timestamp 1730589202
transform 1 0 216 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5846_6
timestamp 1730589202
transform 1 0 264 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5846_6
timestamp 1730589202
transform 1 0 264 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5845_6
timestamp 1730589202
transform 1 0 312 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5845_6
timestamp 1730589202
transform 1 0 312 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5844_6
timestamp 1730589202
transform 1 0 368 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5844_6
timestamp 1730589202
transform 1 0 368 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5360_6
timestamp 1730589202
transform 1 0 424 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5360_6
timestamp 1730589202
transform 1 0 424 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5361_6
timestamp 1730589202
transform 1 0 480 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5361_6
timestamp 1730589202
transform 1 0 480 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5370_6
timestamp 1730589202
transform 1 0 536 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5370_6
timestamp 1730589202
transform 1 0 536 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5371_6
timestamp 1730589202
transform 1 0 584 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5371_6
timestamp 1730589202
transform 1 0 584 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5375_6
timestamp 1730589202
transform 1 0 656 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5372_6
timestamp 1730589202
transform 1 0 624 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5372_6
timestamp 1730589202
transform 1 0 624 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5375_6
timestamp 1730589202
transform 1 0 656 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5376_6
timestamp 1730589202
transform 1 0 680 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5376_6
timestamp 1730589202
transform 1 0 680 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5377_6
timestamp 1730589202
transform 1 0 712 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5377_6
timestamp 1730589202
transform 1 0 712 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5378_6
timestamp 1730589202
transform 1 0 752 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5378_6
timestamp 1730589202
transform 1 0 752 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5379_6
timestamp 1730589202
transform 1 0 792 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5379_6
timestamp 1730589202
transform 1 0 792 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5380_6
timestamp 1730589202
transform 1 0 840 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5380_6
timestamp 1730589202
transform 1 0 840 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5381_6
timestamp 1730589202
transform 1 0 896 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5381_6
timestamp 1730589202
transform 1 0 896 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5382_6
timestamp 1730589202
transform 1 0 944 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5382_6
timestamp 1730589202
transform 1 0 944 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5397_6
timestamp 1730589202
transform 1 0 992 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5397_6
timestamp 1730589202
transform 1 0 992 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5398_6
timestamp 1730589202
transform 1 0 1040 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5398_6
timestamp 1730589202
transform 1 0 1040 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5399_6
timestamp 1730589202
transform 1 0 1088 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5399_6
timestamp 1730589202
transform 1 0 1088 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5400_6
timestamp 1730589202
transform 1 0 1136 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5400_6
timestamp 1730589202
transform 1 0 1136 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5401_6
timestamp 1730589202
transform 1 0 1192 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5401_6
timestamp 1730589202
transform 1 0 1192 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5402_6
timestamp 1730589202
transform 1 0 1248 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5402_6
timestamp 1730589202
transform 1 0 1248 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5403_6
timestamp 1730589202
transform 1 0 1304 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5403_6
timestamp 1730589202
transform 1 0 1304 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5245_6
timestamp 1730589202
transform 1 0 1368 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5245_6
timestamp 1730589202
transform 1 0 1368 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5244_6
timestamp 1730589202
transform 1 0 1408 0 -1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5244_6
timestamp 1730589202
transform 1 0 1408 0 -1 500
box 8 4 20 35
use welltap_svt  __well_tap__19
timestamp 1730589202
transform 1 0 1440 0 -1 496
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730589202
transform 1 0 1440 0 -1 496
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730589202
transform 1 0 104 0 1 504
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730589202
transform 1 0 104 0 1 504
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5843_6
timestamp 1730589202
transform 1 0 216 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5843_6
timestamp 1730589202
transform 1 0 216 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5842_6
timestamp 1730589202
transform 1 0 240 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5841_6
timestamp 1730589202
transform 1 0 264 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5841_6
timestamp 1730589202
transform 1 0 264 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5842_6
timestamp 1730589202
transform 1 0 240 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5840_6
timestamp 1730589202
transform 1 0 288 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5839_6
timestamp 1730589202
transform 1 0 320 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5839_6
timestamp 1730589202
transform 1 0 320 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5840_6
timestamp 1730589202
transform 1 0 288 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5838_6
timestamp 1730589202
transform 1 0 352 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5838_6
timestamp 1730589202
transform 1 0 352 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5837_6
timestamp 1730589202
transform 1 0 384 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5837_6
timestamp 1730589202
transform 1 0 384 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5363_6
timestamp 1730589202
transform 1 0 448 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5362_6
timestamp 1730589202
transform 1 0 416 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5362_6
timestamp 1730589202
transform 1 0 416 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5363_6
timestamp 1730589202
transform 1 0 448 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5364_6
timestamp 1730589202
transform 1 0 480 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5364_6
timestamp 1730589202
transform 1 0 480 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5366_6
timestamp 1730589202
transform 1 0 520 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5366_6
timestamp 1730589202
transform 1 0 520 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5367_6
timestamp 1730589202
transform 1 0 568 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5367_6
timestamp 1730589202
transform 1 0 568 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5368_6
timestamp 1730589202
transform 1 0 616 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5368_6
timestamp 1730589202
transform 1 0 616 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5369_6
timestamp 1730589202
transform 1 0 664 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5369_6
timestamp 1730589202
transform 1 0 664 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5437_6
timestamp 1730589202
transform 1 0 704 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5437_6
timestamp 1730589202
transform 1 0 704 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5436_6
timestamp 1730589202
transform 1 0 752 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5436_6
timestamp 1730589202
transform 1 0 752 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5435_6
timestamp 1730589202
transform 1 0 800 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5435_6
timestamp 1730589202
transform 1 0 800 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5434_6
timestamp 1730589202
transform 1 0 848 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5434_6
timestamp 1730589202
transform 1 0 848 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5433_6
timestamp 1730589202
transform 1 0 904 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5433_6
timestamp 1730589202
transform 1 0 904 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5432_6
timestamp 1730589202
transform 1 0 960 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5432_6
timestamp 1730589202
transform 1 0 960 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5431_6
timestamp 1730589202
transform 1 0 1016 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5431_6
timestamp 1730589202
transform 1 0 1016 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5407_6
timestamp 1730589202
transform 1 0 1072 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5407_6
timestamp 1730589202
transform 1 0 1072 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5406_6
timestamp 1730589202
transform 1 0 1120 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5406_6
timestamp 1730589202
transform 1 0 1120 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5405_6
timestamp 1730589202
transform 1 0 1168 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5405_6
timestamp 1730589202
transform 1 0 1168 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5404_6
timestamp 1730589202
transform 1 0 1216 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5404_6
timestamp 1730589202
transform 1 0 1216 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5239_6
timestamp 1730589202
transform 1 0 1264 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5239_6
timestamp 1730589202
transform 1 0 1264 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5240_6
timestamp 1730589202
transform 1 0 1304 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5240_6
timestamp 1730589202
transform 1 0 1304 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5241_6
timestamp 1730589202
transform 1 0 1344 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5241_6
timestamp 1730589202
transform 1 0 1344 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5243_6
timestamp 1730589202
transform 1 0 1408 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5242_6
timestamp 1730589202
transform 1 0 1384 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5242_6
timestamp 1730589202
transform 1 0 1384 0 1 500
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5243_6
timestamp 1730589202
transform 1 0 1408 0 1 500
box 8 4 20 35
use welltap_svt  __well_tap__21
timestamp 1730589202
transform 1 0 1440 0 1 504
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730589202
transform 1 0 1440 0 1 504
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730589202
transform 1 0 104 0 -1 576
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730589202
transform 1 0 104 0 -1 576
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5836_6
timestamp 1730589202
transform 1 0 256 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5835_6
timestamp 1730589202
transform 1 0 280 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5835_6
timestamp 1730589202
transform 1 0 280 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5836_6
timestamp 1730589202
transform 1 0 256 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5834_6
timestamp 1730589202
transform 1 0 304 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5834_6
timestamp 1730589202
transform 1 0 304 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5833_6
timestamp 1730589202
transform 1 0 328 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5832_6
timestamp 1730589202
transform 1 0 352 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5832_6
timestamp 1730589202
transform 1 0 352 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5833_6
timestamp 1730589202
transform 1 0 328 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5831_6
timestamp 1730589202
transform 1 0 376 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5830_6
timestamp 1730589202
transform 1 0 400 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5830_6
timestamp 1730589202
transform 1 0 400 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5831_6
timestamp 1730589202
transform 1 0 376 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5571_6
timestamp 1730589202
transform 1 0 424 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5571_6
timestamp 1730589202
transform 1 0 424 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5570_6
timestamp 1730589202
transform 1 0 456 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5570_6
timestamp 1730589202
transform 1 0 456 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5365_6
timestamp 1730589202
transform 1 0 496 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5365_6
timestamp 1730589202
transform 1 0 496 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5569_6
timestamp 1730589202
transform 1 0 544 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5569_6
timestamp 1730589202
transform 1 0 544 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5567_6
timestamp 1730589202
transform 1 0 600 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5567_6
timestamp 1730589202
transform 1 0 600 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5568_6
timestamp 1730589202
transform 1 0 656 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5568_6
timestamp 1730589202
transform 1 0 656 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5438_6
timestamp 1730589202
transform 1 0 712 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5438_6
timestamp 1730589202
transform 1 0 712 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5439_6
timestamp 1730589202
transform 1 0 768 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5439_6
timestamp 1730589202
transform 1 0 768 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5430_6
timestamp 1730589202
transform 1 0 824 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5430_6
timestamp 1730589202
transform 1 0 824 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5429_6
timestamp 1730589202
transform 1 0 880 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5429_6
timestamp 1730589202
transform 1 0 880 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5428_6
timestamp 1730589202
transform 1 0 936 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5428_6
timestamp 1730589202
transform 1 0 936 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5427_6
timestamp 1730589202
transform 1 0 1000 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5427_6
timestamp 1730589202
transform 1 0 1000 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5408_6
timestamp 1730589202
transform 1 0 1064 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5408_6
timestamp 1730589202
transform 1 0 1064 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5409_6
timestamp 1730589202
transform 1 0 1120 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5409_6
timestamp 1730589202
transform 1 0 1120 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5410_6
timestamp 1730589202
transform 1 0 1176 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5410_6
timestamp 1730589202
transform 1 0 1176 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5238_6
timestamp 1730589202
transform 1 0 1240 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5238_6
timestamp 1730589202
transform 1 0 1240 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5237_6
timestamp 1730589202
transform 1 0 1304 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5237_6
timestamp 1730589202
transform 1 0 1304 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5236_6
timestamp 1730589202
transform 1 0 1368 0 -1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5236_6
timestamp 1730589202
transform 1 0 1368 0 -1 580
box 8 4 20 35
use welltap_svt  __well_tap__23
timestamp 1730589202
transform 1 0 1440 0 -1 576
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730589202
transform 1 0 1440 0 -1 576
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730589202
transform 1 0 104 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730589202
transform 1 0 104 0 1 584
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5824_6
timestamp 1730589202
transform 1 0 264 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5824_6
timestamp 1730589202
transform 1 0 264 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5826_6
timestamp 1730589202
transform 1 0 312 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5825_6
timestamp 1730589202
transform 1 0 288 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5825_6
timestamp 1730589202
transform 1 0 288 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5826_6
timestamp 1730589202
transform 1 0 312 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5828_6
timestamp 1730589202
transform 1 0 360 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5827_6
timestamp 1730589202
transform 1 0 336 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5827_6
timestamp 1730589202
transform 1 0 336 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5828_6
timestamp 1730589202
transform 1 0 360 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5829_6
timestamp 1730589202
transform 1 0 384 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5829_6
timestamp 1730589202
transform 1 0 384 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5573_6
timestamp 1730589202
transform 1 0 432 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5572_6
timestamp 1730589202
transform 1 0 408 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5572_6
timestamp 1730589202
transform 1 0 408 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5573_6
timestamp 1730589202
transform 1 0 432 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5574_6
timestamp 1730589202
transform 1 0 472 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5574_6
timestamp 1730589202
transform 1 0 472 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5575_6
timestamp 1730589202
transform 1 0 512 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5575_6
timestamp 1730589202
transform 1 0 512 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5566_6
timestamp 1730589202
transform 1 0 560 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5566_6
timestamp 1730589202
transform 1 0 560 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5565_6
timestamp 1730589202
transform 1 0 616 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5565_6
timestamp 1730589202
transform 1 0 616 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5564_6
timestamp 1730589202
transform 1 0 672 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5564_6
timestamp 1730589202
transform 1 0 672 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5441_6
timestamp 1730589202
transform 1 0 728 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5441_6
timestamp 1730589202
transform 1 0 728 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5440_6
timestamp 1730589202
transform 1 0 776 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5440_6
timestamp 1730589202
transform 1 0 776 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5426_6
timestamp 1730589202
transform 1 0 824 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5426_6
timestamp 1730589202
transform 1 0 824 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5425_6
timestamp 1730589202
transform 1 0 872 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5425_6
timestamp 1730589202
transform 1 0 872 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5424_6
timestamp 1730589202
transform 1 0 920 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5424_6
timestamp 1730589202
transform 1 0 920 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5423_6
timestamp 1730589202
transform 1 0 968 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5423_6
timestamp 1730589202
transform 1 0 968 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5414_6
timestamp 1730589202
transform 1 0 1016 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5414_6
timestamp 1730589202
transform 1 0 1016 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5413_6
timestamp 1730589202
transform 1 0 1064 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5413_6
timestamp 1730589202
transform 1 0 1064 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5412_6
timestamp 1730589202
transform 1 0 1104 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5412_6
timestamp 1730589202
transform 1 0 1104 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5411_6
timestamp 1730589202
transform 1 0 1144 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5411_6
timestamp 1730589202
transform 1 0 1144 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5232_6
timestamp 1730589202
transform 1 0 1184 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5232_6
timestamp 1730589202
transform 1 0 1184 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5233_6
timestamp 1730589202
transform 1 0 1232 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5233_6
timestamp 1730589202
transform 1 0 1232 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5234_6
timestamp 1730589202
transform 1 0 1280 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5234_6
timestamp 1730589202
transform 1 0 1280 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5235_6
timestamp 1730589202
transform 1 0 1328 0 1 580
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5235_6
timestamp 1730589202
transform 1 0 1328 0 1 580
box 8 4 20 35
use welltap_svt  __well_tap__25
timestamp 1730589202
transform 1 0 1440 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730589202
transform 1 0 1440 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730589202
transform 1 0 104 0 -1 656
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730589202
transform 1 0 104 0 -1 656
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5817_6
timestamp 1730589202
transform 1 0 184 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5817_6
timestamp 1730589202
transform 1 0 184 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5819_6
timestamp 1730589202
transform 1 0 232 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5818_6
timestamp 1730589202
transform 1 0 208 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5818_6
timestamp 1730589202
transform 1 0 208 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5819_6
timestamp 1730589202
transform 1 0 232 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5820_6
timestamp 1730589202
transform 1 0 256 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5820_6
timestamp 1730589202
transform 1 0 256 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5822_6
timestamp 1730589202
transform 1 0 320 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5821_6
timestamp 1730589202
transform 1 0 288 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5821_6
timestamp 1730589202
transform 1 0 288 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5822_6
timestamp 1730589202
transform 1 0 320 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5823_6
timestamp 1730589202
transform 1 0 360 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5823_6
timestamp 1730589202
transform 1 0 360 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5576_6
timestamp 1730589202
transform 1 0 400 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5576_6
timestamp 1730589202
transform 1 0 400 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5577_6
timestamp 1730589202
transform 1 0 448 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5577_6
timestamp 1730589202
transform 1 0 448 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5578_6
timestamp 1730589202
transform 1 0 496 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5578_6
timestamp 1730589202
transform 1 0 496 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5579_6
timestamp 1730589202
transform 1 0 544 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5579_6
timestamp 1730589202
transform 1 0 544 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5561_6
timestamp 1730589202
transform 1 0 600 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5561_6
timestamp 1730589202
transform 1 0 600 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5562_6
timestamp 1730589202
transform 1 0 656 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5562_6
timestamp 1730589202
transform 1 0 656 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5563_6
timestamp 1730589202
transform 1 0 712 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5563_6
timestamp 1730589202
transform 1 0 712 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5442_6
timestamp 1730589202
transform 1 0 760 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5442_6
timestamp 1730589202
transform 1 0 760 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5443_6
timestamp 1730589202
transform 1 0 808 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5443_6
timestamp 1730589202
transform 1 0 808 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5422_6
timestamp 1730589202
transform 1 0 856 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5422_6
timestamp 1730589202
transform 1 0 856 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5421_6
timestamp 1730589202
transform 1 0 896 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5421_6
timestamp 1730589202
transform 1 0 896 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5420_6
timestamp 1730589202
transform 1 0 928 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5420_6
timestamp 1730589202
transform 1 0 928 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5419_6
timestamp 1730589202
transform 1 0 960 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5419_6
timestamp 1730589202
transform 1 0 960 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5418_6
timestamp 1730589202
transform 1 0 1000 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5418_6
timestamp 1730589202
transform 1 0 1000 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5417_6
timestamp 1730589202
transform 1 0 1040 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5417_6
timestamp 1730589202
transform 1 0 1040 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5416_6
timestamp 1730589202
transform 1 0 1080 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5415_6
timestamp 1730589202
transform 1 0 1120 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5415_6
timestamp 1730589202
transform 1 0 1120 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5416_6
timestamp 1730589202
transform 1 0 1080 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5226_6
timestamp 1730589202
transform 1 0 1152 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5226_6
timestamp 1730589202
transform 1 0 1152 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5227_6
timestamp 1730589202
transform 1 0 1184 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5227_6
timestamp 1730589202
transform 1 0 1184 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5228_6
timestamp 1730589202
transform 1 0 1216 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5228_6
timestamp 1730589202
transform 1 0 1216 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5229_6
timestamp 1730589202
transform 1 0 1256 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5229_6
timestamp 1730589202
transform 1 0 1256 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5230_6
timestamp 1730589202
transform 1 0 1296 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5230_6
timestamp 1730589202
transform 1 0 1296 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5231_6
timestamp 1730589202
transform 1 0 1336 0 -1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5231_6
timestamp 1730589202
transform 1 0 1336 0 -1 660
box 8 4 20 35
use welltap_svt  __well_tap__27
timestamp 1730589202
transform 1 0 1440 0 -1 656
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730589202
transform 1 0 1440 0 -1 656
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730589202
transform 1 0 104 0 1 664
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730589202
transform 1 0 104 0 1 664
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5812_6
timestamp 1730589202
transform 1 0 152 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5811_6
timestamp 1730589202
transform 1 0 128 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5811_6
timestamp 1730589202
transform 1 0 128 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5812_6
timestamp 1730589202
transform 1 0 152 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5813_6
timestamp 1730589202
transform 1 0 192 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5813_6
timestamp 1730589202
transform 1 0 192 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5814_6
timestamp 1730589202
transform 1 0 232 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5814_6
timestamp 1730589202
transform 1 0 232 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5815_6
timestamp 1730589202
transform 1 0 280 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5815_6
timestamp 1730589202
transform 1 0 280 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5816_6
timestamp 1730589202
transform 1 0 328 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5816_6
timestamp 1730589202
transform 1 0 328 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5580_6
timestamp 1730589202
transform 1 0 384 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5580_6
timestamp 1730589202
transform 1 0 384 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5581_6
timestamp 1730589202
transform 1 0 432 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5581_6
timestamp 1730589202
transform 1 0 432 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5582_6
timestamp 1730589202
transform 1 0 480 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5582_6
timestamp 1730589202
transform 1 0 480 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5583_6
timestamp 1730589202
transform 1 0 528 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5583_6
timestamp 1730589202
transform 1 0 528 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5584_6
timestamp 1730589202
transform 1 0 576 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5584_6
timestamp 1730589202
transform 1 0 576 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5560_6
timestamp 1730589202
transform 1 0 632 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5560_6
timestamp 1730589202
transform 1 0 632 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5559_6
timestamp 1730589202
transform 1 0 688 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5559_6
timestamp 1730589202
transform 1 0 688 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5558_6
timestamp 1730589202
transform 1 0 752 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5558_6
timestamp 1730589202
transform 1 0 752 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5446_6
timestamp 1730589202
transform 1 0 824 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5446_6
timestamp 1730589202
transform 1 0 824 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5445_6
timestamp 1730589202
transform 1 0 896 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5445_6
timestamp 1730589202
transform 1 0 896 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5444_6
timestamp 1730589202
transform 1 0 960 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5444_6
timestamp 1730589202
transform 1 0 960 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5225_6
timestamp 1730589202
transform 1 0 1024 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5225_6
timestamp 1730589202
transform 1 0 1024 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5224_6
timestamp 1730589202
transform 1 0 1080 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5224_6
timestamp 1730589202
transform 1 0 1080 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5223_6
timestamp 1730589202
transform 1 0 1128 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5223_6
timestamp 1730589202
transform 1 0 1128 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5222_6
timestamp 1730589202
transform 1 0 1168 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5222_6
timestamp 1730589202
transform 1 0 1168 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5221_6
timestamp 1730589202
transform 1 0 1208 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5220_6
timestamp 1730589202
transform 1 0 1240 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5220_6
timestamp 1730589202
transform 1 0 1240 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5221_6
timestamp 1730589202
transform 1 0 1208 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5219_6
timestamp 1730589202
transform 1 0 1272 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5219_6
timestamp 1730589202
transform 1 0 1272 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5215_6
timestamp 1730589202
transform 1 0 1304 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5215_6
timestamp 1730589202
transform 1 0 1304 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5214_6
timestamp 1730589202
transform 1 0 1336 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5213_6
timestamp 1730589202
transform 1 0 1360 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5213_6
timestamp 1730589202
transform 1 0 1360 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5214_6
timestamp 1730589202
transform 1 0 1336 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5212_6
timestamp 1730589202
transform 1 0 1384 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5211_6
timestamp 1730589202
transform 1 0 1408 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5211_6
timestamp 1730589202
transform 1 0 1408 0 1 660
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5212_6
timestamp 1730589202
transform 1 0 1384 0 1 660
box 8 4 20 35
use welltap_svt  __well_tap__29
timestamp 1730589202
transform 1 0 1440 0 1 664
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730589202
transform 1 0 1440 0 1 664
box 8 4 12 24
use welltap_svt  __well_tap__30
timestamp 1730589202
transform 1 0 104 0 -1 736
box 8 4 12 24
use welltap_svt  __well_tap__30
timestamp 1730589202
transform 1 0 104 0 -1 736
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5805_6
timestamp 1730589202
transform 1 0 152 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5804_6
timestamp 1730589202
transform 1 0 128 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5804_6
timestamp 1730589202
transform 1 0 128 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5805_6
timestamp 1730589202
transform 1 0 152 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5806_6
timestamp 1730589202
transform 1 0 176 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5806_6
timestamp 1730589202
transform 1 0 176 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5807_6
timestamp 1730589202
transform 1 0 208 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5807_6
timestamp 1730589202
transform 1 0 208 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5808_6
timestamp 1730589202
transform 1 0 256 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5808_6
timestamp 1730589202
transform 1 0 256 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5809_6
timestamp 1730589202
transform 1 0 312 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5809_6
timestamp 1730589202
transform 1 0 312 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5810_6
timestamp 1730589202
transform 1 0 368 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5810_6
timestamp 1730589202
transform 1 0 368 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5585_6
timestamp 1730589202
transform 1 0 416 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5585_6
timestamp 1730589202
transform 1 0 416 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5586_6
timestamp 1730589202
transform 1 0 464 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5586_6
timestamp 1730589202
transform 1 0 464 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5587_6
timestamp 1730589202
transform 1 0 512 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5587_6
timestamp 1730589202
transform 1 0 512 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5588_6
timestamp 1730589202
transform 1 0 560 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5588_6
timestamp 1730589202
transform 1 0 560 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5589_6
timestamp 1730589202
transform 1 0 608 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5589_6
timestamp 1730589202
transform 1 0 608 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5590_6
timestamp 1730589202
transform 1 0 656 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5590_6
timestamp 1730589202
transform 1 0 656 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5557_6
timestamp 1730589202
transform 1 0 696 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5557_6
timestamp 1730589202
transform 1 0 696 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5556_6
timestamp 1730589202
transform 1 0 744 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5556_6
timestamp 1730589202
transform 1 0 744 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5447_6
timestamp 1730589202
transform 1 0 800 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5447_6
timestamp 1730589202
transform 1 0 800 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5448_6
timestamp 1730589202
transform 1 0 864 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5448_6
timestamp 1730589202
transform 1 0 864 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5449_6
timestamp 1730589202
transform 1 0 936 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5449_6
timestamp 1730589202
transform 1 0 936 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5450_6
timestamp 1730589202
transform 1 0 1008 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5450_6
timestamp 1730589202
transform 1 0 1008 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5451_6
timestamp 1730589202
transform 1 0 1080 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5451_6
timestamp 1730589202
transform 1 0 1080 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5218_6
timestamp 1730589202
transform 1 0 1144 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5218_6
timestamp 1730589202
transform 1 0 1144 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5217_6
timestamp 1730589202
transform 1 0 1208 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5217_6
timestamp 1730589202
transform 1 0 1208 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5216_6
timestamp 1730589202
transform 1 0 1264 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5216_6
timestamp 1730589202
transform 1 0 1264 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5208_6
timestamp 1730589202
transform 1 0 1320 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5208_6
timestamp 1730589202
transform 1 0 1320 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5210_6
timestamp 1730589202
transform 1 0 1408 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5209_6
timestamp 1730589202
transform 1 0 1376 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5209_6
timestamp 1730589202
transform 1 0 1376 0 -1 740
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5210_6
timestamp 1730589202
transform 1 0 1408 0 -1 740
box 8 4 20 35
use welltap_svt  __well_tap__31
timestamp 1730589202
transform 1 0 1440 0 -1 736
box 8 4 12 24
use welltap_svt  __well_tap__31
timestamp 1730589202
transform 1 0 1440 0 -1 736
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730589202
transform 1 0 104 0 1 748
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730589202
transform 1 0 104 0 1 748
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5803_6
timestamp 1730589202
transform 1 0 128 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5802_6
timestamp 1730589202
transform 1 0 152 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5802_6
timestamp 1730589202
transform 1 0 152 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5803_6
timestamp 1730589202
transform 1 0 128 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5801_6
timestamp 1730589202
transform 1 0 176 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5801_6
timestamp 1730589202
transform 1 0 176 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5800_6
timestamp 1730589202
transform 1 0 216 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5800_6
timestamp 1730589202
transform 1 0 216 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5799_6
timestamp 1730589202
transform 1 0 272 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5799_6
timestamp 1730589202
transform 1 0 272 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5798_6
timestamp 1730589202
transform 1 0 336 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5798_6
timestamp 1730589202
transform 1 0 336 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5797_6
timestamp 1730589202
transform 1 0 400 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5797_6
timestamp 1730589202
transform 1 0 400 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5591_6
timestamp 1730589202
transform 1 0 456 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5591_6
timestamp 1730589202
transform 1 0 456 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5592_6
timestamp 1730589202
transform 1 0 512 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5592_6
timestamp 1730589202
transform 1 0 512 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5593_6
timestamp 1730589202
transform 1 0 568 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5593_6
timestamp 1730589202
transform 1 0 568 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5594_6
timestamp 1730589202
transform 1 0 616 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5594_6
timestamp 1730589202
transform 1 0 616 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5595_6
timestamp 1730589202
transform 1 0 664 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5595_6
timestamp 1730589202
transform 1 0 664 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5596_6
timestamp 1730589202
transform 1 0 712 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5596_6
timestamp 1730589202
transform 1 0 712 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5555_6
timestamp 1730589202
transform 1 0 752 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5555_6
timestamp 1730589202
transform 1 0 752 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5554_6
timestamp 1730589202
transform 1 0 792 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5554_6
timestamp 1730589202
transform 1 0 792 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5452_6
timestamp 1730589202
transform 1 0 832 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5452_6
timestamp 1730589202
transform 1 0 832 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5453_6
timestamp 1730589202
transform 1 0 872 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5453_6
timestamp 1730589202
transform 1 0 872 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5455_6
timestamp 1730589202
transform 1 0 952 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5454_6
timestamp 1730589202
transform 1 0 912 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5454_6
timestamp 1730589202
transform 1 0 912 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5455_6
timestamp 1730589202
transform 1 0 952 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5465_6
timestamp 1730589202
transform 1 0 984 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5465_6
timestamp 1730589202
transform 1 0 984 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5466_6
timestamp 1730589202
transform 1 0 1016 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5466_6
timestamp 1730589202
transform 1 0 1016 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5467_6
timestamp 1730589202
transform 1 0 1048 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5467_6
timestamp 1730589202
transform 1 0 1048 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5469_6
timestamp 1730589202
transform 1 0 1120 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5468_6
timestamp 1730589202
transform 1 0 1080 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5468_6
timestamp 1730589202
transform 1 0 1080 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5469_6
timestamp 1730589202
transform 1 0 1120 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5470_6
timestamp 1730589202
transform 1 0 1168 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5470_6
timestamp 1730589202
transform 1 0 1168 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5471_6
timestamp 1730589202
transform 1 0 1224 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5471_6
timestamp 1730589202
transform 1 0 1224 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5472_6
timestamp 1730589202
transform 1 0 1288 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5472_6
timestamp 1730589202
transform 1 0 1288 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5207_6
timestamp 1730589202
transform 1 0 1360 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5207_6
timestamp 1730589202
transform 1 0 1360 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5206_6
timestamp 1730589202
transform 1 0 1408 0 1 744
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5206_6
timestamp 1730589202
transform 1 0 1408 0 1 744
box 8 4 20 35
use welltap_svt  __well_tap__33
timestamp 1730589202
transform 1 0 1440 0 1 748
box 8 4 12 24
use welltap_svt  __well_tap__33
timestamp 1730589202
transform 1 0 1440 0 1 748
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730589202
transform 1 0 104 0 -1 820
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730589202
transform 1 0 104 0 -1 820
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5796_6
timestamp 1730589202
transform 1 0 128 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5795_6
timestamp 1730589202
transform 1 0 152 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5795_6
timestamp 1730589202
transform 1 0 152 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5796_6
timestamp 1730589202
transform 1 0 128 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5794_6
timestamp 1730589202
transform 1 0 176 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5794_6
timestamp 1730589202
transform 1 0 176 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5793_6
timestamp 1730589202
transform 1 0 208 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5793_6
timestamp 1730589202
transform 1 0 208 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5792_6
timestamp 1730589202
transform 1 0 256 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5792_6
timestamp 1730589202
transform 1 0 256 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5791_6
timestamp 1730589202
transform 1 0 304 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5791_6
timestamp 1730589202
transform 1 0 304 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5790_6
timestamp 1730589202
transform 1 0 360 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5790_6
timestamp 1730589202
transform 1 0 360 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5652_6
timestamp 1730589202
transform 1 0 424 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5652_6
timestamp 1730589202
transform 1 0 424 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5651_6
timestamp 1730589202
transform 1 0 480 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5651_6
timestamp 1730589202
transform 1 0 480 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5650_6
timestamp 1730589202
transform 1 0 536 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5650_6
timestamp 1730589202
transform 1 0 536 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5598_6
timestamp 1730589202
transform 1 0 592 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5598_6
timestamp 1730589202
transform 1 0 592 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5599_6
timestamp 1730589202
transform 1 0 648 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5599_6
timestamp 1730589202
transform 1 0 648 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5597_6
timestamp 1730589202
transform 1 0 704 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5597_6
timestamp 1730589202
transform 1 0 704 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5553_6
timestamp 1730589202
transform 1 0 760 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5553_6
timestamp 1730589202
transform 1 0 760 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5552_6
timestamp 1730589202
transform 1 0 808 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5552_6
timestamp 1730589202
transform 1 0 808 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5456_6
timestamp 1730589202
transform 1 0 856 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5456_6
timestamp 1730589202
transform 1 0 856 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5457_6
timestamp 1730589202
transform 1 0 896 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5457_6
timestamp 1730589202
transform 1 0 896 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5458_6
timestamp 1730589202
transform 1 0 928 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5458_6
timestamp 1730589202
transform 1 0 928 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5460_6
timestamp 1730589202
transform 1 0 984 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5459_6
timestamp 1730589202
transform 1 0 960 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5459_6
timestamp 1730589202
transform 1 0 960 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5460_6
timestamp 1730589202
transform 1 0 984 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5462_6
timestamp 1730589202
transform 1 0 1032 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5461_6
timestamp 1730589202
transform 1 0 1008 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5461_6
timestamp 1730589202
transform 1 0 1008 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5462_6
timestamp 1730589202
transform 1 0 1032 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5463_6
timestamp 1730589202
transform 1 0 1056 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5463_6
timestamp 1730589202
transform 1 0 1056 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5473_6
timestamp 1730589202
transform 1 0 1120 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5464_6
timestamp 1730589202
transform 1 0 1088 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5464_6
timestamp 1730589202
transform 1 0 1088 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5473_6
timestamp 1730589202
transform 1 0 1120 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5474_6
timestamp 1730589202
transform 1 0 1160 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5474_6
timestamp 1730589202
transform 1 0 1160 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5475_6
timestamp 1730589202
transform 1 0 1200 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5475_6
timestamp 1730589202
transform 1 0 1200 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5476_6
timestamp 1730589202
transform 1 0 1248 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5476_6
timestamp 1730589202
transform 1 0 1248 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5477_6
timestamp 1730589202
transform 1 0 1304 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5477_6
timestamp 1730589202
transform 1 0 1304 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5204_6
timestamp 1730589202
transform 1 0 1368 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5204_6
timestamp 1730589202
transform 1 0 1368 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5205_6
timestamp 1730589202
transform 1 0 1408 0 -1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5205_6
timestamp 1730589202
transform 1 0 1408 0 -1 824
box 8 4 20 35
use welltap_svt  __well_tap__35
timestamp 1730589202
transform 1 0 1440 0 -1 820
box 8 4 12 24
use welltap_svt  __well_tap__35
timestamp 1730589202
transform 1 0 1440 0 -1 820
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730589202
transform 1 0 104 0 1 828
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730589202
transform 1 0 104 0 1 828
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5789_6
timestamp 1730589202
transform 1 0 200 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5788_6
timestamp 1730589202
transform 1 0 224 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5783_6
timestamp 1730589202
transform 1 0 224 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5783_6
timestamp 1730589202
transform 1 0 224 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5788_6
timestamp 1730589202
transform 1 0 224 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5789_6
timestamp 1730589202
transform 1 0 200 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5787_6
timestamp 1730589202
transform 1 0 248 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5786_6
timestamp 1730589202
transform 1 0 280 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5782_6
timestamp 1730589202
transform 1 0 248 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5781_6
timestamp 1730589202
transform 1 0 272 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5781_6
timestamp 1730589202
transform 1 0 272 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5782_6
timestamp 1730589202
transform 1 0 248 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5786_6
timestamp 1730589202
transform 1 0 280 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5787_6
timestamp 1730589202
transform 1 0 248 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5785_6
timestamp 1730589202
transform 1 0 312 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5780_6
timestamp 1730589202
transform 1 0 296 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5779_6
timestamp 1730589202
transform 1 0 320 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5779_6
timestamp 1730589202
transform 1 0 320 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5780_6
timestamp 1730589202
transform 1 0 296 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5785_6
timestamp 1730589202
transform 1 0 312 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5784_6
timestamp 1730589202
transform 1 0 344 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5778_6
timestamp 1730589202
transform 1 0 352 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5778_6
timestamp 1730589202
transform 1 0 352 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5784_6
timestamp 1730589202
transform 1 0 344 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5777_6
timestamp 1730589202
transform 1 0 384 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5656_6
timestamp 1730589202
transform 1 0 376 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5656_6
timestamp 1730589202
transform 1 0 376 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5777_6
timestamp 1730589202
transform 1 0 384 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5658_6
timestamp 1730589202
transform 1 0 448 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5657_6
timestamp 1730589202
transform 1 0 416 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5655_6
timestamp 1730589202
transform 1 0 408 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5654_6
timestamp 1730589202
transform 1 0 440 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5654_6
timestamp 1730589202
transform 1 0 440 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5655_6
timestamp 1730589202
transform 1 0 408 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5657_6
timestamp 1730589202
transform 1 0 416 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5658_6
timestamp 1730589202
transform 1 0 448 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5659_6
timestamp 1730589202
transform 1 0 488 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5653_6
timestamp 1730589202
transform 1 0 472 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5653_6
timestamp 1730589202
transform 1 0 472 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5659_6
timestamp 1730589202
transform 1 0 488 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5649_6
timestamp 1730589202
transform 1 0 504 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5645_6
timestamp 1730589202
transform 1 0 528 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5645_6
timestamp 1730589202
transform 1 0 528 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5649_6
timestamp 1730589202
transform 1 0 504 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5648_6
timestamp 1730589202
transform 1 0 544 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5644_6
timestamp 1730589202
transform 1 0 568 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5644_6
timestamp 1730589202
transform 1 0 568 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5648_6
timestamp 1730589202
transform 1 0 544 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5647_6
timestamp 1730589202
transform 1 0 592 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5643_6
timestamp 1730589202
transform 1 0 616 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5643_6
timestamp 1730589202
transform 1 0 616 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5647_6
timestamp 1730589202
transform 1 0 592 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5646_6
timestamp 1730589202
transform 1 0 640 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5642_6
timestamp 1730589202
transform 1 0 656 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5642_6
timestamp 1730589202
transform 1 0 656 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5646_6
timestamp 1730589202
transform 1 0 640 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5602_6
timestamp 1730589202
transform 1 0 696 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5600_6
timestamp 1730589202
transform 1 0 696 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5600_6
timestamp 1730589202
transform 1 0 696 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5602_6
timestamp 1730589202
transform 1 0 696 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5603_6
timestamp 1730589202
transform 1 0 744 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5601_6
timestamp 1730589202
transform 1 0 760 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5601_6
timestamp 1730589202
transform 1 0 760 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5603_6
timestamp 1730589202
transform 1 0 744 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5604_6
timestamp 1730589202
transform 1 0 800 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5604_6
timestamp 1730589202
transform 1 0 800 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5551_6
timestamp 1730589202
transform 1 0 832 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5548_6
timestamp 1730589202
transform 1 0 856 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5548_6
timestamp 1730589202
transform 1 0 856 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5551_6
timestamp 1730589202
transform 1 0 832 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5550_6
timestamp 1730589202
transform 1 0 904 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5550_6
timestamp 1730589202
transform 1 0 904 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5547_6
timestamp 1730589202
transform 1 0 920 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5547_6
timestamp 1730589202
transform 1 0 920 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5549_6
timestamp 1730589202
transform 1 0 976 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5546_6
timestamp 1730589202
transform 1 0 984 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5546_6
timestamp 1730589202
transform 1 0 984 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5549_6
timestamp 1730589202
transform 1 0 976 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5545_6
timestamp 1730589202
transform 1 0 1048 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5478_6
timestamp 1730589202
transform 1 0 1040 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5478_6
timestamp 1730589202
transform 1 0 1040 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5545_6
timestamp 1730589202
transform 1 0 1048 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5485_6
timestamp 1730589202
transform 1 0 1112 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5479_6
timestamp 1730589202
transform 1 0 1096 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5479_6
timestamp 1730589202
transform 1 0 1096 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5485_6
timestamp 1730589202
transform 1 0 1112 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5480_6
timestamp 1730589202
transform 1 0 1152 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5480_6
timestamp 1730589202
transform 1 0 1152 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5486_6
timestamp 1730589202
transform 1 0 1168 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5481_6
timestamp 1730589202
transform 1 0 1200 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5481_6
timestamp 1730589202
transform 1 0 1200 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5486_6
timestamp 1730589202
transform 1 0 1168 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5487_6
timestamp 1730589202
transform 1 0 1224 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5482_6
timestamp 1730589202
transform 1 0 1240 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5482_6
timestamp 1730589202
transform 1 0 1240 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5487_6
timestamp 1730589202
transform 1 0 1224 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5488_6
timestamp 1730589202
transform 1 0 1272 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5483_6
timestamp 1730589202
transform 1 0 1288 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5483_6
timestamp 1730589202
transform 1 0 1288 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5488_6
timestamp 1730589202
transform 1 0 1272 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5489_6
timestamp 1730589202
transform 1 0 1320 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5489_6
timestamp 1730589202
transform 1 0 1320 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5484_6
timestamp 1730589202
transform 1 0 1336 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5484_6
timestamp 1730589202
transform 1 0 1336 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5490_6
timestamp 1730589202
transform 1 0 1376 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5203_6
timestamp 1730589202
transform 1 0 1384 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5202_6
timestamp 1730589202
transform 1 0 1408 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5201_6
timestamp 1730589202
transform 1 0 1408 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5201_6
timestamp 1730589202
transform 1 0 1408 0 -1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5202_6
timestamp 1730589202
transform 1 0 1408 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5203_6
timestamp 1730589202
transform 1 0 1384 0 1 824
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5490_6
timestamp 1730589202
transform 1 0 1376 0 -1 904
box 8 4 20 35
use welltap_svt  __well_tap__37
timestamp 1730589202
transform 1 0 1440 0 1 828
box 8 4 12 24
use welltap_svt  __well_tap__37
timestamp 1730589202
transform 1 0 1440 0 1 828
box 8 4 12 24
use welltap_svt  __well_tap__38
timestamp 1730589202
transform 1 0 104 0 -1 900
box 8 4 12 24
use welltap_svt  __well_tap__38
timestamp 1730589202
transform 1 0 104 0 -1 900
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5771_6
timestamp 1730589202
transform 1 0 232 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5770_6
timestamp 1730589202
transform 1 0 208 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5770_6
timestamp 1730589202
transform 1 0 208 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5771_6
timestamp 1730589202
transform 1 0 232 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5773_6
timestamp 1730589202
transform 1 0 280 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5772_6
timestamp 1730589202
transform 1 0 256 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5772_6
timestamp 1730589202
transform 1 0 256 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5773_6
timestamp 1730589202
transform 1 0 280 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5774_6
timestamp 1730589202
transform 1 0 312 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5774_6
timestamp 1730589202
transform 1 0 312 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5775_6
timestamp 1730589202
transform 1 0 344 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5775_6
timestamp 1730589202
transform 1 0 344 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5776_6
timestamp 1730589202
transform 1 0 384 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5776_6
timestamp 1730589202
transform 1 0 384 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5661_6
timestamp 1730589202
transform 1 0 424 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5661_6
timestamp 1730589202
transform 1 0 424 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5660_6
timestamp 1730589202
transform 1 0 464 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5660_6
timestamp 1730589202
transform 1 0 464 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5662_6
timestamp 1730589202
transform 1 0 512 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5662_6
timestamp 1730589202
transform 1 0 512 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5641_6
timestamp 1730589202
transform 1 0 560 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5641_6
timestamp 1730589202
transform 1 0 560 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5640_6
timestamp 1730589202
transform 1 0 608 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5640_6
timestamp 1730589202
transform 1 0 608 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5639_6
timestamp 1730589202
transform 1 0 664 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5639_6
timestamp 1730589202
transform 1 0 664 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5638_6
timestamp 1730589202
transform 1 0 720 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5638_6
timestamp 1730589202
transform 1 0 720 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5606_6
timestamp 1730589202
transform 1 0 776 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5606_6
timestamp 1730589202
transform 1 0 776 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5605_6
timestamp 1730589202
transform 1 0 840 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5605_6
timestamp 1730589202
transform 1 0 840 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5542_6
timestamp 1730589202
transform 1 0 912 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5542_6
timestamp 1730589202
transform 1 0 912 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5543_6
timestamp 1730589202
transform 1 0 984 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5543_6
timestamp 1730589202
transform 1 0 984 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5544_6
timestamp 1730589202
transform 1 0 1048 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5544_6
timestamp 1730589202
transform 1 0 1048 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5497_6
timestamp 1730589202
transform 1 0 1112 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5497_6
timestamp 1730589202
transform 1 0 1112 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5496_6
timestamp 1730589202
transform 1 0 1168 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5496_6
timestamp 1730589202
transform 1 0 1168 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5495_6
timestamp 1730589202
transform 1 0 1216 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5495_6
timestamp 1730589202
transform 1 0 1216 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5494_6
timestamp 1730589202
transform 1 0 1256 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5493_6
timestamp 1730589202
transform 1 0 1288 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5493_6
timestamp 1730589202
transform 1 0 1288 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5494_6
timestamp 1730589202
transform 1 0 1256 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5492_6
timestamp 1730589202
transform 1 0 1320 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5492_6
timestamp 1730589202
transform 1 0 1320 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5491_6
timestamp 1730589202
transform 1 0 1352 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5491_6
timestamp 1730589202
transform 1 0 1352 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5200_6
timestamp 1730589202
transform 1 0 1384 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5199_6
timestamp 1730589202
transform 1 0 1408 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5199_6
timestamp 1730589202
transform 1 0 1408 0 1 904
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5200_6
timestamp 1730589202
transform 1 0 1384 0 1 904
box 8 4 20 35
use welltap_svt  __well_tap__39
timestamp 1730589202
transform 1 0 1440 0 -1 900
box 8 4 12 24
use welltap_svt  __well_tap__39
timestamp 1730589202
transform 1 0 1440 0 -1 900
box 8 4 12 24
use welltap_svt  __well_tap__40
timestamp 1730589202
transform 1 0 104 0 1 908
box 8 4 12 24
use welltap_svt  __well_tap__40
timestamp 1730589202
transform 1 0 104 0 1 908
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5765_6
timestamp 1730589202
transform 1 0 224 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5764_6
timestamp 1730589202
transform 1 0 200 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5764_6
timestamp 1730589202
transform 1 0 200 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5765_6
timestamp 1730589202
transform 1 0 224 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5767_6
timestamp 1730589202
transform 1 0 280 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5766_6
timestamp 1730589202
transform 1 0 248 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5766_6
timestamp 1730589202
transform 1 0 248 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5767_6
timestamp 1730589202
transform 1 0 280 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5768_6
timestamp 1730589202
transform 1 0 320 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5768_6
timestamp 1730589202
transform 1 0 320 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5769_6
timestamp 1730589202
transform 1 0 368 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5769_6
timestamp 1730589202
transform 1 0 368 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5665_6
timestamp 1730589202
transform 1 0 416 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5665_6
timestamp 1730589202
transform 1 0 416 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5664_6
timestamp 1730589202
transform 1 0 464 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5664_6
timestamp 1730589202
transform 1 0 464 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5663_6
timestamp 1730589202
transform 1 0 512 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5663_6
timestamp 1730589202
transform 1 0 512 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5637_6
timestamp 1730589202
transform 1 0 560 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5637_6
timestamp 1730589202
transform 1 0 560 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5636_6
timestamp 1730589202
transform 1 0 616 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5636_6
timestamp 1730589202
transform 1 0 616 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5635_6
timestamp 1730589202
transform 1 0 672 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5635_6
timestamp 1730589202
transform 1 0 672 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5634_6
timestamp 1730589202
transform 1 0 720 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5634_6
timestamp 1730589202
transform 1 0 720 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5607_6
timestamp 1730589202
transform 1 0 768 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5607_6
timestamp 1730589202
transform 1 0 768 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5608_6
timestamp 1730589202
transform 1 0 824 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5608_6
timestamp 1730589202
transform 1 0 824 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5609_6
timestamp 1730589202
transform 1 0 880 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5609_6
timestamp 1730589202
transform 1 0 880 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5541_6
timestamp 1730589202
transform 1 0 936 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5541_6
timestamp 1730589202
transform 1 0 936 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5540_6
timestamp 1730589202
transform 1 0 992 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5540_6
timestamp 1730589202
transform 1 0 992 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5539_6
timestamp 1730589202
transform 1 0 1040 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5539_6
timestamp 1730589202
transform 1 0 1040 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5538_6
timestamp 1730589202
transform 1 0 1088 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5538_6
timestamp 1730589202
transform 1 0 1088 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5503_6
timestamp 1730589202
transform 1 0 1136 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5503_6
timestamp 1730589202
transform 1 0 1136 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5502_6
timestamp 1730589202
transform 1 0 1184 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5502_6
timestamp 1730589202
transform 1 0 1184 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5501_6
timestamp 1730589202
transform 1 0 1232 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5501_6
timestamp 1730589202
transform 1 0 1232 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5500_6
timestamp 1730589202
transform 1 0 1280 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5500_6
timestamp 1730589202
transform 1 0 1280 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5499_6
timestamp 1730589202
transform 1 0 1328 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5499_6
timestamp 1730589202
transform 1 0 1328 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5498_6
timestamp 1730589202
transform 1 0 1376 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5198_6
timestamp 1730589202
transform 1 0 1408 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5198_6
timestamp 1730589202
transform 1 0 1408 0 -1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5498_6
timestamp 1730589202
transform 1 0 1376 0 -1 984
box 8 4 20 35
use welltap_svt  __well_tap__41
timestamp 1730589202
transform 1 0 1440 0 1 908
box 8 4 12 24
use welltap_svt  __well_tap__41
timestamp 1730589202
transform 1 0 1440 0 1 908
box 8 4 12 24
use welltap_svt  __well_tap__44
timestamp 1730589202
transform 1 0 104 0 1 988
box 8 4 12 24
use welltap_svt  __well_tap__42
timestamp 1730589202
transform 1 0 104 0 -1 980
box 8 4 12 24
use welltap_svt  __well_tap__42
timestamp 1730589202
transform 1 0 104 0 -1 980
box 8 4 12 24
use welltap_svt  __well_tap__44
timestamp 1730589202
transform 1 0 104 0 1 988
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5757_6
timestamp 1730589202
transform 1 0 152 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5757_6
timestamp 1730589202
transform 1 0 152 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5758_6
timestamp 1730589202
transform 1 0 176 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5758_6
timestamp 1730589202
transform 1 0 176 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5760_6
timestamp 1730589202
transform 1 0 224 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5759_6
timestamp 1730589202
transform 1 0 200 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5759_6
timestamp 1730589202
transform 1 0 200 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5760_6
timestamp 1730589202
transform 1 0 224 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5761_6
timestamp 1730589202
transform 1 0 256 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5761_6
timestamp 1730589202
transform 1 0 256 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5762_6
timestamp 1730589202
transform 1 0 296 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5762_6
timestamp 1730589202
transform 1 0 296 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5763_6
timestamp 1730589202
transform 1 0 336 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5763_6
timestamp 1730589202
transform 1 0 336 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5666_6
timestamp 1730589202
transform 1 0 376 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5666_6
timestamp 1730589202
transform 1 0 376 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5667_6
timestamp 1730589202
transform 1 0 424 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5667_6
timestamp 1730589202
transform 1 0 424 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5668_6
timestamp 1730589202
transform 1 0 472 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5668_6
timestamp 1730589202
transform 1 0 472 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5669_6
timestamp 1730589202
transform 1 0 520 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5669_6
timestamp 1730589202
transform 1 0 520 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5670_6
timestamp 1730589202
transform 1 0 568 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5670_6
timestamp 1730589202
transform 1 0 568 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5633_6
timestamp 1730589202
transform 1 0 616 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5633_6
timestamp 1730589202
transform 1 0 616 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5632_6
timestamp 1730589202
transform 1 0 664 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5632_6
timestamp 1730589202
transform 1 0 664 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5631_6
timestamp 1730589202
transform 1 0 712 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5631_6
timestamp 1730589202
transform 1 0 712 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5630_6
timestamp 1730589202
transform 1 0 760 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5630_6
timestamp 1730589202
transform 1 0 760 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5612_6
timestamp 1730589202
transform 1 0 816 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5612_6
timestamp 1730589202
transform 1 0 816 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5611_6
timestamp 1730589202
transform 1 0 872 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5611_6
timestamp 1730589202
transform 1 0 872 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5610_6
timestamp 1730589202
transform 1 0 928 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5610_6
timestamp 1730589202
transform 1 0 928 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5535_6
timestamp 1730589202
transform 1 0 984 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5535_6
timestamp 1730589202
transform 1 0 984 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5536_6
timestamp 1730589202
transform 1 0 1040 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5536_6
timestamp 1730589202
transform 1 0 1040 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5537_6
timestamp 1730589202
transform 1 0 1096 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5537_6
timestamp 1730589202
transform 1 0 1096 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5507_6
timestamp 1730589202
transform 1 0 1152 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5507_6
timestamp 1730589202
transform 1 0 1152 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5506_6
timestamp 1730589202
transform 1 0 1208 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5506_6
timestamp 1730589202
transform 1 0 1208 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5505_6
timestamp 1730589202
transform 1 0 1264 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5505_6
timestamp 1730589202
transform 1 0 1264 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5504_6
timestamp 1730589202
transform 1 0 1320 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5504_6
timestamp 1730589202
transform 1 0 1320 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5197_6
timestamp 1730589202
transform 1 0 1408 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5196_6
timestamp 1730589202
transform 1 0 1376 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5196_6
timestamp 1730589202
transform 1 0 1376 0 1 984
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5197_6
timestamp 1730589202
transform 1 0 1408 0 1 984
box 8 4 20 35
use welltap_svt  __well_tap__45
timestamp 1730589202
transform 1 0 1440 0 1 988
box 8 4 12 24
use welltap_svt  __well_tap__43
timestamp 1730589202
transform 1 0 1440 0 -1 980
box 8 4 12 24
use welltap_svt  __well_tap__43
timestamp 1730589202
transform 1 0 1440 0 -1 980
box 8 4 12 24
use welltap_svt  __well_tap__45
timestamp 1730589202
transform 1 0 1440 0 1 988
box 8 4 12 24
use welltap_svt  __well_tap__46
timestamp 1730589202
transform 1 0 104 0 -1 1060
box 8 4 12 24
use welltap_svt  __well_tap__46
timestamp 1730589202
transform 1 0 104 0 -1 1060
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5751_6
timestamp 1730589202
transform 1 0 152 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5750_6
timestamp 1730589202
transform 1 0 128 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5750_6
timestamp 1730589202
transform 1 0 128 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5751_6
timestamp 1730589202
transform 1 0 152 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5752_6
timestamp 1730589202
transform 1 0 176 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5752_6
timestamp 1730589202
transform 1 0 176 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5754_6
timestamp 1730589202
transform 1 0 224 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5753_6
timestamp 1730589202
transform 1 0 200 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5753_6
timestamp 1730589202
transform 1 0 200 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5754_6
timestamp 1730589202
transform 1 0 224 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5755_6
timestamp 1730589202
transform 1 0 264 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5755_6
timestamp 1730589202
transform 1 0 264 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5756_6
timestamp 1730589202
transform 1 0 304 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5756_6
timestamp 1730589202
transform 1 0 304 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5677_6
timestamp 1730589202
transform 1 0 344 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5677_6
timestamp 1730589202
transform 1 0 344 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5676_6
timestamp 1730589202
transform 1 0 384 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5676_6
timestamp 1730589202
transform 1 0 384 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5675_6
timestamp 1730589202
transform 1 0 424 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5675_6
timestamp 1730589202
transform 1 0 424 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5674_6
timestamp 1730589202
transform 1 0 464 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5674_6
timestamp 1730589202
transform 1 0 464 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5673_6
timestamp 1730589202
transform 1 0 504 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5673_6
timestamp 1730589202
transform 1 0 504 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5672_6
timestamp 1730589202
transform 1 0 544 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5672_6
timestamp 1730589202
transform 1 0 544 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5671_6
timestamp 1730589202
transform 1 0 584 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5671_6
timestamp 1730589202
transform 1 0 584 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5629_6
timestamp 1730589202
transform 1 0 624 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5629_6
timestamp 1730589202
transform 1 0 624 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5628_6
timestamp 1730589202
transform 1 0 664 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5628_6
timestamp 1730589202
transform 1 0 664 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5627_6
timestamp 1730589202
transform 1 0 704 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5626_6
timestamp 1730589202
transform 1 0 736 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5626_6
timestamp 1730589202
transform 1 0 736 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5627_6
timestamp 1730589202
transform 1 0 704 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5625_6
timestamp 1730589202
transform 1 0 776 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5625_6
timestamp 1730589202
transform 1 0 776 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5613_6
timestamp 1730589202
transform 1 0 816 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5613_6
timestamp 1730589202
transform 1 0 816 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5614_6
timestamp 1730589202
transform 1 0 864 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5614_6
timestamp 1730589202
transform 1 0 864 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5615_6
timestamp 1730589202
transform 1 0 912 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5615_6
timestamp 1730589202
transform 1 0 912 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5616_6
timestamp 1730589202
transform 1 0 968 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5616_6
timestamp 1730589202
transform 1 0 968 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5534_6
timestamp 1730589202
transform 1 0 1024 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5534_6
timestamp 1730589202
transform 1 0 1024 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5533_6
timestamp 1730589202
transform 1 0 1072 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5533_6
timestamp 1730589202
transform 1 0 1072 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5532_6
timestamp 1730589202
transform 1 0 1120 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5532_6
timestamp 1730589202
transform 1 0 1120 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5508_6
timestamp 1730589202
transform 1 0 1168 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5508_6
timestamp 1730589202
transform 1 0 1168 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5509_6
timestamp 1730589202
transform 1 0 1216 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5509_6
timestamp 1730589202
transform 1 0 1216 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5510_6
timestamp 1730589202
transform 1 0 1264 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5510_6
timestamp 1730589202
transform 1 0 1264 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5511_6
timestamp 1730589202
transform 1 0 1320 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5511_6
timestamp 1730589202
transform 1 0 1320 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5195_6
timestamp 1730589202
transform 1 0 1376 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5194_6
timestamp 1730589202
transform 1 0 1408 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5194_6
timestamp 1730589202
transform 1 0 1408 0 -1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5195_6
timestamp 1730589202
transform 1 0 1376 0 -1 1064
box 8 4 20 35
use welltap_svt  __well_tap__47
timestamp 1730589202
transform 1 0 1440 0 -1 1060
box 8 4 12 24
use welltap_svt  __well_tap__47
timestamp 1730589202
transform 1 0 1440 0 -1 1060
box 8 4 12 24
use welltap_svt  __well_tap__48
timestamp 1730589202
transform 1 0 104 0 1 1068
box 8 4 12 24
use welltap_svt  __well_tap__48
timestamp 1730589202
transform 1 0 104 0 1 1068
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5746_6
timestamp 1730589202
transform 1 0 128 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5745_6
timestamp 1730589202
transform 1 0 152 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5745_6
timestamp 1730589202
transform 1 0 152 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5746_6
timestamp 1730589202
transform 1 0 128 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5744_6
timestamp 1730589202
transform 1 0 176 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5744_6
timestamp 1730589202
transform 1 0 176 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5747_6
timestamp 1730589202
transform 1 0 200 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5747_6
timestamp 1730589202
transform 1 0 200 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5749_6
timestamp 1730589202
transform 1 0 280 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5748_6
timestamp 1730589202
transform 1 0 240 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5748_6
timestamp 1730589202
transform 1 0 240 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5749_6
timestamp 1730589202
transform 1 0 280 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5683_6
timestamp 1730589202
transform 1 0 320 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5683_6
timestamp 1730589202
transform 1 0 320 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5684_6
timestamp 1730589202
transform 1 0 360 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5684_6
timestamp 1730589202
transform 1 0 360 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5682_6
timestamp 1730589202
transform 1 0 400 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5682_6
timestamp 1730589202
transform 1 0 400 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5681_6
timestamp 1730589202
transform 1 0 448 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5681_6
timestamp 1730589202
transform 1 0 448 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5680_6
timestamp 1730589202
transform 1 0 496 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5680_6
timestamp 1730589202
transform 1 0 496 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5679_6
timestamp 1730589202
transform 1 0 552 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5679_6
timestamp 1730589202
transform 1 0 552 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5678_6
timestamp 1730589202
transform 1 0 600 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5678_6
timestamp 1730589202
transform 1 0 600 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5624_6
timestamp 1730589202
transform 1 0 648 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5624_6
timestamp 1730589202
transform 1 0 648 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5623_6
timestamp 1730589202
transform 1 0 696 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5623_6
timestamp 1730589202
transform 1 0 696 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5622_6
timestamp 1730589202
transform 1 0 736 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5622_6
timestamp 1730589202
transform 1 0 736 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5621_6
timestamp 1730589202
transform 1 0 784 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5621_6
timestamp 1730589202
transform 1 0 784 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5620_6
timestamp 1730589202
transform 1 0 832 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5620_6
timestamp 1730589202
transform 1 0 832 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5619_6
timestamp 1730589202
transform 1 0 880 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5619_6
timestamp 1730589202
transform 1 0 880 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5618_6
timestamp 1730589202
transform 1 0 936 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5618_6
timestamp 1730589202
transform 1 0 936 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5617_6
timestamp 1730589202
transform 1 0 992 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5617_6
timestamp 1730589202
transform 1 0 992 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5529_6
timestamp 1730589202
transform 1 0 1048 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5529_6
timestamp 1730589202
transform 1 0 1048 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5530_6
timestamp 1730589202
transform 1 0 1104 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5530_6
timestamp 1730589202
transform 1 0 1104 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5531_6
timestamp 1730589202
transform 1 0 1160 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5531_6
timestamp 1730589202
transform 1 0 1160 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5512_6
timestamp 1730589202
transform 1 0 1208 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5512_6
timestamp 1730589202
transform 1 0 1208 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5513_6
timestamp 1730589202
transform 1 0 1264 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5513_6
timestamp 1730589202
transform 1 0 1264 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5514_6
timestamp 1730589202
transform 1 0 1320 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5514_6
timestamp 1730589202
transform 1 0 1320 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5515_6
timestamp 1730589202
transform 1 0 1376 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5193_6
timestamp 1730589202
transform 1 0 1408 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5193_6
timestamp 1730589202
transform 1 0 1408 0 1 1064
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5515_6
timestamp 1730589202
transform 1 0 1376 0 1 1064
box 8 4 20 35
use welltap_svt  __well_tap__49
timestamp 1730589202
transform 1 0 1440 0 1 1068
box 8 4 12 24
use welltap_svt  __well_tap__49
timestamp 1730589202
transform 1 0 1440 0 1 1068
box 8 4 12 24
use welltap_svt  __well_tap__50
timestamp 1730589202
transform 1 0 104 0 -1 1144
box 8 4 12 24
use welltap_svt  __well_tap__50
timestamp 1730589202
transform 1 0 104 0 -1 1144
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5742_6
timestamp 1730589202
transform 1 0 152 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5741_6
timestamp 1730589202
transform 1 0 128 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5741_6
timestamp 1730589202
transform 1 0 128 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5742_6
timestamp 1730589202
transform 1 0 152 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5743_6
timestamp 1730589202
transform 1 0 176 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5743_6
timestamp 1730589202
transform 1 0 176 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5732_6
timestamp 1730589202
transform 1 0 208 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5732_6
timestamp 1730589202
transform 1 0 208 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5731_6
timestamp 1730589202
transform 1 0 248 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5731_6
timestamp 1730589202
transform 1 0 248 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5730_6
timestamp 1730589202
transform 1 0 288 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5730_6
timestamp 1730589202
transform 1 0 288 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5729_6
timestamp 1730589202
transform 1 0 328 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5729_6
timestamp 1730589202
transform 1 0 328 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5685_6
timestamp 1730589202
transform 1 0 368 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5685_6
timestamp 1730589202
transform 1 0 368 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5686_6
timestamp 1730589202
transform 1 0 408 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5686_6
timestamp 1730589202
transform 1 0 408 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5687_6
timestamp 1730589202
transform 1 0 456 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5687_6
timestamp 1730589202
transform 1 0 456 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5688_6
timestamp 1730589202
transform 1 0 512 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5688_6
timestamp 1730589202
transform 1 0 512 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5689_6
timestamp 1730589202
transform 1 0 576 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5689_6
timestamp 1730589202
transform 1 0 576 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5690_6
timestamp 1730589202
transform 1 0 640 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5690_6
timestamp 1730589202
transform 1 0 640 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5691_6
timestamp 1730589202
transform 1 0 704 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5691_6
timestamp 1730589202
transform 1 0 704 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5121_6
timestamp 1730589202
transform 1 0 760 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5121_6
timestamp 1730589202
transform 1 0 760 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5122_6
timestamp 1730589202
transform 1 0 824 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5122_6
timestamp 1730589202
transform 1 0 824 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5123_6
timestamp 1730589202
transform 1 0 880 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5123_6
timestamp 1730589202
transform 1 0 880 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5124_6
timestamp 1730589202
transform 1 0 936 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5124_6
timestamp 1730589202
transform 1 0 936 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5125_6
timestamp 1730589202
transform 1 0 992 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5125_6
timestamp 1730589202
transform 1 0 992 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5126_6
timestamp 1730589202
transform 1 0 1048 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5126_6
timestamp 1730589202
transform 1 0 1048 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5528_6
timestamp 1730589202
transform 1 0 1096 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5528_6
timestamp 1730589202
transform 1 0 1096 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5527_6
timestamp 1730589202
transform 1 0 1144 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5527_6
timestamp 1730589202
transform 1 0 1144 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5526_6
timestamp 1730589202
transform 1 0 1184 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5526_6
timestamp 1730589202
transform 1 0 1184 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5525_6
timestamp 1730589202
transform 1 0 1224 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5525_6
timestamp 1730589202
transform 1 0 1224 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5518_6
timestamp 1730589202
transform 1 0 1264 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5518_6
timestamp 1730589202
transform 1 0 1264 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5517_6
timestamp 1730589202
transform 1 0 1304 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5517_6
timestamp 1730589202
transform 1 0 1304 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5516_6
timestamp 1730589202
transform 1 0 1344 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5516_6
timestamp 1730589202
transform 1 0 1344 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5192_6
timestamp 1730589202
transform 1 0 1408 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5191_6
timestamp 1730589202
transform 1 0 1384 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5191_6
timestamp 1730589202
transform 1 0 1384 0 -1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5192_6
timestamp 1730589202
transform 1 0 1408 0 -1 1148
box 8 4 20 35
use welltap_svt  __well_tap__51
timestamp 1730589202
transform 1 0 1440 0 -1 1144
box 8 4 12 24
use welltap_svt  __well_tap__51
timestamp 1730589202
transform 1 0 1440 0 -1 1144
box 8 4 12 24
use welltap_svt  __well_tap__52
timestamp 1730589202
transform 1 0 104 0 1 1152
box 8 4 12 24
use welltap_svt  __well_tap__52
timestamp 1730589202
transform 1 0 104 0 1 1152
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5740_6
timestamp 1730589202
transform 1 0 128 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5739_6
timestamp 1730589202
transform 1 0 152 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5739_6
timestamp 1730589202
transform 1 0 152 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5740_6
timestamp 1730589202
transform 1 0 128 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5738_6
timestamp 1730589202
transform 1 0 176 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5738_6
timestamp 1730589202
transform 1 0 176 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5737_6
timestamp 1730589202
transform 1 0 200 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5736_6
timestamp 1730589202
transform 1 0 224 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5736_6
timestamp 1730589202
transform 1 0 224 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5737_6
timestamp 1730589202
transform 1 0 200 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5735_6
timestamp 1730589202
transform 1 0 248 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5734_6
timestamp 1730589202
transform 1 0 272 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5734_6
timestamp 1730589202
transform 1 0 272 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5735_6
timestamp 1730589202
transform 1 0 248 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5733_6
timestamp 1730589202
transform 1 0 296 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5733_6
timestamp 1730589202
transform 1 0 296 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5726_6
timestamp 1730589202
transform 1 0 328 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5726_6
timestamp 1730589202
transform 1 0 328 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5727_6
timestamp 1730589202
transform 1 0 376 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5727_6
timestamp 1730589202
transform 1 0 376 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5728_6
timestamp 1730589202
transform 1 0 416 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5728_6
timestamp 1730589202
transform 1 0 416 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5692_6
timestamp 1730589202
transform 1 0 456 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5692_6
timestamp 1730589202
transform 1 0 456 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5693_6
timestamp 1730589202
transform 1 0 496 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5693_6
timestamp 1730589202
transform 1 0 496 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5694_6
timestamp 1730589202
transform 1 0 536 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5694_6
timestamp 1730589202
transform 1 0 536 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5696_6
timestamp 1730589202
transform 1 0 616 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5695_6
timestamp 1730589202
transform 1 0 576 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5695_6
timestamp 1730589202
transform 1 0 576 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5696_6
timestamp 1730589202
transform 1 0 616 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5697_6
timestamp 1730589202
transform 1 0 664 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5697_6
timestamp 1730589202
transform 1 0 664 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5698_6
timestamp 1730589202
transform 1 0 712 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5698_6
timestamp 1730589202
transform 1 0 712 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5699_6
timestamp 1730589202
transform 1 0 760 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5699_6
timestamp 1730589202
transform 1 0 760 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5120_6
timestamp 1730589202
transform 1 0 808 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5120_6
timestamp 1730589202
transform 1 0 808 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5119_6
timestamp 1730589202
transform 1 0 856 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5119_6
timestamp 1730589202
transform 1 0 856 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5118_6
timestamp 1730589202
transform 1 0 904 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5118_6
timestamp 1730589202
transform 1 0 904 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5127_6
timestamp 1730589202
transform 1 0 952 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5127_6
timestamp 1730589202
transform 1 0 952 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5128_6
timestamp 1730589202
transform 1 0 1000 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5128_6
timestamp 1730589202
transform 1 0 1000 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5129_6
timestamp 1730589202
transform 1 0 1048 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5129_6
timestamp 1730589202
transform 1 0 1048 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5130_6
timestamp 1730589202
transform 1 0 1096 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5130_6
timestamp 1730589202
transform 1 0 1096 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5524_6
timestamp 1730589202
transform 1 0 1144 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5524_6
timestamp 1730589202
transform 1 0 1144 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5523_6
timestamp 1730589202
transform 1 0 1184 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5523_6
timestamp 1730589202
transform 1 0 1184 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5522_6
timestamp 1730589202
transform 1 0 1224 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5522_6
timestamp 1730589202
transform 1 0 1224 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5521_6
timestamp 1730589202
transform 1 0 1264 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5521_6
timestamp 1730589202
transform 1 0 1264 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5520_6
timestamp 1730589202
transform 1 0 1304 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5520_6
timestamp 1730589202
transform 1 0 1304 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5519_6
timestamp 1730589202
transform 1 0 1344 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5519_6
timestamp 1730589202
transform 1 0 1344 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5190_6
timestamp 1730589202
transform 1 0 1384 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5189_6
timestamp 1730589202
transform 1 0 1408 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5189_6
timestamp 1730589202
transform 1 0 1408 0 1 1148
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5190_6
timestamp 1730589202
transform 1 0 1384 0 1 1148
box 8 4 20 35
use welltap_svt  __well_tap__53
timestamp 1730589202
transform 1 0 1440 0 1 1152
box 8 4 12 24
use welltap_svt  __well_tap__53
timestamp 1730589202
transform 1 0 1440 0 1 1152
box 8 4 12 24
use welltap_svt  __well_tap__54
timestamp 1730589202
transform 1 0 104 0 -1 1224
box 8 4 12 24
use welltap_svt  __well_tap__54
timestamp 1730589202
transform 1 0 104 0 -1 1224
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_5725_6
timestamp 1730589202
transform 1 0 320 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5725_6
timestamp 1730589202
transform 1 0 320 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5724_6
timestamp 1730589202
transform 1 0 360 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5724_6
timestamp 1730589202
transform 1 0 360 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5723_6
timestamp 1730589202
transform 1 0 400 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5723_6
timestamp 1730589202
transform 1 0 400 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5722_6
timestamp 1730589202
transform 1 0 440 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5722_6
timestamp 1730589202
transform 1 0 440 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5705_6
timestamp 1730589202
transform 1 0 480 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5705_6
timestamp 1730589202
transform 1 0 480 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5704_6
timestamp 1730589202
transform 1 0 520 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5704_6
timestamp 1730589202
transform 1 0 520 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5703_6
timestamp 1730589202
transform 1 0 560 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5703_6
timestamp 1730589202
transform 1 0 560 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5702_6
timestamp 1730589202
transform 1 0 600 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5702_6
timestamp 1730589202
transform 1 0 600 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5701_6
timestamp 1730589202
transform 1 0 648 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5701_6
timestamp 1730589202
transform 1 0 648 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5700_6
timestamp 1730589202
transform 1 0 696 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5700_6
timestamp 1730589202
transform 1 0 696 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5114_6
timestamp 1730589202
transform 1 0 744 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5114_6
timestamp 1730589202
transform 1 0 744 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5115_6
timestamp 1730589202
transform 1 0 792 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5115_6
timestamp 1730589202
transform 1 0 792 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5116_6
timestamp 1730589202
transform 1 0 840 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5116_6
timestamp 1730589202
transform 1 0 840 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5117_6
timestamp 1730589202
transform 1 0 888 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5117_6
timestamp 1730589202
transform 1 0 888 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5131_6
timestamp 1730589202
transform 1 0 936 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5131_6
timestamp 1730589202
transform 1 0 936 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5132_6
timestamp 1730589202
transform 1 0 984 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5132_6
timestamp 1730589202
transform 1 0 984 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5133_6
timestamp 1730589202
transform 1 0 1032 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5133_6
timestamp 1730589202
transform 1 0 1032 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5134_6
timestamp 1730589202
transform 1 0 1096 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5134_6
timestamp 1730589202
transform 1 0 1096 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5135_6
timestamp 1730589202
transform 1 0 1168 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5135_6
timestamp 1730589202
transform 1 0 1168 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5136_6
timestamp 1730589202
transform 1 0 1248 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5136_6
timestamp 1730589202
transform 1 0 1248 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5137_6
timestamp 1730589202
transform 1 0 1336 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5137_6
timestamp 1730589202
transform 1 0 1336 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5188_6
timestamp 1730589202
transform 1 0 1408 0 -1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5188_6
timestamp 1730589202
transform 1 0 1408 0 -1 1228
box 8 4 20 35
use welltap_svt  __well_tap__55
timestamp 1730589202
transform 1 0 1440 0 -1 1224
box 8 4 12 24
use welltap_svt  __well_tap__55
timestamp 1730589202
transform 1 0 1440 0 -1 1224
box 8 4 12 24
use welltap_svt  __well_tap__56
timestamp 1730589202
transform 1 0 104 0 1 1232
box 8 4 12 24
use welltap_svt  __well_tap__56
timestamp 1730589202
transform 1 0 104 0 1 1232
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_590_6
timestamp 1730589202
transform 1 0 304 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_590_6
timestamp 1730589202
transform 1 0 304 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_592_6
timestamp 1730589202
transform 1 0 352 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_591_6
timestamp 1730589202
transform 1 0 328 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_591_6
timestamp 1730589202
transform 1 0 328 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_592_6
timestamp 1730589202
transform 1 0 352 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5721_6
timestamp 1730589202
transform 1 0 376 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5721_6
timestamp 1730589202
transform 1 0 376 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5720_6
timestamp 1730589202
transform 1 0 408 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5719_6
timestamp 1730589202
transform 1 0 440 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5719_6
timestamp 1730589202
transform 1 0 440 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5720_6
timestamp 1730589202
transform 1 0 408 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5718_6
timestamp 1730589202
transform 1 0 472 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5718_6
timestamp 1730589202
transform 1 0 472 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5709_6
timestamp 1730589202
transform 1 0 512 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5709_6
timestamp 1730589202
transform 1 0 512 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5708_6
timestamp 1730589202
transform 1 0 552 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5708_6
timestamp 1730589202
transform 1 0 552 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5707_6
timestamp 1730589202
transform 1 0 608 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5707_6
timestamp 1730589202
transform 1 0 608 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5706_6
timestamp 1730589202
transform 1 0 672 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5706_6
timestamp 1730589202
transform 1 0 672 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5113_6
timestamp 1730589202
transform 1 0 744 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5113_6
timestamp 1730589202
transform 1 0 744 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5112_6
timestamp 1730589202
transform 1 0 824 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5112_6
timestamp 1730589202
transform 1 0 824 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5111_6
timestamp 1730589202
transform 1 0 904 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5111_6
timestamp 1730589202
transform 1 0 904 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5139_6
timestamp 1730589202
transform 1 0 984 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5139_6
timestamp 1730589202
transform 1 0 984 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5138_6
timestamp 1730589202
transform 1 0 1056 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5138_6
timestamp 1730589202
transform 1 0 1056 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5167_6
timestamp 1730589202
transform 1 0 1120 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5167_6
timestamp 1730589202
transform 1 0 1120 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5168_6
timestamp 1730589202
transform 1 0 1184 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5168_6
timestamp 1730589202
transform 1 0 1184 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5169_6
timestamp 1730589202
transform 1 0 1240 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5169_6
timestamp 1730589202
transform 1 0 1240 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5170_6
timestamp 1730589202
transform 1 0 1304 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5170_6
timestamp 1730589202
transform 1 0 1304 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5186_6
timestamp 1730589202
transform 1 0 1368 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5186_6
timestamp 1730589202
transform 1 0 1368 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5187_6
timestamp 1730589202
transform 1 0 1408 0 1 1228
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5187_6
timestamp 1730589202
transform 1 0 1408 0 1 1228
box 8 4 20 35
use welltap_svt  __well_tap__57
timestamp 1730589202
transform 1 0 1440 0 1 1232
box 8 4 12 24
use welltap_svt  __well_tap__57
timestamp 1730589202
transform 1 0 1440 0 1 1232
box 8 4 12 24
use welltap_svt  __well_tap__58
timestamp 1730589202
transform 1 0 104 0 -1 1304
box 8 4 12 24
use welltap_svt  __well_tap__58
timestamp 1730589202
transform 1 0 104 0 -1 1304
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_585_6
timestamp 1730589202
transform 1 0 224 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_585_6
timestamp 1730589202
transform 1 0 224 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_587_6
timestamp 1730589202
transform 1 0 272 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_586_6
timestamp 1730589202
transform 1 0 248 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_586_6
timestamp 1730589202
transform 1 0 248 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_587_6
timestamp 1730589202
transform 1 0 272 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_589_6
timestamp 1730589202
transform 1 0 320 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_588_6
timestamp 1730589202
transform 1 0 296 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_588_6
timestamp 1730589202
transform 1 0 296 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_589_6
timestamp 1730589202
transform 1 0 320 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_593_6
timestamp 1730589202
transform 1 0 344 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_593_6
timestamp 1730589202
transform 1 0 344 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5717_6
timestamp 1730589202
transform 1 0 392 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_594_6
timestamp 1730589202
transform 1 0 368 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_594_6
timestamp 1730589202
transform 1 0 368 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5717_6
timestamp 1730589202
transform 1 0 392 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5716_6
timestamp 1730589202
transform 1 0 416 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5715_6
timestamp 1730589202
transform 1 0 440 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5715_6
timestamp 1730589202
transform 1 0 440 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5716_6
timestamp 1730589202
transform 1 0 416 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5714_6
timestamp 1730589202
transform 1 0 464 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5714_6
timestamp 1730589202
transform 1 0 464 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5713_6
timestamp 1730589202
transform 1 0 496 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5713_6
timestamp 1730589202
transform 1 0 496 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5712_6
timestamp 1730589202
transform 1 0 536 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5712_6
timestamp 1730589202
transform 1 0 536 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5711_6
timestamp 1730589202
transform 1 0 584 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5711_6
timestamp 1730589202
transform 1 0 584 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5710_6
timestamp 1730589202
transform 1 0 640 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5710_6
timestamp 1730589202
transform 1 0 640 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5109_6
timestamp 1730589202
transform 1 0 688 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5109_6
timestamp 1730589202
transform 1 0 688 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5110_6
timestamp 1730589202
transform 1 0 736 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5110_6
timestamp 1730589202
transform 1 0 736 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_524_6
timestamp 1730589202
transform 1 0 784 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_524_6
timestamp 1730589202
transform 1 0 784 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_523_6
timestamp 1730589202
transform 1 0 832 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_523_6
timestamp 1730589202
transform 1 0 832 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_522_6
timestamp 1730589202
transform 1 0 872 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_521_6
timestamp 1730589202
transform 1 0 904 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_521_6
timestamp 1730589202
transform 1 0 904 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_522_6
timestamp 1730589202
transform 1 0 872 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_520_6
timestamp 1730589202
transform 1 0 944 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_520_6
timestamp 1730589202
transform 1 0 944 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_519_6
timestamp 1730589202
transform 1 0 984 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_519_6
timestamp 1730589202
transform 1 0 984 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_518_6
timestamp 1730589202
transform 1 0 1024 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_518_6
timestamp 1730589202
transform 1 0 1024 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_517_6
timestamp 1730589202
transform 1 0 1064 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_517_6
timestamp 1730589202
transform 1 0 1064 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5140_6
timestamp 1730589202
transform 1 0 1104 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5140_6
timestamp 1730589202
transform 1 0 1104 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5166_6
timestamp 1730589202
transform 1 0 1144 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5166_6
timestamp 1730589202
transform 1 0 1144 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5165_6
timestamp 1730589202
transform 1 0 1192 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5165_6
timestamp 1730589202
transform 1 0 1192 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5164_6
timestamp 1730589202
transform 1 0 1240 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5164_6
timestamp 1730589202
transform 1 0 1240 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5172_6
timestamp 1730589202
transform 1 0 1296 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5172_6
timestamp 1730589202
transform 1 0 1296 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5171_6
timestamp 1730589202
transform 1 0 1360 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5171_6
timestamp 1730589202
transform 1 0 1360 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5185_6
timestamp 1730589202
transform 1 0 1408 0 -1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5185_6
timestamp 1730589202
transform 1 0 1408 0 -1 1308
box 8 4 20 35
use welltap_svt  __well_tap__59
timestamp 1730589202
transform 1 0 1440 0 -1 1304
box 8 4 12 24
use welltap_svt  __well_tap__59
timestamp 1730589202
transform 1 0 1440 0 -1 1304
box 8 4 12 24
use welltap_svt  __well_tap__60
timestamp 1730589202
transform 1 0 104 0 1 1312
box 8 4 12 24
use welltap_svt  __well_tap__60
timestamp 1730589202
transform 1 0 104 0 1 1312
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_581_6
timestamp 1730589202
transform 1 0 184 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_580_6
timestamp 1730589202
transform 1 0 160 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_580_6
timestamp 1730589202
transform 1 0 160 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_581_6
timestamp 1730589202
transform 1 0 184 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_582_6
timestamp 1730589202
transform 1 0 224 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_582_6
timestamp 1730589202
transform 1 0 224 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_583_6
timestamp 1730589202
transform 1 0 272 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_583_6
timestamp 1730589202
transform 1 0 272 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_584_6
timestamp 1730589202
transform 1 0 328 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_584_6
timestamp 1730589202
transform 1 0 328 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_595_6
timestamp 1730589202
transform 1 0 384 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_595_6
timestamp 1730589202
transform 1 0 384 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_596_6
timestamp 1730589202
transform 1 0 448 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_596_6
timestamp 1730589202
transform 1 0 448 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_597_6
timestamp 1730589202
transform 1 0 512 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_597_6
timestamp 1730589202
transform 1 0 512 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5107_6
timestamp 1730589202
transform 1 0 568 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5107_6
timestamp 1730589202
transform 1 0 568 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5108_6
timestamp 1730589202
transform 1 0 624 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5108_6
timestamp 1730589202
transform 1 0 624 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_533_6
timestamp 1730589202
transform 1 0 672 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_533_6
timestamp 1730589202
transform 1 0 672 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_532_6
timestamp 1730589202
transform 1 0 720 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_532_6
timestamp 1730589202
transform 1 0 720 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_531_6
timestamp 1730589202
transform 1 0 760 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_531_6
timestamp 1730589202
transform 1 0 760 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_530_6
timestamp 1730589202
transform 1 0 792 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_529_6
timestamp 1730589202
transform 1 0 824 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_529_6
timestamp 1730589202
transform 1 0 824 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_530_6
timestamp 1730589202
transform 1 0 792 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_528_6
timestamp 1730589202
transform 1 0 856 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_528_6
timestamp 1730589202
transform 1 0 856 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_527_6
timestamp 1730589202
transform 1 0 888 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_527_6
timestamp 1730589202
transform 1 0 888 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_526_6
timestamp 1730589202
transform 1 0 920 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_526_6
timestamp 1730589202
transform 1 0 920 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_525_6
timestamp 1730589202
transform 1 0 960 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_525_6
timestamp 1730589202
transform 1 0 960 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_515_6
timestamp 1730589202
transform 1 0 1000 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_515_6
timestamp 1730589202
transform 1 0 1000 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_516_6
timestamp 1730589202
transform 1 0 1048 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_516_6
timestamp 1730589202
transform 1 0 1048 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5141_6
timestamp 1730589202
transform 1 0 1096 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5141_6
timestamp 1730589202
transform 1 0 1096 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5162_6
timestamp 1730589202
transform 1 0 1152 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5162_6
timestamp 1730589202
transform 1 0 1152 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5163_6
timestamp 1730589202
transform 1 0 1208 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5163_6
timestamp 1730589202
transform 1 0 1208 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5173_6
timestamp 1730589202
transform 1 0 1264 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5173_6
timestamp 1730589202
transform 1 0 1264 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5174_6
timestamp 1730589202
transform 1 0 1320 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5174_6
timestamp 1730589202
transform 1 0 1320 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5184_6
timestamp 1730589202
transform 1 0 1408 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5175_6
timestamp 1730589202
transform 1 0 1376 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5175_6
timestamp 1730589202
transform 1 0 1376 0 1 1308
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5184_6
timestamp 1730589202
transform 1 0 1408 0 1 1308
box 8 4 20 35
use welltap_svt  __well_tap__61
timestamp 1730589202
transform 1 0 1440 0 1 1312
box 8 4 12 24
use welltap_svt  __well_tap__61
timestamp 1730589202
transform 1 0 1440 0 1 1312
box 8 4 12 24
use welltap_svt  __well_tap__62
timestamp 1730589202
transform 1 0 104 0 -1 1384
box 8 4 12 24
use welltap_svt  __well_tap__62
timestamp 1730589202
transform 1 0 104 0 -1 1384
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_575_6
timestamp 1730589202
transform 1 0 152 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_574_6
timestamp 1730589202
transform 1 0 128 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_574_6
timestamp 1730589202
transform 1 0 128 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_575_6
timestamp 1730589202
transform 1 0 152 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_576_6
timestamp 1730589202
transform 1 0 176 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_576_6
timestamp 1730589202
transform 1 0 176 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_577_6
timestamp 1730589202
transform 1 0 224 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_577_6
timestamp 1730589202
transform 1 0 224 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_578_6
timestamp 1730589202
transform 1 0 272 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_578_6
timestamp 1730589202
transform 1 0 272 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_579_6
timestamp 1730589202
transform 1 0 328 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_579_6
timestamp 1730589202
transform 1 0 328 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_598_6
timestamp 1730589202
transform 1 0 384 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_598_6
timestamp 1730589202
transform 1 0 384 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_599_6
timestamp 1730589202
transform 1 0 432 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_599_6
timestamp 1730589202
transform 1 0 432 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5100_6
timestamp 1730589202
transform 1 0 480 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5100_6
timestamp 1730589202
transform 1 0 480 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5101_6
timestamp 1730589202
transform 1 0 520 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5101_6
timestamp 1730589202
transform 1 0 520 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5103_6
timestamp 1730589202
transform 1 0 560 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5103_6
timestamp 1730589202
transform 1 0 560 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5104_6
timestamp 1730589202
transform 1 0 608 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5104_6
timestamp 1730589202
transform 1 0 608 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5105_6
timestamp 1730589202
transform 1 0 656 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5105_6
timestamp 1730589202
transform 1 0 656 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5106_6
timestamp 1730589202
transform 1 0 704 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5106_6
timestamp 1730589202
transform 1 0 704 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_534_6
timestamp 1730589202
transform 1 0 760 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_534_6
timestamp 1730589202
transform 1 0 760 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_535_6
timestamp 1730589202
transform 1 0 816 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_535_6
timestamp 1730589202
transform 1 0 816 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_536_6
timestamp 1730589202
transform 1 0 872 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_536_6
timestamp 1730589202
transform 1 0 872 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_513_6
timestamp 1730589202
transform 1 0 928 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_513_6
timestamp 1730589202
transform 1 0 928 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_514_6
timestamp 1730589202
transform 1 0 984 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_514_6
timestamp 1730589202
transform 1 0 984 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5143_6
timestamp 1730589202
transform 1 0 1040 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5143_6
timestamp 1730589202
transform 1 0 1040 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5142_6
timestamp 1730589202
transform 1 0 1088 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5142_6
timestamp 1730589202
transform 1 0 1088 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5161_6
timestamp 1730589202
transform 1 0 1136 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5161_6
timestamp 1730589202
transform 1 0 1136 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5160_6
timestamp 1730589202
transform 1 0 1184 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5160_6
timestamp 1730589202
transform 1 0 1184 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5159_6
timestamp 1730589202
transform 1 0 1232 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5159_6
timestamp 1730589202
transform 1 0 1232 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5177_6
timestamp 1730589202
transform 1 0 1280 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5177_6
timestamp 1730589202
transform 1 0 1280 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5176_6
timestamp 1730589202
transform 1 0 1328 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5176_6
timestamp 1730589202
transform 1 0 1328 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5183_6
timestamp 1730589202
transform 1 0 1408 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5182_6
timestamp 1730589202
transform 1 0 1376 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5182_6
timestamp 1730589202
transform 1 0 1376 0 -1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5183_6
timestamp 1730589202
transform 1 0 1408 0 -1 1388
box 8 4 20 35
use welltap_svt  __well_tap__63
timestamp 1730589202
transform 1 0 1440 0 -1 1384
box 8 4 12 24
use welltap_svt  __well_tap__63
timestamp 1730589202
transform 1 0 1440 0 -1 1384
box 8 4 12 24
use welltap_svt  __well_tap__64
timestamp 1730589202
transform 1 0 104 0 1 1392
box 8 4 12 24
use welltap_svt  __well_tap__64
timestamp 1730589202
transform 1 0 104 0 1 1392
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_573_6
timestamp 1730589202
transform 1 0 128 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_572_6
timestamp 1730589202
transform 1 0 152 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_572_6
timestamp 1730589202
transform 1 0 152 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_573_6
timestamp 1730589202
transform 1 0 128 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_571_6
timestamp 1730589202
transform 1 0 176 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_571_6
timestamp 1730589202
transform 1 0 176 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_570_6
timestamp 1730589202
transform 1 0 216 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_570_6
timestamp 1730589202
transform 1 0 216 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_569_6
timestamp 1730589202
transform 1 0 280 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_569_6
timestamp 1730589202
transform 1 0 280 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_568_6
timestamp 1730589202
transform 1 0 344 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_568_6
timestamp 1730589202
transform 1 0 344 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_567_6
timestamp 1730589202
transform 1 0 408 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_567_6
timestamp 1730589202
transform 1 0 408 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5102_6
timestamp 1730589202
transform 1 0 472 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5102_6
timestamp 1730589202
transform 1 0 472 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_543_6
timestamp 1730589202
transform 1 0 528 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_543_6
timestamp 1730589202
transform 1 0 528 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_542_6
timestamp 1730589202
transform 1 0 576 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_542_6
timestamp 1730589202
transform 1 0 576 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_541_6
timestamp 1730589202
transform 1 0 624 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_541_6
timestamp 1730589202
transform 1 0 624 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_540_6
timestamp 1730589202
transform 1 0 680 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_540_6
timestamp 1730589202
transform 1 0 680 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_539_6
timestamp 1730589202
transform 1 0 736 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_539_6
timestamp 1730589202
transform 1 0 736 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_538_6
timestamp 1730589202
transform 1 0 792 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_538_6
timestamp 1730589202
transform 1 0 792 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_537_6
timestamp 1730589202
transform 1 0 848 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_537_6
timestamp 1730589202
transform 1 0 848 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_512_6
timestamp 1730589202
transform 1 0 904 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_512_6
timestamp 1730589202
transform 1 0 904 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_511_6
timestamp 1730589202
transform 1 0 960 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_511_6
timestamp 1730589202
transform 1 0 960 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_510_6
timestamp 1730589202
transform 1 0 1016 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_510_6
timestamp 1730589202
transform 1 0 1016 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5144_6
timestamp 1730589202
transform 1 0 1064 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5144_6
timestamp 1730589202
transform 1 0 1064 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5145_6
timestamp 1730589202
transform 1 0 1112 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5145_6
timestamp 1730589202
transform 1 0 1112 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5158_6
timestamp 1730589202
transform 1 0 1160 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5158_6
timestamp 1730589202
transform 1 0 1160 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5157_6
timestamp 1730589202
transform 1 0 1208 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5157_6
timestamp 1730589202
transform 1 0 1208 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5156_6
timestamp 1730589202
transform 1 0 1256 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5156_6
timestamp 1730589202
transform 1 0 1256 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5178_6
timestamp 1730589202
transform 1 0 1296 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5178_6
timestamp 1730589202
transform 1 0 1296 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5179_6
timestamp 1730589202
transform 1 0 1336 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5179_6
timestamp 1730589202
transform 1 0 1336 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5181_6
timestamp 1730589202
transform 1 0 1408 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5180_6
timestamp 1730589202
transform 1 0 1384 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5180_6
timestamp 1730589202
transform 1 0 1384 0 1 1388
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5181_6
timestamp 1730589202
transform 1 0 1408 0 1 1388
box 8 4 20 35
use welltap_svt  __well_tap__65
timestamp 1730589202
transform 1 0 1440 0 1 1392
box 8 4 12 24
use welltap_svt  __well_tap__65
timestamp 1730589202
transform 1 0 1440 0 1 1392
box 8 4 12 24
use welltap_svt  __well_tap__66
timestamp 1730589202
transform 1 0 104 0 -1 1464
box 8 4 12 24
use welltap_svt  __well_tap__66
timestamp 1730589202
transform 1 0 104 0 -1 1464
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_566_6
timestamp 1730589202
transform 1 0 144 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_566_6
timestamp 1730589202
transform 1 0 144 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_565_6
timestamp 1730589202
transform 1 0 168 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_564_6
timestamp 1730589202
transform 1 0 192 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_564_6
timestamp 1730589202
transform 1 0 192 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_565_6
timestamp 1730589202
transform 1 0 168 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_563_6
timestamp 1730589202
transform 1 0 224 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_563_6
timestamp 1730589202
transform 1 0 224 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_562_6
timestamp 1730589202
transform 1 0 264 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_562_6
timestamp 1730589202
transform 1 0 264 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_561_6
timestamp 1730589202
transform 1 0 312 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_561_6
timestamp 1730589202
transform 1 0 312 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_560_6
timestamp 1730589202
transform 1 0 360 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_560_6
timestamp 1730589202
transform 1 0 360 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_550_6
timestamp 1730589202
transform 1 0 400 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_550_6
timestamp 1730589202
transform 1 0 400 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_549_6
timestamp 1730589202
transform 1 0 448 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_549_6
timestamp 1730589202
transform 1 0 448 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_548_6
timestamp 1730589202
transform 1 0 496 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_548_6
timestamp 1730589202
transform 1 0 496 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_547_6
timestamp 1730589202
transform 1 0 544 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_547_6
timestamp 1730589202
transform 1 0 544 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_546_6
timestamp 1730589202
transform 1 0 600 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_546_6
timestamp 1730589202
transform 1 0 600 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_545_6
timestamp 1730589202
transform 1 0 656 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_545_6
timestamp 1730589202
transform 1 0 656 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_544_6
timestamp 1730589202
transform 1 0 704 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_544_6
timestamp 1730589202
transform 1 0 704 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_54_6
timestamp 1730589202
transform 1 0 752 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_54_6
timestamp 1730589202
transform 1 0 752 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_55_6
timestamp 1730589202
transform 1 0 808 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_55_6
timestamp 1730589202
transform 1 0 808 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_56_6
timestamp 1730589202
transform 1 0 864 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_56_6
timestamp 1730589202
transform 1 0 864 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_57_6
timestamp 1730589202
transform 1 0 920 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_57_6
timestamp 1730589202
transform 1 0 920 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_58_6
timestamp 1730589202
transform 1 0 968 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_58_6
timestamp 1730589202
transform 1 0 968 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_59_6
timestamp 1730589202
transform 1 0 1016 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_59_6
timestamp 1730589202
transform 1 0 1016 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5147_6
timestamp 1730589202
transform 1 0 1064 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5147_6
timestamp 1730589202
transform 1 0 1064 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5146_6
timestamp 1730589202
transform 1 0 1112 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5146_6
timestamp 1730589202
transform 1 0 1112 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5152_6
timestamp 1730589202
transform 1 0 1160 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5152_6
timestamp 1730589202
transform 1 0 1160 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5153_6
timestamp 1730589202
transform 1 0 1208 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5153_6
timestamp 1730589202
transform 1 0 1208 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5154_6
timestamp 1730589202
transform 1 0 1256 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5154_6
timestamp 1730589202
transform 1 0 1256 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5155_6
timestamp 1730589202
transform 1 0 1304 0 -1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5155_6
timestamp 1730589202
transform 1 0 1304 0 -1 1468
box 8 4 20 35
use welltap_svt  __well_tap__67
timestamp 1730589202
transform 1 0 1440 0 -1 1464
box 8 4 12 24
use welltap_svt  __well_tap__67
timestamp 1730589202
transform 1 0 1440 0 -1 1464
box 8 4 12 24
use welltap_svt  __well_tap__68
timestamp 1730589202
transform 1 0 104 0 1 1472
box 8 4 12 24
use welltap_svt  __well_tap__68
timestamp 1730589202
transform 1 0 104 0 1 1472
box 8 4 12 24
use _0_0std_0_0cells_0_0INVX1  inv_559_6
timestamp 1730589202
transform 1 0 288 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_558_6
timestamp 1730589202
transform 1 0 312 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_558_6
timestamp 1730589202
transform 1 0 312 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_559_6
timestamp 1730589202
transform 1 0 288 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_557_6
timestamp 1730589202
transform 1 0 336 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_556_6
timestamp 1730589202
transform 1 0 360 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_556_6
timestamp 1730589202
transform 1 0 360 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_557_6
timestamp 1730589202
transform 1 0 336 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_555_6
timestamp 1730589202
transform 1 0 400 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_555_6
timestamp 1730589202
transform 1 0 400 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_554_6
timestamp 1730589202
transform 1 0 448 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_554_6
timestamp 1730589202
transform 1 0 448 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_553_6
timestamp 1730589202
transform 1 0 504 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_553_6
timestamp 1730589202
transform 1 0 504 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_552_6
timestamp 1730589202
transform 1 0 568 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_552_6
timestamp 1730589202
transform 1 0 568 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_551_6
timestamp 1730589202
transform 1 0 640 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_551_6
timestamp 1730589202
transform 1 0 640 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_50_6
timestamp 1730589202
transform 1 0 720 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_50_6
timestamp 1730589202
transform 1 0 720 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_51_6
timestamp 1730589202
transform 1 0 800 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_51_6
timestamp 1730589202
transform 1 0 800 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_52_6
timestamp 1730589202
transform 1 0 880 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_52_6
timestamp 1730589202
transform 1 0 880 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_53_6
timestamp 1730589202
transform 1 0 952 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_53_6
timestamp 1730589202
transform 1 0 952 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5148_6
timestamp 1730589202
transform 1 0 1024 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5148_6
timestamp 1730589202
transform 1 0 1024 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5149_6
timestamp 1730589202
transform 1 0 1096 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5149_6
timestamp 1730589202
transform 1 0 1096 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5150_6
timestamp 1730589202
transform 1 0 1168 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5150_6
timestamp 1730589202
transform 1 0 1168 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5151_6
timestamp 1730589202
transform 1 0 1240 0 1 1468
box 8 4 20 35
use _0_0std_0_0cells_0_0INVX1  inv_5151_6
timestamp 1730589202
transform 1 0 1240 0 1 1468
box 8 4 20 35
use welltap_svt  __well_tap__69
timestamp 1730589202
transform 1 0 1440 0 1 1472
box 8 4 12 24
use welltap_svt  __well_tap__69
timestamp 1730589202
transform 1 0 1440 0 1 1472
box 8 4 12 24
<< end >>
