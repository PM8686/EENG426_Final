magic
tech sky130l
timestamp 1731220320
<< m1 >>
rect 638 1763 642 1800
rect 1190 1759 1194 1800
rect 240 1723 244 1743
rect 216 1691 220 1707
rect 272 1691 276 1707
rect 440 1691 444 1707
rect 552 1691 556 1707
rect 944 1691 948 1707
rect 1280 1691 1284 1707
rect 1360 1691 1364 1707
rect 1432 1691 1436 1707
rect 1488 1691 1492 1707
rect 1544 1691 1548 1707
rect 1592 1691 1596 1707
rect 80 1631 84 1670
rect 352 1595 356 1611
rect 464 1595 468 1611
rect 1748 1575 1752 1610
rect 80 1507 84 1538
rect 160 1515 164 1531
rect 248 1515 252 1531
rect 488 1515 492 1531
rect 800 1515 804 1531
rect 896 1515 900 1531
rect 1264 1467 1268 1539
rect 456 1443 460 1463
rect 80 1335 84 1402
rect 704 1379 708 1439
rect 728 1435 732 1463
rect 768 1431 772 1463
rect 1384 1415 1388 1463
rect 1748 1411 1752 1418
rect 1608 1379 1612 1395
rect 80 1235 84 1270
rect 608 1203 612 1307
rect 1448 1303 1452 1331
rect 736 1211 740 1291
rect 808 1155 812 1251
rect 1748 1222 1752 1259
rect 1288 1207 1292 1219
rect 80 1083 84 1138
rect 256 1015 260 1111
rect 288 1091 292 1111
rect 928 1019 932 1091
rect 1584 1091 1588 1111
rect 1072 1019 1076 1079
rect 1744 1076 1748 1167
rect 1744 1072 1752 1076
rect 1748 1030 1752 1072
rect 80 911 84 1006
rect 80 907 92 911
rect 88 875 92 907
rect 80 759 84 870
rect 160 807 164 911
rect 1104 883 1108 987
rect 1232 879 1236 987
rect 1544 983 1548 999
rect 208 831 212 871
rect 680 827 684 839
rect 1748 838 1752 879
rect 80 755 92 759
rect 80 699 84 738
rect 88 679 92 755
rect 264 639 268 759
rect 992 683 996 695
rect 264 635 292 639
rect 80 551 84 606
rect 272 527 276 635
rect 288 631 292 635
rect 1016 631 1020 651
rect 1748 646 1752 687
rect 1152 607 1156 627
rect 272 523 284 527
rect 80 470 84 483
rect 80 334 84 399
rect 160 383 164 523
rect 280 423 284 523
rect 768 487 772 547
rect 904 435 908 483
rect 1176 427 1180 595
rect 1504 591 1508 607
rect 1568 591 1572 607
rect 1632 591 1636 607
rect 1748 451 1752 458
rect 288 295 292 375
rect 936 323 940 399
rect 1504 363 1508 379
rect 1544 363 1548 379
rect 80 202 84 279
rect 1056 243 1060 291
rect 1748 262 1752 287
rect 1328 203 1332 219
rect 1464 203 1468 219
rect 1504 203 1508 219
rect 1544 203 1548 219
rect 576 95 580 111
rect 632 95 636 111
rect 696 95 700 111
rect 768 95 772 111
rect 848 95 852 111
rect 1080 95 1084 111
rect 1144 95 1148 111
rect 1200 87 1204 187
rect 638 72 642 83
rect 1190 83 1204 87
rect 1190 72 1194 83
<< m2c >>
rect 638 1759 642 1763
rect 1190 1755 1194 1759
rect 168 1743 172 1747
rect 200 1743 204 1747
rect 232 1743 236 1747
rect 240 1743 244 1747
rect 264 1743 268 1747
rect 296 1743 300 1747
rect 328 1743 332 1747
rect 360 1743 364 1747
rect 392 1743 396 1747
rect 424 1743 428 1747
rect 456 1743 460 1747
rect 488 1743 492 1747
rect 520 1743 524 1747
rect 552 1743 556 1747
rect 584 1743 588 1747
rect 616 1743 620 1747
rect 648 1743 652 1747
rect 680 1743 684 1747
rect 712 1743 716 1747
rect 744 1743 748 1747
rect 776 1743 780 1747
rect 808 1743 812 1747
rect 840 1743 844 1747
rect 872 1743 876 1747
rect 904 1743 908 1747
rect 936 1743 940 1747
rect 968 1743 972 1747
rect 1000 1743 1004 1747
rect 168 1727 172 1731
rect 200 1727 204 1731
rect 232 1727 236 1731
rect 264 1727 268 1731
rect 296 1727 300 1731
rect 328 1727 332 1731
rect 360 1727 364 1731
rect 392 1727 396 1731
rect 424 1727 428 1731
rect 456 1727 460 1731
rect 488 1727 492 1731
rect 520 1727 524 1731
rect 552 1727 556 1731
rect 584 1727 588 1731
rect 616 1727 620 1731
rect 648 1727 652 1731
rect 680 1727 684 1731
rect 712 1727 716 1731
rect 744 1727 748 1731
rect 776 1727 780 1731
rect 808 1727 812 1731
rect 840 1727 844 1731
rect 872 1727 876 1731
rect 904 1727 908 1731
rect 936 1727 940 1731
rect 968 1727 972 1731
rect 1000 1727 1004 1731
rect 240 1719 244 1723
rect 216 1707 220 1711
rect 272 1707 276 1711
rect 440 1707 444 1711
rect 552 1707 556 1711
rect 944 1707 948 1711
rect 1280 1707 1284 1711
rect 1360 1707 1364 1711
rect 1432 1707 1436 1711
rect 1488 1707 1492 1711
rect 1544 1707 1548 1711
rect 1592 1707 1596 1711
rect 208 1703 212 1707
rect 264 1703 268 1707
rect 336 1703 340 1707
rect 432 1703 436 1707
rect 544 1703 548 1707
rect 672 1703 676 1707
rect 808 1703 812 1707
rect 936 1703 940 1707
rect 1064 1703 1068 1707
rect 1176 1703 1180 1707
rect 1272 1703 1276 1707
rect 1352 1703 1356 1707
rect 1424 1703 1428 1707
rect 1480 1703 1484 1707
rect 1536 1703 1540 1707
rect 1584 1703 1588 1707
rect 1640 1703 1644 1707
rect 1672 1703 1676 1707
rect 208 1687 212 1691
rect 216 1687 220 1691
rect 264 1687 268 1691
rect 272 1687 276 1691
rect 336 1687 340 1691
rect 432 1687 436 1691
rect 440 1687 444 1691
rect 544 1687 548 1691
rect 552 1687 556 1691
rect 672 1687 676 1691
rect 808 1687 812 1691
rect 936 1687 940 1691
rect 944 1687 948 1691
rect 1064 1687 1068 1691
rect 1176 1687 1180 1691
rect 1272 1687 1276 1691
rect 1280 1687 1284 1691
rect 1352 1687 1356 1691
rect 1360 1687 1364 1691
rect 1424 1687 1428 1691
rect 1432 1687 1436 1691
rect 1480 1687 1484 1691
rect 1488 1687 1492 1691
rect 1536 1687 1540 1691
rect 1544 1687 1548 1691
rect 1584 1687 1588 1691
rect 1592 1687 1596 1691
rect 1640 1687 1644 1691
rect 1672 1687 1676 1691
rect 152 1651 156 1655
rect 192 1651 196 1655
rect 280 1651 284 1655
rect 408 1651 412 1655
rect 560 1651 564 1655
rect 728 1651 732 1655
rect 896 1651 900 1655
rect 1056 1651 1060 1655
rect 1200 1651 1204 1655
rect 1336 1651 1340 1655
rect 1456 1651 1460 1655
rect 1576 1651 1580 1655
rect 1672 1651 1676 1655
rect 152 1635 156 1639
rect 192 1635 196 1639
rect 280 1635 284 1639
rect 408 1635 412 1639
rect 560 1635 564 1639
rect 728 1635 732 1639
rect 896 1635 900 1639
rect 1056 1635 1060 1639
rect 1200 1635 1204 1639
rect 1336 1635 1340 1639
rect 1456 1635 1460 1639
rect 1576 1635 1580 1639
rect 1672 1635 1676 1639
rect 80 1627 84 1631
rect 352 1611 356 1615
rect 464 1611 468 1615
rect 152 1607 156 1611
rect 184 1607 188 1611
rect 216 1607 220 1611
rect 264 1607 268 1611
rect 344 1607 348 1611
rect 456 1607 460 1611
rect 584 1607 588 1611
rect 728 1607 732 1611
rect 872 1607 876 1611
rect 1016 1607 1020 1611
rect 1144 1607 1148 1611
rect 1264 1607 1268 1611
rect 1376 1607 1380 1611
rect 1480 1607 1484 1611
rect 1584 1607 1588 1611
rect 1672 1607 1676 1611
rect 152 1591 156 1595
rect 184 1591 188 1595
rect 216 1591 220 1595
rect 264 1591 268 1595
rect 344 1591 348 1595
rect 352 1591 356 1595
rect 456 1591 460 1595
rect 464 1591 468 1595
rect 584 1591 588 1595
rect 728 1591 732 1595
rect 872 1591 876 1595
rect 1016 1591 1020 1595
rect 1144 1591 1148 1595
rect 1264 1591 1268 1595
rect 1376 1591 1380 1595
rect 1480 1591 1484 1595
rect 1584 1591 1588 1595
rect 1672 1591 1676 1595
rect 1748 1571 1752 1575
rect 152 1563 156 1567
rect 184 1563 188 1567
rect 248 1563 252 1567
rect 304 1563 308 1567
rect 360 1563 364 1567
rect 416 1563 420 1567
rect 472 1563 476 1567
rect 528 1563 532 1567
rect 592 1563 596 1567
rect 672 1563 676 1567
rect 768 1563 772 1567
rect 872 1563 876 1567
rect 976 1563 980 1567
rect 1080 1563 1084 1567
rect 1176 1563 1180 1567
rect 1264 1563 1268 1567
rect 1344 1563 1348 1567
rect 1416 1563 1420 1567
rect 1488 1563 1492 1567
rect 1552 1563 1556 1567
rect 1624 1563 1628 1567
rect 1672 1563 1676 1567
rect 152 1547 156 1551
rect 184 1547 188 1551
rect 248 1547 252 1551
rect 304 1547 308 1551
rect 360 1547 364 1551
rect 416 1547 420 1551
rect 472 1547 476 1551
rect 528 1547 532 1551
rect 592 1547 596 1551
rect 672 1547 676 1551
rect 768 1547 772 1551
rect 872 1547 876 1551
rect 976 1547 980 1551
rect 1080 1547 1084 1551
rect 1176 1547 1180 1551
rect 1264 1547 1268 1551
rect 1344 1547 1348 1551
rect 1416 1547 1420 1551
rect 1488 1547 1492 1551
rect 1552 1547 1556 1551
rect 1624 1547 1628 1551
rect 1672 1547 1676 1551
rect 1264 1539 1268 1543
rect 160 1531 164 1535
rect 248 1531 252 1535
rect 488 1531 492 1535
rect 800 1531 804 1535
rect 896 1531 900 1535
rect 152 1527 156 1531
rect 192 1527 196 1531
rect 240 1527 244 1531
rect 296 1527 300 1531
rect 352 1527 356 1531
rect 416 1527 420 1531
rect 480 1527 484 1531
rect 552 1527 556 1531
rect 624 1527 628 1531
rect 704 1527 708 1531
rect 792 1527 796 1531
rect 888 1527 892 1531
rect 992 1527 996 1531
rect 1096 1527 1100 1531
rect 1192 1527 1196 1531
rect 152 1511 156 1515
rect 160 1511 164 1515
rect 192 1511 196 1515
rect 240 1511 244 1515
rect 248 1511 252 1515
rect 296 1511 300 1515
rect 352 1511 356 1515
rect 416 1511 420 1515
rect 480 1511 484 1515
rect 488 1511 492 1515
rect 552 1511 556 1515
rect 624 1511 628 1515
rect 704 1511 708 1515
rect 792 1511 796 1515
rect 800 1511 804 1515
rect 888 1511 892 1515
rect 896 1511 900 1515
rect 992 1511 996 1515
rect 1096 1511 1100 1515
rect 1192 1511 1196 1515
rect 80 1503 84 1507
rect 860 1487 864 1491
rect 988 1487 992 1491
rect 1288 1527 1292 1531
rect 1376 1527 1380 1531
rect 1456 1527 1460 1531
rect 1536 1527 1540 1531
rect 1616 1527 1620 1531
rect 1672 1527 1676 1531
rect 1288 1511 1292 1515
rect 1376 1511 1380 1515
rect 1456 1511 1460 1515
rect 1536 1511 1540 1515
rect 1616 1511 1620 1515
rect 1672 1511 1676 1515
rect 192 1463 196 1467
rect 224 1463 228 1467
rect 256 1463 260 1467
rect 288 1463 292 1467
rect 320 1463 324 1467
rect 352 1463 356 1467
rect 384 1463 388 1467
rect 416 1463 420 1467
rect 448 1463 452 1467
rect 456 1463 460 1467
rect 480 1463 484 1467
rect 512 1463 516 1467
rect 544 1463 548 1467
rect 576 1463 580 1467
rect 608 1463 612 1467
rect 640 1463 644 1467
rect 680 1463 684 1467
rect 720 1463 724 1467
rect 728 1463 732 1467
rect 760 1463 764 1467
rect 768 1463 772 1467
rect 792 1463 796 1467
rect 1096 1463 1100 1467
rect 1184 1463 1188 1467
rect 1216 1463 1220 1467
rect 1256 1463 1260 1467
rect 1264 1463 1268 1467
rect 1296 1463 1300 1467
rect 1336 1463 1340 1467
rect 1376 1463 1380 1467
rect 1384 1463 1388 1467
rect 1416 1463 1420 1467
rect 1456 1463 1460 1467
rect 1496 1463 1500 1467
rect 1536 1463 1540 1467
rect 1576 1463 1580 1467
rect 1608 1463 1612 1467
rect 1640 1463 1644 1467
rect 1672 1463 1676 1467
rect 192 1447 196 1451
rect 224 1447 228 1451
rect 256 1447 260 1451
rect 288 1447 292 1451
rect 320 1447 324 1451
rect 352 1447 356 1451
rect 384 1447 388 1451
rect 416 1447 420 1451
rect 448 1447 452 1451
rect 480 1447 484 1451
rect 512 1447 516 1451
rect 544 1447 548 1451
rect 576 1447 580 1451
rect 608 1447 612 1451
rect 640 1447 644 1451
rect 680 1447 684 1451
rect 720 1447 724 1451
rect 456 1439 460 1443
rect 704 1439 708 1443
rect 152 1391 156 1395
rect 184 1391 188 1395
rect 216 1391 220 1395
rect 248 1391 252 1395
rect 280 1391 284 1395
rect 312 1391 316 1395
rect 344 1391 348 1395
rect 376 1391 380 1395
rect 408 1391 412 1395
rect 440 1391 444 1395
rect 472 1391 476 1395
rect 504 1391 508 1395
rect 536 1391 540 1395
rect 568 1391 572 1395
rect 600 1391 604 1395
rect 632 1391 636 1395
rect 664 1391 668 1395
rect 696 1391 700 1395
rect 152 1375 156 1379
rect 184 1375 188 1379
rect 216 1375 220 1379
rect 248 1375 252 1379
rect 280 1375 284 1379
rect 312 1375 316 1379
rect 344 1375 348 1379
rect 376 1375 380 1379
rect 408 1375 412 1379
rect 440 1375 444 1379
rect 472 1375 476 1379
rect 504 1375 508 1379
rect 536 1375 540 1379
rect 568 1376 572 1380
rect 760 1447 764 1451
rect 728 1431 732 1435
rect 920 1455 924 1459
rect 1060 1451 1064 1455
rect 1148 1451 1152 1455
rect 792 1447 796 1451
rect 1096 1447 1100 1451
rect 1184 1447 1188 1451
rect 1216 1447 1220 1451
rect 1256 1447 1260 1451
rect 1296 1447 1300 1451
rect 1336 1447 1340 1451
rect 1376 1447 1380 1451
rect 856 1435 860 1439
rect 920 1435 924 1439
rect 984 1435 988 1439
rect 1044 1435 1048 1439
rect 1132 1435 1136 1439
rect 892 1431 896 1435
rect 1020 1431 1024 1435
rect 1108 1431 1112 1435
rect 768 1427 772 1431
rect 764 1419 768 1423
rect 792 1417 796 1421
rect 836 1419 840 1423
rect 972 1419 976 1423
rect 864 1415 868 1419
rect 888 1415 892 1419
rect 904 1415 908 1419
rect 920 1415 924 1419
rect 1000 1416 1004 1420
rect 1416 1447 1420 1451
rect 1456 1447 1460 1451
rect 1496 1447 1500 1451
rect 1536 1447 1540 1451
rect 1576 1447 1580 1451
rect 1608 1447 1612 1451
rect 1640 1447 1644 1451
rect 1672 1447 1676 1451
rect 1060 1409 1064 1413
rect 1384 1411 1388 1415
rect 1148 1407 1152 1411
rect 1244 1407 1248 1411
rect 1460 1409 1464 1413
rect 1088 1403 1092 1407
rect 1176 1403 1180 1407
rect 1268 1405 1272 1409
rect 1748 1407 1752 1411
rect 1368 1403 1372 1407
rect 1484 1403 1488 1407
rect 720 1399 724 1403
rect 752 1392 756 1396
rect 1040 1391 1044 1395
rect 1128 1391 1132 1395
rect 1216 1393 1220 1397
rect 1432 1393 1436 1397
rect 1608 1395 1612 1399
rect 1284 1389 1288 1393
rect 1552 1391 1556 1395
rect 1600 1391 1604 1395
rect 1500 1387 1504 1391
rect 792 1383 796 1387
rect 864 1383 868 1387
rect 1000 1383 1004 1387
rect 1088 1383 1092 1387
rect 1176 1383 1180 1387
rect 1640 1391 1644 1395
rect 1672 1391 1676 1395
rect 600 1375 604 1379
rect 632 1375 636 1379
rect 664 1375 668 1379
rect 696 1375 700 1379
rect 704 1375 708 1379
rect 1040 1375 1044 1379
rect 1128 1375 1132 1379
rect 1216 1375 1220 1379
rect 1432 1375 1436 1379
rect 1552 1375 1556 1379
rect 1600 1375 1604 1379
rect 1608 1375 1612 1379
rect 1640 1375 1644 1379
rect 1672 1375 1676 1379
rect 824 1371 828 1375
rect 712 1355 716 1359
rect 1372 1351 1376 1355
rect 1116 1339 1120 1343
rect 80 1331 84 1335
rect 1268 1331 1272 1335
rect 1356 1331 1360 1335
rect 1448 1331 1452 1335
rect 152 1307 156 1311
rect 184 1307 188 1311
rect 216 1307 220 1311
rect 248 1307 252 1311
rect 280 1307 284 1311
rect 312 1307 316 1311
rect 344 1307 348 1311
rect 376 1307 380 1311
rect 408 1307 412 1311
rect 440 1307 444 1311
rect 472 1307 476 1311
rect 504 1307 508 1311
rect 536 1307 540 1311
rect 568 1307 572 1311
rect 600 1307 604 1311
rect 608 1307 612 1311
rect 632 1307 636 1311
rect 664 1307 668 1311
rect 696 1307 700 1311
rect 728 1307 732 1311
rect 1408 1307 1412 1311
rect 1440 1307 1444 1311
rect 152 1291 156 1295
rect 184 1291 188 1295
rect 216 1291 220 1295
rect 248 1291 252 1295
rect 280 1291 284 1295
rect 312 1291 316 1295
rect 344 1291 348 1295
rect 376 1291 380 1295
rect 408 1291 412 1295
rect 440 1291 444 1295
rect 472 1291 476 1295
rect 504 1291 508 1295
rect 536 1291 540 1295
rect 568 1291 572 1295
rect 600 1291 604 1295
rect 80 1231 84 1235
rect 1512 1307 1516 1311
rect 1544 1307 1548 1311
rect 1576 1307 1580 1311
rect 1608 1307 1612 1311
rect 1640 1307 1644 1311
rect 1672 1307 1676 1311
rect 1008 1299 1012 1303
rect 1048 1299 1052 1303
rect 1376 1299 1380 1303
rect 1448 1299 1452 1303
rect 1480 1299 1484 1303
rect 1196 1295 1200 1299
rect 632 1291 636 1295
rect 664 1291 668 1295
rect 696 1291 700 1295
rect 728 1291 732 1295
rect 736 1291 740 1295
rect 1408 1291 1412 1295
rect 1440 1291 1444 1295
rect 1512 1291 1516 1295
rect 1544 1291 1548 1295
rect 1576 1291 1580 1295
rect 1608 1291 1612 1295
rect 1640 1291 1644 1295
rect 1672 1291 1676 1295
rect 1048 1279 1052 1283
rect 1100 1279 1104 1283
rect 1180 1279 1184 1283
rect 1264 1279 1268 1283
rect 1352 1279 1356 1283
rect 1480 1279 1484 1283
rect 1020 1275 1024 1279
rect 1128 1275 1132 1279
rect 1156 1275 1160 1279
rect 1452 1275 1456 1279
rect 744 1267 748 1271
rect 760 1267 764 1271
rect 776 1267 780 1271
rect 824 1267 828 1271
rect 840 1267 844 1271
rect 856 1268 860 1272
rect 904 1267 908 1271
rect 920 1267 924 1271
rect 936 1267 940 1271
rect 1008 1267 1012 1271
rect 980 1263 984 1267
rect 1748 1259 1752 1263
rect 808 1251 812 1255
rect 772 1223 776 1227
rect 800 1219 804 1223
rect 736 1207 740 1211
rect 608 1199 612 1203
rect 152 1195 156 1199
rect 184 1195 188 1199
rect 216 1195 220 1199
rect 248 1195 252 1199
rect 280 1195 284 1199
rect 312 1195 316 1199
rect 344 1195 348 1199
rect 376 1195 380 1199
rect 408 1195 412 1199
rect 440 1195 444 1199
rect 472 1195 476 1199
rect 504 1195 508 1199
rect 536 1195 540 1199
rect 568 1195 572 1199
rect 600 1195 604 1199
rect 632 1195 636 1199
rect 664 1195 668 1199
rect 696 1195 700 1199
rect 728 1195 732 1199
rect 760 1195 764 1199
rect 800 1187 804 1191
rect 152 1179 156 1183
rect 184 1179 188 1183
rect 216 1179 220 1183
rect 248 1179 252 1183
rect 280 1179 284 1183
rect 312 1179 316 1183
rect 344 1179 348 1183
rect 376 1179 380 1183
rect 408 1179 412 1183
rect 440 1179 444 1183
rect 472 1179 476 1183
rect 504 1179 508 1183
rect 536 1179 540 1183
rect 568 1179 572 1183
rect 600 1179 604 1183
rect 632 1179 636 1183
rect 664 1179 668 1183
rect 696 1179 700 1183
rect 728 1179 732 1183
rect 760 1179 764 1183
rect 1084 1223 1088 1227
rect 1008 1219 1012 1223
rect 1024 1219 1028 1223
rect 1040 1219 1044 1223
rect 1112 1219 1116 1223
rect 1288 1219 1292 1223
rect 1196 1211 1200 1215
rect 1220 1207 1224 1211
rect 960 1203 964 1207
rect 1288 1203 1292 1207
rect 1296 1203 1300 1207
rect 936 1199 940 1203
rect 992 1195 996 1199
rect 1144 1195 1148 1199
rect 1176 1195 1180 1199
rect 1272 1195 1276 1199
rect 1328 1195 1332 1199
rect 1360 1195 1364 1199
rect 1392 1195 1396 1199
rect 1424 1195 1428 1199
rect 1456 1195 1460 1199
rect 1496 1195 1500 1199
rect 1536 1195 1540 1199
rect 1576 1195 1580 1199
rect 1608 1195 1612 1199
rect 1640 1195 1644 1199
rect 1672 1195 1676 1199
rect 1236 1191 1240 1195
rect 1112 1187 1116 1191
rect 1144 1179 1148 1183
rect 1176 1179 1180 1183
rect 1272 1179 1276 1183
rect 1360 1179 1364 1183
rect 1392 1179 1396 1183
rect 1424 1179 1428 1183
rect 1456 1179 1460 1183
rect 1496 1179 1500 1183
rect 1536 1179 1540 1183
rect 1576 1179 1580 1183
rect 1608 1179 1612 1183
rect 1640 1179 1644 1183
rect 1672 1179 1676 1183
rect 936 1175 940 1179
rect 1744 1167 1748 1171
rect 952 1159 956 1163
rect 1288 1159 1292 1163
rect 808 1151 812 1155
rect 784 1115 788 1119
rect 816 1115 820 1119
rect 1016 1115 1020 1119
rect 152 1111 156 1115
rect 184 1111 188 1115
rect 216 1111 220 1115
rect 248 1111 252 1115
rect 256 1111 260 1115
rect 280 1111 284 1115
rect 288 1111 292 1115
rect 312 1111 316 1115
rect 344 1111 348 1115
rect 376 1111 380 1115
rect 408 1111 412 1115
rect 440 1111 444 1115
rect 472 1111 476 1115
rect 504 1111 508 1115
rect 536 1111 540 1115
rect 568 1111 572 1115
rect 952 1111 956 1115
rect 984 1111 988 1115
rect 1048 1111 1052 1115
rect 1080 1111 1084 1115
rect 1152 1111 1156 1115
rect 1304 1111 1308 1115
rect 1440 1111 1444 1115
rect 1472 1111 1476 1115
rect 1504 1111 1508 1115
rect 1536 1111 1540 1115
rect 1576 1111 1580 1115
rect 1584 1111 1588 1115
rect 1608 1111 1612 1115
rect 1640 1111 1644 1115
rect 1672 1111 1676 1115
rect 152 1095 156 1099
rect 184 1095 188 1099
rect 216 1095 220 1099
rect 248 1095 252 1099
rect 80 1079 84 1083
rect 280 1095 284 1099
rect 1120 1103 1124 1107
rect 1272 1103 1276 1107
rect 312 1095 316 1099
rect 344 1095 348 1099
rect 376 1095 380 1099
rect 408 1095 412 1099
rect 440 1095 444 1099
rect 472 1095 476 1099
rect 504 1095 508 1099
rect 536 1095 540 1099
rect 568 1095 572 1099
rect 952 1095 956 1099
rect 984 1095 988 1099
rect 1048 1095 1052 1099
rect 1080 1095 1084 1099
rect 1152 1095 1156 1099
rect 1304 1095 1308 1099
rect 1440 1095 1444 1099
rect 1472 1095 1476 1099
rect 1504 1095 1508 1099
rect 1536 1095 1540 1099
rect 1576 1095 1580 1099
rect 784 1091 788 1095
rect 928 1091 932 1095
rect 288 1087 292 1091
rect 584 1071 588 1075
rect 600 1071 604 1075
rect 616 1071 620 1075
rect 864 1071 868 1075
rect 920 1073 924 1077
rect 500 1023 504 1027
rect 400 1019 404 1023
rect 416 1019 420 1023
rect 432 1019 436 1023
rect 528 1019 532 1023
rect 600 1019 604 1023
rect 656 1019 660 1023
rect 728 1019 732 1023
rect 784 1019 788 1023
rect 1608 1095 1612 1099
rect 1640 1095 1644 1099
rect 1672 1095 1676 1099
rect 1584 1087 1588 1091
rect 1120 1083 1124 1087
rect 1072 1079 1076 1083
rect 1092 1079 1096 1083
rect 816 1015 820 1019
rect 832 1015 836 1019
rect 852 1015 856 1019
rect 928 1015 932 1019
rect 968 1015 972 1019
rect 984 1015 988 1019
rect 1004 1017 1008 1021
rect 1168 1071 1172 1075
rect 1184 1071 1188 1075
rect 1200 1071 1204 1075
rect 1272 1071 1276 1075
rect 1352 1071 1356 1075
rect 1408 1071 1412 1075
rect 1244 1067 1248 1071
rect 256 1011 260 1015
rect 1060 1013 1064 1017
rect 1072 1015 1076 1019
rect 1196 1013 1200 1017
rect 1324 1013 1328 1017
rect 1364 1013 1368 1017
rect 1088 1007 1092 1011
rect 1224 1007 1228 1011
rect 1352 1007 1356 1011
rect 1392 1007 1396 1011
rect 328 1003 332 1007
rect 1120 1003 1124 1007
rect 1248 1003 1252 1007
rect 1544 999 1548 1003
rect 152 995 156 999
rect 184 995 188 999
rect 216 995 220 999
rect 248 995 252 999
rect 280 995 284 999
rect 360 995 364 999
rect 936 995 940 999
rect 1152 995 1156 999
rect 1184 995 1188 999
rect 1280 995 1284 999
rect 1312 995 1316 999
rect 1424 995 1428 999
rect 1456 995 1460 999
rect 1496 995 1500 999
rect 1536 995 1540 999
rect 528 987 532 991
rect 1088 987 1092 991
rect 1104 987 1108 991
rect 1224 987 1228 991
rect 1232 987 1236 991
rect 1352 987 1356 991
rect 1392 987 1396 991
rect 152 979 156 983
rect 184 979 188 983
rect 216 979 220 983
rect 248 979 252 983
rect 280 979 284 983
rect 936 979 940 983
rect 320 959 324 963
rect 560 915 564 919
rect 696 915 700 919
rect 152 911 156 915
rect 160 911 164 915
rect 184 911 188 915
rect 832 911 836 915
rect 968 911 972 915
rect 1056 911 1060 915
rect 152 895 156 899
rect 88 871 92 875
rect 304 903 308 907
rect 424 903 428 907
rect 1096 903 1100 907
rect 1020 899 1024 903
rect 184 895 188 899
rect 832 895 836 899
rect 968 895 972 899
rect 1056 895 1060 899
rect 560 891 564 895
rect 1004 883 1008 887
rect 980 879 984 883
rect 1068 881 1072 885
rect 1096 883 1100 887
rect 1184 979 1188 983
rect 1112 959 1116 963
rect 1196 941 1200 945
rect 1128 911 1132 915
rect 1128 895 1132 899
rect 1180 883 1184 887
rect 1104 879 1108 883
rect 1208 879 1212 883
rect 1576 995 1580 999
rect 1608 995 1612 999
rect 1640 995 1644 999
rect 1672 995 1676 999
rect 1312 979 1316 983
rect 1424 979 1428 983
rect 1456 979 1460 983
rect 1496 979 1500 983
rect 1536 979 1540 983
rect 1544 979 1548 983
rect 1576 979 1580 983
rect 1608 979 1612 983
rect 1640 979 1644 983
rect 1672 979 1676 983
rect 1240 959 1244 963
rect 1324 943 1328 947
rect 1368 931 1372 935
rect 1256 911 1260 915
rect 1440 911 1444 915
rect 1536 911 1540 915
rect 1576 911 1580 915
rect 1608 911 1612 915
rect 1640 911 1644 915
rect 1672 911 1676 915
rect 1492 899 1496 903
rect 1256 895 1260 899
rect 1408 895 1412 899
rect 1440 895 1444 899
rect 1536 895 1540 899
rect 1576 895 1580 899
rect 1608 895 1612 899
rect 1640 895 1644 899
rect 1672 895 1676 899
rect 1376 887 1380 891
rect 1308 883 1312 887
rect 1476 883 1480 887
rect 1336 879 1340 883
rect 1452 879 1456 883
rect 1748 879 1752 883
rect 1232 875 1236 879
rect 200 871 204 875
rect 208 871 212 875
rect 216 871 220 875
rect 232 871 236 875
rect 304 871 308 875
rect 320 871 324 875
rect 336 871 340 875
rect 352 871 356 875
rect 424 871 428 875
rect 608 871 612 875
rect 664 871 668 875
rect 712 871 716 875
rect 744 871 748 875
rect 800 871 804 875
rect 880 871 884 875
rect 936 871 940 875
rect 276 867 280 871
rect 396 867 400 871
rect 680 839 684 843
rect 208 827 212 831
rect 216 827 220 831
rect 248 827 252 831
rect 304 827 308 831
rect 392 827 396 831
rect 424 827 428 831
rect 480 827 484 831
rect 800 827 804 831
rect 832 827 836 831
rect 888 827 892 831
rect 656 823 660 827
rect 672 823 676 827
rect 680 823 684 827
rect 692 823 696 827
rect 1012 819 1016 823
rect 1036 817 1040 821
rect 1228 819 1232 823
rect 1252 815 1256 819
rect 1364 817 1368 821
rect 1392 819 1396 823
rect 1420 819 1424 823
rect 1468 819 1472 823
rect 1448 815 1452 819
rect 1496 815 1500 819
rect 1168 811 1172 815
rect 152 803 156 807
rect 160 803 164 807
rect 576 803 580 807
rect 1120 803 1124 807
rect 1200 803 1204 807
rect 1312 803 1316 807
rect 1536 803 1540 807
rect 1576 803 1580 807
rect 1608 803 1612 807
rect 1640 803 1644 807
rect 1672 803 1676 807
rect 1052 799 1056 803
rect 1268 799 1272 803
rect 1448 795 1452 799
rect 1496 795 1500 799
rect 152 787 156 791
rect 576 787 580 791
rect 1120 787 1124 791
rect 1312 787 1316 791
rect 1536 787 1540 791
rect 1576 787 1580 791
rect 1608 787 1612 791
rect 1640 787 1644 791
rect 1672 787 1676 791
rect 968 783 972 787
rect 1160 767 1164 771
rect 264 759 268 763
rect 80 695 84 699
rect 240 707 244 711
rect 88 675 92 679
rect 136 675 140 679
rect 152 677 156 681
rect 168 675 172 679
rect 240 675 244 679
rect 212 671 216 675
rect 1380 755 1384 759
rect 568 719 572 723
rect 736 719 740 723
rect 880 715 884 719
rect 1264 715 1268 719
rect 1296 715 1300 719
rect 1328 715 1332 719
rect 1360 715 1364 719
rect 1392 715 1396 719
rect 1424 715 1428 719
rect 1456 715 1460 719
rect 1496 715 1500 719
rect 1536 715 1540 719
rect 1576 715 1580 719
rect 1608 715 1612 719
rect 1640 715 1644 719
rect 1672 715 1676 719
rect 416 707 420 711
rect 1192 707 1196 711
rect 1232 707 1236 711
rect 880 699 884 703
rect 1264 699 1268 703
rect 1296 699 1300 703
rect 1328 699 1332 703
rect 1360 699 1364 703
rect 1392 699 1396 703
rect 1424 699 1428 703
rect 1456 699 1460 703
rect 1496 699 1500 703
rect 1536 699 1540 703
rect 1576 699 1580 703
rect 1608 699 1612 703
rect 1640 699 1644 703
rect 1672 699 1676 703
rect 568 695 572 699
rect 992 695 996 699
rect 600 687 604 691
rect 1232 687 1236 691
rect 1748 687 1752 691
rect 1204 683 1208 687
rect 768 679 772 683
rect 784 679 788 683
rect 804 679 808 683
rect 992 679 996 683
rect 1000 679 1004 683
rect 1016 679 1020 683
rect 1036 679 1040 683
rect 304 675 308 679
rect 360 675 364 679
rect 416 675 420 679
rect 632 675 636 679
rect 688 675 692 679
rect 928 675 932 679
rect 984 675 988 679
rect 1088 675 1092 679
rect 1104 675 1108 679
rect 1120 675 1124 679
rect 1192 675 1196 679
rect 388 671 392 675
rect 1164 671 1168 675
rect 1016 651 1020 655
rect 204 633 208 637
rect 232 627 236 631
rect 152 603 156 607
rect 184 603 188 607
rect 232 595 236 599
rect 152 587 156 591
rect 184 587 188 591
rect 80 547 84 551
rect 900 631 904 635
rect 1116 631 1120 635
rect 1332 631 1336 635
rect 280 627 284 631
rect 288 627 292 631
rect 296 627 300 631
rect 312 627 316 631
rect 400 627 404 631
rect 416 627 420 631
rect 432 627 436 631
rect 552 627 556 631
rect 608 627 612 631
rect 784 627 788 631
rect 840 627 844 631
rect 928 627 932 631
rect 992 627 996 631
rect 1008 627 1012 631
rect 1016 627 1020 631
rect 1024 627 1028 631
rect 1144 627 1148 631
rect 1152 627 1156 631
rect 1208 627 1212 631
rect 1224 627 1228 631
rect 1240 627 1244 631
rect 1360 627 1364 631
rect 1504 607 1508 611
rect 1568 607 1572 611
rect 1632 607 1636 611
rect 688 603 692 607
rect 1152 603 1156 607
rect 1432 603 1436 607
rect 1496 603 1500 607
rect 928 595 932 599
rect 1144 595 1148 599
rect 1176 595 1180 599
rect 1360 595 1364 599
rect 688 587 692 591
rect 768 547 772 551
rect 632 527 636 531
rect 152 523 156 527
rect 160 523 164 527
rect 152 507 156 511
rect 80 483 84 487
rect 80 399 84 403
rect 272 515 276 519
rect 168 483 172 487
rect 184 483 188 487
rect 200 483 204 487
rect 272 483 276 487
rect 244 479 248 483
rect 496 515 500 519
rect 752 515 756 519
rect 632 503 636 507
rect 320 483 324 487
rect 376 483 380 487
rect 392 483 396 487
rect 408 484 412 488
rect 896 515 900 519
rect 1056 515 1060 519
rect 424 483 428 487
rect 496 483 500 487
rect 648 483 652 487
rect 664 483 668 487
rect 680 483 684 487
rect 752 483 756 487
rect 768 483 772 487
rect 776 483 780 487
rect 792 483 796 487
rect 808 483 812 487
rect 896 483 900 487
rect 904 483 908 487
rect 928 483 932 487
rect 944 483 948 487
rect 960 483 964 487
rect 1056 483 1060 487
rect 1096 483 1100 487
rect 1112 483 1116 487
rect 1128 483 1132 487
rect 468 479 472 483
rect 724 479 728 483
rect 868 479 872 483
rect 1028 479 1032 483
rect 904 431 908 435
rect 1560 603 1564 607
rect 1624 603 1628 607
rect 1672 603 1676 607
rect 1432 587 1436 591
rect 1496 587 1500 591
rect 1504 587 1508 591
rect 1560 587 1564 591
rect 1568 587 1572 591
rect 1624 587 1628 591
rect 1632 587 1636 591
rect 1672 587 1676 591
rect 1384 527 1388 531
rect 1440 523 1444 527
rect 1496 523 1500 527
rect 1544 523 1548 527
rect 1592 523 1596 527
rect 1640 523 1644 527
rect 1672 523 1676 527
rect 1224 515 1228 519
rect 1440 507 1444 511
rect 1496 507 1500 511
rect 1544 507 1548 511
rect 1592 507 1596 511
rect 1640 507 1644 511
rect 1672 507 1676 511
rect 1224 483 1228 487
rect 1196 479 1200 483
rect 1748 447 1752 451
rect 1176 423 1180 427
rect 280 419 284 423
rect 372 403 376 407
rect 612 403 616 407
rect 296 399 300 403
rect 312 399 316 403
rect 328 399 332 403
rect 400 399 404 403
rect 536 399 540 403
rect 552 399 556 403
rect 568 399 572 403
rect 640 399 644 403
rect 688 399 692 403
rect 744 399 748 403
rect 936 399 940 403
rect 944 399 948 403
rect 960 399 964 403
rect 976 399 980 403
rect 1248 399 1252 403
rect 1304 399 1308 403
rect 488 385 492 389
rect 160 379 164 383
rect 880 379 884 383
rect 152 375 156 379
rect 184 375 188 379
rect 216 375 220 379
rect 248 375 252 379
rect 280 375 284 379
rect 288 375 292 379
rect 432 375 436 379
rect 464 375 468 379
rect 520 375 524 379
rect 920 375 924 379
rect 152 359 156 363
rect 184 359 188 363
rect 216 359 220 363
rect 248 359 252 363
rect 280 359 284 363
rect 400 367 404 371
rect 640 367 644 371
rect 432 359 436 363
rect 464 359 468 363
rect 920 359 924 363
rect 880 355 884 359
rect 480 339 484 343
rect 1352 395 1356 399
rect 1368 395 1372 399
rect 1388 395 1392 399
rect 1032 383 1036 387
rect 1200 381 1204 385
rect 1504 379 1508 383
rect 1544 379 1548 383
rect 1064 375 1068 379
rect 1336 375 1340 379
rect 1496 375 1500 379
rect 1536 375 1540 379
rect 1576 375 1580 379
rect 1608 375 1612 379
rect 1640 375 1644 379
rect 1672 375 1676 379
rect 1336 359 1340 363
rect 1496 359 1500 363
rect 1504 359 1508 363
rect 1536 359 1540 363
rect 1544 359 1548 363
rect 1576 359 1580 363
rect 1608 359 1612 363
rect 1640 359 1644 363
rect 1672 359 1676 363
rect 1200 355 1204 359
rect 1456 355 1460 359
rect 1024 339 1028 343
rect 936 319 940 323
rect 1304 295 1308 299
rect 152 291 156 295
rect 184 291 188 295
rect 216 291 220 295
rect 248 291 252 295
rect 280 291 284 295
rect 288 291 292 295
rect 312 291 316 295
rect 344 291 348 295
rect 376 291 380 295
rect 408 291 412 295
rect 440 291 444 295
rect 472 291 476 295
rect 504 291 508 295
rect 536 291 540 295
rect 568 291 572 295
rect 1016 291 1020 295
rect 1048 291 1052 295
rect 1056 291 1060 295
rect 1080 291 1084 295
rect 1336 291 1340 295
rect 1368 291 1372 295
rect 1400 291 1404 295
rect 1432 291 1436 295
rect 1464 291 1468 295
rect 1496 291 1500 295
rect 1536 291 1540 295
rect 1576 291 1580 295
rect 1608 291 1612 295
rect 1640 291 1644 295
rect 1672 291 1676 295
rect 80 279 84 283
rect 152 275 156 279
rect 184 275 188 279
rect 216 275 220 279
rect 248 275 252 279
rect 280 275 284 279
rect 312 275 316 279
rect 344 275 348 279
rect 376 275 380 279
rect 408 275 412 279
rect 440 275 444 279
rect 472 275 476 279
rect 504 275 508 279
rect 536 275 540 279
rect 568 275 572 279
rect 1016 275 1020 279
rect 1048 275 1052 279
rect 616 251 620 255
rect 672 251 676 255
rect 688 251 692 255
rect 720 251 724 255
rect 776 251 780 255
rect 824 251 828 255
rect 880 251 884 255
rect 928 251 932 255
rect 984 251 988 255
rect 1748 287 1752 291
rect 1080 275 1084 279
rect 1336 275 1340 279
rect 1368 275 1372 279
rect 1400 275 1404 279
rect 1432 275 1436 279
rect 1464 275 1468 279
rect 1496 275 1500 279
rect 1536 275 1540 279
rect 1576 275 1580 279
rect 1608 275 1612 279
rect 1640 275 1644 279
rect 1672 275 1676 279
rect 1200 255 1204 259
rect 1216 255 1220 259
rect 1236 255 1240 259
rect 1128 251 1132 255
rect 1184 251 1188 255
rect 712 239 716 243
rect 768 239 772 243
rect 984 239 988 243
rect 1040 239 1044 243
rect 1056 239 1060 243
rect 832 235 836 239
rect 848 235 852 239
rect 868 235 872 239
rect 1328 219 1332 223
rect 1464 219 1468 223
rect 1504 219 1508 223
rect 1544 219 1548 223
rect 200 215 204 219
rect 232 215 236 219
rect 264 215 268 219
rect 296 215 300 219
rect 328 215 332 219
rect 360 215 364 219
rect 392 215 396 219
rect 424 215 428 219
rect 456 215 460 219
rect 488 215 492 219
rect 520 215 524 219
rect 552 215 556 219
rect 584 215 588 219
rect 616 215 620 219
rect 656 215 660 219
rect 808 215 812 219
rect 1080 215 1084 219
rect 1120 215 1124 219
rect 1160 215 1164 219
rect 1200 215 1204 219
rect 1240 215 1244 219
rect 1280 215 1284 219
rect 1320 215 1324 219
rect 200 199 204 203
rect 232 199 236 203
rect 264 199 268 203
rect 296 199 300 203
rect 328 199 332 203
rect 360 199 364 203
rect 392 199 396 203
rect 424 199 428 203
rect 456 199 460 203
rect 488 200 492 204
rect 1360 215 1364 219
rect 1392 215 1396 219
rect 1424 215 1428 219
rect 1456 215 1460 219
rect 1496 215 1500 219
rect 1536 215 1540 219
rect 1576 215 1580 219
rect 1608 215 1612 219
rect 1640 215 1644 219
rect 1672 215 1676 219
rect 520 199 524 203
rect 552 199 556 203
rect 584 199 588 203
rect 616 199 620 203
rect 656 199 660 203
rect 808 199 812 203
rect 1080 199 1084 203
rect 1120 199 1124 203
rect 1160 199 1164 203
rect 1200 199 1204 203
rect 1240 199 1244 203
rect 1280 199 1284 203
rect 1320 199 1324 203
rect 1328 199 1332 203
rect 1360 199 1364 203
rect 1392 199 1396 203
rect 1424 199 1428 203
rect 1456 199 1460 203
rect 1464 199 1468 203
rect 1496 199 1500 203
rect 1504 199 1508 203
rect 1536 199 1540 203
rect 1544 199 1548 203
rect 1576 199 1580 203
rect 1608 199 1612 203
rect 1640 199 1644 203
rect 1672 199 1676 203
rect 936 195 940 199
rect 1200 187 1204 191
rect 152 155 156 159
rect 184 155 188 159
rect 232 155 236 159
rect 280 155 284 159
rect 328 155 332 159
rect 384 155 388 159
rect 432 155 436 159
rect 488 155 492 159
rect 552 155 556 159
rect 624 155 628 159
rect 704 155 708 159
rect 792 155 796 159
rect 880 155 884 159
rect 976 155 980 159
rect 1072 155 1076 159
rect 1168 155 1172 159
rect 152 139 156 143
rect 184 139 188 143
rect 232 139 236 143
rect 280 139 284 143
rect 328 139 332 143
rect 384 139 388 143
rect 432 139 436 143
rect 488 139 492 143
rect 552 139 556 143
rect 624 139 628 143
rect 704 139 708 143
rect 792 139 796 143
rect 880 139 884 143
rect 976 139 980 143
rect 1072 139 1076 143
rect 1168 139 1172 143
rect 576 111 580 115
rect 632 111 636 115
rect 696 111 700 115
rect 768 111 772 115
rect 848 111 852 115
rect 1080 111 1084 115
rect 1144 111 1148 115
rect 152 107 156 111
rect 184 107 188 111
rect 216 107 220 111
rect 248 107 252 111
rect 280 107 284 111
rect 312 107 316 111
rect 344 107 348 111
rect 376 107 380 111
rect 408 107 412 111
rect 440 107 444 111
rect 472 107 476 111
rect 504 107 508 111
rect 536 107 540 111
rect 568 107 572 111
rect 624 107 628 111
rect 688 107 692 111
rect 760 107 764 111
rect 840 107 844 111
rect 920 107 924 111
rect 1000 107 1004 111
rect 1072 107 1076 111
rect 1136 107 1140 111
rect 1192 107 1196 111
rect 152 91 156 95
rect 184 91 188 95
rect 216 91 220 95
rect 248 91 252 95
rect 280 91 284 95
rect 312 91 316 95
rect 344 91 348 95
rect 376 91 380 95
rect 408 91 412 95
rect 440 91 444 95
rect 472 91 476 95
rect 504 91 508 95
rect 536 91 540 95
rect 568 91 572 95
rect 576 91 580 95
rect 624 91 628 95
rect 632 91 636 95
rect 688 91 692 95
rect 696 91 700 95
rect 760 91 764 95
rect 768 91 772 95
rect 840 91 844 95
rect 848 91 852 95
rect 920 91 924 95
rect 1000 91 1004 95
rect 1072 91 1076 95
rect 1080 91 1084 95
rect 1136 91 1140 95
rect 1144 91 1148 95
rect 1192 91 1196 95
rect 1256 155 1260 159
rect 1344 155 1348 159
rect 1432 155 1436 159
rect 1520 155 1524 159
rect 1608 155 1612 159
rect 1672 155 1676 159
rect 1256 139 1260 143
rect 1344 139 1348 143
rect 1432 139 1436 143
rect 1520 139 1524 143
rect 1608 139 1612 143
rect 1672 139 1676 143
rect 1240 107 1244 111
rect 1288 107 1292 111
rect 1328 107 1332 111
rect 1360 107 1364 111
rect 1392 107 1396 111
rect 1424 107 1428 111
rect 1456 107 1460 111
rect 1496 107 1500 111
rect 1536 107 1540 111
rect 1576 107 1580 111
rect 1608 107 1612 111
rect 1640 107 1644 111
rect 1672 107 1676 111
rect 1240 91 1244 95
rect 1288 91 1292 95
rect 1328 91 1332 95
rect 1360 91 1364 95
rect 1392 91 1396 95
rect 1424 91 1428 95
rect 1456 91 1460 95
rect 1496 91 1500 95
rect 1536 91 1540 95
rect 1576 91 1580 95
rect 1608 91 1612 95
rect 1640 91 1644 95
rect 1672 91 1676 95
rect 638 83 642 87
<< m2 >>
rect 637 1763 643 1764
rect 637 1759 638 1763
rect 642 1762 643 1763
rect 870 1763 876 1764
rect 870 1762 871 1763
rect 642 1760 871 1762
rect 642 1759 643 1760
rect 637 1758 643 1759
rect 870 1759 871 1760
rect 875 1759 876 1763
rect 870 1758 876 1759
rect 1189 1759 1196 1760
rect 150 1755 156 1756
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 150 1751 151 1755
rect 155 1751 156 1755
rect 150 1750 156 1751
rect 182 1755 188 1756
rect 182 1751 183 1755
rect 187 1751 188 1755
rect 182 1750 188 1751
rect 214 1755 220 1756
rect 214 1751 215 1755
rect 219 1751 220 1755
rect 214 1750 220 1751
rect 246 1755 252 1756
rect 246 1751 247 1755
rect 251 1751 252 1755
rect 246 1750 252 1751
rect 278 1755 284 1756
rect 278 1751 279 1755
rect 283 1751 284 1755
rect 278 1750 284 1751
rect 310 1755 316 1756
rect 310 1751 311 1755
rect 315 1751 316 1755
rect 310 1750 316 1751
rect 342 1755 348 1756
rect 342 1751 343 1755
rect 347 1751 348 1755
rect 342 1750 348 1751
rect 374 1755 380 1756
rect 374 1751 375 1755
rect 379 1751 380 1755
rect 374 1750 380 1751
rect 406 1755 412 1756
rect 406 1751 407 1755
rect 411 1751 412 1755
rect 406 1750 412 1751
rect 438 1755 444 1756
rect 438 1751 439 1755
rect 443 1751 444 1755
rect 438 1750 444 1751
rect 470 1755 476 1756
rect 470 1751 471 1755
rect 475 1751 476 1755
rect 470 1750 476 1751
rect 502 1755 508 1756
rect 502 1751 503 1755
rect 507 1751 508 1755
rect 502 1750 508 1751
rect 534 1755 540 1756
rect 534 1751 535 1755
rect 539 1751 540 1755
rect 534 1750 540 1751
rect 566 1755 572 1756
rect 566 1751 567 1755
rect 571 1751 572 1755
rect 566 1750 572 1751
rect 598 1755 604 1756
rect 598 1751 599 1755
rect 603 1751 604 1755
rect 598 1750 604 1751
rect 630 1755 636 1756
rect 630 1751 631 1755
rect 635 1751 636 1755
rect 630 1750 636 1751
rect 662 1755 668 1756
rect 662 1751 663 1755
rect 667 1751 668 1755
rect 662 1750 668 1751
rect 694 1755 700 1756
rect 694 1751 695 1755
rect 699 1751 700 1755
rect 694 1750 700 1751
rect 726 1755 732 1756
rect 726 1751 727 1755
rect 731 1751 732 1755
rect 726 1750 732 1751
rect 758 1755 764 1756
rect 758 1751 759 1755
rect 763 1751 764 1755
rect 758 1750 764 1751
rect 790 1755 796 1756
rect 790 1751 791 1755
rect 795 1751 796 1755
rect 790 1750 796 1751
rect 822 1755 828 1756
rect 822 1751 823 1755
rect 827 1751 828 1755
rect 822 1750 828 1751
rect 854 1755 860 1756
rect 854 1751 855 1755
rect 859 1751 860 1755
rect 854 1750 860 1751
rect 886 1755 892 1756
rect 886 1751 887 1755
rect 891 1751 892 1755
rect 886 1750 892 1751
rect 918 1755 924 1756
rect 918 1751 919 1755
rect 923 1751 924 1755
rect 918 1750 924 1751
rect 950 1755 956 1756
rect 950 1751 951 1755
rect 955 1751 956 1755
rect 950 1750 956 1751
rect 982 1755 988 1756
rect 982 1751 983 1755
rect 987 1751 988 1755
rect 1189 1755 1190 1759
rect 1195 1755 1196 1759
rect 1189 1754 1196 1755
rect 982 1750 988 1751
rect 1694 1753 1700 1754
rect 110 1748 116 1749
rect 1694 1749 1695 1753
rect 1699 1749 1700 1753
rect 1694 1748 1700 1749
rect 167 1747 173 1748
rect 167 1743 168 1747
rect 172 1746 173 1747
rect 199 1747 205 1748
rect 172 1744 194 1746
rect 172 1743 173 1744
rect 167 1742 173 1743
rect 150 1738 156 1739
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 150 1734 151 1738
rect 155 1734 156 1738
rect 150 1733 156 1734
rect 182 1738 188 1739
rect 182 1734 183 1738
rect 187 1734 188 1738
rect 182 1733 188 1734
rect 110 1731 116 1732
rect 167 1731 173 1732
rect 167 1727 168 1731
rect 172 1730 173 1731
rect 192 1730 194 1744
rect 199 1743 200 1747
rect 204 1746 205 1747
rect 231 1747 237 1748
rect 204 1744 226 1746
rect 204 1743 205 1744
rect 199 1742 205 1743
rect 214 1738 220 1739
rect 214 1734 215 1738
rect 219 1734 220 1738
rect 214 1733 220 1734
rect 199 1731 205 1732
rect 199 1730 200 1731
rect 172 1728 190 1730
rect 192 1728 200 1730
rect 172 1727 173 1728
rect 167 1726 173 1727
rect 188 1722 190 1728
rect 199 1727 200 1728
rect 204 1727 205 1731
rect 224 1730 226 1744
rect 231 1743 232 1747
rect 236 1743 237 1747
rect 231 1742 237 1743
rect 239 1747 245 1748
rect 239 1743 240 1747
rect 244 1746 245 1747
rect 263 1747 269 1748
rect 263 1746 264 1747
rect 244 1744 264 1746
rect 244 1743 245 1744
rect 239 1742 245 1743
rect 263 1743 264 1744
rect 268 1743 269 1747
rect 295 1747 301 1748
rect 295 1746 296 1747
rect 263 1742 269 1743
rect 288 1744 296 1746
rect 232 1738 234 1742
rect 246 1738 252 1739
rect 232 1736 242 1738
rect 231 1731 237 1732
rect 231 1730 232 1731
rect 224 1728 232 1730
rect 199 1726 205 1727
rect 231 1727 232 1728
rect 236 1727 237 1731
rect 240 1730 242 1736
rect 246 1734 247 1738
rect 251 1734 252 1738
rect 246 1733 252 1734
rect 278 1738 284 1739
rect 278 1734 279 1738
rect 283 1734 284 1738
rect 278 1733 284 1734
rect 263 1731 269 1732
rect 240 1728 258 1730
rect 231 1726 237 1727
rect 239 1723 245 1724
rect 239 1722 240 1723
rect 188 1720 240 1722
rect 239 1719 240 1720
rect 244 1719 245 1723
rect 239 1718 245 1719
rect 256 1718 258 1728
rect 263 1727 264 1731
rect 268 1730 269 1731
rect 288 1730 290 1744
rect 295 1743 296 1744
rect 300 1743 301 1747
rect 327 1747 333 1748
rect 327 1746 328 1747
rect 295 1742 301 1743
rect 320 1744 328 1746
rect 310 1738 316 1739
rect 310 1734 311 1738
rect 315 1734 316 1738
rect 310 1733 316 1734
rect 268 1728 290 1730
rect 295 1731 301 1732
rect 268 1727 269 1728
rect 263 1726 269 1727
rect 295 1727 296 1731
rect 300 1730 301 1731
rect 320 1730 322 1744
rect 327 1743 328 1744
rect 332 1743 333 1747
rect 359 1747 365 1748
rect 359 1746 360 1747
rect 327 1742 333 1743
rect 352 1744 360 1746
rect 342 1738 348 1739
rect 342 1734 343 1738
rect 347 1734 348 1738
rect 342 1733 348 1734
rect 300 1728 322 1730
rect 327 1731 333 1732
rect 300 1727 301 1728
rect 295 1726 301 1727
rect 327 1727 328 1731
rect 332 1730 333 1731
rect 352 1730 354 1744
rect 359 1743 360 1744
rect 364 1743 365 1747
rect 391 1747 397 1748
rect 391 1746 392 1747
rect 359 1742 365 1743
rect 384 1744 392 1746
rect 374 1738 380 1739
rect 374 1734 375 1738
rect 379 1734 380 1738
rect 374 1733 380 1734
rect 332 1728 354 1730
rect 359 1731 365 1732
rect 332 1727 333 1728
rect 327 1726 333 1727
rect 359 1727 360 1731
rect 364 1730 365 1731
rect 384 1730 386 1744
rect 391 1743 392 1744
rect 396 1743 397 1747
rect 423 1747 429 1748
rect 423 1746 424 1747
rect 391 1742 397 1743
rect 416 1744 424 1746
rect 406 1738 412 1739
rect 406 1734 407 1738
rect 411 1734 412 1738
rect 406 1733 412 1734
rect 364 1728 386 1730
rect 391 1731 397 1732
rect 364 1727 365 1728
rect 359 1726 365 1727
rect 391 1727 392 1731
rect 396 1730 397 1731
rect 416 1730 418 1744
rect 423 1743 424 1744
rect 428 1743 429 1747
rect 455 1747 461 1748
rect 455 1746 456 1747
rect 423 1742 429 1743
rect 448 1744 456 1746
rect 438 1738 444 1739
rect 438 1734 439 1738
rect 443 1734 444 1738
rect 438 1733 444 1734
rect 396 1728 418 1730
rect 423 1731 429 1732
rect 396 1727 397 1728
rect 391 1726 397 1727
rect 423 1727 424 1731
rect 428 1730 429 1731
rect 448 1730 450 1744
rect 455 1743 456 1744
rect 460 1743 461 1747
rect 487 1747 493 1748
rect 487 1746 488 1747
rect 455 1742 461 1743
rect 480 1744 488 1746
rect 470 1738 476 1739
rect 470 1734 471 1738
rect 475 1734 476 1738
rect 470 1733 476 1734
rect 428 1728 450 1730
rect 455 1731 461 1732
rect 428 1727 429 1728
rect 423 1726 429 1727
rect 455 1727 456 1731
rect 460 1730 461 1731
rect 480 1730 482 1744
rect 487 1743 488 1744
rect 492 1743 493 1747
rect 519 1747 525 1748
rect 519 1746 520 1747
rect 487 1742 493 1743
rect 512 1744 520 1746
rect 502 1738 508 1739
rect 502 1734 503 1738
rect 507 1734 508 1738
rect 502 1733 508 1734
rect 460 1728 482 1730
rect 487 1731 493 1732
rect 460 1727 461 1728
rect 455 1726 461 1727
rect 487 1727 488 1731
rect 492 1730 493 1731
rect 512 1730 514 1744
rect 519 1743 520 1744
rect 524 1743 525 1747
rect 551 1747 557 1748
rect 551 1746 552 1747
rect 519 1742 525 1743
rect 544 1744 552 1746
rect 534 1738 540 1739
rect 534 1734 535 1738
rect 539 1734 540 1738
rect 534 1733 540 1734
rect 492 1728 514 1730
rect 519 1731 525 1732
rect 492 1727 493 1728
rect 487 1726 493 1727
rect 519 1727 520 1731
rect 524 1730 525 1731
rect 544 1730 546 1744
rect 551 1743 552 1744
rect 556 1743 557 1747
rect 583 1747 589 1748
rect 583 1746 584 1747
rect 551 1742 557 1743
rect 576 1744 584 1746
rect 566 1738 572 1739
rect 566 1734 567 1738
rect 571 1734 572 1738
rect 566 1733 572 1734
rect 524 1728 546 1730
rect 551 1731 557 1732
rect 524 1727 525 1728
rect 519 1726 525 1727
rect 551 1727 552 1731
rect 556 1730 557 1731
rect 576 1730 578 1744
rect 583 1743 584 1744
rect 588 1743 589 1747
rect 615 1747 621 1748
rect 615 1746 616 1747
rect 583 1742 589 1743
rect 608 1744 616 1746
rect 598 1738 604 1739
rect 598 1734 599 1738
rect 603 1734 604 1738
rect 598 1733 604 1734
rect 556 1728 578 1730
rect 583 1731 589 1732
rect 556 1727 557 1728
rect 551 1726 557 1727
rect 583 1727 584 1731
rect 588 1730 589 1731
rect 608 1730 610 1744
rect 615 1743 616 1744
rect 620 1743 621 1747
rect 647 1747 653 1748
rect 647 1746 648 1747
rect 615 1742 621 1743
rect 640 1744 648 1746
rect 630 1738 636 1739
rect 630 1734 631 1738
rect 635 1734 636 1738
rect 630 1733 636 1734
rect 588 1728 610 1730
rect 615 1731 621 1732
rect 588 1727 589 1728
rect 583 1726 589 1727
rect 615 1727 616 1731
rect 620 1730 621 1731
rect 640 1730 642 1744
rect 647 1743 648 1744
rect 652 1743 653 1747
rect 679 1747 685 1748
rect 679 1746 680 1747
rect 647 1742 653 1743
rect 656 1744 680 1746
rect 620 1728 642 1730
rect 647 1731 653 1732
rect 620 1727 621 1728
rect 615 1726 621 1727
rect 647 1727 648 1731
rect 652 1730 653 1731
rect 656 1730 658 1744
rect 679 1743 680 1744
rect 684 1743 685 1747
rect 711 1747 717 1748
rect 711 1746 712 1747
rect 679 1742 685 1743
rect 704 1744 712 1746
rect 662 1738 668 1739
rect 662 1734 663 1738
rect 667 1734 668 1738
rect 662 1733 668 1734
rect 694 1738 700 1739
rect 694 1734 695 1738
rect 699 1734 700 1738
rect 694 1733 700 1734
rect 652 1728 658 1730
rect 679 1731 685 1732
rect 652 1727 653 1728
rect 647 1726 653 1727
rect 679 1727 680 1731
rect 684 1730 685 1731
rect 704 1730 706 1744
rect 711 1743 712 1744
rect 716 1743 717 1747
rect 743 1747 749 1748
rect 743 1746 744 1747
rect 711 1742 717 1743
rect 736 1744 744 1746
rect 726 1738 732 1739
rect 726 1734 727 1738
rect 731 1734 732 1738
rect 726 1733 732 1734
rect 684 1728 706 1730
rect 711 1731 717 1732
rect 684 1727 685 1728
rect 679 1726 685 1727
rect 711 1727 712 1731
rect 716 1730 717 1731
rect 736 1730 738 1744
rect 743 1743 744 1744
rect 748 1743 749 1747
rect 775 1747 781 1748
rect 775 1746 776 1747
rect 743 1742 749 1743
rect 768 1744 776 1746
rect 758 1738 764 1739
rect 758 1734 759 1738
rect 763 1734 764 1738
rect 758 1733 764 1734
rect 716 1728 738 1730
rect 743 1731 749 1732
rect 716 1727 717 1728
rect 711 1726 717 1727
rect 743 1727 744 1731
rect 748 1730 749 1731
rect 768 1730 770 1744
rect 775 1743 776 1744
rect 780 1743 781 1747
rect 807 1747 813 1748
rect 807 1746 808 1747
rect 775 1742 781 1743
rect 800 1744 808 1746
rect 790 1738 796 1739
rect 790 1734 791 1738
rect 795 1734 796 1738
rect 790 1733 796 1734
rect 748 1728 770 1730
rect 775 1731 781 1732
rect 748 1727 749 1728
rect 743 1726 749 1727
rect 775 1727 776 1731
rect 780 1730 781 1731
rect 800 1730 802 1744
rect 807 1743 808 1744
rect 812 1743 813 1747
rect 839 1747 845 1748
rect 839 1746 840 1747
rect 807 1742 813 1743
rect 832 1744 840 1746
rect 822 1738 828 1739
rect 822 1734 823 1738
rect 827 1734 828 1738
rect 822 1733 828 1734
rect 780 1728 802 1730
rect 807 1731 813 1732
rect 780 1727 781 1728
rect 775 1726 781 1727
rect 807 1727 808 1731
rect 812 1730 813 1731
rect 832 1730 834 1744
rect 839 1743 840 1744
rect 844 1743 845 1747
rect 871 1747 877 1748
rect 871 1746 872 1747
rect 839 1742 845 1743
rect 864 1744 872 1746
rect 854 1738 860 1739
rect 854 1734 855 1738
rect 859 1734 860 1738
rect 854 1733 860 1734
rect 812 1728 834 1730
rect 839 1731 845 1732
rect 812 1727 813 1728
rect 807 1726 813 1727
rect 839 1727 840 1731
rect 844 1730 845 1731
rect 864 1730 866 1744
rect 871 1743 872 1744
rect 876 1743 877 1747
rect 903 1747 909 1748
rect 903 1746 904 1747
rect 871 1742 877 1743
rect 896 1744 904 1746
rect 886 1738 892 1739
rect 886 1734 887 1738
rect 891 1734 892 1738
rect 886 1733 892 1734
rect 844 1728 866 1730
rect 871 1731 877 1732
rect 844 1727 845 1728
rect 839 1726 845 1727
rect 871 1727 872 1731
rect 876 1730 877 1731
rect 896 1730 898 1744
rect 903 1743 904 1744
rect 908 1743 909 1747
rect 935 1747 941 1748
rect 935 1746 936 1747
rect 903 1742 909 1743
rect 928 1744 936 1746
rect 918 1738 924 1739
rect 918 1734 919 1738
rect 923 1734 924 1738
rect 918 1733 924 1734
rect 876 1728 898 1730
rect 903 1731 909 1732
rect 876 1727 877 1728
rect 871 1726 877 1727
rect 903 1727 904 1731
rect 908 1730 909 1731
rect 928 1730 930 1744
rect 935 1743 936 1744
rect 940 1743 941 1747
rect 967 1747 973 1748
rect 967 1746 968 1747
rect 935 1742 941 1743
rect 960 1744 968 1746
rect 950 1738 956 1739
rect 950 1734 951 1738
rect 955 1734 956 1738
rect 950 1733 956 1734
rect 908 1728 930 1730
rect 935 1731 941 1732
rect 908 1727 909 1728
rect 903 1726 909 1727
rect 935 1727 936 1731
rect 940 1730 941 1731
rect 960 1730 962 1744
rect 967 1743 968 1744
rect 972 1743 973 1747
rect 999 1747 1005 1748
rect 999 1746 1000 1747
rect 967 1742 973 1743
rect 992 1744 1000 1746
rect 982 1738 988 1739
rect 982 1734 983 1738
rect 987 1734 988 1738
rect 982 1733 988 1734
rect 940 1728 962 1730
rect 967 1731 973 1732
rect 940 1727 941 1728
rect 935 1726 941 1727
rect 967 1727 968 1731
rect 972 1730 973 1731
rect 992 1730 994 1744
rect 999 1743 1000 1744
rect 1004 1743 1005 1747
rect 999 1742 1005 1743
rect 1694 1736 1700 1737
rect 1694 1732 1695 1736
rect 1699 1732 1700 1736
rect 972 1728 994 1730
rect 999 1731 1005 1732
rect 972 1727 973 1728
rect 967 1726 973 1727
rect 999 1727 1000 1731
rect 1004 1730 1005 1731
rect 1062 1731 1068 1732
rect 1694 1731 1700 1732
rect 1062 1730 1063 1731
rect 1004 1728 1063 1730
rect 1004 1727 1005 1728
rect 999 1726 1005 1727
rect 1062 1727 1063 1728
rect 1067 1727 1068 1731
rect 1062 1726 1068 1727
rect 256 1716 426 1718
rect 215 1711 221 1712
rect 206 1707 213 1708
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 206 1703 207 1707
rect 212 1703 213 1707
rect 215 1707 216 1711
rect 220 1710 221 1711
rect 271 1711 277 1712
rect 220 1708 258 1710
rect 220 1707 221 1708
rect 215 1706 221 1707
rect 256 1706 258 1708
rect 263 1707 269 1708
rect 263 1706 264 1707
rect 256 1704 264 1706
rect 263 1703 264 1704
rect 268 1703 269 1707
rect 271 1707 272 1711
rect 276 1710 277 1711
rect 276 1708 330 1710
rect 276 1707 277 1708
rect 271 1706 277 1707
rect 328 1706 330 1708
rect 335 1707 341 1708
rect 335 1706 336 1707
rect 328 1704 336 1706
rect 335 1703 336 1704
rect 340 1703 341 1707
rect 424 1706 426 1716
rect 439 1711 445 1712
rect 431 1707 437 1708
rect 431 1706 432 1707
rect 424 1704 432 1706
rect 431 1703 432 1704
rect 436 1703 437 1707
rect 439 1707 440 1711
rect 444 1710 445 1711
rect 551 1711 557 1712
rect 444 1708 547 1710
rect 444 1707 445 1708
rect 439 1706 445 1707
rect 543 1707 549 1708
rect 543 1703 544 1707
rect 548 1703 549 1707
rect 551 1707 552 1711
rect 556 1710 557 1711
rect 902 1711 908 1712
rect 556 1708 675 1710
rect 556 1707 557 1708
rect 551 1706 557 1707
rect 671 1707 677 1708
rect 671 1703 672 1707
rect 676 1703 677 1707
rect 807 1707 813 1708
rect 807 1703 808 1707
rect 812 1706 813 1707
rect 894 1707 900 1708
rect 894 1706 895 1707
rect 812 1704 895 1706
rect 812 1703 813 1704
rect 110 1699 116 1700
rect 190 1702 196 1703
rect 206 1702 213 1703
rect 246 1702 252 1703
rect 263 1702 269 1703
rect 318 1702 324 1703
rect 335 1702 341 1703
rect 414 1702 420 1703
rect 431 1702 437 1703
rect 526 1702 532 1703
rect 543 1702 549 1703
rect 654 1702 660 1703
rect 671 1702 677 1703
rect 790 1702 796 1703
rect 807 1702 813 1703
rect 894 1703 895 1704
rect 899 1703 900 1707
rect 902 1707 903 1711
rect 907 1710 908 1711
rect 943 1711 949 1712
rect 907 1708 930 1710
rect 907 1707 908 1708
rect 902 1706 908 1707
rect 928 1706 930 1708
rect 935 1707 941 1708
rect 935 1706 936 1707
rect 928 1704 936 1706
rect 935 1703 936 1704
rect 940 1703 941 1707
rect 943 1707 944 1711
rect 948 1710 949 1711
rect 1206 1711 1212 1712
rect 948 1708 1058 1710
rect 948 1707 949 1708
rect 943 1706 949 1707
rect 1056 1706 1058 1708
rect 1063 1707 1069 1708
rect 1063 1706 1064 1707
rect 1056 1704 1064 1706
rect 1063 1703 1064 1704
rect 1068 1703 1069 1707
rect 1175 1707 1181 1708
rect 1175 1703 1176 1707
rect 1180 1706 1181 1707
rect 1198 1707 1204 1708
rect 1198 1706 1199 1707
rect 1180 1704 1199 1706
rect 1180 1703 1181 1704
rect 894 1702 900 1703
rect 918 1702 924 1703
rect 935 1702 941 1703
rect 1046 1702 1052 1703
rect 1063 1702 1069 1703
rect 1158 1702 1164 1703
rect 1175 1702 1181 1703
rect 1198 1703 1199 1704
rect 1203 1703 1204 1707
rect 1206 1707 1207 1711
rect 1211 1710 1212 1711
rect 1279 1711 1285 1712
rect 1211 1708 1275 1710
rect 1211 1707 1212 1708
rect 1206 1706 1212 1707
rect 1271 1707 1277 1708
rect 1271 1703 1272 1707
rect 1276 1703 1277 1707
rect 1279 1707 1280 1711
rect 1284 1710 1285 1711
rect 1359 1711 1365 1712
rect 1284 1708 1355 1710
rect 1284 1707 1285 1708
rect 1279 1706 1285 1707
rect 1351 1707 1357 1708
rect 1351 1703 1352 1707
rect 1356 1703 1357 1707
rect 1359 1707 1360 1711
rect 1364 1710 1365 1711
rect 1431 1711 1437 1712
rect 1364 1708 1418 1710
rect 1364 1707 1365 1708
rect 1359 1706 1365 1707
rect 1416 1706 1418 1708
rect 1423 1707 1429 1708
rect 1423 1706 1424 1707
rect 1416 1704 1424 1706
rect 1423 1703 1424 1704
rect 1428 1703 1429 1707
rect 1431 1707 1432 1711
rect 1436 1710 1437 1711
rect 1487 1711 1493 1712
rect 1436 1708 1474 1710
rect 1436 1707 1437 1708
rect 1431 1706 1437 1707
rect 1472 1706 1474 1708
rect 1479 1707 1485 1708
rect 1479 1706 1480 1707
rect 1472 1704 1480 1706
rect 1479 1703 1480 1704
rect 1484 1703 1485 1707
rect 1487 1707 1488 1711
rect 1492 1710 1493 1711
rect 1543 1711 1549 1712
rect 1492 1708 1530 1710
rect 1492 1707 1493 1708
rect 1487 1706 1493 1707
rect 1528 1706 1530 1708
rect 1535 1707 1541 1708
rect 1535 1706 1536 1707
rect 1528 1704 1536 1706
rect 1535 1703 1536 1704
rect 1540 1703 1541 1707
rect 1543 1707 1544 1711
rect 1548 1710 1549 1711
rect 1591 1711 1597 1712
rect 1548 1708 1587 1710
rect 1548 1707 1549 1708
rect 1543 1706 1549 1707
rect 1583 1707 1589 1708
rect 1583 1703 1584 1707
rect 1588 1703 1589 1707
rect 1591 1707 1592 1711
rect 1596 1710 1597 1711
rect 1596 1708 1634 1710
rect 1596 1707 1597 1708
rect 1591 1706 1597 1707
rect 1632 1706 1634 1708
rect 1639 1707 1645 1708
rect 1639 1706 1640 1707
rect 1632 1704 1640 1706
rect 1639 1703 1640 1704
rect 1644 1703 1645 1707
rect 1671 1707 1677 1708
rect 1671 1706 1672 1707
rect 1664 1704 1672 1706
rect 1198 1702 1204 1703
rect 1254 1702 1260 1703
rect 1271 1702 1277 1703
rect 1334 1702 1340 1703
rect 1351 1702 1357 1703
rect 1406 1702 1412 1703
rect 1423 1702 1429 1703
rect 1462 1702 1468 1703
rect 1479 1702 1485 1703
rect 1518 1702 1524 1703
rect 1535 1702 1541 1703
rect 1566 1702 1572 1703
rect 1583 1702 1589 1703
rect 1622 1702 1628 1703
rect 1639 1702 1645 1703
rect 1654 1702 1660 1703
rect 190 1698 191 1702
rect 195 1698 196 1702
rect 190 1697 196 1698
rect 246 1698 247 1702
rect 251 1698 252 1702
rect 246 1697 252 1698
rect 318 1698 319 1702
rect 323 1698 324 1702
rect 318 1697 324 1698
rect 414 1698 415 1702
rect 419 1698 420 1702
rect 414 1697 420 1698
rect 526 1698 527 1702
rect 531 1698 532 1702
rect 526 1697 532 1698
rect 654 1698 655 1702
rect 659 1698 660 1702
rect 654 1697 660 1698
rect 790 1698 791 1702
rect 795 1698 796 1702
rect 790 1697 796 1698
rect 918 1698 919 1702
rect 923 1698 924 1702
rect 918 1697 924 1698
rect 1046 1698 1047 1702
rect 1051 1698 1052 1702
rect 1046 1697 1052 1698
rect 1158 1698 1159 1702
rect 1163 1698 1164 1702
rect 1158 1697 1164 1698
rect 1254 1698 1255 1702
rect 1259 1698 1260 1702
rect 1254 1697 1260 1698
rect 1334 1698 1335 1702
rect 1339 1698 1340 1702
rect 1334 1697 1340 1698
rect 1406 1698 1407 1702
rect 1411 1698 1412 1702
rect 1406 1697 1412 1698
rect 1462 1698 1463 1702
rect 1467 1698 1468 1702
rect 1462 1697 1468 1698
rect 1518 1698 1519 1702
rect 1523 1698 1524 1702
rect 1518 1697 1524 1698
rect 1566 1698 1567 1702
rect 1571 1698 1572 1702
rect 1566 1697 1572 1698
rect 1622 1698 1623 1702
rect 1627 1698 1628 1702
rect 1622 1697 1628 1698
rect 1654 1698 1655 1702
rect 1659 1698 1660 1702
rect 1654 1697 1660 1698
rect 1664 1692 1666 1704
rect 1671 1703 1672 1704
rect 1676 1703 1677 1707
rect 1671 1702 1677 1703
rect 1694 1704 1700 1705
rect 1694 1700 1695 1704
rect 1699 1700 1700 1704
rect 1694 1699 1700 1700
rect 207 1691 213 1692
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 207 1687 208 1691
rect 212 1690 213 1691
rect 215 1691 221 1692
rect 215 1690 216 1691
rect 212 1688 216 1690
rect 212 1687 213 1688
rect 207 1686 213 1687
rect 215 1687 216 1688
rect 220 1687 221 1691
rect 215 1686 221 1687
rect 263 1691 269 1692
rect 263 1687 264 1691
rect 268 1690 269 1691
rect 271 1691 277 1692
rect 271 1690 272 1691
rect 268 1688 272 1690
rect 268 1687 269 1688
rect 263 1686 269 1687
rect 271 1687 272 1688
rect 276 1687 277 1691
rect 271 1686 277 1687
rect 335 1691 341 1692
rect 335 1687 336 1691
rect 340 1690 341 1691
rect 406 1691 412 1692
rect 406 1690 407 1691
rect 340 1688 407 1690
rect 340 1687 341 1688
rect 335 1686 341 1687
rect 406 1687 407 1688
rect 411 1687 412 1691
rect 406 1686 412 1687
rect 431 1691 437 1692
rect 431 1687 432 1691
rect 436 1690 437 1691
rect 439 1691 445 1692
rect 439 1690 440 1691
rect 436 1688 440 1690
rect 436 1687 437 1688
rect 431 1686 437 1687
rect 439 1687 440 1688
rect 444 1687 445 1691
rect 439 1686 445 1687
rect 543 1691 549 1692
rect 543 1687 544 1691
rect 548 1690 549 1691
rect 551 1691 557 1692
rect 551 1690 552 1691
rect 548 1688 552 1690
rect 548 1687 549 1688
rect 543 1686 549 1687
rect 551 1687 552 1688
rect 556 1687 557 1691
rect 551 1686 557 1687
rect 671 1691 677 1692
rect 671 1687 672 1691
rect 676 1687 677 1691
rect 671 1686 677 1687
rect 807 1691 813 1692
rect 807 1687 808 1691
rect 812 1690 813 1691
rect 902 1691 908 1692
rect 902 1690 903 1691
rect 812 1688 903 1690
rect 812 1687 813 1688
rect 807 1686 813 1687
rect 902 1687 903 1688
rect 907 1687 908 1691
rect 902 1686 908 1687
rect 935 1691 941 1692
rect 935 1687 936 1691
rect 940 1690 941 1691
rect 943 1691 949 1692
rect 943 1690 944 1691
rect 940 1688 944 1690
rect 940 1687 941 1688
rect 935 1686 941 1687
rect 943 1687 944 1688
rect 948 1687 949 1691
rect 943 1686 949 1687
rect 1062 1691 1069 1692
rect 1062 1687 1063 1691
rect 1068 1687 1069 1691
rect 1062 1686 1069 1687
rect 1175 1691 1181 1692
rect 1175 1687 1176 1691
rect 1180 1690 1181 1691
rect 1206 1691 1212 1692
rect 1206 1690 1207 1691
rect 1180 1688 1207 1690
rect 1180 1687 1181 1688
rect 1175 1686 1181 1687
rect 1206 1687 1207 1688
rect 1211 1687 1212 1691
rect 1206 1686 1212 1687
rect 1271 1691 1277 1692
rect 1271 1687 1272 1691
rect 1276 1690 1277 1691
rect 1279 1691 1285 1692
rect 1279 1690 1280 1691
rect 1276 1688 1280 1690
rect 1276 1687 1277 1688
rect 1271 1686 1277 1687
rect 1279 1687 1280 1688
rect 1284 1687 1285 1691
rect 1279 1686 1285 1687
rect 1351 1691 1357 1692
rect 1351 1687 1352 1691
rect 1356 1690 1357 1691
rect 1359 1691 1365 1692
rect 1359 1690 1360 1691
rect 1356 1688 1360 1690
rect 1356 1687 1357 1688
rect 1351 1686 1357 1687
rect 1359 1687 1360 1688
rect 1364 1687 1365 1691
rect 1359 1686 1365 1687
rect 1423 1691 1429 1692
rect 1423 1687 1424 1691
rect 1428 1690 1429 1691
rect 1431 1691 1437 1692
rect 1431 1690 1432 1691
rect 1428 1688 1432 1690
rect 1428 1687 1429 1688
rect 1423 1686 1429 1687
rect 1431 1687 1432 1688
rect 1436 1687 1437 1691
rect 1431 1686 1437 1687
rect 1479 1691 1485 1692
rect 1479 1687 1480 1691
rect 1484 1690 1485 1691
rect 1487 1691 1493 1692
rect 1487 1690 1488 1691
rect 1484 1688 1488 1690
rect 1484 1687 1485 1688
rect 1479 1686 1485 1687
rect 1487 1687 1488 1688
rect 1492 1687 1493 1691
rect 1487 1686 1493 1687
rect 1535 1691 1541 1692
rect 1535 1687 1536 1691
rect 1540 1690 1541 1691
rect 1543 1691 1549 1692
rect 1543 1690 1544 1691
rect 1540 1688 1544 1690
rect 1540 1687 1541 1688
rect 1535 1686 1541 1687
rect 1543 1687 1544 1688
rect 1548 1687 1549 1691
rect 1543 1686 1549 1687
rect 1583 1691 1589 1692
rect 1583 1687 1584 1691
rect 1588 1690 1589 1691
rect 1591 1691 1597 1692
rect 1591 1690 1592 1691
rect 1588 1688 1592 1690
rect 1588 1687 1589 1688
rect 1583 1686 1589 1687
rect 1591 1687 1592 1688
rect 1596 1687 1597 1691
rect 1591 1686 1597 1687
rect 1639 1691 1645 1692
rect 1639 1687 1640 1691
rect 1644 1690 1645 1691
rect 1652 1690 1666 1692
rect 1671 1691 1677 1692
rect 1644 1688 1654 1690
rect 1644 1687 1645 1688
rect 1639 1686 1645 1687
rect 1671 1687 1672 1691
rect 1676 1687 1677 1691
rect 1671 1686 1677 1687
rect 1694 1687 1700 1688
rect 110 1682 116 1683
rect 190 1685 196 1686
rect 190 1681 191 1685
rect 195 1681 196 1685
rect 190 1680 196 1681
rect 246 1685 252 1686
rect 246 1681 247 1685
rect 251 1681 252 1685
rect 246 1680 252 1681
rect 318 1685 324 1686
rect 318 1681 319 1685
rect 323 1681 324 1685
rect 318 1680 324 1681
rect 414 1685 420 1686
rect 414 1681 415 1685
rect 419 1681 420 1685
rect 414 1680 420 1681
rect 526 1685 532 1686
rect 526 1681 527 1685
rect 531 1681 532 1685
rect 526 1680 532 1681
rect 654 1685 660 1686
rect 654 1681 655 1685
rect 659 1681 660 1685
rect 654 1680 660 1681
rect 206 1679 212 1680
rect 206 1675 207 1679
rect 211 1678 212 1679
rect 673 1678 675 1686
rect 790 1685 796 1686
rect 790 1681 791 1685
rect 795 1681 796 1685
rect 790 1680 796 1681
rect 918 1685 924 1686
rect 918 1681 919 1685
rect 923 1681 924 1685
rect 918 1680 924 1681
rect 1046 1685 1052 1686
rect 1046 1681 1047 1685
rect 1051 1681 1052 1685
rect 1046 1680 1052 1681
rect 1158 1685 1164 1686
rect 1158 1681 1159 1685
rect 1163 1681 1164 1685
rect 1158 1680 1164 1681
rect 1254 1685 1260 1686
rect 1254 1681 1255 1685
rect 1259 1681 1260 1685
rect 1254 1680 1260 1681
rect 1334 1685 1340 1686
rect 1334 1681 1335 1685
rect 1339 1681 1340 1685
rect 1334 1680 1340 1681
rect 1406 1685 1412 1686
rect 1406 1681 1407 1685
rect 1411 1681 1412 1685
rect 1406 1680 1412 1681
rect 1462 1685 1468 1686
rect 1462 1681 1463 1685
rect 1467 1681 1468 1685
rect 1462 1680 1468 1681
rect 1518 1685 1524 1686
rect 1518 1681 1519 1685
rect 1523 1681 1524 1685
rect 1518 1680 1524 1681
rect 1566 1685 1572 1686
rect 1566 1681 1567 1685
rect 1571 1681 1572 1685
rect 1566 1680 1572 1681
rect 1622 1685 1628 1686
rect 1622 1681 1623 1685
rect 1627 1681 1628 1685
rect 1622 1680 1628 1681
rect 1654 1685 1660 1686
rect 1654 1681 1655 1685
rect 1659 1681 1660 1685
rect 1654 1680 1660 1681
rect 211 1676 675 1678
rect 1470 1679 1476 1680
rect 211 1675 212 1676
rect 206 1674 212 1675
rect 1470 1675 1471 1679
rect 1475 1678 1476 1679
rect 1672 1678 1674 1686
rect 1694 1683 1695 1687
rect 1699 1683 1700 1687
rect 1694 1682 1700 1683
rect 1475 1676 1674 1678
rect 1475 1675 1476 1676
rect 1470 1674 1476 1675
rect 154 1671 160 1672
rect 154 1667 155 1671
rect 159 1670 160 1671
rect 159 1668 731 1670
rect 159 1667 160 1668
rect 154 1666 160 1667
rect 134 1663 140 1664
rect 110 1661 116 1662
rect 110 1657 111 1661
rect 115 1657 116 1661
rect 134 1659 135 1663
rect 139 1659 140 1663
rect 134 1658 140 1659
rect 174 1663 180 1664
rect 174 1659 175 1663
rect 179 1659 180 1663
rect 174 1658 180 1659
rect 262 1663 268 1664
rect 262 1659 263 1663
rect 267 1659 268 1663
rect 262 1658 268 1659
rect 390 1663 396 1664
rect 390 1659 391 1663
rect 395 1659 396 1663
rect 390 1658 396 1659
rect 542 1663 548 1664
rect 542 1659 543 1663
rect 547 1659 548 1663
rect 542 1658 548 1659
rect 710 1663 716 1664
rect 710 1659 711 1663
rect 715 1659 716 1663
rect 710 1658 716 1659
rect 110 1656 116 1657
rect 729 1656 731 1668
rect 878 1663 884 1664
rect 878 1659 879 1663
rect 883 1659 884 1663
rect 878 1658 884 1659
rect 1038 1663 1044 1664
rect 1038 1659 1039 1663
rect 1043 1659 1044 1663
rect 1038 1658 1044 1659
rect 1182 1663 1188 1664
rect 1182 1659 1183 1663
rect 1187 1659 1188 1663
rect 1182 1658 1188 1659
rect 1318 1663 1324 1664
rect 1318 1659 1319 1663
rect 1323 1659 1324 1663
rect 1318 1658 1324 1659
rect 1438 1663 1444 1664
rect 1438 1659 1439 1663
rect 1443 1659 1444 1663
rect 1438 1658 1444 1659
rect 1558 1663 1564 1664
rect 1558 1659 1559 1663
rect 1563 1659 1564 1663
rect 1558 1658 1564 1659
rect 1654 1663 1660 1664
rect 1654 1659 1655 1663
rect 1659 1659 1660 1663
rect 1654 1658 1660 1659
rect 1694 1661 1700 1662
rect 1694 1657 1695 1661
rect 1699 1657 1700 1661
rect 1694 1656 1700 1657
rect 151 1655 157 1656
rect 151 1651 152 1655
rect 156 1654 157 1655
rect 191 1655 197 1656
rect 156 1652 186 1654
rect 156 1651 157 1652
rect 151 1650 157 1651
rect 134 1646 140 1647
rect 110 1644 116 1645
rect 110 1640 111 1644
rect 115 1640 116 1644
rect 134 1642 135 1646
rect 139 1642 140 1646
rect 134 1641 140 1642
rect 174 1646 180 1647
rect 174 1642 175 1646
rect 179 1642 180 1646
rect 174 1641 180 1642
rect 110 1639 116 1640
rect 151 1639 160 1640
rect 151 1635 152 1639
rect 159 1635 160 1639
rect 184 1638 186 1652
rect 191 1651 192 1655
rect 196 1654 197 1655
rect 279 1655 285 1656
rect 196 1652 238 1654
rect 196 1651 197 1652
rect 191 1650 197 1651
rect 191 1639 197 1640
rect 191 1638 192 1639
rect 184 1636 192 1638
rect 151 1634 160 1635
rect 191 1635 192 1636
rect 196 1635 197 1639
rect 236 1638 238 1652
rect 279 1651 280 1655
rect 284 1654 285 1655
rect 342 1655 348 1656
rect 342 1654 343 1655
rect 284 1652 343 1654
rect 284 1651 285 1652
rect 279 1650 285 1651
rect 342 1651 343 1652
rect 347 1651 348 1655
rect 342 1650 348 1651
rect 407 1655 413 1656
rect 407 1651 408 1655
rect 412 1654 413 1655
rect 559 1655 565 1656
rect 412 1652 486 1654
rect 412 1651 413 1652
rect 407 1650 413 1651
rect 262 1646 268 1647
rect 262 1642 263 1646
rect 267 1642 268 1646
rect 262 1641 268 1642
rect 390 1646 396 1647
rect 390 1642 391 1646
rect 395 1642 396 1646
rect 390 1641 396 1642
rect 279 1639 285 1640
rect 279 1638 280 1639
rect 236 1636 280 1638
rect 191 1634 197 1635
rect 279 1635 280 1636
rect 284 1635 285 1639
rect 279 1634 285 1635
rect 406 1639 413 1640
rect 406 1635 407 1639
rect 412 1635 413 1639
rect 484 1638 486 1652
rect 559 1651 560 1655
rect 564 1654 565 1655
rect 727 1655 733 1656
rect 564 1652 622 1654
rect 564 1651 565 1652
rect 559 1650 565 1651
rect 542 1646 548 1647
rect 542 1642 543 1646
rect 547 1642 548 1646
rect 542 1641 548 1642
rect 559 1639 565 1640
rect 559 1638 560 1639
rect 484 1636 560 1638
rect 406 1634 413 1635
rect 559 1635 560 1636
rect 564 1635 565 1639
rect 620 1638 622 1652
rect 727 1651 728 1655
rect 732 1651 733 1655
rect 727 1650 733 1651
rect 894 1655 901 1656
rect 894 1651 895 1655
rect 900 1651 901 1655
rect 1055 1655 1061 1656
rect 1055 1654 1056 1655
rect 894 1650 901 1651
rect 976 1652 1056 1654
rect 710 1646 716 1647
rect 710 1642 711 1646
rect 715 1642 716 1646
rect 710 1641 716 1642
rect 878 1646 884 1647
rect 878 1642 879 1646
rect 883 1642 884 1646
rect 878 1641 884 1642
rect 727 1639 733 1640
rect 727 1638 728 1639
rect 620 1636 728 1638
rect 559 1634 565 1635
rect 727 1635 728 1636
rect 732 1635 733 1639
rect 727 1634 733 1635
rect 895 1639 901 1640
rect 895 1635 896 1639
rect 900 1638 901 1639
rect 976 1638 978 1652
rect 1055 1651 1056 1652
rect 1060 1651 1061 1655
rect 1055 1650 1061 1651
rect 1198 1655 1205 1656
rect 1198 1651 1199 1655
rect 1204 1651 1205 1655
rect 1335 1655 1341 1656
rect 1335 1654 1336 1655
rect 1198 1650 1205 1651
rect 1272 1652 1336 1654
rect 1038 1646 1044 1647
rect 1038 1642 1039 1646
rect 1043 1642 1044 1646
rect 1038 1641 1044 1642
rect 1182 1646 1188 1647
rect 1182 1642 1183 1646
rect 1187 1642 1188 1646
rect 1182 1641 1188 1642
rect 900 1636 978 1638
rect 1018 1639 1024 1640
rect 900 1635 901 1636
rect 895 1634 901 1635
rect 1018 1635 1019 1639
rect 1023 1638 1024 1639
rect 1055 1639 1061 1640
rect 1055 1638 1056 1639
rect 1023 1636 1056 1638
rect 1023 1635 1024 1636
rect 1018 1634 1024 1635
rect 1055 1635 1056 1636
rect 1060 1635 1061 1639
rect 1055 1634 1061 1635
rect 1199 1639 1205 1640
rect 1199 1635 1200 1639
rect 1204 1638 1205 1639
rect 1272 1638 1274 1652
rect 1335 1651 1336 1652
rect 1340 1651 1341 1655
rect 1335 1650 1341 1651
rect 1455 1655 1461 1656
rect 1455 1651 1456 1655
rect 1460 1654 1461 1655
rect 1575 1655 1581 1656
rect 1460 1652 1518 1654
rect 1460 1651 1461 1652
rect 1455 1650 1461 1651
rect 1318 1646 1324 1647
rect 1318 1642 1319 1646
rect 1323 1642 1324 1646
rect 1318 1641 1324 1642
rect 1438 1646 1444 1647
rect 1438 1642 1439 1646
rect 1443 1642 1444 1646
rect 1438 1641 1444 1642
rect 1204 1636 1274 1638
rect 1335 1639 1341 1640
rect 1204 1635 1205 1636
rect 1199 1634 1205 1635
rect 1335 1635 1336 1639
rect 1340 1638 1341 1639
rect 1374 1639 1380 1640
rect 1374 1638 1375 1639
rect 1340 1636 1375 1638
rect 1340 1635 1341 1636
rect 1335 1634 1341 1635
rect 1374 1635 1375 1636
rect 1379 1635 1380 1639
rect 1374 1634 1380 1635
rect 1455 1639 1461 1640
rect 1455 1635 1456 1639
rect 1460 1638 1461 1639
rect 1470 1639 1476 1640
rect 1470 1638 1471 1639
rect 1460 1636 1471 1638
rect 1460 1635 1461 1636
rect 1455 1634 1461 1635
rect 1470 1635 1471 1636
rect 1475 1635 1476 1639
rect 1516 1638 1518 1652
rect 1575 1651 1576 1655
rect 1580 1654 1581 1655
rect 1670 1655 1677 1656
rect 1580 1652 1626 1654
rect 1580 1651 1581 1652
rect 1575 1650 1581 1651
rect 1558 1646 1564 1647
rect 1558 1642 1559 1646
rect 1563 1642 1564 1646
rect 1558 1641 1564 1642
rect 1575 1639 1581 1640
rect 1575 1638 1576 1639
rect 1516 1636 1576 1638
rect 1470 1634 1476 1635
rect 1575 1635 1576 1636
rect 1580 1635 1581 1639
rect 1624 1638 1626 1652
rect 1670 1651 1671 1655
rect 1676 1651 1677 1655
rect 1670 1650 1677 1651
rect 1654 1646 1660 1647
rect 1654 1642 1655 1646
rect 1659 1642 1660 1646
rect 1654 1641 1660 1642
rect 1694 1644 1700 1645
rect 1694 1640 1695 1644
rect 1699 1640 1700 1644
rect 1671 1639 1677 1640
rect 1694 1639 1700 1640
rect 1671 1638 1672 1639
rect 1624 1636 1672 1638
rect 1575 1634 1581 1635
rect 1671 1635 1672 1636
rect 1676 1635 1677 1639
rect 1671 1634 1677 1635
rect 79 1631 85 1632
rect 79 1627 80 1631
rect 84 1630 85 1631
rect 186 1631 192 1632
rect 186 1630 187 1631
rect 84 1628 187 1630
rect 84 1627 85 1628
rect 79 1626 85 1627
rect 186 1627 187 1628
rect 191 1627 192 1631
rect 186 1626 192 1627
rect 582 1623 588 1624
rect 582 1622 583 1623
rect 321 1620 583 1622
rect 153 1612 178 1614
rect 151 1611 157 1612
rect 110 1608 116 1609
rect 110 1604 111 1608
rect 115 1604 116 1608
rect 151 1607 152 1611
rect 156 1607 157 1611
rect 110 1603 116 1604
rect 134 1606 140 1607
rect 151 1606 157 1607
rect 166 1606 172 1607
rect 134 1602 135 1606
rect 139 1602 140 1606
rect 134 1601 140 1602
rect 166 1602 167 1606
rect 171 1602 172 1606
rect 166 1601 172 1602
rect 150 1595 157 1596
rect 110 1591 116 1592
rect 110 1587 111 1591
rect 115 1587 116 1591
rect 150 1591 151 1595
rect 156 1591 157 1595
rect 176 1594 178 1612
rect 183 1611 189 1612
rect 183 1607 184 1611
rect 188 1610 189 1611
rect 215 1611 221 1612
rect 188 1608 194 1610
rect 188 1607 189 1608
rect 183 1606 189 1607
rect 192 1598 194 1608
rect 215 1607 216 1611
rect 220 1610 221 1611
rect 263 1611 269 1612
rect 220 1608 242 1610
rect 220 1607 221 1608
rect 198 1606 204 1607
rect 215 1606 221 1607
rect 198 1602 199 1606
rect 203 1602 204 1606
rect 198 1601 204 1602
rect 240 1598 242 1608
rect 263 1607 264 1611
rect 268 1610 269 1611
rect 321 1610 323 1620
rect 582 1619 583 1620
rect 587 1619 588 1623
rect 582 1618 588 1619
rect 351 1615 357 1616
rect 268 1608 323 1610
rect 342 1611 349 1612
rect 268 1607 269 1608
rect 342 1607 343 1611
rect 348 1607 349 1611
rect 351 1611 352 1615
rect 356 1614 357 1615
rect 463 1615 469 1616
rect 356 1612 459 1614
rect 356 1611 357 1612
rect 351 1610 357 1611
rect 455 1611 461 1612
rect 455 1607 456 1611
rect 460 1607 461 1611
rect 463 1611 464 1615
rect 468 1614 469 1615
rect 1210 1615 1216 1616
rect 468 1612 578 1614
rect 729 1612 866 1614
rect 468 1611 469 1612
rect 463 1610 469 1611
rect 576 1610 578 1612
rect 583 1611 589 1612
rect 583 1610 584 1611
rect 576 1608 584 1610
rect 583 1607 584 1608
rect 588 1607 589 1611
rect 727 1611 733 1612
rect 727 1607 728 1611
rect 732 1607 733 1611
rect 246 1606 252 1607
rect 263 1606 269 1607
rect 326 1606 332 1607
rect 342 1606 349 1607
rect 438 1606 444 1607
rect 455 1606 461 1607
rect 566 1606 572 1607
rect 583 1606 589 1607
rect 710 1606 716 1607
rect 727 1606 733 1607
rect 854 1606 860 1607
rect 246 1602 247 1606
rect 251 1602 252 1606
rect 246 1601 252 1602
rect 326 1602 327 1606
rect 331 1602 332 1606
rect 326 1601 332 1602
rect 438 1602 439 1606
rect 443 1602 444 1606
rect 438 1601 444 1602
rect 566 1602 567 1606
rect 571 1602 572 1606
rect 566 1601 572 1602
rect 710 1602 711 1606
rect 715 1602 716 1606
rect 710 1601 716 1602
rect 854 1602 855 1606
rect 859 1602 860 1606
rect 854 1601 860 1602
rect 192 1596 198 1598
rect 240 1596 246 1598
rect 183 1595 189 1596
rect 183 1594 184 1595
rect 176 1592 184 1594
rect 150 1590 157 1591
rect 183 1591 184 1592
rect 188 1591 189 1595
rect 196 1594 210 1596
rect 215 1595 221 1596
rect 215 1594 216 1595
rect 208 1592 216 1594
rect 183 1590 189 1591
rect 215 1591 216 1592
rect 220 1591 221 1595
rect 244 1594 258 1596
rect 263 1595 269 1596
rect 263 1594 264 1595
rect 256 1592 264 1594
rect 215 1590 221 1591
rect 263 1591 264 1592
rect 268 1591 269 1595
rect 263 1590 269 1591
rect 343 1595 349 1596
rect 343 1591 344 1595
rect 348 1594 349 1595
rect 351 1595 357 1596
rect 351 1594 352 1595
rect 348 1592 352 1594
rect 348 1591 349 1592
rect 343 1590 349 1591
rect 351 1591 352 1592
rect 356 1591 357 1595
rect 351 1590 357 1591
rect 455 1595 461 1596
rect 455 1591 456 1595
rect 460 1594 461 1595
rect 463 1595 469 1596
rect 463 1594 464 1595
rect 460 1592 464 1594
rect 460 1591 461 1592
rect 455 1590 461 1591
rect 463 1591 464 1592
rect 468 1591 469 1595
rect 463 1590 469 1591
rect 582 1595 589 1596
rect 582 1591 583 1595
rect 588 1591 589 1595
rect 582 1590 589 1591
rect 722 1595 733 1596
rect 722 1591 723 1595
rect 727 1591 728 1595
rect 732 1591 733 1595
rect 864 1594 866 1612
rect 871 1611 877 1612
rect 871 1607 872 1611
rect 876 1610 877 1611
rect 974 1611 980 1612
rect 974 1610 975 1611
rect 876 1608 975 1610
rect 876 1607 877 1608
rect 871 1606 877 1607
rect 974 1607 975 1608
rect 979 1607 980 1611
rect 1015 1611 1021 1612
rect 1015 1607 1016 1611
rect 1020 1610 1021 1611
rect 1078 1611 1084 1612
rect 1078 1610 1079 1611
rect 1020 1608 1079 1610
rect 1020 1607 1021 1608
rect 974 1606 980 1607
rect 998 1606 1004 1607
rect 1015 1606 1021 1607
rect 1078 1607 1079 1608
rect 1083 1607 1084 1611
rect 1143 1611 1149 1612
rect 1143 1607 1144 1611
rect 1148 1610 1149 1611
rect 1174 1611 1180 1612
rect 1174 1610 1175 1611
rect 1148 1608 1175 1610
rect 1148 1607 1149 1608
rect 1078 1606 1084 1607
rect 1126 1606 1132 1607
rect 1143 1606 1149 1607
rect 1174 1607 1175 1608
rect 1179 1607 1180 1611
rect 1210 1611 1211 1615
rect 1215 1614 1216 1615
rect 1215 1612 1258 1614
rect 1456 1612 1474 1614
rect 1585 1612 1666 1614
rect 1215 1611 1216 1612
rect 1210 1610 1216 1611
rect 1256 1610 1258 1612
rect 1263 1611 1269 1612
rect 1263 1610 1264 1611
rect 1256 1608 1264 1610
rect 1263 1607 1264 1608
rect 1268 1607 1269 1611
rect 1375 1611 1381 1612
rect 1375 1607 1376 1611
rect 1380 1610 1381 1611
rect 1456 1610 1458 1612
rect 1380 1608 1458 1610
rect 1380 1607 1381 1608
rect 1174 1606 1180 1607
rect 1246 1606 1252 1607
rect 1263 1606 1269 1607
rect 1358 1606 1364 1607
rect 1375 1606 1381 1607
rect 1462 1606 1468 1607
rect 998 1602 999 1606
rect 1003 1602 1004 1606
rect 998 1601 1004 1602
rect 1126 1602 1127 1606
rect 1131 1602 1132 1606
rect 1126 1601 1132 1602
rect 1246 1602 1247 1606
rect 1251 1602 1252 1606
rect 1246 1601 1252 1602
rect 1358 1602 1359 1606
rect 1363 1602 1364 1606
rect 1358 1601 1364 1602
rect 1462 1602 1463 1606
rect 1467 1602 1468 1606
rect 1462 1601 1468 1602
rect 871 1595 877 1596
rect 871 1594 872 1595
rect 864 1592 872 1594
rect 722 1590 733 1591
rect 871 1591 872 1592
rect 876 1591 877 1595
rect 871 1590 877 1591
rect 1015 1595 1024 1596
rect 1015 1591 1016 1595
rect 1023 1591 1024 1595
rect 1015 1590 1024 1591
rect 1143 1595 1149 1596
rect 1143 1591 1144 1595
rect 1148 1594 1149 1595
rect 1210 1595 1216 1596
rect 1210 1594 1211 1595
rect 1148 1592 1211 1594
rect 1148 1591 1149 1592
rect 1143 1590 1149 1591
rect 1210 1591 1211 1592
rect 1215 1591 1216 1595
rect 1210 1590 1216 1591
rect 1263 1595 1269 1596
rect 1263 1591 1264 1595
rect 1268 1594 1269 1595
rect 1342 1595 1348 1596
rect 1342 1594 1343 1595
rect 1268 1592 1343 1594
rect 1268 1591 1269 1592
rect 1263 1590 1269 1591
rect 1342 1591 1343 1592
rect 1347 1591 1348 1595
rect 1342 1590 1348 1591
rect 1374 1595 1381 1596
rect 1374 1591 1375 1595
rect 1380 1591 1381 1595
rect 1472 1594 1474 1612
rect 1478 1611 1485 1612
rect 1478 1607 1479 1611
rect 1484 1607 1485 1611
rect 1583 1611 1589 1612
rect 1583 1607 1584 1611
rect 1588 1607 1589 1611
rect 1478 1606 1485 1607
rect 1566 1606 1572 1607
rect 1583 1606 1589 1607
rect 1654 1606 1660 1607
rect 1566 1602 1567 1606
rect 1571 1602 1572 1606
rect 1566 1601 1572 1602
rect 1654 1602 1655 1606
rect 1659 1602 1660 1606
rect 1654 1601 1660 1602
rect 1479 1595 1485 1596
rect 1479 1594 1480 1595
rect 1472 1592 1480 1594
rect 1374 1590 1381 1591
rect 1479 1591 1480 1592
rect 1484 1591 1485 1595
rect 1479 1590 1485 1591
rect 1583 1595 1589 1596
rect 1583 1591 1584 1595
rect 1588 1594 1589 1595
rect 1622 1595 1628 1596
rect 1622 1594 1623 1595
rect 1588 1592 1623 1594
rect 1588 1591 1589 1592
rect 1583 1590 1589 1591
rect 1622 1591 1623 1592
rect 1627 1591 1628 1595
rect 1664 1594 1666 1612
rect 1670 1611 1677 1612
rect 1670 1607 1671 1611
rect 1676 1607 1677 1611
rect 1670 1606 1677 1607
rect 1694 1608 1700 1609
rect 1694 1604 1695 1608
rect 1699 1604 1700 1608
rect 1694 1603 1700 1604
rect 1671 1595 1677 1596
rect 1671 1594 1672 1595
rect 1664 1592 1672 1594
rect 1622 1590 1628 1591
rect 1671 1591 1672 1592
rect 1676 1591 1677 1595
rect 1671 1590 1677 1591
rect 1694 1591 1700 1592
rect 110 1586 116 1587
rect 134 1589 140 1590
rect 134 1585 135 1589
rect 139 1585 140 1589
rect 134 1584 140 1585
rect 166 1589 172 1590
rect 166 1585 167 1589
rect 171 1585 172 1589
rect 166 1584 172 1585
rect 198 1589 204 1590
rect 198 1585 199 1589
rect 203 1585 204 1589
rect 198 1584 204 1585
rect 246 1589 252 1590
rect 246 1585 247 1589
rect 251 1585 252 1589
rect 246 1584 252 1585
rect 326 1589 332 1590
rect 326 1585 327 1589
rect 331 1585 332 1589
rect 326 1584 332 1585
rect 438 1589 444 1590
rect 438 1585 439 1589
rect 443 1585 444 1589
rect 438 1584 444 1585
rect 566 1589 572 1590
rect 566 1585 567 1589
rect 571 1585 572 1589
rect 566 1584 572 1585
rect 710 1589 716 1590
rect 710 1585 711 1589
rect 715 1585 716 1589
rect 710 1584 716 1585
rect 854 1589 860 1590
rect 854 1585 855 1589
rect 859 1585 860 1589
rect 854 1584 860 1585
rect 998 1589 1004 1590
rect 998 1585 999 1589
rect 1003 1585 1004 1589
rect 998 1584 1004 1585
rect 1126 1589 1132 1590
rect 1126 1585 1127 1589
rect 1131 1585 1132 1589
rect 1126 1584 1132 1585
rect 1246 1589 1252 1590
rect 1246 1585 1247 1589
rect 1251 1585 1252 1589
rect 1246 1584 1252 1585
rect 1358 1589 1364 1590
rect 1358 1585 1359 1589
rect 1363 1585 1364 1589
rect 1358 1584 1364 1585
rect 1462 1589 1468 1590
rect 1462 1585 1463 1589
rect 1467 1585 1468 1589
rect 1462 1584 1468 1585
rect 1566 1589 1572 1590
rect 1566 1585 1567 1589
rect 1571 1585 1572 1589
rect 1566 1584 1572 1585
rect 1654 1589 1660 1590
rect 1654 1585 1655 1589
rect 1659 1585 1660 1589
rect 1694 1587 1695 1591
rect 1699 1587 1700 1591
rect 1694 1586 1700 1587
rect 1654 1584 1660 1585
rect 134 1575 140 1576
rect 110 1573 116 1574
rect 110 1569 111 1573
rect 115 1569 116 1573
rect 134 1571 135 1575
rect 139 1571 140 1575
rect 134 1570 140 1571
rect 166 1575 172 1576
rect 166 1571 167 1575
rect 171 1571 172 1575
rect 166 1570 172 1571
rect 230 1575 236 1576
rect 230 1571 231 1575
rect 235 1571 236 1575
rect 230 1570 236 1571
rect 286 1575 292 1576
rect 286 1571 287 1575
rect 291 1571 292 1575
rect 286 1570 292 1571
rect 342 1575 348 1576
rect 342 1571 343 1575
rect 347 1571 348 1575
rect 342 1570 348 1571
rect 398 1575 404 1576
rect 398 1571 399 1575
rect 403 1571 404 1575
rect 398 1570 404 1571
rect 454 1575 460 1576
rect 454 1571 455 1575
rect 459 1571 460 1575
rect 454 1570 460 1571
rect 510 1575 516 1576
rect 510 1571 511 1575
rect 515 1571 516 1575
rect 510 1570 516 1571
rect 574 1575 580 1576
rect 574 1571 575 1575
rect 579 1571 580 1575
rect 574 1570 580 1571
rect 654 1575 660 1576
rect 654 1571 655 1575
rect 659 1571 660 1575
rect 654 1570 660 1571
rect 750 1575 756 1576
rect 750 1571 751 1575
rect 755 1571 756 1575
rect 750 1570 756 1571
rect 854 1575 860 1576
rect 854 1571 855 1575
rect 859 1571 860 1575
rect 854 1570 860 1571
rect 958 1575 964 1576
rect 958 1571 959 1575
rect 963 1571 964 1575
rect 958 1570 964 1571
rect 1062 1575 1068 1576
rect 1062 1571 1063 1575
rect 1067 1571 1068 1575
rect 1062 1570 1068 1571
rect 1158 1575 1164 1576
rect 1158 1571 1159 1575
rect 1163 1571 1164 1575
rect 1158 1570 1164 1571
rect 1246 1575 1252 1576
rect 1246 1571 1247 1575
rect 1251 1571 1252 1575
rect 1246 1570 1252 1571
rect 1326 1575 1332 1576
rect 1326 1571 1327 1575
rect 1331 1571 1332 1575
rect 1326 1570 1332 1571
rect 1398 1575 1404 1576
rect 1398 1571 1399 1575
rect 1403 1571 1404 1575
rect 1398 1570 1404 1571
rect 1470 1575 1476 1576
rect 1470 1571 1471 1575
rect 1475 1571 1476 1575
rect 1470 1570 1476 1571
rect 1534 1575 1540 1576
rect 1534 1571 1535 1575
rect 1539 1571 1540 1575
rect 1534 1570 1540 1571
rect 1606 1575 1612 1576
rect 1606 1571 1607 1575
rect 1611 1571 1612 1575
rect 1606 1570 1612 1571
rect 1654 1575 1660 1576
rect 1654 1571 1655 1575
rect 1659 1571 1660 1575
rect 1702 1575 1708 1576
rect 1654 1570 1660 1571
rect 1694 1573 1700 1574
rect 110 1568 116 1569
rect 1694 1569 1695 1573
rect 1699 1569 1700 1573
rect 1702 1571 1703 1575
rect 1707 1574 1708 1575
rect 1747 1575 1753 1576
rect 1747 1574 1748 1575
rect 1707 1572 1748 1574
rect 1707 1571 1708 1572
rect 1702 1570 1708 1571
rect 1747 1571 1748 1572
rect 1752 1571 1753 1575
rect 1747 1570 1753 1571
rect 1694 1568 1700 1569
rect 151 1567 157 1568
rect 151 1563 152 1567
rect 156 1566 157 1567
rect 183 1567 189 1568
rect 156 1564 178 1566
rect 156 1563 157 1564
rect 151 1562 157 1563
rect 134 1558 140 1559
rect 110 1556 116 1557
rect 110 1552 111 1556
rect 115 1552 116 1556
rect 134 1554 135 1558
rect 139 1554 140 1558
rect 134 1553 140 1554
rect 166 1558 172 1559
rect 166 1554 167 1558
rect 171 1554 172 1558
rect 166 1553 172 1554
rect 110 1551 116 1552
rect 150 1551 157 1552
rect 150 1547 151 1551
rect 156 1547 157 1551
rect 176 1550 178 1564
rect 183 1563 184 1567
rect 188 1566 189 1567
rect 247 1567 253 1568
rect 188 1564 218 1566
rect 188 1563 189 1564
rect 183 1562 189 1563
rect 183 1551 189 1552
rect 183 1550 184 1551
rect 176 1548 184 1550
rect 150 1546 157 1547
rect 183 1547 184 1548
rect 188 1547 189 1551
rect 216 1550 218 1564
rect 247 1563 248 1567
rect 252 1566 253 1567
rect 298 1567 309 1568
rect 252 1564 278 1566
rect 252 1563 253 1564
rect 247 1562 253 1563
rect 230 1558 236 1559
rect 230 1554 231 1558
rect 235 1554 236 1558
rect 230 1553 236 1554
rect 247 1551 253 1552
rect 247 1550 248 1551
rect 216 1548 248 1550
rect 183 1546 189 1547
rect 247 1547 248 1548
rect 252 1547 253 1551
rect 276 1550 278 1564
rect 298 1563 299 1567
rect 303 1563 304 1567
rect 308 1563 309 1567
rect 298 1562 309 1563
rect 359 1567 365 1568
rect 359 1563 360 1567
rect 364 1566 365 1567
rect 378 1567 384 1568
rect 378 1566 379 1567
rect 364 1564 379 1566
rect 364 1563 365 1564
rect 359 1562 365 1563
rect 378 1563 379 1564
rect 383 1563 384 1567
rect 415 1567 421 1568
rect 415 1566 416 1567
rect 378 1562 384 1563
rect 388 1564 416 1566
rect 286 1558 292 1559
rect 286 1554 287 1558
rect 291 1554 292 1558
rect 286 1553 292 1554
rect 342 1558 348 1559
rect 342 1554 343 1558
rect 347 1554 348 1558
rect 342 1553 348 1554
rect 303 1551 309 1552
rect 303 1550 304 1551
rect 276 1548 304 1550
rect 247 1546 253 1547
rect 303 1547 304 1548
rect 308 1547 309 1551
rect 303 1546 309 1547
rect 359 1551 365 1552
rect 359 1547 360 1551
rect 364 1550 365 1551
rect 388 1550 390 1564
rect 415 1563 416 1564
rect 420 1563 421 1567
rect 471 1567 477 1568
rect 471 1566 472 1567
rect 415 1562 421 1563
rect 448 1564 472 1566
rect 398 1558 404 1559
rect 398 1554 399 1558
rect 403 1554 404 1558
rect 398 1553 404 1554
rect 364 1548 390 1550
rect 415 1551 421 1552
rect 364 1547 365 1548
rect 359 1546 365 1547
rect 415 1547 416 1551
rect 420 1550 421 1551
rect 448 1550 450 1564
rect 471 1563 472 1564
rect 476 1563 477 1567
rect 527 1567 533 1568
rect 527 1566 528 1567
rect 471 1562 477 1563
rect 500 1564 528 1566
rect 454 1558 460 1559
rect 454 1554 455 1558
rect 459 1554 460 1558
rect 454 1553 460 1554
rect 420 1548 450 1550
rect 471 1551 477 1552
rect 420 1547 421 1548
rect 415 1546 421 1547
rect 471 1547 472 1551
rect 476 1550 477 1551
rect 500 1550 502 1564
rect 527 1563 528 1564
rect 532 1563 533 1567
rect 591 1567 597 1568
rect 591 1566 592 1567
rect 527 1562 533 1563
rect 564 1564 592 1566
rect 510 1558 516 1559
rect 510 1554 511 1558
rect 515 1554 516 1558
rect 510 1553 516 1554
rect 476 1548 502 1550
rect 527 1551 533 1552
rect 476 1547 477 1548
rect 471 1546 477 1547
rect 527 1547 528 1551
rect 532 1550 533 1551
rect 564 1550 566 1564
rect 591 1563 592 1564
rect 596 1563 597 1567
rect 591 1562 597 1563
rect 671 1567 677 1568
rect 671 1563 672 1567
rect 676 1566 677 1567
rect 730 1567 736 1568
rect 730 1566 731 1567
rect 676 1564 731 1566
rect 676 1563 677 1564
rect 671 1562 677 1563
rect 730 1563 731 1564
rect 735 1563 736 1567
rect 730 1562 736 1563
rect 767 1567 773 1568
rect 767 1563 768 1567
rect 772 1566 773 1567
rect 871 1567 877 1568
rect 772 1564 866 1566
rect 772 1563 773 1564
rect 767 1562 773 1563
rect 722 1559 728 1560
rect 574 1558 580 1559
rect 574 1554 575 1558
rect 579 1554 580 1558
rect 574 1553 580 1554
rect 654 1558 660 1559
rect 722 1558 723 1559
rect 654 1554 655 1558
rect 659 1554 660 1558
rect 654 1553 660 1554
rect 664 1556 723 1558
rect 532 1548 566 1550
rect 591 1551 597 1552
rect 532 1547 533 1548
rect 527 1546 533 1547
rect 591 1547 592 1551
rect 596 1550 597 1551
rect 664 1550 666 1556
rect 722 1555 723 1556
rect 727 1555 728 1559
rect 722 1554 728 1555
rect 750 1558 756 1559
rect 750 1554 751 1558
rect 755 1554 756 1558
rect 750 1553 756 1554
rect 854 1558 860 1559
rect 854 1554 855 1558
rect 859 1554 860 1558
rect 854 1553 860 1554
rect 596 1548 666 1550
rect 671 1551 677 1552
rect 596 1547 597 1548
rect 591 1546 597 1547
rect 671 1547 672 1551
rect 676 1547 677 1551
rect 671 1546 677 1547
rect 758 1551 764 1552
rect 758 1547 759 1551
rect 763 1550 764 1551
rect 767 1551 773 1552
rect 767 1550 768 1551
rect 763 1548 768 1550
rect 763 1547 764 1548
rect 758 1546 764 1547
rect 767 1547 768 1548
rect 772 1547 773 1551
rect 864 1550 866 1564
rect 871 1563 872 1567
rect 876 1566 877 1567
rect 974 1567 981 1568
rect 876 1564 926 1566
rect 876 1563 877 1564
rect 871 1562 877 1563
rect 871 1551 877 1552
rect 871 1550 872 1551
rect 864 1548 872 1550
rect 767 1546 773 1547
rect 871 1547 872 1548
rect 876 1547 877 1551
rect 924 1550 926 1564
rect 974 1563 975 1567
rect 980 1563 981 1567
rect 974 1562 981 1563
rect 1078 1567 1085 1568
rect 1078 1563 1079 1567
rect 1084 1563 1085 1567
rect 1078 1562 1085 1563
rect 1174 1567 1181 1568
rect 1174 1563 1175 1567
rect 1180 1563 1181 1567
rect 1174 1562 1181 1563
rect 1263 1567 1269 1568
rect 1263 1563 1264 1567
rect 1268 1566 1269 1567
rect 1343 1567 1349 1568
rect 1268 1564 1338 1566
rect 1268 1563 1269 1564
rect 1263 1562 1269 1563
rect 958 1558 964 1559
rect 958 1554 959 1558
rect 963 1554 964 1558
rect 958 1553 964 1554
rect 1062 1558 1068 1559
rect 1062 1554 1063 1558
rect 1067 1554 1068 1558
rect 1062 1553 1068 1554
rect 1158 1558 1164 1559
rect 1158 1554 1159 1558
rect 1163 1554 1164 1558
rect 1158 1553 1164 1554
rect 1246 1558 1252 1559
rect 1246 1554 1247 1558
rect 1251 1554 1252 1558
rect 1246 1553 1252 1554
rect 1326 1558 1332 1559
rect 1326 1554 1327 1558
rect 1331 1554 1332 1558
rect 1336 1558 1338 1564
rect 1343 1563 1344 1567
rect 1348 1566 1349 1567
rect 1374 1567 1380 1568
rect 1374 1566 1375 1567
rect 1348 1564 1375 1566
rect 1348 1563 1349 1564
rect 1343 1562 1349 1563
rect 1374 1563 1375 1564
rect 1379 1563 1380 1567
rect 1374 1562 1380 1563
rect 1415 1567 1421 1568
rect 1415 1563 1416 1567
rect 1420 1566 1421 1567
rect 1487 1567 1493 1568
rect 1420 1564 1454 1566
rect 1420 1563 1421 1564
rect 1415 1562 1421 1563
rect 1398 1558 1404 1559
rect 1336 1556 1354 1558
rect 1326 1553 1332 1554
rect 975 1551 981 1552
rect 975 1550 976 1551
rect 924 1548 976 1550
rect 871 1546 877 1547
rect 975 1547 976 1548
rect 980 1547 981 1551
rect 975 1546 981 1547
rect 1079 1551 1085 1552
rect 1079 1547 1080 1551
rect 1084 1550 1085 1551
rect 1102 1551 1108 1552
rect 1102 1550 1103 1551
rect 1084 1548 1103 1550
rect 1084 1547 1085 1548
rect 1079 1546 1085 1547
rect 1102 1547 1103 1548
rect 1107 1547 1108 1551
rect 1102 1546 1108 1547
rect 1175 1551 1181 1552
rect 1175 1547 1176 1551
rect 1180 1550 1181 1551
rect 1194 1551 1200 1552
rect 1180 1548 1190 1550
rect 1180 1547 1181 1548
rect 1175 1546 1181 1547
rect 298 1543 304 1544
rect 298 1542 299 1543
rect 153 1540 299 1542
rect 153 1532 155 1540
rect 298 1539 299 1540
rect 303 1539 304 1543
rect 298 1538 304 1539
rect 378 1543 384 1544
rect 378 1539 379 1543
rect 383 1542 384 1543
rect 554 1543 560 1544
rect 383 1540 419 1542
rect 383 1539 384 1540
rect 378 1538 384 1539
rect 159 1535 165 1536
rect 151 1531 157 1532
rect 110 1528 116 1529
rect 110 1524 111 1528
rect 115 1524 116 1528
rect 151 1527 152 1531
rect 156 1527 157 1531
rect 159 1531 160 1535
rect 164 1534 165 1535
rect 210 1535 216 1536
rect 164 1532 186 1534
rect 164 1531 165 1532
rect 159 1530 165 1531
rect 184 1530 186 1532
rect 191 1531 197 1532
rect 191 1530 192 1531
rect 184 1528 192 1530
rect 191 1527 192 1528
rect 196 1527 197 1531
rect 210 1531 211 1535
rect 215 1534 216 1535
rect 247 1535 253 1536
rect 215 1532 234 1534
rect 215 1531 216 1532
rect 210 1530 216 1531
rect 232 1530 234 1532
rect 239 1531 245 1532
rect 239 1530 240 1531
rect 232 1528 240 1530
rect 239 1527 240 1528
rect 244 1527 245 1531
rect 247 1531 248 1535
rect 252 1534 253 1535
rect 252 1532 290 1534
rect 353 1532 410 1534
rect 417 1532 419 1540
rect 554 1539 555 1543
rect 559 1542 560 1543
rect 673 1542 675 1546
rect 559 1540 675 1542
rect 1030 1543 1036 1544
rect 559 1539 560 1540
rect 554 1538 560 1539
rect 1030 1539 1031 1543
rect 1035 1542 1036 1543
rect 1188 1542 1190 1548
rect 1194 1547 1195 1551
rect 1199 1550 1200 1551
rect 1263 1551 1269 1552
rect 1263 1550 1264 1551
rect 1199 1548 1264 1550
rect 1199 1547 1200 1548
rect 1194 1546 1200 1547
rect 1263 1547 1264 1548
rect 1268 1547 1269 1551
rect 1263 1546 1269 1547
rect 1342 1551 1349 1552
rect 1342 1547 1343 1551
rect 1348 1547 1349 1551
rect 1352 1550 1354 1556
rect 1398 1554 1399 1558
rect 1403 1554 1404 1558
rect 1398 1553 1404 1554
rect 1415 1551 1421 1552
rect 1415 1550 1416 1551
rect 1352 1548 1416 1550
rect 1342 1546 1349 1547
rect 1415 1547 1416 1548
rect 1420 1547 1421 1551
rect 1452 1550 1454 1564
rect 1487 1563 1488 1567
rect 1492 1566 1493 1567
rect 1546 1567 1557 1568
rect 1492 1564 1522 1566
rect 1492 1563 1493 1564
rect 1487 1562 1493 1563
rect 1470 1558 1476 1559
rect 1470 1554 1471 1558
rect 1475 1554 1476 1558
rect 1470 1553 1476 1554
rect 1487 1551 1493 1552
rect 1487 1550 1488 1551
rect 1452 1548 1488 1550
rect 1415 1546 1421 1547
rect 1487 1547 1488 1548
rect 1492 1547 1493 1551
rect 1520 1550 1522 1564
rect 1546 1563 1547 1567
rect 1551 1563 1552 1567
rect 1556 1563 1557 1567
rect 1546 1562 1557 1563
rect 1623 1567 1629 1568
rect 1623 1563 1624 1567
rect 1628 1566 1629 1567
rect 1670 1567 1677 1568
rect 1628 1564 1650 1566
rect 1628 1563 1629 1564
rect 1623 1562 1629 1563
rect 1534 1558 1540 1559
rect 1534 1554 1535 1558
rect 1539 1554 1540 1558
rect 1534 1553 1540 1554
rect 1606 1558 1612 1559
rect 1606 1554 1607 1558
rect 1611 1554 1612 1558
rect 1606 1553 1612 1554
rect 1551 1551 1557 1552
rect 1551 1550 1552 1551
rect 1520 1548 1552 1550
rect 1487 1546 1493 1547
rect 1551 1547 1552 1548
rect 1556 1547 1557 1551
rect 1551 1546 1557 1547
rect 1622 1551 1629 1552
rect 1622 1547 1623 1551
rect 1628 1547 1629 1551
rect 1648 1550 1650 1564
rect 1670 1563 1671 1567
rect 1676 1563 1677 1567
rect 1670 1562 1677 1563
rect 1654 1558 1660 1559
rect 1654 1554 1655 1558
rect 1659 1554 1660 1558
rect 1654 1553 1660 1554
rect 1694 1556 1700 1557
rect 1694 1552 1695 1556
rect 1699 1552 1700 1556
rect 1671 1551 1677 1552
rect 1694 1551 1700 1552
rect 1671 1550 1672 1551
rect 1648 1548 1672 1550
rect 1622 1546 1629 1547
rect 1671 1547 1672 1548
rect 1676 1547 1677 1551
rect 1671 1546 1677 1547
rect 1263 1543 1269 1544
rect 1263 1542 1264 1543
rect 1035 1540 1264 1542
rect 1035 1539 1036 1540
rect 1030 1538 1036 1539
rect 1263 1539 1264 1540
rect 1268 1539 1269 1543
rect 1263 1538 1269 1539
rect 487 1535 493 1536
rect 252 1531 253 1532
rect 247 1530 253 1531
rect 288 1530 290 1532
rect 295 1531 301 1532
rect 295 1530 296 1531
rect 288 1528 296 1530
rect 295 1527 296 1528
rect 300 1527 301 1531
rect 351 1531 357 1532
rect 351 1527 352 1531
rect 356 1527 357 1531
rect 110 1523 116 1524
rect 134 1526 140 1527
rect 151 1526 157 1527
rect 174 1526 180 1527
rect 191 1526 197 1527
rect 222 1526 228 1527
rect 239 1526 245 1527
rect 278 1526 284 1527
rect 295 1526 301 1527
rect 334 1526 340 1527
rect 351 1526 357 1527
rect 398 1526 404 1527
rect 134 1522 135 1526
rect 139 1522 140 1526
rect 134 1521 140 1522
rect 174 1522 175 1526
rect 179 1522 180 1526
rect 174 1521 180 1522
rect 222 1522 223 1526
rect 227 1522 228 1526
rect 222 1521 228 1522
rect 278 1522 279 1526
rect 283 1522 284 1526
rect 278 1521 284 1522
rect 334 1522 335 1526
rect 339 1522 340 1526
rect 334 1521 340 1522
rect 398 1522 399 1526
rect 403 1522 404 1526
rect 398 1521 404 1522
rect 151 1515 157 1516
rect 110 1511 116 1512
rect 79 1507 85 1508
rect 79 1503 80 1507
rect 84 1506 85 1507
rect 102 1507 108 1508
rect 102 1506 103 1507
rect 84 1504 103 1506
rect 84 1503 85 1504
rect 79 1502 85 1503
rect 102 1503 103 1504
rect 107 1503 108 1507
rect 110 1507 111 1511
rect 115 1507 116 1511
rect 151 1511 152 1515
rect 156 1514 157 1515
rect 159 1515 165 1516
rect 159 1514 160 1515
rect 156 1512 160 1514
rect 156 1511 157 1512
rect 151 1510 157 1511
rect 159 1511 160 1512
rect 164 1511 165 1515
rect 159 1510 165 1511
rect 191 1515 197 1516
rect 191 1511 192 1515
rect 196 1514 197 1515
rect 210 1515 216 1516
rect 210 1514 211 1515
rect 196 1512 211 1514
rect 196 1511 197 1512
rect 191 1510 197 1511
rect 210 1511 211 1512
rect 215 1511 216 1515
rect 210 1510 216 1511
rect 239 1515 245 1516
rect 239 1511 240 1515
rect 244 1514 245 1515
rect 247 1515 253 1516
rect 247 1514 248 1515
rect 244 1512 248 1514
rect 244 1511 245 1512
rect 239 1510 245 1511
rect 247 1511 248 1512
rect 252 1511 253 1515
rect 247 1510 253 1511
rect 295 1515 301 1516
rect 295 1511 296 1515
rect 300 1514 301 1515
rect 318 1515 324 1516
rect 318 1514 319 1515
rect 300 1512 319 1514
rect 300 1511 301 1512
rect 295 1510 301 1511
rect 318 1511 319 1512
rect 323 1511 324 1515
rect 318 1510 324 1511
rect 350 1515 357 1516
rect 350 1511 351 1515
rect 356 1511 357 1515
rect 408 1514 410 1532
rect 415 1531 421 1532
rect 415 1527 416 1531
rect 420 1527 421 1531
rect 470 1531 476 1532
rect 470 1527 471 1531
rect 475 1530 476 1531
rect 479 1531 485 1532
rect 479 1530 480 1531
rect 475 1528 480 1530
rect 475 1527 476 1528
rect 415 1526 421 1527
rect 462 1526 468 1527
rect 470 1526 476 1527
rect 479 1527 480 1528
rect 484 1527 485 1531
rect 487 1531 488 1535
rect 492 1534 493 1535
rect 646 1535 652 1536
rect 492 1532 546 1534
rect 492 1531 493 1532
rect 487 1530 493 1531
rect 544 1530 546 1532
rect 551 1531 557 1532
rect 551 1530 552 1531
rect 544 1528 552 1530
rect 551 1527 552 1528
rect 556 1527 557 1531
rect 623 1531 629 1532
rect 623 1527 624 1531
rect 628 1530 629 1531
rect 638 1531 644 1532
rect 638 1530 639 1531
rect 628 1528 639 1530
rect 628 1527 629 1528
rect 479 1526 485 1527
rect 534 1526 540 1527
rect 551 1526 557 1527
rect 606 1526 612 1527
rect 623 1526 629 1527
rect 638 1527 639 1528
rect 643 1527 644 1531
rect 646 1531 647 1535
rect 651 1534 652 1535
rect 730 1535 736 1536
rect 651 1532 707 1534
rect 651 1531 652 1532
rect 646 1530 652 1531
rect 703 1531 709 1532
rect 703 1527 704 1531
rect 708 1527 709 1531
rect 730 1531 731 1535
rect 735 1534 736 1535
rect 799 1535 805 1536
rect 735 1532 795 1534
rect 735 1531 736 1532
rect 730 1530 736 1531
rect 791 1531 797 1532
rect 791 1527 792 1531
rect 796 1527 797 1531
rect 799 1531 800 1535
rect 804 1534 805 1535
rect 895 1535 901 1536
rect 804 1532 882 1534
rect 804 1531 805 1532
rect 799 1530 805 1531
rect 880 1530 882 1532
rect 887 1531 893 1532
rect 887 1530 888 1531
rect 880 1528 888 1530
rect 887 1527 888 1528
rect 892 1527 893 1531
rect 895 1531 896 1535
rect 900 1534 901 1535
rect 1254 1535 1260 1536
rect 900 1532 986 1534
rect 900 1531 901 1532
rect 895 1530 901 1531
rect 984 1530 986 1532
rect 991 1531 997 1532
rect 991 1530 992 1531
rect 984 1528 992 1530
rect 991 1527 992 1528
rect 996 1527 997 1531
rect 1094 1531 1101 1532
rect 1094 1527 1095 1531
rect 1100 1527 1101 1531
rect 1186 1531 1197 1532
rect 1186 1527 1187 1531
rect 1191 1527 1192 1531
rect 1196 1530 1197 1531
rect 1214 1531 1220 1532
rect 1214 1530 1215 1531
rect 1196 1528 1215 1530
rect 1196 1527 1197 1528
rect 638 1526 644 1527
rect 686 1526 692 1527
rect 703 1526 709 1527
rect 774 1526 780 1527
rect 791 1526 797 1527
rect 870 1526 876 1527
rect 887 1526 893 1527
rect 974 1526 980 1527
rect 991 1526 997 1527
rect 1078 1526 1084 1527
rect 1094 1526 1101 1527
rect 1174 1526 1180 1527
rect 1186 1526 1197 1527
rect 1214 1527 1215 1528
rect 1219 1527 1220 1531
rect 1254 1531 1255 1535
rect 1259 1534 1260 1535
rect 1259 1532 1282 1534
rect 1259 1531 1260 1532
rect 1254 1530 1260 1531
rect 1280 1530 1282 1532
rect 1287 1531 1293 1532
rect 1287 1530 1288 1531
rect 1280 1528 1288 1530
rect 1287 1527 1288 1528
rect 1292 1527 1293 1531
rect 1374 1531 1381 1532
rect 1374 1527 1375 1531
rect 1380 1527 1381 1531
rect 1446 1531 1452 1532
rect 1446 1527 1447 1531
rect 1451 1530 1452 1531
rect 1455 1531 1461 1532
rect 1455 1530 1456 1531
rect 1451 1528 1456 1530
rect 1451 1527 1452 1528
rect 1214 1526 1220 1527
rect 1270 1526 1276 1527
rect 1287 1526 1293 1527
rect 1358 1526 1364 1527
rect 1374 1526 1381 1527
rect 1438 1526 1444 1527
rect 1446 1526 1452 1527
rect 1455 1527 1456 1528
rect 1460 1527 1461 1531
rect 1535 1531 1541 1532
rect 1535 1527 1536 1531
rect 1540 1530 1541 1531
rect 1546 1531 1552 1532
rect 1546 1530 1547 1531
rect 1540 1528 1547 1530
rect 1540 1527 1541 1528
rect 1455 1526 1461 1527
rect 1518 1526 1524 1527
rect 1535 1526 1541 1527
rect 1546 1527 1547 1528
rect 1551 1527 1552 1531
rect 1615 1531 1621 1532
rect 1615 1527 1616 1531
rect 1620 1530 1621 1531
rect 1670 1531 1677 1532
rect 1620 1528 1650 1530
rect 1620 1527 1621 1528
rect 1546 1526 1552 1527
rect 1598 1526 1604 1527
rect 1615 1526 1621 1527
rect 462 1522 463 1526
rect 467 1522 468 1526
rect 462 1521 468 1522
rect 534 1522 535 1526
rect 539 1522 540 1526
rect 534 1521 540 1522
rect 606 1522 607 1526
rect 611 1522 612 1526
rect 606 1521 612 1522
rect 686 1522 687 1526
rect 691 1522 692 1526
rect 686 1521 692 1522
rect 774 1522 775 1526
rect 779 1522 780 1526
rect 774 1521 780 1522
rect 870 1522 871 1526
rect 875 1522 876 1526
rect 870 1521 876 1522
rect 974 1522 975 1526
rect 979 1522 980 1526
rect 974 1521 980 1522
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1102 1523 1108 1524
rect 1102 1522 1103 1523
rect 1078 1521 1084 1522
rect 1097 1520 1103 1522
rect 1097 1516 1099 1520
rect 1102 1519 1103 1520
rect 1107 1519 1108 1523
rect 1174 1522 1175 1526
rect 1179 1522 1180 1526
rect 1174 1521 1180 1522
rect 1270 1522 1271 1526
rect 1275 1522 1276 1526
rect 1270 1521 1276 1522
rect 1358 1522 1359 1526
rect 1363 1522 1364 1526
rect 1358 1521 1364 1522
rect 1438 1522 1439 1526
rect 1443 1522 1444 1526
rect 1438 1521 1444 1522
rect 1518 1522 1519 1526
rect 1523 1522 1524 1526
rect 1518 1521 1524 1522
rect 1598 1522 1599 1526
rect 1603 1522 1604 1526
rect 1598 1521 1604 1522
rect 1102 1518 1108 1519
rect 1648 1518 1650 1528
rect 1670 1527 1671 1531
rect 1676 1527 1677 1531
rect 1654 1526 1660 1527
rect 1670 1526 1677 1527
rect 1694 1528 1700 1529
rect 1654 1522 1655 1526
rect 1659 1522 1660 1526
rect 1694 1524 1695 1528
rect 1699 1524 1700 1528
rect 1694 1523 1700 1524
rect 1654 1521 1660 1522
rect 1648 1516 1654 1518
rect 415 1515 421 1516
rect 415 1514 416 1515
rect 408 1512 416 1514
rect 350 1510 357 1511
rect 415 1511 416 1512
rect 420 1511 421 1515
rect 415 1510 421 1511
rect 479 1515 485 1516
rect 479 1511 480 1515
rect 484 1514 485 1515
rect 487 1515 493 1516
rect 487 1514 488 1515
rect 484 1512 488 1514
rect 484 1511 485 1512
rect 479 1510 485 1511
rect 487 1511 488 1512
rect 492 1511 493 1515
rect 487 1510 493 1511
rect 551 1515 560 1516
rect 551 1511 552 1515
rect 559 1511 560 1515
rect 551 1510 560 1511
rect 623 1515 629 1516
rect 623 1511 624 1515
rect 628 1514 629 1515
rect 646 1515 652 1516
rect 646 1514 647 1515
rect 628 1512 647 1514
rect 628 1511 629 1512
rect 623 1510 629 1511
rect 646 1511 647 1512
rect 651 1511 652 1515
rect 646 1510 652 1511
rect 703 1515 709 1516
rect 703 1511 704 1515
rect 708 1514 709 1515
rect 718 1515 724 1516
rect 718 1514 719 1515
rect 708 1512 719 1514
rect 708 1511 709 1512
rect 703 1510 709 1511
rect 718 1511 719 1512
rect 723 1511 724 1515
rect 718 1510 724 1511
rect 791 1515 797 1516
rect 791 1511 792 1515
rect 796 1514 797 1515
rect 799 1515 805 1516
rect 799 1514 800 1515
rect 796 1512 800 1514
rect 796 1511 797 1512
rect 791 1510 797 1511
rect 799 1511 800 1512
rect 804 1511 805 1515
rect 799 1510 805 1511
rect 887 1515 893 1516
rect 887 1511 888 1515
rect 892 1514 893 1515
rect 895 1515 901 1516
rect 895 1514 896 1515
rect 892 1512 896 1514
rect 892 1511 893 1512
rect 887 1510 893 1511
rect 895 1511 896 1512
rect 900 1511 901 1515
rect 895 1510 901 1511
rect 990 1515 997 1516
rect 990 1511 991 1515
rect 996 1511 997 1515
rect 990 1510 997 1511
rect 1095 1515 1101 1516
rect 1095 1511 1096 1515
rect 1100 1511 1101 1515
rect 1095 1510 1101 1511
rect 1191 1515 1200 1516
rect 1191 1511 1192 1515
rect 1199 1511 1200 1515
rect 1191 1510 1200 1511
rect 1287 1515 1293 1516
rect 1287 1511 1288 1515
rect 1292 1514 1293 1515
rect 1334 1515 1340 1516
rect 1334 1514 1335 1515
rect 1292 1512 1335 1514
rect 1292 1511 1293 1512
rect 1287 1510 1293 1511
rect 1334 1511 1335 1512
rect 1339 1511 1340 1515
rect 1334 1510 1340 1511
rect 1374 1515 1381 1516
rect 1374 1511 1375 1515
rect 1380 1511 1381 1515
rect 1374 1510 1381 1511
rect 1455 1515 1461 1516
rect 1455 1511 1456 1515
rect 1460 1514 1461 1515
rect 1478 1515 1484 1516
rect 1478 1514 1479 1515
rect 1460 1512 1479 1514
rect 1460 1511 1461 1512
rect 1455 1510 1461 1511
rect 1478 1511 1479 1512
rect 1483 1511 1484 1515
rect 1535 1515 1541 1516
rect 1535 1514 1536 1515
rect 1478 1510 1484 1511
rect 1528 1512 1536 1514
rect 110 1506 116 1507
rect 134 1509 140 1510
rect 134 1505 135 1509
rect 139 1505 140 1509
rect 134 1504 140 1505
rect 174 1509 180 1510
rect 174 1505 175 1509
rect 179 1505 180 1509
rect 174 1504 180 1505
rect 222 1509 228 1510
rect 222 1505 223 1509
rect 227 1505 228 1509
rect 222 1504 228 1505
rect 278 1509 284 1510
rect 278 1505 279 1509
rect 283 1505 284 1509
rect 278 1504 284 1505
rect 334 1509 340 1510
rect 334 1505 335 1509
rect 339 1505 340 1509
rect 334 1504 340 1505
rect 398 1509 404 1510
rect 398 1505 399 1509
rect 403 1505 404 1509
rect 398 1504 404 1505
rect 462 1509 468 1510
rect 462 1505 463 1509
rect 467 1505 468 1509
rect 462 1504 468 1505
rect 534 1509 540 1510
rect 534 1505 535 1509
rect 539 1505 540 1509
rect 534 1504 540 1505
rect 606 1509 612 1510
rect 606 1505 607 1509
rect 611 1505 612 1509
rect 606 1504 612 1505
rect 686 1509 692 1510
rect 686 1505 687 1509
rect 691 1505 692 1509
rect 686 1504 692 1505
rect 774 1509 780 1510
rect 774 1505 775 1509
rect 779 1505 780 1509
rect 774 1504 780 1505
rect 870 1509 876 1510
rect 870 1505 871 1509
rect 875 1505 876 1509
rect 870 1504 876 1505
rect 974 1509 980 1510
rect 974 1505 975 1509
rect 979 1505 980 1509
rect 974 1504 980 1505
rect 1078 1509 1084 1510
rect 1078 1505 1079 1509
rect 1083 1505 1084 1509
rect 1078 1504 1084 1505
rect 1174 1509 1180 1510
rect 1174 1505 1175 1509
rect 1179 1505 1180 1509
rect 1174 1504 1180 1505
rect 1270 1509 1276 1510
rect 1270 1505 1271 1509
rect 1275 1505 1276 1509
rect 1270 1504 1276 1505
rect 1358 1509 1364 1510
rect 1358 1505 1359 1509
rect 1363 1505 1364 1509
rect 1358 1504 1364 1505
rect 1438 1509 1444 1510
rect 1438 1505 1439 1509
rect 1443 1505 1444 1509
rect 1438 1504 1444 1505
rect 1518 1509 1524 1510
rect 1518 1505 1519 1509
rect 1523 1505 1524 1509
rect 1518 1504 1524 1505
rect 102 1502 108 1503
rect 1498 1503 1504 1504
rect 1498 1499 1499 1503
rect 1503 1502 1504 1503
rect 1528 1502 1530 1512
rect 1535 1511 1536 1512
rect 1540 1511 1541 1515
rect 1535 1510 1541 1511
rect 1615 1515 1621 1516
rect 1615 1511 1616 1515
rect 1620 1514 1621 1515
rect 1638 1515 1644 1516
rect 1638 1514 1639 1515
rect 1620 1512 1639 1514
rect 1620 1511 1621 1512
rect 1615 1510 1621 1511
rect 1638 1511 1639 1512
rect 1643 1511 1644 1515
rect 1652 1514 1666 1516
rect 1671 1515 1677 1516
rect 1671 1514 1672 1515
rect 1664 1512 1672 1514
rect 1638 1510 1644 1511
rect 1671 1511 1672 1512
rect 1676 1511 1677 1515
rect 1671 1510 1677 1511
rect 1694 1511 1700 1512
rect 1598 1509 1604 1510
rect 1598 1505 1599 1509
rect 1603 1505 1604 1509
rect 1598 1504 1604 1505
rect 1654 1509 1660 1510
rect 1654 1505 1655 1509
rect 1659 1505 1660 1509
rect 1694 1507 1695 1511
rect 1699 1507 1700 1511
rect 1694 1506 1700 1507
rect 1654 1504 1660 1505
rect 1503 1500 1530 1502
rect 1503 1499 1504 1500
rect 1498 1498 1504 1499
rect 859 1491 865 1492
rect 859 1487 860 1491
rect 864 1490 865 1491
rect 918 1491 924 1492
rect 918 1490 919 1491
rect 864 1488 919 1490
rect 864 1487 865 1488
rect 859 1486 865 1487
rect 918 1487 919 1488
rect 923 1487 924 1491
rect 918 1486 924 1487
rect 987 1491 993 1492
rect 987 1487 988 1491
rect 992 1490 993 1491
rect 1146 1491 1152 1492
rect 1146 1490 1147 1491
rect 992 1488 1147 1490
rect 992 1487 993 1488
rect 987 1486 993 1487
rect 1146 1487 1147 1488
rect 1151 1487 1152 1491
rect 1146 1486 1152 1487
rect 382 1483 388 1484
rect 382 1482 383 1483
rect 321 1480 383 1482
rect 174 1475 180 1476
rect 110 1473 116 1474
rect 110 1469 111 1473
rect 115 1469 116 1473
rect 174 1471 175 1475
rect 179 1471 180 1475
rect 174 1470 180 1471
rect 206 1475 212 1476
rect 206 1471 207 1475
rect 211 1471 212 1475
rect 206 1470 212 1471
rect 238 1475 244 1476
rect 238 1471 239 1475
rect 243 1471 244 1475
rect 238 1470 244 1471
rect 270 1475 276 1476
rect 270 1471 271 1475
rect 275 1471 276 1475
rect 270 1470 276 1471
rect 302 1475 308 1476
rect 302 1471 303 1475
rect 307 1471 308 1475
rect 302 1470 308 1471
rect 110 1468 116 1469
rect 321 1468 323 1480
rect 382 1479 383 1480
rect 387 1479 388 1483
rect 470 1483 476 1484
rect 470 1482 471 1483
rect 382 1478 388 1479
rect 408 1480 471 1482
rect 334 1475 340 1476
rect 334 1471 335 1475
rect 339 1471 340 1475
rect 334 1470 340 1471
rect 366 1475 372 1476
rect 366 1471 367 1475
rect 371 1471 372 1475
rect 366 1470 372 1471
rect 398 1475 404 1476
rect 398 1471 399 1475
rect 403 1471 404 1475
rect 398 1470 404 1471
rect 150 1467 156 1468
rect 150 1463 151 1467
rect 155 1466 156 1467
rect 191 1467 197 1468
rect 191 1466 192 1467
rect 155 1464 192 1466
rect 155 1463 156 1464
rect 150 1462 156 1463
rect 191 1463 192 1464
rect 196 1463 197 1467
rect 223 1467 229 1468
rect 223 1466 224 1467
rect 191 1462 197 1463
rect 216 1464 224 1466
rect 174 1458 180 1459
rect 110 1456 116 1457
rect 110 1452 111 1456
rect 115 1452 116 1456
rect 174 1454 175 1458
rect 179 1454 180 1458
rect 174 1453 180 1454
rect 206 1458 212 1459
rect 206 1454 207 1458
rect 211 1454 212 1458
rect 206 1453 212 1454
rect 110 1451 116 1452
rect 191 1451 197 1452
rect 191 1447 192 1451
rect 196 1450 197 1451
rect 216 1450 218 1464
rect 223 1463 224 1464
rect 228 1463 229 1467
rect 255 1467 261 1468
rect 255 1466 256 1467
rect 223 1462 229 1463
rect 248 1464 256 1466
rect 238 1458 244 1459
rect 238 1454 239 1458
rect 243 1454 244 1458
rect 238 1453 244 1454
rect 196 1448 218 1450
rect 223 1451 229 1452
rect 196 1447 197 1448
rect 191 1446 197 1447
rect 223 1447 224 1451
rect 228 1450 229 1451
rect 248 1450 250 1464
rect 255 1463 256 1464
rect 260 1463 261 1467
rect 287 1467 293 1468
rect 287 1466 288 1467
rect 255 1462 261 1463
rect 280 1464 288 1466
rect 270 1458 276 1459
rect 270 1454 271 1458
rect 275 1454 276 1458
rect 270 1453 276 1454
rect 228 1448 250 1450
rect 255 1451 261 1452
rect 228 1447 229 1448
rect 223 1446 229 1447
rect 255 1447 256 1451
rect 260 1450 261 1451
rect 280 1450 282 1464
rect 287 1463 288 1464
rect 292 1463 293 1467
rect 287 1462 293 1463
rect 319 1467 325 1468
rect 319 1463 320 1467
rect 324 1463 325 1467
rect 351 1467 357 1468
rect 351 1466 352 1467
rect 319 1462 325 1463
rect 328 1464 352 1466
rect 302 1458 308 1459
rect 328 1458 330 1464
rect 351 1463 352 1464
rect 356 1463 357 1467
rect 351 1462 357 1463
rect 383 1467 389 1468
rect 383 1463 384 1467
rect 388 1466 389 1467
rect 408 1466 410 1480
rect 470 1479 471 1480
rect 475 1479 476 1483
rect 470 1478 476 1479
rect 806 1476 812 1477
rect 430 1475 436 1476
rect 430 1471 431 1475
rect 435 1471 436 1475
rect 430 1470 436 1471
rect 462 1475 468 1476
rect 462 1471 463 1475
rect 467 1471 468 1475
rect 462 1470 468 1471
rect 494 1475 500 1476
rect 494 1471 495 1475
rect 499 1471 500 1475
rect 494 1470 500 1471
rect 526 1475 532 1476
rect 526 1471 527 1475
rect 531 1471 532 1475
rect 526 1470 532 1471
rect 558 1475 564 1476
rect 558 1471 559 1475
rect 563 1471 564 1475
rect 558 1470 564 1471
rect 590 1475 596 1476
rect 590 1471 591 1475
rect 595 1471 596 1475
rect 590 1470 596 1471
rect 622 1475 628 1476
rect 622 1471 623 1475
rect 627 1471 628 1475
rect 622 1470 628 1471
rect 662 1475 668 1476
rect 662 1471 663 1475
rect 667 1471 668 1475
rect 662 1470 668 1471
rect 702 1475 708 1476
rect 702 1471 703 1475
rect 707 1471 708 1475
rect 702 1470 708 1471
rect 742 1475 748 1476
rect 742 1471 743 1475
rect 747 1471 748 1475
rect 742 1470 748 1471
rect 774 1475 780 1476
rect 774 1471 775 1475
rect 779 1471 780 1475
rect 806 1472 807 1476
rect 811 1472 812 1476
rect 806 1471 812 1472
rect 894 1476 900 1477
rect 894 1472 895 1476
rect 899 1472 900 1476
rect 894 1471 900 1472
rect 934 1476 940 1477
rect 934 1472 935 1476
rect 939 1472 940 1476
rect 934 1471 940 1472
rect 1022 1476 1028 1477
rect 1110 1476 1116 1477
rect 1022 1472 1023 1476
rect 1027 1472 1028 1476
rect 1022 1471 1028 1472
rect 1078 1475 1084 1476
rect 1078 1471 1079 1475
rect 1083 1471 1084 1475
rect 1110 1472 1111 1476
rect 1115 1472 1116 1476
rect 1110 1471 1116 1472
rect 1166 1475 1172 1476
rect 1166 1471 1167 1475
rect 1171 1471 1172 1475
rect 774 1470 780 1471
rect 1078 1470 1084 1471
rect 1166 1470 1172 1471
rect 1198 1475 1204 1476
rect 1198 1471 1199 1475
rect 1203 1471 1204 1475
rect 1198 1470 1204 1471
rect 1238 1475 1244 1476
rect 1238 1471 1239 1475
rect 1243 1471 1244 1475
rect 1238 1470 1244 1471
rect 1278 1475 1284 1476
rect 1278 1471 1279 1475
rect 1283 1471 1284 1475
rect 1278 1470 1284 1471
rect 1318 1475 1324 1476
rect 1318 1471 1319 1475
rect 1323 1471 1324 1475
rect 1318 1470 1324 1471
rect 1358 1475 1364 1476
rect 1358 1471 1359 1475
rect 1363 1471 1364 1475
rect 1358 1470 1364 1471
rect 1398 1475 1404 1476
rect 1398 1471 1399 1475
rect 1403 1471 1404 1475
rect 1398 1470 1404 1471
rect 1438 1475 1444 1476
rect 1438 1471 1439 1475
rect 1443 1471 1444 1475
rect 1438 1470 1444 1471
rect 1478 1475 1484 1476
rect 1478 1471 1479 1475
rect 1483 1471 1484 1475
rect 1478 1470 1484 1471
rect 1518 1475 1524 1476
rect 1518 1471 1519 1475
rect 1523 1471 1524 1475
rect 1518 1470 1524 1471
rect 1558 1475 1564 1476
rect 1558 1471 1559 1475
rect 1563 1471 1564 1475
rect 1558 1470 1564 1471
rect 1590 1475 1596 1476
rect 1590 1471 1591 1475
rect 1595 1471 1596 1475
rect 1590 1470 1596 1471
rect 1622 1475 1628 1476
rect 1622 1471 1623 1475
rect 1627 1471 1628 1475
rect 1622 1470 1628 1471
rect 1654 1475 1660 1476
rect 1654 1471 1655 1475
rect 1659 1471 1660 1475
rect 1654 1470 1660 1471
rect 1694 1473 1700 1474
rect 1694 1469 1695 1473
rect 1699 1469 1700 1473
rect 1694 1468 1700 1469
rect 388 1464 410 1466
rect 415 1467 421 1468
rect 388 1463 389 1464
rect 383 1462 389 1463
rect 415 1463 416 1467
rect 420 1466 421 1467
rect 446 1467 453 1468
rect 420 1464 442 1466
rect 420 1463 421 1464
rect 415 1462 421 1463
rect 302 1454 303 1458
rect 307 1454 308 1458
rect 302 1453 308 1454
rect 312 1456 330 1458
rect 334 1458 340 1459
rect 260 1448 282 1450
rect 287 1451 293 1452
rect 260 1447 261 1448
rect 255 1446 261 1447
rect 287 1447 288 1451
rect 292 1450 293 1451
rect 312 1450 314 1456
rect 334 1454 335 1458
rect 339 1454 340 1458
rect 334 1453 340 1454
rect 366 1458 372 1459
rect 366 1454 367 1458
rect 371 1454 372 1458
rect 366 1453 372 1454
rect 398 1458 404 1459
rect 398 1454 399 1458
rect 403 1454 404 1458
rect 398 1453 404 1454
rect 430 1458 436 1459
rect 430 1454 431 1458
rect 435 1454 436 1458
rect 430 1453 436 1454
rect 292 1448 314 1450
rect 318 1451 325 1452
rect 292 1447 293 1448
rect 287 1446 293 1447
rect 318 1447 319 1451
rect 324 1447 325 1451
rect 318 1446 325 1447
rect 350 1451 357 1452
rect 350 1447 351 1451
rect 356 1447 357 1451
rect 350 1446 357 1447
rect 382 1451 389 1452
rect 382 1447 383 1451
rect 388 1447 389 1451
rect 382 1446 389 1447
rect 415 1451 421 1452
rect 415 1447 416 1451
rect 420 1447 421 1451
rect 440 1450 442 1464
rect 446 1463 447 1467
rect 452 1463 453 1467
rect 446 1462 453 1463
rect 455 1467 461 1468
rect 455 1463 456 1467
rect 460 1466 461 1467
rect 479 1467 485 1468
rect 479 1466 480 1467
rect 460 1464 480 1466
rect 460 1463 461 1464
rect 455 1462 461 1463
rect 479 1463 480 1464
rect 484 1463 485 1467
rect 511 1467 517 1468
rect 511 1466 512 1467
rect 479 1462 485 1463
rect 504 1464 512 1466
rect 462 1458 468 1459
rect 462 1454 463 1458
rect 467 1454 468 1458
rect 462 1453 468 1454
rect 494 1458 500 1459
rect 494 1454 495 1458
rect 499 1454 500 1458
rect 494 1453 500 1454
rect 447 1451 453 1452
rect 447 1450 448 1451
rect 440 1448 448 1450
rect 415 1446 421 1447
rect 447 1447 448 1448
rect 452 1447 453 1451
rect 447 1446 453 1447
rect 479 1451 485 1452
rect 479 1447 480 1451
rect 484 1450 485 1451
rect 504 1450 506 1464
rect 511 1463 512 1464
rect 516 1463 517 1467
rect 511 1462 517 1463
rect 542 1467 549 1468
rect 542 1463 543 1467
rect 548 1463 549 1467
rect 575 1467 581 1468
rect 575 1466 576 1467
rect 542 1462 549 1463
rect 568 1464 576 1466
rect 526 1458 532 1459
rect 526 1454 527 1458
rect 531 1454 532 1458
rect 526 1453 532 1454
rect 558 1458 564 1459
rect 558 1454 559 1458
rect 563 1454 564 1458
rect 558 1453 564 1454
rect 484 1448 506 1450
rect 511 1451 517 1452
rect 484 1447 485 1448
rect 479 1446 485 1447
rect 511 1447 512 1451
rect 516 1450 517 1451
rect 534 1451 540 1452
rect 534 1450 535 1451
rect 516 1448 535 1450
rect 516 1447 517 1448
rect 511 1446 517 1447
rect 534 1447 535 1448
rect 539 1447 540 1451
rect 534 1446 540 1447
rect 543 1451 549 1452
rect 543 1447 544 1451
rect 548 1450 549 1451
rect 568 1450 570 1464
rect 575 1463 576 1464
rect 580 1463 581 1467
rect 607 1467 613 1468
rect 607 1466 608 1467
rect 575 1462 581 1463
rect 600 1464 608 1466
rect 590 1458 596 1459
rect 590 1454 591 1458
rect 595 1454 596 1458
rect 590 1453 596 1454
rect 548 1448 570 1450
rect 575 1451 581 1452
rect 548 1447 549 1448
rect 543 1446 549 1447
rect 575 1447 576 1451
rect 580 1450 581 1451
rect 600 1450 602 1464
rect 607 1463 608 1464
rect 612 1463 613 1467
rect 607 1462 613 1463
rect 638 1467 645 1468
rect 638 1463 639 1467
rect 644 1463 645 1467
rect 638 1462 645 1463
rect 679 1467 688 1468
rect 679 1463 680 1467
rect 687 1463 688 1467
rect 719 1467 725 1468
rect 719 1466 720 1467
rect 679 1462 688 1463
rect 696 1464 720 1466
rect 622 1458 628 1459
rect 622 1454 623 1458
rect 627 1454 628 1458
rect 622 1453 628 1454
rect 662 1458 668 1459
rect 662 1454 663 1458
rect 667 1454 668 1458
rect 662 1453 668 1454
rect 580 1448 602 1450
rect 607 1451 613 1452
rect 580 1447 581 1448
rect 575 1446 581 1447
rect 607 1447 608 1451
rect 612 1447 613 1451
rect 607 1446 613 1447
rect 639 1451 645 1452
rect 639 1447 640 1451
rect 644 1447 645 1451
rect 639 1446 645 1447
rect 679 1451 685 1452
rect 679 1447 680 1451
rect 684 1450 685 1451
rect 696 1450 698 1464
rect 719 1463 720 1464
rect 724 1463 725 1467
rect 719 1462 725 1463
rect 727 1467 733 1468
rect 727 1463 728 1467
rect 732 1466 733 1467
rect 759 1467 765 1468
rect 759 1466 760 1467
rect 732 1464 760 1466
rect 732 1463 733 1464
rect 727 1462 733 1463
rect 759 1463 760 1464
rect 764 1463 765 1467
rect 759 1462 765 1463
rect 767 1467 773 1468
rect 767 1463 768 1467
rect 772 1466 773 1467
rect 791 1467 797 1468
rect 791 1466 792 1467
rect 772 1464 792 1466
rect 772 1463 773 1464
rect 767 1462 773 1463
rect 791 1463 792 1464
rect 796 1463 797 1467
rect 886 1467 892 1468
rect 791 1462 797 1463
rect 801 1464 849 1466
rect 702 1458 708 1459
rect 702 1454 703 1458
rect 707 1454 708 1458
rect 702 1453 708 1454
rect 742 1458 748 1459
rect 742 1454 743 1458
rect 747 1454 748 1458
rect 742 1453 748 1454
rect 774 1457 780 1458
rect 774 1453 775 1457
rect 779 1453 780 1457
rect 774 1452 780 1453
rect 684 1448 698 1450
rect 718 1451 725 1452
rect 684 1447 685 1448
rect 679 1446 685 1447
rect 718 1447 719 1451
rect 724 1447 725 1451
rect 718 1446 725 1447
rect 759 1451 765 1452
rect 759 1447 760 1451
rect 764 1447 765 1451
rect 759 1446 765 1447
rect 791 1451 797 1452
rect 791 1447 792 1451
rect 796 1450 797 1451
rect 801 1450 803 1464
rect 886 1463 887 1467
rect 891 1466 892 1467
rect 1094 1467 1101 1468
rect 891 1464 977 1466
rect 891 1463 892 1464
rect 886 1462 892 1463
rect 1094 1463 1095 1467
rect 1100 1463 1101 1467
rect 1094 1462 1101 1463
rect 1183 1467 1189 1468
rect 1183 1463 1184 1467
rect 1188 1466 1189 1467
rect 1215 1467 1221 1468
rect 1188 1464 1210 1466
rect 1188 1463 1189 1464
rect 1183 1462 1189 1463
rect 918 1459 925 1460
rect 806 1457 812 1458
rect 806 1453 807 1457
rect 811 1453 812 1457
rect 918 1455 919 1459
rect 924 1455 925 1459
rect 1078 1458 1084 1459
rect 918 1454 925 1455
rect 934 1457 940 1458
rect 806 1452 812 1453
rect 934 1453 935 1457
rect 939 1453 940 1457
rect 934 1452 940 1453
rect 1038 1455 1044 1456
rect 1038 1451 1039 1455
rect 1043 1451 1044 1455
rect 1059 1455 1065 1456
rect 1059 1454 1060 1455
rect 1038 1450 1044 1451
rect 1048 1452 1060 1454
rect 796 1448 803 1450
rect 894 1448 900 1449
rect 796 1447 797 1448
rect 791 1446 797 1447
rect 417 1442 419 1446
rect 455 1443 461 1444
rect 455 1442 456 1443
rect 417 1440 456 1442
rect 455 1439 456 1440
rect 460 1439 461 1443
rect 455 1438 461 1439
rect 609 1434 611 1446
rect 641 1442 643 1446
rect 703 1443 709 1444
rect 703 1442 704 1443
rect 641 1440 704 1442
rect 703 1439 704 1440
rect 708 1439 709 1443
rect 761 1442 763 1446
rect 894 1444 895 1448
rect 899 1444 900 1448
rect 1048 1446 1050 1452
rect 1059 1451 1060 1452
rect 1064 1451 1065 1455
rect 1078 1454 1079 1458
rect 1083 1454 1084 1458
rect 1166 1458 1172 1459
rect 1078 1453 1084 1454
rect 1126 1455 1132 1456
rect 1059 1450 1065 1451
rect 1095 1451 1101 1452
rect 1095 1447 1096 1451
rect 1100 1447 1101 1451
rect 1126 1451 1127 1455
rect 1131 1451 1132 1455
rect 1126 1450 1132 1451
rect 1146 1455 1153 1456
rect 1146 1451 1147 1455
rect 1152 1451 1153 1455
rect 1166 1454 1167 1458
rect 1171 1454 1172 1458
rect 1166 1453 1172 1454
rect 1198 1458 1204 1459
rect 1198 1454 1199 1458
rect 1203 1454 1204 1458
rect 1208 1458 1210 1464
rect 1215 1463 1216 1467
rect 1220 1466 1221 1467
rect 1230 1467 1236 1468
rect 1230 1466 1231 1467
rect 1220 1464 1231 1466
rect 1220 1463 1221 1464
rect 1215 1462 1221 1463
rect 1230 1463 1231 1464
rect 1235 1463 1236 1467
rect 1230 1462 1236 1463
rect 1254 1467 1261 1468
rect 1254 1463 1255 1467
rect 1260 1463 1261 1467
rect 1254 1462 1261 1463
rect 1263 1467 1269 1468
rect 1263 1463 1264 1467
rect 1268 1466 1269 1467
rect 1295 1467 1301 1468
rect 1295 1466 1296 1467
rect 1268 1464 1296 1466
rect 1268 1463 1269 1464
rect 1263 1462 1269 1463
rect 1295 1463 1296 1464
rect 1300 1463 1301 1467
rect 1295 1462 1301 1463
rect 1335 1467 1341 1468
rect 1335 1463 1336 1467
rect 1340 1466 1341 1467
rect 1375 1467 1381 1468
rect 1340 1464 1370 1466
rect 1340 1463 1341 1464
rect 1335 1462 1341 1463
rect 1238 1458 1244 1459
rect 1318 1458 1324 1459
rect 1208 1456 1226 1458
rect 1198 1453 1204 1454
rect 1146 1450 1153 1451
rect 1182 1451 1189 1452
rect 1095 1446 1101 1447
rect 1138 1447 1144 1448
rect 1138 1446 1139 1447
rect 814 1443 820 1444
rect 814 1442 815 1443
rect 761 1440 815 1442
rect 703 1438 709 1439
rect 814 1439 815 1440
rect 819 1439 820 1443
rect 886 1443 892 1444
rect 894 1443 900 1444
rect 1012 1444 1050 1446
rect 1097 1444 1139 1446
rect 886 1442 887 1443
rect 872 1440 887 1442
rect 814 1438 820 1439
rect 855 1439 861 1440
rect 727 1435 733 1436
rect 727 1434 728 1435
rect 609 1432 728 1434
rect 727 1431 728 1432
rect 732 1431 733 1435
rect 855 1435 856 1439
rect 860 1438 861 1439
rect 872 1438 874 1440
rect 886 1439 887 1440
rect 891 1439 892 1443
rect 886 1438 892 1439
rect 919 1439 925 1440
rect 860 1436 874 1438
rect 860 1435 861 1436
rect 855 1434 861 1435
rect 891 1435 897 1436
rect 727 1430 733 1431
rect 767 1431 773 1432
rect 767 1430 768 1431
rect 736 1428 768 1430
rect 534 1427 540 1428
rect 534 1423 535 1427
rect 539 1426 540 1427
rect 670 1427 676 1428
rect 670 1426 671 1427
rect 539 1424 671 1426
rect 539 1423 540 1424
rect 534 1422 540 1423
rect 670 1423 671 1424
rect 675 1426 676 1427
rect 736 1426 738 1428
rect 767 1427 768 1428
rect 772 1427 773 1431
rect 891 1431 892 1435
rect 896 1434 897 1435
rect 910 1435 916 1436
rect 910 1434 911 1435
rect 896 1432 911 1434
rect 896 1431 897 1432
rect 891 1430 897 1431
rect 910 1431 911 1432
rect 915 1431 916 1435
rect 919 1435 920 1439
rect 924 1435 925 1439
rect 919 1434 925 1435
rect 983 1439 989 1440
rect 983 1435 984 1439
rect 988 1438 989 1439
rect 1012 1438 1014 1444
rect 1138 1443 1139 1444
rect 1143 1443 1144 1447
rect 1182 1447 1183 1451
rect 1188 1447 1189 1451
rect 1182 1446 1189 1447
rect 1214 1451 1221 1452
rect 1214 1447 1215 1451
rect 1220 1447 1221 1451
rect 1224 1450 1226 1456
rect 1238 1454 1239 1458
rect 1243 1454 1244 1458
rect 1238 1453 1244 1454
rect 1278 1457 1284 1458
rect 1278 1453 1279 1457
rect 1283 1453 1284 1457
rect 1318 1454 1319 1458
rect 1323 1454 1324 1458
rect 1318 1453 1324 1454
rect 1358 1458 1364 1459
rect 1358 1454 1359 1458
rect 1363 1454 1364 1458
rect 1368 1458 1370 1464
rect 1375 1463 1376 1467
rect 1380 1466 1381 1467
rect 1383 1467 1389 1468
rect 1383 1466 1384 1467
rect 1380 1464 1384 1466
rect 1380 1463 1381 1464
rect 1375 1462 1381 1463
rect 1383 1463 1384 1464
rect 1388 1463 1389 1467
rect 1383 1462 1389 1463
rect 1415 1467 1421 1468
rect 1415 1463 1416 1467
rect 1420 1466 1421 1467
rect 1455 1467 1464 1468
rect 1420 1464 1434 1466
rect 1420 1463 1421 1464
rect 1415 1462 1421 1463
rect 1398 1458 1404 1459
rect 1368 1456 1386 1458
rect 1358 1453 1364 1454
rect 1278 1452 1284 1453
rect 1255 1451 1261 1452
rect 1255 1450 1256 1451
rect 1224 1448 1256 1450
rect 1214 1446 1221 1447
rect 1255 1447 1256 1448
rect 1260 1447 1261 1451
rect 1255 1446 1261 1447
rect 1295 1451 1304 1452
rect 1295 1447 1296 1451
rect 1303 1447 1304 1451
rect 1295 1446 1304 1447
rect 1334 1451 1341 1452
rect 1334 1447 1335 1451
rect 1340 1447 1341 1451
rect 1334 1446 1341 1447
rect 1374 1451 1381 1452
rect 1374 1447 1375 1451
rect 1380 1447 1381 1451
rect 1384 1450 1386 1456
rect 1398 1454 1399 1458
rect 1403 1454 1404 1458
rect 1398 1453 1404 1454
rect 1415 1451 1421 1452
rect 1415 1450 1416 1451
rect 1384 1448 1416 1450
rect 1374 1446 1381 1447
rect 1415 1447 1416 1448
rect 1420 1447 1421 1451
rect 1432 1450 1434 1464
rect 1455 1463 1456 1467
rect 1463 1463 1464 1467
rect 1455 1462 1464 1463
rect 1495 1467 1501 1468
rect 1495 1463 1496 1467
rect 1500 1466 1501 1467
rect 1535 1467 1541 1468
rect 1500 1464 1514 1466
rect 1500 1463 1501 1464
rect 1495 1462 1501 1463
rect 1438 1458 1444 1459
rect 1438 1454 1439 1458
rect 1443 1454 1444 1458
rect 1438 1453 1444 1454
rect 1478 1458 1484 1459
rect 1478 1454 1479 1458
rect 1483 1454 1484 1458
rect 1478 1453 1484 1454
rect 1455 1451 1461 1452
rect 1455 1450 1456 1451
rect 1432 1448 1456 1450
rect 1415 1446 1421 1447
rect 1455 1447 1456 1448
rect 1460 1447 1461 1451
rect 1455 1446 1461 1447
rect 1495 1451 1504 1452
rect 1495 1447 1496 1451
rect 1503 1447 1504 1451
rect 1512 1450 1514 1464
rect 1535 1463 1536 1467
rect 1540 1466 1541 1467
rect 1550 1467 1556 1468
rect 1550 1466 1551 1467
rect 1540 1464 1551 1466
rect 1540 1463 1541 1464
rect 1535 1462 1541 1463
rect 1550 1463 1551 1464
rect 1555 1463 1556 1467
rect 1550 1462 1556 1463
rect 1574 1467 1581 1468
rect 1574 1463 1575 1467
rect 1580 1463 1581 1467
rect 1607 1467 1613 1468
rect 1607 1466 1608 1467
rect 1574 1462 1581 1463
rect 1600 1464 1608 1466
rect 1518 1458 1524 1459
rect 1518 1454 1519 1458
rect 1523 1454 1524 1458
rect 1518 1453 1524 1454
rect 1558 1458 1564 1459
rect 1558 1454 1559 1458
rect 1563 1454 1564 1458
rect 1558 1453 1564 1454
rect 1590 1458 1596 1459
rect 1590 1454 1591 1458
rect 1595 1454 1596 1458
rect 1590 1453 1596 1454
rect 1535 1451 1541 1452
rect 1535 1450 1536 1451
rect 1512 1448 1536 1450
rect 1495 1446 1504 1447
rect 1535 1447 1536 1448
rect 1540 1447 1541 1451
rect 1535 1446 1541 1447
rect 1575 1451 1581 1452
rect 1575 1447 1576 1451
rect 1580 1450 1581 1451
rect 1600 1450 1602 1464
rect 1607 1463 1608 1464
rect 1612 1463 1613 1467
rect 1607 1462 1613 1463
rect 1639 1467 1645 1468
rect 1639 1463 1640 1467
rect 1644 1466 1645 1467
rect 1670 1467 1677 1468
rect 1644 1464 1666 1466
rect 1644 1463 1645 1464
rect 1639 1462 1645 1463
rect 1622 1458 1628 1459
rect 1622 1454 1623 1458
rect 1627 1454 1628 1458
rect 1622 1453 1628 1454
rect 1654 1458 1660 1459
rect 1654 1454 1655 1458
rect 1659 1454 1660 1458
rect 1654 1453 1660 1454
rect 1580 1448 1602 1450
rect 1607 1451 1613 1452
rect 1580 1447 1581 1448
rect 1575 1446 1581 1447
rect 1607 1447 1608 1451
rect 1612 1447 1613 1451
rect 1607 1446 1613 1447
rect 1638 1451 1645 1452
rect 1638 1447 1639 1451
rect 1644 1447 1645 1451
rect 1664 1450 1666 1464
rect 1670 1463 1671 1467
rect 1676 1463 1677 1467
rect 1670 1462 1677 1463
rect 1694 1456 1700 1457
rect 1694 1452 1695 1456
rect 1699 1452 1700 1456
rect 1671 1451 1677 1452
rect 1694 1451 1700 1452
rect 1671 1450 1672 1451
rect 1664 1448 1672 1450
rect 1638 1446 1645 1447
rect 1671 1447 1672 1448
rect 1676 1447 1677 1451
rect 1671 1446 1677 1447
rect 1138 1442 1144 1443
rect 1190 1443 1196 1444
rect 988 1436 1014 1438
rect 1043 1439 1052 1440
rect 988 1435 989 1436
rect 983 1434 989 1435
rect 1019 1435 1025 1436
rect 1019 1434 1020 1435
rect 910 1430 916 1431
rect 921 1430 923 1434
rect 1000 1432 1020 1434
rect 990 1431 996 1432
rect 990 1430 991 1431
rect 767 1426 773 1427
rect 796 1428 867 1430
rect 675 1424 738 1426
rect 796 1424 798 1428
rect 865 1426 867 1428
rect 893 1426 895 1430
rect 921 1428 991 1430
rect 990 1427 991 1428
rect 995 1427 996 1431
rect 990 1426 996 1427
rect 998 1431 1004 1432
rect 998 1427 999 1431
rect 1003 1427 1004 1431
rect 1019 1431 1020 1432
rect 1024 1434 1025 1435
rect 1030 1435 1036 1436
rect 1030 1434 1031 1435
rect 1024 1432 1031 1434
rect 1024 1431 1025 1432
rect 1019 1430 1025 1431
rect 1030 1431 1031 1432
rect 1035 1431 1036 1435
rect 1043 1435 1044 1439
rect 1051 1435 1052 1439
rect 1131 1439 1137 1440
rect 1043 1434 1052 1435
rect 1107 1435 1113 1436
rect 1030 1430 1036 1431
rect 1107 1431 1108 1435
rect 1112 1434 1113 1435
rect 1131 1435 1132 1439
rect 1136 1438 1137 1439
rect 1190 1439 1191 1443
rect 1195 1439 1196 1443
rect 1609 1442 1611 1446
rect 1670 1443 1676 1444
rect 1670 1442 1671 1443
rect 1609 1440 1671 1442
rect 1190 1438 1196 1439
rect 1670 1439 1671 1440
rect 1675 1439 1676 1443
rect 1670 1438 1676 1439
rect 1136 1436 1194 1438
rect 1136 1435 1137 1436
rect 1131 1434 1137 1435
rect 1702 1435 1708 1436
rect 1702 1434 1703 1435
rect 1112 1432 1126 1434
rect 1112 1431 1113 1432
rect 1107 1430 1113 1431
rect 1124 1430 1126 1432
rect 1159 1432 1703 1434
rect 1159 1430 1161 1432
rect 1702 1431 1703 1432
rect 1707 1431 1708 1435
rect 1702 1430 1708 1431
rect 1124 1428 1161 1430
rect 998 1426 1004 1427
rect 1190 1427 1196 1428
rect 865 1424 895 1426
rect 675 1423 676 1424
rect 670 1422 676 1423
rect 750 1423 756 1424
rect 750 1419 751 1423
rect 755 1422 756 1423
rect 763 1423 769 1424
rect 763 1422 764 1423
rect 755 1420 764 1422
rect 755 1419 756 1420
rect 750 1418 756 1419
rect 763 1419 764 1420
rect 768 1419 769 1423
rect 794 1423 800 1424
rect 794 1422 795 1423
rect 763 1418 769 1419
rect 791 1421 795 1422
rect 791 1417 792 1421
rect 799 1419 800 1423
rect 796 1418 800 1419
rect 830 1423 841 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 840 1419 841 1423
rect 865 1420 867 1424
rect 946 1423 952 1424
rect 830 1418 841 1419
rect 863 1419 869 1420
rect 796 1417 797 1418
rect 791 1416 797 1417
rect 766 1415 772 1416
rect 766 1411 767 1415
rect 771 1411 772 1415
rect 766 1410 772 1411
rect 838 1415 844 1416
rect 838 1411 839 1415
rect 843 1411 844 1415
rect 863 1415 864 1419
rect 868 1415 869 1419
rect 863 1414 869 1415
rect 878 1419 884 1420
rect 878 1415 879 1419
rect 883 1418 884 1419
rect 887 1419 893 1420
rect 887 1418 888 1419
rect 883 1416 888 1418
rect 883 1415 884 1416
rect 878 1414 884 1415
rect 887 1415 888 1416
rect 892 1415 893 1419
rect 887 1414 893 1415
rect 902 1419 909 1420
rect 902 1415 903 1419
rect 908 1415 909 1419
rect 902 1414 909 1415
rect 918 1419 925 1420
rect 918 1415 919 1419
rect 924 1415 925 1419
rect 946 1419 947 1423
rect 951 1422 952 1423
rect 971 1423 977 1424
rect 971 1422 972 1423
rect 951 1420 972 1422
rect 951 1419 952 1420
rect 946 1418 952 1419
rect 971 1419 972 1420
rect 976 1419 977 1423
rect 1190 1423 1191 1427
rect 1195 1426 1196 1427
rect 1195 1424 1274 1426
rect 1195 1423 1196 1424
rect 1190 1422 1196 1423
rect 1272 1422 1274 1424
rect 1470 1423 1476 1424
rect 1470 1422 1471 1423
rect 999 1420 1005 1421
rect 1272 1420 1471 1422
rect 971 1418 977 1419
rect 990 1419 996 1420
rect 918 1414 925 1415
rect 966 1415 972 1416
rect 966 1414 967 1415
rect 921 1412 967 1414
rect 966 1411 967 1412
rect 971 1411 972 1415
rect 838 1410 844 1411
rect 894 1410 900 1411
rect 966 1410 972 1411
rect 974 1415 980 1416
rect 974 1411 975 1415
rect 979 1411 980 1415
rect 990 1415 991 1419
rect 995 1418 996 1419
rect 999 1418 1000 1420
rect 995 1416 1000 1418
rect 1004 1418 1005 1420
rect 1122 1419 1128 1420
rect 1004 1416 1050 1418
rect 995 1415 996 1416
rect 999 1415 1005 1416
rect 1046 1415 1052 1416
rect 990 1414 996 1415
rect 974 1410 980 1411
rect 1046 1411 1047 1415
rect 1051 1414 1052 1415
rect 1122 1415 1123 1419
rect 1127 1418 1128 1419
rect 1214 1419 1220 1420
rect 1214 1418 1215 1419
rect 1127 1416 1215 1418
rect 1127 1415 1128 1416
rect 1122 1414 1128 1415
rect 1214 1415 1215 1416
rect 1219 1415 1220 1419
rect 1214 1414 1220 1415
rect 1051 1413 1098 1414
rect 1051 1412 1060 1413
rect 1051 1411 1052 1412
rect 1046 1410 1052 1411
rect 758 1407 764 1408
rect 446 1403 452 1404
rect 446 1399 447 1403
rect 451 1402 452 1403
rect 542 1403 548 1404
rect 451 1400 498 1402
rect 451 1399 452 1400
rect 446 1398 452 1399
rect 150 1395 157 1396
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 150 1391 151 1395
rect 156 1391 157 1395
rect 183 1395 189 1396
rect 183 1394 184 1395
rect 176 1392 184 1394
rect 110 1387 116 1388
rect 134 1390 140 1391
rect 150 1390 157 1391
rect 166 1390 172 1391
rect 134 1386 135 1390
rect 139 1386 140 1390
rect 134 1385 140 1386
rect 166 1386 167 1390
rect 171 1386 172 1390
rect 166 1385 172 1386
rect 176 1380 178 1392
rect 183 1391 184 1392
rect 188 1391 189 1395
rect 215 1395 221 1396
rect 215 1394 216 1395
rect 208 1392 216 1394
rect 183 1390 189 1391
rect 198 1390 204 1391
rect 198 1386 199 1390
rect 203 1386 204 1390
rect 198 1385 204 1386
rect 208 1380 210 1392
rect 215 1391 216 1392
rect 220 1391 221 1395
rect 247 1395 253 1396
rect 247 1394 248 1395
rect 240 1392 248 1394
rect 215 1390 221 1391
rect 230 1390 236 1391
rect 230 1386 231 1390
rect 235 1386 236 1390
rect 230 1385 236 1386
rect 240 1380 242 1392
rect 247 1391 248 1392
rect 252 1391 253 1395
rect 279 1395 285 1396
rect 279 1394 280 1395
rect 272 1392 280 1394
rect 247 1390 253 1391
rect 262 1390 268 1391
rect 262 1386 263 1390
rect 267 1386 268 1390
rect 262 1385 268 1386
rect 272 1380 274 1392
rect 279 1391 280 1392
rect 284 1391 285 1395
rect 311 1395 317 1396
rect 311 1394 312 1395
rect 304 1392 312 1394
rect 279 1390 285 1391
rect 294 1390 300 1391
rect 294 1386 295 1390
rect 299 1386 300 1390
rect 294 1385 300 1386
rect 304 1380 306 1392
rect 311 1391 312 1392
rect 316 1391 317 1395
rect 343 1395 349 1396
rect 343 1394 344 1395
rect 336 1392 344 1394
rect 311 1390 317 1391
rect 326 1390 332 1391
rect 326 1386 327 1390
rect 331 1386 332 1390
rect 326 1385 332 1386
rect 336 1380 338 1392
rect 343 1391 344 1392
rect 348 1391 349 1395
rect 375 1395 384 1396
rect 375 1391 376 1395
rect 383 1391 384 1395
rect 407 1395 413 1396
rect 407 1394 408 1395
rect 400 1392 408 1394
rect 343 1390 349 1391
rect 358 1390 364 1391
rect 375 1390 384 1391
rect 390 1390 396 1391
rect 358 1386 359 1390
rect 363 1386 364 1390
rect 358 1385 364 1386
rect 390 1386 391 1390
rect 395 1386 396 1390
rect 390 1385 396 1386
rect 400 1380 402 1392
rect 407 1391 408 1392
rect 412 1391 413 1395
rect 439 1395 445 1396
rect 439 1394 440 1395
rect 432 1392 440 1394
rect 407 1390 413 1391
rect 422 1390 428 1391
rect 422 1386 423 1390
rect 427 1386 428 1390
rect 422 1385 428 1386
rect 432 1380 434 1392
rect 439 1391 440 1392
rect 444 1391 445 1395
rect 471 1395 477 1396
rect 471 1394 472 1395
rect 464 1392 472 1394
rect 439 1390 445 1391
rect 454 1390 460 1391
rect 454 1386 455 1390
rect 459 1386 460 1390
rect 454 1385 460 1386
rect 464 1380 466 1392
rect 471 1391 472 1392
rect 476 1391 477 1395
rect 496 1394 498 1400
rect 542 1399 543 1403
rect 547 1402 548 1403
rect 719 1403 725 1404
rect 547 1400 594 1402
rect 547 1399 548 1400
rect 542 1398 548 1399
rect 503 1395 509 1396
rect 503 1394 504 1395
rect 496 1392 504 1394
rect 503 1391 504 1392
rect 508 1391 509 1395
rect 535 1395 541 1396
rect 535 1394 536 1395
rect 528 1392 536 1394
rect 471 1390 477 1391
rect 486 1390 492 1391
rect 503 1390 509 1391
rect 518 1390 524 1391
rect 486 1386 487 1390
rect 491 1386 492 1390
rect 486 1385 492 1386
rect 518 1386 519 1390
rect 523 1386 524 1390
rect 518 1385 524 1386
rect 528 1380 530 1392
rect 535 1391 536 1392
rect 540 1391 541 1395
rect 567 1395 573 1396
rect 567 1394 568 1395
rect 560 1392 568 1394
rect 535 1390 541 1391
rect 550 1390 556 1391
rect 550 1386 551 1390
rect 555 1386 556 1390
rect 550 1385 556 1386
rect 560 1380 562 1392
rect 567 1391 568 1392
rect 572 1391 573 1395
rect 592 1394 594 1400
rect 719 1399 720 1403
rect 724 1402 725 1403
rect 758 1403 759 1407
rect 763 1403 764 1407
rect 894 1406 895 1410
rect 899 1406 900 1410
rect 1059 1409 1060 1412
rect 1064 1412 1098 1413
rect 1064 1409 1065 1412
rect 1059 1408 1065 1409
rect 1096 1410 1098 1412
rect 1147 1411 1153 1412
rect 1147 1410 1148 1411
rect 1096 1408 1148 1410
rect 894 1405 900 1406
rect 1070 1407 1076 1408
rect 758 1402 764 1403
rect 1070 1403 1071 1407
rect 1075 1406 1076 1407
rect 1087 1407 1093 1408
rect 1087 1406 1088 1407
rect 1075 1404 1088 1406
rect 1075 1403 1076 1404
rect 1070 1402 1076 1403
rect 1087 1403 1088 1404
rect 1092 1403 1093 1407
rect 1147 1407 1148 1408
rect 1152 1410 1153 1411
rect 1230 1411 1236 1412
rect 1152 1408 1161 1410
rect 1152 1407 1153 1408
rect 1147 1406 1153 1407
rect 1087 1402 1093 1403
rect 724 1400 882 1402
rect 724 1399 725 1400
rect 719 1398 725 1399
rect 751 1396 757 1397
rect 599 1395 605 1396
rect 599 1394 600 1395
rect 592 1392 600 1394
rect 599 1391 600 1392
rect 604 1391 605 1395
rect 631 1395 637 1396
rect 631 1394 632 1395
rect 624 1392 632 1394
rect 567 1390 573 1391
rect 582 1390 588 1391
rect 599 1390 605 1391
rect 614 1390 620 1391
rect 582 1386 583 1390
rect 587 1386 588 1390
rect 582 1385 588 1386
rect 614 1386 615 1390
rect 619 1386 620 1390
rect 614 1385 620 1386
rect 567 1380 573 1381
rect 624 1380 626 1392
rect 631 1391 632 1392
rect 636 1391 637 1395
rect 663 1395 669 1396
rect 663 1394 664 1395
rect 656 1392 664 1394
rect 631 1390 637 1391
rect 646 1390 652 1391
rect 646 1386 647 1390
rect 651 1386 652 1390
rect 646 1385 652 1386
rect 656 1380 658 1392
rect 663 1391 664 1392
rect 668 1391 669 1395
rect 694 1395 701 1396
rect 694 1391 695 1395
rect 700 1391 701 1395
rect 663 1390 669 1391
rect 678 1390 684 1391
rect 694 1390 701 1391
rect 718 1393 724 1394
rect 678 1386 679 1390
rect 683 1386 684 1390
rect 718 1389 719 1393
rect 723 1389 724 1393
rect 751 1392 752 1396
rect 756 1394 757 1396
rect 762 1395 768 1396
rect 762 1394 763 1395
rect 756 1392 763 1394
rect 751 1391 757 1392
rect 762 1391 763 1392
rect 767 1391 768 1395
rect 762 1390 768 1391
rect 806 1395 812 1396
rect 806 1391 807 1395
rect 811 1391 812 1395
rect 806 1390 812 1391
rect 718 1388 724 1389
rect 678 1385 684 1386
rect 786 1387 797 1388
rect 786 1383 787 1387
rect 791 1383 792 1387
rect 796 1383 797 1387
rect 786 1382 797 1383
rect 863 1387 872 1388
rect 863 1383 864 1387
rect 871 1383 872 1387
rect 880 1386 882 1400
rect 1062 1400 1068 1401
rect 1062 1396 1063 1400
rect 1067 1396 1068 1400
rect 1150 1400 1156 1401
rect 1150 1396 1151 1400
rect 1155 1396 1156 1400
rect 1159 1398 1161 1408
rect 1175 1407 1181 1408
rect 1175 1403 1176 1407
rect 1180 1406 1181 1407
rect 1214 1407 1220 1408
rect 1214 1406 1215 1407
rect 1180 1404 1215 1406
rect 1180 1403 1181 1404
rect 1175 1402 1181 1403
rect 1214 1403 1215 1404
rect 1219 1403 1220 1407
rect 1230 1407 1231 1411
rect 1235 1410 1236 1411
rect 1243 1411 1249 1412
rect 1243 1410 1244 1411
rect 1235 1408 1244 1410
rect 1235 1407 1236 1408
rect 1230 1406 1236 1407
rect 1243 1407 1244 1408
rect 1248 1407 1249 1411
rect 1272 1410 1274 1420
rect 1470 1419 1471 1420
rect 1475 1419 1476 1423
rect 1470 1418 1476 1419
rect 1383 1415 1389 1416
rect 1383 1414 1384 1415
rect 1243 1406 1249 1407
rect 1267 1409 1274 1410
rect 1267 1405 1268 1409
rect 1272 1408 1274 1409
rect 1280 1412 1384 1414
rect 1272 1405 1273 1408
rect 1267 1404 1273 1405
rect 1214 1402 1220 1403
rect 1190 1399 1196 1400
rect 1190 1398 1191 1399
rect 1159 1396 1191 1398
rect 998 1395 1004 1396
rect 998 1394 999 1395
rect 948 1392 999 1394
rect 948 1388 950 1392
rect 998 1391 999 1392
rect 1003 1391 1004 1395
rect 1039 1395 1045 1396
rect 1039 1391 1040 1395
rect 1044 1394 1045 1395
rect 1054 1395 1060 1396
rect 1062 1395 1068 1396
rect 1127 1395 1136 1396
rect 1150 1395 1156 1396
rect 1190 1395 1191 1396
rect 1195 1395 1196 1399
rect 1280 1398 1282 1412
rect 1383 1411 1384 1412
rect 1388 1411 1389 1415
rect 1383 1410 1389 1411
rect 1458 1415 1464 1416
rect 1458 1411 1459 1415
rect 1463 1414 1464 1415
rect 1463 1413 1522 1414
rect 1464 1412 1522 1413
rect 1458 1410 1460 1411
rect 1459 1409 1460 1410
rect 1464 1409 1465 1412
rect 1459 1408 1465 1409
rect 1520 1410 1522 1412
rect 1747 1411 1753 1412
rect 1747 1410 1748 1411
rect 1520 1408 1748 1410
rect 1367 1407 1373 1408
rect 1367 1406 1368 1407
rect 1054 1394 1055 1395
rect 1044 1392 1055 1394
rect 1044 1391 1045 1392
rect 998 1390 1004 1391
rect 1022 1390 1028 1391
rect 1039 1390 1045 1391
rect 1054 1391 1055 1392
rect 1059 1391 1060 1395
rect 1054 1390 1060 1391
rect 1110 1391 1116 1392
rect 940 1386 950 1388
rect 966 1387 972 1388
rect 880 1384 942 1386
rect 863 1382 872 1383
rect 946 1383 952 1384
rect 151 1379 157 1380
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 151 1375 152 1379
rect 156 1378 157 1379
rect 164 1378 178 1380
rect 183 1379 189 1380
rect 156 1376 166 1378
rect 156 1375 157 1376
rect 151 1374 157 1375
rect 183 1375 184 1379
rect 188 1378 189 1379
rect 196 1378 210 1380
rect 215 1379 221 1380
rect 188 1376 198 1378
rect 188 1375 189 1376
rect 183 1374 189 1375
rect 215 1375 216 1379
rect 220 1378 221 1379
rect 228 1378 242 1380
rect 247 1379 253 1380
rect 220 1376 230 1378
rect 220 1375 221 1376
rect 215 1374 221 1375
rect 247 1375 248 1379
rect 252 1378 253 1379
rect 260 1378 274 1380
rect 279 1379 285 1380
rect 252 1376 262 1378
rect 252 1375 253 1376
rect 247 1374 253 1375
rect 279 1375 280 1379
rect 284 1378 285 1379
rect 292 1378 306 1380
rect 311 1379 317 1380
rect 284 1376 294 1378
rect 284 1375 285 1376
rect 279 1374 285 1375
rect 311 1375 312 1379
rect 316 1378 317 1379
rect 324 1378 338 1380
rect 343 1379 352 1380
rect 316 1376 326 1378
rect 316 1375 317 1376
rect 311 1374 317 1375
rect 343 1375 344 1379
rect 351 1375 352 1379
rect 343 1374 352 1375
rect 375 1379 381 1380
rect 375 1375 376 1379
rect 380 1378 381 1379
rect 388 1378 402 1380
rect 407 1379 413 1380
rect 380 1376 390 1378
rect 380 1375 381 1376
rect 375 1374 381 1375
rect 407 1375 408 1379
rect 412 1378 413 1379
rect 420 1378 434 1380
rect 439 1379 445 1380
rect 412 1376 422 1378
rect 412 1375 413 1376
rect 407 1374 413 1375
rect 439 1375 440 1379
rect 444 1378 445 1379
rect 452 1378 466 1380
rect 470 1379 477 1380
rect 444 1376 454 1378
rect 444 1375 445 1376
rect 439 1374 445 1375
rect 470 1375 471 1379
rect 476 1375 477 1379
rect 470 1374 477 1375
rect 503 1379 509 1380
rect 503 1375 504 1379
rect 508 1378 509 1379
rect 516 1378 530 1380
rect 535 1379 541 1380
rect 508 1376 518 1378
rect 508 1375 509 1376
rect 503 1374 509 1375
rect 535 1375 536 1379
rect 540 1378 541 1379
rect 548 1378 562 1380
rect 566 1379 568 1380
rect 540 1376 550 1378
rect 540 1375 541 1376
rect 535 1374 541 1375
rect 566 1375 567 1379
rect 572 1376 573 1380
rect 571 1375 573 1376
rect 599 1379 605 1380
rect 599 1375 600 1379
rect 604 1378 605 1379
rect 612 1378 626 1380
rect 631 1379 637 1380
rect 604 1376 614 1378
rect 604 1375 605 1376
rect 566 1374 572 1375
rect 599 1374 605 1375
rect 631 1375 632 1379
rect 636 1378 637 1379
rect 644 1378 658 1380
rect 662 1379 669 1380
rect 636 1376 646 1378
rect 636 1375 637 1376
rect 631 1374 637 1375
rect 662 1375 663 1379
rect 668 1375 669 1379
rect 662 1374 669 1375
rect 695 1379 701 1380
rect 695 1375 696 1379
rect 700 1378 701 1379
rect 703 1379 709 1380
rect 703 1378 704 1379
rect 700 1376 704 1378
rect 700 1375 701 1376
rect 695 1374 701 1375
rect 703 1375 704 1376
rect 708 1375 709 1379
rect 846 1379 852 1380
rect 846 1378 847 1379
rect 828 1376 847 1378
rect 703 1374 709 1375
rect 823 1375 830 1376
rect 110 1370 116 1371
rect 134 1373 140 1374
rect 134 1369 135 1373
rect 139 1369 140 1373
rect 134 1368 140 1369
rect 166 1373 172 1374
rect 166 1369 167 1373
rect 171 1369 172 1373
rect 166 1368 172 1369
rect 198 1373 204 1374
rect 198 1369 199 1373
rect 203 1369 204 1373
rect 198 1368 204 1369
rect 230 1373 236 1374
rect 230 1369 231 1373
rect 235 1369 236 1373
rect 230 1368 236 1369
rect 262 1373 268 1374
rect 262 1369 263 1373
rect 267 1369 268 1373
rect 262 1368 268 1369
rect 294 1373 300 1374
rect 294 1369 295 1373
rect 299 1369 300 1373
rect 294 1368 300 1369
rect 326 1373 332 1374
rect 326 1369 327 1373
rect 331 1369 332 1373
rect 326 1368 332 1369
rect 358 1373 364 1374
rect 358 1369 359 1373
rect 363 1369 364 1373
rect 358 1368 364 1369
rect 390 1373 396 1374
rect 390 1369 391 1373
rect 395 1369 396 1373
rect 390 1368 396 1369
rect 422 1373 428 1374
rect 422 1369 423 1373
rect 427 1369 428 1373
rect 422 1368 428 1369
rect 454 1373 460 1374
rect 454 1369 455 1373
rect 459 1369 460 1373
rect 454 1368 460 1369
rect 486 1373 492 1374
rect 486 1369 487 1373
rect 491 1369 492 1373
rect 486 1368 492 1369
rect 518 1373 524 1374
rect 518 1369 519 1373
rect 523 1369 524 1373
rect 518 1368 524 1369
rect 550 1373 556 1374
rect 550 1369 551 1373
rect 555 1369 556 1373
rect 550 1368 556 1369
rect 582 1373 588 1374
rect 582 1369 583 1373
rect 587 1369 588 1373
rect 582 1368 588 1369
rect 614 1373 620 1374
rect 614 1369 615 1373
rect 619 1369 620 1373
rect 614 1368 620 1369
rect 646 1373 652 1374
rect 646 1369 647 1373
rect 651 1369 652 1373
rect 646 1368 652 1369
rect 678 1373 684 1374
rect 678 1369 679 1373
rect 683 1369 684 1373
rect 806 1372 812 1373
rect 678 1368 684 1369
rect 766 1368 772 1369
rect 378 1367 384 1368
rect 378 1363 379 1367
rect 383 1366 384 1367
rect 566 1367 572 1368
rect 566 1366 567 1367
rect 383 1364 567 1366
rect 383 1363 384 1364
rect 378 1362 384 1363
rect 566 1363 567 1364
rect 571 1363 572 1367
rect 566 1362 572 1363
rect 734 1366 740 1367
rect 734 1362 735 1366
rect 739 1362 740 1366
rect 766 1364 767 1368
rect 771 1364 772 1368
rect 806 1368 807 1372
rect 811 1368 812 1372
rect 823 1371 824 1375
rect 828 1372 830 1375
rect 846 1375 847 1376
rect 851 1375 852 1379
rect 946 1379 947 1383
rect 951 1379 952 1383
rect 966 1383 967 1387
rect 971 1386 972 1387
rect 999 1387 1005 1388
rect 999 1386 1000 1387
rect 971 1384 1000 1386
rect 971 1383 972 1384
rect 966 1382 972 1383
rect 999 1383 1000 1384
rect 1004 1383 1005 1387
rect 1022 1386 1023 1390
rect 1027 1386 1028 1390
rect 1022 1385 1028 1386
rect 1087 1387 1093 1388
rect 999 1382 1005 1383
rect 1070 1383 1076 1384
rect 1070 1382 1071 1383
rect 1060 1380 1071 1382
rect 946 1378 952 1379
rect 1039 1379 1045 1380
rect 846 1374 852 1375
rect 1039 1375 1040 1379
rect 1044 1378 1045 1379
rect 1060 1378 1062 1380
rect 1070 1379 1071 1380
rect 1075 1379 1076 1383
rect 1087 1383 1088 1387
rect 1092 1386 1093 1387
rect 1102 1387 1108 1388
rect 1102 1386 1103 1387
rect 1092 1384 1103 1386
rect 1092 1383 1093 1384
rect 1087 1382 1093 1383
rect 1102 1383 1103 1384
rect 1107 1383 1108 1387
rect 1110 1387 1111 1391
rect 1115 1387 1116 1391
rect 1127 1391 1128 1395
rect 1135 1391 1136 1395
rect 1190 1394 1196 1395
rect 1215 1397 1282 1398
rect 1215 1393 1216 1397
rect 1220 1396 1282 1397
rect 1284 1404 1368 1406
rect 1220 1393 1221 1396
rect 1284 1394 1286 1404
rect 1367 1403 1368 1404
rect 1372 1403 1373 1407
rect 1367 1402 1373 1403
rect 1470 1407 1476 1408
rect 1470 1403 1471 1407
rect 1475 1406 1476 1407
rect 1483 1407 1489 1408
rect 1483 1406 1484 1407
rect 1475 1404 1484 1406
rect 1475 1403 1476 1404
rect 1470 1402 1476 1403
rect 1483 1403 1484 1404
rect 1488 1403 1489 1407
rect 1747 1407 1748 1408
rect 1752 1407 1753 1411
rect 1747 1406 1753 1407
rect 1483 1402 1489 1403
rect 1406 1399 1412 1400
rect 1406 1395 1407 1399
rect 1411 1398 1412 1399
rect 1574 1399 1580 1400
rect 1411 1397 1437 1398
rect 1411 1396 1432 1397
rect 1411 1395 1412 1396
rect 1406 1394 1412 1395
rect 1215 1392 1221 1393
rect 1262 1393 1268 1394
rect 1127 1390 1136 1391
rect 1198 1390 1204 1391
rect 1110 1386 1116 1387
rect 1166 1387 1172 1388
rect 1102 1382 1108 1383
rect 1166 1383 1167 1387
rect 1171 1386 1172 1387
rect 1175 1387 1181 1388
rect 1175 1386 1176 1387
rect 1171 1384 1176 1386
rect 1171 1383 1172 1384
rect 1166 1382 1172 1383
rect 1175 1383 1176 1384
rect 1180 1383 1181 1387
rect 1198 1386 1199 1390
rect 1203 1386 1204 1390
rect 1262 1389 1263 1393
rect 1267 1389 1268 1393
rect 1262 1388 1268 1389
rect 1283 1393 1289 1394
rect 1283 1389 1284 1393
rect 1288 1389 1289 1393
rect 1431 1393 1432 1396
rect 1436 1393 1437 1397
rect 1550 1395 1557 1396
rect 1431 1392 1437 1393
rect 1478 1393 1484 1394
rect 1283 1388 1289 1389
rect 1318 1391 1324 1392
rect 1318 1387 1319 1391
rect 1323 1387 1324 1391
rect 1318 1386 1324 1387
rect 1414 1390 1420 1391
rect 1414 1386 1415 1390
rect 1419 1386 1420 1390
rect 1478 1389 1479 1393
rect 1483 1389 1484 1393
rect 1478 1388 1484 1389
rect 1486 1391 1492 1392
rect 1486 1387 1487 1391
rect 1491 1390 1492 1391
rect 1499 1391 1505 1392
rect 1550 1391 1551 1395
rect 1556 1391 1557 1395
rect 1574 1395 1575 1399
rect 1579 1398 1580 1399
rect 1607 1399 1613 1400
rect 1579 1396 1594 1398
rect 1579 1395 1580 1396
rect 1574 1394 1580 1395
rect 1592 1394 1594 1396
rect 1599 1395 1605 1396
rect 1599 1394 1600 1395
rect 1592 1392 1600 1394
rect 1599 1391 1600 1392
rect 1604 1391 1605 1395
rect 1607 1395 1608 1399
rect 1612 1398 1613 1399
rect 1612 1396 1634 1398
rect 1612 1395 1613 1396
rect 1607 1394 1613 1395
rect 1632 1394 1634 1396
rect 1639 1395 1645 1396
rect 1639 1394 1640 1395
rect 1632 1392 1640 1394
rect 1639 1391 1640 1392
rect 1644 1391 1645 1395
rect 1671 1395 1677 1396
rect 1671 1394 1672 1395
rect 1664 1392 1672 1394
rect 1499 1390 1500 1391
rect 1491 1388 1500 1390
rect 1491 1387 1492 1388
rect 1486 1386 1492 1387
rect 1499 1387 1500 1388
rect 1504 1387 1505 1391
rect 1499 1386 1505 1387
rect 1534 1390 1540 1391
rect 1550 1390 1557 1391
rect 1582 1390 1588 1391
rect 1599 1390 1605 1391
rect 1622 1390 1628 1391
rect 1639 1390 1645 1391
rect 1654 1390 1660 1391
rect 1534 1386 1535 1390
rect 1539 1386 1540 1390
rect 1198 1385 1204 1386
rect 1414 1385 1420 1386
rect 1534 1385 1540 1386
rect 1582 1386 1583 1390
rect 1587 1386 1588 1390
rect 1582 1385 1588 1386
rect 1622 1386 1623 1390
rect 1627 1386 1628 1390
rect 1622 1385 1628 1386
rect 1654 1386 1655 1390
rect 1659 1386 1660 1390
rect 1654 1385 1660 1386
rect 1175 1382 1181 1383
rect 1298 1383 1304 1384
rect 1070 1378 1076 1379
rect 1122 1379 1133 1380
rect 1044 1376 1062 1378
rect 1044 1375 1045 1376
rect 1039 1374 1045 1375
rect 1122 1375 1123 1379
rect 1127 1375 1128 1379
rect 1132 1375 1133 1379
rect 1122 1374 1133 1375
rect 1214 1379 1221 1380
rect 1214 1375 1215 1379
rect 1220 1375 1221 1379
rect 1298 1379 1299 1383
rect 1303 1382 1304 1383
rect 1303 1380 1361 1382
rect 1664 1380 1666 1392
rect 1671 1391 1672 1392
rect 1676 1391 1677 1395
rect 1671 1390 1677 1391
rect 1694 1392 1700 1393
rect 1694 1388 1695 1392
rect 1699 1388 1700 1392
rect 1694 1387 1700 1388
rect 1303 1379 1304 1380
rect 1298 1378 1304 1379
rect 1431 1379 1437 1380
rect 1214 1374 1221 1375
rect 1431 1375 1432 1379
rect 1436 1378 1437 1379
rect 1446 1379 1452 1380
rect 1446 1378 1447 1379
rect 1436 1376 1447 1378
rect 1436 1375 1437 1376
rect 1431 1374 1437 1375
rect 1446 1375 1447 1376
rect 1451 1375 1452 1379
rect 1446 1374 1452 1375
rect 1546 1379 1557 1380
rect 1546 1375 1547 1379
rect 1551 1375 1552 1379
rect 1556 1375 1557 1379
rect 1546 1374 1557 1375
rect 1599 1379 1605 1380
rect 1599 1375 1600 1379
rect 1604 1378 1605 1379
rect 1607 1379 1613 1380
rect 1607 1378 1608 1379
rect 1604 1376 1608 1378
rect 1604 1375 1605 1376
rect 1599 1374 1605 1375
rect 1607 1375 1608 1376
rect 1612 1375 1613 1379
rect 1607 1374 1613 1375
rect 1639 1379 1645 1380
rect 1639 1375 1640 1379
rect 1644 1378 1645 1379
rect 1652 1378 1666 1380
rect 1671 1379 1677 1380
rect 1644 1376 1654 1378
rect 1644 1375 1645 1376
rect 1639 1374 1645 1375
rect 1671 1375 1672 1379
rect 1676 1375 1677 1379
rect 1671 1374 1677 1375
rect 1694 1375 1700 1376
rect 1022 1373 1028 1374
rect 1110 1373 1116 1374
rect 1198 1373 1204 1374
rect 1414 1373 1420 1374
rect 1534 1373 1540 1374
rect 886 1372 892 1373
rect 828 1371 829 1372
rect 823 1370 829 1371
rect 806 1367 812 1368
rect 838 1368 844 1369
rect 766 1363 772 1364
rect 838 1364 839 1368
rect 843 1364 844 1368
rect 886 1368 887 1372
rect 891 1368 892 1372
rect 1022 1369 1023 1373
rect 1027 1369 1028 1373
rect 886 1367 892 1368
rect 974 1368 980 1369
rect 1022 1368 1028 1369
rect 1062 1372 1068 1373
rect 1062 1368 1063 1372
rect 1067 1368 1068 1372
rect 1110 1369 1111 1373
rect 1115 1369 1116 1373
rect 1110 1368 1116 1369
rect 1150 1372 1156 1373
rect 1150 1368 1151 1372
rect 1155 1368 1156 1372
rect 1198 1369 1199 1373
rect 1203 1369 1204 1373
rect 1198 1368 1204 1369
rect 1246 1372 1252 1373
rect 1246 1368 1247 1372
rect 1251 1368 1252 1372
rect 838 1363 844 1364
rect 974 1364 975 1368
rect 979 1364 980 1368
rect 1062 1367 1068 1368
rect 1150 1367 1156 1368
rect 1246 1367 1252 1368
rect 1318 1372 1324 1373
rect 1318 1368 1319 1372
rect 1323 1368 1324 1372
rect 1414 1369 1415 1373
rect 1419 1369 1420 1373
rect 1414 1368 1420 1369
rect 1462 1372 1468 1373
rect 1462 1368 1463 1372
rect 1467 1368 1468 1372
rect 1534 1369 1535 1373
rect 1539 1369 1540 1373
rect 1534 1368 1540 1369
rect 1582 1373 1588 1374
rect 1582 1369 1583 1373
rect 1587 1369 1588 1373
rect 1582 1368 1588 1369
rect 1622 1373 1628 1374
rect 1622 1369 1623 1373
rect 1627 1369 1628 1373
rect 1622 1368 1628 1369
rect 1654 1373 1660 1374
rect 1654 1369 1655 1373
rect 1659 1369 1660 1373
rect 1654 1368 1660 1369
rect 1318 1367 1324 1368
rect 1462 1367 1468 1368
rect 1574 1367 1580 1368
rect 974 1363 980 1364
rect 1574 1363 1575 1367
rect 1579 1366 1580 1367
rect 1672 1366 1674 1374
rect 1694 1371 1695 1375
rect 1699 1371 1700 1375
rect 1694 1370 1700 1371
rect 1579 1364 1674 1366
rect 1579 1363 1580 1364
rect 1574 1362 1580 1363
rect 734 1361 740 1362
rect 686 1359 692 1360
rect 686 1355 687 1359
rect 691 1358 692 1359
rect 711 1359 717 1360
rect 711 1358 712 1359
rect 691 1356 712 1358
rect 691 1355 692 1356
rect 686 1354 692 1355
rect 711 1355 712 1356
rect 716 1355 717 1359
rect 711 1354 717 1355
rect 814 1355 820 1356
rect 814 1351 815 1355
rect 819 1354 820 1355
rect 950 1355 956 1356
rect 950 1354 951 1355
rect 819 1352 951 1354
rect 819 1351 820 1352
rect 814 1350 820 1351
rect 950 1351 951 1352
rect 955 1354 956 1355
rect 1122 1355 1128 1356
rect 1122 1354 1123 1355
rect 955 1352 1123 1354
rect 955 1351 956 1352
rect 950 1350 956 1351
rect 1122 1351 1123 1352
rect 1127 1351 1128 1355
rect 1122 1350 1128 1351
rect 1371 1355 1377 1356
rect 1371 1351 1372 1355
rect 1376 1354 1377 1355
rect 1486 1355 1492 1356
rect 1486 1354 1487 1355
rect 1376 1352 1487 1354
rect 1376 1351 1377 1352
rect 1371 1350 1377 1351
rect 1486 1351 1487 1352
rect 1491 1351 1492 1355
rect 1486 1350 1492 1351
rect 1115 1343 1121 1344
rect 1115 1339 1116 1343
rect 1120 1342 1121 1343
rect 1166 1343 1172 1344
rect 1166 1342 1167 1343
rect 1120 1340 1167 1342
rect 1120 1339 1121 1340
rect 1115 1338 1121 1339
rect 1166 1339 1167 1340
rect 1171 1339 1172 1343
rect 1166 1338 1172 1339
rect 79 1335 85 1336
rect 79 1331 80 1335
rect 84 1334 85 1335
rect 178 1335 184 1336
rect 178 1334 179 1335
rect 84 1332 179 1334
rect 84 1331 85 1332
rect 79 1330 85 1331
rect 178 1331 179 1332
rect 183 1331 184 1335
rect 178 1330 184 1331
rect 1238 1335 1244 1336
rect 1238 1331 1239 1335
rect 1243 1334 1244 1335
rect 1267 1335 1273 1336
rect 1267 1334 1268 1335
rect 1243 1332 1268 1334
rect 1243 1331 1244 1332
rect 1238 1330 1244 1331
rect 1267 1331 1268 1332
rect 1272 1331 1273 1335
rect 1267 1330 1273 1331
rect 1355 1335 1361 1336
rect 1355 1331 1356 1335
rect 1360 1334 1361 1335
rect 1447 1335 1453 1336
rect 1447 1334 1448 1335
rect 1360 1332 1448 1334
rect 1360 1331 1361 1332
rect 1355 1330 1361 1331
rect 1447 1331 1448 1332
rect 1452 1331 1453 1335
rect 1447 1330 1453 1331
rect 982 1324 988 1325
rect 742 1320 748 1321
rect 134 1319 140 1320
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1315 135 1319
rect 139 1315 140 1319
rect 134 1314 140 1315
rect 166 1319 172 1320
rect 166 1315 167 1319
rect 171 1315 172 1319
rect 166 1314 172 1315
rect 198 1319 204 1320
rect 198 1315 199 1319
rect 203 1315 204 1319
rect 198 1314 204 1315
rect 230 1319 236 1320
rect 230 1315 231 1319
rect 235 1315 236 1319
rect 230 1314 236 1315
rect 262 1319 268 1320
rect 262 1315 263 1319
rect 267 1315 268 1319
rect 262 1314 268 1315
rect 294 1319 300 1320
rect 294 1315 295 1319
rect 299 1315 300 1319
rect 294 1314 300 1315
rect 326 1319 332 1320
rect 326 1315 327 1319
rect 331 1315 332 1319
rect 326 1314 332 1315
rect 358 1319 364 1320
rect 358 1315 359 1319
rect 363 1315 364 1319
rect 358 1314 364 1315
rect 390 1319 396 1320
rect 390 1315 391 1319
rect 395 1315 396 1319
rect 390 1314 396 1315
rect 422 1319 428 1320
rect 422 1315 423 1319
rect 427 1315 428 1319
rect 422 1314 428 1315
rect 454 1319 460 1320
rect 454 1315 455 1319
rect 459 1315 460 1319
rect 454 1314 460 1315
rect 486 1319 492 1320
rect 486 1315 487 1319
rect 491 1315 492 1319
rect 486 1314 492 1315
rect 518 1319 524 1320
rect 518 1315 519 1319
rect 523 1315 524 1319
rect 518 1314 524 1315
rect 550 1319 556 1320
rect 550 1315 551 1319
rect 555 1315 556 1319
rect 550 1314 556 1315
rect 582 1319 588 1320
rect 582 1315 583 1319
rect 587 1315 588 1319
rect 582 1314 588 1315
rect 614 1319 620 1320
rect 614 1315 615 1319
rect 619 1315 620 1319
rect 614 1314 620 1315
rect 646 1319 652 1320
rect 646 1315 647 1319
rect 651 1315 652 1319
rect 646 1314 652 1315
rect 678 1319 684 1320
rect 678 1315 679 1319
rect 683 1315 684 1319
rect 678 1314 684 1315
rect 710 1319 716 1320
rect 710 1315 711 1319
rect 715 1315 716 1319
rect 742 1316 743 1320
rect 747 1316 748 1320
rect 742 1315 748 1316
rect 822 1320 828 1321
rect 822 1316 823 1320
rect 827 1316 828 1320
rect 822 1315 828 1316
rect 902 1320 908 1321
rect 902 1316 903 1320
rect 907 1316 908 1320
rect 982 1320 983 1324
rect 987 1320 988 1324
rect 982 1319 988 1320
rect 1022 1320 1028 1321
rect 902 1315 908 1316
rect 1022 1316 1023 1320
rect 1027 1316 1028 1320
rect 1022 1315 1028 1316
rect 1062 1320 1068 1321
rect 1062 1316 1063 1320
rect 1067 1316 1068 1320
rect 1062 1315 1068 1316
rect 1158 1320 1164 1321
rect 1158 1316 1159 1320
rect 1163 1316 1164 1320
rect 1158 1315 1164 1316
rect 1214 1320 1220 1321
rect 1214 1316 1215 1320
rect 1219 1316 1220 1320
rect 1214 1315 1220 1316
rect 1302 1320 1308 1321
rect 1454 1320 1460 1321
rect 1302 1316 1303 1320
rect 1307 1316 1308 1320
rect 1302 1315 1308 1316
rect 1390 1319 1396 1320
rect 1390 1315 1391 1319
rect 1395 1315 1396 1319
rect 710 1314 716 1315
rect 1390 1314 1396 1315
rect 1422 1319 1428 1320
rect 1422 1315 1423 1319
rect 1427 1315 1428 1319
rect 1454 1316 1455 1320
rect 1459 1316 1460 1320
rect 1454 1315 1460 1316
rect 1494 1319 1500 1320
rect 1494 1315 1495 1319
rect 1499 1315 1500 1319
rect 1422 1314 1428 1315
rect 1494 1314 1500 1315
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1558 1319 1564 1320
rect 1558 1315 1559 1319
rect 1563 1315 1564 1319
rect 1558 1314 1564 1315
rect 1590 1319 1596 1320
rect 1590 1315 1591 1319
rect 1595 1315 1596 1319
rect 1590 1314 1596 1315
rect 1622 1319 1628 1320
rect 1622 1315 1623 1319
rect 1627 1315 1628 1319
rect 1622 1314 1628 1315
rect 1654 1319 1660 1320
rect 1654 1315 1655 1319
rect 1659 1315 1660 1319
rect 1654 1314 1660 1315
rect 1694 1317 1700 1318
rect 110 1312 116 1313
rect 1694 1313 1695 1317
rect 1699 1313 1700 1317
rect 1694 1312 1700 1313
rect 150 1311 157 1312
rect 150 1307 151 1311
rect 156 1307 157 1311
rect 183 1311 189 1312
rect 183 1310 184 1311
rect 150 1306 157 1307
rect 176 1308 184 1310
rect 134 1302 140 1303
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 134 1298 135 1302
rect 139 1298 140 1302
rect 134 1297 140 1298
rect 166 1302 172 1303
rect 166 1298 167 1302
rect 171 1298 172 1302
rect 166 1297 172 1298
rect 110 1295 116 1296
rect 151 1295 157 1296
rect 151 1291 152 1295
rect 156 1294 157 1295
rect 176 1294 178 1308
rect 183 1307 184 1308
rect 188 1307 189 1311
rect 215 1311 221 1312
rect 215 1310 216 1311
rect 183 1306 189 1307
rect 208 1308 216 1310
rect 198 1302 204 1303
rect 198 1298 199 1302
rect 203 1298 204 1302
rect 198 1297 204 1298
rect 156 1292 178 1294
rect 183 1295 189 1296
rect 156 1291 157 1292
rect 151 1290 157 1291
rect 183 1291 184 1295
rect 188 1294 189 1295
rect 208 1294 210 1308
rect 215 1307 216 1308
rect 220 1307 221 1311
rect 247 1311 253 1312
rect 247 1310 248 1311
rect 215 1306 221 1307
rect 240 1308 248 1310
rect 230 1302 236 1303
rect 230 1298 231 1302
rect 235 1298 236 1302
rect 230 1297 236 1298
rect 188 1292 210 1294
rect 215 1295 221 1296
rect 188 1291 189 1292
rect 183 1290 189 1291
rect 215 1291 216 1295
rect 220 1294 221 1295
rect 240 1294 242 1308
rect 247 1307 248 1308
rect 252 1307 253 1311
rect 279 1311 285 1312
rect 279 1310 280 1311
rect 247 1306 253 1307
rect 272 1308 280 1310
rect 262 1302 268 1303
rect 262 1298 263 1302
rect 267 1298 268 1302
rect 262 1297 268 1298
rect 220 1292 242 1294
rect 247 1295 253 1296
rect 220 1291 221 1292
rect 215 1290 221 1291
rect 247 1291 248 1295
rect 252 1294 253 1295
rect 272 1294 274 1308
rect 279 1307 280 1308
rect 284 1307 285 1311
rect 311 1311 317 1312
rect 311 1310 312 1311
rect 279 1306 285 1307
rect 304 1308 312 1310
rect 294 1302 300 1303
rect 294 1298 295 1302
rect 299 1298 300 1302
rect 294 1297 300 1298
rect 252 1292 274 1294
rect 279 1295 285 1296
rect 252 1291 253 1292
rect 247 1290 253 1291
rect 279 1291 280 1295
rect 284 1294 285 1295
rect 304 1294 306 1308
rect 311 1307 312 1308
rect 316 1307 317 1311
rect 343 1311 349 1312
rect 343 1310 344 1311
rect 311 1306 317 1307
rect 336 1308 344 1310
rect 326 1302 332 1303
rect 326 1298 327 1302
rect 331 1298 332 1302
rect 326 1297 332 1298
rect 284 1292 306 1294
rect 311 1295 317 1296
rect 284 1291 285 1292
rect 279 1290 285 1291
rect 311 1291 312 1295
rect 316 1294 317 1295
rect 336 1294 338 1308
rect 343 1307 344 1308
rect 348 1307 349 1311
rect 343 1306 349 1307
rect 375 1311 381 1312
rect 375 1307 376 1311
rect 380 1310 381 1311
rect 407 1311 413 1312
rect 380 1308 402 1310
rect 380 1307 381 1308
rect 375 1306 381 1307
rect 346 1303 352 1304
rect 346 1299 347 1303
rect 351 1302 352 1303
rect 358 1302 364 1303
rect 351 1299 354 1302
rect 346 1298 354 1299
rect 316 1292 338 1294
rect 343 1295 349 1296
rect 316 1291 317 1292
rect 311 1290 317 1291
rect 343 1291 344 1295
rect 348 1294 349 1295
rect 352 1294 354 1298
rect 358 1298 359 1302
rect 363 1298 364 1302
rect 358 1297 364 1298
rect 390 1302 396 1303
rect 390 1298 391 1302
rect 395 1298 396 1302
rect 390 1297 396 1298
rect 375 1295 381 1296
rect 375 1294 376 1295
rect 348 1291 350 1294
rect 352 1292 376 1294
rect 343 1290 350 1291
rect 375 1291 376 1292
rect 380 1291 381 1295
rect 400 1294 402 1308
rect 407 1307 408 1311
rect 412 1310 413 1311
rect 439 1311 445 1312
rect 412 1308 434 1310
rect 412 1307 413 1308
rect 407 1306 413 1307
rect 422 1302 428 1303
rect 422 1298 423 1302
rect 427 1298 428 1302
rect 422 1297 428 1298
rect 407 1295 413 1296
rect 407 1294 408 1295
rect 400 1292 408 1294
rect 375 1290 381 1291
rect 407 1291 408 1292
rect 412 1291 413 1295
rect 432 1294 434 1308
rect 439 1307 440 1311
rect 444 1310 445 1311
rect 471 1311 477 1312
rect 444 1308 466 1310
rect 444 1307 445 1308
rect 439 1306 445 1307
rect 454 1302 460 1303
rect 454 1298 455 1302
rect 459 1298 460 1302
rect 454 1297 460 1298
rect 439 1295 445 1296
rect 439 1294 440 1295
rect 432 1292 440 1294
rect 407 1290 413 1291
rect 439 1291 440 1292
rect 444 1291 445 1295
rect 464 1294 466 1308
rect 471 1307 472 1311
rect 476 1310 477 1311
rect 503 1311 509 1312
rect 476 1308 498 1310
rect 476 1307 477 1308
rect 471 1306 477 1307
rect 486 1302 492 1303
rect 486 1298 487 1302
rect 491 1298 492 1302
rect 486 1297 492 1298
rect 471 1295 477 1296
rect 471 1294 472 1295
rect 464 1292 472 1294
rect 439 1290 445 1291
rect 471 1291 472 1292
rect 476 1291 477 1295
rect 496 1294 498 1308
rect 503 1307 504 1311
rect 508 1310 509 1311
rect 535 1311 541 1312
rect 508 1308 530 1310
rect 508 1307 509 1308
rect 503 1306 509 1307
rect 518 1302 524 1303
rect 518 1298 519 1302
rect 523 1298 524 1302
rect 518 1297 524 1298
rect 503 1295 509 1296
rect 503 1294 504 1295
rect 496 1292 504 1294
rect 471 1290 477 1291
rect 503 1291 504 1292
rect 508 1291 509 1295
rect 528 1294 530 1308
rect 535 1307 536 1311
rect 540 1310 541 1311
rect 567 1311 573 1312
rect 540 1308 562 1310
rect 540 1307 541 1308
rect 535 1306 541 1307
rect 550 1302 556 1303
rect 550 1298 551 1302
rect 555 1298 556 1302
rect 550 1297 556 1298
rect 535 1295 541 1296
rect 535 1294 536 1295
rect 528 1292 536 1294
rect 503 1290 509 1291
rect 535 1291 536 1292
rect 540 1291 541 1295
rect 560 1294 562 1308
rect 567 1307 568 1311
rect 572 1310 573 1311
rect 599 1311 605 1312
rect 572 1308 594 1310
rect 572 1307 573 1308
rect 567 1306 573 1307
rect 582 1302 588 1303
rect 582 1298 583 1302
rect 587 1298 588 1302
rect 582 1297 588 1298
rect 567 1295 573 1296
rect 567 1294 568 1295
rect 560 1292 568 1294
rect 535 1290 541 1291
rect 567 1291 568 1292
rect 572 1291 573 1295
rect 592 1294 594 1308
rect 599 1307 600 1311
rect 604 1310 605 1311
rect 607 1311 613 1312
rect 607 1310 608 1311
rect 604 1308 608 1310
rect 604 1307 605 1308
rect 599 1306 605 1307
rect 607 1307 608 1308
rect 612 1307 613 1311
rect 607 1306 613 1307
rect 626 1311 637 1312
rect 626 1307 627 1311
rect 631 1307 632 1311
rect 636 1307 637 1311
rect 663 1311 669 1312
rect 663 1310 664 1311
rect 626 1306 637 1307
rect 656 1308 664 1310
rect 614 1302 620 1303
rect 614 1298 615 1302
rect 619 1298 620 1302
rect 614 1297 620 1298
rect 646 1302 652 1303
rect 646 1298 647 1302
rect 651 1298 652 1302
rect 646 1297 652 1298
rect 599 1295 605 1296
rect 599 1294 600 1295
rect 592 1292 600 1294
rect 567 1290 573 1291
rect 599 1291 600 1292
rect 604 1291 605 1295
rect 599 1290 605 1291
rect 631 1295 637 1296
rect 631 1291 632 1295
rect 636 1294 637 1295
rect 656 1294 658 1308
rect 663 1307 664 1308
rect 668 1307 669 1311
rect 663 1306 669 1307
rect 694 1311 701 1312
rect 694 1307 695 1311
rect 700 1307 701 1311
rect 727 1311 733 1312
rect 727 1310 728 1311
rect 694 1306 701 1307
rect 720 1308 728 1310
rect 678 1302 684 1303
rect 678 1298 679 1302
rect 683 1298 684 1302
rect 678 1297 684 1298
rect 710 1302 716 1303
rect 710 1298 711 1302
rect 715 1298 716 1302
rect 710 1297 716 1298
rect 636 1292 658 1294
rect 662 1295 669 1296
rect 636 1291 637 1292
rect 631 1290 637 1291
rect 662 1291 663 1295
rect 668 1291 669 1295
rect 662 1290 669 1291
rect 695 1295 701 1296
rect 695 1291 696 1295
rect 700 1294 701 1295
rect 720 1294 722 1308
rect 727 1307 728 1308
rect 732 1307 733 1311
rect 970 1311 976 1312
rect 970 1310 971 1311
rect 752 1308 761 1310
rect 832 1308 841 1310
rect 965 1308 971 1310
rect 727 1306 733 1307
rect 750 1307 756 1308
rect 750 1303 751 1307
rect 755 1303 756 1307
rect 750 1302 756 1303
rect 830 1307 836 1308
rect 830 1303 831 1307
rect 835 1303 836 1307
rect 970 1307 971 1308
rect 975 1307 976 1311
rect 970 1306 976 1307
rect 1130 1311 1136 1312
rect 1130 1307 1131 1311
rect 1135 1307 1136 1311
rect 1130 1306 1136 1307
rect 1286 1311 1292 1312
rect 1286 1307 1287 1311
rect 1291 1307 1292 1311
rect 1286 1306 1292 1307
rect 1407 1311 1416 1312
rect 1407 1307 1408 1311
rect 1415 1307 1416 1311
rect 1407 1306 1416 1307
rect 1434 1311 1445 1312
rect 1434 1307 1435 1311
rect 1439 1307 1440 1311
rect 1444 1307 1445 1311
rect 1434 1306 1445 1307
rect 1482 1311 1488 1312
rect 1482 1307 1483 1311
rect 1487 1310 1488 1311
rect 1511 1311 1517 1312
rect 1511 1310 1512 1311
rect 1487 1308 1512 1310
rect 1487 1307 1488 1308
rect 1482 1306 1488 1307
rect 1511 1307 1512 1308
rect 1516 1307 1517 1311
rect 1511 1306 1517 1307
rect 1538 1311 1549 1312
rect 1538 1307 1539 1311
rect 1543 1307 1544 1311
rect 1548 1307 1549 1311
rect 1538 1306 1549 1307
rect 1575 1311 1581 1312
rect 1575 1307 1576 1311
rect 1580 1310 1581 1311
rect 1607 1311 1613 1312
rect 1580 1308 1602 1310
rect 1580 1307 1581 1308
rect 1575 1306 1581 1307
rect 830 1302 836 1303
rect 962 1303 968 1304
rect 962 1299 963 1303
rect 967 1302 968 1303
rect 1007 1303 1013 1304
rect 1007 1302 1008 1303
rect 967 1300 1008 1302
rect 967 1299 968 1300
rect 962 1298 968 1299
rect 1007 1299 1008 1300
rect 1012 1299 1013 1303
rect 1007 1298 1013 1299
rect 1047 1303 1053 1304
rect 1047 1299 1048 1303
rect 1052 1302 1053 1303
rect 1375 1303 1381 1304
rect 1447 1303 1453 1304
rect 1052 1300 1058 1302
rect 1052 1299 1053 1300
rect 1047 1298 1053 1299
rect 700 1292 722 1294
rect 727 1295 733 1296
rect 700 1291 701 1292
rect 695 1290 701 1291
rect 727 1291 728 1295
rect 732 1294 733 1295
rect 735 1295 741 1296
rect 735 1294 736 1295
rect 732 1292 736 1294
rect 732 1291 733 1292
rect 727 1290 733 1291
rect 735 1291 736 1292
rect 740 1291 741 1295
rect 735 1290 741 1291
rect 1022 1292 1028 1293
rect 348 1286 350 1290
rect 1022 1288 1023 1292
rect 1027 1288 1028 1292
rect 470 1287 476 1288
rect 1022 1287 1028 1288
rect 470 1286 471 1287
rect 348 1284 471 1286
rect 470 1283 471 1284
rect 475 1283 476 1287
rect 1047 1283 1053 1284
rect 470 1282 476 1283
rect 750 1282 756 1283
rect 186 1279 192 1280
rect 186 1275 187 1279
rect 191 1278 192 1279
rect 734 1279 740 1280
rect 734 1278 735 1279
rect 191 1276 735 1278
rect 191 1275 192 1276
rect 186 1274 192 1275
rect 734 1275 735 1276
rect 739 1275 740 1279
rect 750 1278 751 1282
rect 755 1278 756 1282
rect 750 1277 756 1278
rect 830 1282 836 1283
rect 830 1278 831 1282
rect 835 1278 836 1282
rect 830 1277 836 1278
rect 910 1282 916 1283
rect 910 1278 911 1282
rect 915 1278 916 1282
rect 1019 1279 1025 1280
rect 910 1277 916 1278
rect 982 1277 988 1278
rect 734 1274 740 1275
rect 982 1273 983 1277
rect 987 1273 988 1277
rect 1019 1275 1020 1279
rect 1024 1278 1025 1279
rect 1038 1279 1044 1280
rect 1038 1278 1039 1279
rect 1024 1276 1039 1278
rect 1024 1275 1025 1276
rect 1019 1274 1025 1275
rect 1038 1275 1039 1276
rect 1043 1275 1044 1279
rect 1047 1279 1048 1283
rect 1052 1282 1053 1283
rect 1056 1282 1058 1300
rect 1062 1301 1068 1302
rect 1062 1297 1063 1301
rect 1067 1297 1068 1301
rect 1214 1301 1220 1302
rect 1062 1296 1068 1297
rect 1174 1299 1180 1300
rect 1174 1295 1175 1299
rect 1179 1295 1180 1299
rect 1174 1294 1180 1295
rect 1195 1299 1201 1300
rect 1195 1295 1196 1299
rect 1200 1298 1201 1299
rect 1200 1296 1210 1298
rect 1214 1297 1215 1301
rect 1219 1297 1220 1301
rect 1214 1296 1220 1297
rect 1302 1301 1308 1302
rect 1302 1297 1303 1301
rect 1307 1297 1308 1301
rect 1375 1299 1376 1303
rect 1380 1302 1381 1303
rect 1422 1302 1428 1303
rect 1380 1299 1382 1302
rect 1375 1298 1382 1299
rect 1302 1296 1308 1297
rect 1200 1295 1201 1296
rect 1195 1294 1201 1295
rect 1099 1283 1105 1284
rect 1099 1282 1100 1283
rect 1052 1279 1054 1282
rect 1056 1280 1100 1282
rect 1047 1278 1054 1279
rect 1099 1279 1100 1280
rect 1104 1279 1105 1283
rect 1179 1283 1185 1284
rect 1099 1278 1105 1279
rect 1110 1279 1116 1280
rect 1038 1274 1044 1275
rect 855 1272 861 1273
rect 982 1272 988 1273
rect 102 1271 108 1272
rect 102 1267 103 1271
rect 107 1270 108 1271
rect 574 1271 580 1272
rect 574 1270 575 1271
rect 107 1268 575 1270
rect 107 1267 108 1268
rect 102 1266 108 1267
rect 574 1267 575 1268
rect 579 1270 580 1271
rect 743 1271 749 1272
rect 743 1270 744 1271
rect 579 1268 744 1270
rect 579 1267 580 1268
rect 574 1266 580 1267
rect 743 1267 744 1268
rect 748 1267 749 1271
rect 743 1266 749 1267
rect 758 1271 765 1272
rect 758 1267 759 1271
rect 764 1267 765 1271
rect 758 1266 765 1267
rect 775 1271 781 1272
rect 775 1267 776 1271
rect 780 1270 781 1271
rect 786 1271 792 1272
rect 786 1270 787 1271
rect 780 1268 787 1270
rect 780 1267 781 1268
rect 775 1266 781 1267
rect 786 1267 787 1268
rect 791 1270 792 1271
rect 823 1271 829 1272
rect 823 1270 824 1271
rect 791 1268 824 1270
rect 791 1267 792 1268
rect 786 1266 792 1267
rect 823 1267 824 1268
rect 828 1267 829 1271
rect 823 1266 829 1267
rect 838 1271 845 1272
rect 838 1267 839 1271
rect 844 1267 845 1271
rect 855 1268 856 1272
rect 860 1270 861 1272
rect 866 1271 872 1272
rect 866 1270 867 1271
rect 860 1268 867 1270
rect 855 1267 861 1268
rect 866 1267 867 1268
rect 871 1270 872 1271
rect 894 1271 900 1272
rect 894 1270 895 1271
rect 871 1268 895 1270
rect 871 1267 872 1268
rect 838 1266 845 1267
rect 866 1266 872 1267
rect 894 1267 895 1268
rect 899 1267 900 1271
rect 894 1266 900 1267
rect 903 1271 909 1272
rect 903 1267 904 1271
rect 908 1267 909 1271
rect 903 1266 909 1267
rect 919 1271 925 1272
rect 919 1267 920 1271
rect 924 1267 925 1271
rect 919 1266 925 1267
rect 930 1271 941 1272
rect 930 1267 931 1271
rect 935 1267 936 1271
rect 940 1270 941 1271
rect 962 1271 968 1272
rect 962 1270 963 1271
rect 940 1268 963 1270
rect 940 1267 941 1268
rect 930 1266 941 1267
rect 962 1267 963 1268
rect 967 1267 968 1271
rect 1007 1271 1013 1272
rect 962 1266 968 1267
rect 970 1267 976 1268
rect 734 1263 740 1264
rect 734 1259 735 1263
rect 739 1262 740 1263
rect 904 1262 906 1266
rect 739 1260 906 1262
rect 739 1259 740 1260
rect 734 1258 740 1259
rect 606 1255 612 1256
rect 606 1251 607 1255
rect 611 1254 612 1255
rect 758 1255 764 1256
rect 758 1254 759 1255
rect 611 1252 759 1254
rect 611 1251 612 1252
rect 606 1250 612 1251
rect 758 1251 759 1252
rect 763 1251 764 1255
rect 758 1250 764 1251
rect 807 1255 813 1256
rect 807 1251 808 1255
rect 812 1254 813 1255
rect 838 1255 844 1256
rect 838 1254 839 1255
rect 812 1252 839 1254
rect 812 1251 813 1252
rect 807 1250 813 1251
rect 838 1251 839 1252
rect 843 1254 844 1255
rect 886 1255 892 1256
rect 886 1254 887 1255
rect 843 1252 887 1254
rect 843 1251 844 1252
rect 838 1250 844 1251
rect 886 1251 887 1252
rect 891 1254 892 1255
rect 921 1254 923 1266
rect 970 1263 971 1267
rect 975 1266 976 1267
rect 979 1267 985 1268
rect 979 1266 980 1267
rect 975 1264 980 1266
rect 975 1263 976 1264
rect 970 1262 976 1263
rect 979 1263 980 1264
rect 984 1263 985 1267
rect 1007 1267 1008 1271
rect 1012 1270 1013 1271
rect 1021 1270 1023 1274
rect 1012 1268 1023 1270
rect 1052 1270 1054 1278
rect 1110 1275 1111 1279
rect 1115 1278 1116 1279
rect 1127 1279 1133 1280
rect 1127 1278 1128 1279
rect 1115 1276 1128 1278
rect 1115 1275 1116 1276
rect 1110 1274 1116 1275
rect 1127 1275 1128 1276
rect 1132 1275 1133 1279
rect 1127 1274 1133 1275
rect 1138 1279 1144 1280
rect 1138 1275 1139 1279
rect 1143 1278 1144 1279
rect 1154 1279 1161 1280
rect 1154 1278 1155 1279
rect 1143 1276 1155 1278
rect 1143 1275 1144 1276
rect 1138 1274 1144 1275
rect 1154 1275 1155 1276
rect 1160 1275 1161 1279
rect 1179 1279 1180 1283
rect 1184 1282 1185 1283
rect 1190 1283 1196 1284
rect 1190 1282 1191 1283
rect 1184 1280 1191 1282
rect 1184 1279 1185 1280
rect 1179 1278 1185 1279
rect 1190 1279 1191 1280
rect 1195 1279 1196 1283
rect 1208 1282 1210 1296
rect 1380 1294 1382 1298
rect 1390 1301 1396 1302
rect 1390 1297 1391 1301
rect 1395 1297 1396 1301
rect 1422 1298 1423 1302
rect 1427 1298 1428 1302
rect 1447 1299 1448 1303
rect 1452 1302 1453 1303
rect 1479 1303 1485 1304
rect 1479 1302 1480 1303
rect 1452 1300 1480 1302
rect 1452 1299 1453 1300
rect 1447 1298 1453 1299
rect 1479 1299 1480 1300
rect 1484 1299 1485 1303
rect 1479 1298 1485 1299
rect 1494 1302 1500 1303
rect 1494 1298 1495 1302
rect 1499 1298 1500 1302
rect 1422 1297 1428 1298
rect 1494 1297 1500 1298
rect 1526 1302 1532 1303
rect 1526 1298 1527 1302
rect 1531 1298 1532 1302
rect 1526 1297 1532 1298
rect 1558 1302 1564 1303
rect 1558 1298 1559 1302
rect 1563 1298 1564 1302
rect 1558 1297 1564 1298
rect 1590 1302 1596 1303
rect 1590 1298 1591 1302
rect 1595 1298 1596 1302
rect 1590 1297 1596 1298
rect 1390 1296 1396 1297
rect 1407 1295 1413 1296
rect 1407 1294 1408 1295
rect 1380 1292 1408 1294
rect 1407 1291 1408 1292
rect 1412 1291 1413 1295
rect 1407 1290 1413 1291
rect 1438 1295 1445 1296
rect 1438 1291 1439 1295
rect 1444 1291 1445 1295
rect 1511 1295 1520 1296
rect 1438 1290 1445 1291
rect 1454 1292 1460 1293
rect 1454 1288 1455 1292
rect 1459 1288 1460 1292
rect 1511 1291 1512 1295
rect 1519 1291 1520 1295
rect 1511 1290 1520 1291
rect 1543 1295 1552 1296
rect 1543 1291 1544 1295
rect 1551 1291 1552 1295
rect 1543 1290 1552 1291
rect 1574 1295 1581 1296
rect 1574 1291 1575 1295
rect 1580 1291 1581 1295
rect 1600 1294 1602 1308
rect 1607 1307 1608 1311
rect 1612 1310 1613 1311
rect 1639 1311 1645 1312
rect 1612 1308 1634 1310
rect 1612 1307 1613 1308
rect 1607 1306 1613 1307
rect 1622 1302 1628 1303
rect 1622 1298 1623 1302
rect 1627 1298 1628 1302
rect 1622 1297 1628 1298
rect 1607 1295 1613 1296
rect 1607 1294 1608 1295
rect 1600 1292 1608 1294
rect 1574 1290 1581 1291
rect 1607 1291 1608 1292
rect 1612 1291 1613 1295
rect 1632 1294 1634 1308
rect 1639 1307 1640 1311
rect 1644 1310 1645 1311
rect 1670 1311 1677 1312
rect 1644 1308 1666 1310
rect 1644 1307 1645 1308
rect 1639 1306 1645 1307
rect 1654 1302 1660 1303
rect 1654 1298 1655 1302
rect 1659 1298 1660 1302
rect 1654 1297 1660 1298
rect 1639 1295 1645 1296
rect 1639 1294 1640 1295
rect 1632 1292 1640 1294
rect 1607 1290 1613 1291
rect 1639 1291 1640 1292
rect 1644 1291 1645 1295
rect 1664 1294 1666 1308
rect 1670 1307 1671 1311
rect 1676 1307 1677 1311
rect 1670 1306 1677 1307
rect 1694 1300 1700 1301
rect 1694 1296 1695 1300
rect 1699 1296 1700 1300
rect 1671 1295 1677 1296
rect 1694 1295 1700 1296
rect 1671 1294 1672 1295
rect 1664 1292 1672 1294
rect 1639 1290 1645 1291
rect 1671 1291 1672 1292
rect 1676 1291 1677 1295
rect 1671 1290 1677 1291
rect 1410 1287 1416 1288
rect 1263 1283 1269 1284
rect 1263 1282 1264 1283
rect 1208 1280 1264 1282
rect 1190 1278 1196 1279
rect 1263 1279 1264 1280
rect 1268 1279 1269 1283
rect 1263 1278 1269 1279
rect 1286 1283 1292 1284
rect 1286 1279 1287 1283
rect 1291 1282 1292 1283
rect 1351 1283 1357 1284
rect 1351 1282 1352 1283
rect 1291 1280 1352 1282
rect 1291 1279 1292 1280
rect 1286 1278 1292 1279
rect 1351 1279 1352 1280
rect 1356 1279 1357 1283
rect 1410 1283 1411 1287
rect 1415 1286 1416 1287
rect 1438 1287 1444 1288
rect 1438 1286 1439 1287
rect 1415 1284 1439 1286
rect 1415 1283 1416 1284
rect 1410 1282 1416 1283
rect 1438 1283 1439 1284
rect 1443 1286 1444 1287
rect 1446 1287 1452 1288
rect 1454 1287 1460 1288
rect 1446 1286 1447 1287
rect 1443 1284 1447 1286
rect 1443 1283 1444 1284
rect 1438 1282 1444 1283
rect 1446 1283 1447 1284
rect 1451 1283 1452 1287
rect 1446 1282 1452 1283
rect 1479 1283 1488 1284
rect 1351 1278 1357 1279
rect 1451 1279 1457 1280
rect 1154 1274 1161 1275
rect 1451 1275 1452 1279
rect 1456 1278 1457 1279
rect 1470 1279 1476 1280
rect 1470 1278 1471 1279
rect 1456 1276 1471 1278
rect 1456 1275 1457 1276
rect 1451 1274 1457 1275
rect 1470 1275 1471 1276
rect 1475 1275 1476 1279
rect 1479 1279 1480 1283
rect 1487 1279 1488 1283
rect 1479 1278 1488 1279
rect 1470 1274 1476 1275
rect 1198 1271 1204 1272
rect 1198 1270 1199 1271
rect 1052 1268 1199 1270
rect 1012 1267 1013 1268
rect 1007 1266 1013 1267
rect 1198 1267 1199 1268
rect 1203 1267 1204 1271
rect 1198 1266 1204 1267
rect 979 1262 985 1263
rect 1054 1263 1060 1264
rect 1054 1259 1055 1263
rect 1059 1262 1060 1263
rect 1747 1263 1753 1264
rect 1747 1262 1748 1263
rect 1059 1260 1748 1262
rect 1059 1259 1060 1260
rect 1054 1258 1060 1259
rect 1747 1259 1748 1260
rect 1752 1259 1753 1263
rect 1747 1258 1753 1259
rect 990 1255 996 1256
rect 990 1254 991 1255
rect 891 1252 991 1254
rect 891 1251 892 1252
rect 886 1250 892 1251
rect 990 1251 991 1252
rect 995 1251 996 1255
rect 990 1250 996 1251
rect 918 1247 924 1248
rect 918 1246 919 1247
rect 909 1244 919 1246
rect 918 1243 919 1244
rect 923 1243 924 1247
rect 918 1242 924 1243
rect 79 1235 85 1236
rect 79 1231 80 1235
rect 84 1234 85 1235
rect 190 1235 196 1236
rect 190 1234 191 1235
rect 84 1232 191 1234
rect 84 1231 85 1232
rect 79 1230 85 1231
rect 190 1231 191 1232
rect 195 1231 196 1235
rect 190 1230 196 1231
rect 898 1235 904 1236
rect 898 1231 899 1235
rect 903 1231 904 1235
rect 898 1230 904 1231
rect 990 1231 996 1232
rect 654 1227 660 1228
rect 654 1223 655 1227
rect 659 1226 660 1227
rect 771 1227 777 1228
rect 771 1226 772 1227
rect 659 1224 772 1226
rect 659 1223 660 1224
rect 654 1222 660 1223
rect 771 1223 772 1224
rect 776 1223 777 1227
rect 846 1227 852 1228
rect 771 1222 777 1223
rect 794 1223 805 1224
rect 774 1219 780 1220
rect 590 1215 596 1216
rect 590 1211 591 1215
rect 595 1214 596 1215
rect 626 1215 632 1216
rect 626 1214 627 1215
rect 595 1212 627 1214
rect 595 1211 596 1212
rect 590 1210 596 1211
rect 626 1211 627 1212
rect 631 1211 632 1215
rect 774 1215 775 1219
rect 779 1215 780 1219
rect 794 1219 795 1223
rect 799 1219 800 1223
rect 804 1219 805 1223
rect 846 1223 847 1227
rect 851 1223 852 1227
rect 990 1227 991 1231
rect 995 1230 996 1231
rect 995 1228 1018 1230
rect 995 1227 996 1228
rect 990 1226 996 1227
rect 846 1222 852 1223
rect 1007 1223 1013 1224
rect 1007 1222 1008 1223
rect 794 1218 805 1219
rect 856 1220 1008 1222
rect 774 1214 780 1215
rect 790 1215 796 1216
rect 626 1210 632 1211
rect 735 1211 741 1212
rect 598 1207 604 1208
rect 598 1206 599 1207
rect 545 1204 599 1206
rect 150 1199 157 1200
rect 110 1196 116 1197
rect 110 1192 111 1196
rect 115 1192 116 1196
rect 150 1195 151 1199
rect 156 1195 157 1199
rect 183 1199 189 1200
rect 183 1198 184 1199
rect 176 1196 184 1198
rect 110 1191 116 1192
rect 134 1194 140 1195
rect 150 1194 157 1195
rect 166 1194 172 1195
rect 134 1190 135 1194
rect 139 1190 140 1194
rect 134 1189 140 1190
rect 166 1190 167 1194
rect 171 1190 172 1194
rect 166 1189 172 1190
rect 176 1184 178 1196
rect 183 1195 184 1196
rect 188 1195 189 1199
rect 215 1199 221 1200
rect 215 1198 216 1199
rect 208 1196 216 1198
rect 183 1194 189 1195
rect 198 1194 204 1195
rect 198 1190 199 1194
rect 203 1190 204 1194
rect 198 1189 204 1190
rect 208 1184 210 1196
rect 215 1195 216 1196
rect 220 1195 221 1199
rect 247 1199 253 1200
rect 247 1198 248 1199
rect 240 1196 248 1198
rect 215 1194 221 1195
rect 230 1194 236 1195
rect 230 1190 231 1194
rect 235 1190 236 1194
rect 230 1189 236 1190
rect 240 1184 242 1196
rect 247 1195 248 1196
rect 252 1195 253 1199
rect 279 1199 285 1200
rect 279 1198 280 1199
rect 272 1196 280 1198
rect 247 1194 253 1195
rect 262 1194 268 1195
rect 262 1190 263 1194
rect 267 1190 268 1194
rect 262 1189 268 1190
rect 272 1184 274 1196
rect 279 1195 280 1196
rect 284 1195 285 1199
rect 311 1199 317 1200
rect 311 1198 312 1199
rect 304 1196 312 1198
rect 279 1194 285 1195
rect 294 1194 300 1195
rect 294 1190 295 1194
rect 299 1190 300 1194
rect 294 1189 300 1190
rect 304 1184 306 1196
rect 311 1195 312 1196
rect 316 1195 317 1199
rect 343 1199 349 1200
rect 343 1198 344 1199
rect 336 1196 344 1198
rect 311 1194 317 1195
rect 326 1194 332 1195
rect 326 1190 327 1194
rect 331 1190 332 1194
rect 326 1189 332 1190
rect 336 1184 338 1196
rect 343 1195 344 1196
rect 348 1195 349 1199
rect 375 1199 381 1200
rect 375 1198 376 1199
rect 368 1196 376 1198
rect 343 1194 349 1195
rect 358 1194 364 1195
rect 358 1190 359 1194
rect 363 1190 364 1194
rect 358 1189 364 1190
rect 368 1184 370 1196
rect 375 1195 376 1196
rect 380 1195 381 1199
rect 407 1199 413 1200
rect 407 1198 408 1199
rect 400 1196 408 1198
rect 375 1194 381 1195
rect 390 1194 396 1195
rect 390 1190 391 1194
rect 395 1190 396 1194
rect 390 1189 396 1190
rect 400 1184 402 1196
rect 407 1195 408 1196
rect 412 1195 413 1199
rect 439 1199 445 1200
rect 439 1198 440 1199
rect 432 1196 440 1198
rect 407 1194 413 1195
rect 422 1194 428 1195
rect 422 1190 423 1194
rect 427 1190 428 1194
rect 422 1189 428 1190
rect 432 1184 434 1196
rect 439 1195 440 1196
rect 444 1195 445 1199
rect 471 1199 477 1200
rect 471 1198 472 1199
rect 464 1196 472 1198
rect 439 1194 445 1195
rect 454 1194 460 1195
rect 454 1190 455 1194
rect 459 1190 460 1194
rect 454 1189 460 1190
rect 464 1184 466 1196
rect 471 1195 472 1196
rect 476 1195 477 1199
rect 503 1199 509 1200
rect 503 1198 504 1199
rect 496 1196 504 1198
rect 471 1194 477 1195
rect 486 1194 492 1195
rect 486 1190 487 1194
rect 491 1190 492 1194
rect 486 1189 492 1190
rect 496 1184 498 1196
rect 503 1195 504 1196
rect 508 1195 509 1199
rect 535 1199 541 1200
rect 535 1195 536 1199
rect 540 1198 541 1199
rect 545 1198 547 1204
rect 598 1203 599 1204
rect 603 1203 604 1207
rect 735 1207 736 1211
rect 740 1210 741 1211
rect 758 1211 764 1212
rect 758 1210 759 1211
rect 740 1208 759 1210
rect 740 1207 741 1208
rect 735 1206 741 1207
rect 758 1207 759 1208
rect 763 1207 764 1211
rect 790 1211 791 1215
rect 795 1214 796 1215
rect 856 1214 858 1220
rect 1007 1219 1008 1220
rect 1012 1219 1013 1223
rect 1016 1222 1018 1228
rect 1066 1227 1072 1228
rect 1023 1223 1029 1224
rect 1023 1222 1024 1223
rect 1016 1220 1024 1222
rect 1007 1218 1013 1219
rect 1023 1219 1024 1220
rect 1028 1219 1029 1223
rect 1023 1218 1029 1219
rect 1038 1223 1045 1224
rect 1038 1219 1039 1223
rect 1044 1222 1045 1223
rect 1066 1223 1067 1227
rect 1071 1226 1072 1227
rect 1083 1227 1089 1228
rect 1083 1226 1084 1227
rect 1071 1224 1084 1226
rect 1071 1223 1072 1224
rect 1066 1222 1072 1223
rect 1083 1223 1084 1224
rect 1088 1223 1089 1227
rect 1083 1222 1089 1223
rect 1102 1223 1108 1224
rect 1044 1220 1062 1222
rect 1044 1219 1045 1220
rect 1038 1218 1045 1219
rect 1060 1218 1062 1220
rect 1078 1219 1084 1220
rect 1078 1218 1079 1219
rect 1060 1216 1079 1218
rect 1078 1215 1079 1216
rect 1083 1215 1084 1219
rect 795 1212 858 1214
rect 1014 1214 1020 1215
rect 1078 1214 1084 1215
rect 1086 1219 1092 1220
rect 1086 1215 1087 1219
rect 1091 1215 1092 1219
rect 1102 1219 1103 1223
rect 1107 1222 1108 1223
rect 1111 1223 1117 1224
rect 1111 1222 1112 1223
rect 1107 1220 1112 1222
rect 1107 1219 1108 1220
rect 1102 1218 1108 1219
rect 1111 1219 1112 1220
rect 1116 1222 1117 1223
rect 1190 1223 1196 1224
rect 1190 1222 1191 1223
rect 1116 1220 1191 1222
rect 1116 1219 1117 1220
rect 1111 1218 1117 1219
rect 1190 1219 1191 1220
rect 1195 1219 1196 1223
rect 1190 1218 1196 1219
rect 1287 1223 1293 1224
rect 1287 1219 1288 1223
rect 1292 1222 1293 1223
rect 1446 1223 1452 1224
rect 1446 1222 1447 1223
rect 1292 1220 1447 1222
rect 1292 1219 1293 1220
rect 1287 1218 1293 1219
rect 1446 1219 1447 1220
rect 1451 1219 1452 1223
rect 1446 1218 1452 1219
rect 1086 1214 1092 1215
rect 1195 1215 1204 1216
rect 795 1211 796 1212
rect 790 1210 796 1211
rect 1014 1210 1015 1214
rect 1019 1210 1020 1214
rect 1195 1211 1196 1215
rect 1203 1211 1204 1215
rect 1454 1215 1460 1216
rect 1454 1214 1455 1215
rect 1273 1212 1455 1214
rect 1195 1210 1204 1211
rect 1219 1211 1225 1212
rect 1014 1209 1020 1210
rect 758 1206 764 1207
rect 950 1207 956 1208
rect 598 1202 604 1203
rect 607 1203 613 1204
rect 567 1199 573 1200
rect 567 1198 568 1199
rect 540 1196 547 1198
rect 560 1196 568 1198
rect 540 1195 541 1196
rect 503 1194 509 1195
rect 518 1194 524 1195
rect 535 1194 541 1195
rect 550 1194 556 1195
rect 518 1190 519 1194
rect 523 1190 524 1194
rect 518 1189 524 1190
rect 550 1190 551 1194
rect 555 1190 556 1194
rect 550 1189 556 1190
rect 560 1184 562 1196
rect 567 1195 568 1196
rect 572 1195 573 1199
rect 590 1199 596 1200
rect 590 1195 591 1199
rect 595 1198 596 1199
rect 599 1199 605 1200
rect 599 1198 600 1199
rect 595 1196 600 1198
rect 595 1195 596 1196
rect 567 1194 573 1195
rect 582 1194 588 1195
rect 590 1194 596 1195
rect 599 1195 600 1196
rect 604 1195 605 1199
rect 607 1199 608 1203
rect 612 1202 613 1203
rect 822 1203 828 1204
rect 612 1200 626 1202
rect 704 1200 731 1202
rect 736 1200 763 1202
rect 612 1199 613 1200
rect 607 1198 613 1199
rect 624 1198 626 1200
rect 631 1199 637 1200
rect 631 1198 632 1199
rect 624 1196 632 1198
rect 631 1195 632 1196
rect 636 1195 637 1199
rect 663 1199 669 1200
rect 663 1198 664 1199
rect 656 1196 664 1198
rect 599 1194 605 1195
rect 614 1194 620 1195
rect 631 1194 637 1195
rect 646 1194 652 1195
rect 582 1190 583 1194
rect 587 1190 588 1194
rect 582 1189 588 1190
rect 614 1190 615 1194
rect 619 1190 620 1194
rect 614 1189 620 1190
rect 646 1190 647 1194
rect 651 1190 652 1194
rect 646 1189 652 1190
rect 656 1184 658 1196
rect 663 1195 664 1196
rect 668 1195 669 1199
rect 695 1199 701 1200
rect 695 1198 696 1199
rect 688 1196 696 1198
rect 663 1194 669 1195
rect 678 1194 684 1195
rect 678 1190 679 1194
rect 683 1190 684 1194
rect 678 1189 684 1190
rect 688 1184 690 1196
rect 695 1195 696 1196
rect 700 1195 701 1199
rect 695 1194 701 1195
rect 151 1183 157 1184
rect 110 1179 116 1180
rect 110 1175 111 1179
rect 115 1175 116 1179
rect 151 1179 152 1183
rect 156 1182 157 1183
rect 164 1182 178 1184
rect 183 1183 189 1184
rect 156 1180 166 1182
rect 156 1179 157 1180
rect 151 1178 157 1179
rect 183 1179 184 1183
rect 188 1182 189 1183
rect 196 1182 210 1184
rect 215 1183 221 1184
rect 188 1180 198 1182
rect 188 1179 189 1180
rect 183 1178 189 1179
rect 215 1179 216 1183
rect 220 1182 221 1183
rect 228 1182 242 1184
rect 247 1183 253 1184
rect 220 1180 230 1182
rect 220 1179 221 1180
rect 215 1178 221 1179
rect 247 1179 248 1183
rect 252 1182 253 1183
rect 260 1182 274 1184
rect 279 1183 285 1184
rect 252 1180 262 1182
rect 252 1179 253 1180
rect 247 1178 253 1179
rect 279 1179 280 1183
rect 284 1182 285 1183
rect 292 1182 306 1184
rect 311 1183 317 1184
rect 284 1180 294 1182
rect 284 1179 285 1180
rect 279 1178 285 1179
rect 311 1179 312 1183
rect 316 1182 317 1183
rect 324 1182 338 1184
rect 343 1183 349 1184
rect 316 1180 326 1182
rect 316 1179 317 1180
rect 311 1178 317 1179
rect 343 1179 344 1183
rect 348 1182 349 1183
rect 356 1182 370 1184
rect 375 1183 381 1184
rect 348 1180 358 1182
rect 348 1179 349 1180
rect 343 1178 349 1179
rect 375 1179 376 1183
rect 380 1182 381 1183
rect 388 1182 402 1184
rect 407 1183 413 1184
rect 380 1180 390 1182
rect 380 1179 381 1180
rect 375 1178 381 1179
rect 407 1179 408 1183
rect 412 1182 413 1183
rect 420 1182 434 1184
rect 439 1183 445 1184
rect 412 1180 422 1182
rect 412 1179 413 1180
rect 407 1178 413 1179
rect 439 1179 440 1183
rect 444 1182 445 1183
rect 452 1182 466 1184
rect 471 1183 477 1184
rect 444 1180 454 1182
rect 444 1179 445 1180
rect 439 1178 445 1179
rect 471 1179 472 1183
rect 476 1182 477 1183
rect 484 1182 498 1184
rect 503 1183 509 1184
rect 476 1180 486 1182
rect 476 1179 477 1180
rect 471 1178 477 1179
rect 503 1179 504 1183
rect 508 1179 509 1183
rect 503 1178 509 1179
rect 535 1183 541 1184
rect 535 1179 536 1183
rect 540 1182 541 1183
rect 548 1182 562 1184
rect 566 1183 573 1184
rect 540 1180 550 1182
rect 540 1179 541 1180
rect 535 1178 541 1179
rect 566 1179 567 1183
rect 572 1179 573 1183
rect 566 1178 573 1179
rect 598 1183 605 1184
rect 598 1179 599 1183
rect 604 1179 605 1183
rect 598 1178 605 1179
rect 631 1183 637 1184
rect 631 1179 632 1183
rect 636 1182 637 1183
rect 644 1182 658 1184
rect 663 1183 669 1184
rect 636 1180 646 1182
rect 636 1179 637 1180
rect 631 1178 637 1179
rect 663 1179 664 1183
rect 668 1182 669 1183
rect 676 1182 690 1184
rect 695 1183 701 1184
rect 668 1180 678 1182
rect 668 1179 669 1180
rect 663 1178 669 1179
rect 695 1179 696 1183
rect 700 1182 701 1183
rect 704 1182 706 1200
rect 727 1199 733 1200
rect 727 1195 728 1199
rect 732 1195 733 1199
rect 710 1194 716 1195
rect 727 1194 733 1195
rect 710 1190 711 1194
rect 715 1190 716 1194
rect 710 1189 716 1190
rect 700 1180 706 1182
rect 727 1183 733 1184
rect 700 1179 701 1180
rect 695 1178 701 1179
rect 727 1179 728 1183
rect 732 1182 733 1183
rect 736 1182 738 1200
rect 759 1199 765 1200
rect 759 1195 760 1199
rect 764 1195 765 1199
rect 822 1199 823 1203
rect 827 1202 828 1203
rect 935 1203 941 1204
rect 935 1202 936 1203
rect 827 1200 936 1202
rect 827 1199 828 1200
rect 822 1198 828 1199
rect 935 1199 936 1200
rect 940 1199 941 1203
rect 950 1203 951 1207
rect 955 1206 956 1207
rect 959 1207 965 1208
rect 959 1206 960 1207
rect 955 1204 960 1206
rect 955 1203 956 1204
rect 950 1202 956 1203
rect 959 1203 960 1204
rect 964 1203 965 1207
rect 959 1202 965 1203
rect 1190 1207 1196 1208
rect 1190 1203 1191 1207
rect 1195 1206 1196 1207
rect 1219 1207 1220 1211
rect 1224 1207 1225 1211
rect 1219 1206 1225 1207
rect 1262 1207 1268 1208
rect 1262 1206 1263 1207
rect 1195 1204 1263 1206
rect 1195 1203 1196 1204
rect 1190 1202 1196 1203
rect 1262 1203 1263 1204
rect 1267 1203 1268 1207
rect 1262 1202 1268 1203
rect 1145 1200 1170 1202
rect 1273 1200 1275 1212
rect 1454 1211 1455 1212
rect 1459 1211 1460 1215
rect 1454 1210 1460 1211
rect 1287 1207 1293 1208
rect 1287 1203 1288 1207
rect 1292 1206 1293 1207
rect 1295 1207 1301 1208
rect 1295 1206 1296 1207
rect 1292 1204 1296 1206
rect 1292 1203 1293 1204
rect 1287 1202 1293 1203
rect 1295 1203 1296 1204
rect 1300 1203 1301 1207
rect 1414 1207 1420 1208
rect 1414 1206 1415 1207
rect 1368 1204 1415 1206
rect 1295 1202 1301 1203
rect 1350 1203 1356 1204
rect 1350 1202 1351 1203
rect 1336 1200 1351 1202
rect 935 1198 941 1199
rect 990 1199 997 1200
rect 958 1197 964 1198
rect 742 1194 748 1195
rect 759 1194 765 1195
rect 810 1195 816 1196
rect 742 1190 743 1194
rect 747 1190 748 1194
rect 742 1189 748 1190
rect 790 1191 796 1192
rect 790 1187 791 1191
rect 795 1190 796 1191
rect 799 1191 805 1192
rect 799 1190 800 1191
rect 795 1188 800 1190
rect 795 1187 796 1188
rect 790 1186 796 1187
rect 799 1187 800 1188
rect 804 1187 805 1191
rect 810 1191 811 1195
rect 815 1191 816 1195
rect 958 1193 959 1197
rect 963 1193 964 1197
rect 990 1195 991 1199
rect 996 1195 997 1199
rect 1143 1199 1149 1200
rect 1143 1195 1144 1199
rect 1148 1195 1149 1199
rect 990 1194 997 1195
rect 1126 1194 1132 1195
rect 1143 1194 1149 1195
rect 1158 1194 1164 1195
rect 958 1192 964 1193
rect 810 1190 816 1191
rect 1078 1191 1084 1192
rect 799 1186 805 1187
rect 1066 1187 1072 1188
rect 732 1180 738 1182
rect 758 1183 765 1184
rect 732 1179 733 1180
rect 727 1178 733 1179
rect 758 1179 759 1183
rect 764 1179 765 1183
rect 1066 1183 1067 1187
rect 1071 1183 1072 1187
rect 1078 1187 1079 1191
rect 1083 1190 1084 1191
rect 1111 1191 1117 1192
rect 1111 1190 1112 1191
rect 1083 1188 1112 1190
rect 1083 1187 1084 1188
rect 1078 1186 1084 1187
rect 1111 1187 1112 1188
rect 1116 1187 1117 1191
rect 1126 1190 1127 1194
rect 1131 1190 1132 1194
rect 1126 1189 1132 1190
rect 1158 1190 1159 1194
rect 1163 1190 1164 1194
rect 1158 1189 1164 1190
rect 1111 1186 1117 1187
rect 1066 1182 1072 1183
rect 1142 1183 1149 1184
rect 758 1178 765 1179
rect 838 1180 844 1181
rect 110 1174 116 1175
rect 134 1177 140 1178
rect 134 1173 135 1177
rect 139 1173 140 1177
rect 134 1172 140 1173
rect 166 1177 172 1178
rect 166 1173 167 1177
rect 171 1173 172 1177
rect 166 1172 172 1173
rect 198 1177 204 1178
rect 198 1173 199 1177
rect 203 1173 204 1177
rect 198 1172 204 1173
rect 230 1177 236 1178
rect 230 1173 231 1177
rect 235 1173 236 1177
rect 230 1172 236 1173
rect 262 1177 268 1178
rect 262 1173 263 1177
rect 267 1173 268 1177
rect 262 1172 268 1173
rect 294 1177 300 1178
rect 294 1173 295 1177
rect 299 1173 300 1177
rect 294 1172 300 1173
rect 326 1177 332 1178
rect 326 1173 327 1177
rect 331 1173 332 1177
rect 326 1172 332 1173
rect 358 1177 364 1178
rect 358 1173 359 1177
rect 363 1173 364 1177
rect 358 1172 364 1173
rect 390 1177 396 1178
rect 390 1173 391 1177
rect 395 1173 396 1177
rect 390 1172 396 1173
rect 422 1177 428 1178
rect 422 1173 423 1177
rect 427 1173 428 1177
rect 422 1172 428 1173
rect 454 1177 460 1178
rect 454 1173 455 1177
rect 459 1173 460 1177
rect 454 1172 460 1173
rect 486 1177 492 1178
rect 486 1173 487 1177
rect 491 1173 492 1177
rect 486 1172 492 1173
rect 442 1171 448 1172
rect 442 1167 443 1171
rect 447 1170 448 1171
rect 504 1170 506 1178
rect 518 1177 524 1178
rect 518 1173 519 1177
rect 523 1173 524 1177
rect 518 1172 524 1173
rect 550 1177 556 1178
rect 550 1173 551 1177
rect 555 1173 556 1177
rect 550 1172 556 1173
rect 582 1177 588 1178
rect 582 1173 583 1177
rect 587 1173 588 1177
rect 582 1172 588 1173
rect 614 1177 620 1178
rect 614 1173 615 1177
rect 619 1173 620 1177
rect 614 1172 620 1173
rect 646 1177 652 1178
rect 646 1173 647 1177
rect 651 1173 652 1177
rect 646 1172 652 1173
rect 678 1177 684 1178
rect 678 1173 679 1177
rect 683 1173 684 1177
rect 678 1172 684 1173
rect 710 1177 716 1178
rect 710 1173 711 1177
rect 715 1173 716 1177
rect 710 1172 716 1173
rect 742 1177 748 1178
rect 742 1173 743 1177
rect 747 1173 748 1177
rect 838 1176 839 1180
rect 843 1176 844 1180
rect 838 1175 844 1176
rect 930 1179 941 1180
rect 930 1175 931 1179
rect 935 1175 936 1179
rect 940 1175 941 1179
rect 1142 1179 1143 1183
rect 1148 1179 1149 1183
rect 1168 1182 1170 1200
rect 1175 1199 1181 1200
rect 1175 1195 1176 1199
rect 1180 1198 1181 1199
rect 1198 1199 1204 1200
rect 1198 1198 1199 1199
rect 1180 1196 1199 1198
rect 1180 1195 1181 1196
rect 1175 1194 1181 1195
rect 1198 1195 1199 1196
rect 1203 1195 1204 1199
rect 1271 1199 1277 1200
rect 1198 1194 1204 1195
rect 1214 1197 1220 1198
rect 1214 1193 1215 1197
rect 1219 1193 1220 1197
rect 1214 1192 1220 1193
rect 1235 1195 1244 1196
rect 1271 1195 1272 1199
rect 1276 1195 1277 1199
rect 1327 1199 1333 1200
rect 1235 1191 1236 1195
rect 1243 1191 1244 1195
rect 1235 1190 1244 1191
rect 1254 1194 1260 1195
rect 1271 1194 1277 1195
rect 1294 1197 1300 1198
rect 1254 1190 1255 1194
rect 1259 1190 1260 1194
rect 1294 1193 1295 1197
rect 1299 1193 1300 1197
rect 1327 1195 1328 1199
rect 1332 1198 1333 1199
rect 1336 1198 1338 1200
rect 1350 1199 1351 1200
rect 1355 1199 1356 1203
rect 1350 1198 1356 1199
rect 1359 1199 1365 1200
rect 1332 1196 1338 1198
rect 1332 1195 1333 1196
rect 1359 1195 1360 1199
rect 1364 1198 1365 1199
rect 1368 1198 1370 1204
rect 1414 1203 1415 1204
rect 1419 1203 1420 1207
rect 1414 1202 1420 1203
rect 1546 1203 1552 1204
rect 1391 1199 1397 1200
rect 1391 1198 1392 1199
rect 1364 1196 1370 1198
rect 1384 1196 1392 1198
rect 1364 1195 1365 1196
rect 1327 1194 1333 1195
rect 1342 1194 1348 1195
rect 1359 1194 1365 1195
rect 1374 1194 1380 1195
rect 1294 1192 1300 1193
rect 1254 1189 1260 1190
rect 1342 1190 1343 1194
rect 1347 1190 1348 1194
rect 1342 1189 1348 1190
rect 1374 1190 1375 1194
rect 1379 1190 1380 1194
rect 1374 1189 1380 1190
rect 1384 1184 1386 1196
rect 1391 1195 1392 1196
rect 1396 1195 1397 1199
rect 1423 1199 1429 1200
rect 1423 1195 1424 1199
rect 1428 1195 1429 1199
rect 1455 1199 1461 1200
rect 1455 1195 1456 1199
rect 1460 1198 1461 1199
rect 1495 1199 1504 1200
rect 1460 1196 1474 1198
rect 1460 1195 1461 1196
rect 1391 1194 1397 1195
rect 1406 1194 1412 1195
rect 1423 1194 1429 1195
rect 1438 1194 1444 1195
rect 1455 1194 1461 1195
rect 1406 1190 1407 1194
rect 1411 1190 1412 1194
rect 1406 1189 1412 1190
rect 1438 1190 1439 1194
rect 1443 1190 1444 1194
rect 1438 1189 1444 1190
rect 1472 1186 1474 1196
rect 1495 1195 1496 1199
rect 1503 1195 1504 1199
rect 1535 1199 1544 1200
rect 1535 1195 1536 1199
rect 1543 1195 1544 1199
rect 1546 1199 1547 1203
rect 1551 1202 1552 1203
rect 1551 1200 1570 1202
rect 1609 1200 1634 1202
rect 1551 1199 1552 1200
rect 1546 1198 1552 1199
rect 1568 1198 1570 1200
rect 1575 1199 1581 1200
rect 1575 1198 1576 1199
rect 1568 1196 1576 1198
rect 1575 1195 1576 1196
rect 1580 1195 1581 1199
rect 1607 1199 1613 1200
rect 1607 1195 1608 1199
rect 1612 1195 1613 1199
rect 1478 1194 1484 1195
rect 1495 1194 1504 1195
rect 1518 1194 1524 1195
rect 1535 1194 1544 1195
rect 1558 1194 1564 1195
rect 1575 1194 1581 1195
rect 1590 1194 1596 1195
rect 1607 1194 1613 1195
rect 1622 1194 1628 1195
rect 1478 1190 1479 1194
rect 1483 1190 1484 1194
rect 1478 1189 1484 1190
rect 1518 1190 1519 1194
rect 1523 1190 1524 1194
rect 1518 1189 1524 1190
rect 1558 1190 1559 1194
rect 1563 1190 1564 1194
rect 1558 1189 1564 1190
rect 1590 1190 1591 1194
rect 1595 1190 1596 1194
rect 1590 1189 1596 1190
rect 1622 1190 1623 1194
rect 1627 1190 1628 1194
rect 1622 1189 1628 1190
rect 1472 1184 1478 1186
rect 1175 1183 1181 1184
rect 1175 1182 1176 1183
rect 1168 1180 1176 1182
rect 1142 1178 1149 1179
rect 1175 1179 1176 1180
rect 1180 1179 1181 1183
rect 1175 1178 1181 1179
rect 1271 1183 1277 1184
rect 1271 1179 1272 1183
rect 1276 1182 1277 1183
rect 1286 1183 1292 1184
rect 1286 1182 1287 1183
rect 1276 1180 1287 1182
rect 1276 1179 1277 1180
rect 1271 1178 1277 1179
rect 1286 1179 1287 1180
rect 1291 1179 1292 1183
rect 1286 1178 1292 1179
rect 1359 1183 1365 1184
rect 1359 1179 1360 1183
rect 1364 1182 1365 1183
rect 1372 1182 1386 1184
rect 1391 1183 1397 1184
rect 1364 1180 1374 1182
rect 1364 1179 1365 1180
rect 1359 1178 1365 1179
rect 1391 1179 1392 1183
rect 1396 1182 1397 1183
rect 1418 1183 1429 1184
rect 1396 1180 1402 1182
rect 1396 1179 1397 1180
rect 1391 1178 1397 1179
rect 1126 1177 1132 1178
rect 930 1174 941 1175
rect 1006 1176 1012 1177
rect 742 1172 748 1173
rect 774 1172 780 1173
rect 447 1168 506 1170
rect 774 1168 775 1172
rect 779 1168 780 1172
rect 1006 1172 1007 1176
rect 1011 1172 1012 1176
rect 1126 1173 1127 1177
rect 1131 1173 1132 1177
rect 1006 1171 1012 1172
rect 1086 1172 1092 1173
rect 1126 1172 1132 1173
rect 1158 1177 1164 1178
rect 1254 1177 1260 1178
rect 1158 1173 1159 1177
rect 1163 1173 1164 1177
rect 1158 1172 1164 1173
rect 1198 1176 1204 1177
rect 1198 1172 1199 1176
rect 1203 1172 1204 1176
rect 1254 1173 1255 1177
rect 1259 1173 1260 1177
rect 1254 1172 1260 1173
rect 1342 1177 1348 1178
rect 1342 1173 1343 1177
rect 1347 1173 1348 1177
rect 1342 1172 1348 1173
rect 1374 1177 1380 1178
rect 1374 1173 1375 1177
rect 1379 1173 1380 1177
rect 1374 1172 1380 1173
rect 447 1167 448 1168
rect 774 1167 780 1168
rect 974 1170 980 1171
rect 442 1166 448 1167
rect 974 1166 975 1170
rect 979 1166 980 1170
rect 1086 1168 1087 1172
rect 1091 1168 1092 1172
rect 1198 1171 1204 1172
rect 1086 1167 1092 1168
rect 1310 1170 1316 1171
rect 974 1165 980 1166
rect 1310 1166 1311 1170
rect 1315 1166 1316 1170
rect 1400 1170 1402 1180
rect 1418 1179 1419 1183
rect 1423 1179 1424 1183
rect 1428 1179 1429 1183
rect 1418 1178 1429 1179
rect 1454 1183 1461 1184
rect 1454 1179 1455 1183
rect 1460 1179 1461 1183
rect 1476 1182 1490 1184
rect 1495 1183 1501 1184
rect 1495 1182 1496 1183
rect 1488 1180 1496 1182
rect 1454 1178 1461 1179
rect 1495 1179 1496 1180
rect 1500 1179 1501 1183
rect 1495 1178 1501 1179
rect 1535 1183 1541 1184
rect 1535 1179 1536 1183
rect 1540 1182 1541 1183
rect 1546 1183 1552 1184
rect 1546 1182 1547 1183
rect 1540 1180 1547 1182
rect 1540 1179 1541 1180
rect 1535 1178 1541 1179
rect 1546 1179 1547 1180
rect 1551 1179 1552 1183
rect 1546 1178 1552 1179
rect 1574 1183 1581 1184
rect 1574 1179 1575 1183
rect 1580 1179 1581 1183
rect 1574 1178 1581 1179
rect 1607 1183 1616 1184
rect 1607 1179 1608 1183
rect 1615 1179 1616 1183
rect 1632 1182 1634 1200
rect 1639 1199 1645 1200
rect 1639 1195 1640 1199
rect 1644 1198 1645 1199
rect 1670 1199 1677 1200
rect 1644 1196 1650 1198
rect 1644 1195 1645 1196
rect 1639 1194 1645 1195
rect 1648 1186 1650 1196
rect 1670 1195 1671 1199
rect 1676 1195 1677 1199
rect 1654 1194 1660 1195
rect 1670 1194 1677 1195
rect 1694 1196 1700 1197
rect 1654 1190 1655 1194
rect 1659 1190 1660 1194
rect 1694 1192 1695 1196
rect 1699 1192 1700 1196
rect 1694 1191 1700 1192
rect 1654 1189 1660 1190
rect 1648 1184 1654 1186
rect 1639 1183 1645 1184
rect 1639 1182 1640 1183
rect 1632 1180 1640 1182
rect 1607 1178 1616 1179
rect 1639 1179 1640 1180
rect 1644 1179 1645 1183
rect 1652 1182 1666 1184
rect 1671 1183 1677 1184
rect 1671 1182 1672 1183
rect 1664 1180 1672 1182
rect 1639 1178 1645 1179
rect 1671 1179 1672 1180
rect 1676 1179 1677 1183
rect 1671 1178 1677 1179
rect 1694 1179 1700 1180
rect 1406 1177 1412 1178
rect 1406 1173 1407 1177
rect 1411 1173 1412 1177
rect 1406 1172 1412 1173
rect 1438 1177 1444 1178
rect 1438 1173 1439 1177
rect 1443 1173 1444 1177
rect 1438 1172 1444 1173
rect 1478 1177 1484 1178
rect 1478 1173 1479 1177
rect 1483 1173 1484 1177
rect 1478 1172 1484 1173
rect 1518 1177 1524 1178
rect 1518 1173 1519 1177
rect 1523 1173 1524 1177
rect 1518 1172 1524 1173
rect 1558 1177 1564 1178
rect 1558 1173 1559 1177
rect 1563 1173 1564 1177
rect 1558 1172 1564 1173
rect 1590 1177 1596 1178
rect 1590 1173 1591 1177
rect 1595 1173 1596 1177
rect 1590 1172 1596 1173
rect 1622 1177 1628 1178
rect 1622 1173 1623 1177
rect 1627 1173 1628 1177
rect 1622 1172 1628 1173
rect 1654 1177 1660 1178
rect 1654 1173 1655 1177
rect 1659 1173 1660 1177
rect 1694 1175 1695 1179
rect 1699 1175 1700 1179
rect 1694 1174 1700 1175
rect 1654 1172 1660 1173
rect 1430 1171 1436 1172
rect 1430 1170 1431 1171
rect 1400 1168 1431 1170
rect 1430 1167 1431 1168
rect 1435 1167 1436 1171
rect 1430 1166 1436 1167
rect 1446 1171 1452 1172
rect 1446 1167 1447 1171
rect 1451 1170 1452 1171
rect 1743 1171 1749 1172
rect 1743 1170 1744 1171
rect 1451 1168 1744 1170
rect 1451 1167 1452 1168
rect 1446 1166 1452 1167
rect 1743 1167 1744 1168
rect 1748 1167 1749 1171
rect 1743 1166 1749 1167
rect 1310 1165 1316 1166
rect 542 1163 548 1164
rect 542 1159 543 1163
rect 547 1162 548 1163
rect 798 1163 804 1164
rect 798 1162 799 1163
rect 547 1160 799 1162
rect 547 1159 548 1160
rect 542 1158 548 1159
rect 798 1159 799 1160
rect 803 1159 804 1163
rect 798 1158 804 1159
rect 814 1163 820 1164
rect 814 1159 815 1163
rect 819 1162 820 1163
rect 951 1163 957 1164
rect 951 1162 952 1163
rect 819 1160 952 1162
rect 819 1159 820 1160
rect 814 1158 820 1159
rect 951 1159 952 1160
rect 956 1159 957 1163
rect 951 1158 957 1159
rect 1286 1163 1293 1164
rect 1286 1159 1287 1163
rect 1292 1159 1293 1163
rect 1286 1158 1293 1159
rect 807 1155 813 1156
rect 807 1154 808 1155
rect 740 1152 808 1154
rect 414 1151 420 1152
rect 414 1147 415 1151
rect 419 1150 420 1151
rect 740 1150 742 1152
rect 807 1151 808 1152
rect 812 1151 813 1155
rect 807 1150 813 1151
rect 419 1148 742 1150
rect 419 1147 420 1148
rect 414 1146 420 1147
rect 954 1143 960 1144
rect 954 1139 955 1143
rect 959 1142 960 1143
rect 1142 1143 1148 1144
rect 1142 1142 1143 1143
rect 959 1140 1143 1142
rect 959 1139 960 1140
rect 954 1138 960 1139
rect 1142 1139 1143 1140
rect 1147 1139 1148 1143
rect 1142 1138 1148 1139
rect 282 1131 288 1132
rect 282 1127 283 1131
rect 287 1130 288 1131
rect 287 1128 546 1130
rect 287 1127 288 1128
rect 282 1126 288 1127
rect 134 1123 140 1124
rect 110 1121 116 1122
rect 110 1117 111 1121
rect 115 1117 116 1121
rect 134 1119 135 1123
rect 139 1119 140 1123
rect 134 1118 140 1119
rect 166 1123 172 1124
rect 166 1119 167 1123
rect 171 1119 172 1123
rect 166 1118 172 1119
rect 198 1123 204 1124
rect 198 1119 199 1123
rect 203 1119 204 1123
rect 198 1118 204 1119
rect 230 1123 236 1124
rect 230 1119 231 1123
rect 235 1119 236 1123
rect 230 1118 236 1119
rect 262 1123 268 1124
rect 262 1119 263 1123
rect 267 1119 268 1123
rect 262 1118 268 1119
rect 294 1123 300 1124
rect 294 1119 295 1123
rect 299 1119 300 1123
rect 294 1118 300 1119
rect 326 1123 332 1124
rect 326 1119 327 1123
rect 331 1119 332 1123
rect 326 1118 332 1119
rect 358 1123 364 1124
rect 358 1119 359 1123
rect 363 1119 364 1123
rect 358 1118 364 1119
rect 390 1123 396 1124
rect 390 1119 391 1123
rect 395 1119 396 1123
rect 390 1118 396 1119
rect 422 1123 428 1124
rect 422 1119 423 1123
rect 427 1119 428 1123
rect 422 1118 428 1119
rect 454 1123 460 1124
rect 454 1119 455 1123
rect 459 1119 460 1123
rect 454 1118 460 1119
rect 486 1123 492 1124
rect 486 1119 487 1123
rect 491 1119 492 1123
rect 486 1118 492 1119
rect 518 1123 524 1124
rect 518 1119 519 1123
rect 523 1119 524 1123
rect 518 1118 524 1119
rect 110 1116 116 1117
rect 151 1115 157 1116
rect 151 1111 152 1115
rect 156 1114 157 1115
rect 183 1115 189 1116
rect 156 1112 178 1114
rect 156 1111 157 1112
rect 151 1110 157 1111
rect 134 1106 140 1107
rect 110 1104 116 1105
rect 110 1100 111 1104
rect 115 1100 116 1104
rect 134 1102 135 1106
rect 139 1102 140 1106
rect 134 1101 140 1102
rect 166 1106 172 1107
rect 166 1102 167 1106
rect 171 1102 172 1106
rect 166 1101 172 1102
rect 110 1099 116 1100
rect 151 1099 157 1100
rect 151 1095 152 1099
rect 156 1095 157 1099
rect 176 1098 178 1112
rect 183 1111 184 1115
rect 188 1114 189 1115
rect 215 1115 221 1116
rect 188 1112 210 1114
rect 188 1111 189 1112
rect 183 1110 189 1111
rect 198 1106 204 1107
rect 198 1102 199 1106
rect 203 1102 204 1106
rect 198 1101 204 1102
rect 183 1099 189 1100
rect 183 1098 184 1099
rect 176 1096 184 1098
rect 151 1094 157 1095
rect 183 1095 184 1096
rect 188 1095 189 1099
rect 208 1098 210 1112
rect 215 1111 216 1115
rect 220 1114 221 1115
rect 246 1115 253 1116
rect 220 1112 242 1114
rect 220 1111 221 1112
rect 215 1110 221 1111
rect 230 1106 236 1107
rect 230 1102 231 1106
rect 235 1102 236 1106
rect 230 1101 236 1102
rect 215 1099 221 1100
rect 215 1098 216 1099
rect 208 1096 216 1098
rect 183 1094 189 1095
rect 215 1095 216 1096
rect 220 1095 221 1099
rect 240 1098 242 1112
rect 246 1111 247 1115
rect 252 1111 253 1115
rect 246 1110 253 1111
rect 255 1115 261 1116
rect 255 1111 256 1115
rect 260 1114 261 1115
rect 279 1115 285 1116
rect 279 1114 280 1115
rect 260 1112 280 1114
rect 260 1111 261 1112
rect 255 1110 261 1111
rect 279 1111 280 1112
rect 284 1111 285 1115
rect 279 1110 285 1111
rect 287 1115 293 1116
rect 287 1111 288 1115
rect 292 1114 293 1115
rect 311 1115 317 1116
rect 311 1114 312 1115
rect 292 1112 312 1114
rect 292 1111 293 1112
rect 287 1110 293 1111
rect 311 1111 312 1112
rect 316 1111 317 1115
rect 343 1115 349 1116
rect 343 1114 344 1115
rect 311 1110 317 1111
rect 336 1112 344 1114
rect 262 1106 268 1107
rect 262 1102 263 1106
rect 267 1102 268 1106
rect 262 1101 268 1102
rect 294 1106 300 1107
rect 294 1102 295 1106
rect 299 1102 300 1106
rect 294 1101 300 1102
rect 326 1106 332 1107
rect 326 1102 327 1106
rect 331 1102 332 1106
rect 326 1101 332 1102
rect 247 1099 253 1100
rect 247 1098 248 1099
rect 240 1096 248 1098
rect 215 1094 221 1095
rect 247 1095 248 1096
rect 252 1095 253 1099
rect 247 1094 253 1095
rect 279 1099 288 1100
rect 279 1095 280 1099
rect 287 1095 288 1099
rect 279 1094 288 1095
rect 311 1099 317 1100
rect 311 1095 312 1099
rect 316 1098 317 1099
rect 336 1098 338 1112
rect 343 1111 344 1112
rect 348 1111 349 1115
rect 375 1115 381 1116
rect 375 1114 376 1115
rect 343 1110 349 1111
rect 368 1112 376 1114
rect 358 1106 364 1107
rect 358 1102 359 1106
rect 363 1102 364 1106
rect 358 1101 364 1102
rect 316 1096 338 1098
rect 343 1099 349 1100
rect 316 1095 317 1096
rect 311 1094 317 1095
rect 343 1095 344 1099
rect 348 1098 349 1099
rect 368 1098 370 1112
rect 375 1111 376 1112
rect 380 1111 381 1115
rect 407 1115 413 1116
rect 407 1114 408 1115
rect 375 1110 381 1111
rect 400 1112 408 1114
rect 390 1106 396 1107
rect 390 1102 391 1106
rect 395 1102 396 1106
rect 390 1101 396 1102
rect 348 1096 370 1098
rect 375 1099 381 1100
rect 348 1095 349 1096
rect 343 1094 349 1095
rect 375 1095 376 1099
rect 380 1098 381 1099
rect 400 1098 402 1112
rect 407 1111 408 1112
rect 412 1111 413 1115
rect 407 1110 413 1111
rect 439 1115 445 1116
rect 439 1111 440 1115
rect 444 1114 445 1115
rect 471 1115 477 1116
rect 444 1112 466 1114
rect 444 1111 445 1112
rect 439 1110 445 1111
rect 422 1106 428 1107
rect 422 1102 423 1106
rect 427 1102 428 1106
rect 422 1101 428 1102
rect 454 1106 460 1107
rect 454 1102 455 1106
rect 459 1102 460 1106
rect 454 1101 460 1102
rect 380 1096 402 1098
rect 407 1099 413 1100
rect 380 1095 381 1096
rect 375 1094 381 1095
rect 407 1095 408 1099
rect 412 1098 413 1099
rect 439 1099 448 1100
rect 412 1096 434 1098
rect 412 1095 413 1096
rect 407 1094 413 1095
rect 153 1090 155 1094
rect 287 1091 293 1092
rect 287 1090 288 1091
rect 153 1088 288 1090
rect 287 1087 288 1088
rect 292 1087 293 1091
rect 432 1090 434 1096
rect 439 1095 440 1099
rect 447 1095 448 1099
rect 464 1098 466 1112
rect 471 1111 472 1115
rect 476 1114 477 1115
rect 503 1115 509 1116
rect 476 1112 498 1114
rect 476 1111 477 1112
rect 471 1110 477 1111
rect 486 1106 492 1107
rect 486 1102 487 1106
rect 491 1102 492 1106
rect 486 1101 492 1102
rect 471 1099 477 1100
rect 471 1098 472 1099
rect 464 1096 472 1098
rect 439 1094 448 1095
rect 471 1095 472 1096
rect 476 1095 477 1099
rect 496 1098 498 1112
rect 503 1111 504 1115
rect 508 1114 509 1115
rect 534 1115 541 1116
rect 508 1112 530 1114
rect 508 1111 509 1112
rect 503 1110 509 1111
rect 518 1106 524 1107
rect 518 1102 519 1106
rect 523 1102 524 1106
rect 518 1101 524 1102
rect 503 1099 509 1100
rect 503 1098 504 1099
rect 496 1096 504 1098
rect 471 1094 477 1095
rect 503 1095 504 1096
rect 508 1095 509 1099
rect 528 1098 530 1112
rect 534 1111 535 1115
rect 540 1111 541 1115
rect 544 1114 546 1128
rect 1246 1128 1252 1129
rect 846 1126 852 1127
rect 582 1124 588 1125
rect 550 1123 556 1124
rect 550 1119 551 1123
rect 555 1119 556 1123
rect 582 1120 583 1124
rect 587 1120 588 1124
rect 798 1124 804 1125
rect 582 1119 588 1120
rect 686 1120 692 1121
rect 798 1120 799 1124
rect 803 1120 804 1124
rect 846 1122 847 1126
rect 851 1122 852 1126
rect 998 1124 1004 1125
rect 1094 1124 1100 1125
rect 1166 1124 1172 1125
rect 846 1121 852 1122
rect 934 1123 940 1124
rect 550 1118 556 1119
rect 686 1116 687 1120
rect 691 1116 692 1120
rect 567 1115 573 1116
rect 567 1114 568 1115
rect 544 1112 568 1114
rect 534 1110 541 1111
rect 567 1111 568 1112
rect 572 1111 573 1115
rect 654 1115 660 1116
rect 686 1115 692 1116
rect 782 1119 789 1120
rect 798 1119 804 1120
rect 815 1119 821 1120
rect 782 1115 783 1119
rect 788 1115 789 1119
rect 654 1114 655 1115
rect 645 1112 655 1114
rect 567 1110 573 1111
rect 654 1111 655 1112
rect 659 1111 660 1115
rect 782 1114 789 1115
rect 815 1115 816 1119
rect 820 1118 821 1119
rect 854 1119 860 1120
rect 854 1118 855 1119
rect 820 1116 855 1118
rect 820 1115 821 1116
rect 815 1114 821 1115
rect 854 1115 855 1116
rect 859 1115 860 1119
rect 934 1119 935 1123
rect 939 1119 940 1123
rect 934 1118 940 1119
rect 966 1123 972 1124
rect 966 1119 967 1123
rect 971 1119 972 1123
rect 998 1120 999 1124
rect 1003 1120 1004 1124
rect 1030 1123 1036 1124
rect 998 1119 1004 1120
rect 1014 1119 1021 1120
rect 966 1118 972 1119
rect 854 1114 860 1115
rect 951 1115 957 1116
rect 654 1110 660 1111
rect 951 1111 952 1115
rect 956 1114 957 1115
rect 983 1115 989 1116
rect 956 1112 978 1114
rect 956 1111 957 1112
rect 951 1110 957 1111
rect 550 1106 556 1107
rect 934 1106 940 1107
rect 550 1102 551 1106
rect 555 1102 556 1106
rect 550 1101 556 1102
rect 658 1105 664 1106
rect 658 1101 659 1105
rect 663 1101 664 1105
rect 934 1102 935 1106
rect 939 1102 940 1106
rect 658 1100 664 1101
rect 798 1101 804 1102
rect 934 1101 940 1102
rect 966 1106 972 1107
rect 966 1102 967 1106
rect 971 1102 972 1106
rect 966 1101 972 1102
rect 535 1099 541 1100
rect 535 1098 536 1099
rect 528 1096 536 1098
rect 503 1094 509 1095
rect 535 1095 536 1096
rect 540 1095 541 1099
rect 535 1094 541 1095
rect 566 1099 573 1100
rect 566 1095 567 1099
rect 572 1095 573 1099
rect 798 1097 799 1101
rect 803 1097 804 1101
rect 798 1096 804 1097
rect 951 1099 960 1100
rect 566 1094 573 1095
rect 702 1095 708 1096
rect 534 1091 540 1092
rect 534 1090 535 1091
rect 432 1088 535 1090
rect 287 1086 293 1087
rect 534 1087 535 1088
rect 539 1087 540 1091
rect 702 1091 703 1095
rect 707 1094 708 1095
rect 783 1095 789 1096
rect 783 1094 784 1095
rect 707 1092 784 1094
rect 707 1091 708 1092
rect 702 1090 708 1091
rect 783 1091 784 1092
rect 788 1091 789 1095
rect 927 1095 933 1096
rect 927 1094 928 1095
rect 897 1092 928 1094
rect 783 1090 789 1091
rect 927 1091 928 1092
rect 932 1091 933 1095
rect 951 1095 952 1099
rect 959 1095 960 1099
rect 976 1098 978 1112
rect 983 1111 984 1115
rect 988 1114 989 1115
rect 1014 1115 1015 1119
rect 1020 1115 1021 1119
rect 1030 1119 1031 1123
rect 1035 1119 1036 1123
rect 1030 1118 1036 1119
rect 1062 1123 1068 1124
rect 1062 1119 1063 1123
rect 1067 1119 1068 1123
rect 1094 1120 1095 1124
rect 1099 1120 1100 1124
rect 1094 1119 1100 1120
rect 1134 1123 1140 1124
rect 1134 1119 1135 1123
rect 1139 1119 1140 1123
rect 1166 1120 1167 1124
rect 1171 1120 1172 1124
rect 1246 1124 1247 1128
rect 1251 1124 1252 1128
rect 1334 1126 1340 1127
rect 1246 1123 1252 1124
rect 1286 1123 1292 1124
rect 1166 1119 1172 1120
rect 1286 1119 1287 1123
rect 1291 1119 1292 1123
rect 1334 1122 1335 1126
rect 1339 1122 1340 1126
rect 1334 1121 1340 1122
rect 1422 1123 1428 1124
rect 1062 1118 1068 1119
rect 1134 1118 1140 1119
rect 1286 1118 1292 1119
rect 1422 1119 1423 1123
rect 1427 1119 1428 1123
rect 1422 1118 1428 1119
rect 1454 1123 1460 1124
rect 1454 1119 1455 1123
rect 1459 1119 1460 1123
rect 1454 1118 1460 1119
rect 1486 1123 1492 1124
rect 1486 1119 1487 1123
rect 1491 1119 1492 1123
rect 1486 1118 1492 1119
rect 1518 1123 1524 1124
rect 1518 1119 1519 1123
rect 1523 1119 1524 1123
rect 1518 1118 1524 1119
rect 1558 1123 1564 1124
rect 1558 1119 1559 1123
rect 1563 1119 1564 1123
rect 1558 1118 1564 1119
rect 1590 1123 1596 1124
rect 1590 1119 1591 1123
rect 1595 1119 1596 1123
rect 1590 1118 1596 1119
rect 1622 1123 1628 1124
rect 1622 1119 1623 1123
rect 1627 1119 1628 1123
rect 1622 1118 1628 1119
rect 1654 1123 1660 1124
rect 1654 1119 1655 1123
rect 1659 1119 1660 1123
rect 1654 1118 1660 1119
rect 1694 1121 1700 1122
rect 1694 1117 1695 1121
rect 1699 1117 1700 1121
rect 1694 1116 1700 1117
rect 1014 1114 1021 1115
rect 1047 1115 1053 1116
rect 988 1112 1006 1114
rect 988 1111 989 1112
rect 983 1110 989 1111
rect 1004 1110 1006 1112
rect 1047 1111 1048 1115
rect 1052 1114 1053 1115
rect 1079 1115 1088 1116
rect 1052 1112 1074 1114
rect 1052 1111 1053 1112
rect 1047 1110 1053 1111
rect 1004 1108 1018 1110
rect 998 1101 1004 1102
rect 983 1099 989 1100
rect 983 1098 984 1099
rect 976 1096 984 1098
rect 951 1094 960 1095
rect 983 1095 984 1096
rect 988 1095 989 1099
rect 998 1097 999 1101
rect 1003 1097 1004 1101
rect 998 1096 1004 1097
rect 1016 1098 1018 1108
rect 1030 1106 1036 1107
rect 1030 1102 1031 1106
rect 1035 1102 1036 1106
rect 1030 1101 1036 1102
rect 1062 1106 1068 1107
rect 1062 1102 1063 1106
rect 1067 1102 1068 1106
rect 1062 1101 1068 1102
rect 1047 1099 1053 1100
rect 1047 1098 1048 1099
rect 1016 1096 1048 1098
rect 983 1094 989 1095
rect 1047 1095 1048 1096
rect 1052 1095 1053 1099
rect 1072 1098 1074 1112
rect 1079 1111 1080 1115
rect 1087 1111 1088 1115
rect 1079 1110 1088 1111
rect 1122 1115 1128 1116
rect 1122 1111 1123 1115
rect 1127 1114 1128 1115
rect 1151 1115 1157 1116
rect 1151 1114 1152 1115
rect 1127 1112 1152 1114
rect 1127 1111 1128 1112
rect 1122 1110 1128 1111
rect 1151 1111 1152 1112
rect 1156 1111 1157 1115
rect 1234 1115 1240 1116
rect 1234 1114 1235 1115
rect 1229 1112 1235 1114
rect 1151 1110 1157 1111
rect 1234 1111 1235 1112
rect 1239 1111 1240 1115
rect 1234 1110 1240 1111
rect 1278 1115 1284 1116
rect 1278 1111 1279 1115
rect 1283 1114 1284 1115
rect 1303 1115 1309 1116
rect 1303 1114 1304 1115
rect 1283 1112 1304 1114
rect 1283 1111 1284 1112
rect 1278 1110 1284 1111
rect 1303 1111 1304 1112
rect 1308 1111 1309 1115
rect 1303 1110 1309 1111
rect 1439 1115 1445 1116
rect 1439 1111 1440 1115
rect 1444 1114 1445 1115
rect 1470 1115 1477 1116
rect 1444 1112 1466 1114
rect 1444 1111 1445 1112
rect 1439 1110 1445 1111
rect 1110 1107 1116 1108
rect 1110 1103 1111 1107
rect 1115 1106 1116 1107
rect 1119 1107 1125 1108
rect 1226 1107 1232 1108
rect 1119 1106 1120 1107
rect 1115 1104 1120 1106
rect 1115 1103 1116 1104
rect 1110 1102 1116 1103
rect 1119 1103 1120 1104
rect 1124 1103 1125 1107
rect 1119 1102 1125 1103
rect 1134 1106 1140 1107
rect 1134 1102 1135 1106
rect 1139 1102 1140 1106
rect 1226 1103 1227 1107
rect 1231 1106 1232 1107
rect 1271 1107 1277 1108
rect 1271 1106 1272 1107
rect 1231 1104 1272 1106
rect 1231 1103 1232 1104
rect 1226 1102 1232 1103
rect 1271 1103 1272 1104
rect 1276 1103 1277 1107
rect 1271 1102 1277 1103
rect 1286 1106 1292 1107
rect 1286 1102 1287 1106
rect 1291 1102 1292 1106
rect 1134 1101 1140 1102
rect 1079 1099 1085 1100
rect 1079 1098 1080 1099
rect 1072 1096 1080 1098
rect 1047 1094 1053 1095
rect 1079 1095 1080 1096
rect 1084 1095 1085 1099
rect 1151 1099 1157 1100
rect 1079 1094 1085 1095
rect 1094 1096 1100 1097
rect 1094 1092 1095 1096
rect 1099 1092 1100 1096
rect 1151 1095 1152 1099
rect 1156 1095 1157 1099
rect 1273 1098 1275 1102
rect 1286 1101 1292 1102
rect 1422 1106 1428 1107
rect 1422 1102 1423 1106
rect 1427 1102 1428 1106
rect 1422 1101 1428 1102
rect 1454 1106 1460 1107
rect 1454 1102 1455 1106
rect 1459 1102 1460 1106
rect 1454 1101 1460 1102
rect 1303 1099 1309 1100
rect 1303 1098 1304 1099
rect 1273 1096 1304 1098
rect 1151 1094 1157 1095
rect 1303 1095 1304 1096
rect 1308 1095 1309 1099
rect 1303 1094 1309 1095
rect 1430 1099 1436 1100
rect 1430 1095 1431 1099
rect 1435 1098 1436 1099
rect 1439 1099 1445 1100
rect 1439 1098 1440 1099
rect 1435 1096 1440 1098
rect 1435 1095 1436 1096
rect 1430 1094 1436 1095
rect 1439 1095 1440 1096
rect 1444 1095 1445 1099
rect 1464 1098 1466 1112
rect 1470 1111 1471 1115
rect 1476 1111 1477 1115
rect 1470 1110 1477 1111
rect 1498 1115 1509 1116
rect 1498 1111 1499 1115
rect 1503 1111 1504 1115
rect 1508 1111 1509 1115
rect 1498 1110 1509 1111
rect 1534 1115 1541 1116
rect 1534 1111 1535 1115
rect 1540 1111 1541 1115
rect 1575 1115 1581 1116
rect 1575 1114 1576 1115
rect 1534 1110 1541 1111
rect 1552 1112 1576 1114
rect 1486 1106 1492 1107
rect 1486 1102 1487 1106
rect 1491 1102 1492 1106
rect 1486 1101 1492 1102
rect 1518 1106 1524 1107
rect 1518 1102 1519 1106
rect 1523 1102 1524 1106
rect 1518 1101 1524 1102
rect 1471 1099 1477 1100
rect 1471 1098 1472 1099
rect 1464 1096 1472 1098
rect 1439 1094 1445 1095
rect 1471 1095 1472 1096
rect 1476 1095 1477 1099
rect 1471 1094 1477 1095
rect 1503 1099 1509 1100
rect 1503 1095 1504 1099
rect 1508 1098 1509 1099
rect 1535 1099 1541 1100
rect 1508 1096 1521 1098
rect 1508 1095 1509 1096
rect 1503 1094 1509 1095
rect 1153 1092 1219 1094
rect 1094 1091 1100 1092
rect 927 1090 933 1091
rect 1119 1087 1128 1088
rect 534 1086 540 1087
rect 590 1086 596 1087
rect 79 1083 85 1084
rect 79 1079 80 1083
rect 84 1082 85 1083
rect 306 1083 312 1084
rect 306 1082 307 1083
rect 84 1080 307 1082
rect 84 1079 85 1080
rect 79 1078 85 1079
rect 306 1079 307 1080
rect 311 1079 312 1083
rect 590 1082 591 1086
rect 595 1082 596 1086
rect 590 1081 596 1082
rect 846 1085 852 1086
rect 846 1081 847 1085
rect 851 1081 852 1085
rect 846 1080 852 1081
rect 1071 1083 1077 1084
rect 306 1078 312 1079
rect 790 1079 796 1080
rect 790 1078 791 1079
rect 664 1076 791 1078
rect 190 1075 196 1076
rect 190 1071 191 1075
rect 195 1074 196 1075
rect 583 1075 589 1076
rect 583 1074 584 1075
rect 195 1072 584 1074
rect 195 1071 196 1072
rect 190 1070 196 1071
rect 583 1071 584 1072
rect 588 1074 589 1075
rect 598 1075 605 1076
rect 588 1071 590 1074
rect 583 1070 590 1071
rect 598 1071 599 1075
rect 604 1071 605 1075
rect 598 1070 605 1071
rect 615 1075 621 1076
rect 615 1071 616 1075
rect 620 1074 621 1075
rect 664 1074 666 1076
rect 790 1075 791 1076
rect 795 1075 796 1079
rect 922 1079 928 1080
rect 922 1078 923 1079
rect 919 1077 923 1078
rect 790 1074 796 1075
rect 862 1075 869 1076
rect 620 1072 666 1074
rect 620 1071 621 1072
rect 615 1070 621 1071
rect 822 1071 828 1072
rect 822 1070 823 1071
rect 588 1066 590 1070
rect 741 1068 823 1070
rect 606 1067 612 1068
rect 606 1066 607 1067
rect 588 1064 607 1066
rect 606 1063 607 1064
rect 611 1063 612 1067
rect 822 1067 823 1068
rect 827 1067 828 1071
rect 862 1071 863 1075
rect 868 1074 869 1075
rect 868 1072 914 1074
rect 919 1073 920 1077
rect 927 1075 928 1079
rect 1071 1079 1072 1083
rect 1076 1082 1077 1083
rect 1091 1083 1097 1084
rect 1091 1082 1092 1083
rect 1076 1080 1092 1082
rect 1076 1079 1077 1080
rect 1071 1078 1077 1079
rect 1091 1079 1092 1080
rect 1096 1082 1097 1083
rect 1102 1083 1108 1084
rect 1102 1082 1103 1083
rect 1096 1080 1103 1082
rect 1096 1079 1097 1080
rect 1091 1078 1097 1079
rect 1102 1079 1103 1080
rect 1107 1079 1108 1083
rect 1119 1083 1120 1087
rect 1127 1083 1128 1087
rect 1119 1082 1128 1083
rect 1102 1078 1108 1079
rect 1168 1076 1170 1092
rect 1217 1090 1219 1092
rect 1328 1090 1330 1093
rect 1217 1088 1330 1090
rect 1519 1090 1521 1096
rect 1535 1095 1536 1099
rect 1540 1098 1541 1099
rect 1552 1098 1554 1112
rect 1575 1111 1576 1112
rect 1580 1111 1581 1115
rect 1575 1110 1581 1111
rect 1583 1115 1589 1116
rect 1583 1111 1584 1115
rect 1588 1114 1589 1115
rect 1607 1115 1613 1116
rect 1607 1114 1608 1115
rect 1588 1112 1608 1114
rect 1588 1111 1589 1112
rect 1583 1110 1589 1111
rect 1607 1111 1608 1112
rect 1612 1111 1613 1115
rect 1607 1110 1613 1111
rect 1639 1115 1645 1116
rect 1639 1111 1640 1115
rect 1644 1114 1645 1115
rect 1670 1115 1677 1116
rect 1644 1112 1666 1114
rect 1644 1111 1645 1112
rect 1639 1110 1645 1111
rect 1610 1107 1616 1108
rect 1558 1106 1564 1107
rect 1558 1102 1559 1106
rect 1563 1102 1564 1106
rect 1558 1101 1564 1102
rect 1590 1106 1596 1107
rect 1590 1102 1591 1106
rect 1595 1102 1596 1106
rect 1610 1103 1611 1107
rect 1615 1106 1616 1107
rect 1622 1106 1628 1107
rect 1615 1103 1618 1106
rect 1610 1102 1618 1103
rect 1590 1101 1596 1102
rect 1540 1096 1554 1098
rect 1574 1099 1581 1100
rect 1540 1095 1541 1096
rect 1535 1094 1541 1095
rect 1574 1095 1575 1099
rect 1580 1095 1581 1099
rect 1574 1094 1581 1095
rect 1607 1099 1613 1100
rect 1607 1095 1608 1099
rect 1612 1095 1613 1099
rect 1616 1098 1618 1102
rect 1622 1102 1623 1106
rect 1627 1102 1628 1106
rect 1622 1101 1628 1102
rect 1654 1106 1660 1107
rect 1654 1102 1655 1106
rect 1659 1102 1660 1106
rect 1654 1101 1660 1102
rect 1639 1099 1645 1100
rect 1639 1098 1640 1099
rect 1616 1096 1640 1098
rect 1607 1094 1613 1095
rect 1639 1095 1640 1096
rect 1644 1095 1645 1099
rect 1664 1098 1666 1112
rect 1670 1111 1671 1115
rect 1676 1111 1677 1115
rect 1670 1110 1677 1111
rect 1694 1104 1700 1105
rect 1694 1100 1695 1104
rect 1699 1100 1700 1104
rect 1671 1099 1677 1100
rect 1694 1099 1700 1100
rect 1671 1098 1672 1099
rect 1664 1096 1672 1098
rect 1639 1094 1645 1095
rect 1671 1095 1672 1096
rect 1676 1095 1677 1099
rect 1671 1094 1677 1095
rect 1583 1091 1589 1092
rect 1583 1090 1584 1091
rect 1519 1088 1584 1090
rect 1583 1087 1584 1088
rect 1588 1087 1589 1091
rect 1609 1090 1611 1094
rect 1670 1091 1676 1092
rect 1670 1090 1671 1091
rect 1609 1088 1671 1090
rect 1174 1086 1180 1087
rect 1583 1086 1589 1087
rect 1670 1087 1671 1088
rect 1675 1087 1676 1091
rect 1670 1086 1676 1087
rect 1174 1082 1175 1086
rect 1179 1082 1180 1086
rect 1334 1085 1340 1086
rect 1174 1081 1180 1082
rect 1246 1081 1252 1082
rect 1246 1077 1247 1081
rect 1251 1077 1252 1081
rect 1334 1081 1335 1085
rect 1339 1081 1340 1085
rect 1334 1080 1340 1081
rect 1246 1076 1252 1077
rect 924 1074 928 1075
rect 1167 1075 1173 1076
rect 924 1073 925 1074
rect 919 1072 925 1073
rect 868 1071 869 1072
rect 862 1070 869 1071
rect 912 1070 914 1072
rect 1167 1071 1168 1075
rect 1172 1071 1173 1075
rect 1167 1070 1173 1071
rect 1183 1075 1189 1076
rect 1183 1071 1184 1075
rect 1188 1071 1189 1075
rect 1183 1070 1189 1071
rect 1194 1075 1205 1076
rect 1194 1071 1195 1075
rect 1199 1071 1200 1075
rect 1204 1074 1205 1075
rect 1226 1075 1232 1076
rect 1226 1074 1227 1075
rect 1204 1072 1227 1074
rect 1204 1071 1205 1072
rect 1194 1070 1205 1071
rect 1226 1071 1227 1072
rect 1231 1071 1232 1075
rect 1262 1075 1268 1076
rect 1226 1070 1232 1071
rect 1234 1071 1240 1072
rect 912 1068 922 1070
rect 822 1066 828 1067
rect 920 1066 922 1068
rect 928 1068 1050 1070
rect 928 1066 930 1068
rect 920 1064 930 1066
rect 1048 1066 1050 1068
rect 1185 1066 1187 1070
rect 1234 1067 1235 1071
rect 1239 1070 1240 1071
rect 1243 1071 1249 1072
rect 1243 1070 1244 1071
rect 1239 1068 1244 1070
rect 1239 1067 1240 1068
rect 1234 1066 1240 1067
rect 1243 1067 1244 1068
rect 1248 1067 1249 1071
rect 1262 1071 1263 1075
rect 1267 1074 1268 1075
rect 1271 1075 1277 1076
rect 1271 1074 1272 1075
rect 1267 1072 1272 1074
rect 1267 1071 1268 1072
rect 1262 1070 1268 1071
rect 1271 1071 1272 1072
rect 1276 1071 1277 1075
rect 1271 1070 1277 1071
rect 1350 1075 1357 1076
rect 1350 1071 1351 1075
rect 1356 1071 1357 1075
rect 1350 1070 1357 1071
rect 1407 1075 1413 1076
rect 1407 1071 1408 1075
rect 1412 1074 1413 1075
rect 1446 1075 1452 1076
rect 1446 1074 1447 1075
rect 1412 1072 1447 1074
rect 1412 1071 1413 1072
rect 1407 1070 1413 1071
rect 1446 1071 1447 1072
rect 1451 1071 1452 1075
rect 1446 1070 1452 1071
rect 1243 1066 1249 1067
rect 1048 1064 1187 1066
rect 606 1062 612 1063
rect 1038 1063 1044 1064
rect 1038 1062 1039 1063
rect 749 1060 1039 1062
rect 1038 1059 1039 1060
rect 1043 1059 1044 1063
rect 1038 1058 1044 1059
rect 914 1055 920 1056
rect 914 1054 915 1055
rect 757 1052 915 1054
rect 914 1051 915 1052
rect 919 1051 920 1055
rect 914 1050 920 1051
rect 830 1031 836 1032
rect 830 1030 831 1031
rect 776 1028 831 1030
rect 494 1027 505 1028
rect 398 1023 405 1024
rect 398 1019 399 1023
rect 404 1019 405 1023
rect 398 1018 405 1019
rect 414 1023 421 1024
rect 414 1019 415 1023
rect 420 1019 421 1023
rect 414 1018 421 1019
rect 431 1023 437 1024
rect 431 1019 432 1023
rect 436 1022 437 1023
rect 458 1023 464 1024
rect 458 1022 459 1023
rect 436 1020 459 1022
rect 436 1019 437 1020
rect 431 1018 437 1019
rect 458 1019 459 1020
rect 463 1019 464 1023
rect 494 1023 495 1027
rect 499 1023 500 1027
rect 504 1023 505 1027
rect 494 1022 505 1023
rect 527 1023 533 1024
rect 458 1018 464 1019
rect 502 1019 508 1020
rect 255 1015 261 1016
rect 502 1015 503 1019
rect 507 1015 508 1019
rect 527 1019 528 1023
rect 532 1022 533 1023
rect 542 1023 548 1024
rect 542 1022 543 1023
rect 532 1020 543 1022
rect 532 1019 533 1020
rect 527 1018 533 1019
rect 542 1019 543 1020
rect 547 1019 548 1023
rect 542 1018 548 1019
rect 599 1023 605 1024
rect 599 1019 600 1023
rect 604 1022 605 1023
rect 614 1023 620 1024
rect 614 1022 615 1023
rect 604 1020 615 1022
rect 604 1019 605 1020
rect 599 1018 605 1019
rect 614 1019 615 1020
rect 619 1019 620 1023
rect 614 1018 620 1019
rect 655 1023 664 1024
rect 655 1019 656 1023
rect 663 1019 664 1023
rect 655 1018 664 1019
rect 727 1023 733 1024
rect 727 1019 728 1023
rect 732 1022 733 1023
rect 776 1022 778 1028
rect 830 1027 831 1028
rect 835 1030 836 1031
rect 862 1031 868 1032
rect 862 1030 863 1031
rect 835 1028 863 1030
rect 835 1027 836 1028
rect 830 1026 836 1027
rect 862 1027 863 1028
rect 867 1027 868 1031
rect 862 1026 868 1027
rect 844 1024 858 1026
rect 920 1024 987 1026
rect 732 1020 778 1022
rect 782 1023 789 1024
rect 732 1019 733 1020
rect 727 1018 733 1019
rect 782 1019 783 1023
rect 788 1019 789 1023
rect 844 1020 846 1024
rect 856 1022 866 1024
rect 920 1022 922 1024
rect 864 1020 922 1022
rect 985 1020 987 1024
rect 1014 1023 1020 1024
rect 1014 1022 1015 1023
rect 1003 1021 1015 1022
rect 782 1018 789 1019
rect 815 1019 821 1020
rect 255 1014 256 1015
rect 185 1012 256 1014
rect 153 1000 178 1002
rect 185 1000 187 1012
rect 255 1011 256 1012
rect 260 1011 261 1015
rect 255 1010 261 1011
rect 406 1014 412 1015
rect 502 1014 508 1015
rect 582 1015 588 1016
rect 406 1010 407 1014
rect 411 1010 412 1014
rect 582 1011 583 1015
rect 587 1011 588 1015
rect 582 1010 588 1011
rect 710 1015 716 1016
rect 710 1011 711 1015
rect 715 1011 716 1015
rect 815 1015 816 1019
rect 820 1015 821 1019
rect 815 1014 821 1015
rect 831 1019 837 1020
rect 831 1015 832 1019
rect 836 1018 837 1019
rect 842 1019 848 1020
rect 842 1018 843 1019
rect 836 1016 843 1018
rect 836 1015 837 1016
rect 831 1014 837 1015
rect 842 1015 843 1016
rect 847 1015 848 1019
rect 842 1014 848 1015
rect 851 1019 860 1020
rect 851 1015 852 1019
rect 859 1015 860 1019
rect 851 1014 860 1015
rect 927 1019 933 1020
rect 927 1015 928 1019
rect 932 1018 933 1019
rect 967 1019 973 1020
rect 967 1018 968 1019
rect 932 1016 968 1018
rect 932 1015 933 1016
rect 927 1014 933 1015
rect 967 1015 968 1016
rect 972 1015 973 1019
rect 967 1014 973 1015
rect 983 1019 989 1020
rect 983 1015 984 1019
rect 988 1015 989 1019
rect 1003 1017 1004 1021
rect 1008 1020 1015 1021
rect 1008 1017 1009 1020
rect 1014 1019 1015 1020
rect 1019 1019 1020 1023
rect 1014 1018 1020 1019
rect 1046 1019 1052 1020
rect 1003 1016 1009 1017
rect 983 1014 989 1015
rect 1046 1015 1047 1019
rect 1051 1018 1052 1019
rect 1071 1019 1077 1020
rect 1071 1018 1072 1019
rect 1051 1017 1072 1018
rect 1051 1016 1060 1017
rect 1051 1015 1052 1016
rect 1046 1014 1052 1015
rect 710 1010 716 1011
rect 406 1009 412 1010
rect 246 1007 252 1008
rect 246 1006 247 1007
rect 217 1004 247 1006
rect 217 1000 219 1004
rect 246 1003 247 1004
rect 251 1003 252 1007
rect 246 1002 252 1003
rect 327 1007 333 1008
rect 327 1003 328 1007
rect 332 1006 333 1007
rect 382 1007 388 1008
rect 382 1006 383 1007
rect 332 1004 383 1006
rect 332 1003 333 1004
rect 327 1002 333 1003
rect 382 1003 383 1004
rect 387 1003 388 1007
rect 382 1002 388 1003
rect 574 1007 580 1008
rect 574 1003 575 1007
rect 579 1003 580 1007
rect 817 1006 819 1014
rect 1059 1013 1060 1016
rect 1064 1016 1072 1017
rect 1064 1013 1065 1016
rect 1071 1015 1072 1016
rect 1076 1015 1077 1019
rect 1262 1019 1268 1020
rect 1262 1018 1263 1019
rect 1195 1017 1263 1018
rect 1071 1014 1077 1015
rect 1182 1015 1188 1016
rect 1182 1014 1183 1015
rect 1059 1012 1065 1013
rect 1092 1012 1183 1014
rect 1074 1011 1080 1012
rect 761 1004 819 1006
rect 822 1009 828 1010
rect 822 1005 823 1009
rect 827 1005 828 1009
rect 822 1004 828 1005
rect 974 1009 980 1010
rect 974 1005 975 1009
rect 979 1005 980 1009
rect 1074 1007 1075 1011
rect 1079 1010 1080 1011
rect 1087 1011 1094 1012
rect 1087 1010 1088 1011
rect 1079 1008 1088 1010
rect 1079 1007 1080 1008
rect 1074 1006 1080 1007
rect 1087 1007 1088 1008
rect 1092 1008 1094 1011
rect 1182 1011 1183 1012
rect 1187 1011 1188 1015
rect 1195 1013 1196 1017
rect 1200 1016 1263 1017
rect 1200 1013 1201 1016
rect 1262 1015 1263 1016
rect 1267 1018 1268 1019
rect 1267 1017 1369 1018
rect 1267 1016 1324 1017
rect 1267 1015 1268 1016
rect 1262 1014 1268 1015
rect 1195 1012 1201 1013
rect 1323 1013 1324 1016
rect 1328 1016 1364 1017
rect 1328 1013 1329 1016
rect 1323 1012 1329 1013
rect 1363 1013 1364 1016
rect 1368 1013 1369 1017
rect 1363 1012 1369 1013
rect 1182 1010 1188 1011
rect 1206 1011 1212 1012
rect 1092 1007 1093 1008
rect 1087 1006 1093 1007
rect 1119 1007 1125 1008
rect 974 1004 980 1005
rect 1062 1004 1068 1005
rect 574 1002 580 1003
rect 257 1000 283 1002
rect 1062 1000 1063 1004
rect 1067 1000 1068 1004
rect 1119 1003 1120 1007
rect 1124 1006 1125 1007
rect 1190 1007 1196 1008
rect 1190 1006 1191 1007
rect 1124 1004 1191 1006
rect 1124 1003 1125 1004
rect 1119 1002 1125 1003
rect 1190 1003 1191 1004
rect 1195 1003 1196 1007
rect 1206 1007 1207 1011
rect 1211 1010 1212 1011
rect 1223 1011 1229 1012
rect 1223 1010 1224 1011
rect 1211 1008 1224 1010
rect 1211 1007 1212 1008
rect 1206 1006 1212 1007
rect 1223 1007 1224 1008
rect 1228 1007 1229 1011
rect 1334 1011 1340 1012
rect 1223 1006 1229 1007
rect 1247 1007 1253 1008
rect 1190 1002 1196 1003
rect 1198 1004 1204 1005
rect 1153 1000 1178 1002
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1247 1003 1248 1007
rect 1252 1006 1253 1007
rect 1278 1007 1284 1008
rect 1278 1006 1279 1007
rect 1252 1004 1279 1006
rect 1252 1003 1253 1004
rect 1247 1002 1253 1003
rect 1278 1003 1279 1004
rect 1283 1003 1284 1007
rect 1334 1007 1335 1011
rect 1339 1010 1340 1011
rect 1351 1011 1357 1012
rect 1351 1010 1352 1011
rect 1339 1008 1352 1010
rect 1339 1007 1340 1008
rect 1334 1006 1340 1007
rect 1351 1007 1352 1008
rect 1356 1007 1357 1011
rect 1351 1006 1357 1007
rect 1391 1011 1397 1012
rect 1391 1007 1392 1011
rect 1396 1010 1397 1011
rect 1454 1011 1460 1012
rect 1454 1010 1455 1011
rect 1396 1008 1455 1010
rect 1396 1007 1397 1008
rect 1391 1006 1397 1007
rect 1454 1007 1455 1008
rect 1459 1007 1460 1011
rect 1454 1006 1460 1007
rect 1278 1002 1284 1003
rect 1326 1004 1332 1005
rect 1288 1000 1306 1002
rect 1326 1000 1327 1004
rect 1331 1000 1332 1004
rect 151 999 157 1000
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 151 995 152 999
rect 156 995 157 999
rect 110 991 116 992
rect 134 994 140 995
rect 151 994 157 995
rect 166 994 172 995
rect 134 990 135 994
rect 139 990 140 994
rect 134 989 140 990
rect 166 990 167 994
rect 171 990 172 994
rect 166 989 172 990
rect 150 983 157 984
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 150 979 151 983
rect 156 979 157 983
rect 176 982 178 1000
rect 183 999 189 1000
rect 183 995 184 999
rect 188 995 189 999
rect 215 999 221 1000
rect 215 995 216 999
rect 220 995 221 999
rect 247 999 253 1000
rect 247 998 248 999
rect 240 996 248 998
rect 183 994 189 995
rect 198 994 204 995
rect 215 994 221 995
rect 230 994 236 995
rect 198 990 199 994
rect 203 990 204 994
rect 198 989 204 990
rect 230 990 231 994
rect 235 990 236 994
rect 230 989 236 990
rect 240 984 242 996
rect 247 995 248 996
rect 252 995 253 999
rect 247 994 253 995
rect 183 983 189 984
rect 183 982 184 983
rect 176 980 184 982
rect 150 978 157 979
rect 183 979 184 980
rect 188 979 189 983
rect 183 978 189 979
rect 215 983 221 984
rect 215 979 216 983
rect 220 982 221 983
rect 228 982 242 984
rect 247 983 253 984
rect 220 980 230 982
rect 220 979 221 980
rect 215 978 221 979
rect 247 979 248 983
rect 252 982 253 983
rect 257 982 259 1000
rect 279 999 285 1000
rect 279 995 280 999
rect 284 995 285 999
rect 358 999 365 1000
rect 262 994 268 995
rect 279 994 285 995
rect 326 997 332 998
rect 262 990 263 994
rect 267 990 268 994
rect 326 993 327 997
rect 331 993 332 997
rect 358 995 359 999
rect 364 995 365 999
rect 935 999 941 1000
rect 1062 999 1068 1000
rect 1151 999 1157 1000
rect 358 994 365 995
rect 458 995 464 996
rect 935 995 936 999
rect 940 998 941 999
rect 940 996 962 998
rect 940 995 941 996
rect 326 992 332 993
rect 458 991 459 995
rect 463 994 464 995
rect 918 994 924 995
rect 935 994 941 995
rect 463 992 506 994
rect 463 991 464 992
rect 458 990 464 991
rect 504 990 506 992
rect 527 991 536 992
rect 527 990 528 991
rect 262 989 268 990
rect 504 988 528 990
rect 494 987 500 988
rect 494 986 495 987
rect 461 984 495 986
rect 252 980 259 982
rect 279 983 285 984
rect 252 979 253 980
rect 247 978 253 979
rect 279 979 280 983
rect 284 982 285 983
rect 318 983 324 984
rect 318 982 319 983
rect 284 980 319 982
rect 284 979 285 980
rect 279 978 285 979
rect 318 979 319 980
rect 323 979 324 983
rect 494 983 495 984
rect 499 983 500 987
rect 527 987 528 988
rect 535 987 536 991
rect 918 990 919 994
rect 923 990 924 994
rect 918 989 924 990
rect 960 990 962 996
rect 1118 997 1124 998
rect 1118 993 1119 997
rect 1123 993 1124 997
rect 1151 995 1152 999
rect 1156 995 1157 999
rect 1176 998 1178 1000
rect 1183 999 1189 1000
rect 1198 999 1204 1000
rect 1279 999 1285 1000
rect 1183 998 1184 999
rect 1176 996 1184 998
rect 1183 995 1184 996
rect 1188 995 1189 999
rect 1151 994 1157 995
rect 1166 994 1172 995
rect 1183 994 1189 995
rect 1246 997 1252 998
rect 1118 992 1124 993
rect 1087 991 1093 992
rect 960 988 993 990
rect 527 986 536 987
rect 1087 987 1088 991
rect 1092 990 1093 991
rect 1103 991 1109 992
rect 1103 990 1104 991
rect 1092 988 1104 990
rect 1092 987 1093 988
rect 1087 986 1093 987
rect 1103 987 1104 988
rect 1108 987 1109 991
rect 1166 990 1167 994
rect 1171 990 1172 994
rect 1246 993 1247 997
rect 1251 993 1252 997
rect 1279 995 1280 999
rect 1284 998 1285 999
rect 1288 998 1290 1000
rect 1284 996 1290 998
rect 1304 998 1306 1000
rect 1311 999 1317 1000
rect 1326 999 1332 1000
rect 1366 1004 1372 1005
rect 1366 1000 1367 1004
rect 1371 1000 1372 1004
rect 1543 1003 1549 1004
rect 1366 999 1372 1000
rect 1400 1000 1418 1002
rect 1472 1000 1490 1002
rect 1311 998 1312 999
rect 1304 996 1312 998
rect 1284 995 1285 996
rect 1311 995 1312 996
rect 1316 995 1317 999
rect 1279 994 1285 995
rect 1294 994 1300 995
rect 1311 994 1317 995
rect 1246 992 1252 993
rect 1166 989 1172 990
rect 1223 991 1229 992
rect 1103 986 1109 987
rect 1206 987 1212 988
rect 1206 986 1207 987
rect 1196 984 1207 986
rect 494 982 500 983
rect 934 983 941 984
rect 318 978 324 979
rect 822 979 828 980
rect 110 974 116 975
rect 134 977 140 978
rect 134 973 135 977
rect 139 973 140 977
rect 134 972 140 973
rect 166 977 172 978
rect 166 973 167 977
rect 171 973 172 977
rect 166 972 172 973
rect 198 977 204 978
rect 198 973 199 977
rect 203 973 204 977
rect 198 972 204 973
rect 230 977 236 978
rect 230 973 231 977
rect 235 973 236 977
rect 230 972 236 973
rect 262 977 268 978
rect 262 973 263 977
rect 267 973 268 977
rect 262 972 268 973
rect 398 976 404 977
rect 398 972 399 976
rect 403 972 404 976
rect 822 975 823 979
rect 827 978 828 979
rect 934 979 935 983
rect 940 979 941 983
rect 934 978 941 979
rect 1183 983 1189 984
rect 1183 979 1184 983
rect 1188 982 1189 983
rect 1196 982 1198 984
rect 1206 983 1207 984
rect 1211 983 1212 987
rect 1223 987 1224 991
rect 1228 990 1229 991
rect 1231 991 1237 992
rect 1231 990 1232 991
rect 1228 988 1232 990
rect 1228 987 1229 988
rect 1223 986 1229 987
rect 1231 987 1232 988
rect 1236 987 1237 991
rect 1294 990 1295 994
rect 1299 990 1300 994
rect 1294 989 1300 990
rect 1351 991 1357 992
rect 1231 986 1237 987
rect 1334 987 1340 988
rect 1334 986 1335 987
rect 1324 984 1335 986
rect 1206 982 1212 983
rect 1311 983 1317 984
rect 1188 980 1198 982
rect 1188 979 1189 980
rect 1183 978 1189 979
rect 1311 979 1312 983
rect 1316 982 1317 983
rect 1324 982 1326 984
rect 1334 983 1335 984
rect 1339 983 1340 987
rect 1351 987 1352 991
rect 1356 990 1357 991
rect 1382 991 1388 992
rect 1382 990 1383 991
rect 1356 988 1383 990
rect 1356 987 1357 988
rect 1351 986 1357 987
rect 1382 987 1383 988
rect 1387 987 1388 991
rect 1382 986 1388 987
rect 1391 991 1397 992
rect 1391 987 1392 991
rect 1396 990 1397 991
rect 1400 990 1402 1000
rect 1416 998 1418 1000
rect 1423 999 1429 1000
rect 1423 998 1424 999
rect 1416 996 1424 998
rect 1423 995 1424 996
rect 1428 995 1429 999
rect 1455 999 1461 1000
rect 1455 995 1456 999
rect 1460 998 1461 999
rect 1470 999 1476 1000
rect 1470 998 1471 999
rect 1460 996 1471 998
rect 1460 995 1461 996
rect 1396 988 1402 990
rect 1406 994 1412 995
rect 1423 994 1429 995
rect 1438 994 1444 995
rect 1455 994 1461 995
rect 1470 995 1471 996
rect 1475 995 1476 999
rect 1488 998 1490 1000
rect 1495 999 1501 1000
rect 1495 998 1496 999
rect 1488 996 1496 998
rect 1495 995 1496 996
rect 1500 995 1501 999
rect 1534 999 1541 1000
rect 1534 995 1535 999
rect 1540 995 1541 999
rect 1543 999 1544 1003
rect 1548 1002 1549 1003
rect 1548 1000 1579 1002
rect 1585 1000 1611 1002
rect 1616 1000 1643 1002
rect 1648 1000 1675 1002
rect 1548 999 1549 1000
rect 1543 998 1549 999
rect 1575 999 1581 1000
rect 1575 995 1576 999
rect 1580 995 1581 999
rect 1470 994 1476 995
rect 1478 994 1484 995
rect 1495 994 1501 995
rect 1518 994 1524 995
rect 1534 994 1541 995
rect 1558 994 1564 995
rect 1575 994 1581 995
rect 1406 990 1407 994
rect 1411 990 1412 994
rect 1406 989 1412 990
rect 1438 990 1439 994
rect 1443 990 1444 994
rect 1438 989 1444 990
rect 1478 990 1479 994
rect 1483 990 1484 994
rect 1478 989 1484 990
rect 1518 990 1519 994
rect 1523 990 1524 994
rect 1518 989 1524 990
rect 1558 990 1559 994
rect 1563 990 1564 994
rect 1558 989 1564 990
rect 1396 987 1397 988
rect 1391 986 1397 987
rect 1334 982 1340 983
rect 1423 983 1432 984
rect 1316 980 1326 982
rect 1316 979 1317 980
rect 1311 978 1317 979
rect 1423 979 1424 983
rect 1431 979 1432 983
rect 1423 978 1432 979
rect 1454 983 1461 984
rect 1454 979 1455 983
rect 1460 979 1461 983
rect 1454 978 1461 979
rect 1494 983 1501 984
rect 1494 979 1495 983
rect 1500 979 1501 983
rect 1494 978 1501 979
rect 1535 983 1541 984
rect 1535 979 1536 983
rect 1540 982 1541 983
rect 1543 983 1549 984
rect 1543 982 1544 983
rect 1540 980 1544 982
rect 1540 979 1541 980
rect 1535 978 1541 979
rect 1543 979 1544 980
rect 1548 979 1549 983
rect 1543 978 1549 979
rect 1575 983 1581 984
rect 1575 979 1576 983
rect 1580 982 1581 983
rect 1585 982 1587 1000
rect 1607 999 1613 1000
rect 1607 995 1608 999
rect 1612 995 1613 999
rect 1590 994 1596 995
rect 1607 994 1613 995
rect 1590 990 1591 994
rect 1595 990 1596 994
rect 1590 989 1596 990
rect 1580 980 1587 982
rect 1607 983 1613 984
rect 1580 979 1581 980
rect 1575 978 1581 979
rect 1607 979 1608 983
rect 1612 982 1613 983
rect 1616 982 1618 1000
rect 1639 999 1645 1000
rect 1639 995 1640 999
rect 1644 995 1645 999
rect 1622 994 1628 995
rect 1639 994 1645 995
rect 1622 990 1623 994
rect 1627 990 1628 994
rect 1622 989 1628 990
rect 1612 980 1618 982
rect 1639 983 1645 984
rect 1612 979 1613 980
rect 1607 978 1613 979
rect 1639 979 1640 983
rect 1644 982 1645 983
rect 1648 982 1650 1000
rect 1671 999 1677 1000
rect 1671 995 1672 999
rect 1676 995 1677 999
rect 1654 994 1660 995
rect 1671 994 1677 995
rect 1694 996 1700 997
rect 1654 990 1655 994
rect 1659 990 1660 994
rect 1694 992 1695 996
rect 1699 992 1700 996
rect 1694 991 1700 992
rect 1654 989 1660 990
rect 1644 980 1650 982
rect 1671 983 1677 984
rect 1644 979 1645 980
rect 1639 978 1645 979
rect 1671 979 1672 983
rect 1676 979 1677 983
rect 1671 978 1677 979
rect 1694 979 1700 980
rect 827 976 833 978
rect 918 977 924 978
rect 1166 977 1172 978
rect 1294 977 1300 978
rect 1406 977 1412 978
rect 827 975 828 976
rect 582 974 588 975
rect 398 971 404 972
rect 502 972 508 973
rect 342 970 348 971
rect 342 966 343 970
rect 347 966 348 970
rect 502 968 503 972
rect 507 968 508 972
rect 582 970 583 974
rect 587 970 588 974
rect 582 969 588 970
rect 710 974 716 975
rect 822 974 828 975
rect 710 970 711 974
rect 715 970 716 974
rect 918 973 919 977
rect 923 973 924 977
rect 918 972 924 973
rect 1062 976 1068 977
rect 1062 972 1063 976
rect 1067 972 1068 976
rect 1166 973 1167 977
rect 1171 973 1172 977
rect 1166 972 1172 973
rect 1198 976 1204 977
rect 1198 972 1199 976
rect 1203 972 1204 976
rect 1294 973 1295 977
rect 1299 973 1300 977
rect 1294 972 1300 973
rect 1326 976 1332 977
rect 1326 972 1327 976
rect 1331 972 1332 976
rect 1062 971 1068 972
rect 1198 971 1204 972
rect 1326 971 1332 972
rect 1366 976 1372 977
rect 1366 972 1367 976
rect 1371 972 1372 976
rect 1406 973 1407 977
rect 1411 973 1412 977
rect 1406 972 1412 973
rect 1438 977 1444 978
rect 1438 973 1439 977
rect 1443 973 1444 977
rect 1438 972 1444 973
rect 1478 977 1484 978
rect 1478 973 1479 977
rect 1483 973 1484 977
rect 1478 972 1484 973
rect 1518 977 1524 978
rect 1518 973 1519 977
rect 1523 973 1524 977
rect 1518 972 1524 973
rect 1558 977 1564 978
rect 1558 973 1559 977
rect 1563 973 1564 977
rect 1558 972 1564 973
rect 1590 977 1596 978
rect 1590 973 1591 977
rect 1595 973 1596 977
rect 1590 972 1596 973
rect 1622 977 1628 978
rect 1622 973 1623 977
rect 1627 973 1628 977
rect 1622 972 1628 973
rect 1654 977 1660 978
rect 1654 973 1655 977
rect 1659 973 1660 977
rect 1654 972 1660 973
rect 1366 971 1372 972
rect 1538 971 1544 972
rect 1134 970 1140 971
rect 710 969 716 970
rect 814 969 820 970
rect 502 967 508 968
rect 342 965 348 966
rect 814 965 815 969
rect 819 965 820 969
rect 814 964 820 965
rect 966 969 972 970
rect 966 965 967 969
rect 971 965 972 969
rect 1134 966 1135 970
rect 1139 966 1140 970
rect 1134 965 1140 966
rect 1262 970 1268 971
rect 1262 966 1263 970
rect 1267 966 1268 970
rect 1538 967 1539 971
rect 1543 970 1544 971
rect 1673 970 1675 978
rect 1694 975 1695 979
rect 1699 975 1700 979
rect 1694 974 1700 975
rect 1543 968 1675 970
rect 1543 967 1544 968
rect 1538 966 1544 967
rect 1262 965 1268 966
rect 966 964 972 965
rect 318 963 325 964
rect 318 959 319 963
rect 324 959 325 963
rect 318 958 325 959
rect 1082 963 1088 964
rect 1082 959 1083 963
rect 1087 962 1088 963
rect 1111 963 1117 964
rect 1111 962 1112 963
rect 1087 960 1112 962
rect 1087 959 1088 960
rect 1082 958 1088 959
rect 1111 959 1112 960
rect 1116 962 1117 963
rect 1239 963 1245 964
rect 1239 962 1240 963
rect 1116 960 1240 962
rect 1116 959 1117 960
rect 1111 958 1117 959
rect 1239 959 1240 960
rect 1244 959 1245 963
rect 1239 958 1245 959
rect 218 955 224 956
rect 218 951 219 955
rect 223 954 224 955
rect 598 955 604 956
rect 598 954 599 955
rect 223 952 599 954
rect 223 951 224 952
rect 218 950 224 951
rect 598 951 599 952
rect 603 951 604 955
rect 598 950 604 951
rect 658 955 664 956
rect 658 951 659 955
rect 663 954 664 955
rect 854 955 860 956
rect 854 954 855 955
rect 663 952 855 954
rect 663 951 664 952
rect 658 950 664 951
rect 854 951 855 952
rect 859 951 860 955
rect 854 950 860 951
rect 1323 947 1329 948
rect 1195 945 1201 946
rect 1195 944 1196 945
rect 338 943 344 944
rect 338 939 339 943
rect 343 942 344 943
rect 414 943 420 944
rect 414 942 415 943
rect 343 940 415 942
rect 343 939 344 940
rect 338 938 344 939
rect 414 939 415 940
rect 419 939 420 943
rect 414 938 420 939
rect 1194 943 1196 944
rect 1194 939 1195 943
rect 1200 941 1201 945
rect 1323 943 1324 947
rect 1328 946 1329 947
rect 1398 947 1404 948
rect 1398 946 1399 947
rect 1328 944 1399 946
rect 1328 943 1329 944
rect 1323 942 1329 943
rect 1398 943 1399 944
rect 1403 943 1404 947
rect 1398 942 1404 943
rect 1199 940 1201 941
rect 1199 939 1200 940
rect 1194 938 1200 939
rect 1122 935 1128 936
rect 990 931 996 932
rect 278 928 284 929
rect 198 924 204 925
rect 134 923 140 924
rect 110 921 116 922
rect 110 917 111 921
rect 115 917 116 921
rect 134 919 135 923
rect 139 919 140 923
rect 134 918 140 919
rect 166 923 172 924
rect 166 919 167 923
rect 171 919 172 923
rect 198 920 199 924
rect 203 920 204 924
rect 278 924 279 928
rect 283 924 284 928
rect 398 928 404 929
rect 278 923 284 924
rect 318 924 324 925
rect 198 919 204 920
rect 318 920 319 924
rect 323 920 324 924
rect 398 924 399 928
rect 403 924 404 928
rect 990 927 991 931
rect 995 930 996 931
rect 1122 931 1123 935
rect 1127 934 1128 935
rect 1367 935 1373 936
rect 1367 934 1368 935
rect 1127 932 1368 934
rect 1127 931 1128 932
rect 1122 930 1128 931
rect 1367 931 1368 932
rect 1372 931 1373 935
rect 1367 930 1373 931
rect 1390 930 1396 931
rect 995 928 1106 930
rect 995 927 996 928
rect 398 923 404 924
rect 590 926 596 927
rect 590 922 591 926
rect 595 922 596 926
rect 726 926 732 927
rect 590 921 596 922
rect 678 924 684 925
rect 318 919 324 920
rect 462 920 468 921
rect 678 920 679 924
rect 683 920 684 924
rect 726 922 727 926
rect 731 922 732 926
rect 862 926 868 927
rect 990 926 996 927
rect 726 921 732 922
rect 814 923 820 924
rect 166 918 172 919
rect 110 916 116 917
rect 462 916 463 920
rect 467 916 468 920
rect 151 915 157 916
rect 151 911 152 915
rect 156 914 157 915
rect 159 915 165 916
rect 159 914 160 915
rect 156 912 160 914
rect 156 911 157 912
rect 151 910 157 911
rect 159 911 160 912
rect 164 911 165 915
rect 159 910 165 911
rect 183 915 192 916
rect 183 911 184 915
rect 191 911 192 915
rect 266 915 272 916
rect 266 914 267 915
rect 261 912 267 914
rect 183 910 192 911
rect 266 911 267 912
rect 271 911 272 915
rect 386 915 392 916
rect 462 915 468 916
rect 559 919 565 920
rect 559 915 560 919
rect 564 918 565 919
rect 598 919 604 920
rect 678 919 684 920
rect 694 919 701 920
rect 598 918 599 919
rect 564 916 599 918
rect 564 915 565 916
rect 386 914 387 915
rect 381 912 387 914
rect 266 910 272 911
rect 386 911 387 912
rect 391 911 392 915
rect 559 914 565 915
rect 598 915 599 916
rect 603 915 604 919
rect 598 914 604 915
rect 694 915 695 919
rect 700 915 701 919
rect 814 919 815 923
rect 819 919 820 923
rect 862 922 863 926
rect 867 922 868 926
rect 982 924 988 925
rect 1070 924 1076 925
rect 862 921 868 922
rect 950 923 956 924
rect 814 918 820 919
rect 950 919 951 923
rect 955 919 956 923
rect 982 920 983 924
rect 987 920 988 924
rect 982 919 988 920
rect 1038 923 1044 924
rect 1038 919 1039 923
rect 1043 919 1044 923
rect 1070 920 1071 924
rect 1075 920 1076 924
rect 1070 919 1076 920
rect 950 918 956 919
rect 1038 918 1044 919
rect 694 914 701 915
rect 802 915 808 916
rect 386 910 392 911
rect 802 911 803 915
rect 807 914 808 915
rect 831 915 837 916
rect 831 914 832 915
rect 807 912 832 914
rect 807 911 808 912
rect 802 910 808 911
rect 831 911 832 912
rect 836 911 837 915
rect 831 910 837 911
rect 967 915 976 916
rect 967 911 968 915
rect 975 911 976 915
rect 967 910 976 911
rect 1055 915 1061 916
rect 1055 911 1056 915
rect 1060 914 1061 915
rect 1094 915 1100 916
rect 1094 914 1095 915
rect 1060 912 1095 914
rect 1060 911 1061 912
rect 1055 910 1061 911
rect 1094 911 1095 912
rect 1099 911 1100 915
rect 1104 914 1106 928
rect 1390 926 1391 930
rect 1395 926 1396 930
rect 1390 925 1396 926
rect 1142 924 1148 925
rect 1270 924 1276 925
rect 1454 924 1460 925
rect 1110 923 1116 924
rect 1110 919 1111 923
rect 1115 919 1116 923
rect 1142 920 1143 924
rect 1147 920 1148 924
rect 1142 919 1148 920
rect 1238 923 1244 924
rect 1238 919 1239 923
rect 1243 919 1244 923
rect 1270 920 1271 924
rect 1275 920 1276 924
rect 1270 919 1276 920
rect 1422 923 1428 924
rect 1422 919 1423 923
rect 1427 919 1428 923
rect 1454 920 1455 924
rect 1459 920 1460 924
rect 1454 919 1460 920
rect 1518 923 1524 924
rect 1518 919 1519 923
rect 1523 919 1524 923
rect 1110 918 1116 919
rect 1238 918 1244 919
rect 1422 918 1428 919
rect 1518 918 1524 919
rect 1558 923 1564 924
rect 1558 919 1559 923
rect 1563 919 1564 923
rect 1558 918 1564 919
rect 1590 923 1596 924
rect 1590 919 1591 923
rect 1595 919 1596 923
rect 1590 918 1596 919
rect 1622 923 1628 924
rect 1622 919 1623 923
rect 1627 919 1628 923
rect 1622 918 1628 919
rect 1654 923 1660 924
rect 1654 919 1655 923
rect 1659 919 1660 923
rect 1654 918 1660 919
rect 1694 921 1700 922
rect 1694 917 1695 921
rect 1699 917 1700 921
rect 1694 916 1700 917
rect 1127 915 1133 916
rect 1127 914 1128 915
rect 1104 912 1128 914
rect 1094 910 1100 911
rect 1127 911 1128 912
rect 1132 911 1133 915
rect 1230 915 1236 916
rect 1127 910 1133 911
rect 1136 912 1185 914
rect 258 907 264 908
rect 134 906 140 907
rect 110 904 116 905
rect 110 900 111 904
rect 115 900 116 904
rect 134 902 135 906
rect 139 902 140 906
rect 134 901 140 902
rect 166 906 172 907
rect 166 902 167 906
rect 171 902 172 906
rect 258 903 259 907
rect 263 906 264 907
rect 303 907 309 908
rect 303 906 304 907
rect 263 904 304 906
rect 263 903 264 904
rect 258 902 264 903
rect 303 903 304 904
rect 308 903 309 907
rect 303 902 309 903
rect 423 907 432 908
rect 1095 907 1101 908
rect 423 903 424 907
rect 431 903 432 907
rect 814 906 820 907
rect 423 902 432 903
rect 434 905 440 906
rect 166 901 172 902
rect 434 901 435 905
rect 439 901 440 905
rect 814 902 815 906
rect 819 902 820 906
rect 434 900 440 901
rect 678 901 684 902
rect 814 901 820 902
rect 950 906 956 907
rect 950 902 951 906
rect 955 902 956 906
rect 1038 906 1044 907
rect 950 901 956 902
rect 998 903 1004 904
rect 110 899 116 900
rect 150 899 157 900
rect 150 895 151 899
rect 156 895 157 899
rect 150 894 157 895
rect 182 899 189 900
rect 182 895 183 899
rect 188 895 189 899
rect 678 897 679 901
rect 683 897 684 901
rect 678 896 684 897
rect 822 899 828 900
rect 182 894 189 895
rect 522 895 528 896
rect 522 891 523 895
rect 527 894 528 895
rect 559 895 565 896
rect 559 894 560 895
rect 527 892 560 894
rect 527 891 528 892
rect 522 890 528 891
rect 559 891 560 892
rect 564 891 565 895
rect 559 890 565 891
rect 606 895 612 896
rect 606 891 607 895
rect 611 891 612 895
rect 822 895 823 899
rect 827 898 828 899
rect 831 899 837 900
rect 831 898 832 899
rect 827 896 832 898
rect 827 895 828 896
rect 822 894 828 895
rect 831 895 832 896
rect 836 895 837 899
rect 967 899 973 900
rect 831 894 837 895
rect 854 895 860 896
rect 606 890 612 891
rect 854 891 855 895
rect 859 891 860 895
rect 967 895 968 899
rect 972 898 973 899
rect 990 899 996 900
rect 990 898 991 899
rect 972 896 991 898
rect 972 895 973 896
rect 967 894 973 895
rect 990 895 991 896
rect 995 895 996 899
rect 998 899 999 903
rect 1003 899 1004 903
rect 998 898 1004 899
rect 1019 903 1025 904
rect 1019 899 1020 903
rect 1024 902 1025 903
rect 1038 902 1039 906
rect 1043 902 1044 906
rect 1095 903 1096 907
rect 1100 906 1101 907
rect 1100 904 1106 906
rect 1100 903 1101 904
rect 1095 902 1101 903
rect 1024 900 1034 902
rect 1038 901 1044 902
rect 1024 899 1025 900
rect 1019 898 1025 899
rect 1032 898 1034 900
rect 1055 899 1061 900
rect 1055 898 1056 899
rect 1032 896 1056 898
rect 990 894 996 895
rect 1055 895 1056 896
rect 1060 895 1061 899
rect 1055 894 1061 895
rect 1070 896 1076 897
rect 1070 892 1071 896
rect 1075 892 1076 896
rect 1070 891 1076 892
rect 854 890 860 891
rect 1104 890 1106 904
rect 1110 905 1116 906
rect 1110 901 1111 905
rect 1115 901 1116 905
rect 1110 900 1116 901
rect 1127 899 1133 900
rect 1127 895 1128 899
rect 1132 898 1133 899
rect 1136 898 1138 912
rect 1230 911 1231 915
rect 1235 914 1236 915
rect 1255 915 1261 916
rect 1255 914 1256 915
rect 1235 912 1256 914
rect 1235 911 1236 912
rect 1230 910 1236 911
rect 1255 911 1256 912
rect 1260 911 1261 915
rect 1439 915 1445 916
rect 1439 914 1440 915
rect 1255 910 1261 911
rect 1264 912 1313 914
rect 1412 912 1440 914
rect 1142 905 1148 906
rect 1142 901 1143 905
rect 1147 901 1148 905
rect 1142 900 1148 901
rect 1238 905 1244 906
rect 1238 901 1239 905
rect 1243 901 1244 905
rect 1238 900 1244 901
rect 1206 899 1212 900
rect 1206 898 1207 899
rect 1132 896 1138 898
rect 1159 896 1207 898
rect 1132 895 1133 896
rect 1127 894 1133 895
rect 1159 890 1161 896
rect 1206 895 1207 896
rect 1211 895 1212 899
rect 1206 894 1212 895
rect 1255 899 1261 900
rect 1255 895 1256 899
rect 1260 898 1261 899
rect 1264 898 1266 912
rect 1354 911 1360 912
rect 1354 907 1355 911
rect 1359 910 1360 911
rect 1412 910 1414 912
rect 1439 911 1440 912
rect 1444 911 1445 915
rect 1439 910 1445 911
rect 1535 915 1541 916
rect 1535 911 1536 915
rect 1540 914 1541 915
rect 1575 915 1581 916
rect 1540 912 1570 914
rect 1540 911 1541 912
rect 1535 910 1541 911
rect 1359 908 1414 910
rect 1359 907 1360 908
rect 1354 906 1360 907
rect 1422 906 1428 907
rect 1270 905 1276 906
rect 1270 901 1271 905
rect 1275 901 1276 905
rect 1270 900 1276 901
rect 1374 903 1380 904
rect 1374 899 1375 903
rect 1379 899 1380 903
rect 1422 902 1423 906
rect 1427 902 1428 906
rect 1518 906 1524 907
rect 1422 901 1428 902
rect 1470 903 1476 904
rect 1374 898 1380 899
rect 1398 899 1404 900
rect 1260 896 1266 898
rect 1260 895 1261 896
rect 1255 894 1261 895
rect 1398 895 1399 899
rect 1403 898 1404 899
rect 1407 899 1413 900
rect 1407 898 1408 899
rect 1403 896 1408 898
rect 1403 895 1404 896
rect 1398 894 1404 895
rect 1407 895 1408 896
rect 1412 895 1413 899
rect 1407 894 1413 895
rect 1430 899 1436 900
rect 1430 895 1431 899
rect 1435 898 1436 899
rect 1439 899 1445 900
rect 1439 898 1440 899
rect 1435 896 1440 898
rect 1435 895 1436 896
rect 1430 894 1436 895
rect 1439 895 1440 896
rect 1444 895 1445 899
rect 1470 899 1471 903
rect 1475 899 1476 903
rect 1491 903 1497 904
rect 1491 902 1492 903
rect 1470 898 1476 899
rect 1480 900 1492 902
rect 1439 894 1445 895
rect 1480 894 1482 900
rect 1491 899 1492 900
rect 1496 899 1497 903
rect 1518 902 1519 906
rect 1523 902 1524 906
rect 1518 901 1524 902
rect 1558 906 1564 907
rect 1558 902 1559 906
rect 1563 902 1564 906
rect 1558 901 1564 902
rect 1491 898 1497 899
rect 1535 899 1544 900
rect 1535 895 1536 899
rect 1543 895 1544 899
rect 1568 898 1570 912
rect 1575 911 1576 915
rect 1580 914 1581 915
rect 1607 915 1613 916
rect 1580 912 1602 914
rect 1580 911 1581 912
rect 1575 910 1581 911
rect 1590 906 1596 907
rect 1590 902 1591 906
rect 1595 902 1596 906
rect 1590 901 1596 902
rect 1575 899 1581 900
rect 1575 898 1576 899
rect 1568 896 1576 898
rect 1535 894 1544 895
rect 1575 895 1576 896
rect 1580 895 1581 899
rect 1600 898 1602 912
rect 1607 911 1608 915
rect 1612 914 1613 915
rect 1639 915 1645 916
rect 1612 912 1634 914
rect 1612 911 1613 912
rect 1607 910 1613 911
rect 1622 906 1628 907
rect 1622 902 1623 906
rect 1627 902 1628 906
rect 1622 901 1628 902
rect 1607 899 1613 900
rect 1607 898 1608 899
rect 1600 896 1608 898
rect 1575 894 1581 895
rect 1607 895 1608 896
rect 1612 895 1613 899
rect 1632 898 1634 912
rect 1639 911 1640 915
rect 1644 914 1645 915
rect 1670 915 1677 916
rect 1644 912 1666 914
rect 1644 911 1645 912
rect 1639 910 1645 911
rect 1654 906 1660 907
rect 1654 902 1655 906
rect 1659 902 1660 906
rect 1654 901 1660 902
rect 1639 899 1645 900
rect 1639 898 1640 899
rect 1632 896 1640 898
rect 1607 894 1613 895
rect 1639 895 1640 896
rect 1644 895 1645 899
rect 1664 898 1666 912
rect 1670 911 1671 915
rect 1676 911 1677 915
rect 1670 910 1677 911
rect 1694 904 1700 905
rect 1694 900 1695 904
rect 1699 900 1700 904
rect 1671 899 1677 900
rect 1694 899 1700 900
rect 1671 898 1672 899
rect 1664 896 1672 898
rect 1639 894 1645 895
rect 1671 895 1672 896
rect 1676 895 1677 899
rect 1671 894 1677 895
rect 1460 892 1482 894
rect 1354 891 1360 892
rect 1104 888 1161 890
rect 1200 888 1219 890
rect 1003 887 1009 888
rect 206 886 212 887
rect 206 882 207 886
rect 211 882 212 886
rect 326 886 332 887
rect 326 882 327 886
rect 331 882 332 886
rect 590 885 596 886
rect 206 881 212 882
rect 278 881 284 882
rect 326 881 332 882
rect 398 881 404 882
rect 278 877 279 881
rect 283 877 284 881
rect 278 876 284 877
rect 398 877 399 881
rect 403 877 404 881
rect 590 881 591 885
rect 595 881 596 885
rect 590 880 596 881
rect 726 885 732 886
rect 726 881 727 885
rect 731 881 732 885
rect 726 880 732 881
rect 862 885 868 886
rect 862 881 863 885
rect 867 881 868 885
rect 862 880 868 881
rect 970 883 976 884
rect 542 879 548 880
rect 542 878 543 879
rect 398 876 404 877
rect 425 876 543 878
rect 87 875 93 876
rect 87 871 88 875
rect 92 874 93 875
rect 199 875 205 876
rect 199 874 200 875
rect 92 872 200 874
rect 92 871 93 872
rect 87 870 93 871
rect 199 871 200 872
rect 204 874 205 875
rect 207 875 213 876
rect 207 874 208 875
rect 204 872 208 874
rect 204 871 205 872
rect 199 870 205 871
rect 207 871 208 872
rect 212 871 213 875
rect 207 870 213 871
rect 215 875 224 876
rect 215 871 216 875
rect 223 871 224 875
rect 215 870 224 871
rect 231 875 237 876
rect 231 871 232 875
rect 236 874 237 875
rect 258 875 264 876
rect 258 874 259 875
rect 236 872 259 874
rect 236 871 237 872
rect 231 870 237 871
rect 258 871 259 872
rect 263 871 264 875
rect 303 875 312 876
rect 258 870 264 871
rect 266 871 272 872
rect 266 867 267 871
rect 271 870 272 871
rect 275 871 281 872
rect 275 870 276 871
rect 271 868 276 870
rect 271 867 272 868
rect 266 866 272 867
rect 275 867 276 868
rect 280 867 281 871
rect 303 871 304 875
rect 311 871 312 875
rect 303 870 312 871
rect 319 875 325 876
rect 319 871 320 875
rect 324 871 325 875
rect 319 870 325 871
rect 335 875 344 876
rect 335 871 336 875
rect 343 871 344 875
rect 335 870 344 871
rect 351 875 357 876
rect 351 871 352 875
rect 356 874 357 875
rect 414 875 420 876
rect 356 872 382 874
rect 356 871 357 872
rect 351 870 357 871
rect 275 866 281 867
rect 258 863 264 864
rect 258 859 259 863
rect 263 862 264 863
rect 319 862 321 870
rect 263 860 321 862
rect 380 862 382 872
rect 386 871 392 872
rect 386 867 387 871
rect 391 870 392 871
rect 395 871 401 872
rect 395 870 396 871
rect 391 868 396 870
rect 391 867 392 868
rect 386 866 392 867
rect 395 867 396 868
rect 400 867 401 871
rect 414 871 415 875
rect 419 874 420 875
rect 423 875 429 876
rect 423 874 424 875
rect 419 872 424 874
rect 419 871 420 872
rect 414 870 420 871
rect 423 871 424 872
rect 428 871 429 875
rect 542 875 543 876
rect 547 875 548 879
rect 970 879 971 883
rect 975 882 976 883
rect 979 883 985 884
rect 979 882 980 883
rect 975 880 980 882
rect 975 879 976 880
rect 970 878 976 879
rect 979 879 980 880
rect 984 879 985 883
rect 1003 883 1004 887
rect 1008 886 1009 887
rect 1046 887 1052 888
rect 1046 886 1047 887
rect 1008 884 1047 886
rect 1008 883 1009 884
rect 1003 882 1009 883
rect 1046 883 1047 884
rect 1051 886 1052 887
rect 1078 887 1084 888
rect 1078 886 1079 887
rect 1051 885 1079 886
rect 1051 884 1068 885
rect 1051 883 1052 884
rect 1046 882 1052 883
rect 1067 881 1068 884
rect 1072 884 1079 885
rect 1072 881 1073 884
rect 1078 883 1079 884
rect 1083 883 1084 887
rect 1078 882 1084 883
rect 1094 887 1101 888
rect 1094 883 1095 887
rect 1100 883 1101 887
rect 1179 887 1185 888
rect 1179 886 1180 887
rect 1159 884 1180 886
rect 1094 882 1101 883
rect 1103 883 1109 884
rect 1067 880 1073 881
rect 979 878 985 879
rect 1103 879 1104 883
rect 1108 882 1109 883
rect 1159 882 1161 884
rect 1179 883 1180 884
rect 1184 886 1185 887
rect 1200 886 1202 888
rect 1184 884 1202 886
rect 1217 886 1219 888
rect 1307 887 1313 888
rect 1307 886 1308 887
rect 1217 884 1308 886
rect 1184 883 1185 884
rect 1179 882 1185 883
rect 1206 883 1213 884
rect 1108 880 1161 882
rect 1108 879 1109 880
rect 1103 878 1109 879
rect 1206 879 1207 883
rect 1212 879 1213 883
rect 1307 883 1308 884
rect 1312 883 1313 887
rect 1354 887 1355 891
rect 1359 890 1360 891
rect 1375 891 1381 892
rect 1375 890 1376 891
rect 1359 888 1376 890
rect 1359 887 1360 888
rect 1354 886 1360 887
rect 1375 887 1376 888
rect 1380 887 1381 891
rect 1375 886 1381 887
rect 1414 891 1420 892
rect 1414 887 1415 891
rect 1419 890 1420 891
rect 1460 890 1462 892
rect 1419 888 1462 890
rect 1419 887 1420 888
rect 1414 886 1420 887
rect 1475 887 1484 888
rect 1307 882 1313 883
rect 1335 883 1341 884
rect 1335 882 1336 883
rect 1316 880 1336 882
rect 1206 878 1213 879
rect 1231 879 1237 880
rect 542 874 548 875
rect 607 875 613 876
rect 423 870 429 871
rect 607 871 608 875
rect 612 871 613 875
rect 607 870 613 871
rect 663 875 669 876
rect 663 871 664 875
rect 668 874 669 875
rect 711 875 717 876
rect 711 874 712 875
rect 668 872 712 874
rect 668 871 669 872
rect 663 870 669 871
rect 711 871 712 872
rect 716 871 717 875
rect 711 870 717 871
rect 743 875 749 876
rect 743 871 744 875
rect 748 874 749 875
rect 799 875 808 876
rect 748 871 750 874
rect 743 870 750 871
rect 799 871 800 875
rect 807 871 808 875
rect 879 875 885 876
rect 879 874 880 875
rect 799 870 808 871
rect 812 872 880 874
rect 517 868 578 870
rect 748 868 750 870
rect 395 866 401 867
rect 576 866 578 868
rect 702 867 708 868
rect 702 866 703 867
rect 576 864 703 866
rect 426 863 432 864
rect 426 862 427 863
rect 380 860 427 862
rect 263 859 264 860
rect 258 858 264 859
rect 426 859 427 860
rect 431 862 432 863
rect 702 863 703 864
rect 707 863 708 867
rect 702 862 708 863
rect 746 867 752 868
rect 746 863 747 867
rect 751 866 752 867
rect 812 866 814 872
rect 879 871 880 872
rect 884 871 885 875
rect 879 870 885 871
rect 934 875 941 876
rect 934 871 935 875
rect 940 871 941 875
rect 1231 875 1232 879
rect 1236 878 1237 879
rect 1316 878 1318 880
rect 1335 879 1336 880
rect 1340 879 1341 883
rect 1335 878 1341 879
rect 1382 883 1388 884
rect 1382 879 1383 883
rect 1387 882 1388 883
rect 1451 883 1457 884
rect 1451 882 1452 883
rect 1387 880 1452 882
rect 1387 879 1388 880
rect 1382 878 1388 879
rect 1451 879 1452 880
rect 1456 879 1457 883
rect 1475 883 1476 887
rect 1483 883 1484 887
rect 1475 882 1484 883
rect 1662 883 1668 884
rect 1451 878 1457 879
rect 1662 879 1663 883
rect 1667 882 1668 883
rect 1747 883 1753 884
rect 1747 882 1748 883
rect 1667 880 1748 882
rect 1667 879 1668 880
rect 1662 878 1668 879
rect 1747 879 1748 880
rect 1752 879 1753 883
rect 1747 878 1753 879
rect 1236 876 1318 878
rect 1236 875 1237 876
rect 1231 874 1237 875
rect 934 870 941 871
rect 751 864 814 866
rect 751 863 752 864
rect 746 862 752 863
rect 431 860 453 862
rect 431 859 432 860
rect 426 858 432 859
rect 598 859 604 860
rect 306 855 312 856
rect 306 851 307 855
rect 311 854 312 855
rect 414 855 420 856
rect 414 854 415 855
rect 311 852 415 854
rect 311 851 312 852
rect 306 850 312 851
rect 414 851 415 852
rect 419 851 420 855
rect 414 850 420 851
rect 530 855 536 856
rect 530 851 531 855
rect 535 851 536 855
rect 598 855 599 859
rect 603 858 604 859
rect 886 859 892 860
rect 886 858 887 859
rect 603 856 887 858
rect 603 855 604 856
rect 598 854 604 855
rect 886 855 887 856
rect 891 855 892 859
rect 886 854 892 855
rect 530 850 536 851
rect 679 843 685 844
rect 302 839 308 840
rect 302 838 303 839
rect 249 836 303 838
rect 249 832 251 836
rect 302 835 303 836
rect 307 838 308 839
rect 358 839 364 840
rect 358 838 359 839
rect 307 836 359 838
rect 307 835 308 836
rect 302 834 308 835
rect 358 835 359 836
rect 363 838 364 839
rect 606 839 612 840
rect 606 838 607 839
rect 363 836 607 838
rect 363 835 364 836
rect 358 834 364 835
rect 606 835 607 836
rect 611 835 612 839
rect 679 839 680 843
rect 684 842 685 843
rect 850 843 856 844
rect 850 842 851 843
rect 684 840 851 842
rect 684 839 685 840
rect 679 838 685 839
rect 850 839 851 840
rect 855 839 856 843
rect 850 838 856 839
rect 1254 839 1260 840
rect 606 834 612 835
rect 1254 835 1255 839
rect 1259 838 1260 839
rect 1478 839 1484 840
rect 1478 838 1479 839
rect 1259 836 1479 838
rect 1259 835 1260 836
rect 1254 834 1260 835
rect 1478 835 1479 836
rect 1483 835 1484 839
rect 1478 834 1484 835
rect 664 832 706 834
rect 207 831 213 832
rect 207 827 208 831
rect 212 830 213 831
rect 215 831 221 832
rect 215 830 216 831
rect 212 828 216 830
rect 212 827 213 828
rect 207 826 213 827
rect 215 827 216 828
rect 220 827 221 831
rect 215 826 221 827
rect 247 831 253 832
rect 247 827 248 831
rect 252 827 253 831
rect 247 826 253 827
rect 303 831 309 832
rect 303 827 304 831
rect 308 830 309 831
rect 391 831 397 832
rect 391 830 392 831
rect 308 828 392 830
rect 308 827 309 828
rect 303 826 309 827
rect 391 827 392 828
rect 396 827 397 831
rect 391 826 397 827
rect 423 831 432 832
rect 423 827 424 831
rect 431 827 432 831
rect 423 826 432 827
rect 479 831 485 832
rect 479 827 480 831
rect 484 830 485 831
rect 574 831 580 832
rect 574 830 575 831
rect 484 828 575 830
rect 484 827 485 828
rect 479 826 485 827
rect 574 827 575 828
rect 579 827 580 831
rect 574 826 580 827
rect 655 827 661 828
rect 230 823 236 824
rect 230 819 231 823
rect 235 819 236 823
rect 230 818 236 819
rect 406 823 412 824
rect 406 819 407 823
rect 411 819 412 823
rect 655 823 656 827
rect 660 826 661 827
rect 664 826 666 832
rect 704 830 706 832
rect 799 831 805 832
rect 799 830 800 831
rect 704 828 800 830
rect 660 824 666 826
rect 671 827 677 828
rect 660 823 661 824
rect 655 822 661 823
rect 671 823 672 827
rect 676 826 677 827
rect 679 827 685 828
rect 679 826 680 827
rect 676 824 680 826
rect 676 823 677 824
rect 671 822 677 823
rect 679 823 680 824
rect 684 823 685 827
rect 679 822 685 823
rect 691 827 700 828
rect 691 823 692 827
rect 699 823 700 827
rect 799 827 800 828
rect 804 827 805 831
rect 799 826 805 827
rect 830 831 837 832
rect 830 827 831 831
rect 836 827 837 831
rect 830 826 837 827
rect 886 831 893 832
rect 886 827 887 831
rect 892 827 893 831
rect 886 826 893 827
rect 1278 831 1284 832
rect 1278 827 1279 831
rect 1283 830 1284 831
rect 1283 828 1430 830
rect 1283 827 1284 828
rect 1278 826 1284 827
rect 691 822 700 823
rect 814 823 820 824
rect 406 818 412 819
rect 814 819 815 823
rect 819 819 820 823
rect 814 818 820 819
rect 990 823 996 824
rect 990 819 991 823
rect 995 822 996 823
rect 1011 823 1017 824
rect 1011 822 1012 823
rect 995 820 1012 822
rect 995 819 996 820
rect 990 818 996 819
rect 1011 819 1012 820
rect 1016 819 1017 823
rect 1227 823 1236 824
rect 1227 822 1228 823
rect 1011 818 1017 819
rect 1035 821 1228 822
rect 662 817 668 818
rect 662 813 663 817
rect 667 813 668 817
rect 1035 817 1036 821
rect 1040 820 1228 821
rect 1040 817 1041 820
rect 1227 819 1228 820
rect 1235 819 1236 823
rect 1391 823 1397 824
rect 1363 821 1369 822
rect 1227 818 1236 819
rect 1251 819 1260 820
rect 1035 816 1041 817
rect 662 812 668 813
rect 1167 815 1173 816
rect 1167 811 1168 815
rect 1172 814 1173 815
rect 1251 815 1252 819
rect 1259 815 1260 819
rect 1363 817 1364 821
rect 1368 817 1369 821
rect 1391 819 1392 823
rect 1396 822 1397 823
rect 1414 823 1425 824
rect 1396 820 1410 822
rect 1396 819 1397 820
rect 1391 818 1397 819
rect 1363 816 1369 817
rect 1251 814 1260 815
rect 1354 815 1360 816
rect 1354 814 1355 815
rect 1172 812 1246 814
rect 1172 811 1173 812
rect 1167 810 1173 811
rect 1244 810 1246 812
rect 1305 812 1355 814
rect 1305 810 1307 812
rect 1354 811 1355 812
rect 1359 811 1360 815
rect 1354 810 1360 811
rect 1244 808 1307 810
rect 151 807 157 808
rect 110 804 116 805
rect 110 800 111 804
rect 115 800 116 804
rect 151 803 152 807
rect 156 806 157 807
rect 159 807 165 808
rect 159 806 160 807
rect 156 804 160 806
rect 156 803 157 804
rect 110 799 116 800
rect 134 802 140 803
rect 151 802 157 803
rect 159 803 160 804
rect 164 803 165 807
rect 575 807 581 808
rect 575 803 576 807
rect 580 806 581 807
rect 950 807 956 808
rect 580 804 630 806
rect 580 803 581 804
rect 159 802 165 803
rect 558 802 564 803
rect 575 802 581 803
rect 134 798 135 802
rect 139 798 140 802
rect 134 797 140 798
rect 558 798 559 802
rect 563 798 564 802
rect 558 797 564 798
rect 628 798 630 804
rect 950 803 951 807
rect 955 803 956 807
rect 1110 807 1116 808
rect 950 802 956 803
rect 1030 805 1036 806
rect 1030 801 1031 805
rect 1035 801 1036 805
rect 1030 800 1036 801
rect 1042 803 1048 804
rect 1042 799 1043 803
rect 1047 802 1048 803
rect 1051 803 1060 804
rect 1110 803 1111 807
rect 1115 806 1116 807
rect 1119 807 1128 808
rect 1119 806 1120 807
rect 1115 804 1120 806
rect 1115 803 1116 804
rect 1051 802 1052 803
rect 1047 800 1052 802
rect 1047 799 1048 800
rect 1042 798 1048 799
rect 1051 799 1052 800
rect 1059 799 1060 803
rect 1051 798 1060 799
rect 1102 802 1108 803
rect 1110 802 1116 803
rect 1119 803 1120 804
rect 1127 803 1128 807
rect 1194 807 1205 808
rect 1119 802 1128 803
rect 1166 805 1172 806
rect 1102 798 1103 802
rect 1107 798 1108 802
rect 1166 801 1167 805
rect 1171 801 1172 805
rect 1194 803 1195 807
rect 1199 803 1200 807
rect 1204 803 1205 807
rect 1311 807 1317 808
rect 1194 802 1205 803
rect 1246 805 1252 806
rect 1166 800 1172 801
rect 1246 801 1247 805
rect 1251 801 1252 805
rect 1246 800 1252 801
rect 1267 803 1273 804
rect 1267 799 1268 803
rect 1272 802 1273 803
rect 1278 803 1284 804
rect 1278 802 1279 803
rect 1272 800 1279 802
rect 1272 799 1273 800
rect 1267 798 1273 799
rect 1278 799 1279 800
rect 1283 799 1284 803
rect 1278 798 1284 799
rect 1294 803 1300 804
rect 1294 799 1295 803
rect 1299 799 1300 803
rect 1311 803 1312 807
rect 1316 806 1317 807
rect 1364 806 1366 816
rect 1408 810 1410 820
rect 1414 819 1415 823
rect 1419 819 1420 823
rect 1424 819 1425 823
rect 1414 818 1425 819
rect 1428 818 1430 828
rect 1467 823 1473 824
rect 1447 819 1453 820
rect 1447 818 1448 819
rect 1428 816 1448 818
rect 1447 815 1448 816
rect 1452 815 1453 819
rect 1467 819 1468 823
rect 1472 822 1473 823
rect 1478 823 1484 824
rect 1478 822 1479 823
rect 1472 820 1479 822
rect 1472 819 1473 820
rect 1467 818 1473 819
rect 1478 819 1479 820
rect 1483 819 1484 823
rect 1478 818 1484 819
rect 1494 819 1501 820
rect 1447 814 1453 815
rect 1494 815 1495 819
rect 1500 815 1501 819
rect 1494 814 1501 815
rect 1422 812 1428 813
rect 1408 808 1418 810
rect 1316 804 1322 806
rect 1364 804 1410 806
rect 1316 803 1317 804
rect 1311 802 1317 803
rect 1294 798 1300 799
rect 628 796 681 798
rect 1102 797 1108 798
rect 1270 795 1276 796
rect 150 791 157 792
rect 110 787 116 788
rect 110 783 111 787
rect 115 783 116 787
rect 150 787 151 791
rect 156 787 157 791
rect 150 786 157 787
rect 574 791 581 792
rect 574 787 575 791
rect 580 787 581 791
rect 1119 791 1125 792
rect 574 786 581 787
rect 967 787 973 788
rect 110 782 116 783
rect 134 785 140 786
rect 134 781 135 785
rect 139 781 140 785
rect 558 785 564 786
rect 134 780 140 781
rect 230 782 236 783
rect 230 778 231 782
rect 235 778 236 782
rect 230 777 236 778
rect 406 782 412 783
rect 406 778 407 782
rect 411 778 412 782
rect 558 781 559 785
rect 563 781 564 785
rect 950 784 956 785
rect 558 780 564 781
rect 814 782 820 783
rect 814 778 815 782
rect 819 778 820 782
rect 950 780 951 784
rect 955 780 956 784
rect 967 783 968 787
rect 972 786 973 787
rect 1119 787 1120 791
rect 1124 790 1125 791
rect 1158 791 1164 792
rect 1158 790 1159 791
rect 1124 788 1159 790
rect 1124 787 1125 788
rect 1119 786 1125 787
rect 1158 787 1159 788
rect 1163 787 1164 791
rect 1270 791 1271 795
rect 1275 794 1276 795
rect 1320 794 1322 804
rect 1326 803 1332 804
rect 1326 799 1327 803
rect 1331 799 1332 803
rect 1326 798 1332 799
rect 1408 798 1410 804
rect 1416 802 1418 808
rect 1422 808 1423 812
rect 1427 808 1428 812
rect 1422 807 1428 808
rect 1470 812 1476 813
rect 1470 808 1471 812
rect 1475 808 1476 812
rect 1537 808 1570 810
rect 1577 808 1602 810
rect 1609 808 1634 810
rect 1641 808 1666 810
rect 1470 807 1476 808
rect 1535 807 1541 808
rect 1441 804 1458 806
rect 1441 802 1443 804
rect 1416 800 1443 802
rect 1447 799 1453 800
rect 1447 798 1448 799
rect 1408 796 1448 798
rect 1447 795 1448 796
rect 1452 795 1453 799
rect 1456 798 1458 804
rect 1535 803 1536 807
rect 1540 803 1541 807
rect 1518 802 1524 803
rect 1535 802 1541 803
rect 1558 802 1564 803
rect 1495 799 1501 800
rect 1495 798 1496 799
rect 1456 796 1496 798
rect 1447 794 1453 795
rect 1495 795 1496 796
rect 1500 795 1501 799
rect 1518 798 1519 802
rect 1523 798 1524 802
rect 1518 797 1524 798
rect 1558 798 1559 802
rect 1563 798 1564 802
rect 1558 797 1564 798
rect 1495 794 1501 795
rect 1275 792 1306 794
rect 1320 792 1369 794
rect 1275 791 1276 792
rect 1270 790 1276 791
rect 1304 790 1306 792
rect 1311 791 1317 792
rect 1311 790 1312 791
rect 1304 788 1312 790
rect 1158 786 1164 787
rect 1311 787 1312 788
rect 1316 787 1317 791
rect 1311 786 1317 787
rect 1535 791 1541 792
rect 1535 787 1536 791
rect 1540 787 1541 791
rect 1568 790 1570 808
rect 1575 807 1581 808
rect 1575 803 1576 807
rect 1580 803 1581 807
rect 1575 802 1581 803
rect 1590 802 1596 803
rect 1590 798 1591 802
rect 1595 798 1596 802
rect 1590 797 1596 798
rect 1575 791 1581 792
rect 1575 790 1576 791
rect 1568 788 1576 790
rect 1535 786 1541 787
rect 1575 787 1576 788
rect 1580 787 1581 791
rect 1600 790 1602 808
rect 1607 807 1613 808
rect 1607 803 1608 807
rect 1612 803 1613 807
rect 1607 802 1613 803
rect 1622 802 1628 803
rect 1622 798 1623 802
rect 1627 798 1628 802
rect 1622 797 1628 798
rect 1607 791 1613 792
rect 1607 790 1608 791
rect 1600 788 1608 790
rect 1575 786 1581 787
rect 1607 787 1608 788
rect 1612 787 1613 791
rect 1632 790 1634 808
rect 1639 807 1645 808
rect 1639 803 1640 807
rect 1644 803 1645 807
rect 1639 802 1645 803
rect 1654 802 1660 803
rect 1654 798 1655 802
rect 1659 798 1660 802
rect 1654 797 1660 798
rect 1639 791 1645 792
rect 1639 790 1640 791
rect 1632 788 1640 790
rect 1607 786 1613 787
rect 1639 787 1640 788
rect 1644 787 1645 791
rect 1664 790 1666 808
rect 1670 807 1677 808
rect 1670 803 1671 807
rect 1676 803 1677 807
rect 1670 802 1677 803
rect 1694 804 1700 805
rect 1694 800 1695 804
rect 1699 800 1700 804
rect 1694 799 1700 800
rect 1671 791 1677 792
rect 1671 790 1672 791
rect 1664 788 1672 790
rect 1639 786 1645 787
rect 1671 787 1672 788
rect 1676 787 1677 791
rect 1671 786 1677 787
rect 1694 787 1700 788
rect 972 784 1010 786
rect 1102 785 1108 786
rect 1294 785 1300 786
rect 1518 785 1524 786
rect 972 783 973 784
rect 967 782 973 783
rect 950 779 956 780
rect 406 777 412 778
rect 654 777 660 778
rect 814 777 820 778
rect 654 773 655 777
rect 659 773 660 777
rect 654 772 660 773
rect 1008 774 1010 784
rect 1014 784 1020 785
rect 1014 780 1015 784
rect 1019 780 1020 784
rect 1102 781 1103 785
rect 1107 781 1108 785
rect 1102 780 1108 781
rect 1230 784 1236 785
rect 1230 780 1231 784
rect 1235 780 1236 784
rect 1294 781 1295 785
rect 1299 781 1300 785
rect 1294 780 1300 781
rect 1326 784 1332 785
rect 1326 780 1327 784
rect 1331 780 1332 784
rect 1014 779 1020 780
rect 1230 779 1236 780
rect 1326 779 1332 780
rect 1422 784 1428 785
rect 1422 780 1423 784
rect 1427 780 1428 784
rect 1422 779 1428 780
rect 1470 784 1476 785
rect 1470 780 1471 784
rect 1475 780 1476 784
rect 1518 781 1519 785
rect 1523 781 1524 785
rect 1518 780 1524 781
rect 1470 779 1476 780
rect 1498 779 1504 780
rect 1182 778 1188 779
rect 1034 775 1040 776
rect 1034 774 1035 775
rect 1008 772 1035 774
rect 1034 771 1035 772
rect 1039 771 1040 775
rect 1182 774 1183 778
rect 1187 774 1188 778
rect 1498 775 1499 779
rect 1503 778 1504 779
rect 1537 778 1539 786
rect 1558 785 1564 786
rect 1558 781 1559 785
rect 1563 781 1564 785
rect 1558 780 1564 781
rect 1590 785 1596 786
rect 1590 781 1591 785
rect 1595 781 1596 785
rect 1590 780 1596 781
rect 1622 785 1628 786
rect 1622 781 1623 785
rect 1627 781 1628 785
rect 1622 780 1628 781
rect 1654 785 1660 786
rect 1654 781 1655 785
rect 1659 781 1660 785
rect 1694 783 1695 787
rect 1699 783 1700 787
rect 1694 782 1700 783
rect 1654 780 1660 781
rect 1503 776 1539 778
rect 1503 775 1504 776
rect 1498 774 1504 775
rect 1182 773 1188 774
rect 1034 770 1040 771
rect 1158 771 1165 772
rect 1158 767 1159 771
rect 1164 767 1165 771
rect 1158 766 1165 767
rect 218 763 224 764
rect 218 759 219 763
rect 223 762 224 763
rect 263 763 269 764
rect 263 762 264 763
rect 223 760 264 762
rect 223 759 224 760
rect 218 758 224 759
rect 263 759 264 760
rect 268 759 269 763
rect 263 758 269 759
rect 1222 759 1228 760
rect 1222 755 1223 759
rect 1227 758 1228 759
rect 1379 759 1385 760
rect 1379 758 1380 759
rect 1227 756 1380 758
rect 1227 755 1228 756
rect 1222 754 1228 755
rect 1379 755 1380 756
rect 1384 755 1385 759
rect 1379 754 1385 755
rect 766 735 772 736
rect 214 732 220 733
rect 134 728 140 729
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 134 724 135 728
rect 139 724 140 728
rect 214 728 215 732
rect 219 728 220 732
rect 390 732 396 733
rect 214 727 220 728
rect 286 730 292 731
rect 286 726 287 730
rect 291 726 292 730
rect 390 728 391 732
rect 395 728 396 732
rect 766 731 767 735
rect 771 731 772 735
rect 998 735 1004 736
rect 998 731 999 735
rect 1003 731 1004 735
rect 390 727 396 728
rect 614 730 620 731
rect 766 730 772 731
rect 910 730 916 731
rect 998 730 1004 731
rect 1166 732 1172 733
rect 286 725 292 726
rect 614 726 615 730
rect 619 726 620 730
rect 614 725 620 726
rect 718 728 724 729
rect 134 723 140 724
rect 470 724 476 725
rect 718 724 719 728
rect 723 724 724 728
rect 862 727 868 728
rect 110 720 116 721
rect 470 720 471 724
rect 475 720 476 724
rect 202 719 208 720
rect 470 719 476 720
rect 567 723 573 724
rect 567 719 568 723
rect 572 722 573 723
rect 622 723 628 724
rect 718 723 724 724
rect 735 723 741 724
rect 622 722 623 723
rect 572 720 623 722
rect 572 719 573 720
rect 202 718 203 719
rect 197 716 203 718
rect 202 715 203 716
rect 207 715 208 719
rect 567 718 573 719
rect 622 719 623 720
rect 627 719 628 723
rect 622 718 628 719
rect 735 719 736 723
rect 740 722 741 723
rect 766 723 772 724
rect 766 722 767 723
rect 740 720 767 722
rect 740 719 741 720
rect 735 718 741 719
rect 766 719 767 720
rect 771 719 772 723
rect 862 723 863 727
rect 867 723 868 727
rect 910 726 911 730
rect 915 726 916 730
rect 1086 728 1092 729
rect 910 725 916 726
rect 862 722 868 723
rect 980 724 1017 726
rect 1086 724 1087 728
rect 1091 724 1092 728
rect 1166 728 1167 732
rect 1171 728 1172 732
rect 1166 727 1172 728
rect 1206 728 1212 729
rect 766 718 772 719
rect 842 719 848 720
rect 202 714 208 715
rect 842 715 843 719
rect 847 718 848 719
rect 879 719 885 720
rect 879 718 880 719
rect 847 716 880 718
rect 847 715 848 716
rect 842 714 848 715
rect 879 715 880 716
rect 884 715 885 719
rect 980 718 982 724
rect 1086 723 1092 724
rect 1206 724 1207 728
rect 1211 724 1212 728
rect 1206 723 1212 724
rect 1246 727 1252 728
rect 1246 723 1247 727
rect 1251 723 1252 727
rect 1246 722 1252 723
rect 1278 727 1284 728
rect 1278 723 1279 727
rect 1283 723 1284 727
rect 1278 722 1284 723
rect 1310 727 1316 728
rect 1310 723 1311 727
rect 1315 723 1316 727
rect 1310 722 1316 723
rect 1342 727 1348 728
rect 1342 723 1343 727
rect 1347 723 1348 727
rect 1342 722 1348 723
rect 1374 727 1380 728
rect 1374 723 1375 727
rect 1379 723 1380 727
rect 1374 722 1380 723
rect 1406 727 1412 728
rect 1406 723 1407 727
rect 1411 723 1412 727
rect 1406 722 1412 723
rect 1438 727 1444 728
rect 1438 723 1439 727
rect 1443 723 1444 727
rect 1438 722 1444 723
rect 1478 727 1484 728
rect 1478 723 1479 727
rect 1483 723 1484 727
rect 1478 722 1484 723
rect 1518 727 1524 728
rect 1518 723 1519 727
rect 1523 723 1524 727
rect 1518 722 1524 723
rect 1558 727 1564 728
rect 1558 723 1559 727
rect 1563 723 1564 727
rect 1558 722 1564 723
rect 1590 727 1596 728
rect 1590 723 1591 727
rect 1595 723 1596 727
rect 1590 722 1596 723
rect 1622 727 1628 728
rect 1622 723 1623 727
rect 1627 723 1628 727
rect 1622 722 1628 723
rect 1654 727 1660 728
rect 1654 723 1655 727
rect 1659 723 1660 727
rect 1654 722 1660 723
rect 1694 725 1700 726
rect 1694 721 1695 725
rect 1699 721 1700 725
rect 1694 720 1700 721
rect 1154 719 1160 720
rect 1154 718 1155 719
rect 879 714 885 715
rect 892 716 982 718
rect 1149 716 1155 718
rect 239 711 248 712
rect 110 708 116 709
rect 110 704 111 708
rect 115 704 116 708
rect 239 707 240 711
rect 247 707 248 711
rect 239 706 248 707
rect 415 711 424 712
rect 415 707 416 711
rect 423 707 424 711
rect 730 711 736 712
rect 415 706 424 707
rect 442 709 448 710
rect 442 705 443 709
rect 447 705 448 709
rect 730 707 731 711
rect 735 710 736 711
rect 862 710 868 711
rect 735 708 793 710
rect 735 707 736 708
rect 730 706 736 707
rect 862 706 863 710
rect 867 706 868 710
rect 442 704 448 705
rect 718 705 724 706
rect 862 705 868 706
rect 110 703 116 704
rect 718 701 719 705
rect 723 701 724 705
rect 718 700 724 701
rect 879 703 885 704
rect 79 699 85 700
rect 79 695 80 699
rect 84 698 85 699
rect 278 699 284 700
rect 278 698 279 699
rect 84 696 279 698
rect 84 695 85 696
rect 79 694 85 695
rect 278 695 279 696
rect 283 695 284 699
rect 278 694 284 695
rect 566 699 573 700
rect 566 695 567 699
rect 572 695 573 699
rect 879 699 880 703
rect 884 702 885 703
rect 892 702 894 716
rect 1154 715 1155 716
rect 1159 715 1160 719
rect 1154 714 1160 715
rect 1234 719 1240 720
rect 1234 715 1235 719
rect 1239 718 1240 719
rect 1263 719 1269 720
rect 1263 718 1264 719
rect 1239 716 1264 718
rect 1239 715 1240 716
rect 1234 714 1240 715
rect 1263 715 1264 716
rect 1268 715 1269 719
rect 1295 719 1301 720
rect 1295 718 1296 719
rect 1263 714 1269 715
rect 1288 716 1296 718
rect 1146 711 1152 712
rect 1146 707 1147 711
rect 1151 710 1152 711
rect 1191 711 1197 712
rect 1191 710 1192 711
rect 1151 708 1192 710
rect 1151 707 1152 708
rect 1146 706 1152 707
rect 1191 707 1192 708
rect 1196 710 1197 711
rect 1222 711 1228 712
rect 1196 708 1218 710
rect 1196 707 1197 708
rect 1191 706 1197 707
rect 884 700 894 702
rect 1216 702 1218 708
rect 1222 707 1223 711
rect 1227 710 1228 711
rect 1231 711 1237 712
rect 1231 710 1232 711
rect 1227 708 1232 710
rect 1227 707 1228 708
rect 1222 706 1228 707
rect 1231 707 1232 708
rect 1236 707 1237 711
rect 1231 706 1237 707
rect 1246 710 1252 711
rect 1246 706 1247 710
rect 1251 706 1252 710
rect 1246 705 1252 706
rect 1278 710 1284 711
rect 1278 706 1279 710
rect 1283 706 1284 710
rect 1278 705 1284 706
rect 1226 703 1232 704
rect 1226 702 1227 703
rect 1206 700 1212 701
rect 1216 700 1227 702
rect 884 699 885 700
rect 879 698 885 699
rect 991 699 997 700
rect 991 698 992 699
rect 961 696 992 698
rect 566 694 573 695
rect 774 695 780 696
rect 380 692 402 694
rect 142 690 148 691
rect 142 686 143 690
rect 147 686 148 690
rect 286 689 292 690
rect 190 687 196 688
rect 190 686 191 687
rect 142 685 148 686
rect 153 684 191 686
rect 153 682 155 684
rect 190 683 191 684
rect 195 683 196 687
rect 190 682 196 683
rect 214 685 220 686
rect 151 681 157 682
rect 87 679 93 680
rect 87 675 88 679
rect 92 678 93 679
rect 135 679 141 680
rect 135 678 136 679
rect 92 676 136 678
rect 92 675 93 676
rect 87 674 93 675
rect 135 675 136 676
rect 140 675 141 679
rect 151 677 152 681
rect 156 677 157 681
rect 214 681 215 685
rect 219 681 220 685
rect 286 685 287 689
rect 291 685 292 689
rect 286 684 292 685
rect 214 680 220 681
rect 151 676 157 677
rect 167 679 173 680
rect 135 674 141 675
rect 167 675 168 679
rect 172 678 173 679
rect 234 679 245 680
rect 172 676 198 678
rect 172 675 173 676
rect 167 674 173 675
rect 196 666 198 676
rect 202 675 208 676
rect 202 671 203 675
rect 207 674 208 675
rect 211 675 217 676
rect 211 674 212 675
rect 207 672 212 674
rect 207 671 208 672
rect 202 670 208 671
rect 211 671 212 672
rect 216 671 217 675
rect 234 675 235 679
rect 239 675 240 679
rect 244 675 245 679
rect 234 674 245 675
rect 302 679 309 680
rect 302 675 303 679
rect 308 678 309 679
rect 322 679 328 680
rect 322 678 323 679
rect 308 676 323 678
rect 308 675 309 676
rect 302 674 309 675
rect 322 675 323 676
rect 327 675 328 679
rect 322 674 328 675
rect 359 679 365 680
rect 359 675 360 679
rect 364 678 365 679
rect 380 678 382 692
rect 400 690 402 692
rect 599 691 605 692
rect 599 690 600 691
rect 400 688 600 690
rect 599 687 600 688
rect 604 687 605 691
rect 774 691 775 695
rect 779 691 780 695
rect 991 695 992 696
rect 996 695 997 699
rect 1206 696 1207 700
rect 1211 696 1212 700
rect 1226 699 1227 700
rect 1231 699 1232 703
rect 1226 698 1232 699
rect 1263 703 1269 704
rect 1263 699 1264 703
rect 1268 702 1269 703
rect 1288 702 1290 716
rect 1295 715 1296 716
rect 1300 715 1301 719
rect 1327 719 1333 720
rect 1327 718 1328 719
rect 1295 714 1301 715
rect 1320 716 1328 718
rect 1310 710 1316 711
rect 1310 706 1311 710
rect 1315 706 1316 710
rect 1310 705 1316 706
rect 1268 700 1290 702
rect 1295 703 1301 704
rect 1268 699 1269 700
rect 1263 698 1269 699
rect 1295 699 1296 703
rect 1300 702 1301 703
rect 1320 702 1322 716
rect 1327 715 1328 716
rect 1332 715 1333 719
rect 1359 719 1365 720
rect 1359 718 1360 719
rect 1327 714 1333 715
rect 1352 716 1360 718
rect 1342 710 1348 711
rect 1342 706 1343 710
rect 1347 706 1348 710
rect 1342 705 1348 706
rect 1300 700 1322 702
rect 1327 703 1333 704
rect 1300 699 1301 700
rect 1295 698 1301 699
rect 1327 699 1328 703
rect 1332 702 1333 703
rect 1352 702 1354 716
rect 1359 715 1360 716
rect 1364 715 1365 719
rect 1391 719 1397 720
rect 1391 718 1392 719
rect 1359 714 1365 715
rect 1384 716 1392 718
rect 1374 710 1380 711
rect 1374 706 1375 710
rect 1379 706 1380 710
rect 1374 705 1380 706
rect 1332 700 1354 702
rect 1359 703 1365 704
rect 1332 699 1333 700
rect 1327 698 1333 699
rect 1359 699 1360 703
rect 1364 702 1365 703
rect 1384 702 1386 716
rect 1391 715 1392 716
rect 1396 715 1397 719
rect 1423 719 1429 720
rect 1423 718 1424 719
rect 1391 714 1397 715
rect 1416 716 1424 718
rect 1406 710 1412 711
rect 1406 706 1407 710
rect 1411 706 1412 710
rect 1406 705 1412 706
rect 1364 700 1386 702
rect 1391 703 1397 704
rect 1364 699 1365 700
rect 1359 698 1365 699
rect 1391 699 1392 703
rect 1396 702 1397 703
rect 1416 702 1418 716
rect 1423 715 1424 716
rect 1428 715 1429 719
rect 1455 719 1461 720
rect 1455 718 1456 719
rect 1423 714 1429 715
rect 1432 716 1456 718
rect 1396 700 1418 702
rect 1423 703 1429 704
rect 1396 699 1397 700
rect 1391 698 1397 699
rect 1423 699 1424 703
rect 1428 702 1429 703
rect 1432 702 1434 716
rect 1455 715 1456 716
rect 1460 715 1461 719
rect 1455 714 1461 715
rect 1495 719 1501 720
rect 1495 715 1496 719
rect 1500 718 1501 719
rect 1535 719 1541 720
rect 1500 716 1514 718
rect 1500 715 1501 716
rect 1495 714 1501 715
rect 1438 710 1444 711
rect 1438 706 1439 710
rect 1443 706 1444 710
rect 1438 705 1444 706
rect 1478 710 1484 711
rect 1478 706 1479 710
rect 1483 706 1484 710
rect 1478 705 1484 706
rect 1428 700 1434 702
rect 1446 703 1452 704
rect 1428 699 1429 700
rect 1423 698 1429 699
rect 1446 699 1447 703
rect 1451 702 1452 703
rect 1455 703 1461 704
rect 1455 702 1456 703
rect 1451 700 1456 702
rect 1451 699 1452 700
rect 1446 698 1452 699
rect 1455 699 1456 700
rect 1460 699 1461 703
rect 1455 698 1461 699
rect 1495 703 1504 704
rect 1495 699 1496 703
rect 1503 699 1504 703
rect 1512 702 1514 716
rect 1535 715 1536 719
rect 1540 718 1541 719
rect 1575 719 1581 720
rect 1540 716 1570 718
rect 1540 715 1541 716
rect 1535 714 1541 715
rect 1518 710 1524 711
rect 1518 706 1519 710
rect 1523 706 1524 710
rect 1518 705 1524 706
rect 1558 710 1564 711
rect 1558 706 1559 710
rect 1563 706 1564 710
rect 1558 705 1564 706
rect 1535 703 1541 704
rect 1535 702 1536 703
rect 1512 700 1536 702
rect 1495 698 1504 699
rect 1535 699 1536 700
rect 1540 699 1541 703
rect 1568 702 1570 716
rect 1575 715 1576 719
rect 1580 718 1581 719
rect 1607 719 1613 720
rect 1580 716 1602 718
rect 1580 715 1581 716
rect 1575 714 1581 715
rect 1590 710 1596 711
rect 1590 706 1591 710
rect 1595 706 1596 710
rect 1590 705 1596 706
rect 1575 703 1581 704
rect 1575 702 1576 703
rect 1568 700 1576 702
rect 1535 698 1541 699
rect 1575 699 1576 700
rect 1580 699 1581 703
rect 1600 702 1602 716
rect 1607 715 1608 719
rect 1612 718 1613 719
rect 1639 719 1645 720
rect 1612 716 1634 718
rect 1612 715 1613 716
rect 1607 714 1613 715
rect 1622 710 1628 711
rect 1622 706 1623 710
rect 1627 706 1628 710
rect 1622 705 1628 706
rect 1607 703 1613 704
rect 1607 702 1608 703
rect 1600 700 1608 702
rect 1575 698 1581 699
rect 1607 699 1608 700
rect 1612 699 1613 703
rect 1632 702 1634 716
rect 1639 715 1640 719
rect 1644 718 1645 719
rect 1670 719 1677 720
rect 1644 716 1666 718
rect 1644 715 1645 716
rect 1639 714 1645 715
rect 1654 710 1660 711
rect 1654 706 1655 710
rect 1659 706 1660 710
rect 1654 705 1660 706
rect 1639 703 1645 704
rect 1639 702 1640 703
rect 1632 700 1640 702
rect 1607 698 1613 699
rect 1639 699 1640 700
rect 1644 699 1645 703
rect 1664 702 1666 716
rect 1670 715 1671 719
rect 1676 715 1677 719
rect 1670 714 1677 715
rect 1694 708 1700 709
rect 1694 704 1695 708
rect 1699 704 1700 708
rect 1671 703 1677 704
rect 1694 703 1700 704
rect 1671 702 1672 703
rect 1664 700 1672 702
rect 1639 698 1645 699
rect 1671 699 1672 700
rect 1676 699 1677 703
rect 1671 698 1677 699
rect 991 694 997 695
rect 1006 695 1012 696
rect 1206 695 1212 696
rect 774 690 780 691
rect 850 691 856 692
rect 850 690 851 691
rect 599 686 605 687
rect 614 689 620 690
rect 390 685 396 686
rect 390 681 391 685
rect 395 681 396 685
rect 614 685 615 689
rect 619 685 620 689
rect 785 688 851 690
rect 746 687 752 688
rect 746 686 747 687
rect 614 684 620 685
rect 676 684 747 686
rect 390 680 396 681
rect 426 683 432 684
rect 364 676 382 678
rect 410 679 421 680
rect 364 675 365 676
rect 359 674 365 675
rect 387 675 393 676
rect 211 670 217 671
rect 387 671 388 675
rect 392 674 393 675
rect 398 675 404 676
rect 398 674 399 675
rect 392 672 399 674
rect 392 671 393 672
rect 387 670 393 671
rect 398 671 399 672
rect 403 671 404 675
rect 410 675 411 679
rect 415 675 416 679
rect 420 675 421 679
rect 426 679 427 683
rect 431 682 432 683
rect 431 680 558 682
rect 431 679 432 680
rect 426 678 432 679
rect 554 679 560 680
rect 410 674 421 675
rect 522 675 528 676
rect 398 670 404 671
rect 522 671 523 675
rect 527 671 528 675
rect 554 675 555 679
rect 559 678 560 679
rect 631 679 637 680
rect 631 678 632 679
rect 559 676 632 678
rect 559 675 560 676
rect 554 674 560 675
rect 631 675 632 676
rect 636 678 637 679
rect 676 678 678 684
rect 746 683 747 684
rect 751 683 752 687
rect 785 684 787 688
rect 850 687 851 688
rect 855 687 856 691
rect 1006 691 1007 695
rect 1011 691 1012 695
rect 1231 691 1240 692
rect 1006 690 1012 691
rect 1094 690 1100 691
rect 850 686 856 687
rect 910 689 916 690
rect 910 685 911 689
rect 915 685 916 689
rect 1094 686 1095 690
rect 1099 686 1100 690
rect 1203 687 1209 688
rect 1094 685 1100 686
rect 1166 685 1172 686
rect 910 684 916 685
rect 746 682 752 683
rect 758 683 764 684
rect 636 676 678 678
rect 687 679 693 680
rect 636 675 637 676
rect 631 674 637 675
rect 687 675 688 679
rect 692 678 693 679
rect 758 679 759 683
rect 763 682 764 683
rect 767 683 773 684
rect 767 682 768 683
rect 763 680 768 682
rect 763 679 764 680
rect 758 678 764 679
rect 767 679 768 680
rect 772 679 773 683
rect 767 678 773 679
rect 783 683 789 684
rect 783 679 784 683
rect 788 679 789 683
rect 803 683 809 684
rect 803 682 804 683
rect 783 678 789 679
rect 792 680 804 682
rect 692 676 754 678
rect 692 675 693 676
rect 687 674 693 675
rect 522 670 528 671
rect 242 667 248 668
rect 242 666 243 667
rect 196 664 243 666
rect 242 663 243 664
rect 247 663 248 667
rect 242 662 248 663
rect 314 667 320 668
rect 314 663 315 667
rect 319 666 320 667
rect 410 667 416 668
rect 410 666 411 667
rect 319 664 411 666
rect 319 663 320 664
rect 314 662 320 663
rect 410 663 411 664
rect 415 663 416 667
rect 410 662 416 663
rect 418 667 424 668
rect 418 663 419 667
rect 423 666 424 667
rect 458 667 464 668
rect 458 666 459 667
rect 423 664 459 666
rect 423 663 424 664
rect 418 662 424 663
rect 458 663 459 664
rect 463 663 464 667
rect 752 666 754 676
rect 766 675 772 676
rect 766 671 767 675
rect 771 674 772 675
rect 792 674 794 680
rect 803 679 804 680
rect 808 679 809 683
rect 991 683 997 684
rect 803 678 809 679
rect 830 679 836 680
rect 830 675 831 679
rect 835 678 836 679
rect 927 679 933 680
rect 927 678 928 679
rect 835 676 928 678
rect 835 675 836 676
rect 830 674 836 675
rect 927 675 928 676
rect 932 675 933 679
rect 927 674 933 675
rect 982 679 989 680
rect 982 675 983 679
rect 988 675 989 679
rect 991 679 992 683
rect 996 682 997 683
rect 999 683 1005 684
rect 999 682 1000 683
rect 996 680 1000 682
rect 996 679 997 680
rect 991 678 997 679
rect 999 679 1000 680
rect 1004 679 1005 683
rect 999 678 1005 679
rect 1014 683 1021 684
rect 1014 679 1015 683
rect 1020 679 1021 683
rect 1014 678 1021 679
rect 1034 683 1041 684
rect 1034 679 1035 683
rect 1040 679 1041 683
rect 1166 681 1167 685
rect 1171 681 1172 685
rect 1203 683 1204 687
rect 1208 683 1209 687
rect 1231 687 1232 691
rect 1239 687 1240 691
rect 1231 686 1240 687
rect 1454 691 1460 692
rect 1454 687 1455 691
rect 1459 690 1460 691
rect 1747 691 1753 692
rect 1747 690 1748 691
rect 1459 688 1748 690
rect 1459 687 1460 688
rect 1454 686 1460 687
rect 1747 687 1748 688
rect 1752 687 1753 691
rect 1747 686 1753 687
rect 1203 682 1209 683
rect 1166 680 1172 681
rect 1034 678 1041 679
rect 1086 679 1093 680
rect 982 674 989 675
rect 1086 675 1087 679
rect 1092 675 1093 679
rect 1086 674 1093 675
rect 1102 679 1109 680
rect 1102 675 1103 679
rect 1108 675 1109 679
rect 1102 674 1109 675
rect 1119 679 1125 680
rect 1119 675 1120 679
rect 1124 678 1125 679
rect 1146 679 1152 680
rect 1146 678 1147 679
rect 1124 676 1147 678
rect 1124 675 1125 676
rect 1119 674 1125 675
rect 1146 675 1147 676
rect 1151 675 1152 679
rect 1182 679 1188 680
rect 1146 674 1152 675
rect 1154 675 1160 676
rect 771 672 794 674
rect 771 671 772 672
rect 766 670 772 671
rect 929 670 931 674
rect 1062 671 1068 672
rect 1062 670 1063 671
rect 929 668 1063 670
rect 842 667 848 668
rect 842 666 843 667
rect 752 664 843 666
rect 458 662 464 663
rect 842 663 843 664
rect 847 663 848 667
rect 1062 667 1063 668
rect 1067 667 1068 671
rect 1154 671 1155 675
rect 1159 674 1160 675
rect 1163 675 1169 676
rect 1163 674 1164 675
rect 1159 672 1164 674
rect 1159 671 1160 672
rect 1154 670 1160 671
rect 1163 671 1164 672
rect 1168 671 1169 675
rect 1182 675 1183 679
rect 1187 678 1188 679
rect 1191 679 1197 680
rect 1191 678 1192 679
rect 1187 676 1192 678
rect 1187 675 1188 676
rect 1182 674 1188 675
rect 1191 675 1192 676
rect 1196 678 1197 679
rect 1204 678 1206 682
rect 1254 679 1260 680
rect 1254 678 1255 679
rect 1196 676 1255 678
rect 1196 675 1197 676
rect 1191 674 1197 675
rect 1254 675 1255 676
rect 1259 678 1260 679
rect 1358 679 1364 680
rect 1358 678 1359 679
rect 1259 676 1359 678
rect 1259 675 1260 676
rect 1254 674 1260 675
rect 1358 675 1359 676
rect 1363 675 1364 679
rect 1358 674 1364 675
rect 1163 670 1169 671
rect 1062 666 1068 667
rect 842 662 848 663
rect 850 663 856 664
rect 242 659 248 660
rect 242 655 243 659
rect 247 658 248 659
rect 850 659 851 663
rect 855 662 856 663
rect 1014 663 1020 664
rect 1014 662 1015 663
rect 855 660 1015 662
rect 855 659 856 660
rect 850 658 856 659
rect 1014 659 1015 660
rect 1019 662 1020 663
rect 1110 663 1116 664
rect 1110 662 1111 663
rect 1019 660 1111 662
rect 1019 659 1020 660
rect 1014 658 1020 659
rect 1110 659 1111 660
rect 1115 662 1116 663
rect 1115 660 1161 662
rect 1115 659 1116 660
rect 1110 658 1116 659
rect 1159 658 1161 660
rect 1174 659 1180 660
rect 1174 658 1175 659
rect 247 656 449 658
rect 1159 656 1175 658
rect 247 655 248 656
rect 242 654 248 655
rect 1015 655 1021 656
rect 1015 651 1016 655
rect 1020 654 1021 655
rect 1102 655 1108 656
rect 1102 654 1103 655
rect 1020 652 1103 654
rect 1020 651 1021 652
rect 1015 650 1021 651
rect 1102 651 1103 652
rect 1107 651 1108 655
rect 1174 655 1175 656
rect 1179 655 1180 659
rect 1174 654 1180 655
rect 1102 650 1108 651
rect 234 647 240 648
rect 234 643 235 647
rect 239 646 240 647
rect 314 647 320 648
rect 314 646 315 647
rect 239 644 315 646
rect 239 643 240 644
rect 234 642 240 643
rect 314 643 315 644
rect 319 643 320 647
rect 314 642 320 643
rect 1078 643 1084 644
rect 294 639 300 640
rect 294 638 295 639
rect 203 637 295 638
rect 203 633 204 637
rect 208 636 295 637
rect 208 633 209 636
rect 294 635 295 636
rect 299 635 300 639
rect 294 634 300 635
rect 338 639 344 640
rect 338 635 339 639
rect 343 638 344 639
rect 634 639 640 640
rect 343 636 418 638
rect 343 635 344 636
rect 338 634 344 635
rect 203 632 209 633
rect 416 632 418 636
rect 634 635 635 639
rect 639 638 640 639
rect 1078 639 1079 643
rect 1083 642 1084 643
rect 1083 640 1146 642
rect 1083 639 1084 640
rect 1078 638 1084 639
rect 1144 638 1146 640
rect 1182 639 1188 640
rect 1182 638 1183 639
rect 639 636 794 638
rect 1144 636 1183 638
rect 639 635 640 636
rect 634 634 640 635
rect 231 631 240 632
rect 206 627 212 628
rect 206 623 207 627
rect 211 623 212 627
rect 231 627 232 631
rect 239 627 240 631
rect 231 626 240 627
rect 278 631 285 632
rect 278 627 279 631
rect 284 627 285 631
rect 278 626 285 627
rect 287 631 293 632
rect 287 627 288 631
rect 292 630 293 631
rect 295 631 301 632
rect 295 630 296 631
rect 292 628 296 630
rect 292 627 293 628
rect 287 626 293 627
rect 295 627 296 628
rect 300 627 301 631
rect 295 626 301 627
rect 306 631 317 632
rect 306 627 307 631
rect 311 627 312 631
rect 316 630 317 631
rect 399 631 405 632
rect 399 630 400 631
rect 316 628 400 630
rect 316 627 317 628
rect 306 626 317 627
rect 399 627 400 628
rect 404 627 405 631
rect 399 626 405 627
rect 414 631 421 632
rect 414 627 415 631
rect 420 627 421 631
rect 414 626 421 627
rect 431 631 437 632
rect 431 627 432 631
rect 436 630 437 631
rect 458 631 464 632
rect 458 630 459 631
rect 436 628 459 630
rect 436 627 437 628
rect 431 626 437 627
rect 458 627 459 628
rect 463 627 464 631
rect 458 626 464 627
rect 518 631 524 632
rect 518 627 519 631
rect 523 630 524 631
rect 551 631 560 632
rect 551 630 552 631
rect 523 628 552 630
rect 523 627 524 628
rect 518 626 524 627
rect 551 627 552 628
rect 559 627 560 631
rect 551 626 560 627
rect 607 631 613 632
rect 607 627 608 631
rect 612 630 613 631
rect 686 631 692 632
rect 686 630 687 631
rect 612 628 687 630
rect 612 627 613 628
rect 607 626 613 627
rect 686 627 687 628
rect 691 627 692 631
rect 686 626 692 627
rect 783 631 789 632
rect 783 627 784 631
rect 788 627 789 631
rect 792 630 794 636
rect 899 635 905 636
rect 839 631 845 632
rect 839 630 840 631
rect 792 628 840 630
rect 783 626 789 627
rect 839 627 840 628
rect 844 627 845 631
rect 899 631 900 635
rect 904 634 905 635
rect 918 635 924 636
rect 918 634 919 635
rect 904 632 919 634
rect 904 631 905 632
rect 899 630 905 631
rect 918 631 919 632
rect 923 631 924 635
rect 1050 635 1056 636
rect 918 630 924 631
rect 927 631 933 632
rect 839 626 845 627
rect 902 627 908 628
rect 785 624 834 626
rect 534 623 540 624
rect 206 622 212 623
rect 286 622 292 623
rect 286 618 287 622
rect 291 618 292 622
rect 286 617 292 618
rect 406 622 412 623
rect 406 618 407 622
rect 411 618 412 622
rect 534 619 535 623
rect 539 619 540 623
rect 534 618 540 619
rect 766 623 772 624
rect 766 619 767 623
rect 771 619 772 623
rect 766 618 772 619
rect 830 623 836 624
rect 830 619 831 623
rect 835 619 836 623
rect 902 623 903 627
rect 907 623 908 627
rect 927 627 928 631
rect 932 630 933 631
rect 950 631 956 632
rect 950 630 951 631
rect 932 628 951 630
rect 932 627 933 628
rect 927 626 933 627
rect 950 627 951 628
rect 955 627 956 631
rect 950 626 956 627
rect 982 631 988 632
rect 982 627 983 631
rect 987 630 988 631
rect 991 631 997 632
rect 991 630 992 631
rect 987 628 992 630
rect 987 627 988 628
rect 982 626 988 627
rect 991 627 992 628
rect 996 627 997 631
rect 991 626 997 627
rect 1006 631 1013 632
rect 1006 627 1007 631
rect 1012 630 1013 631
rect 1015 631 1021 632
rect 1015 630 1016 631
rect 1012 628 1016 630
rect 1012 627 1013 628
rect 1006 626 1013 627
rect 1015 627 1016 628
rect 1020 627 1021 631
rect 1015 626 1021 627
rect 1023 631 1029 632
rect 1023 627 1024 631
rect 1028 630 1029 631
rect 1050 631 1051 635
rect 1055 634 1056 635
rect 1115 635 1121 636
rect 1115 634 1116 635
rect 1055 632 1116 634
rect 1055 631 1056 632
rect 1050 630 1056 631
rect 1115 631 1116 632
rect 1120 631 1121 635
rect 1144 632 1146 636
rect 1182 635 1183 636
rect 1187 635 1188 639
rect 1182 634 1188 635
rect 1266 635 1272 636
rect 1115 630 1121 631
rect 1142 631 1149 632
rect 1028 628 1046 630
rect 1028 627 1029 628
rect 1023 626 1029 627
rect 1044 626 1046 628
rect 1110 627 1116 628
rect 1110 626 1111 627
rect 1044 624 1111 626
rect 1110 623 1111 624
rect 1115 623 1116 627
rect 902 622 908 623
rect 998 622 1004 623
rect 1110 622 1116 623
rect 1118 627 1124 628
rect 1118 623 1119 627
rect 1123 623 1124 627
rect 1142 627 1143 631
rect 1148 627 1149 631
rect 1142 626 1149 627
rect 1151 631 1157 632
rect 1151 627 1152 631
rect 1156 630 1157 631
rect 1207 631 1213 632
rect 1207 630 1208 631
rect 1156 628 1208 630
rect 1156 627 1157 628
rect 1151 626 1157 627
rect 1207 627 1208 628
rect 1212 627 1213 631
rect 1207 626 1213 627
rect 1222 631 1229 632
rect 1222 627 1223 631
rect 1228 627 1229 631
rect 1222 626 1229 627
rect 1239 631 1245 632
rect 1239 627 1240 631
rect 1244 630 1245 631
rect 1266 631 1267 635
rect 1271 634 1272 635
rect 1331 635 1337 636
rect 1331 634 1332 635
rect 1271 632 1332 634
rect 1271 631 1272 632
rect 1266 630 1272 631
rect 1331 631 1332 632
rect 1336 631 1337 635
rect 1331 630 1337 631
rect 1358 631 1365 632
rect 1244 628 1258 630
rect 1244 627 1245 628
rect 1239 626 1245 627
rect 1118 622 1124 623
rect 1214 622 1220 623
rect 830 618 836 619
rect 998 618 999 622
rect 1003 618 1004 622
rect 406 617 412 618
rect 998 617 1004 618
rect 1214 618 1215 622
rect 1219 618 1220 622
rect 1214 617 1220 618
rect 1256 618 1258 628
rect 1334 627 1340 628
rect 1334 623 1335 627
rect 1339 623 1340 627
rect 1358 627 1359 631
rect 1364 627 1365 631
rect 1358 626 1365 627
rect 1334 622 1340 623
rect 1346 619 1352 620
rect 1346 618 1347 619
rect 1256 616 1347 618
rect 758 615 764 616
rect 526 611 532 612
rect 150 607 157 608
rect 110 604 116 605
rect 110 600 111 604
rect 115 600 116 604
rect 150 603 151 607
rect 156 603 157 607
rect 183 607 189 608
rect 183 603 184 607
rect 188 606 189 607
rect 254 607 260 608
rect 254 606 255 607
rect 188 604 255 606
rect 188 603 189 604
rect 110 599 116 600
rect 134 602 140 603
rect 150 602 157 603
rect 166 602 172 603
rect 183 602 189 603
rect 254 603 255 604
rect 259 603 260 607
rect 526 607 527 611
rect 531 607 532 611
rect 758 611 759 615
rect 763 611 764 615
rect 1346 615 1347 616
rect 1351 615 1352 619
rect 1670 619 1676 620
rect 1670 618 1671 619
rect 1346 614 1352 615
rect 1496 616 1671 618
rect 758 610 764 611
rect 1496 608 1498 616
rect 1670 615 1671 616
rect 1675 615 1676 619
rect 1670 614 1676 615
rect 1503 611 1509 612
rect 526 606 532 607
rect 687 607 693 608
rect 687 603 688 607
rect 692 606 693 607
rect 730 607 736 608
rect 730 606 731 607
rect 692 604 731 606
rect 692 603 693 604
rect 254 602 260 603
rect 670 602 676 603
rect 687 602 693 603
rect 730 603 731 604
rect 735 603 736 607
rect 1151 607 1157 608
rect 1151 606 1152 607
rect 730 602 736 603
rect 1049 604 1152 606
rect 134 598 135 602
rect 139 598 140 602
rect 134 597 140 598
rect 166 598 167 602
rect 171 598 172 602
rect 166 597 172 598
rect 231 599 237 600
rect 231 595 232 599
rect 236 598 237 599
rect 286 599 292 600
rect 286 598 287 599
rect 236 596 287 598
rect 236 595 237 596
rect 231 594 237 595
rect 286 595 287 596
rect 291 595 292 599
rect 670 598 671 602
rect 675 598 676 602
rect 1049 600 1051 604
rect 1151 603 1152 604
rect 1156 603 1157 607
rect 1431 607 1440 608
rect 1431 603 1432 607
rect 1439 603 1440 607
rect 1495 607 1501 608
rect 1495 603 1496 607
rect 1500 603 1501 607
rect 1503 607 1504 611
rect 1508 610 1509 611
rect 1567 611 1573 612
rect 1508 608 1554 610
rect 1508 607 1509 608
rect 1503 606 1509 607
rect 1552 606 1554 608
rect 1559 607 1565 608
rect 1559 606 1560 607
rect 1552 604 1560 606
rect 1559 603 1560 604
rect 1564 603 1565 607
rect 1567 607 1568 611
rect 1572 610 1573 611
rect 1631 611 1637 612
rect 1572 608 1618 610
rect 1572 607 1573 608
rect 1567 606 1573 607
rect 1616 606 1618 608
rect 1623 607 1629 608
rect 1623 606 1624 607
rect 1616 604 1624 606
rect 1623 603 1624 604
rect 1628 603 1629 607
rect 1631 607 1632 611
rect 1636 610 1637 611
rect 1636 608 1675 610
rect 1636 607 1637 608
rect 1631 606 1637 607
rect 1671 607 1677 608
rect 1671 603 1672 607
rect 1676 603 1677 607
rect 1151 602 1157 603
rect 1414 602 1420 603
rect 1431 602 1440 603
rect 1478 602 1484 603
rect 1495 602 1501 603
rect 1542 602 1548 603
rect 1559 602 1565 603
rect 1606 602 1612 603
rect 1623 602 1629 603
rect 1654 602 1660 603
rect 1671 602 1677 603
rect 1694 604 1700 605
rect 670 597 676 598
rect 927 599 933 600
rect 286 594 292 595
rect 294 595 300 596
rect 150 591 157 592
rect 110 587 116 588
rect 110 583 111 587
rect 115 583 116 587
rect 150 587 151 591
rect 156 587 157 591
rect 150 586 157 587
rect 182 591 189 592
rect 182 587 183 591
rect 188 587 189 591
rect 294 591 295 595
rect 299 591 300 595
rect 294 590 300 591
rect 398 595 404 596
rect 398 591 399 595
rect 403 594 404 595
rect 927 595 928 599
rect 932 598 933 599
rect 958 599 964 600
rect 958 598 959 599
rect 932 596 959 598
rect 932 595 933 596
rect 927 594 933 595
rect 958 595 959 596
rect 963 598 964 599
rect 1044 598 1051 600
rect 1110 599 1116 600
rect 963 596 1046 598
rect 963 595 964 596
rect 958 594 964 595
rect 1050 595 1056 596
rect 403 592 417 594
rect 403 591 404 592
rect 398 590 404 591
rect 686 591 693 592
rect 182 586 189 587
rect 686 587 687 591
rect 692 587 693 591
rect 1050 591 1051 595
rect 1055 591 1056 595
rect 1110 595 1111 599
rect 1115 598 1116 599
rect 1143 599 1149 600
rect 1143 598 1144 599
rect 1115 596 1144 598
rect 1115 595 1116 596
rect 1110 594 1116 595
rect 1143 595 1144 596
rect 1148 598 1149 599
rect 1175 599 1181 600
rect 1175 598 1176 599
rect 1148 596 1176 598
rect 1148 595 1149 596
rect 1143 594 1149 595
rect 1175 595 1176 596
rect 1180 595 1181 599
rect 1346 599 1352 600
rect 1175 594 1181 595
rect 1266 595 1272 596
rect 1050 590 1056 591
rect 1266 591 1267 595
rect 1271 591 1272 595
rect 1346 595 1347 599
rect 1351 598 1352 599
rect 1359 599 1365 600
rect 1359 598 1360 599
rect 1351 596 1360 598
rect 1351 595 1352 596
rect 1346 594 1352 595
rect 1359 595 1360 596
rect 1364 595 1365 599
rect 1414 598 1415 602
rect 1419 598 1420 602
rect 1414 597 1420 598
rect 1478 598 1479 602
rect 1483 598 1484 602
rect 1478 597 1484 598
rect 1542 598 1543 602
rect 1547 598 1548 602
rect 1542 597 1548 598
rect 1606 598 1607 602
rect 1611 598 1612 602
rect 1606 597 1612 598
rect 1654 598 1655 602
rect 1659 598 1660 602
rect 1694 600 1695 604
rect 1699 600 1700 604
rect 1694 599 1700 600
rect 1654 597 1660 598
rect 1359 594 1365 595
rect 1266 590 1272 591
rect 1431 591 1437 592
rect 686 586 693 587
rect 1431 587 1432 591
rect 1436 590 1437 591
rect 1446 591 1452 592
rect 1446 590 1447 591
rect 1436 588 1447 590
rect 1436 587 1437 588
rect 1431 586 1437 587
rect 1446 587 1447 588
rect 1451 587 1452 591
rect 1446 586 1452 587
rect 1495 591 1501 592
rect 1495 587 1496 591
rect 1500 590 1501 591
rect 1503 591 1509 592
rect 1503 590 1504 591
rect 1500 588 1504 590
rect 1500 587 1501 588
rect 1495 586 1501 587
rect 1503 587 1504 588
rect 1508 587 1509 591
rect 1503 586 1509 587
rect 1559 591 1565 592
rect 1559 587 1560 591
rect 1564 590 1565 591
rect 1567 591 1573 592
rect 1567 590 1568 591
rect 1564 588 1568 590
rect 1564 587 1565 588
rect 1559 586 1565 587
rect 1567 587 1568 588
rect 1572 587 1573 591
rect 1567 586 1573 587
rect 1623 591 1629 592
rect 1623 587 1624 591
rect 1628 590 1629 591
rect 1631 591 1637 592
rect 1631 590 1632 591
rect 1628 588 1632 590
rect 1628 587 1629 588
rect 1623 586 1629 587
rect 1631 587 1632 588
rect 1636 587 1637 591
rect 1631 586 1637 587
rect 1670 591 1677 592
rect 1670 587 1671 591
rect 1676 587 1677 591
rect 1670 586 1677 587
rect 1694 587 1700 588
rect 110 582 116 583
rect 134 585 140 586
rect 134 581 135 585
rect 139 581 140 585
rect 134 580 140 581
rect 166 585 172 586
rect 670 585 676 586
rect 1414 585 1420 586
rect 166 581 167 585
rect 171 581 172 585
rect 278 584 284 585
rect 166 580 172 581
rect 206 580 212 581
rect 206 576 207 580
rect 211 576 212 580
rect 278 580 279 584
rect 283 580 284 584
rect 278 579 284 580
rect 398 584 404 585
rect 398 580 399 584
rect 403 580 404 584
rect 398 579 404 580
rect 534 582 540 583
rect 534 578 535 582
rect 539 578 540 582
rect 670 581 671 585
rect 675 581 676 585
rect 990 584 996 585
rect 670 580 676 581
rect 766 582 772 583
rect 534 577 540 578
rect 766 578 767 582
rect 771 578 772 582
rect 766 577 772 578
rect 902 580 908 581
rect 206 575 212 576
rect 902 576 903 580
rect 907 576 908 580
rect 990 580 991 584
rect 995 580 996 584
rect 1206 584 1212 585
rect 990 579 996 580
rect 1118 580 1124 581
rect 902 575 908 576
rect 1118 576 1119 580
rect 1123 576 1124 580
rect 1206 580 1207 584
rect 1211 580 1212 584
rect 1414 581 1415 585
rect 1419 581 1420 585
rect 1206 579 1212 580
rect 1334 580 1340 581
rect 1414 580 1420 581
rect 1478 585 1484 586
rect 1478 581 1479 585
rect 1483 581 1484 585
rect 1478 580 1484 581
rect 1542 585 1548 586
rect 1542 581 1543 585
rect 1547 581 1548 585
rect 1542 580 1548 581
rect 1606 585 1612 586
rect 1606 581 1607 585
rect 1611 581 1612 585
rect 1606 580 1612 581
rect 1654 585 1660 586
rect 1654 581 1655 585
rect 1659 581 1660 585
rect 1694 583 1695 587
rect 1699 583 1700 587
rect 1694 582 1700 583
rect 1654 580 1660 581
rect 1118 575 1124 576
rect 1334 576 1335 580
rect 1339 576 1340 580
rect 1334 575 1340 576
rect 1102 567 1108 568
rect 378 563 384 564
rect 378 559 379 563
rect 383 562 384 563
rect 526 563 532 564
rect 526 562 527 563
rect 383 560 527 562
rect 383 559 384 560
rect 378 558 384 559
rect 526 559 527 560
rect 531 559 532 563
rect 526 558 532 559
rect 794 563 800 564
rect 794 559 795 563
rect 799 562 800 563
rect 1006 563 1012 564
rect 1006 562 1007 563
rect 799 560 1007 562
rect 799 559 800 560
rect 794 558 800 559
rect 1006 559 1007 560
rect 1011 559 1012 563
rect 1102 563 1103 567
rect 1107 566 1108 567
rect 1222 567 1228 568
rect 1222 566 1223 567
rect 1107 564 1223 566
rect 1107 563 1108 564
rect 1102 562 1108 563
rect 1222 563 1223 564
rect 1227 563 1228 567
rect 1222 562 1228 563
rect 1006 558 1012 559
rect 292 552 342 554
rect 79 551 85 552
rect 79 547 80 551
rect 84 550 85 551
rect 292 550 294 552
rect 84 548 294 550
rect 340 550 342 552
rect 767 551 773 552
rect 767 550 768 551
rect 340 548 518 550
rect 84 547 85 548
rect 79 546 85 547
rect 516 546 518 548
rect 652 548 768 550
rect 652 546 654 548
rect 767 547 768 548
rect 772 547 773 551
rect 767 546 773 547
rect 516 544 654 546
rect 246 540 252 541
rect 166 536 172 537
rect 134 535 140 536
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 134 531 135 535
rect 139 531 140 535
rect 166 532 167 536
rect 171 532 172 536
rect 246 536 247 540
rect 251 536 252 540
rect 470 540 476 541
rect 246 535 252 536
rect 302 538 308 539
rect 302 534 303 538
rect 307 534 308 538
rect 302 533 308 534
rect 390 536 396 537
rect 166 531 172 532
rect 390 532 391 536
rect 395 532 396 536
rect 470 536 471 540
rect 475 536 476 540
rect 726 540 732 541
rect 470 535 476 536
rect 646 536 652 537
rect 390 531 396 532
rect 534 532 540 533
rect 646 532 647 536
rect 651 532 652 536
rect 726 536 727 540
rect 731 536 732 540
rect 870 540 876 541
rect 726 535 732 536
rect 774 536 780 537
rect 134 530 140 531
rect 110 528 116 529
rect 534 528 535 532
rect 539 528 540 532
rect 151 527 157 528
rect 151 523 152 527
rect 156 526 157 527
rect 159 527 165 528
rect 159 526 160 527
rect 156 524 160 526
rect 156 523 157 524
rect 151 522 157 523
rect 159 523 160 524
rect 164 523 165 527
rect 234 527 240 528
rect 234 526 235 527
rect 229 524 235 526
rect 159 522 165 523
rect 234 523 235 524
rect 239 523 240 527
rect 458 527 464 528
rect 534 527 540 528
rect 631 531 640 532
rect 646 531 652 532
rect 774 532 775 536
rect 779 532 780 536
rect 870 536 871 540
rect 875 536 876 540
rect 1030 540 1036 541
rect 870 535 876 536
rect 926 536 932 537
rect 774 531 780 532
rect 926 532 927 536
rect 931 532 932 536
rect 1030 536 1031 540
rect 1035 536 1036 540
rect 1198 540 1204 541
rect 1030 535 1036 536
rect 1094 536 1100 537
rect 926 531 932 532
rect 1094 532 1095 536
rect 1099 532 1100 536
rect 1198 536 1199 540
rect 1203 536 1204 540
rect 1198 535 1204 536
rect 1422 535 1428 536
rect 1094 531 1100 532
rect 1286 532 1292 533
rect 631 527 632 531
rect 639 527 640 531
rect 1286 528 1287 532
rect 1291 528 1292 532
rect 458 526 459 527
rect 453 524 459 526
rect 234 522 240 523
rect 458 523 459 524
rect 463 523 464 527
rect 631 526 640 527
rect 714 527 720 528
rect 714 526 715 527
rect 709 524 715 526
rect 458 522 464 523
rect 714 523 715 524
rect 719 523 720 527
rect 842 527 848 528
rect 842 526 843 527
rect 837 524 843 526
rect 714 522 720 523
rect 842 523 843 524
rect 847 523 848 527
rect 842 522 848 523
rect 918 527 924 528
rect 918 523 919 527
rect 923 526 924 527
rect 1190 527 1196 528
rect 1286 527 1292 528
rect 1378 531 1389 532
rect 1378 527 1379 531
rect 1383 527 1384 531
rect 1388 527 1389 531
rect 1422 531 1423 535
rect 1427 531 1428 535
rect 1422 530 1428 531
rect 1478 535 1484 536
rect 1478 531 1479 535
rect 1483 531 1484 535
rect 1478 530 1484 531
rect 1526 535 1532 536
rect 1526 531 1527 535
rect 1531 531 1532 535
rect 1526 530 1532 531
rect 1574 535 1580 536
rect 1574 531 1575 535
rect 1579 531 1580 535
rect 1574 530 1580 531
rect 1622 535 1628 536
rect 1622 531 1623 535
rect 1627 531 1628 535
rect 1622 530 1628 531
rect 1654 535 1660 536
rect 1654 531 1655 535
rect 1659 531 1660 535
rect 1654 530 1660 531
rect 1694 533 1700 534
rect 1694 529 1695 533
rect 1699 529 1700 533
rect 1694 528 1700 529
rect 1190 526 1191 527
rect 923 524 945 526
rect 1157 524 1191 526
rect 923 523 924 524
rect 918 522 924 523
rect 1190 523 1191 524
rect 1195 523 1196 527
rect 1378 526 1389 527
rect 1434 527 1445 528
rect 1190 522 1196 523
rect 1434 523 1435 527
rect 1439 523 1440 527
rect 1444 523 1445 527
rect 1495 527 1501 528
rect 1495 526 1496 527
rect 1434 522 1445 523
rect 1468 524 1496 526
rect 271 519 280 520
rect 134 518 140 519
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 134 514 135 518
rect 139 514 140 518
rect 271 515 272 519
rect 279 515 280 519
rect 271 514 280 515
rect 495 519 504 520
rect 495 515 496 519
rect 503 515 504 519
rect 746 519 757 520
rect 495 514 504 515
rect 506 517 512 518
rect 134 513 140 514
rect 506 513 507 517
rect 511 513 512 517
rect 746 515 747 519
rect 751 515 752 519
rect 756 515 757 519
rect 746 514 757 515
rect 834 519 840 520
rect 834 515 835 519
rect 839 518 840 519
rect 895 519 901 520
rect 895 518 896 519
rect 839 516 896 518
rect 839 515 840 516
rect 834 514 840 515
rect 895 515 896 516
rect 900 515 901 519
rect 895 514 901 515
rect 1054 519 1061 520
rect 1054 515 1055 519
rect 1060 515 1061 519
rect 1054 514 1061 515
rect 1154 519 1160 520
rect 1154 515 1155 519
rect 1159 518 1160 519
rect 1223 519 1229 520
rect 1223 518 1224 519
rect 1159 516 1224 518
rect 1159 515 1160 516
rect 1154 514 1160 515
rect 1223 515 1224 516
rect 1228 515 1229 519
rect 1422 518 1428 519
rect 1223 514 1229 515
rect 1258 517 1264 518
rect 506 512 512 513
rect 1258 513 1259 517
rect 1263 513 1264 517
rect 1422 514 1423 518
rect 1427 514 1428 518
rect 1422 513 1428 514
rect 1258 512 1264 513
rect 110 511 116 512
rect 150 511 157 512
rect 150 507 151 511
rect 156 507 157 511
rect 1439 511 1445 512
rect 150 506 157 507
rect 294 507 300 508
rect 294 503 295 507
rect 299 503 300 507
rect 631 507 637 508
rect 294 502 300 503
rect 610 503 616 504
rect 610 502 611 503
rect 440 500 611 502
rect 174 498 180 499
rect 398 498 404 499
rect 174 494 175 498
rect 179 494 180 498
rect 302 497 308 498
rect 174 493 180 494
rect 246 493 252 494
rect 246 489 247 493
rect 251 489 252 493
rect 302 493 303 497
rect 307 493 308 497
rect 398 494 399 498
rect 403 494 404 498
rect 440 494 442 500
rect 610 499 611 500
rect 615 499 616 503
rect 631 503 632 507
rect 636 506 637 507
rect 766 507 772 508
rect 766 506 767 507
rect 636 504 767 506
rect 636 503 637 504
rect 631 502 637 503
rect 766 503 767 504
rect 771 503 772 507
rect 1222 507 1228 508
rect 1222 506 1223 507
rect 766 502 772 503
rect 1057 504 1223 506
rect 610 498 616 499
rect 654 498 660 499
rect 654 494 655 498
rect 659 494 660 498
rect 782 498 788 499
rect 782 494 783 498
rect 787 494 788 498
rect 934 498 940 499
rect 934 494 935 498
rect 939 494 940 498
rect 398 493 404 494
rect 302 492 308 493
rect 408 492 442 494
rect 470 493 476 494
rect 654 493 660 494
rect 726 493 732 494
rect 782 493 788 494
rect 870 493 876 494
rect 934 493 940 494
rect 1030 493 1036 494
rect 246 488 252 489
rect 406 491 412 492
rect 79 487 85 488
rect 79 483 80 487
rect 84 486 85 487
rect 167 487 173 488
rect 167 486 168 487
rect 84 484 168 486
rect 84 483 85 484
rect 79 482 85 483
rect 167 483 168 484
rect 172 483 173 487
rect 167 482 173 483
rect 183 487 192 488
rect 183 483 184 487
rect 191 483 192 487
rect 183 482 192 483
rect 199 487 205 488
rect 199 483 200 487
rect 204 486 205 487
rect 271 487 277 488
rect 204 484 230 486
rect 204 483 205 484
rect 199 482 205 483
rect 228 474 230 484
rect 234 483 240 484
rect 234 479 235 483
rect 239 482 240 483
rect 243 483 249 484
rect 243 482 244 483
rect 239 480 244 482
rect 239 479 240 480
rect 234 478 240 479
rect 243 479 244 480
rect 248 479 249 483
rect 271 483 272 487
rect 276 486 277 487
rect 319 487 328 488
rect 276 484 286 486
rect 276 483 277 484
rect 271 482 277 483
rect 243 478 249 479
rect 284 478 286 484
rect 319 483 320 487
rect 327 483 328 487
rect 319 482 328 483
rect 375 487 384 488
rect 375 483 376 487
rect 383 483 384 487
rect 375 482 384 483
rect 390 487 397 488
rect 390 483 391 487
rect 396 483 397 487
rect 406 487 407 491
rect 411 489 412 491
rect 470 489 471 493
rect 475 489 476 493
rect 626 491 632 492
rect 626 490 627 491
rect 411 488 413 489
rect 470 488 476 489
rect 512 488 627 490
rect 406 486 408 487
rect 407 484 408 486
rect 412 484 413 488
rect 407 483 413 484
rect 423 487 429 488
rect 423 483 424 487
rect 428 486 429 487
rect 478 487 484 488
rect 428 484 454 486
rect 428 483 429 484
rect 390 482 397 483
rect 423 482 429 483
rect 314 479 320 480
rect 314 478 315 479
rect 284 476 315 478
rect 274 475 280 476
rect 274 474 275 475
rect 228 472 275 474
rect 274 471 275 472
rect 279 471 280 475
rect 314 475 315 476
rect 319 478 320 479
rect 382 479 388 480
rect 382 478 383 479
rect 319 476 383 478
rect 319 475 320 476
rect 314 474 320 475
rect 382 475 383 476
rect 387 475 388 479
rect 382 474 388 475
rect 452 474 454 484
rect 458 483 464 484
rect 458 479 459 483
rect 463 482 464 483
rect 467 483 473 484
rect 467 482 468 483
rect 463 480 468 482
rect 463 479 464 480
rect 458 478 464 479
rect 467 479 468 480
rect 472 479 473 483
rect 478 483 479 487
rect 483 486 484 487
rect 495 487 501 488
rect 495 486 496 487
rect 483 484 496 486
rect 483 483 484 484
rect 478 482 484 483
rect 495 483 496 484
rect 500 486 501 487
rect 512 486 514 488
rect 626 487 627 488
rect 631 487 632 491
rect 726 489 727 493
rect 731 489 732 493
rect 726 488 732 489
rect 870 489 871 493
rect 875 489 876 493
rect 870 488 876 489
rect 1030 489 1031 493
rect 1035 489 1036 493
rect 1030 488 1036 489
rect 1057 488 1059 504
rect 1142 503 1148 504
rect 1142 499 1143 503
rect 1147 499 1148 503
rect 1222 503 1223 504
rect 1227 503 1228 507
rect 1439 507 1440 511
rect 1444 510 1445 511
rect 1468 510 1470 524
rect 1495 523 1496 524
rect 1500 523 1501 527
rect 1543 527 1549 528
rect 1543 526 1544 527
rect 1495 522 1501 523
rect 1520 524 1544 526
rect 1478 518 1484 519
rect 1478 514 1479 518
rect 1483 514 1484 518
rect 1478 513 1484 514
rect 1444 508 1470 510
rect 1495 511 1501 512
rect 1444 507 1445 508
rect 1439 506 1445 507
rect 1495 507 1496 511
rect 1500 510 1501 511
rect 1520 510 1522 524
rect 1543 523 1544 524
rect 1548 523 1549 527
rect 1591 527 1597 528
rect 1591 526 1592 527
rect 1543 522 1549 523
rect 1568 524 1592 526
rect 1526 518 1532 519
rect 1526 514 1527 518
rect 1531 514 1532 518
rect 1526 513 1532 514
rect 1500 508 1522 510
rect 1543 511 1549 512
rect 1500 507 1501 508
rect 1495 506 1501 507
rect 1543 507 1544 511
rect 1548 510 1549 511
rect 1568 510 1570 524
rect 1591 523 1592 524
rect 1596 523 1597 527
rect 1591 522 1597 523
rect 1606 527 1612 528
rect 1606 523 1607 527
rect 1611 526 1612 527
rect 1639 527 1645 528
rect 1639 526 1640 527
rect 1611 524 1640 526
rect 1611 523 1612 524
rect 1606 522 1612 523
rect 1639 523 1640 524
rect 1644 523 1645 527
rect 1671 527 1677 528
rect 1671 526 1672 527
rect 1639 522 1645 523
rect 1664 524 1672 526
rect 1574 518 1580 519
rect 1574 514 1575 518
rect 1579 514 1580 518
rect 1574 513 1580 514
rect 1622 518 1628 519
rect 1622 514 1623 518
rect 1627 514 1628 518
rect 1622 513 1628 514
rect 1654 518 1660 519
rect 1654 514 1655 518
rect 1659 514 1660 518
rect 1654 513 1660 514
rect 1548 508 1570 510
rect 1582 511 1588 512
rect 1548 507 1549 508
rect 1543 506 1549 507
rect 1582 507 1583 511
rect 1587 510 1588 511
rect 1591 511 1597 512
rect 1591 510 1592 511
rect 1587 508 1592 510
rect 1587 507 1588 508
rect 1582 506 1588 507
rect 1591 507 1592 508
rect 1596 507 1597 511
rect 1591 506 1597 507
rect 1639 511 1645 512
rect 1639 507 1640 511
rect 1644 510 1645 511
rect 1664 510 1666 524
rect 1671 523 1672 524
rect 1676 523 1677 527
rect 1671 522 1677 523
rect 1694 516 1700 517
rect 1694 512 1695 516
rect 1699 512 1700 516
rect 1644 508 1666 510
rect 1670 511 1677 512
rect 1694 511 1700 512
rect 1644 507 1645 508
rect 1639 506 1645 507
rect 1670 507 1671 511
rect 1676 507 1677 511
rect 1670 506 1677 507
rect 1222 502 1228 503
rect 1102 498 1108 499
rect 1142 498 1148 499
rect 1102 494 1103 498
rect 1107 494 1108 498
rect 1102 493 1108 494
rect 1198 493 1204 494
rect 1198 489 1199 493
rect 1203 489 1204 493
rect 1198 488 1204 489
rect 626 486 632 487
rect 642 487 653 488
rect 500 484 514 486
rect 500 483 501 484
rect 495 482 501 483
rect 566 483 572 484
rect 467 478 473 479
rect 566 479 567 483
rect 571 479 572 483
rect 642 483 643 487
rect 647 483 648 487
rect 652 483 653 487
rect 642 482 653 483
rect 663 487 672 488
rect 663 483 664 487
rect 671 483 672 487
rect 663 482 672 483
rect 679 487 685 488
rect 679 483 680 487
rect 684 486 685 487
rect 734 487 740 488
rect 684 484 710 486
rect 684 483 685 484
rect 679 482 685 483
rect 566 478 572 479
rect 498 475 504 476
rect 498 474 499 475
rect 452 472 499 474
rect 274 470 280 471
rect 498 471 499 472
rect 503 474 504 475
rect 708 474 710 484
rect 714 483 720 484
rect 714 479 715 483
rect 719 482 720 483
rect 723 483 729 484
rect 723 482 724 483
rect 719 480 724 482
rect 719 479 720 480
rect 714 478 720 479
rect 723 479 724 480
rect 728 479 729 483
rect 734 483 735 487
rect 739 486 740 487
rect 751 487 757 488
rect 751 486 752 487
rect 739 484 752 486
rect 739 483 740 484
rect 734 482 740 483
rect 751 483 752 484
rect 756 483 757 487
rect 751 482 757 483
rect 767 487 773 488
rect 767 483 768 487
rect 772 486 773 487
rect 775 487 781 488
rect 775 486 776 487
rect 772 484 776 486
rect 772 483 773 484
rect 767 482 773 483
rect 775 483 776 484
rect 780 483 781 487
rect 775 482 781 483
rect 791 487 800 488
rect 791 483 792 487
rect 799 483 800 487
rect 791 482 800 483
rect 806 487 813 488
rect 806 483 807 487
rect 812 486 813 487
rect 834 487 840 488
rect 834 486 835 487
rect 812 484 835 486
rect 812 483 813 484
rect 806 482 813 483
rect 834 483 835 484
rect 839 483 840 487
rect 895 487 901 488
rect 834 482 840 483
rect 842 483 848 484
rect 723 478 729 479
rect 842 479 843 483
rect 847 482 848 483
rect 867 483 873 484
rect 867 482 868 483
rect 847 480 868 482
rect 847 479 848 480
rect 842 478 848 479
rect 867 479 868 480
rect 872 479 873 483
rect 895 483 896 487
rect 900 483 901 487
rect 895 482 901 483
rect 903 487 909 488
rect 903 483 904 487
rect 908 486 909 487
rect 927 487 933 488
rect 927 486 928 487
rect 908 484 928 486
rect 908 483 909 484
rect 903 482 909 483
rect 927 483 928 484
rect 932 483 933 487
rect 927 482 933 483
rect 942 487 949 488
rect 942 483 943 487
rect 948 483 949 487
rect 942 482 949 483
rect 958 487 965 488
rect 958 483 959 487
rect 964 483 965 487
rect 1055 487 1061 488
rect 1055 486 1056 487
rect 1049 484 1056 486
rect 958 482 965 483
rect 1002 483 1008 484
rect 867 478 873 479
rect 746 475 752 476
rect 746 474 747 475
rect 503 472 525 474
rect 708 472 747 474
rect 503 471 504 472
rect 498 470 504 471
rect 746 471 747 472
rect 751 471 752 475
rect 896 474 898 482
rect 1002 479 1003 483
rect 1007 482 1008 483
rect 1027 483 1033 484
rect 1027 482 1028 483
rect 1007 480 1028 482
rect 1007 479 1008 480
rect 1002 478 1008 479
rect 1027 479 1028 480
rect 1032 479 1033 483
rect 1027 478 1033 479
rect 950 475 956 476
rect 950 474 951 475
rect 896 472 951 474
rect 746 470 752 471
rect 950 471 951 472
rect 955 474 956 475
rect 1049 474 1051 484
rect 1055 483 1056 484
rect 1060 483 1061 487
rect 1095 487 1101 488
rect 1095 486 1096 487
rect 1055 482 1061 483
rect 1064 484 1096 486
rect 1054 479 1060 480
rect 1054 475 1055 479
rect 1059 478 1060 479
rect 1064 478 1066 484
rect 1095 483 1096 484
rect 1100 483 1101 487
rect 1095 482 1101 483
rect 1110 487 1117 488
rect 1110 483 1111 487
rect 1116 483 1117 487
rect 1110 482 1117 483
rect 1127 487 1133 488
rect 1127 483 1128 487
rect 1132 486 1133 487
rect 1154 487 1160 488
rect 1154 486 1155 487
rect 1132 484 1155 486
rect 1132 483 1133 484
rect 1127 482 1133 483
rect 1154 483 1155 484
rect 1159 483 1160 487
rect 1222 487 1229 488
rect 1154 482 1160 483
rect 1190 483 1201 484
rect 1190 479 1191 483
rect 1195 479 1196 483
rect 1200 479 1201 483
rect 1222 483 1223 487
rect 1228 483 1229 487
rect 1222 482 1229 483
rect 1190 478 1201 479
rect 1214 479 1220 480
rect 1059 476 1066 478
rect 1059 475 1060 476
rect 1054 474 1060 475
rect 1214 475 1215 479
rect 1219 478 1220 479
rect 1272 478 1274 481
rect 1219 476 1274 478
rect 1219 475 1220 476
rect 1214 474 1220 475
rect 1346 475 1352 476
rect 955 472 1051 474
rect 955 471 956 472
rect 950 470 956 471
rect 1346 471 1347 475
rect 1351 471 1352 475
rect 1346 470 1352 471
rect 274 467 280 468
rect 274 463 275 467
rect 279 466 280 467
rect 610 467 616 468
rect 279 464 513 466
rect 279 463 280 464
rect 274 462 280 463
rect 610 463 611 467
rect 615 466 616 467
rect 666 467 672 468
rect 666 466 667 467
rect 615 464 667 466
rect 615 463 616 464
rect 610 462 616 463
rect 666 463 667 464
rect 671 466 672 467
rect 794 467 800 468
rect 794 466 795 467
rect 671 464 795 466
rect 671 463 672 464
rect 666 462 672 463
rect 794 463 795 464
rect 799 463 800 467
rect 794 462 800 463
rect 1230 467 1236 468
rect 1230 463 1231 467
rect 1235 466 1236 467
rect 1235 464 1265 466
rect 1235 463 1236 464
rect 1230 462 1236 463
rect 186 459 192 460
rect 186 455 187 459
rect 191 458 192 459
rect 406 459 412 460
rect 406 458 407 459
rect 191 456 407 458
rect 191 455 192 456
rect 186 454 192 455
rect 406 455 407 456
rect 411 455 412 459
rect 406 454 412 455
rect 534 459 540 460
rect 534 455 535 459
rect 539 458 540 459
rect 1042 459 1048 460
rect 1042 458 1043 459
rect 539 456 1043 458
rect 539 455 540 456
rect 534 454 540 455
rect 1042 455 1043 456
rect 1047 455 1048 459
rect 1042 454 1048 455
rect 322 451 328 452
rect 322 447 323 451
rect 327 450 328 451
rect 606 451 612 452
rect 606 450 607 451
rect 327 448 607 450
rect 327 447 328 448
rect 322 446 328 447
rect 606 447 607 448
rect 611 450 612 451
rect 686 451 692 452
rect 686 450 687 451
rect 611 448 687 450
rect 611 447 612 448
rect 606 446 612 447
rect 686 447 687 448
rect 691 447 692 451
rect 686 446 692 447
rect 1086 451 1092 452
rect 1086 447 1087 451
rect 1091 450 1092 451
rect 1747 451 1753 452
rect 1747 450 1748 451
rect 1091 448 1748 450
rect 1091 447 1092 448
rect 1086 446 1092 447
rect 1747 447 1748 448
rect 1752 447 1753 451
rect 1747 446 1753 447
rect 550 443 556 444
rect 550 439 551 443
rect 555 442 556 443
rect 942 443 948 444
rect 942 442 943 443
rect 555 440 943 442
rect 555 439 556 440
rect 550 438 556 439
rect 942 439 943 440
rect 947 442 948 443
rect 958 443 964 444
rect 958 442 959 443
rect 947 440 959 442
rect 947 439 948 440
rect 942 438 948 439
rect 958 439 959 440
rect 963 439 964 443
rect 958 438 964 439
rect 678 435 684 436
rect 678 431 679 435
rect 683 434 684 435
rect 903 435 909 436
rect 903 434 904 435
rect 683 432 904 434
rect 683 431 684 432
rect 678 430 684 431
rect 903 431 904 432
rect 908 431 909 435
rect 903 430 909 431
rect 922 435 928 436
rect 922 431 923 435
rect 927 434 928 435
rect 1330 435 1336 436
rect 1330 434 1331 435
rect 927 432 1331 434
rect 927 431 928 432
rect 922 430 928 431
rect 1330 431 1331 432
rect 1335 431 1336 435
rect 1330 430 1336 431
rect 806 427 812 428
rect 279 423 285 424
rect 279 419 280 423
rect 284 422 285 423
rect 310 423 316 424
rect 310 422 311 423
rect 284 420 311 422
rect 284 419 285 420
rect 279 418 285 419
rect 310 419 311 420
rect 315 422 316 423
rect 550 423 556 424
rect 550 422 551 423
rect 315 420 551 422
rect 315 419 316 420
rect 310 418 316 419
rect 550 419 551 420
rect 555 419 556 423
rect 806 423 807 427
rect 811 423 812 427
rect 1175 427 1181 428
rect 1175 426 1176 427
rect 1173 424 1176 426
rect 806 422 812 423
rect 1175 423 1176 424
rect 1180 423 1181 427
rect 1175 422 1181 423
rect 1190 423 1196 424
rect 550 418 556 419
rect 1190 419 1191 423
rect 1195 422 1196 423
rect 1266 423 1272 424
rect 1266 422 1267 423
rect 1195 420 1267 422
rect 1195 419 1196 420
rect 1190 418 1196 419
rect 1266 419 1267 420
rect 1271 422 1272 423
rect 1338 423 1344 424
rect 1338 422 1339 423
rect 1271 420 1339 422
rect 1271 419 1272 420
rect 1266 418 1272 419
rect 1338 419 1339 420
rect 1343 419 1344 423
rect 1338 418 1344 419
rect 768 416 773 418
rect 390 415 396 416
rect 390 414 391 415
rect 348 412 391 414
rect 79 403 85 404
rect 79 399 80 403
rect 84 402 85 403
rect 294 403 301 404
rect 294 402 295 403
rect 84 400 295 402
rect 84 399 85 400
rect 79 398 85 399
rect 294 399 295 400
rect 300 399 301 403
rect 294 398 301 399
rect 310 403 317 404
rect 310 399 311 403
rect 316 399 317 403
rect 310 398 317 399
rect 327 403 333 404
rect 327 399 328 403
rect 332 402 333 403
rect 348 402 350 412
rect 390 411 391 412
rect 395 411 396 415
rect 642 415 648 416
rect 642 414 643 415
rect 390 410 396 411
rect 569 412 643 414
rect 354 407 360 408
rect 354 403 355 407
rect 359 406 360 407
rect 371 407 377 408
rect 371 406 372 407
rect 359 404 372 406
rect 359 403 360 404
rect 354 402 360 403
rect 371 403 372 404
rect 376 403 377 407
rect 371 402 377 403
rect 382 407 388 408
rect 382 403 383 407
rect 387 406 388 407
rect 478 407 484 408
rect 478 406 479 407
rect 387 404 479 406
rect 387 403 388 404
rect 382 402 388 403
rect 399 403 405 404
rect 332 400 350 402
rect 332 399 333 400
rect 327 398 333 399
rect 374 399 380 400
rect 374 395 375 399
rect 379 395 380 399
rect 399 399 400 403
rect 404 399 405 403
rect 478 403 479 404
rect 483 403 484 407
rect 569 404 571 412
rect 642 411 643 412
rect 647 411 648 415
rect 746 415 752 416
rect 642 410 648 411
rect 734 411 740 412
rect 734 410 735 411
rect 652 408 735 410
rect 594 407 600 408
rect 478 402 484 403
rect 526 403 532 404
rect 399 398 405 399
rect 526 399 527 403
rect 531 402 532 403
rect 535 403 541 404
rect 535 402 536 403
rect 531 400 536 402
rect 531 399 532 400
rect 526 398 532 399
rect 535 399 536 400
rect 540 399 541 403
rect 535 398 541 399
rect 550 403 557 404
rect 550 399 551 403
rect 556 399 557 403
rect 550 398 557 399
rect 567 403 573 404
rect 567 399 568 403
rect 572 399 573 403
rect 594 403 595 407
rect 599 406 600 407
rect 611 407 617 408
rect 611 406 612 407
rect 599 404 612 406
rect 599 403 600 404
rect 594 402 600 403
rect 611 403 612 404
rect 616 403 617 407
rect 611 402 617 403
rect 626 403 632 404
rect 567 398 573 399
rect 614 399 620 400
rect 614 395 615 399
rect 619 395 620 399
rect 626 399 627 403
rect 631 402 632 403
rect 639 403 645 404
rect 639 402 640 403
rect 631 400 640 402
rect 631 399 632 400
rect 626 398 632 399
rect 639 399 640 400
rect 644 402 645 403
rect 652 402 654 408
rect 734 407 735 408
rect 739 407 740 411
rect 746 411 747 415
rect 751 414 752 415
rect 768 414 770 416
rect 751 412 770 414
rect 1162 415 1168 416
rect 751 411 752 412
rect 746 410 752 411
rect 882 411 888 412
rect 734 406 740 407
rect 766 407 772 408
rect 644 400 654 402
rect 686 403 693 404
rect 644 399 645 400
rect 639 398 645 399
rect 686 399 687 403
rect 692 399 693 403
rect 686 398 693 399
rect 718 403 724 404
rect 718 399 719 403
rect 723 402 724 403
rect 743 403 749 404
rect 743 402 744 403
rect 723 400 744 402
rect 723 399 724 400
rect 718 398 724 399
rect 743 399 744 400
rect 748 399 749 403
rect 766 403 767 407
rect 771 403 772 407
rect 882 407 883 411
rect 887 410 888 411
rect 1162 411 1163 415
rect 1167 411 1168 415
rect 1162 410 1168 411
rect 1174 415 1180 416
rect 1174 411 1175 415
rect 1179 414 1180 415
rect 1366 415 1372 416
rect 1366 414 1367 415
rect 1179 412 1367 414
rect 1179 411 1180 412
rect 1174 410 1180 411
rect 1366 411 1367 412
rect 1371 411 1372 415
rect 1366 410 1372 411
rect 887 408 1089 410
rect 887 407 888 408
rect 882 406 888 407
rect 1378 407 1384 408
rect 1378 406 1379 407
rect 1305 404 1379 406
rect 766 402 772 403
rect 935 403 941 404
rect 743 398 749 399
rect 935 399 936 403
rect 940 402 941 403
rect 943 403 949 404
rect 943 402 944 403
rect 940 400 944 402
rect 940 399 941 400
rect 935 398 941 399
rect 943 399 944 400
rect 948 399 949 403
rect 943 398 949 399
rect 958 403 965 404
rect 958 399 959 403
rect 964 399 965 403
rect 958 398 965 399
rect 975 403 981 404
rect 975 399 976 403
rect 980 402 981 403
rect 1054 403 1060 404
rect 1054 402 1055 403
rect 980 400 1055 402
rect 980 399 981 400
rect 975 398 981 399
rect 1054 399 1055 400
rect 1059 399 1060 403
rect 1054 398 1060 399
rect 1062 403 1068 404
rect 1062 399 1063 403
rect 1067 402 1068 403
rect 1247 403 1253 404
rect 1247 402 1248 403
rect 1067 400 1248 402
rect 1067 399 1068 400
rect 1062 398 1068 399
rect 1126 399 1132 400
rect 302 394 308 395
rect 374 394 380 395
rect 542 394 548 395
rect 614 394 620 395
rect 670 395 676 396
rect 1126 395 1127 399
rect 1131 395 1132 399
rect 1247 399 1248 400
rect 1252 399 1253 403
rect 1247 398 1253 399
rect 1303 403 1309 404
rect 1303 399 1304 403
rect 1308 399 1309 403
rect 1378 403 1379 404
rect 1383 403 1384 407
rect 1378 402 1384 403
rect 1303 398 1309 399
rect 1351 399 1357 400
rect 1351 398 1352 399
rect 1324 396 1352 398
rect 302 390 303 394
rect 307 390 308 394
rect 534 391 540 392
rect 534 390 535 391
rect 302 389 308 390
rect 487 389 535 390
rect 487 386 488 389
rect 465 385 488 386
rect 492 388 535 389
rect 492 385 493 388
rect 534 387 535 388
rect 539 387 540 391
rect 542 390 543 394
rect 547 390 548 394
rect 670 391 671 395
rect 675 391 676 395
rect 670 390 676 391
rect 950 394 956 395
rect 1126 394 1132 395
rect 1230 395 1236 396
rect 950 390 951 394
rect 955 390 956 394
rect 1230 391 1231 395
rect 1235 391 1236 395
rect 1230 390 1236 391
rect 542 389 548 390
rect 950 389 956 390
rect 534 386 540 387
rect 1031 387 1037 388
rect 465 384 493 385
rect 159 383 165 384
rect 159 382 160 383
rect 153 380 160 382
rect 151 379 157 380
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 151 375 152 379
rect 156 375 157 379
rect 159 379 160 380
rect 164 379 165 383
rect 192 380 219 382
rect 249 380 274 382
rect 433 380 458 382
rect 465 380 467 384
rect 879 383 888 384
rect 159 378 165 379
rect 183 379 189 380
rect 183 378 184 379
rect 176 376 184 378
rect 110 371 116 372
rect 134 374 140 375
rect 151 374 157 375
rect 166 374 172 375
rect 134 370 135 374
rect 139 370 140 374
rect 134 369 140 370
rect 166 370 167 374
rect 171 370 172 374
rect 166 369 172 370
rect 176 364 178 376
rect 183 375 184 376
rect 188 375 189 379
rect 183 374 189 375
rect 151 363 157 364
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 151 359 152 363
rect 156 362 157 363
rect 164 362 178 364
rect 183 363 189 364
rect 156 360 166 362
rect 156 359 157 360
rect 151 358 157 359
rect 183 359 184 363
rect 188 362 189 363
rect 192 362 194 380
rect 215 379 221 380
rect 215 375 216 379
rect 220 375 221 379
rect 247 379 253 380
rect 247 375 248 379
rect 252 375 253 379
rect 198 374 204 375
rect 215 374 221 375
rect 230 374 236 375
rect 247 374 253 375
rect 262 374 268 375
rect 198 370 199 374
rect 203 370 204 374
rect 198 369 204 370
rect 230 370 231 374
rect 235 370 236 374
rect 230 369 236 370
rect 262 370 263 374
rect 267 370 268 374
rect 262 369 268 370
rect 188 360 194 362
rect 215 363 221 364
rect 188 359 189 360
rect 183 358 189 359
rect 215 359 216 363
rect 220 359 221 363
rect 215 358 221 359
rect 247 363 253 364
rect 247 359 248 363
rect 252 359 253 363
rect 272 362 274 380
rect 279 379 285 380
rect 279 375 280 379
rect 284 378 285 379
rect 287 379 293 380
rect 287 378 288 379
rect 284 376 288 378
rect 284 375 285 376
rect 279 374 285 375
rect 287 375 288 376
rect 292 375 293 379
rect 431 379 437 380
rect 431 375 432 379
rect 436 375 437 379
rect 287 374 293 375
rect 414 374 420 375
rect 431 374 437 375
rect 446 374 452 375
rect 390 371 396 372
rect 354 367 360 368
rect 279 363 285 364
rect 279 362 280 363
rect 272 360 280 362
rect 247 358 253 359
rect 279 359 280 360
rect 284 359 285 363
rect 354 363 355 367
rect 359 363 360 367
rect 390 367 391 371
rect 395 370 396 371
rect 399 371 405 372
rect 399 370 400 371
rect 395 368 400 370
rect 395 367 396 368
rect 390 366 396 367
rect 399 367 400 368
rect 404 367 405 371
rect 414 370 415 374
rect 419 370 420 374
rect 414 369 420 370
rect 446 370 447 374
rect 451 370 452 374
rect 446 369 452 370
rect 399 366 405 367
rect 354 362 360 363
rect 430 363 437 364
rect 279 358 285 359
rect 430 359 431 363
rect 436 359 437 363
rect 456 362 458 380
rect 463 379 469 380
rect 463 375 464 379
rect 468 375 469 379
rect 518 379 525 380
rect 463 374 469 375
rect 486 377 492 378
rect 486 373 487 377
rect 491 373 492 377
rect 518 375 519 379
rect 524 375 525 379
rect 664 378 666 381
rect 879 379 880 383
rect 887 379 888 383
rect 1031 383 1032 387
rect 1036 386 1037 387
rect 1190 387 1196 388
rect 1190 386 1191 387
rect 1036 384 1191 386
rect 1036 383 1037 384
rect 1031 382 1037 383
rect 1190 383 1191 384
rect 1195 383 1196 387
rect 1214 387 1220 388
rect 1214 386 1215 387
rect 1190 382 1196 383
rect 1199 385 1215 386
rect 1199 381 1200 385
rect 1204 384 1215 385
rect 1204 381 1205 384
rect 1214 383 1215 384
rect 1219 383 1220 387
rect 1324 386 1326 396
rect 1351 395 1352 396
rect 1356 395 1357 399
rect 1351 394 1357 395
rect 1366 399 1373 400
rect 1366 395 1367 399
rect 1372 395 1373 399
rect 1366 394 1373 395
rect 1387 399 1393 400
rect 1387 395 1388 399
rect 1392 398 1393 399
rect 1454 399 1460 400
rect 1454 398 1455 399
rect 1392 396 1455 398
rect 1392 395 1393 396
rect 1387 394 1393 395
rect 1454 395 1455 396
rect 1459 395 1460 399
rect 1454 394 1460 395
rect 1281 384 1326 386
rect 1358 389 1364 390
rect 1358 385 1359 389
rect 1363 385 1364 389
rect 1358 384 1364 385
rect 1214 382 1220 383
rect 1503 383 1509 384
rect 1199 380 1205 381
rect 879 378 888 379
rect 919 379 928 380
rect 518 374 525 375
rect 596 376 666 378
rect 486 372 492 373
rect 596 372 598 376
rect 754 375 760 376
rect 919 375 920 379
rect 927 375 928 379
rect 1062 379 1069 380
rect 526 371 532 372
rect 526 367 527 371
rect 531 370 532 371
rect 588 370 598 372
rect 639 371 648 372
rect 531 368 590 370
rect 531 367 532 368
rect 526 366 532 367
rect 594 367 600 368
rect 463 363 469 364
rect 463 362 464 363
rect 456 360 464 362
rect 430 358 437 359
rect 463 359 464 360
rect 468 359 469 363
rect 594 363 595 367
rect 599 363 600 367
rect 639 367 640 371
rect 647 367 648 371
rect 754 371 755 375
rect 759 371 760 375
rect 754 370 760 371
rect 902 374 908 375
rect 919 374 928 375
rect 1030 377 1036 378
rect 902 370 903 374
rect 907 370 908 374
rect 1030 373 1031 377
rect 1035 373 1036 377
rect 1062 375 1063 379
rect 1068 375 1069 379
rect 1335 379 1344 380
rect 1062 374 1069 375
rect 1074 375 1080 376
rect 1335 375 1336 379
rect 1343 375 1344 379
rect 1030 372 1036 373
rect 1074 371 1075 375
rect 1079 371 1080 375
rect 1074 370 1080 371
rect 1318 374 1324 375
rect 1335 374 1344 375
rect 1438 379 1444 380
rect 1438 375 1439 379
rect 1443 375 1444 379
rect 1494 379 1501 380
rect 1494 375 1495 379
rect 1500 375 1501 379
rect 1503 379 1504 383
rect 1508 382 1509 383
rect 1543 383 1549 384
rect 1508 380 1539 382
rect 1508 379 1509 380
rect 1503 378 1509 379
rect 1535 379 1541 380
rect 1535 375 1536 379
rect 1540 375 1541 379
rect 1543 379 1544 383
rect 1548 382 1549 383
rect 1548 380 1579 382
rect 1616 380 1643 382
rect 1648 380 1675 382
rect 1548 379 1549 380
rect 1543 378 1549 379
rect 1575 379 1581 380
rect 1575 375 1576 379
rect 1580 375 1581 379
rect 1606 379 1613 380
rect 1606 375 1607 379
rect 1612 375 1613 379
rect 1438 374 1444 375
rect 1478 374 1484 375
rect 1494 374 1501 375
rect 1518 374 1524 375
rect 1535 374 1541 375
rect 1558 374 1564 375
rect 1575 374 1581 375
rect 1590 374 1596 375
rect 1606 374 1613 375
rect 1318 370 1319 374
rect 1323 370 1324 374
rect 902 369 908 370
rect 1318 369 1324 370
rect 1330 371 1336 372
rect 639 366 648 367
rect 1002 367 1008 368
rect 594 362 600 363
rect 918 363 925 364
rect 463 358 469 359
rect 782 360 788 361
rect 110 354 116 355
rect 134 357 140 358
rect 134 353 135 357
rect 139 353 140 357
rect 134 352 140 353
rect 166 357 172 358
rect 166 353 167 357
rect 171 353 172 357
rect 166 352 172 353
rect 198 357 204 358
rect 198 353 199 357
rect 203 353 204 357
rect 198 352 204 353
rect 154 351 160 352
rect 154 347 155 351
rect 159 350 160 351
rect 217 350 219 358
rect 230 357 236 358
rect 230 353 231 357
rect 235 353 236 357
rect 230 352 236 353
rect 262 357 268 358
rect 414 357 420 358
rect 262 353 263 357
rect 267 353 268 357
rect 262 352 268 353
rect 294 356 300 357
rect 294 352 295 356
rect 299 352 300 356
rect 414 353 415 357
rect 419 353 420 357
rect 294 351 300 352
rect 374 352 380 353
rect 414 352 420 353
rect 446 357 452 358
rect 446 353 447 357
rect 451 353 452 357
rect 446 352 452 353
rect 534 356 540 357
rect 534 352 535 356
rect 539 352 540 356
rect 782 356 783 360
rect 787 356 788 360
rect 782 355 788 356
rect 878 359 885 360
rect 878 355 879 359
rect 884 355 885 359
rect 918 359 919 363
rect 924 359 925 363
rect 1002 363 1003 367
rect 1007 363 1008 367
rect 1330 367 1331 371
rect 1335 370 1336 371
rect 1478 370 1479 374
rect 1483 370 1484 374
rect 1335 368 1377 370
rect 1478 369 1484 370
rect 1518 370 1519 374
rect 1523 370 1524 374
rect 1518 369 1524 370
rect 1558 370 1559 374
rect 1563 370 1564 374
rect 1558 369 1564 370
rect 1590 370 1591 374
rect 1595 370 1596 374
rect 1590 369 1596 370
rect 1335 367 1336 368
rect 1330 366 1336 367
rect 1002 362 1008 363
rect 1334 363 1341 364
rect 918 358 925 359
rect 1102 360 1108 361
rect 670 354 676 355
rect 878 354 885 355
rect 902 357 908 358
rect 159 348 219 350
rect 374 348 375 352
rect 379 348 380 352
rect 534 351 540 352
rect 614 352 620 353
rect 159 347 160 348
rect 374 347 380 348
rect 502 350 508 351
rect 154 346 160 347
rect 502 346 503 350
rect 507 346 508 350
rect 614 348 615 352
rect 619 348 620 352
rect 670 350 671 354
rect 675 350 676 354
rect 902 353 903 357
rect 907 353 908 357
rect 902 352 908 353
rect 942 356 948 357
rect 942 352 943 356
rect 947 352 948 356
rect 1102 356 1103 360
rect 1107 356 1108 360
rect 1102 355 1108 356
rect 1194 359 1205 360
rect 1194 355 1195 359
rect 1199 355 1200 359
rect 1204 355 1205 359
rect 1334 359 1335 363
rect 1340 359 1341 363
rect 1495 363 1501 364
rect 1334 358 1341 359
rect 1454 359 1461 360
rect 1318 357 1324 358
rect 1194 354 1205 355
rect 1230 354 1236 355
rect 942 351 948 352
rect 670 349 676 350
rect 1046 350 1052 351
rect 614 347 620 348
rect 502 345 508 346
rect 1046 346 1047 350
rect 1051 346 1052 350
rect 1230 350 1231 354
rect 1235 350 1236 354
rect 1318 353 1319 357
rect 1323 353 1324 357
rect 1318 352 1324 353
rect 1438 356 1444 357
rect 1438 352 1439 356
rect 1443 352 1444 356
rect 1454 355 1455 359
rect 1460 355 1461 359
rect 1495 359 1496 363
rect 1500 362 1501 363
rect 1503 363 1509 364
rect 1503 362 1504 363
rect 1500 360 1504 362
rect 1500 359 1501 360
rect 1495 358 1501 359
rect 1503 359 1504 360
rect 1508 359 1509 363
rect 1503 358 1509 359
rect 1535 363 1541 364
rect 1535 359 1536 363
rect 1540 362 1541 363
rect 1543 363 1549 364
rect 1543 362 1544 363
rect 1540 360 1544 362
rect 1540 359 1541 360
rect 1535 358 1541 359
rect 1543 359 1544 360
rect 1548 359 1549 363
rect 1543 358 1549 359
rect 1575 363 1581 364
rect 1575 359 1576 363
rect 1580 359 1581 363
rect 1575 358 1581 359
rect 1607 363 1613 364
rect 1607 359 1608 363
rect 1612 362 1613 363
rect 1616 362 1618 380
rect 1639 379 1645 380
rect 1639 375 1640 379
rect 1644 375 1645 379
rect 1622 374 1628 375
rect 1639 374 1645 375
rect 1622 370 1623 374
rect 1627 370 1628 374
rect 1622 369 1628 370
rect 1612 360 1618 362
rect 1639 363 1645 364
rect 1612 359 1613 360
rect 1607 358 1613 359
rect 1639 359 1640 363
rect 1644 362 1645 363
rect 1648 362 1650 380
rect 1671 379 1677 380
rect 1671 375 1672 379
rect 1676 375 1677 379
rect 1654 374 1660 375
rect 1671 374 1677 375
rect 1694 376 1700 377
rect 1654 370 1655 374
rect 1659 370 1660 374
rect 1694 372 1695 376
rect 1699 372 1700 376
rect 1694 371 1700 372
rect 1654 369 1660 370
rect 1644 360 1650 362
rect 1671 363 1677 364
rect 1644 359 1645 360
rect 1639 358 1645 359
rect 1671 359 1672 363
rect 1676 359 1677 363
rect 1671 358 1677 359
rect 1694 359 1700 360
rect 1454 354 1461 355
rect 1478 357 1484 358
rect 1478 353 1479 357
rect 1483 353 1484 357
rect 1478 352 1484 353
rect 1518 357 1524 358
rect 1518 353 1519 357
rect 1523 353 1524 357
rect 1518 352 1524 353
rect 1558 357 1564 358
rect 1558 353 1559 357
rect 1563 353 1564 357
rect 1558 352 1564 353
rect 1590 357 1596 358
rect 1590 353 1591 357
rect 1595 353 1596 357
rect 1590 352 1596 353
rect 1622 357 1628 358
rect 1622 353 1623 357
rect 1627 353 1628 357
rect 1622 352 1628 353
rect 1654 357 1660 358
rect 1654 353 1655 357
rect 1659 353 1660 357
rect 1654 352 1660 353
rect 1438 351 1444 352
rect 1642 351 1648 352
rect 1230 349 1236 350
rect 1350 349 1356 350
rect 1046 345 1052 346
rect 1350 345 1351 349
rect 1355 345 1356 349
rect 1642 347 1643 351
rect 1647 350 1648 351
rect 1673 350 1675 358
rect 1694 355 1695 359
rect 1699 355 1700 359
rect 1694 354 1700 355
rect 1647 348 1675 350
rect 1647 347 1648 348
rect 1642 346 1648 347
rect 1350 344 1356 345
rect 479 343 485 344
rect 479 339 480 343
rect 484 342 485 343
rect 1023 343 1029 344
rect 484 340 530 342
rect 484 339 485 340
rect 479 338 485 339
rect 528 338 530 340
rect 566 339 572 340
rect 566 338 567 339
rect 528 336 567 338
rect 566 335 567 336
rect 571 335 572 339
rect 1023 339 1024 343
rect 1028 342 1029 343
rect 1038 343 1044 344
rect 1038 342 1039 343
rect 1028 340 1039 342
rect 1028 339 1029 340
rect 1023 338 1029 339
rect 1038 339 1039 340
rect 1043 339 1044 343
rect 1038 338 1044 339
rect 566 334 572 335
rect 518 331 524 332
rect 518 327 519 331
rect 523 330 524 331
rect 710 331 716 332
rect 710 330 711 331
rect 523 328 711 330
rect 523 327 524 328
rect 518 326 524 327
rect 710 327 711 328
rect 715 327 716 331
rect 710 326 716 327
rect 935 323 941 324
rect 935 319 936 323
rect 940 322 941 323
rect 982 323 988 324
rect 982 322 983 323
rect 940 320 983 322
rect 940 319 941 320
rect 935 318 941 319
rect 982 319 983 320
rect 987 319 988 323
rect 982 318 988 319
rect 1174 319 1180 320
rect 1174 315 1175 319
rect 1179 318 1180 319
rect 1214 319 1220 320
rect 1214 318 1215 319
rect 1179 316 1215 318
rect 1179 315 1180 316
rect 1174 314 1180 315
rect 1214 315 1215 316
rect 1219 315 1220 319
rect 1214 314 1220 315
rect 1198 311 1204 312
rect 1198 307 1199 311
rect 1203 307 1204 311
rect 598 306 604 307
rect 134 303 140 304
rect 110 301 116 302
rect 110 297 111 301
rect 115 297 116 301
rect 134 299 135 303
rect 139 299 140 303
rect 134 298 140 299
rect 166 303 172 304
rect 166 299 167 303
rect 171 299 172 303
rect 166 298 172 299
rect 198 303 204 304
rect 198 299 199 303
rect 203 299 204 303
rect 198 298 204 299
rect 230 303 236 304
rect 230 299 231 303
rect 235 299 236 303
rect 230 298 236 299
rect 262 303 268 304
rect 262 299 263 303
rect 267 299 268 303
rect 262 298 268 299
rect 294 303 300 304
rect 294 299 295 303
rect 299 299 300 303
rect 294 298 300 299
rect 326 303 332 304
rect 326 299 327 303
rect 331 299 332 303
rect 326 298 332 299
rect 358 303 364 304
rect 358 299 359 303
rect 363 299 364 303
rect 358 298 364 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 422 303 428 304
rect 422 299 423 303
rect 427 299 428 303
rect 422 298 428 299
rect 454 303 460 304
rect 454 299 455 303
rect 459 299 460 303
rect 454 298 460 299
rect 486 303 492 304
rect 486 299 487 303
rect 491 299 492 303
rect 486 298 492 299
rect 518 303 524 304
rect 518 299 519 303
rect 523 299 524 303
rect 518 298 524 299
rect 550 303 556 304
rect 550 299 551 303
rect 555 299 556 303
rect 598 302 599 306
rect 603 302 604 306
rect 598 301 604 302
rect 702 306 708 307
rect 702 302 703 306
rect 707 302 708 306
rect 702 301 708 302
rect 806 306 812 307
rect 806 302 807 306
rect 811 302 812 306
rect 806 301 812 302
rect 910 306 916 307
rect 910 302 911 306
rect 915 302 916 306
rect 1110 306 1116 307
rect 1198 306 1204 307
rect 1494 311 1500 312
rect 1494 307 1495 311
rect 1499 310 1500 311
rect 1499 308 1579 310
rect 1499 307 1500 308
rect 1494 306 1500 307
rect 910 301 916 302
rect 998 303 1004 304
rect 550 298 556 299
rect 998 299 999 303
rect 1003 299 1004 303
rect 998 298 1004 299
rect 1030 303 1036 304
rect 1030 299 1031 303
rect 1035 299 1036 303
rect 1030 298 1036 299
rect 1062 303 1068 304
rect 1062 299 1063 303
rect 1067 299 1068 303
rect 1110 302 1111 306
rect 1115 302 1116 306
rect 1286 304 1292 305
rect 1110 301 1116 302
rect 1062 298 1068 299
rect 1192 300 1217 302
rect 1286 300 1287 304
rect 1291 300 1292 304
rect 1318 303 1324 304
rect 110 296 116 297
rect 151 295 157 296
rect 151 291 152 295
rect 156 294 157 295
rect 183 295 189 296
rect 156 292 178 294
rect 156 291 157 292
rect 151 290 157 291
rect 134 286 140 287
rect 110 284 116 285
rect 79 283 88 284
rect 79 279 80 283
rect 87 279 88 283
rect 110 280 111 284
rect 115 280 116 284
rect 134 282 135 286
rect 139 282 140 286
rect 134 281 140 282
rect 166 286 172 287
rect 166 282 167 286
rect 171 282 172 286
rect 166 281 172 282
rect 110 279 116 280
rect 151 279 160 280
rect 79 278 88 279
rect 151 275 152 279
rect 159 275 160 279
rect 176 278 178 292
rect 183 291 184 295
rect 188 294 189 295
rect 215 295 221 296
rect 188 292 210 294
rect 188 291 189 292
rect 183 290 189 291
rect 198 286 204 287
rect 198 282 199 286
rect 203 282 204 286
rect 198 281 204 282
rect 183 279 189 280
rect 183 278 184 279
rect 176 276 184 278
rect 151 274 160 275
rect 183 275 184 276
rect 188 275 189 279
rect 208 278 210 292
rect 215 291 216 295
rect 220 294 221 295
rect 247 295 253 296
rect 220 292 242 294
rect 220 291 221 292
rect 215 290 221 291
rect 230 286 236 287
rect 230 282 231 286
rect 235 282 236 286
rect 230 281 236 282
rect 215 279 221 280
rect 215 278 216 279
rect 208 276 216 278
rect 183 274 189 275
rect 215 275 216 276
rect 220 275 221 279
rect 240 278 242 292
rect 247 291 248 295
rect 252 294 253 295
rect 274 295 285 296
rect 252 292 259 294
rect 252 291 253 292
rect 247 290 253 291
rect 247 279 253 280
rect 247 278 248 279
rect 240 276 248 278
rect 215 274 221 275
rect 247 275 248 276
rect 252 275 253 279
rect 257 278 259 292
rect 274 291 275 295
rect 279 291 280 295
rect 284 291 285 295
rect 274 290 285 291
rect 287 295 293 296
rect 287 291 288 295
rect 292 294 293 295
rect 311 295 317 296
rect 311 294 312 295
rect 292 292 312 294
rect 292 291 293 292
rect 287 290 293 291
rect 311 291 312 292
rect 316 291 317 295
rect 343 295 349 296
rect 343 294 344 295
rect 311 290 317 291
rect 319 292 344 294
rect 262 286 268 287
rect 262 282 263 286
rect 267 282 268 286
rect 262 281 268 282
rect 294 286 300 287
rect 294 282 295 286
rect 299 282 300 286
rect 294 281 300 282
rect 279 279 285 280
rect 279 278 280 279
rect 257 276 280 278
rect 247 274 253 275
rect 279 275 280 276
rect 284 275 285 279
rect 279 274 285 275
rect 311 279 317 280
rect 311 275 312 279
rect 316 278 317 279
rect 319 278 321 292
rect 343 291 344 292
rect 348 291 349 295
rect 375 295 381 296
rect 375 294 376 295
rect 343 290 349 291
rect 352 292 376 294
rect 326 286 332 287
rect 326 282 327 286
rect 331 282 332 286
rect 326 281 332 282
rect 316 276 321 278
rect 343 279 349 280
rect 316 275 317 276
rect 311 274 317 275
rect 343 275 344 279
rect 348 278 349 279
rect 352 278 354 292
rect 375 291 376 292
rect 380 291 381 295
rect 375 290 381 291
rect 407 295 413 296
rect 407 291 408 295
rect 412 294 413 295
rect 439 295 445 296
rect 412 292 434 294
rect 412 291 413 292
rect 407 290 413 291
rect 358 286 364 287
rect 358 282 359 286
rect 363 282 364 286
rect 358 281 364 282
rect 390 286 396 287
rect 390 282 391 286
rect 395 282 396 286
rect 390 281 396 282
rect 422 286 428 287
rect 422 282 423 286
rect 427 282 428 286
rect 432 286 434 292
rect 439 291 440 295
rect 444 294 445 295
rect 471 295 477 296
rect 444 292 466 294
rect 444 291 445 292
rect 439 290 445 291
rect 454 286 460 287
rect 432 284 443 286
rect 422 281 428 282
rect 441 280 443 284
rect 454 282 455 286
rect 459 282 460 286
rect 454 281 460 282
rect 348 276 354 278
rect 366 279 372 280
rect 348 275 349 276
rect 343 274 349 275
rect 366 275 367 279
rect 371 278 372 279
rect 375 279 381 280
rect 375 278 376 279
rect 371 276 376 278
rect 371 275 372 276
rect 366 274 372 275
rect 375 275 376 276
rect 380 275 381 279
rect 375 274 381 275
rect 407 279 413 280
rect 407 275 408 279
rect 412 278 413 279
rect 430 279 436 280
rect 430 278 431 279
rect 412 276 431 278
rect 412 275 413 276
rect 407 274 413 275
rect 430 275 431 276
rect 435 275 436 279
rect 430 274 436 275
rect 439 279 445 280
rect 439 275 440 279
rect 444 275 445 279
rect 464 278 466 292
rect 471 291 472 295
rect 476 294 477 295
rect 503 295 509 296
rect 476 292 498 294
rect 476 291 477 292
rect 471 290 477 291
rect 486 286 492 287
rect 486 282 487 286
rect 491 282 492 286
rect 486 281 492 282
rect 471 279 477 280
rect 471 278 472 279
rect 464 276 472 278
rect 439 274 445 275
rect 471 275 472 276
rect 476 275 477 279
rect 496 278 498 292
rect 503 291 504 295
rect 508 291 509 295
rect 503 290 509 291
rect 530 295 541 296
rect 530 291 531 295
rect 535 291 536 295
rect 540 291 541 295
rect 530 290 541 291
rect 566 295 573 296
rect 566 291 567 295
rect 572 291 573 295
rect 566 290 573 291
rect 778 295 784 296
rect 778 291 779 295
rect 783 294 784 295
rect 918 295 924 296
rect 918 294 919 295
rect 783 292 919 294
rect 783 291 784 292
rect 778 290 784 291
rect 918 291 919 292
rect 923 291 924 295
rect 918 290 924 291
rect 1015 295 1021 296
rect 1015 291 1016 295
rect 1020 291 1021 295
rect 1015 290 1021 291
rect 1042 295 1053 296
rect 1042 291 1043 295
rect 1047 291 1048 295
rect 1052 291 1053 295
rect 1042 290 1053 291
rect 1055 295 1061 296
rect 1055 291 1056 295
rect 1060 294 1061 295
rect 1079 295 1085 296
rect 1079 294 1080 295
rect 1060 292 1080 294
rect 1060 291 1061 292
rect 1055 290 1061 291
rect 1079 291 1080 292
rect 1084 291 1085 295
rect 1192 294 1194 300
rect 1286 299 1292 300
rect 1298 299 1309 300
rect 1298 295 1299 299
rect 1303 295 1304 299
rect 1308 295 1309 299
rect 1318 299 1319 303
rect 1323 299 1324 303
rect 1318 298 1324 299
rect 1350 303 1356 304
rect 1350 299 1351 303
rect 1355 299 1356 303
rect 1350 298 1356 299
rect 1382 303 1388 304
rect 1382 299 1383 303
rect 1387 299 1388 303
rect 1382 298 1388 299
rect 1414 303 1420 304
rect 1414 299 1415 303
rect 1419 299 1420 303
rect 1414 298 1420 299
rect 1446 303 1452 304
rect 1446 299 1447 303
rect 1451 299 1452 303
rect 1446 298 1452 299
rect 1478 303 1484 304
rect 1478 299 1479 303
rect 1483 299 1484 303
rect 1478 298 1484 299
rect 1518 303 1524 304
rect 1518 299 1519 303
rect 1523 299 1524 303
rect 1518 298 1524 299
rect 1558 303 1564 304
rect 1558 299 1559 303
rect 1563 299 1564 303
rect 1558 298 1564 299
rect 1577 296 1579 308
rect 1590 303 1596 304
rect 1590 299 1591 303
rect 1595 299 1596 303
rect 1590 298 1596 299
rect 1622 303 1628 304
rect 1622 299 1623 303
rect 1627 299 1628 303
rect 1622 298 1628 299
rect 1654 303 1660 304
rect 1654 299 1655 303
rect 1659 299 1660 303
rect 1654 298 1660 299
rect 1694 301 1700 302
rect 1694 297 1695 301
rect 1699 297 1700 301
rect 1694 296 1700 297
rect 1298 294 1309 295
rect 1335 295 1341 296
rect 1079 290 1085 291
rect 1096 292 1194 294
rect 505 286 507 290
rect 518 286 524 287
rect 505 284 514 286
rect 503 279 509 280
rect 503 278 504 279
rect 496 276 504 278
rect 471 274 477 275
rect 503 275 504 276
rect 508 275 509 279
rect 512 278 514 284
rect 518 282 519 286
rect 523 282 524 286
rect 518 281 524 282
rect 550 286 556 287
rect 550 282 551 286
rect 555 282 556 286
rect 550 281 556 282
rect 998 286 1004 287
rect 998 282 999 286
rect 1003 282 1004 286
rect 1017 286 1019 290
rect 1030 286 1036 287
rect 1017 284 1026 286
rect 998 281 1004 282
rect 535 279 541 280
rect 535 278 536 279
rect 512 276 536 278
rect 503 274 509 275
rect 535 275 536 276
rect 540 275 541 279
rect 535 274 541 275
rect 567 279 573 280
rect 567 275 568 279
rect 572 278 573 279
rect 582 279 588 280
rect 582 278 583 279
rect 572 276 583 278
rect 572 275 573 276
rect 567 274 573 275
rect 582 275 583 276
rect 587 275 588 279
rect 1015 279 1021 280
rect 582 274 588 275
rect 622 275 628 276
rect 622 271 623 275
rect 627 271 628 275
rect 622 270 628 271
rect 830 275 836 276
rect 830 271 831 275
rect 835 271 836 275
rect 982 275 988 276
rect 982 274 983 275
rect 961 272 983 274
rect 830 270 836 271
rect 982 271 983 272
rect 987 274 988 275
rect 1006 275 1012 276
rect 1006 274 1007 275
rect 987 272 1007 274
rect 987 271 988 272
rect 982 270 988 271
rect 1006 271 1007 272
rect 1011 271 1012 275
rect 1015 275 1016 279
rect 1020 275 1021 279
rect 1024 278 1026 284
rect 1030 282 1031 286
rect 1035 282 1036 286
rect 1030 281 1036 282
rect 1062 286 1068 287
rect 1062 282 1063 286
rect 1067 282 1068 286
rect 1062 281 1068 282
rect 1047 279 1053 280
rect 1047 278 1048 279
rect 1024 276 1048 278
rect 1015 274 1021 275
rect 1047 275 1048 276
rect 1052 275 1053 279
rect 1047 274 1053 275
rect 1079 279 1085 280
rect 1079 275 1080 279
rect 1084 278 1085 279
rect 1096 278 1098 292
rect 1335 291 1336 295
rect 1340 294 1341 295
rect 1367 295 1373 296
rect 1340 292 1362 294
rect 1340 291 1341 292
rect 1335 290 1341 291
rect 1318 286 1324 287
rect 1318 282 1319 286
rect 1323 282 1324 286
rect 1084 276 1098 278
rect 1286 281 1292 282
rect 1318 281 1324 282
rect 1350 286 1356 287
rect 1350 282 1351 286
rect 1355 282 1356 286
rect 1350 281 1356 282
rect 1286 277 1287 281
rect 1291 277 1292 281
rect 1286 276 1292 277
rect 1334 279 1341 280
rect 1084 275 1085 276
rect 1079 274 1085 275
rect 1334 275 1335 279
rect 1340 275 1341 279
rect 1360 278 1362 292
rect 1367 291 1368 295
rect 1372 294 1373 295
rect 1399 295 1405 296
rect 1372 292 1394 294
rect 1372 291 1373 292
rect 1367 290 1373 291
rect 1382 286 1388 287
rect 1382 282 1383 286
rect 1387 282 1388 286
rect 1382 281 1388 282
rect 1367 279 1373 280
rect 1367 278 1368 279
rect 1360 276 1368 278
rect 1334 274 1341 275
rect 1367 275 1368 276
rect 1372 275 1373 279
rect 1392 278 1394 292
rect 1399 291 1400 295
rect 1404 294 1405 295
rect 1431 295 1437 296
rect 1404 292 1426 294
rect 1404 291 1405 292
rect 1399 290 1405 291
rect 1414 286 1420 287
rect 1414 282 1415 286
rect 1419 282 1420 286
rect 1414 281 1420 282
rect 1399 279 1405 280
rect 1399 278 1400 279
rect 1392 276 1400 278
rect 1367 274 1373 275
rect 1399 275 1400 276
rect 1404 275 1405 279
rect 1424 278 1426 292
rect 1431 291 1432 295
rect 1436 294 1437 295
rect 1463 295 1469 296
rect 1436 292 1458 294
rect 1436 291 1437 292
rect 1431 290 1437 291
rect 1446 286 1452 287
rect 1446 282 1447 286
rect 1451 282 1452 286
rect 1446 281 1452 282
rect 1431 279 1437 280
rect 1431 278 1432 279
rect 1424 276 1432 278
rect 1399 274 1405 275
rect 1431 275 1432 276
rect 1436 275 1437 279
rect 1456 278 1458 292
rect 1463 291 1464 295
rect 1468 294 1469 295
rect 1495 295 1501 296
rect 1468 292 1490 294
rect 1468 291 1469 292
rect 1463 290 1469 291
rect 1478 286 1484 287
rect 1478 282 1479 286
rect 1483 282 1484 286
rect 1478 281 1484 282
rect 1463 279 1469 280
rect 1463 278 1464 279
rect 1456 276 1464 278
rect 1431 274 1437 275
rect 1463 275 1464 276
rect 1468 275 1469 279
rect 1488 278 1490 292
rect 1495 291 1496 295
rect 1500 294 1501 295
rect 1530 295 1541 296
rect 1500 292 1514 294
rect 1500 291 1501 292
rect 1495 290 1501 291
rect 1495 279 1501 280
rect 1495 278 1496 279
rect 1488 276 1496 278
rect 1463 274 1469 275
rect 1495 275 1496 276
rect 1500 275 1501 279
rect 1512 278 1514 292
rect 1530 291 1531 295
rect 1535 291 1536 295
rect 1540 291 1541 295
rect 1530 290 1541 291
rect 1575 295 1581 296
rect 1575 291 1576 295
rect 1580 291 1581 295
rect 1607 295 1613 296
rect 1607 294 1608 295
rect 1575 290 1581 291
rect 1600 292 1608 294
rect 1518 286 1524 287
rect 1518 282 1519 286
rect 1523 282 1524 286
rect 1518 281 1524 282
rect 1558 286 1564 287
rect 1558 282 1559 286
rect 1563 282 1564 286
rect 1558 281 1564 282
rect 1590 286 1596 287
rect 1590 282 1591 286
rect 1595 282 1596 286
rect 1590 281 1596 282
rect 1535 279 1541 280
rect 1535 278 1536 279
rect 1512 276 1536 278
rect 1495 274 1501 275
rect 1535 275 1536 276
rect 1540 275 1541 279
rect 1535 274 1541 275
rect 1575 279 1581 280
rect 1575 275 1576 279
rect 1580 278 1581 279
rect 1600 278 1602 292
rect 1607 291 1608 292
rect 1612 291 1613 295
rect 1607 290 1613 291
rect 1639 295 1645 296
rect 1639 291 1640 295
rect 1644 294 1645 295
rect 1670 295 1677 296
rect 1644 292 1666 294
rect 1644 291 1645 292
rect 1639 290 1645 291
rect 1622 286 1628 287
rect 1622 282 1623 286
rect 1627 282 1628 286
rect 1622 281 1628 282
rect 1654 286 1660 287
rect 1654 282 1655 286
rect 1659 282 1660 286
rect 1654 281 1660 282
rect 1580 276 1602 278
rect 1606 279 1613 280
rect 1580 275 1581 276
rect 1575 274 1581 275
rect 1606 275 1607 279
rect 1612 275 1613 279
rect 1606 274 1613 275
rect 1639 279 1648 280
rect 1639 275 1640 279
rect 1647 275 1648 279
rect 1664 278 1666 292
rect 1670 291 1671 295
rect 1676 291 1677 295
rect 1670 290 1677 291
rect 1722 291 1728 292
rect 1722 287 1723 291
rect 1727 290 1728 291
rect 1747 291 1753 292
rect 1747 290 1748 291
rect 1727 288 1748 290
rect 1727 287 1728 288
rect 1722 286 1728 287
rect 1747 287 1748 288
rect 1752 287 1753 291
rect 1747 286 1753 287
rect 1694 284 1700 285
rect 1694 280 1695 284
rect 1699 280 1700 284
rect 1671 279 1677 280
rect 1694 279 1700 280
rect 1671 278 1672 279
rect 1664 276 1672 278
rect 1639 274 1648 275
rect 1671 275 1672 276
rect 1676 275 1677 279
rect 1671 274 1677 275
rect 1006 270 1012 271
rect 1017 270 1019 274
rect 1161 272 1194 274
rect 1082 271 1088 272
rect 1082 270 1083 271
rect 1017 268 1083 270
rect 1082 267 1083 268
rect 1087 267 1088 271
rect 1082 266 1088 267
rect 598 265 604 266
rect 598 261 599 265
rect 603 261 604 265
rect 598 260 604 261
rect 702 265 708 266
rect 702 261 703 265
rect 707 261 708 265
rect 806 265 812 266
rect 702 260 708 261
rect 769 260 790 262
rect 806 261 807 265
rect 811 261 812 265
rect 806 260 812 261
rect 910 265 916 266
rect 910 261 911 265
rect 915 261 916 265
rect 910 260 916 261
rect 1110 265 1116 266
rect 1110 261 1111 265
rect 1115 261 1116 265
rect 1110 260 1116 261
rect 606 255 612 256
rect 606 251 607 255
rect 611 254 612 255
rect 615 255 621 256
rect 615 254 616 255
rect 611 252 616 254
rect 611 251 612 252
rect 606 250 612 251
rect 615 251 616 252
rect 620 251 621 255
rect 615 250 621 251
rect 671 255 677 256
rect 671 251 672 255
rect 676 254 677 255
rect 687 255 693 256
rect 687 254 688 255
rect 676 252 688 254
rect 676 251 677 252
rect 671 250 677 251
rect 687 251 688 252
rect 692 251 693 255
rect 687 250 693 251
rect 710 255 716 256
rect 710 251 711 255
rect 715 254 716 255
rect 719 255 725 256
rect 719 254 720 255
rect 715 252 720 254
rect 715 251 716 252
rect 710 250 716 251
rect 719 251 720 252
rect 724 254 725 255
rect 769 254 771 260
rect 724 252 771 254
rect 775 255 784 256
rect 724 251 725 252
rect 719 250 725 251
rect 775 251 776 255
rect 783 251 784 255
rect 775 250 784 251
rect 622 247 628 248
rect 622 243 623 247
rect 627 246 628 247
rect 670 247 676 248
rect 670 246 671 247
rect 627 244 671 246
rect 627 243 628 244
rect 622 242 628 243
rect 670 243 671 244
rect 675 243 676 247
rect 670 242 676 243
rect 711 243 717 244
rect 711 239 712 243
rect 716 242 717 243
rect 720 242 722 250
rect 788 246 790 260
rect 1182 259 1188 260
rect 822 255 829 256
rect 822 251 823 255
rect 828 251 829 255
rect 822 250 829 251
rect 878 255 885 256
rect 878 251 879 255
rect 884 251 885 255
rect 878 250 885 251
rect 926 255 933 256
rect 926 251 927 255
rect 932 251 933 255
rect 926 250 933 251
rect 982 255 989 256
rect 982 251 983 255
rect 988 251 989 255
rect 1126 255 1133 256
rect 982 250 989 251
rect 1006 251 1012 252
rect 1006 247 1007 251
rect 1011 250 1012 251
rect 1118 251 1124 252
rect 1118 250 1119 251
rect 1011 248 1119 250
rect 1011 247 1012 248
rect 1006 246 1012 247
rect 1118 247 1119 248
rect 1123 247 1124 251
rect 1126 251 1127 255
rect 1132 251 1133 255
rect 1182 255 1183 259
rect 1187 256 1188 259
rect 1192 258 1194 272
rect 1206 271 1212 272
rect 1206 267 1207 271
rect 1211 267 1212 271
rect 1206 266 1212 267
rect 1199 259 1205 260
rect 1199 258 1200 259
rect 1192 256 1200 258
rect 1187 255 1189 256
rect 1182 254 1184 255
rect 1126 250 1133 251
rect 1183 251 1184 254
rect 1188 251 1189 255
rect 1199 255 1200 256
rect 1204 255 1205 259
rect 1199 254 1205 255
rect 1214 259 1221 260
rect 1214 255 1215 259
rect 1220 255 1221 259
rect 1214 254 1221 255
rect 1235 259 1241 260
rect 1235 255 1236 259
rect 1240 258 1241 259
rect 1298 259 1304 260
rect 1298 258 1299 259
rect 1240 256 1299 258
rect 1240 255 1241 256
rect 1235 254 1241 255
rect 1298 255 1299 256
rect 1303 255 1304 259
rect 1298 254 1304 255
rect 1183 250 1189 251
rect 1118 246 1124 247
rect 788 244 987 246
rect 716 240 722 242
rect 767 243 773 244
rect 716 239 717 240
rect 711 238 717 239
rect 767 239 768 243
rect 772 242 773 243
rect 983 243 989 244
rect 772 240 810 242
rect 772 239 773 240
rect 767 238 773 239
rect 806 239 812 240
rect 694 235 700 236
rect 582 231 588 232
rect 270 227 276 228
rect 270 226 271 227
rect 208 224 271 226
rect 199 219 205 220
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 199 215 200 219
rect 204 218 205 219
rect 208 218 210 224
rect 270 223 271 224
rect 275 223 276 227
rect 270 222 276 223
rect 330 227 336 228
rect 330 223 331 227
rect 335 226 336 227
rect 582 227 583 231
rect 587 230 588 231
rect 654 231 660 232
rect 654 230 655 231
rect 587 228 655 230
rect 587 227 588 228
rect 582 226 588 227
rect 654 227 655 228
rect 659 227 660 231
rect 694 231 695 235
rect 699 231 700 235
rect 806 235 807 239
rect 811 235 812 239
rect 806 234 812 235
rect 830 239 837 240
rect 830 235 831 239
rect 836 235 837 239
rect 830 234 837 235
rect 847 239 856 240
rect 847 235 848 239
rect 855 235 856 239
rect 847 234 856 235
rect 867 239 873 240
rect 867 235 868 239
rect 872 238 873 239
rect 934 239 940 240
rect 934 238 935 239
rect 872 236 935 238
rect 872 235 873 236
rect 867 234 873 235
rect 934 235 935 236
rect 939 235 940 239
rect 983 239 984 243
rect 988 239 989 243
rect 983 238 989 239
rect 1039 243 1045 244
rect 1039 239 1040 243
rect 1044 242 1045 243
rect 1055 243 1061 244
rect 1055 242 1056 243
rect 1044 240 1056 242
rect 1044 239 1045 240
rect 1039 238 1045 239
rect 1055 239 1056 240
rect 1060 239 1061 243
rect 1055 238 1061 239
rect 934 234 940 235
rect 966 235 972 236
rect 694 230 700 231
rect 966 231 967 235
rect 971 231 972 235
rect 966 230 972 231
rect 1198 231 1204 232
rect 1198 230 1199 231
rect 654 226 660 227
rect 838 229 844 230
rect 335 224 386 226
rect 838 225 839 229
rect 843 225 844 229
rect 1159 228 1199 230
rect 1159 226 1161 228
rect 1198 227 1199 228
rect 1203 227 1204 231
rect 1530 231 1536 232
rect 1530 230 1531 231
rect 1198 226 1204 227
rect 1320 228 1531 230
rect 838 224 844 225
rect 1136 224 1161 226
rect 335 223 336 224
rect 330 222 336 223
rect 231 219 237 220
rect 231 218 232 219
rect 204 216 210 218
rect 224 216 232 218
rect 204 215 205 216
rect 110 211 116 212
rect 182 214 188 215
rect 199 214 205 215
rect 214 214 220 215
rect 182 210 183 214
rect 187 210 188 214
rect 182 209 188 210
rect 214 210 215 214
rect 219 210 220 214
rect 214 209 220 210
rect 224 204 226 216
rect 231 215 232 216
rect 236 215 237 219
rect 263 219 269 220
rect 263 218 264 219
rect 256 216 264 218
rect 231 214 237 215
rect 246 214 252 215
rect 246 210 247 214
rect 251 210 252 214
rect 246 209 252 210
rect 256 204 258 216
rect 263 215 264 216
rect 268 215 269 219
rect 295 219 301 220
rect 295 218 296 219
rect 288 216 296 218
rect 263 214 269 215
rect 278 214 284 215
rect 278 210 279 214
rect 283 210 284 214
rect 278 209 284 210
rect 288 204 290 216
rect 295 215 296 216
rect 300 215 301 219
rect 327 219 333 220
rect 327 218 328 219
rect 319 216 328 218
rect 295 214 301 215
rect 310 214 316 215
rect 310 210 311 214
rect 315 210 316 214
rect 310 209 316 210
rect 319 204 321 216
rect 327 215 328 216
rect 332 215 333 219
rect 358 219 365 220
rect 358 215 359 219
rect 364 215 365 219
rect 384 218 386 224
rect 718 223 724 224
rect 592 220 619 222
rect 391 219 397 220
rect 391 218 392 219
rect 384 216 392 218
rect 391 215 392 216
rect 396 215 397 219
rect 423 219 429 220
rect 423 218 424 219
rect 416 216 424 218
rect 327 214 333 215
rect 342 214 348 215
rect 358 214 365 215
rect 374 214 380 215
rect 391 214 397 215
rect 406 214 412 215
rect 342 210 343 214
rect 347 210 348 214
rect 366 211 372 212
rect 366 210 367 211
rect 342 209 348 210
rect 360 208 367 210
rect 360 204 362 208
rect 366 207 367 208
rect 371 207 372 211
rect 374 210 375 214
rect 379 210 380 214
rect 374 209 380 210
rect 406 210 407 214
rect 411 210 412 214
rect 406 209 412 210
rect 366 206 372 207
rect 416 204 418 216
rect 423 215 424 216
rect 428 215 429 219
rect 455 219 461 220
rect 455 218 456 219
rect 448 216 456 218
rect 423 214 429 215
rect 438 214 444 215
rect 438 210 439 214
rect 443 210 444 214
rect 438 209 444 210
rect 448 204 450 216
rect 455 215 456 216
rect 460 215 461 219
rect 487 219 493 220
rect 487 218 488 219
rect 480 216 488 218
rect 455 214 461 215
rect 470 214 476 215
rect 470 210 471 214
rect 475 210 476 214
rect 470 209 476 210
rect 480 204 482 216
rect 487 215 488 216
rect 492 215 493 219
rect 519 219 525 220
rect 519 215 520 219
rect 524 215 525 219
rect 551 219 557 220
rect 551 218 552 219
rect 544 216 552 218
rect 487 214 493 215
rect 502 214 508 215
rect 519 214 525 215
rect 534 214 540 215
rect 502 210 503 214
rect 507 210 508 214
rect 502 209 508 210
rect 534 210 535 214
rect 539 210 540 214
rect 534 209 540 210
rect 487 204 493 205
rect 544 204 546 216
rect 551 215 552 216
rect 556 215 557 219
rect 583 219 589 220
rect 583 218 584 219
rect 576 216 584 218
rect 551 214 557 215
rect 566 214 572 215
rect 566 210 567 214
rect 571 210 572 214
rect 566 209 572 210
rect 576 204 578 216
rect 583 215 584 216
rect 588 215 589 219
rect 583 214 589 215
rect 199 203 205 204
rect 110 199 116 200
rect 110 195 111 199
rect 115 195 116 199
rect 199 199 200 203
rect 204 202 205 203
rect 212 202 226 204
rect 231 203 237 204
rect 204 200 214 202
rect 204 199 205 200
rect 199 198 205 199
rect 231 199 232 203
rect 236 202 237 203
rect 244 202 258 204
rect 263 203 269 204
rect 236 200 246 202
rect 236 199 237 200
rect 231 198 237 199
rect 263 199 264 203
rect 268 202 269 203
rect 276 202 290 204
rect 295 203 301 204
rect 268 200 278 202
rect 268 199 269 200
rect 263 198 269 199
rect 295 199 296 203
rect 300 202 301 203
rect 308 202 321 204
rect 327 203 336 204
rect 300 200 310 202
rect 300 199 301 200
rect 295 198 301 199
rect 327 199 328 203
rect 335 199 336 203
rect 327 198 336 199
rect 359 203 365 204
rect 359 199 360 203
rect 364 199 365 203
rect 359 198 365 199
rect 391 203 397 204
rect 391 199 392 203
rect 396 202 397 203
rect 404 202 418 204
rect 423 203 429 204
rect 396 200 406 202
rect 396 199 397 200
rect 391 198 397 199
rect 423 199 424 203
rect 428 202 429 203
rect 436 202 450 204
rect 455 203 461 204
rect 428 200 438 202
rect 428 199 429 200
rect 423 198 429 199
rect 455 199 456 203
rect 460 202 461 203
rect 468 202 482 204
rect 486 203 488 204
rect 460 200 470 202
rect 460 199 461 200
rect 455 198 461 199
rect 486 199 487 203
rect 492 200 493 204
rect 491 199 493 200
rect 519 203 525 204
rect 519 199 520 203
rect 524 202 525 203
rect 532 202 546 204
rect 551 203 557 204
rect 524 200 534 202
rect 524 199 525 200
rect 486 198 492 199
rect 519 198 525 199
rect 551 199 552 203
rect 556 202 557 203
rect 564 202 578 204
rect 583 203 589 204
rect 556 200 566 202
rect 556 199 557 200
rect 551 198 557 199
rect 583 199 584 203
rect 588 202 589 203
rect 592 202 594 220
rect 615 219 621 220
rect 615 215 616 219
rect 620 215 621 219
rect 646 219 652 220
rect 646 215 647 219
rect 651 218 652 219
rect 655 219 661 220
rect 655 218 656 219
rect 651 216 656 218
rect 651 215 652 216
rect 598 214 604 215
rect 615 214 621 215
rect 638 214 644 215
rect 646 214 652 215
rect 655 215 656 216
rect 660 215 661 219
rect 718 219 719 223
rect 723 219 724 223
rect 982 223 988 224
rect 718 218 724 219
rect 807 219 813 220
rect 807 215 808 219
rect 812 218 813 219
rect 918 219 924 220
rect 812 216 830 218
rect 812 215 813 216
rect 655 214 661 215
rect 790 214 796 215
rect 807 214 813 215
rect 598 210 599 214
rect 603 210 604 214
rect 598 209 604 210
rect 638 210 639 214
rect 643 210 644 214
rect 638 209 644 210
rect 790 210 791 214
rect 795 210 796 214
rect 790 209 796 210
rect 828 210 830 216
rect 918 215 919 219
rect 923 215 924 219
rect 982 219 983 223
rect 987 219 988 223
rect 982 218 988 219
rect 1074 219 1085 220
rect 1074 215 1075 219
rect 1079 215 1080 219
rect 1084 215 1085 219
rect 1119 219 1125 220
rect 1119 215 1120 219
rect 1124 218 1125 219
rect 1136 218 1138 224
rect 1310 223 1316 224
rect 1310 222 1311 223
rect 1201 220 1234 222
rect 1296 220 1311 222
rect 1159 219 1165 220
rect 1159 218 1160 219
rect 1124 216 1138 218
rect 1152 216 1160 218
rect 1124 215 1125 216
rect 918 214 924 215
rect 1062 214 1068 215
rect 1074 214 1085 215
rect 1102 214 1108 215
rect 1119 214 1125 215
rect 1142 214 1148 215
rect 1062 210 1063 214
rect 1067 210 1068 214
rect 828 208 857 210
rect 1062 209 1068 210
rect 1102 210 1103 214
rect 1107 210 1108 214
rect 1102 209 1108 210
rect 1142 210 1143 214
rect 1147 210 1148 214
rect 1142 209 1148 210
rect 1152 204 1154 216
rect 1159 215 1160 216
rect 1164 215 1165 219
rect 1199 219 1205 220
rect 1199 215 1200 219
rect 1204 215 1205 219
rect 1159 214 1165 215
rect 1182 214 1188 215
rect 1199 214 1205 215
rect 1222 214 1228 215
rect 1182 210 1183 214
rect 1187 210 1188 214
rect 1182 209 1188 210
rect 1222 210 1223 214
rect 1227 210 1228 214
rect 1222 209 1228 210
rect 588 200 594 202
rect 614 203 621 204
rect 588 199 589 200
rect 583 198 589 199
rect 614 199 615 203
rect 620 199 621 203
rect 614 198 621 199
rect 654 203 661 204
rect 654 199 655 203
rect 660 199 661 203
rect 654 198 661 199
rect 806 203 813 204
rect 806 199 807 203
rect 812 199 813 203
rect 1079 203 1088 204
rect 806 198 813 199
rect 934 199 941 200
rect 110 194 116 195
rect 182 197 188 198
rect 182 193 183 197
rect 187 193 188 197
rect 182 192 188 193
rect 214 197 220 198
rect 214 193 215 197
rect 219 193 220 197
rect 214 192 220 193
rect 246 197 252 198
rect 246 193 247 197
rect 251 193 252 197
rect 246 192 252 193
rect 278 197 284 198
rect 278 193 279 197
rect 283 193 284 197
rect 278 192 284 193
rect 310 197 316 198
rect 310 193 311 197
rect 315 193 316 197
rect 310 192 316 193
rect 342 197 348 198
rect 342 193 343 197
rect 347 193 348 197
rect 342 192 348 193
rect 374 197 380 198
rect 374 193 375 197
rect 379 193 380 197
rect 374 192 380 193
rect 406 197 412 198
rect 406 193 407 197
rect 411 193 412 197
rect 406 192 412 193
rect 438 197 444 198
rect 438 193 439 197
rect 443 193 444 197
rect 438 192 444 193
rect 470 197 476 198
rect 470 193 471 197
rect 475 193 476 197
rect 470 192 476 193
rect 502 197 508 198
rect 502 193 503 197
rect 507 193 508 197
rect 502 192 508 193
rect 534 197 540 198
rect 534 193 535 197
rect 539 193 540 197
rect 534 192 540 193
rect 566 197 572 198
rect 566 193 567 197
rect 571 193 572 197
rect 566 192 572 193
rect 598 197 604 198
rect 598 193 599 197
rect 603 193 604 197
rect 598 192 604 193
rect 638 197 644 198
rect 638 193 639 197
rect 643 193 644 197
rect 790 197 796 198
rect 638 192 644 193
rect 694 194 700 195
rect 358 191 364 192
rect 358 187 359 191
rect 363 190 364 191
rect 486 191 492 192
rect 486 190 487 191
rect 363 188 487 190
rect 363 187 364 188
rect 358 186 364 187
rect 486 187 487 188
rect 491 187 492 191
rect 694 190 695 194
rect 699 190 700 194
rect 790 193 791 197
rect 795 193 796 197
rect 790 192 796 193
rect 918 196 924 197
rect 918 192 919 196
rect 923 192 924 196
rect 934 195 935 199
rect 940 195 941 199
rect 1079 199 1080 203
rect 1087 199 1088 203
rect 1079 198 1088 199
rect 1119 203 1125 204
rect 1119 199 1120 203
rect 1124 202 1125 203
rect 1140 202 1154 204
rect 1159 203 1168 204
rect 1124 200 1142 202
rect 1124 199 1125 200
rect 1119 198 1125 199
rect 1159 199 1160 203
rect 1167 199 1168 203
rect 1159 198 1168 199
rect 1198 203 1205 204
rect 1198 199 1199 203
rect 1204 199 1205 203
rect 1232 202 1234 220
rect 1239 219 1245 220
rect 1239 215 1240 219
rect 1244 218 1245 219
rect 1279 219 1285 220
rect 1244 216 1258 218
rect 1244 215 1245 216
rect 1239 214 1245 215
rect 1256 206 1258 216
rect 1279 215 1280 219
rect 1284 218 1285 219
rect 1296 218 1298 220
rect 1310 219 1311 220
rect 1315 219 1316 223
rect 1320 220 1322 228
rect 1530 227 1531 228
rect 1535 227 1536 231
rect 1530 226 1536 227
rect 1327 223 1333 224
rect 1310 218 1316 219
rect 1319 219 1325 220
rect 1284 216 1298 218
rect 1284 215 1285 216
rect 1319 215 1320 219
rect 1324 215 1325 219
rect 1327 219 1328 223
rect 1332 222 1333 223
rect 1463 223 1469 224
rect 1332 220 1354 222
rect 1332 219 1333 220
rect 1327 218 1333 219
rect 1352 218 1354 220
rect 1359 219 1365 220
rect 1359 218 1360 219
rect 1352 216 1360 218
rect 1359 215 1360 216
rect 1364 215 1365 219
rect 1391 219 1397 220
rect 1391 218 1392 219
rect 1384 216 1392 218
rect 1262 214 1268 215
rect 1279 214 1285 215
rect 1302 214 1308 215
rect 1319 214 1325 215
rect 1342 214 1348 215
rect 1359 214 1365 215
rect 1374 214 1380 215
rect 1262 210 1263 214
rect 1267 210 1268 214
rect 1262 209 1268 210
rect 1302 210 1303 214
rect 1307 210 1308 214
rect 1302 209 1308 210
rect 1342 210 1343 214
rect 1347 210 1348 214
rect 1342 209 1348 210
rect 1374 210 1375 214
rect 1379 210 1380 214
rect 1374 209 1380 210
rect 1256 204 1262 206
rect 1384 204 1386 216
rect 1391 215 1392 216
rect 1396 215 1397 219
rect 1423 219 1429 220
rect 1423 218 1424 219
rect 1416 216 1424 218
rect 1391 214 1397 215
rect 1406 214 1412 215
rect 1406 210 1407 214
rect 1411 210 1412 214
rect 1406 209 1412 210
rect 1416 204 1418 216
rect 1423 215 1424 216
rect 1428 215 1429 219
rect 1455 219 1461 220
rect 1455 218 1456 219
rect 1448 216 1456 218
rect 1423 214 1429 215
rect 1438 214 1444 215
rect 1438 210 1439 214
rect 1443 210 1444 214
rect 1438 209 1444 210
rect 1448 204 1450 216
rect 1455 215 1456 216
rect 1460 215 1461 219
rect 1463 219 1464 223
rect 1468 222 1469 223
rect 1503 223 1509 224
rect 1468 220 1499 222
rect 1468 219 1469 220
rect 1463 218 1469 219
rect 1495 219 1501 220
rect 1495 215 1496 219
rect 1500 215 1501 219
rect 1503 219 1504 223
rect 1508 222 1509 223
rect 1543 223 1549 224
rect 1508 220 1539 222
rect 1508 219 1509 220
rect 1503 218 1509 219
rect 1535 219 1541 220
rect 1535 215 1536 219
rect 1540 215 1541 219
rect 1543 219 1544 223
rect 1548 222 1549 223
rect 1548 220 1579 222
rect 1641 220 1666 222
rect 1548 219 1549 220
rect 1543 218 1549 219
rect 1575 219 1581 220
rect 1575 215 1576 219
rect 1580 215 1581 219
rect 1598 219 1604 220
rect 1598 215 1599 219
rect 1603 218 1604 219
rect 1607 219 1613 220
rect 1607 218 1608 219
rect 1603 216 1608 218
rect 1603 215 1604 216
rect 1455 214 1461 215
rect 1478 214 1484 215
rect 1495 214 1501 215
rect 1518 214 1524 215
rect 1535 214 1541 215
rect 1558 214 1564 215
rect 1575 214 1581 215
rect 1590 214 1596 215
rect 1598 214 1604 215
rect 1607 215 1608 216
rect 1612 215 1613 219
rect 1639 219 1645 220
rect 1639 215 1640 219
rect 1644 215 1645 219
rect 1607 214 1613 215
rect 1622 214 1628 215
rect 1639 214 1645 215
rect 1654 214 1660 215
rect 1478 210 1479 214
rect 1483 210 1484 214
rect 1478 209 1484 210
rect 1518 210 1519 214
rect 1523 210 1524 214
rect 1518 209 1524 210
rect 1558 210 1559 214
rect 1563 210 1564 214
rect 1558 209 1564 210
rect 1590 210 1591 214
rect 1595 210 1596 214
rect 1590 209 1596 210
rect 1622 210 1623 214
rect 1627 210 1628 214
rect 1622 209 1628 210
rect 1654 210 1655 214
rect 1659 210 1660 214
rect 1654 209 1660 210
rect 1239 203 1245 204
rect 1239 202 1240 203
rect 1232 200 1240 202
rect 1198 198 1205 199
rect 1239 199 1240 200
rect 1244 199 1245 203
rect 1260 202 1274 204
rect 1279 203 1285 204
rect 1279 202 1280 203
rect 1272 200 1280 202
rect 1239 198 1245 199
rect 1279 199 1280 200
rect 1284 199 1285 203
rect 1279 198 1285 199
rect 1319 203 1325 204
rect 1319 199 1320 203
rect 1324 202 1325 203
rect 1327 203 1333 204
rect 1327 202 1328 203
rect 1324 200 1328 202
rect 1324 199 1325 200
rect 1319 198 1325 199
rect 1327 199 1328 200
rect 1332 199 1333 203
rect 1327 198 1333 199
rect 1359 203 1365 204
rect 1359 199 1360 203
rect 1364 202 1365 203
rect 1372 202 1386 204
rect 1391 203 1397 204
rect 1364 200 1374 202
rect 1364 199 1365 200
rect 1359 198 1365 199
rect 1391 199 1392 203
rect 1396 202 1397 203
rect 1404 202 1418 204
rect 1423 203 1429 204
rect 1396 200 1406 202
rect 1396 199 1397 200
rect 1391 198 1397 199
rect 1423 199 1424 203
rect 1428 202 1429 203
rect 1436 202 1450 204
rect 1455 203 1461 204
rect 1428 200 1438 202
rect 1428 199 1429 200
rect 1423 198 1429 199
rect 1455 199 1456 203
rect 1460 202 1461 203
rect 1463 203 1469 204
rect 1463 202 1464 203
rect 1460 200 1464 202
rect 1460 199 1461 200
rect 1455 198 1461 199
rect 1463 199 1464 200
rect 1468 199 1469 203
rect 1463 198 1469 199
rect 1495 203 1501 204
rect 1495 199 1496 203
rect 1500 202 1501 203
rect 1503 203 1509 204
rect 1503 202 1504 203
rect 1500 200 1504 202
rect 1500 199 1501 200
rect 1495 198 1501 199
rect 1503 199 1504 200
rect 1508 199 1509 203
rect 1503 198 1509 199
rect 1535 203 1541 204
rect 1535 199 1536 203
rect 1540 202 1541 203
rect 1543 203 1549 204
rect 1543 202 1544 203
rect 1540 200 1544 202
rect 1540 199 1541 200
rect 1535 198 1541 199
rect 1543 199 1544 200
rect 1548 199 1549 203
rect 1543 198 1549 199
rect 1575 203 1584 204
rect 1575 199 1576 203
rect 1583 199 1584 203
rect 1575 198 1584 199
rect 1606 203 1613 204
rect 1606 199 1607 203
rect 1612 199 1613 203
rect 1606 198 1613 199
rect 1639 203 1648 204
rect 1639 199 1640 203
rect 1647 199 1648 203
rect 1664 202 1666 220
rect 1670 219 1677 220
rect 1670 215 1671 219
rect 1676 215 1677 219
rect 1670 214 1677 215
rect 1694 216 1700 217
rect 1694 212 1695 216
rect 1699 212 1700 216
rect 1694 211 1700 212
rect 1671 203 1677 204
rect 1671 202 1672 203
rect 1664 200 1672 202
rect 1639 198 1648 199
rect 1671 199 1672 200
rect 1676 199 1677 203
rect 1671 198 1677 199
rect 1694 199 1700 200
rect 1062 197 1068 198
rect 934 194 941 195
rect 966 194 972 195
rect 918 191 924 192
rect 966 190 967 194
rect 971 190 972 194
rect 1062 193 1063 197
rect 1067 193 1068 197
rect 1062 192 1068 193
rect 1102 197 1108 198
rect 1102 193 1103 197
rect 1107 193 1108 197
rect 1102 192 1108 193
rect 1142 197 1148 198
rect 1142 193 1143 197
rect 1147 193 1148 197
rect 1142 192 1148 193
rect 1182 197 1188 198
rect 1182 193 1183 197
rect 1187 193 1188 197
rect 1182 192 1188 193
rect 1222 197 1228 198
rect 1222 193 1223 197
rect 1227 193 1228 197
rect 1222 192 1228 193
rect 1262 197 1268 198
rect 1262 193 1263 197
rect 1267 193 1268 197
rect 1262 192 1268 193
rect 1302 197 1308 198
rect 1302 193 1303 197
rect 1307 193 1308 197
rect 1302 192 1308 193
rect 1342 197 1348 198
rect 1342 193 1343 197
rect 1347 193 1348 197
rect 1342 192 1348 193
rect 1374 197 1380 198
rect 1374 193 1375 197
rect 1379 193 1380 197
rect 1374 192 1380 193
rect 1406 197 1412 198
rect 1406 193 1407 197
rect 1411 193 1412 197
rect 1406 192 1412 193
rect 1438 197 1444 198
rect 1438 193 1439 197
rect 1443 193 1444 197
rect 1438 192 1444 193
rect 1478 197 1484 198
rect 1478 193 1479 197
rect 1483 193 1484 197
rect 1478 192 1484 193
rect 1518 197 1524 198
rect 1518 193 1519 197
rect 1523 193 1524 197
rect 1518 192 1524 193
rect 1558 197 1564 198
rect 1558 193 1559 197
rect 1563 193 1564 197
rect 1558 192 1564 193
rect 1590 197 1596 198
rect 1590 193 1591 197
rect 1595 193 1596 197
rect 1590 192 1596 193
rect 1622 197 1628 198
rect 1622 193 1623 197
rect 1627 193 1628 197
rect 1622 192 1628 193
rect 1654 197 1660 198
rect 1654 193 1655 197
rect 1659 193 1660 197
rect 1694 195 1695 199
rect 1699 195 1700 199
rect 1694 194 1700 195
rect 1654 192 1660 193
rect 694 189 700 190
rect 830 189 836 190
rect 966 189 972 190
rect 1118 191 1124 192
rect 486 186 492 187
rect 830 185 831 189
rect 835 185 836 189
rect 1118 187 1119 191
rect 1123 190 1124 191
rect 1199 191 1205 192
rect 1199 190 1200 191
rect 1123 188 1200 190
rect 1123 187 1124 188
rect 1118 186 1124 187
rect 1199 187 1200 188
rect 1204 187 1205 191
rect 1199 186 1205 187
rect 830 184 836 185
rect 134 167 140 168
rect 110 165 116 166
rect 110 161 111 165
rect 115 161 116 165
rect 134 163 135 167
rect 139 163 140 167
rect 134 162 140 163
rect 166 167 172 168
rect 166 163 167 167
rect 171 163 172 167
rect 166 162 172 163
rect 214 167 220 168
rect 214 163 215 167
rect 219 163 220 167
rect 214 162 220 163
rect 262 167 268 168
rect 262 163 263 167
rect 267 163 268 167
rect 262 162 268 163
rect 310 167 316 168
rect 310 163 311 167
rect 315 163 316 167
rect 310 162 316 163
rect 366 167 372 168
rect 366 163 367 167
rect 371 163 372 167
rect 366 162 372 163
rect 414 167 420 168
rect 414 163 415 167
rect 419 163 420 167
rect 414 162 420 163
rect 470 167 476 168
rect 470 163 471 167
rect 475 163 476 167
rect 470 162 476 163
rect 534 167 540 168
rect 534 163 535 167
rect 539 163 540 167
rect 534 162 540 163
rect 606 167 612 168
rect 606 163 607 167
rect 611 163 612 167
rect 606 162 612 163
rect 686 167 692 168
rect 686 163 687 167
rect 691 163 692 167
rect 686 162 692 163
rect 774 167 780 168
rect 774 163 775 167
rect 779 163 780 167
rect 774 162 780 163
rect 862 167 868 168
rect 862 163 863 167
rect 867 163 868 167
rect 862 162 868 163
rect 958 167 964 168
rect 958 163 959 167
rect 963 163 964 167
rect 958 162 964 163
rect 1054 167 1060 168
rect 1054 163 1055 167
rect 1059 163 1060 167
rect 1054 162 1060 163
rect 1150 167 1156 168
rect 1150 163 1151 167
rect 1155 163 1156 167
rect 1150 162 1156 163
rect 1238 167 1244 168
rect 1238 163 1239 167
rect 1243 163 1244 167
rect 1238 162 1244 163
rect 1326 167 1332 168
rect 1326 163 1327 167
rect 1331 163 1332 167
rect 1326 162 1332 163
rect 1414 167 1420 168
rect 1414 163 1415 167
rect 1419 163 1420 167
rect 1414 162 1420 163
rect 1502 167 1508 168
rect 1502 163 1503 167
rect 1507 163 1508 167
rect 1502 162 1508 163
rect 1590 167 1596 168
rect 1590 163 1591 167
rect 1595 163 1596 167
rect 1590 162 1596 163
rect 1654 167 1660 168
rect 1654 163 1655 167
rect 1659 163 1660 167
rect 1654 162 1660 163
rect 1694 165 1700 166
rect 110 160 116 161
rect 1694 161 1695 165
rect 1699 161 1700 165
rect 1694 160 1700 161
rect 150 159 157 160
rect 150 155 151 159
rect 156 155 157 159
rect 183 159 189 160
rect 183 158 184 159
rect 150 154 157 155
rect 176 156 184 158
rect 134 150 140 151
rect 110 148 116 149
rect 110 144 111 148
rect 115 144 116 148
rect 134 146 135 150
rect 139 146 140 150
rect 134 145 140 146
rect 166 150 172 151
rect 166 146 167 150
rect 171 146 172 150
rect 166 145 172 146
rect 110 143 116 144
rect 151 143 157 144
rect 151 139 152 143
rect 156 142 157 143
rect 176 142 178 156
rect 183 155 184 156
rect 188 155 189 159
rect 231 159 237 160
rect 231 158 232 159
rect 183 154 189 155
rect 208 156 232 158
rect 156 140 178 142
rect 183 143 189 144
rect 156 139 157 140
rect 151 138 157 139
rect 183 139 184 143
rect 188 142 189 143
rect 208 142 210 156
rect 231 155 232 156
rect 236 155 237 159
rect 279 159 285 160
rect 279 158 280 159
rect 231 154 237 155
rect 256 156 280 158
rect 214 150 220 151
rect 214 146 215 150
rect 219 146 220 150
rect 214 145 220 146
rect 188 140 210 142
rect 231 143 237 144
rect 188 139 189 140
rect 183 138 189 139
rect 231 139 232 143
rect 236 142 237 143
rect 256 142 258 156
rect 279 155 280 156
rect 284 155 285 159
rect 327 159 333 160
rect 327 158 328 159
rect 279 154 285 155
rect 319 156 328 158
rect 262 150 268 151
rect 262 146 263 150
rect 267 146 268 150
rect 262 145 268 146
rect 310 150 316 151
rect 310 146 311 150
rect 315 146 316 150
rect 310 145 316 146
rect 236 140 258 142
rect 279 143 285 144
rect 236 139 237 140
rect 231 138 237 139
rect 279 139 280 143
rect 284 142 285 143
rect 319 142 321 156
rect 327 155 328 156
rect 332 155 333 159
rect 383 159 389 160
rect 383 158 384 159
rect 327 154 333 155
rect 356 156 384 158
rect 284 140 321 142
rect 327 143 333 144
rect 284 139 285 140
rect 279 138 285 139
rect 327 139 328 143
rect 332 142 333 143
rect 356 142 358 156
rect 383 155 384 156
rect 388 155 389 159
rect 431 159 437 160
rect 431 158 432 159
rect 383 154 389 155
rect 409 156 432 158
rect 366 150 372 151
rect 366 146 367 150
rect 371 146 372 150
rect 366 145 372 146
rect 332 140 358 142
rect 383 143 389 144
rect 332 139 333 140
rect 327 138 333 139
rect 383 139 384 143
rect 388 142 389 143
rect 409 142 411 156
rect 431 155 432 156
rect 436 155 437 159
rect 487 159 493 160
rect 487 158 488 159
rect 431 154 437 155
rect 460 156 488 158
rect 414 150 420 151
rect 414 146 415 150
rect 419 146 420 150
rect 414 145 420 146
rect 388 140 411 142
rect 431 143 437 144
rect 388 139 389 140
rect 383 138 389 139
rect 431 139 432 143
rect 436 142 437 143
rect 460 142 462 156
rect 487 155 488 156
rect 492 155 493 159
rect 551 159 557 160
rect 551 158 552 159
rect 487 154 493 155
rect 524 156 552 158
rect 470 150 476 151
rect 470 146 471 150
rect 475 146 476 150
rect 470 145 476 146
rect 436 140 462 142
rect 487 143 493 144
rect 436 139 437 140
rect 431 138 437 139
rect 487 139 488 143
rect 492 142 493 143
rect 524 142 526 156
rect 551 155 552 156
rect 556 155 557 159
rect 551 154 557 155
rect 623 159 629 160
rect 623 155 624 159
rect 628 158 629 159
rect 646 159 652 160
rect 646 158 647 159
rect 628 156 647 158
rect 628 155 629 156
rect 623 154 629 155
rect 646 155 647 156
rect 651 155 652 159
rect 703 159 709 160
rect 703 158 704 159
rect 646 154 652 155
rect 668 156 704 158
rect 534 150 540 151
rect 534 146 535 150
rect 539 146 540 150
rect 534 145 540 146
rect 606 150 612 151
rect 606 146 607 150
rect 611 146 612 150
rect 606 145 612 146
rect 492 140 526 142
rect 551 143 557 144
rect 492 139 493 140
rect 487 138 493 139
rect 551 139 552 143
rect 556 142 557 143
rect 614 143 620 144
rect 614 142 615 143
rect 556 140 615 142
rect 556 139 557 140
rect 551 138 557 139
rect 614 139 615 140
rect 619 139 620 143
rect 614 138 620 139
rect 623 143 629 144
rect 623 139 624 143
rect 628 142 629 143
rect 668 142 670 156
rect 703 155 704 156
rect 708 155 709 159
rect 791 159 797 160
rect 791 158 792 159
rect 703 154 709 155
rect 716 156 792 158
rect 686 150 692 151
rect 686 146 687 150
rect 691 146 692 150
rect 686 145 692 146
rect 628 140 670 142
rect 703 143 709 144
rect 628 139 629 140
rect 623 138 629 139
rect 703 139 704 143
rect 708 142 709 143
rect 716 142 718 156
rect 791 155 792 156
rect 796 155 797 159
rect 879 159 885 160
rect 879 158 880 159
rect 791 154 797 155
rect 836 156 880 158
rect 774 150 780 151
rect 774 146 775 150
rect 779 146 780 150
rect 774 145 780 146
rect 708 140 718 142
rect 791 143 797 144
rect 708 139 709 140
rect 703 138 709 139
rect 791 139 792 143
rect 796 142 797 143
rect 836 142 838 156
rect 879 155 880 156
rect 884 155 885 159
rect 879 154 885 155
rect 975 159 981 160
rect 975 155 976 159
rect 980 158 981 159
rect 998 159 1004 160
rect 998 158 999 159
rect 980 156 999 158
rect 980 155 981 156
rect 975 154 981 155
rect 998 155 999 156
rect 1003 155 1004 159
rect 998 154 1004 155
rect 1071 159 1080 160
rect 1071 155 1072 159
rect 1079 155 1080 159
rect 1167 159 1173 160
rect 1167 158 1168 159
rect 1071 154 1080 155
rect 1084 156 1168 158
rect 862 150 868 151
rect 862 146 863 150
rect 867 146 868 150
rect 862 145 868 146
rect 958 150 964 151
rect 958 146 959 150
rect 963 146 964 150
rect 958 145 964 146
rect 1054 150 1060 151
rect 1084 150 1086 156
rect 1167 155 1168 156
rect 1172 155 1173 159
rect 1167 154 1173 155
rect 1255 159 1261 160
rect 1255 155 1256 159
rect 1260 158 1261 159
rect 1310 159 1316 160
rect 1260 156 1302 158
rect 1260 155 1261 156
rect 1255 154 1261 155
rect 1054 146 1055 150
rect 1059 146 1060 150
rect 1054 145 1060 146
rect 1064 148 1086 150
rect 1150 150 1156 151
rect 796 140 838 142
rect 879 143 885 144
rect 796 139 797 140
rect 791 138 797 139
rect 879 139 880 143
rect 884 142 885 143
rect 918 143 924 144
rect 918 142 919 143
rect 884 140 919 142
rect 884 139 885 140
rect 879 138 885 139
rect 918 139 919 140
rect 923 139 924 143
rect 918 138 924 139
rect 975 143 981 144
rect 975 139 976 143
rect 980 142 981 143
rect 1064 142 1066 148
rect 1150 146 1151 150
rect 1155 146 1156 150
rect 1150 145 1156 146
rect 1238 150 1244 151
rect 1238 146 1239 150
rect 1243 146 1244 150
rect 1238 145 1244 146
rect 980 140 1066 142
rect 1071 143 1077 144
rect 980 139 981 140
rect 975 138 981 139
rect 1071 139 1072 143
rect 1076 139 1077 143
rect 1071 138 1077 139
rect 1162 143 1173 144
rect 1162 139 1163 143
rect 1167 139 1168 143
rect 1172 139 1173 143
rect 1162 138 1173 139
rect 1194 143 1200 144
rect 1194 139 1195 143
rect 1199 142 1200 143
rect 1255 143 1261 144
rect 1255 142 1256 143
rect 1199 140 1256 142
rect 1199 139 1200 140
rect 1194 138 1200 139
rect 1255 139 1256 140
rect 1260 139 1261 143
rect 1300 142 1302 156
rect 1310 155 1311 159
rect 1315 158 1316 159
rect 1343 159 1349 160
rect 1343 158 1344 159
rect 1315 156 1344 158
rect 1315 155 1316 156
rect 1310 154 1316 155
rect 1343 155 1344 156
rect 1348 155 1349 159
rect 1343 154 1349 155
rect 1431 159 1437 160
rect 1431 155 1432 159
rect 1436 158 1437 159
rect 1519 159 1525 160
rect 1436 156 1499 158
rect 1436 155 1437 156
rect 1431 154 1437 155
rect 1326 150 1332 151
rect 1326 146 1327 150
rect 1331 146 1332 150
rect 1326 145 1332 146
rect 1414 150 1420 151
rect 1414 146 1415 150
rect 1419 146 1420 150
rect 1414 145 1420 146
rect 1343 143 1349 144
rect 1343 142 1344 143
rect 1300 140 1344 142
rect 1255 138 1261 139
rect 1343 139 1344 140
rect 1348 139 1349 143
rect 1343 138 1349 139
rect 1431 143 1437 144
rect 1431 139 1432 143
rect 1436 139 1437 143
rect 1497 142 1499 156
rect 1519 155 1520 159
rect 1524 158 1525 159
rect 1534 159 1540 160
rect 1534 158 1535 159
rect 1524 156 1535 158
rect 1524 155 1525 156
rect 1519 154 1525 155
rect 1534 155 1535 156
rect 1539 155 1540 159
rect 1534 154 1540 155
rect 1542 159 1548 160
rect 1542 155 1543 159
rect 1547 158 1548 159
rect 1607 159 1613 160
rect 1607 158 1608 159
rect 1547 156 1608 158
rect 1547 155 1548 156
rect 1542 154 1548 155
rect 1607 155 1608 156
rect 1612 155 1613 159
rect 1607 154 1613 155
rect 1670 159 1677 160
rect 1670 155 1671 159
rect 1676 155 1677 159
rect 1670 154 1677 155
rect 1502 150 1508 151
rect 1502 146 1503 150
rect 1507 146 1508 150
rect 1502 145 1508 146
rect 1590 150 1596 151
rect 1590 146 1591 150
rect 1595 146 1596 150
rect 1590 145 1596 146
rect 1654 150 1660 151
rect 1654 146 1655 150
rect 1659 146 1660 150
rect 1654 145 1660 146
rect 1694 148 1700 149
rect 1694 144 1695 148
rect 1699 144 1700 148
rect 1519 143 1525 144
rect 1519 142 1520 143
rect 1497 140 1520 142
rect 1431 138 1437 139
rect 1519 139 1520 140
rect 1524 139 1525 143
rect 1519 138 1525 139
rect 1578 143 1584 144
rect 1578 139 1579 143
rect 1583 142 1584 143
rect 1607 143 1613 144
rect 1607 142 1608 143
rect 1583 140 1608 142
rect 1583 139 1584 140
rect 1578 138 1584 139
rect 1607 139 1608 140
rect 1612 139 1613 143
rect 1607 138 1613 139
rect 1642 143 1648 144
rect 1642 139 1643 143
rect 1647 142 1648 143
rect 1671 143 1677 144
rect 1694 143 1700 144
rect 1671 142 1672 143
rect 1647 140 1672 142
rect 1647 139 1648 140
rect 1642 138 1648 139
rect 1671 139 1672 140
rect 1676 139 1677 143
rect 1671 138 1677 139
rect 1026 135 1032 136
rect 1026 131 1027 135
rect 1031 134 1032 135
rect 1072 134 1074 138
rect 1031 132 1074 134
rect 1433 134 1435 138
rect 1542 135 1548 136
rect 1542 134 1543 135
rect 1433 132 1543 134
rect 1031 131 1032 132
rect 1026 130 1032 131
rect 1542 131 1543 132
rect 1547 131 1548 135
rect 1542 130 1548 131
rect 1577 116 1634 118
rect 575 115 581 116
rect 160 112 187 114
rect 192 112 219 114
rect 224 112 251 114
rect 256 112 283 114
rect 288 112 315 114
rect 319 112 347 114
rect 352 112 379 114
rect 384 112 411 114
rect 416 112 443 114
rect 448 112 475 114
rect 480 112 507 114
rect 512 112 539 114
rect 544 112 571 114
rect 150 111 157 112
rect 110 108 116 109
rect 110 104 111 108
rect 115 104 116 108
rect 150 107 151 111
rect 156 107 157 111
rect 110 103 116 104
rect 134 106 140 107
rect 150 106 157 107
rect 134 102 135 106
rect 139 102 140 106
rect 134 101 140 102
rect 151 95 157 96
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 151 91 152 95
rect 156 94 157 95
rect 160 94 162 112
rect 183 111 189 112
rect 183 107 184 111
rect 188 107 189 111
rect 166 106 172 107
rect 183 106 189 107
rect 166 102 167 106
rect 171 102 172 106
rect 166 101 172 102
rect 156 92 162 94
rect 183 95 189 96
rect 156 91 157 92
rect 151 90 157 91
rect 183 91 184 95
rect 188 94 189 95
rect 192 94 194 112
rect 215 111 221 112
rect 215 107 216 111
rect 220 107 221 111
rect 198 106 204 107
rect 215 106 221 107
rect 198 102 199 106
rect 203 102 204 106
rect 198 101 204 102
rect 188 92 194 94
rect 215 95 221 96
rect 188 91 189 92
rect 183 90 189 91
rect 215 91 216 95
rect 220 94 221 95
rect 224 94 226 112
rect 247 111 253 112
rect 247 107 248 111
rect 252 107 253 111
rect 230 106 236 107
rect 247 106 253 107
rect 230 102 231 106
rect 235 102 236 106
rect 230 101 236 102
rect 220 92 226 94
rect 247 95 253 96
rect 220 91 221 92
rect 215 90 221 91
rect 247 91 248 95
rect 252 94 253 95
rect 256 94 258 112
rect 279 111 285 112
rect 279 107 280 111
rect 284 107 285 111
rect 262 106 268 107
rect 279 106 285 107
rect 262 102 263 106
rect 267 102 268 106
rect 262 101 268 102
rect 252 92 258 94
rect 279 95 285 96
rect 252 91 253 92
rect 247 90 253 91
rect 279 91 280 95
rect 284 94 285 95
rect 288 94 290 112
rect 311 111 317 112
rect 311 107 312 111
rect 316 107 317 111
rect 294 106 300 107
rect 311 106 317 107
rect 294 102 295 106
rect 299 102 300 106
rect 294 101 300 102
rect 284 92 290 94
rect 311 95 317 96
rect 284 91 285 92
rect 279 90 285 91
rect 311 91 312 95
rect 316 94 317 95
rect 319 94 321 112
rect 343 111 349 112
rect 343 107 344 111
rect 348 107 349 111
rect 326 106 332 107
rect 343 106 349 107
rect 326 102 327 106
rect 331 102 332 106
rect 326 101 332 102
rect 316 92 321 94
rect 343 95 349 96
rect 316 91 317 92
rect 311 90 317 91
rect 343 91 344 95
rect 348 94 349 95
rect 352 94 354 112
rect 375 111 381 112
rect 375 107 376 111
rect 380 107 381 111
rect 358 106 364 107
rect 375 106 381 107
rect 358 102 359 106
rect 363 102 364 106
rect 358 101 364 102
rect 348 92 354 94
rect 375 95 381 96
rect 348 91 349 92
rect 343 90 349 91
rect 375 91 376 95
rect 380 94 381 95
rect 384 94 386 112
rect 407 111 413 112
rect 407 107 408 111
rect 412 107 413 111
rect 390 106 396 107
rect 407 106 413 107
rect 390 102 391 106
rect 395 102 396 106
rect 390 101 396 102
rect 380 92 386 94
rect 407 95 413 96
rect 380 91 381 92
rect 375 90 381 91
rect 407 91 408 95
rect 412 94 413 95
rect 416 94 418 112
rect 439 111 445 112
rect 439 107 440 111
rect 444 107 445 111
rect 422 106 428 107
rect 439 106 445 107
rect 422 102 423 106
rect 427 102 428 106
rect 422 101 428 102
rect 412 92 418 94
rect 439 95 445 96
rect 412 91 413 92
rect 407 90 413 91
rect 439 91 440 95
rect 444 94 445 95
rect 448 94 450 112
rect 471 111 477 112
rect 471 107 472 111
rect 476 107 477 111
rect 454 106 460 107
rect 471 106 477 107
rect 454 102 455 106
rect 459 102 460 106
rect 454 101 460 102
rect 444 92 450 94
rect 471 95 477 96
rect 444 91 445 92
rect 439 90 445 91
rect 471 91 472 95
rect 476 94 477 95
rect 480 94 482 112
rect 503 111 509 112
rect 503 107 504 111
rect 508 107 509 111
rect 486 106 492 107
rect 503 106 509 107
rect 486 102 487 106
rect 491 102 492 106
rect 486 101 492 102
rect 476 92 482 94
rect 503 95 509 96
rect 476 91 477 92
rect 471 90 477 91
rect 503 91 504 95
rect 508 94 509 95
rect 512 94 514 112
rect 535 111 541 112
rect 535 107 536 111
rect 540 107 541 111
rect 518 106 524 107
rect 535 106 541 107
rect 518 102 519 106
rect 523 102 524 106
rect 518 101 524 102
rect 508 92 514 94
rect 535 95 541 96
rect 508 91 509 92
rect 503 90 509 91
rect 535 91 536 95
rect 540 94 541 95
rect 544 94 546 112
rect 567 111 573 112
rect 567 107 568 111
rect 572 107 573 111
rect 575 111 576 115
rect 580 114 581 115
rect 631 115 637 116
rect 580 112 618 114
rect 580 111 581 112
rect 575 110 581 111
rect 616 110 618 112
rect 623 111 629 112
rect 623 110 624 111
rect 616 108 624 110
rect 623 107 624 108
rect 628 107 629 111
rect 631 111 632 115
rect 636 114 637 115
rect 695 115 701 116
rect 636 112 691 114
rect 636 111 637 112
rect 631 110 637 111
rect 687 111 693 112
rect 687 107 688 111
rect 692 107 693 111
rect 695 111 696 115
rect 700 114 701 115
rect 767 115 773 116
rect 700 112 754 114
rect 700 111 701 112
rect 695 110 701 111
rect 752 110 754 112
rect 759 111 765 112
rect 759 110 760 111
rect 752 108 760 110
rect 759 107 760 108
rect 764 107 765 111
rect 767 111 768 115
rect 772 114 773 115
rect 847 115 853 116
rect 772 112 834 114
rect 772 111 773 112
rect 767 110 773 111
rect 832 110 834 112
rect 839 111 845 112
rect 839 110 840 111
rect 832 108 840 110
rect 839 107 840 108
rect 844 107 845 111
rect 847 111 848 115
rect 852 114 853 115
rect 1079 115 1085 116
rect 852 112 914 114
rect 852 111 853 112
rect 847 110 853 111
rect 912 110 914 112
rect 919 111 925 112
rect 919 110 920 111
rect 912 108 920 110
rect 919 107 920 108
rect 924 107 925 111
rect 998 111 1005 112
rect 998 107 999 111
rect 1004 107 1005 111
rect 1070 111 1077 112
rect 1070 107 1071 111
rect 1076 107 1077 111
rect 1079 111 1080 115
rect 1084 114 1085 115
rect 1143 115 1149 116
rect 1084 112 1130 114
rect 1084 111 1085 112
rect 1079 110 1085 111
rect 1128 110 1130 112
rect 1135 111 1141 112
rect 1135 110 1136 111
rect 1128 108 1136 110
rect 1135 107 1136 108
rect 1140 107 1141 111
rect 1143 111 1144 115
rect 1148 114 1149 115
rect 1148 112 1187 114
rect 1264 112 1282 114
rect 1304 112 1322 114
rect 1337 112 1354 114
rect 1369 112 1386 114
rect 1401 112 1418 114
rect 1433 112 1450 114
rect 1472 112 1490 114
rect 1497 112 1530 114
rect 1577 112 1579 116
rect 1584 112 1611 114
rect 1148 111 1149 112
rect 1143 110 1149 111
rect 1185 110 1187 112
rect 1191 111 1197 112
rect 1191 110 1192 111
rect 1185 108 1192 110
rect 1191 107 1192 108
rect 1196 107 1197 111
rect 1239 111 1245 112
rect 1239 107 1240 111
rect 1244 110 1245 111
rect 1264 110 1266 112
rect 1244 108 1266 110
rect 1244 107 1245 108
rect 550 106 556 107
rect 567 106 573 107
rect 606 106 612 107
rect 623 106 629 107
rect 670 106 676 107
rect 687 106 693 107
rect 742 106 748 107
rect 759 106 765 107
rect 822 106 828 107
rect 839 106 845 107
rect 902 106 908 107
rect 919 106 925 107
rect 982 106 988 107
rect 998 106 1005 107
rect 1054 106 1060 107
rect 1070 106 1077 107
rect 1118 106 1124 107
rect 1135 106 1141 107
rect 1174 106 1180 107
rect 1191 106 1197 107
rect 1222 106 1228 107
rect 1239 106 1245 107
rect 1270 106 1276 107
rect 550 102 551 106
rect 555 102 556 106
rect 550 101 556 102
rect 606 102 607 106
rect 611 102 612 106
rect 606 101 612 102
rect 670 102 671 106
rect 675 102 676 106
rect 670 101 676 102
rect 742 102 743 106
rect 747 102 748 106
rect 742 101 748 102
rect 822 102 823 106
rect 827 102 828 106
rect 822 101 828 102
rect 902 102 903 106
rect 907 102 908 106
rect 902 101 908 102
rect 982 102 983 106
rect 987 102 988 106
rect 982 101 988 102
rect 1054 102 1055 106
rect 1059 102 1060 106
rect 1054 101 1060 102
rect 1118 102 1119 106
rect 1123 102 1124 106
rect 1118 101 1124 102
rect 1174 102 1175 106
rect 1179 102 1180 106
rect 1174 101 1180 102
rect 1222 102 1223 106
rect 1227 102 1228 106
rect 1222 101 1228 102
rect 1270 102 1271 106
rect 1275 102 1276 106
rect 1270 101 1276 102
rect 540 92 546 94
rect 567 95 573 96
rect 540 91 541 92
rect 535 90 541 91
rect 567 91 568 95
rect 572 94 573 95
rect 575 95 581 96
rect 575 94 576 95
rect 572 92 576 94
rect 572 91 573 92
rect 567 90 573 91
rect 575 91 576 92
rect 580 91 581 95
rect 575 90 581 91
rect 623 95 629 96
rect 623 91 624 95
rect 628 94 629 95
rect 631 95 637 96
rect 631 94 632 95
rect 628 92 632 94
rect 628 91 629 92
rect 623 90 629 91
rect 631 91 632 92
rect 636 91 637 95
rect 631 90 637 91
rect 687 95 693 96
rect 687 91 688 95
rect 692 94 693 95
rect 695 95 701 96
rect 695 94 696 95
rect 692 92 696 94
rect 692 91 693 92
rect 687 90 693 91
rect 695 91 696 92
rect 700 91 701 95
rect 695 90 701 91
rect 759 95 765 96
rect 759 91 760 95
rect 764 94 765 95
rect 767 95 773 96
rect 767 94 768 95
rect 764 92 768 94
rect 764 91 765 92
rect 759 90 765 91
rect 767 91 768 92
rect 772 91 773 95
rect 767 90 773 91
rect 839 95 845 96
rect 839 91 840 95
rect 844 94 845 95
rect 847 95 853 96
rect 847 94 848 95
rect 844 92 848 94
rect 844 91 845 92
rect 839 90 845 91
rect 847 91 848 92
rect 852 91 853 95
rect 847 90 853 91
rect 918 95 925 96
rect 918 91 919 95
rect 924 91 925 95
rect 918 90 925 91
rect 999 95 1005 96
rect 999 91 1000 95
rect 1004 94 1005 95
rect 1026 95 1032 96
rect 1026 94 1027 95
rect 1004 92 1027 94
rect 1004 91 1005 92
rect 999 90 1005 91
rect 1026 91 1027 92
rect 1031 91 1032 95
rect 1026 90 1032 91
rect 1071 95 1077 96
rect 1071 91 1072 95
rect 1076 94 1077 95
rect 1079 95 1085 96
rect 1079 94 1080 95
rect 1076 92 1080 94
rect 1076 91 1077 92
rect 1071 90 1077 91
rect 1079 91 1080 92
rect 1084 91 1085 95
rect 1079 90 1085 91
rect 1135 95 1141 96
rect 1135 91 1136 95
rect 1140 94 1141 95
rect 1143 95 1149 96
rect 1143 94 1144 95
rect 1140 92 1144 94
rect 1140 91 1141 92
rect 1135 90 1141 91
rect 1143 91 1144 92
rect 1148 91 1149 95
rect 1143 90 1149 91
rect 1191 95 1200 96
rect 1191 91 1192 95
rect 1199 91 1200 95
rect 1239 95 1245 96
rect 1239 94 1240 95
rect 1191 90 1200 91
rect 1232 92 1240 94
rect 110 86 116 87
rect 134 89 140 90
rect 134 85 135 89
rect 139 85 140 89
rect 134 84 140 85
rect 166 89 172 90
rect 166 85 167 89
rect 171 85 172 89
rect 166 84 172 85
rect 198 89 204 90
rect 198 85 199 89
rect 203 85 204 89
rect 198 84 204 85
rect 230 89 236 90
rect 230 85 231 89
rect 235 85 236 89
rect 230 84 236 85
rect 262 89 268 90
rect 262 85 263 89
rect 267 85 268 89
rect 262 84 268 85
rect 294 89 300 90
rect 294 85 295 89
rect 299 85 300 89
rect 294 84 300 85
rect 326 89 332 90
rect 326 85 327 89
rect 331 85 332 89
rect 326 84 332 85
rect 358 89 364 90
rect 358 85 359 89
rect 363 85 364 89
rect 358 84 364 85
rect 390 89 396 90
rect 390 85 391 89
rect 395 85 396 89
rect 390 84 396 85
rect 422 89 428 90
rect 422 85 423 89
rect 427 85 428 89
rect 422 84 428 85
rect 454 89 460 90
rect 454 85 455 89
rect 459 85 460 89
rect 454 84 460 85
rect 486 89 492 90
rect 486 85 487 89
rect 491 85 492 89
rect 486 84 492 85
rect 518 89 524 90
rect 518 85 519 89
rect 523 85 524 89
rect 518 84 524 85
rect 550 89 556 90
rect 550 85 551 89
rect 555 85 556 89
rect 550 84 556 85
rect 606 89 612 90
rect 606 85 607 89
rect 611 85 612 89
rect 670 89 676 90
rect 606 84 612 85
rect 622 87 628 88
rect 622 83 623 87
rect 627 86 628 87
rect 637 87 643 88
rect 637 86 638 87
rect 627 84 638 86
rect 627 83 628 84
rect 622 82 628 83
rect 637 83 638 84
rect 642 83 643 87
rect 670 85 671 89
rect 675 85 676 89
rect 670 84 676 85
rect 742 89 748 90
rect 742 85 743 89
rect 747 85 748 89
rect 742 84 748 85
rect 822 89 828 90
rect 822 85 823 89
rect 827 85 828 89
rect 822 84 828 85
rect 902 89 908 90
rect 902 85 903 89
rect 907 85 908 89
rect 902 84 908 85
rect 982 89 988 90
rect 982 85 983 89
rect 987 85 988 89
rect 982 84 988 85
rect 1054 89 1060 90
rect 1054 85 1055 89
rect 1059 85 1060 89
rect 1054 84 1060 85
rect 1118 89 1124 90
rect 1118 85 1119 89
rect 1123 85 1124 89
rect 1118 84 1124 85
rect 1174 89 1180 90
rect 1174 85 1175 89
rect 1179 85 1180 89
rect 1174 84 1180 85
rect 1222 89 1228 90
rect 1222 85 1223 89
rect 1227 85 1228 89
rect 1222 84 1228 85
rect 637 82 643 83
rect 1070 83 1076 84
rect 1070 79 1071 83
rect 1075 82 1076 83
rect 1232 82 1234 92
rect 1239 91 1240 92
rect 1244 91 1245 95
rect 1280 94 1282 112
rect 1287 111 1293 112
rect 1287 107 1288 111
rect 1292 110 1293 111
rect 1304 110 1306 112
rect 1292 108 1306 110
rect 1292 107 1293 108
rect 1287 106 1293 107
rect 1310 106 1316 107
rect 1310 102 1311 106
rect 1315 102 1316 106
rect 1310 101 1316 102
rect 1287 95 1293 96
rect 1287 94 1288 95
rect 1280 92 1288 94
rect 1239 90 1245 91
rect 1287 91 1288 92
rect 1292 91 1293 95
rect 1320 94 1322 112
rect 1327 111 1333 112
rect 1327 107 1328 111
rect 1332 110 1333 111
rect 1337 110 1339 112
rect 1332 108 1339 110
rect 1332 107 1333 108
rect 1327 106 1333 107
rect 1342 106 1348 107
rect 1342 102 1343 106
rect 1347 102 1348 106
rect 1342 101 1348 102
rect 1327 95 1333 96
rect 1327 94 1328 95
rect 1320 92 1328 94
rect 1287 90 1293 91
rect 1327 91 1328 92
rect 1332 91 1333 95
rect 1352 94 1354 112
rect 1359 111 1365 112
rect 1359 107 1360 111
rect 1364 110 1365 111
rect 1369 110 1371 112
rect 1364 108 1371 110
rect 1364 107 1365 108
rect 1359 106 1365 107
rect 1374 106 1380 107
rect 1374 102 1375 106
rect 1379 102 1380 106
rect 1374 101 1380 102
rect 1359 95 1365 96
rect 1359 94 1360 95
rect 1352 92 1360 94
rect 1327 90 1333 91
rect 1359 91 1360 92
rect 1364 91 1365 95
rect 1384 94 1386 112
rect 1391 111 1397 112
rect 1391 107 1392 111
rect 1396 110 1397 111
rect 1401 110 1403 112
rect 1396 108 1403 110
rect 1396 107 1397 108
rect 1391 106 1397 107
rect 1406 106 1412 107
rect 1406 102 1407 106
rect 1411 102 1412 106
rect 1406 101 1412 102
rect 1391 95 1397 96
rect 1391 94 1392 95
rect 1384 92 1392 94
rect 1359 90 1365 91
rect 1391 91 1392 92
rect 1396 91 1397 95
rect 1416 94 1418 112
rect 1423 111 1429 112
rect 1423 107 1424 111
rect 1428 110 1429 111
rect 1433 110 1435 112
rect 1428 108 1435 110
rect 1428 107 1429 108
rect 1423 106 1429 107
rect 1438 106 1444 107
rect 1438 102 1439 106
rect 1443 102 1444 106
rect 1438 101 1444 102
rect 1423 95 1429 96
rect 1423 94 1424 95
rect 1416 92 1424 94
rect 1391 90 1397 91
rect 1423 91 1424 92
rect 1428 91 1429 95
rect 1448 94 1450 112
rect 1455 111 1461 112
rect 1455 107 1456 111
rect 1460 110 1461 111
rect 1472 110 1474 112
rect 1460 108 1474 110
rect 1460 107 1461 108
rect 1455 106 1461 107
rect 1478 106 1484 107
rect 1478 102 1479 106
rect 1483 102 1484 106
rect 1478 101 1484 102
rect 1488 98 1490 112
rect 1495 111 1501 112
rect 1495 107 1496 111
rect 1500 107 1501 111
rect 1495 106 1501 107
rect 1518 106 1524 107
rect 1518 102 1519 106
rect 1523 102 1524 106
rect 1518 101 1524 102
rect 1488 96 1499 98
rect 1455 95 1461 96
rect 1455 94 1456 95
rect 1448 92 1456 94
rect 1423 90 1429 91
rect 1455 91 1456 92
rect 1460 91 1461 95
rect 1455 90 1461 91
rect 1495 95 1501 96
rect 1495 91 1496 95
rect 1500 91 1501 95
rect 1528 94 1530 112
rect 1534 111 1541 112
rect 1534 107 1535 111
rect 1540 107 1541 111
rect 1575 111 1581 112
rect 1575 107 1576 111
rect 1580 107 1581 111
rect 1534 106 1541 107
rect 1558 106 1564 107
rect 1575 106 1581 107
rect 1558 102 1559 106
rect 1563 102 1564 106
rect 1558 101 1564 102
rect 1535 95 1541 96
rect 1535 94 1536 95
rect 1528 92 1536 94
rect 1495 90 1501 91
rect 1535 91 1536 92
rect 1540 91 1541 95
rect 1535 90 1541 91
rect 1575 95 1581 96
rect 1575 91 1576 95
rect 1580 94 1581 95
rect 1584 94 1586 112
rect 1607 111 1613 112
rect 1607 107 1608 111
rect 1612 107 1613 111
rect 1590 106 1596 107
rect 1607 106 1613 107
rect 1622 106 1628 107
rect 1590 102 1591 106
rect 1595 102 1596 106
rect 1590 101 1596 102
rect 1622 102 1623 106
rect 1627 102 1628 106
rect 1622 101 1628 102
rect 1580 92 1586 94
rect 1602 95 1613 96
rect 1580 91 1581 92
rect 1575 90 1581 91
rect 1602 91 1603 95
rect 1607 91 1608 95
rect 1612 91 1613 95
rect 1632 94 1634 116
rect 1641 112 1666 114
rect 1639 111 1645 112
rect 1639 107 1640 111
rect 1644 107 1645 111
rect 1639 106 1645 107
rect 1654 106 1660 107
rect 1654 102 1655 106
rect 1659 102 1660 106
rect 1654 101 1660 102
rect 1639 95 1645 96
rect 1639 94 1640 95
rect 1632 92 1640 94
rect 1602 90 1613 91
rect 1639 91 1640 92
rect 1644 91 1645 95
rect 1664 94 1666 112
rect 1670 111 1677 112
rect 1670 107 1671 111
rect 1676 107 1677 111
rect 1670 106 1677 107
rect 1694 108 1700 109
rect 1694 104 1695 108
rect 1699 104 1700 108
rect 1694 103 1700 104
rect 1671 95 1677 96
rect 1671 94 1672 95
rect 1664 92 1672 94
rect 1639 90 1645 91
rect 1671 91 1672 92
rect 1676 91 1677 95
rect 1671 90 1677 91
rect 1694 91 1700 92
rect 1270 89 1276 90
rect 1270 85 1271 89
rect 1275 85 1276 89
rect 1270 84 1276 85
rect 1310 89 1316 90
rect 1310 85 1311 89
rect 1315 85 1316 89
rect 1310 84 1316 85
rect 1342 89 1348 90
rect 1342 85 1343 89
rect 1347 85 1348 89
rect 1342 84 1348 85
rect 1374 89 1380 90
rect 1374 85 1375 89
rect 1379 85 1380 89
rect 1374 84 1380 85
rect 1406 89 1412 90
rect 1406 85 1407 89
rect 1411 85 1412 89
rect 1406 84 1412 85
rect 1438 89 1444 90
rect 1438 85 1439 89
rect 1443 85 1444 89
rect 1438 84 1444 85
rect 1478 89 1484 90
rect 1478 85 1479 89
rect 1483 85 1484 89
rect 1478 84 1484 85
rect 1518 89 1524 90
rect 1518 85 1519 89
rect 1523 85 1524 89
rect 1518 84 1524 85
rect 1558 89 1564 90
rect 1558 85 1559 89
rect 1563 85 1564 89
rect 1558 84 1564 85
rect 1590 89 1596 90
rect 1590 85 1591 89
rect 1595 85 1596 89
rect 1590 84 1596 85
rect 1622 89 1628 90
rect 1622 85 1623 89
rect 1627 85 1628 89
rect 1622 84 1628 85
rect 1654 89 1660 90
rect 1654 85 1655 89
rect 1659 85 1660 89
rect 1694 87 1695 91
rect 1699 87 1700 91
rect 1694 86 1700 87
rect 1654 84 1660 85
rect 1075 80 1234 82
rect 1075 79 1076 80
rect 1070 78 1076 79
<< m3c >>
rect 871 1759 875 1763
rect 111 1749 115 1753
rect 151 1751 155 1755
rect 183 1751 187 1755
rect 215 1751 219 1755
rect 247 1751 251 1755
rect 279 1751 283 1755
rect 311 1751 315 1755
rect 343 1751 347 1755
rect 375 1751 379 1755
rect 407 1751 411 1755
rect 439 1751 443 1755
rect 471 1751 475 1755
rect 503 1751 507 1755
rect 535 1751 539 1755
rect 567 1751 571 1755
rect 599 1751 603 1755
rect 631 1751 635 1755
rect 663 1751 667 1755
rect 695 1751 699 1755
rect 727 1751 731 1755
rect 759 1751 763 1755
rect 791 1751 795 1755
rect 823 1751 827 1755
rect 855 1751 859 1755
rect 887 1751 891 1755
rect 919 1751 923 1755
rect 951 1751 955 1755
rect 983 1751 987 1755
rect 1191 1755 1194 1759
rect 1194 1755 1195 1759
rect 1695 1749 1699 1753
rect 111 1732 115 1736
rect 151 1734 155 1738
rect 183 1734 187 1738
rect 215 1734 219 1738
rect 247 1734 251 1738
rect 279 1734 283 1738
rect 311 1734 315 1738
rect 343 1734 347 1738
rect 375 1734 379 1738
rect 407 1734 411 1738
rect 439 1734 443 1738
rect 471 1734 475 1738
rect 503 1734 507 1738
rect 535 1734 539 1738
rect 567 1734 571 1738
rect 599 1734 603 1738
rect 631 1734 635 1738
rect 663 1734 667 1738
rect 695 1734 699 1738
rect 727 1734 731 1738
rect 759 1734 763 1738
rect 791 1734 795 1738
rect 823 1734 827 1738
rect 855 1734 859 1738
rect 887 1734 891 1738
rect 919 1734 923 1738
rect 951 1734 955 1738
rect 983 1734 987 1738
rect 1695 1732 1699 1736
rect 1063 1727 1067 1731
rect 111 1700 115 1704
rect 207 1703 208 1707
rect 208 1703 211 1707
rect 895 1703 899 1707
rect 903 1707 907 1711
rect 1199 1703 1203 1707
rect 1207 1707 1211 1711
rect 191 1698 195 1702
rect 247 1698 251 1702
rect 319 1698 323 1702
rect 415 1698 419 1702
rect 527 1698 531 1702
rect 655 1698 659 1702
rect 791 1698 795 1702
rect 919 1698 923 1702
rect 1047 1698 1051 1702
rect 1159 1698 1163 1702
rect 1255 1698 1259 1702
rect 1335 1698 1339 1702
rect 1407 1698 1411 1702
rect 1463 1698 1467 1702
rect 1519 1698 1523 1702
rect 1567 1698 1571 1702
rect 1623 1698 1627 1702
rect 1655 1698 1659 1702
rect 1695 1700 1699 1704
rect 111 1683 115 1687
rect 407 1687 411 1691
rect 903 1687 907 1691
rect 1063 1687 1064 1691
rect 1064 1687 1067 1691
rect 1207 1687 1211 1691
rect 191 1681 195 1685
rect 247 1681 251 1685
rect 319 1681 323 1685
rect 415 1681 419 1685
rect 527 1681 531 1685
rect 655 1681 659 1685
rect 207 1675 211 1679
rect 791 1681 795 1685
rect 919 1681 923 1685
rect 1047 1681 1051 1685
rect 1159 1681 1163 1685
rect 1255 1681 1259 1685
rect 1335 1681 1339 1685
rect 1407 1681 1411 1685
rect 1463 1681 1467 1685
rect 1519 1681 1523 1685
rect 1567 1681 1571 1685
rect 1623 1681 1627 1685
rect 1655 1681 1659 1685
rect 1471 1675 1475 1679
rect 1695 1683 1699 1687
rect 155 1667 159 1671
rect 111 1657 115 1661
rect 135 1659 139 1663
rect 175 1659 179 1663
rect 263 1659 267 1663
rect 391 1659 395 1663
rect 543 1659 547 1663
rect 711 1659 715 1663
rect 879 1659 883 1663
rect 1039 1659 1043 1663
rect 1183 1659 1187 1663
rect 1319 1659 1323 1663
rect 1439 1659 1443 1663
rect 1559 1659 1563 1663
rect 1655 1659 1659 1663
rect 1695 1657 1699 1661
rect 111 1640 115 1644
rect 135 1642 139 1646
rect 175 1642 179 1646
rect 155 1635 156 1639
rect 156 1635 159 1639
rect 343 1651 347 1655
rect 263 1642 267 1646
rect 391 1642 395 1646
rect 407 1635 408 1639
rect 408 1635 411 1639
rect 543 1642 547 1646
rect 895 1651 896 1655
rect 896 1651 899 1655
rect 711 1642 715 1646
rect 879 1642 883 1646
rect 1199 1651 1200 1655
rect 1200 1651 1203 1655
rect 1039 1642 1043 1646
rect 1183 1642 1187 1646
rect 1019 1635 1023 1639
rect 1319 1642 1323 1646
rect 1439 1642 1443 1646
rect 1375 1635 1379 1639
rect 1471 1635 1475 1639
rect 1559 1642 1563 1646
rect 1671 1651 1672 1655
rect 1672 1651 1675 1655
rect 1655 1642 1659 1646
rect 1695 1640 1699 1644
rect 187 1627 191 1631
rect 111 1604 115 1608
rect 135 1602 139 1606
rect 167 1602 171 1606
rect 111 1587 115 1591
rect 151 1591 152 1595
rect 152 1591 155 1595
rect 199 1602 203 1606
rect 583 1619 587 1623
rect 343 1607 344 1611
rect 344 1607 347 1611
rect 247 1602 251 1606
rect 327 1602 331 1606
rect 439 1602 443 1606
rect 567 1602 571 1606
rect 711 1602 715 1606
rect 855 1602 859 1606
rect 583 1591 584 1595
rect 584 1591 587 1595
rect 723 1591 727 1595
rect 975 1607 979 1611
rect 1079 1607 1083 1611
rect 1175 1607 1179 1611
rect 1211 1611 1215 1615
rect 999 1602 1003 1606
rect 1127 1602 1131 1606
rect 1247 1602 1251 1606
rect 1359 1602 1363 1606
rect 1463 1602 1467 1606
rect 1019 1591 1020 1595
rect 1020 1591 1023 1595
rect 1211 1591 1215 1595
rect 1343 1591 1347 1595
rect 1375 1591 1376 1595
rect 1376 1591 1379 1595
rect 1479 1607 1480 1611
rect 1480 1607 1483 1611
rect 1567 1602 1571 1606
rect 1655 1602 1659 1606
rect 1623 1591 1627 1595
rect 1671 1607 1672 1611
rect 1672 1607 1675 1611
rect 1695 1604 1699 1608
rect 135 1585 139 1589
rect 167 1585 171 1589
rect 199 1585 203 1589
rect 247 1585 251 1589
rect 327 1585 331 1589
rect 439 1585 443 1589
rect 567 1585 571 1589
rect 711 1585 715 1589
rect 855 1585 859 1589
rect 999 1585 1003 1589
rect 1127 1585 1131 1589
rect 1247 1585 1251 1589
rect 1359 1585 1363 1589
rect 1463 1585 1467 1589
rect 1567 1585 1571 1589
rect 1655 1585 1659 1589
rect 1695 1587 1699 1591
rect 111 1569 115 1573
rect 135 1571 139 1575
rect 167 1571 171 1575
rect 231 1571 235 1575
rect 287 1571 291 1575
rect 343 1571 347 1575
rect 399 1571 403 1575
rect 455 1571 459 1575
rect 511 1571 515 1575
rect 575 1571 579 1575
rect 655 1571 659 1575
rect 751 1571 755 1575
rect 855 1571 859 1575
rect 959 1571 963 1575
rect 1063 1571 1067 1575
rect 1159 1571 1163 1575
rect 1247 1571 1251 1575
rect 1327 1571 1331 1575
rect 1399 1571 1403 1575
rect 1471 1571 1475 1575
rect 1535 1571 1539 1575
rect 1607 1571 1611 1575
rect 1655 1571 1659 1575
rect 1695 1569 1699 1573
rect 1703 1571 1707 1575
rect 111 1552 115 1556
rect 135 1554 139 1558
rect 167 1554 171 1558
rect 151 1547 152 1551
rect 152 1547 155 1551
rect 231 1554 235 1558
rect 299 1563 303 1567
rect 379 1563 383 1567
rect 287 1554 291 1558
rect 343 1554 347 1558
rect 399 1554 403 1558
rect 455 1554 459 1558
rect 511 1554 515 1558
rect 731 1563 735 1567
rect 575 1554 579 1558
rect 655 1554 659 1558
rect 723 1555 727 1559
rect 751 1554 755 1558
rect 855 1554 859 1558
rect 759 1547 763 1551
rect 975 1563 976 1567
rect 976 1563 979 1567
rect 1079 1563 1080 1567
rect 1080 1563 1083 1567
rect 1175 1563 1176 1567
rect 1176 1563 1179 1567
rect 959 1554 963 1558
rect 1063 1554 1067 1558
rect 1159 1554 1163 1558
rect 1247 1554 1251 1558
rect 1327 1554 1331 1558
rect 1375 1563 1379 1567
rect 1103 1547 1107 1551
rect 299 1539 303 1543
rect 379 1539 383 1543
rect 111 1524 115 1528
rect 211 1531 215 1535
rect 555 1539 559 1543
rect 1031 1539 1035 1543
rect 1195 1547 1199 1551
rect 1343 1547 1344 1551
rect 1344 1547 1347 1551
rect 1399 1554 1403 1558
rect 1471 1554 1475 1558
rect 1547 1563 1551 1567
rect 1535 1554 1539 1558
rect 1607 1554 1611 1558
rect 1623 1547 1624 1551
rect 1624 1547 1627 1551
rect 1671 1563 1672 1567
rect 1672 1563 1675 1567
rect 1655 1554 1659 1558
rect 1695 1552 1699 1556
rect 135 1522 139 1526
rect 175 1522 179 1526
rect 223 1522 227 1526
rect 279 1522 283 1526
rect 335 1522 339 1526
rect 399 1522 403 1526
rect 103 1503 107 1507
rect 111 1507 115 1511
rect 211 1511 215 1515
rect 319 1511 323 1515
rect 351 1511 352 1515
rect 352 1511 355 1515
rect 471 1527 475 1531
rect 639 1527 643 1531
rect 647 1531 651 1535
rect 731 1531 735 1535
rect 1095 1527 1096 1531
rect 1096 1527 1099 1531
rect 1187 1527 1191 1531
rect 1215 1527 1219 1531
rect 1255 1531 1259 1535
rect 1375 1527 1376 1531
rect 1376 1527 1379 1531
rect 1447 1527 1451 1531
rect 1547 1527 1551 1531
rect 463 1522 467 1526
rect 535 1522 539 1526
rect 607 1522 611 1526
rect 687 1522 691 1526
rect 775 1522 779 1526
rect 871 1522 875 1526
rect 975 1522 979 1526
rect 1079 1522 1083 1526
rect 1103 1519 1107 1523
rect 1175 1522 1179 1526
rect 1271 1522 1275 1526
rect 1359 1522 1363 1526
rect 1439 1522 1443 1526
rect 1519 1522 1523 1526
rect 1599 1522 1603 1526
rect 1671 1527 1672 1531
rect 1672 1527 1675 1531
rect 1655 1522 1659 1526
rect 1695 1524 1699 1528
rect 555 1511 556 1515
rect 556 1511 559 1515
rect 647 1511 651 1515
rect 719 1511 723 1515
rect 991 1511 992 1515
rect 992 1511 995 1515
rect 1195 1511 1196 1515
rect 1196 1511 1199 1515
rect 1335 1511 1339 1515
rect 1375 1511 1376 1515
rect 1376 1511 1379 1515
rect 1479 1511 1483 1515
rect 135 1505 139 1509
rect 175 1505 179 1509
rect 223 1505 227 1509
rect 279 1505 283 1509
rect 335 1505 339 1509
rect 399 1505 403 1509
rect 463 1505 467 1509
rect 535 1505 539 1509
rect 607 1505 611 1509
rect 687 1505 691 1509
rect 775 1505 779 1509
rect 871 1505 875 1509
rect 975 1505 979 1509
rect 1079 1505 1083 1509
rect 1175 1505 1179 1509
rect 1271 1505 1275 1509
rect 1359 1505 1363 1509
rect 1439 1505 1443 1509
rect 1519 1505 1523 1509
rect 1499 1499 1503 1503
rect 1639 1511 1643 1515
rect 1599 1505 1603 1509
rect 1655 1505 1659 1509
rect 1695 1507 1699 1511
rect 919 1487 923 1491
rect 1147 1487 1151 1491
rect 111 1469 115 1473
rect 175 1471 179 1475
rect 207 1471 211 1475
rect 239 1471 243 1475
rect 271 1471 275 1475
rect 303 1471 307 1475
rect 383 1479 387 1483
rect 335 1471 339 1475
rect 367 1471 371 1475
rect 399 1471 403 1475
rect 151 1463 155 1467
rect 111 1452 115 1456
rect 175 1454 179 1458
rect 207 1454 211 1458
rect 239 1454 243 1458
rect 271 1454 275 1458
rect 471 1479 475 1483
rect 431 1471 435 1475
rect 463 1471 467 1475
rect 495 1471 499 1475
rect 527 1471 531 1475
rect 559 1471 563 1475
rect 591 1471 595 1475
rect 623 1471 627 1475
rect 663 1471 667 1475
rect 703 1471 707 1475
rect 743 1471 747 1475
rect 775 1471 779 1475
rect 807 1472 811 1476
rect 895 1472 899 1476
rect 935 1472 939 1476
rect 1023 1472 1027 1476
rect 1079 1471 1083 1475
rect 1111 1472 1115 1476
rect 1167 1471 1171 1475
rect 1199 1471 1203 1475
rect 1239 1471 1243 1475
rect 1279 1471 1283 1475
rect 1319 1471 1323 1475
rect 1359 1471 1363 1475
rect 1399 1471 1403 1475
rect 1439 1471 1443 1475
rect 1479 1471 1483 1475
rect 1519 1471 1523 1475
rect 1559 1471 1563 1475
rect 1591 1471 1595 1475
rect 1623 1471 1627 1475
rect 1655 1471 1659 1475
rect 1695 1469 1699 1473
rect 303 1454 307 1458
rect 335 1454 339 1458
rect 367 1454 371 1458
rect 399 1454 403 1458
rect 431 1454 435 1458
rect 319 1447 320 1451
rect 320 1447 323 1451
rect 351 1447 352 1451
rect 352 1447 355 1451
rect 383 1447 384 1451
rect 384 1447 387 1451
rect 447 1463 448 1467
rect 448 1463 451 1467
rect 463 1454 467 1458
rect 495 1454 499 1458
rect 543 1463 544 1467
rect 544 1463 547 1467
rect 527 1454 531 1458
rect 559 1454 563 1458
rect 535 1447 539 1451
rect 591 1454 595 1458
rect 639 1463 640 1467
rect 640 1463 643 1467
rect 683 1463 684 1467
rect 684 1463 687 1467
rect 623 1454 627 1458
rect 663 1454 667 1458
rect 703 1454 707 1458
rect 743 1454 747 1458
rect 775 1453 779 1457
rect 719 1447 720 1451
rect 720 1447 723 1451
rect 887 1463 891 1467
rect 1095 1463 1096 1467
rect 1096 1463 1099 1467
rect 807 1453 811 1457
rect 919 1455 920 1459
rect 920 1455 923 1459
rect 935 1453 939 1457
rect 1039 1451 1043 1455
rect 895 1444 899 1448
rect 1079 1454 1083 1458
rect 1127 1451 1131 1455
rect 1147 1451 1148 1455
rect 1148 1451 1151 1455
rect 1167 1454 1171 1458
rect 1199 1454 1203 1458
rect 1231 1463 1235 1467
rect 1255 1463 1256 1467
rect 1256 1463 1259 1467
rect 815 1439 819 1443
rect 887 1439 891 1443
rect 535 1423 539 1427
rect 671 1423 675 1427
rect 911 1431 915 1435
rect 1139 1443 1143 1447
rect 1183 1447 1184 1451
rect 1184 1447 1187 1451
rect 1215 1447 1216 1451
rect 1216 1447 1219 1451
rect 1239 1454 1243 1458
rect 1279 1453 1283 1457
rect 1319 1454 1323 1458
rect 1359 1454 1363 1458
rect 1299 1447 1300 1451
rect 1300 1447 1303 1451
rect 1335 1447 1336 1451
rect 1336 1447 1339 1451
rect 1375 1447 1376 1451
rect 1376 1447 1379 1451
rect 1399 1454 1403 1458
rect 1459 1463 1460 1467
rect 1460 1463 1463 1467
rect 1439 1454 1443 1458
rect 1479 1454 1483 1458
rect 1499 1447 1500 1451
rect 1500 1447 1503 1451
rect 1551 1463 1555 1467
rect 1575 1463 1576 1467
rect 1576 1463 1579 1467
rect 1519 1454 1523 1458
rect 1559 1454 1563 1458
rect 1591 1454 1595 1458
rect 1623 1454 1627 1458
rect 1655 1454 1659 1458
rect 1639 1447 1640 1451
rect 1640 1447 1643 1451
rect 1671 1463 1672 1467
rect 1672 1463 1675 1467
rect 1695 1452 1699 1456
rect 991 1427 995 1431
rect 999 1427 1003 1431
rect 1031 1431 1035 1435
rect 1047 1435 1048 1439
rect 1048 1435 1051 1439
rect 1191 1439 1195 1443
rect 1671 1439 1675 1443
rect 1703 1431 1707 1435
rect 751 1419 755 1423
rect 795 1421 799 1423
rect 795 1419 796 1421
rect 796 1419 799 1421
rect 831 1419 835 1423
rect 767 1411 771 1415
rect 839 1411 843 1415
rect 879 1415 883 1419
rect 903 1415 904 1419
rect 904 1415 907 1419
rect 919 1415 920 1419
rect 920 1415 923 1419
rect 947 1419 951 1423
rect 1191 1423 1195 1427
rect 967 1411 971 1415
rect 975 1411 979 1415
rect 991 1415 995 1419
rect 1047 1411 1051 1415
rect 1123 1415 1127 1419
rect 1215 1415 1219 1419
rect 447 1399 451 1403
rect 111 1388 115 1392
rect 151 1391 152 1395
rect 152 1391 155 1395
rect 135 1386 139 1390
rect 167 1386 171 1390
rect 199 1386 203 1390
rect 231 1386 235 1390
rect 263 1386 267 1390
rect 295 1386 299 1390
rect 327 1386 331 1390
rect 379 1391 380 1395
rect 380 1391 383 1395
rect 359 1386 363 1390
rect 391 1386 395 1390
rect 423 1386 427 1390
rect 455 1386 459 1390
rect 543 1399 547 1403
rect 487 1386 491 1390
rect 519 1386 523 1390
rect 551 1386 555 1390
rect 759 1403 763 1407
rect 895 1406 899 1410
rect 1071 1403 1075 1407
rect 583 1386 587 1390
rect 615 1386 619 1390
rect 647 1386 651 1390
rect 695 1391 696 1395
rect 696 1391 699 1395
rect 679 1386 683 1390
rect 719 1389 723 1393
rect 763 1391 767 1395
rect 807 1391 811 1395
rect 787 1383 791 1387
rect 867 1383 868 1387
rect 868 1383 871 1387
rect 1063 1396 1067 1400
rect 1151 1396 1155 1400
rect 1215 1403 1219 1407
rect 1231 1407 1235 1411
rect 1471 1419 1475 1423
rect 999 1391 1003 1395
rect 1191 1395 1195 1399
rect 1459 1413 1463 1415
rect 1459 1411 1460 1413
rect 1460 1411 1463 1413
rect 1055 1391 1059 1395
rect 111 1371 115 1375
rect 347 1375 348 1379
rect 348 1375 351 1379
rect 471 1375 472 1379
rect 472 1375 475 1379
rect 567 1376 568 1379
rect 568 1376 571 1379
rect 567 1375 571 1376
rect 663 1375 664 1379
rect 664 1375 667 1379
rect 135 1369 139 1373
rect 167 1369 171 1373
rect 199 1369 203 1373
rect 231 1369 235 1373
rect 263 1369 267 1373
rect 295 1369 299 1373
rect 327 1369 331 1373
rect 359 1369 363 1373
rect 391 1369 395 1373
rect 423 1369 427 1373
rect 455 1369 459 1373
rect 487 1369 491 1373
rect 519 1369 523 1373
rect 551 1369 555 1373
rect 583 1369 587 1373
rect 615 1369 619 1373
rect 647 1369 651 1373
rect 679 1369 683 1373
rect 379 1363 383 1367
rect 567 1363 571 1367
rect 735 1362 739 1366
rect 767 1364 771 1368
rect 807 1368 811 1372
rect 847 1375 851 1379
rect 947 1379 951 1383
rect 967 1383 971 1387
rect 1023 1386 1027 1390
rect 1071 1379 1075 1383
rect 1103 1383 1107 1387
rect 1111 1387 1115 1391
rect 1131 1391 1132 1395
rect 1132 1391 1135 1395
rect 1471 1403 1475 1407
rect 1407 1395 1411 1399
rect 1167 1383 1171 1387
rect 1199 1386 1203 1390
rect 1263 1389 1267 1393
rect 1319 1387 1323 1391
rect 1415 1386 1419 1390
rect 1479 1389 1483 1393
rect 1487 1387 1491 1391
rect 1551 1391 1552 1395
rect 1552 1391 1555 1395
rect 1575 1395 1579 1399
rect 1535 1386 1539 1390
rect 1583 1386 1587 1390
rect 1623 1386 1627 1390
rect 1655 1386 1659 1390
rect 1123 1375 1127 1379
rect 1215 1375 1216 1379
rect 1216 1375 1219 1379
rect 1299 1379 1303 1383
rect 1695 1388 1699 1392
rect 1447 1375 1451 1379
rect 1547 1375 1551 1379
rect 839 1364 843 1368
rect 887 1368 891 1372
rect 1023 1369 1027 1373
rect 1063 1368 1067 1372
rect 1111 1369 1115 1373
rect 1151 1368 1155 1372
rect 1199 1369 1203 1373
rect 1247 1368 1251 1372
rect 975 1364 979 1368
rect 1319 1368 1323 1372
rect 1415 1369 1419 1373
rect 1463 1368 1467 1372
rect 1535 1369 1539 1373
rect 1583 1369 1587 1373
rect 1623 1369 1627 1373
rect 1655 1369 1659 1373
rect 1575 1363 1579 1367
rect 1695 1371 1699 1375
rect 687 1355 691 1359
rect 815 1351 819 1355
rect 951 1351 955 1355
rect 1123 1351 1127 1355
rect 1487 1351 1491 1355
rect 1167 1339 1171 1343
rect 179 1331 183 1335
rect 1239 1331 1243 1335
rect 111 1313 115 1317
rect 135 1315 139 1319
rect 167 1315 171 1319
rect 199 1315 203 1319
rect 231 1315 235 1319
rect 263 1315 267 1319
rect 295 1315 299 1319
rect 327 1315 331 1319
rect 359 1315 363 1319
rect 391 1315 395 1319
rect 423 1315 427 1319
rect 455 1315 459 1319
rect 487 1315 491 1319
rect 519 1315 523 1319
rect 551 1315 555 1319
rect 583 1315 587 1319
rect 615 1315 619 1319
rect 647 1315 651 1319
rect 679 1315 683 1319
rect 711 1315 715 1319
rect 743 1316 747 1320
rect 823 1316 827 1320
rect 903 1316 907 1320
rect 983 1320 987 1324
rect 1023 1316 1027 1320
rect 1063 1316 1067 1320
rect 1159 1316 1163 1320
rect 1215 1316 1219 1320
rect 1303 1316 1307 1320
rect 1391 1315 1395 1319
rect 1423 1315 1427 1319
rect 1455 1316 1459 1320
rect 1495 1315 1499 1319
rect 1527 1315 1531 1319
rect 1559 1315 1563 1319
rect 1591 1315 1595 1319
rect 1623 1315 1627 1319
rect 1655 1315 1659 1319
rect 1695 1313 1699 1317
rect 151 1307 152 1311
rect 152 1307 155 1311
rect 111 1296 115 1300
rect 135 1298 139 1302
rect 167 1298 171 1302
rect 199 1298 203 1302
rect 231 1298 235 1302
rect 263 1298 267 1302
rect 295 1298 299 1302
rect 327 1298 331 1302
rect 347 1299 351 1303
rect 359 1298 363 1302
rect 391 1298 395 1302
rect 423 1298 427 1302
rect 455 1298 459 1302
rect 487 1298 491 1302
rect 519 1298 523 1302
rect 551 1298 555 1302
rect 583 1298 587 1302
rect 627 1307 631 1311
rect 615 1298 619 1302
rect 647 1298 651 1302
rect 695 1307 696 1311
rect 696 1307 699 1311
rect 679 1298 683 1302
rect 711 1298 715 1302
rect 663 1291 664 1295
rect 664 1291 667 1295
rect 751 1303 755 1307
rect 831 1303 835 1307
rect 971 1307 975 1311
rect 1131 1307 1135 1311
rect 1287 1307 1291 1311
rect 1411 1307 1412 1311
rect 1412 1307 1415 1311
rect 1435 1307 1439 1311
rect 1483 1307 1487 1311
rect 1539 1307 1543 1311
rect 963 1299 967 1303
rect 1023 1288 1027 1292
rect 471 1283 475 1287
rect 187 1275 191 1279
rect 735 1275 739 1279
rect 751 1278 755 1282
rect 831 1278 835 1282
rect 911 1278 915 1282
rect 983 1273 987 1277
rect 1039 1275 1043 1279
rect 1063 1297 1067 1301
rect 1175 1295 1179 1299
rect 1215 1297 1219 1301
rect 1303 1297 1307 1301
rect 103 1267 107 1271
rect 575 1267 579 1271
rect 759 1267 760 1271
rect 760 1267 763 1271
rect 787 1267 791 1271
rect 839 1267 840 1271
rect 840 1267 843 1271
rect 867 1267 871 1271
rect 895 1267 899 1271
rect 931 1267 935 1271
rect 963 1267 967 1271
rect 735 1259 739 1263
rect 607 1251 611 1255
rect 759 1251 763 1255
rect 839 1251 843 1255
rect 887 1251 891 1255
rect 971 1263 975 1267
rect 1111 1275 1115 1279
rect 1139 1275 1143 1279
rect 1155 1275 1156 1279
rect 1156 1275 1159 1279
rect 1191 1279 1195 1283
rect 1391 1297 1395 1301
rect 1423 1298 1427 1302
rect 1495 1298 1499 1302
rect 1527 1298 1531 1302
rect 1559 1298 1563 1302
rect 1591 1298 1595 1302
rect 1439 1291 1440 1295
rect 1440 1291 1443 1295
rect 1455 1288 1459 1292
rect 1515 1291 1516 1295
rect 1516 1291 1519 1295
rect 1547 1291 1548 1295
rect 1548 1291 1551 1295
rect 1575 1291 1576 1295
rect 1576 1291 1579 1295
rect 1623 1298 1627 1302
rect 1655 1298 1659 1302
rect 1671 1307 1672 1311
rect 1672 1307 1675 1311
rect 1695 1296 1699 1300
rect 1287 1279 1291 1283
rect 1411 1283 1415 1287
rect 1439 1283 1443 1287
rect 1447 1283 1451 1287
rect 1471 1275 1475 1279
rect 1483 1279 1484 1283
rect 1484 1279 1487 1283
rect 1199 1267 1203 1271
rect 1055 1259 1059 1263
rect 991 1251 995 1255
rect 919 1243 923 1247
rect 191 1231 195 1235
rect 899 1231 903 1235
rect 655 1223 659 1227
rect 591 1211 595 1215
rect 627 1211 631 1215
rect 775 1215 779 1219
rect 795 1219 799 1223
rect 847 1223 851 1227
rect 991 1227 995 1231
rect 111 1192 115 1196
rect 151 1195 152 1199
rect 152 1195 155 1199
rect 135 1190 139 1194
rect 167 1190 171 1194
rect 199 1190 203 1194
rect 231 1190 235 1194
rect 263 1190 267 1194
rect 295 1190 299 1194
rect 327 1190 331 1194
rect 359 1190 363 1194
rect 391 1190 395 1194
rect 423 1190 427 1194
rect 455 1190 459 1194
rect 487 1190 491 1194
rect 599 1203 603 1207
rect 759 1207 763 1211
rect 791 1211 795 1215
rect 1039 1219 1040 1223
rect 1040 1219 1043 1223
rect 1067 1223 1071 1227
rect 1079 1215 1083 1219
rect 1087 1215 1091 1219
rect 1103 1219 1107 1223
rect 1191 1219 1195 1223
rect 1447 1219 1451 1223
rect 1015 1210 1019 1214
rect 1199 1211 1200 1215
rect 1200 1211 1203 1215
rect 519 1190 523 1194
rect 551 1190 555 1194
rect 591 1195 595 1199
rect 583 1190 587 1194
rect 615 1190 619 1194
rect 647 1190 651 1194
rect 679 1190 683 1194
rect 111 1175 115 1179
rect 567 1179 568 1183
rect 568 1179 571 1183
rect 599 1179 600 1183
rect 600 1179 603 1183
rect 711 1190 715 1194
rect 823 1199 827 1203
rect 951 1203 955 1207
rect 1191 1203 1195 1207
rect 1263 1203 1267 1207
rect 1455 1211 1459 1215
rect 743 1190 747 1194
rect 791 1187 795 1191
rect 811 1191 815 1195
rect 959 1193 963 1197
rect 991 1195 992 1199
rect 992 1195 995 1199
rect 759 1179 760 1183
rect 760 1179 763 1183
rect 1067 1183 1071 1187
rect 1079 1187 1083 1191
rect 1127 1190 1131 1194
rect 1159 1190 1163 1194
rect 135 1173 139 1177
rect 167 1173 171 1177
rect 199 1173 203 1177
rect 231 1173 235 1177
rect 263 1173 267 1177
rect 295 1173 299 1177
rect 327 1173 331 1177
rect 359 1173 363 1177
rect 391 1173 395 1177
rect 423 1173 427 1177
rect 455 1173 459 1177
rect 487 1173 491 1177
rect 443 1167 447 1171
rect 519 1173 523 1177
rect 551 1173 555 1177
rect 583 1173 587 1177
rect 615 1173 619 1177
rect 647 1173 651 1177
rect 679 1173 683 1177
rect 711 1173 715 1177
rect 743 1173 747 1177
rect 839 1176 843 1180
rect 931 1175 935 1179
rect 1143 1179 1144 1183
rect 1144 1179 1147 1183
rect 1199 1195 1203 1199
rect 1215 1193 1219 1197
rect 1239 1191 1240 1195
rect 1240 1191 1243 1195
rect 1255 1190 1259 1194
rect 1295 1193 1299 1197
rect 1351 1199 1355 1203
rect 1415 1203 1419 1207
rect 1343 1190 1347 1194
rect 1375 1190 1379 1194
rect 1424 1195 1428 1199
rect 1407 1190 1411 1194
rect 1439 1190 1443 1194
rect 1499 1195 1500 1199
rect 1500 1195 1503 1199
rect 1539 1195 1540 1199
rect 1540 1195 1543 1199
rect 1547 1199 1551 1203
rect 1479 1190 1483 1194
rect 1519 1190 1523 1194
rect 1559 1190 1563 1194
rect 1591 1190 1595 1194
rect 1623 1190 1627 1194
rect 1287 1179 1291 1183
rect 775 1168 779 1172
rect 1007 1172 1011 1176
rect 1127 1173 1131 1177
rect 1159 1173 1163 1177
rect 1199 1172 1203 1176
rect 1255 1173 1259 1177
rect 1343 1173 1347 1177
rect 1375 1173 1379 1177
rect 975 1166 979 1170
rect 1087 1168 1091 1172
rect 1311 1166 1315 1170
rect 1419 1179 1423 1183
rect 1455 1179 1456 1183
rect 1456 1179 1459 1183
rect 1547 1179 1551 1183
rect 1575 1179 1576 1183
rect 1576 1179 1579 1183
rect 1611 1179 1612 1183
rect 1612 1179 1615 1183
rect 1671 1195 1672 1199
rect 1672 1195 1675 1199
rect 1655 1190 1659 1194
rect 1695 1192 1699 1196
rect 1407 1173 1411 1177
rect 1439 1173 1443 1177
rect 1479 1173 1483 1177
rect 1519 1173 1523 1177
rect 1559 1173 1563 1177
rect 1591 1173 1595 1177
rect 1623 1173 1627 1177
rect 1655 1173 1659 1177
rect 1695 1175 1699 1179
rect 1431 1167 1435 1171
rect 1447 1167 1451 1171
rect 543 1159 547 1163
rect 799 1159 803 1163
rect 815 1159 819 1163
rect 1287 1159 1288 1163
rect 1288 1159 1291 1163
rect 415 1147 419 1151
rect 955 1139 959 1143
rect 1143 1139 1147 1143
rect 283 1127 287 1131
rect 111 1117 115 1121
rect 135 1119 139 1123
rect 167 1119 171 1123
rect 199 1119 203 1123
rect 231 1119 235 1123
rect 263 1119 267 1123
rect 295 1119 299 1123
rect 327 1119 331 1123
rect 359 1119 363 1123
rect 391 1119 395 1123
rect 423 1119 427 1123
rect 455 1119 459 1123
rect 487 1119 491 1123
rect 519 1119 523 1123
rect 111 1100 115 1104
rect 135 1102 139 1106
rect 167 1102 171 1106
rect 199 1102 203 1106
rect 231 1102 235 1106
rect 247 1111 248 1115
rect 248 1111 251 1115
rect 263 1102 267 1106
rect 295 1102 299 1106
rect 327 1102 331 1106
rect 283 1095 284 1099
rect 284 1095 287 1099
rect 359 1102 363 1106
rect 391 1102 395 1106
rect 423 1102 427 1106
rect 455 1102 459 1106
rect 443 1095 444 1099
rect 444 1095 447 1099
rect 487 1102 491 1106
rect 519 1102 523 1106
rect 535 1111 536 1115
rect 536 1111 539 1115
rect 551 1119 555 1123
rect 583 1120 587 1124
rect 799 1120 803 1124
rect 847 1122 851 1126
rect 687 1116 691 1120
rect 783 1115 784 1119
rect 784 1115 787 1119
rect 655 1111 659 1115
rect 855 1115 859 1119
rect 935 1119 939 1123
rect 967 1119 971 1123
rect 999 1120 1003 1124
rect 551 1102 555 1106
rect 659 1101 663 1105
rect 935 1102 939 1106
rect 967 1102 971 1106
rect 567 1095 568 1099
rect 568 1095 571 1099
rect 799 1097 803 1101
rect 535 1087 539 1091
rect 703 1091 707 1095
rect 955 1095 956 1099
rect 956 1095 959 1099
rect 1015 1115 1016 1119
rect 1016 1115 1019 1119
rect 1031 1119 1035 1123
rect 1063 1119 1067 1123
rect 1095 1120 1099 1124
rect 1135 1119 1139 1123
rect 1167 1120 1171 1124
rect 1247 1124 1251 1128
rect 1287 1119 1291 1123
rect 1335 1122 1339 1126
rect 1423 1119 1427 1123
rect 1455 1119 1459 1123
rect 1487 1119 1491 1123
rect 1519 1119 1523 1123
rect 1559 1119 1563 1123
rect 1591 1119 1595 1123
rect 1623 1119 1627 1123
rect 1655 1119 1659 1123
rect 1695 1117 1699 1121
rect 999 1097 1003 1101
rect 1031 1102 1035 1106
rect 1063 1102 1067 1106
rect 1083 1111 1084 1115
rect 1084 1111 1087 1115
rect 1123 1111 1127 1115
rect 1235 1111 1239 1115
rect 1279 1111 1283 1115
rect 1111 1103 1115 1107
rect 1135 1102 1139 1106
rect 1227 1103 1231 1107
rect 1287 1102 1291 1106
rect 1095 1092 1099 1096
rect 1423 1102 1427 1106
rect 1455 1102 1459 1106
rect 1431 1095 1435 1099
rect 1471 1111 1472 1115
rect 1472 1111 1475 1115
rect 1499 1111 1503 1115
rect 1535 1111 1536 1115
rect 1536 1111 1539 1115
rect 1487 1102 1491 1106
rect 1519 1102 1523 1106
rect 307 1079 311 1083
rect 591 1082 595 1086
rect 847 1081 851 1085
rect 191 1071 195 1075
rect 599 1071 600 1075
rect 600 1071 603 1075
rect 791 1075 795 1079
rect 923 1077 927 1079
rect 607 1063 611 1067
rect 823 1067 827 1071
rect 863 1071 864 1075
rect 864 1071 867 1075
rect 923 1075 924 1077
rect 924 1075 927 1077
rect 1103 1079 1107 1083
rect 1123 1083 1124 1087
rect 1124 1083 1127 1087
rect 1559 1102 1563 1106
rect 1591 1102 1595 1106
rect 1611 1103 1615 1107
rect 1575 1095 1576 1099
rect 1576 1095 1579 1099
rect 1623 1102 1627 1106
rect 1655 1102 1659 1106
rect 1671 1111 1672 1115
rect 1672 1111 1675 1115
rect 1695 1100 1699 1104
rect 1671 1087 1675 1091
rect 1175 1082 1179 1086
rect 1247 1077 1251 1081
rect 1335 1081 1339 1085
rect 1195 1071 1199 1075
rect 1227 1071 1231 1075
rect 1235 1067 1239 1071
rect 1263 1071 1267 1075
rect 1351 1071 1352 1075
rect 1352 1071 1355 1075
rect 1447 1071 1451 1075
rect 1039 1059 1043 1063
rect 915 1051 919 1055
rect 399 1019 400 1023
rect 400 1019 403 1023
rect 415 1019 416 1023
rect 416 1019 419 1023
rect 459 1019 463 1023
rect 495 1023 499 1027
rect 503 1015 507 1019
rect 543 1019 547 1023
rect 615 1019 619 1023
rect 659 1019 660 1023
rect 660 1019 663 1023
rect 831 1027 835 1031
rect 863 1027 867 1031
rect 783 1019 784 1023
rect 784 1019 787 1023
rect 407 1010 411 1014
rect 583 1011 587 1015
rect 711 1011 715 1015
rect 843 1015 847 1019
rect 855 1015 856 1019
rect 856 1015 859 1019
rect 1015 1019 1019 1023
rect 1047 1015 1051 1019
rect 247 1003 251 1007
rect 383 1003 387 1007
rect 575 1003 579 1007
rect 823 1005 827 1009
rect 975 1005 979 1009
rect 1075 1007 1079 1011
rect 1183 1011 1187 1015
rect 1263 1015 1267 1019
rect 1063 1000 1067 1004
rect 1191 1003 1195 1007
rect 1207 1007 1211 1011
rect 1199 1000 1203 1004
rect 1279 1003 1283 1007
rect 1335 1007 1339 1011
rect 1455 1007 1459 1011
rect 1327 1000 1331 1004
rect 111 992 115 996
rect 135 990 139 994
rect 167 990 171 994
rect 111 975 115 979
rect 151 979 152 983
rect 152 979 155 983
rect 199 990 203 994
rect 231 990 235 994
rect 263 990 267 994
rect 327 993 331 997
rect 359 995 360 999
rect 360 995 363 999
rect 459 991 463 995
rect 319 979 323 983
rect 495 983 499 987
rect 531 987 532 991
rect 532 987 535 991
rect 919 990 923 994
rect 1119 993 1123 997
rect 1167 990 1171 994
rect 1247 993 1251 997
rect 1367 1000 1371 1004
rect 135 973 139 977
rect 167 973 171 977
rect 199 973 203 977
rect 231 973 235 977
rect 263 973 267 977
rect 399 972 403 976
rect 823 975 827 979
rect 935 979 936 983
rect 936 979 939 983
rect 1207 983 1211 987
rect 1295 990 1299 994
rect 1335 983 1339 987
rect 1383 987 1387 991
rect 1471 995 1475 999
rect 1535 995 1536 999
rect 1536 995 1539 999
rect 1407 990 1411 994
rect 1439 990 1443 994
rect 1479 990 1483 994
rect 1519 990 1523 994
rect 1559 990 1563 994
rect 1427 979 1428 983
rect 1428 979 1431 983
rect 1455 979 1456 983
rect 1456 979 1459 983
rect 1495 979 1496 983
rect 1496 979 1499 983
rect 1591 990 1595 994
rect 1623 990 1627 994
rect 1655 990 1659 994
rect 1695 992 1699 996
rect 343 966 347 970
rect 503 968 507 972
rect 583 970 587 974
rect 711 970 715 974
rect 919 973 923 977
rect 1063 972 1067 976
rect 1167 973 1171 977
rect 1199 972 1203 976
rect 1295 973 1299 977
rect 1327 972 1331 976
rect 1367 972 1371 976
rect 1407 973 1411 977
rect 1439 973 1443 977
rect 1479 973 1483 977
rect 1519 973 1523 977
rect 1559 973 1563 977
rect 1591 973 1595 977
rect 1623 973 1627 977
rect 1655 973 1659 977
rect 815 965 819 969
rect 967 965 971 969
rect 1135 966 1139 970
rect 1263 966 1267 970
rect 1539 967 1543 971
rect 1695 975 1699 979
rect 319 959 320 963
rect 320 959 323 963
rect 1083 959 1087 963
rect 219 951 223 955
rect 599 951 603 955
rect 659 951 663 955
rect 855 951 859 955
rect 339 939 343 943
rect 415 939 419 943
rect 1195 941 1196 943
rect 1196 941 1199 943
rect 1399 943 1403 947
rect 1195 939 1199 941
rect 111 917 115 921
rect 135 919 139 923
rect 167 919 171 923
rect 199 920 203 924
rect 279 924 283 928
rect 319 920 323 924
rect 399 924 403 928
rect 991 927 995 931
rect 1123 931 1127 935
rect 591 922 595 926
rect 679 920 683 924
rect 727 922 731 926
rect 463 916 467 920
rect 187 911 188 915
rect 188 911 191 915
rect 267 911 271 915
rect 387 911 391 915
rect 599 915 603 919
rect 695 915 696 919
rect 696 915 699 919
rect 815 919 819 923
rect 863 922 867 926
rect 951 919 955 923
rect 983 920 987 924
rect 1039 919 1043 923
rect 1071 920 1075 924
rect 803 911 807 915
rect 971 911 972 915
rect 972 911 975 915
rect 1095 911 1099 915
rect 1391 926 1395 930
rect 1111 919 1115 923
rect 1143 920 1147 924
rect 1239 919 1243 923
rect 1271 920 1275 924
rect 1423 919 1427 923
rect 1455 920 1459 924
rect 1519 919 1523 923
rect 1559 919 1563 923
rect 1591 919 1595 923
rect 1623 919 1627 923
rect 1655 919 1659 923
rect 1695 917 1699 921
rect 111 900 115 904
rect 135 902 139 906
rect 167 902 171 906
rect 259 903 263 907
rect 427 903 428 907
rect 428 903 431 907
rect 435 901 439 905
rect 815 902 819 906
rect 951 902 955 906
rect 151 895 152 899
rect 152 895 155 899
rect 183 895 184 899
rect 184 895 187 899
rect 679 897 683 901
rect 523 891 527 895
rect 607 891 611 895
rect 823 895 827 899
rect 855 891 859 895
rect 991 895 995 899
rect 999 899 1003 903
rect 1039 902 1043 906
rect 1071 892 1075 896
rect 1111 901 1115 905
rect 1231 911 1235 915
rect 1143 901 1147 905
rect 1239 901 1243 905
rect 1207 895 1211 899
rect 1355 907 1359 911
rect 1271 901 1275 905
rect 1375 899 1379 903
rect 1423 902 1427 906
rect 1399 895 1403 899
rect 1431 895 1435 899
rect 1471 899 1475 903
rect 1519 902 1523 906
rect 1559 902 1563 906
rect 1539 895 1540 899
rect 1540 895 1543 899
rect 1591 902 1595 906
rect 1623 902 1627 906
rect 1655 902 1659 906
rect 1671 911 1672 915
rect 1672 911 1675 915
rect 1695 900 1699 904
rect 207 882 211 886
rect 327 882 331 886
rect 279 877 283 881
rect 399 877 403 881
rect 591 881 595 885
rect 727 881 731 885
rect 863 881 867 885
rect 219 871 220 875
rect 220 871 223 875
rect 259 871 263 875
rect 267 867 271 871
rect 307 871 308 875
rect 308 871 311 875
rect 339 871 340 875
rect 340 871 343 875
rect 259 859 263 863
rect 387 867 391 871
rect 415 871 419 875
rect 543 875 547 879
rect 971 879 975 883
rect 1047 883 1051 887
rect 1079 883 1083 887
rect 1095 883 1096 887
rect 1096 883 1099 887
rect 1207 879 1208 883
rect 1208 879 1211 883
rect 1355 887 1359 891
rect 1415 887 1419 891
rect 608 871 612 875
rect 803 871 804 875
rect 804 871 807 875
rect 427 859 431 863
rect 703 863 707 867
rect 747 863 751 867
rect 935 871 936 875
rect 936 871 939 875
rect 1383 879 1387 883
rect 1479 883 1480 887
rect 1480 883 1483 887
rect 1663 879 1667 883
rect 307 851 311 855
rect 415 851 419 855
rect 531 851 535 855
rect 599 855 603 859
rect 887 855 891 859
rect 303 835 307 839
rect 359 835 363 839
rect 607 835 611 839
rect 851 839 855 843
rect 1255 835 1259 839
rect 1479 835 1483 839
rect 427 827 428 831
rect 428 827 431 831
rect 575 827 579 831
rect 231 819 235 823
rect 407 819 411 823
rect 695 823 696 827
rect 696 823 699 827
rect 831 827 832 831
rect 832 827 835 831
rect 887 827 888 831
rect 888 827 891 831
rect 1279 827 1283 831
rect 815 819 819 823
rect 991 819 995 823
rect 663 813 667 817
rect 1231 819 1232 823
rect 1232 819 1235 823
rect 1255 815 1256 819
rect 1256 815 1259 819
rect 1355 811 1359 815
rect 111 800 115 804
rect 135 798 139 802
rect 559 798 563 802
rect 951 803 955 807
rect 1031 801 1035 805
rect 1043 799 1047 803
rect 1111 803 1115 807
rect 1055 799 1056 803
rect 1056 799 1059 803
rect 1123 803 1124 807
rect 1124 803 1127 807
rect 1103 798 1107 802
rect 1167 801 1171 805
rect 1195 803 1199 807
rect 1247 801 1251 805
rect 1279 799 1283 803
rect 1295 799 1299 803
rect 1415 819 1419 823
rect 1479 819 1483 823
rect 1495 815 1496 819
rect 1496 815 1499 819
rect 111 783 115 787
rect 151 787 152 791
rect 152 787 155 791
rect 575 787 576 791
rect 576 787 579 791
rect 135 781 139 785
rect 231 778 235 782
rect 407 778 411 782
rect 559 781 563 785
rect 815 778 819 782
rect 951 780 955 784
rect 1159 787 1163 791
rect 1271 791 1275 795
rect 1327 799 1331 803
rect 1423 808 1427 812
rect 1471 808 1475 812
rect 1519 798 1523 802
rect 1559 798 1563 802
rect 1591 798 1595 802
rect 1623 798 1627 802
rect 1655 798 1659 802
rect 1671 803 1672 807
rect 1672 803 1675 807
rect 1695 800 1699 804
rect 655 773 659 777
rect 1015 780 1019 784
rect 1103 781 1107 785
rect 1231 780 1235 784
rect 1295 781 1299 785
rect 1327 780 1331 784
rect 1423 780 1427 784
rect 1471 780 1475 784
rect 1519 781 1523 785
rect 1035 771 1039 775
rect 1183 774 1187 778
rect 1499 775 1503 779
rect 1559 781 1563 785
rect 1591 781 1595 785
rect 1623 781 1627 785
rect 1655 781 1659 785
rect 1695 783 1699 787
rect 1159 767 1160 771
rect 1160 767 1163 771
rect 219 759 223 763
rect 1223 755 1227 759
rect 111 721 115 725
rect 135 724 139 728
rect 215 728 219 732
rect 287 726 291 730
rect 391 728 395 732
rect 767 731 771 735
rect 999 731 1003 735
rect 615 726 619 730
rect 719 724 723 728
rect 471 720 475 724
rect 203 715 207 719
rect 623 719 627 723
rect 767 719 771 723
rect 863 723 867 727
rect 911 726 915 730
rect 1087 724 1091 728
rect 1167 728 1171 732
rect 843 715 847 719
rect 1207 724 1211 728
rect 1247 723 1251 727
rect 1279 723 1283 727
rect 1311 723 1315 727
rect 1343 723 1347 727
rect 1375 723 1379 727
rect 1407 723 1411 727
rect 1439 723 1443 727
rect 1479 723 1483 727
rect 1519 723 1523 727
rect 1559 723 1563 727
rect 1591 723 1595 727
rect 1623 723 1627 727
rect 1655 723 1659 727
rect 1695 721 1699 725
rect 111 704 115 708
rect 243 707 244 711
rect 244 707 247 711
rect 419 707 420 711
rect 420 707 423 711
rect 443 705 447 709
rect 731 707 735 711
rect 863 706 867 710
rect 719 701 723 705
rect 279 695 283 699
rect 567 695 568 699
rect 568 695 571 699
rect 1155 715 1159 719
rect 1235 715 1239 719
rect 1147 707 1151 711
rect 1223 707 1227 711
rect 1247 706 1251 710
rect 1279 706 1283 710
rect 143 686 147 690
rect 191 683 195 687
rect 215 681 219 685
rect 287 685 291 689
rect 203 671 207 675
rect 235 675 239 679
rect 303 675 304 679
rect 304 675 307 679
rect 323 675 327 679
rect 775 691 779 695
rect 1207 696 1211 700
rect 1227 699 1231 703
rect 1311 706 1315 710
rect 1343 706 1347 710
rect 1375 706 1379 710
rect 1407 706 1411 710
rect 1439 706 1443 710
rect 1479 706 1483 710
rect 1447 699 1451 703
rect 1499 699 1500 703
rect 1500 699 1503 703
rect 1519 706 1523 710
rect 1559 706 1563 710
rect 1591 706 1595 710
rect 1623 706 1627 710
rect 1655 706 1659 710
rect 1671 715 1672 719
rect 1672 715 1675 719
rect 1695 704 1699 708
rect 391 681 395 685
rect 615 685 619 689
rect 399 671 403 675
rect 411 675 415 679
rect 427 679 431 683
rect 523 671 527 675
rect 555 675 559 679
rect 747 683 751 687
rect 851 687 855 691
rect 1007 691 1011 695
rect 911 685 915 689
rect 1095 686 1099 690
rect 759 679 763 683
rect 243 663 247 667
rect 315 663 319 667
rect 411 663 415 667
rect 419 663 423 667
rect 459 663 463 667
rect 767 671 771 675
rect 831 675 835 679
rect 983 675 984 679
rect 984 675 987 679
rect 1015 679 1016 683
rect 1016 679 1019 683
rect 1035 679 1036 683
rect 1036 679 1039 683
rect 1167 681 1171 685
rect 1235 687 1236 691
rect 1236 687 1239 691
rect 1455 687 1459 691
rect 1087 675 1088 679
rect 1088 675 1091 679
rect 1103 675 1104 679
rect 1104 675 1107 679
rect 1147 675 1151 679
rect 843 663 847 667
rect 1063 667 1067 671
rect 1155 671 1159 675
rect 1183 675 1187 679
rect 1255 675 1259 679
rect 1359 675 1363 679
rect 243 655 247 659
rect 851 659 855 663
rect 1015 659 1019 663
rect 1111 659 1115 663
rect 1103 651 1107 655
rect 1175 655 1179 659
rect 235 643 239 647
rect 315 643 319 647
rect 295 635 299 639
rect 339 635 343 639
rect 635 635 639 639
rect 1079 639 1083 643
rect 207 623 211 627
rect 235 627 236 631
rect 236 627 239 631
rect 279 627 280 631
rect 280 627 283 631
rect 307 627 311 631
rect 415 627 416 631
rect 416 627 419 631
rect 459 627 463 631
rect 519 627 523 631
rect 555 627 556 631
rect 556 627 559 631
rect 687 627 691 631
rect 919 631 923 635
rect 287 618 291 622
rect 407 618 411 622
rect 535 619 539 623
rect 767 619 771 623
rect 831 619 835 623
rect 903 623 907 627
rect 951 627 955 631
rect 983 627 987 631
rect 1007 627 1008 631
rect 1008 627 1011 631
rect 1051 631 1055 635
rect 1183 635 1187 639
rect 1111 623 1115 627
rect 1119 623 1123 627
rect 1143 627 1144 631
rect 1144 627 1147 631
rect 1223 627 1224 631
rect 1224 627 1227 631
rect 1267 631 1271 635
rect 999 618 1003 622
rect 1215 618 1219 622
rect 1335 623 1339 627
rect 1359 627 1360 631
rect 1360 627 1363 631
rect 111 600 115 604
rect 151 603 152 607
rect 152 603 155 607
rect 255 603 259 607
rect 527 607 531 611
rect 759 611 763 615
rect 1347 615 1351 619
rect 1671 615 1675 619
rect 731 603 735 607
rect 135 598 139 602
rect 167 598 171 602
rect 287 595 291 599
rect 671 598 675 602
rect 1435 603 1436 607
rect 1436 603 1439 607
rect 111 583 115 587
rect 151 587 152 591
rect 152 587 155 591
rect 183 587 184 591
rect 184 587 187 591
rect 295 591 299 595
rect 399 591 403 595
rect 959 595 963 599
rect 687 587 688 591
rect 688 587 691 591
rect 1051 591 1055 595
rect 1111 595 1115 599
rect 1267 591 1271 595
rect 1347 595 1351 599
rect 1415 598 1419 602
rect 1479 598 1483 602
rect 1543 598 1547 602
rect 1607 598 1611 602
rect 1655 598 1659 602
rect 1695 600 1699 604
rect 1447 587 1451 591
rect 1671 587 1672 591
rect 1672 587 1675 591
rect 135 581 139 585
rect 167 581 171 585
rect 207 576 211 580
rect 279 580 283 584
rect 399 580 403 584
rect 535 578 539 582
rect 671 581 675 585
rect 767 578 771 582
rect 903 576 907 580
rect 991 580 995 584
rect 1119 576 1123 580
rect 1207 580 1211 584
rect 1415 581 1419 585
rect 1479 581 1483 585
rect 1543 581 1547 585
rect 1607 581 1611 585
rect 1655 581 1659 585
rect 1695 583 1699 587
rect 1335 576 1339 580
rect 379 559 383 563
rect 527 559 531 563
rect 795 559 799 563
rect 1007 559 1011 563
rect 1103 563 1107 567
rect 1223 563 1227 567
rect 111 529 115 533
rect 135 531 139 535
rect 167 532 171 536
rect 247 536 251 540
rect 303 534 307 538
rect 391 532 395 536
rect 471 536 475 540
rect 647 532 651 536
rect 727 536 731 540
rect 535 528 539 532
rect 235 523 239 527
rect 775 532 779 536
rect 871 536 875 540
rect 927 532 931 536
rect 1031 536 1035 540
rect 1095 532 1099 536
rect 1199 536 1203 540
rect 635 527 636 531
rect 636 527 639 531
rect 1287 528 1291 532
rect 459 523 463 527
rect 715 523 719 527
rect 843 523 847 527
rect 919 523 923 527
rect 1379 527 1383 531
rect 1423 531 1427 535
rect 1479 531 1483 535
rect 1527 531 1531 535
rect 1575 531 1579 535
rect 1623 531 1627 535
rect 1655 531 1659 535
rect 1695 529 1699 533
rect 1191 523 1195 527
rect 1435 523 1439 527
rect 111 512 115 516
rect 135 514 139 518
rect 275 515 276 519
rect 276 515 279 519
rect 499 515 500 519
rect 500 515 503 519
rect 507 513 511 517
rect 747 515 751 519
rect 835 515 839 519
rect 1055 515 1056 519
rect 1056 515 1059 519
rect 1155 515 1159 519
rect 1259 513 1263 517
rect 1423 514 1427 518
rect 151 507 152 511
rect 152 507 155 511
rect 295 503 299 507
rect 175 494 179 498
rect 247 489 251 493
rect 303 493 307 497
rect 399 494 403 498
rect 611 499 615 503
rect 767 503 771 507
rect 655 494 659 498
rect 783 494 787 498
rect 935 494 939 498
rect 187 483 188 487
rect 188 483 191 487
rect 235 479 239 483
rect 323 483 324 487
rect 324 483 327 487
rect 379 483 380 487
rect 380 483 383 487
rect 391 483 392 487
rect 392 483 395 487
rect 407 488 411 491
rect 471 489 475 493
rect 407 487 408 488
rect 408 487 411 488
rect 275 471 279 475
rect 315 475 319 479
rect 383 475 387 479
rect 459 479 463 483
rect 479 483 483 487
rect 627 487 631 491
rect 727 489 731 493
rect 871 489 875 493
rect 1031 489 1035 493
rect 1143 499 1147 503
rect 1223 503 1227 507
rect 1479 514 1483 518
rect 1527 514 1531 518
rect 1607 523 1611 527
rect 1575 514 1579 518
rect 1623 514 1627 518
rect 1655 514 1659 518
rect 1583 507 1587 511
rect 1695 512 1699 516
rect 1671 507 1672 511
rect 1672 507 1675 511
rect 1103 494 1107 498
rect 1199 489 1203 493
rect 567 479 571 483
rect 643 483 647 487
rect 667 483 668 487
rect 668 483 671 487
rect 499 471 503 475
rect 715 479 719 483
rect 735 483 739 487
rect 795 483 796 487
rect 796 483 799 487
rect 807 483 808 487
rect 808 483 811 487
rect 835 483 839 487
rect 843 479 847 483
rect 943 483 944 487
rect 944 483 947 487
rect 959 483 960 487
rect 960 483 963 487
rect 747 471 751 475
rect 1003 479 1007 483
rect 951 471 955 475
rect 1055 475 1059 479
rect 1111 483 1112 487
rect 1112 483 1115 487
rect 1155 483 1159 487
rect 1191 479 1195 483
rect 1223 483 1224 487
rect 1224 483 1227 487
rect 1215 475 1219 479
rect 1347 471 1351 475
rect 275 463 279 467
rect 611 463 615 467
rect 667 463 671 467
rect 795 463 799 467
rect 1231 463 1235 467
rect 187 455 191 459
rect 407 455 411 459
rect 535 455 539 459
rect 1043 455 1047 459
rect 323 447 327 451
rect 607 447 611 451
rect 687 447 691 451
rect 1087 447 1091 451
rect 551 439 555 443
rect 943 439 947 443
rect 959 439 963 443
rect 679 431 683 435
rect 923 431 927 435
rect 1331 431 1335 435
rect 311 419 315 423
rect 551 419 555 423
rect 807 423 811 427
rect 1191 419 1195 423
rect 1267 419 1271 423
rect 1339 419 1343 423
rect 295 399 296 403
rect 296 399 299 403
rect 311 399 312 403
rect 312 399 315 403
rect 391 411 395 415
rect 355 403 359 407
rect 383 403 387 407
rect 375 395 379 399
rect 479 403 483 407
rect 643 411 647 415
rect 527 399 531 403
rect 551 399 552 403
rect 552 399 555 403
rect 595 403 599 407
rect 615 395 619 399
rect 627 399 631 403
rect 735 407 739 411
rect 747 411 751 415
rect 687 399 688 403
rect 688 399 691 403
rect 719 399 723 403
rect 767 403 771 407
rect 883 407 887 411
rect 1163 411 1167 415
rect 1175 411 1179 415
rect 1367 411 1371 415
rect 959 399 960 403
rect 960 399 963 403
rect 1055 399 1059 403
rect 1063 399 1067 403
rect 1127 395 1131 399
rect 1379 403 1383 407
rect 303 390 307 394
rect 535 387 539 391
rect 543 390 547 394
rect 671 391 675 395
rect 951 390 955 394
rect 1231 391 1235 395
rect 111 372 115 376
rect 135 370 139 374
rect 167 370 171 374
rect 111 355 115 359
rect 199 370 203 374
rect 231 370 235 374
rect 263 370 267 374
rect 248 359 252 363
rect 355 363 359 367
rect 391 367 395 371
rect 415 370 419 374
rect 447 370 451 374
rect 431 359 432 363
rect 432 359 435 363
rect 487 373 491 377
rect 519 375 520 379
rect 520 375 523 379
rect 883 379 884 383
rect 884 379 887 383
rect 1191 383 1195 387
rect 1215 383 1219 387
rect 1367 395 1368 399
rect 1368 395 1371 399
rect 1455 395 1459 399
rect 1359 385 1363 389
rect 923 375 924 379
rect 924 375 927 379
rect 527 367 531 371
rect 595 363 599 367
rect 643 367 644 371
rect 644 367 647 371
rect 755 371 759 375
rect 903 370 907 374
rect 1031 373 1035 377
rect 1063 375 1064 379
rect 1064 375 1067 379
rect 1339 375 1340 379
rect 1340 375 1343 379
rect 1075 371 1079 375
rect 1439 375 1443 379
rect 1495 375 1496 379
rect 1496 375 1499 379
rect 1607 375 1608 379
rect 1608 375 1611 379
rect 1319 370 1323 374
rect 135 353 139 357
rect 167 353 171 357
rect 199 353 203 357
rect 155 347 159 351
rect 231 353 235 357
rect 263 353 267 357
rect 295 352 299 356
rect 415 353 419 357
rect 447 353 451 357
rect 535 352 539 356
rect 783 356 787 360
rect 879 355 880 359
rect 880 355 883 359
rect 919 359 920 363
rect 920 359 923 363
rect 1003 363 1007 367
rect 1331 367 1335 371
rect 1479 370 1483 374
rect 1519 370 1523 374
rect 1559 370 1563 374
rect 1591 370 1595 374
rect 375 348 379 352
rect 503 346 507 350
rect 615 348 619 352
rect 671 350 675 354
rect 903 353 907 357
rect 943 352 947 356
rect 1103 356 1107 360
rect 1195 355 1199 359
rect 1335 359 1336 363
rect 1336 359 1339 363
rect 1047 346 1051 350
rect 1231 350 1235 354
rect 1319 353 1323 357
rect 1439 352 1443 356
rect 1455 355 1456 359
rect 1456 355 1459 359
rect 1576 359 1580 363
rect 1623 370 1627 374
rect 1655 370 1659 374
rect 1695 372 1699 376
rect 1479 353 1483 357
rect 1519 353 1523 357
rect 1559 353 1563 357
rect 1591 353 1595 357
rect 1623 353 1627 357
rect 1655 353 1659 357
rect 1351 345 1355 349
rect 1643 347 1647 351
rect 1695 355 1699 359
rect 567 335 571 339
rect 1039 339 1043 343
rect 519 327 523 331
rect 711 327 715 331
rect 983 319 987 323
rect 1175 315 1179 319
rect 1215 315 1219 319
rect 1199 307 1203 311
rect 111 297 115 301
rect 135 299 139 303
rect 167 299 171 303
rect 199 299 203 303
rect 231 299 235 303
rect 263 299 267 303
rect 295 299 299 303
rect 327 299 331 303
rect 359 299 363 303
rect 391 299 395 303
rect 423 299 427 303
rect 455 299 459 303
rect 487 299 491 303
rect 519 299 523 303
rect 551 299 555 303
rect 599 302 603 306
rect 703 302 707 306
rect 807 302 811 306
rect 911 302 915 306
rect 1495 307 1499 311
rect 999 299 1003 303
rect 1031 299 1035 303
rect 1063 299 1067 303
rect 1111 302 1115 306
rect 1287 300 1291 304
rect 83 279 84 283
rect 84 279 87 283
rect 111 280 115 284
rect 135 282 139 286
rect 167 282 171 286
rect 155 275 156 279
rect 156 275 159 279
rect 199 282 203 286
rect 231 282 235 286
rect 275 291 279 295
rect 263 282 267 286
rect 295 282 299 286
rect 327 282 331 286
rect 359 282 363 286
rect 391 282 395 286
rect 423 282 427 286
rect 455 282 459 286
rect 367 275 371 279
rect 431 275 435 279
rect 487 282 491 286
rect 531 291 535 295
rect 567 291 568 295
rect 568 291 571 295
rect 779 291 783 295
rect 919 291 923 295
rect 1043 291 1047 295
rect 1299 295 1303 299
rect 1319 299 1323 303
rect 1351 299 1355 303
rect 1383 299 1387 303
rect 1415 299 1419 303
rect 1447 299 1451 303
rect 1479 299 1483 303
rect 1519 299 1523 303
rect 1559 299 1563 303
rect 1591 299 1595 303
rect 1623 299 1627 303
rect 1655 299 1659 303
rect 1695 297 1699 301
rect 519 282 523 286
rect 551 282 555 286
rect 999 282 1003 286
rect 583 275 587 279
rect 623 271 627 275
rect 831 271 835 275
rect 983 271 987 275
rect 1007 271 1011 275
rect 1031 282 1035 286
rect 1063 282 1067 286
rect 1319 282 1323 286
rect 1351 282 1355 286
rect 1287 277 1291 281
rect 1335 275 1336 279
rect 1336 275 1339 279
rect 1383 282 1387 286
rect 1415 282 1419 286
rect 1447 282 1451 286
rect 1479 282 1483 286
rect 1531 291 1535 295
rect 1519 282 1523 286
rect 1559 282 1563 286
rect 1591 282 1595 286
rect 1623 282 1627 286
rect 1655 282 1659 286
rect 1607 275 1608 279
rect 1608 275 1611 279
rect 1643 275 1644 279
rect 1644 275 1647 279
rect 1671 291 1672 295
rect 1672 291 1675 295
rect 1723 287 1727 291
rect 1695 280 1699 284
rect 1083 267 1087 271
rect 599 261 603 265
rect 703 261 707 265
rect 807 261 811 265
rect 911 261 915 265
rect 1111 261 1115 265
rect 607 251 611 255
rect 711 251 715 255
rect 779 251 780 255
rect 780 251 783 255
rect 623 243 627 247
rect 671 243 675 247
rect 823 251 824 255
rect 824 251 827 255
rect 879 251 880 255
rect 880 251 883 255
rect 927 251 928 255
rect 928 251 931 255
rect 983 251 984 255
rect 984 251 987 255
rect 1007 247 1011 251
rect 1119 247 1123 251
rect 1127 251 1128 255
rect 1128 251 1131 255
rect 1183 255 1187 259
rect 1207 267 1211 271
rect 1215 255 1216 259
rect 1216 255 1219 259
rect 1299 255 1303 259
rect 111 212 115 216
rect 271 223 275 227
rect 331 223 335 227
rect 583 227 587 231
rect 655 227 659 231
rect 695 231 699 235
rect 807 235 811 239
rect 831 235 832 239
rect 832 235 835 239
rect 851 235 852 239
rect 852 235 855 239
rect 935 235 939 239
rect 967 231 971 235
rect 839 225 843 229
rect 1199 227 1203 231
rect 183 210 187 214
rect 215 210 219 214
rect 247 210 251 214
rect 279 210 283 214
rect 311 210 315 214
rect 359 215 360 219
rect 360 215 363 219
rect 343 210 347 214
rect 367 207 371 211
rect 375 210 379 214
rect 407 210 411 214
rect 439 210 443 214
rect 471 210 475 214
rect 520 215 524 219
rect 503 210 507 214
rect 535 210 539 214
rect 567 210 571 214
rect 111 195 115 199
rect 331 199 332 203
rect 332 199 335 203
rect 487 200 488 203
rect 488 200 491 203
rect 487 199 491 200
rect 647 215 651 219
rect 719 219 723 223
rect 599 210 603 214
rect 639 210 643 214
rect 791 210 795 214
rect 919 215 923 219
rect 983 219 987 223
rect 1075 215 1079 219
rect 1063 210 1067 214
rect 1103 210 1107 214
rect 1143 210 1147 214
rect 1183 210 1187 214
rect 1223 210 1227 214
rect 615 199 616 203
rect 616 199 619 203
rect 655 199 656 203
rect 656 199 659 203
rect 807 199 808 203
rect 808 199 811 203
rect 183 193 187 197
rect 215 193 219 197
rect 247 193 251 197
rect 279 193 283 197
rect 311 193 315 197
rect 343 193 347 197
rect 375 193 379 197
rect 407 193 411 197
rect 439 193 443 197
rect 471 193 475 197
rect 503 193 507 197
rect 535 193 539 197
rect 567 193 571 197
rect 599 193 603 197
rect 639 193 643 197
rect 359 187 363 191
rect 487 187 491 191
rect 695 190 699 194
rect 791 193 795 197
rect 919 192 923 196
rect 935 195 936 199
rect 936 195 939 199
rect 1083 199 1084 203
rect 1084 199 1087 203
rect 1163 199 1164 203
rect 1164 199 1167 203
rect 1199 199 1200 203
rect 1200 199 1203 203
rect 1311 219 1315 223
rect 1531 227 1535 231
rect 1263 210 1267 214
rect 1303 210 1307 214
rect 1343 210 1347 214
rect 1375 210 1379 214
rect 1407 210 1411 214
rect 1439 210 1443 214
rect 1599 215 1603 219
rect 1479 210 1483 214
rect 1519 210 1523 214
rect 1559 210 1563 214
rect 1591 210 1595 214
rect 1623 210 1627 214
rect 1655 210 1659 214
rect 1579 199 1580 203
rect 1580 199 1583 203
rect 1607 199 1608 203
rect 1608 199 1611 203
rect 1643 199 1644 203
rect 1644 199 1647 203
rect 1671 215 1672 219
rect 1672 215 1675 219
rect 1695 212 1699 216
rect 967 190 971 194
rect 1063 193 1067 197
rect 1103 193 1107 197
rect 1143 193 1147 197
rect 1183 193 1187 197
rect 1223 193 1227 197
rect 1263 193 1267 197
rect 1303 193 1307 197
rect 1343 193 1347 197
rect 1375 193 1379 197
rect 1407 193 1411 197
rect 1439 193 1443 197
rect 1479 193 1483 197
rect 1519 193 1523 197
rect 1559 193 1563 197
rect 1591 193 1595 197
rect 1623 193 1627 197
rect 1655 193 1659 197
rect 1695 195 1699 199
rect 831 185 835 189
rect 1119 187 1123 191
rect 111 161 115 165
rect 135 163 139 167
rect 167 163 171 167
rect 215 163 219 167
rect 263 163 267 167
rect 311 163 315 167
rect 367 163 371 167
rect 415 163 419 167
rect 471 163 475 167
rect 535 163 539 167
rect 607 163 611 167
rect 687 163 691 167
rect 775 163 779 167
rect 863 163 867 167
rect 959 163 963 167
rect 1055 163 1059 167
rect 1151 163 1155 167
rect 1239 163 1243 167
rect 1327 163 1331 167
rect 1415 163 1419 167
rect 1503 163 1507 167
rect 1591 163 1595 167
rect 1655 163 1659 167
rect 1695 161 1699 165
rect 151 155 152 159
rect 152 155 155 159
rect 111 144 115 148
rect 135 146 139 150
rect 167 146 171 150
rect 215 146 219 150
rect 263 146 267 150
rect 311 146 315 150
rect 367 146 371 150
rect 415 146 419 150
rect 471 146 475 150
rect 647 155 651 159
rect 535 146 539 150
rect 607 146 611 150
rect 615 139 619 143
rect 687 146 691 150
rect 775 146 779 150
rect 999 155 1003 159
rect 1075 155 1076 159
rect 1076 155 1079 159
rect 863 146 867 150
rect 959 146 963 150
rect 1055 146 1059 150
rect 919 139 923 143
rect 1151 146 1155 150
rect 1239 146 1243 150
rect 1163 139 1167 143
rect 1195 139 1199 143
rect 1311 155 1315 159
rect 1327 146 1331 150
rect 1415 146 1419 150
rect 1535 155 1539 159
rect 1543 155 1547 159
rect 1671 155 1672 159
rect 1672 155 1675 159
rect 1503 146 1507 150
rect 1591 146 1595 150
rect 1655 146 1659 150
rect 1695 144 1699 148
rect 1579 139 1583 143
rect 1643 139 1647 143
rect 1027 131 1031 135
rect 1543 131 1547 135
rect 111 104 115 108
rect 151 107 152 111
rect 152 107 155 111
rect 135 102 139 106
rect 111 87 115 91
rect 167 102 171 106
rect 199 102 203 106
rect 231 102 235 106
rect 263 102 267 106
rect 295 102 299 106
rect 327 102 331 106
rect 359 102 363 106
rect 391 102 395 106
rect 423 102 427 106
rect 455 102 459 106
rect 487 102 491 106
rect 519 102 523 106
rect 999 107 1000 111
rect 1000 107 1003 111
rect 1071 107 1072 111
rect 1072 107 1075 111
rect 551 102 555 106
rect 607 102 611 106
rect 671 102 675 106
rect 743 102 747 106
rect 823 102 827 106
rect 903 102 907 106
rect 983 102 987 106
rect 1055 102 1059 106
rect 1119 102 1123 106
rect 1175 102 1179 106
rect 1223 102 1227 106
rect 1271 102 1275 106
rect 919 91 920 95
rect 920 91 923 95
rect 1027 91 1031 95
rect 1195 91 1196 95
rect 1196 91 1199 95
rect 135 85 139 89
rect 167 85 171 89
rect 199 85 203 89
rect 231 85 235 89
rect 263 85 267 89
rect 295 85 299 89
rect 327 85 331 89
rect 359 85 363 89
rect 391 85 395 89
rect 423 85 427 89
rect 455 85 459 89
rect 487 85 491 89
rect 519 85 523 89
rect 551 85 555 89
rect 607 85 611 89
rect 623 83 627 87
rect 671 85 675 89
rect 743 85 747 89
rect 823 85 827 89
rect 903 85 907 89
rect 983 85 987 89
rect 1055 85 1059 89
rect 1119 85 1123 89
rect 1175 85 1179 89
rect 1223 85 1227 89
rect 1071 79 1075 83
rect 1311 102 1315 106
rect 1343 102 1347 106
rect 1375 102 1379 106
rect 1407 102 1411 106
rect 1439 102 1443 106
rect 1479 102 1483 106
rect 1519 102 1523 106
rect 1535 107 1536 111
rect 1536 107 1539 111
rect 1559 102 1563 106
rect 1591 102 1595 106
rect 1623 102 1627 106
rect 1603 91 1607 95
rect 1655 102 1659 106
rect 1671 107 1672 111
rect 1672 107 1675 111
rect 1695 104 1699 108
rect 1271 85 1275 89
rect 1311 85 1315 89
rect 1343 85 1347 89
rect 1375 85 1379 89
rect 1407 85 1411 89
rect 1439 85 1443 89
rect 1479 85 1483 89
rect 1519 85 1523 89
rect 1559 85 1563 89
rect 1591 85 1595 89
rect 1623 85 1627 89
rect 1655 85 1659 89
rect 1695 87 1699 91
<< m3 >>
rect 870 1763 876 1764
rect 111 1762 115 1763
rect 111 1757 115 1758
rect 151 1762 155 1763
rect 112 1754 114 1757
rect 151 1756 155 1758
rect 183 1762 187 1763
rect 183 1756 187 1758
rect 215 1762 219 1763
rect 215 1756 219 1758
rect 247 1762 251 1763
rect 247 1756 251 1758
rect 279 1762 283 1763
rect 279 1756 283 1758
rect 311 1762 315 1763
rect 311 1756 315 1758
rect 343 1762 347 1763
rect 343 1756 347 1758
rect 375 1762 379 1763
rect 375 1756 379 1758
rect 407 1762 411 1763
rect 407 1756 411 1758
rect 439 1762 443 1763
rect 439 1756 443 1758
rect 471 1762 475 1763
rect 471 1756 475 1758
rect 503 1762 507 1763
rect 503 1756 507 1758
rect 535 1762 539 1763
rect 535 1756 539 1758
rect 567 1762 571 1763
rect 567 1756 571 1758
rect 599 1762 603 1763
rect 599 1756 603 1758
rect 631 1762 635 1763
rect 631 1756 635 1758
rect 663 1762 667 1763
rect 663 1756 667 1758
rect 695 1762 699 1763
rect 695 1756 699 1758
rect 727 1762 731 1763
rect 727 1756 731 1758
rect 759 1762 763 1763
rect 759 1756 763 1758
rect 791 1762 795 1763
rect 791 1756 795 1758
rect 823 1762 827 1763
rect 823 1756 827 1758
rect 855 1762 859 1763
rect 870 1759 871 1763
rect 875 1759 876 1763
rect 870 1758 876 1759
rect 887 1762 891 1763
rect 855 1756 859 1758
rect 150 1755 156 1756
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 150 1751 151 1755
rect 155 1751 156 1755
rect 150 1750 156 1751
rect 182 1755 188 1756
rect 182 1751 183 1755
rect 187 1751 188 1755
rect 182 1750 188 1751
rect 214 1755 220 1756
rect 214 1751 215 1755
rect 219 1751 220 1755
rect 214 1750 220 1751
rect 246 1755 252 1756
rect 246 1751 247 1755
rect 251 1751 252 1755
rect 246 1750 252 1751
rect 278 1755 284 1756
rect 278 1751 279 1755
rect 283 1751 284 1755
rect 278 1750 284 1751
rect 310 1755 316 1756
rect 310 1751 311 1755
rect 315 1751 316 1755
rect 310 1750 316 1751
rect 342 1755 348 1756
rect 342 1751 343 1755
rect 347 1751 348 1755
rect 342 1750 348 1751
rect 374 1755 380 1756
rect 374 1751 375 1755
rect 379 1751 380 1755
rect 374 1750 380 1751
rect 406 1755 412 1756
rect 406 1751 407 1755
rect 411 1751 412 1755
rect 406 1750 412 1751
rect 438 1755 444 1756
rect 438 1751 439 1755
rect 443 1751 444 1755
rect 438 1750 444 1751
rect 470 1755 476 1756
rect 470 1751 471 1755
rect 475 1751 476 1755
rect 470 1750 476 1751
rect 502 1755 508 1756
rect 502 1751 503 1755
rect 507 1751 508 1755
rect 502 1750 508 1751
rect 534 1755 540 1756
rect 534 1751 535 1755
rect 539 1751 540 1755
rect 534 1750 540 1751
rect 566 1755 572 1756
rect 566 1751 567 1755
rect 571 1751 572 1755
rect 566 1750 572 1751
rect 598 1755 604 1756
rect 598 1751 599 1755
rect 603 1751 604 1755
rect 598 1750 604 1751
rect 630 1755 636 1756
rect 630 1751 631 1755
rect 635 1751 636 1755
rect 630 1750 636 1751
rect 662 1755 668 1756
rect 662 1751 663 1755
rect 667 1751 668 1755
rect 662 1750 668 1751
rect 694 1755 700 1756
rect 694 1751 695 1755
rect 699 1751 700 1755
rect 694 1750 700 1751
rect 726 1755 732 1756
rect 726 1751 727 1755
rect 731 1751 732 1755
rect 726 1750 732 1751
rect 758 1755 764 1756
rect 758 1751 759 1755
rect 763 1751 764 1755
rect 758 1750 764 1751
rect 790 1755 796 1756
rect 790 1751 791 1755
rect 795 1751 796 1755
rect 790 1750 796 1751
rect 822 1755 828 1756
rect 822 1751 823 1755
rect 827 1751 828 1755
rect 822 1750 828 1751
rect 854 1755 860 1756
rect 854 1751 855 1755
rect 859 1751 860 1755
rect 854 1750 860 1751
rect 110 1748 116 1749
rect 150 1738 156 1739
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 150 1734 151 1738
rect 155 1734 156 1738
rect 150 1733 156 1734
rect 182 1738 188 1739
rect 182 1734 183 1738
rect 187 1734 188 1738
rect 182 1733 188 1734
rect 214 1738 220 1739
rect 214 1734 215 1738
rect 219 1734 220 1738
rect 214 1733 220 1734
rect 246 1738 252 1739
rect 246 1734 247 1738
rect 251 1734 252 1738
rect 246 1733 252 1734
rect 278 1738 284 1739
rect 278 1734 279 1738
rect 283 1734 284 1738
rect 278 1733 284 1734
rect 310 1738 316 1739
rect 310 1734 311 1738
rect 315 1734 316 1738
rect 310 1733 316 1734
rect 342 1738 348 1739
rect 342 1734 343 1738
rect 347 1734 348 1738
rect 342 1733 348 1734
rect 374 1738 380 1739
rect 374 1734 375 1738
rect 379 1734 380 1738
rect 374 1733 380 1734
rect 406 1738 412 1739
rect 406 1734 407 1738
rect 411 1734 412 1738
rect 406 1733 412 1734
rect 438 1738 444 1739
rect 438 1734 439 1738
rect 443 1734 444 1738
rect 438 1733 444 1734
rect 470 1738 476 1739
rect 470 1734 471 1738
rect 475 1734 476 1738
rect 470 1733 476 1734
rect 502 1738 508 1739
rect 502 1734 503 1738
rect 507 1734 508 1738
rect 502 1733 508 1734
rect 534 1738 540 1739
rect 534 1734 535 1738
rect 539 1734 540 1738
rect 534 1733 540 1734
rect 566 1738 572 1739
rect 566 1734 567 1738
rect 571 1734 572 1738
rect 566 1733 572 1734
rect 598 1738 604 1739
rect 598 1734 599 1738
rect 603 1734 604 1738
rect 598 1733 604 1734
rect 630 1738 636 1739
rect 630 1734 631 1738
rect 635 1734 636 1738
rect 630 1733 636 1734
rect 662 1738 668 1739
rect 662 1734 663 1738
rect 667 1734 668 1738
rect 662 1733 668 1734
rect 694 1738 700 1739
rect 694 1734 695 1738
rect 699 1734 700 1738
rect 694 1733 700 1734
rect 726 1738 732 1739
rect 726 1734 727 1738
rect 731 1734 732 1738
rect 726 1733 732 1734
rect 758 1738 764 1739
rect 758 1734 759 1738
rect 763 1734 764 1738
rect 758 1733 764 1734
rect 790 1738 796 1739
rect 790 1734 791 1738
rect 795 1734 796 1738
rect 790 1733 796 1734
rect 822 1738 828 1739
rect 822 1734 823 1738
rect 827 1734 828 1738
rect 822 1733 828 1734
rect 854 1738 860 1739
rect 854 1734 855 1738
rect 859 1734 860 1738
rect 854 1733 860 1734
rect 110 1731 116 1732
rect 112 1719 114 1731
rect 152 1719 154 1733
rect 184 1719 186 1733
rect 216 1719 218 1733
rect 248 1719 250 1733
rect 280 1719 282 1733
rect 312 1719 314 1733
rect 344 1719 346 1733
rect 376 1719 378 1733
rect 408 1719 410 1733
rect 440 1719 442 1733
rect 472 1719 474 1733
rect 504 1719 506 1733
rect 536 1719 538 1733
rect 568 1719 570 1733
rect 600 1719 602 1733
rect 632 1719 634 1733
rect 664 1719 666 1733
rect 696 1719 698 1733
rect 728 1719 730 1733
rect 760 1719 762 1733
rect 792 1719 794 1733
rect 824 1719 826 1733
rect 856 1719 858 1733
rect 111 1718 115 1719
rect 111 1713 115 1714
rect 151 1718 155 1719
rect 151 1713 155 1714
rect 183 1718 187 1719
rect 183 1713 187 1714
rect 191 1718 195 1719
rect 191 1713 195 1714
rect 215 1718 219 1719
rect 215 1713 219 1714
rect 247 1718 251 1719
rect 247 1713 251 1714
rect 279 1718 283 1719
rect 279 1713 283 1714
rect 311 1718 315 1719
rect 311 1713 315 1714
rect 319 1718 323 1719
rect 319 1713 323 1714
rect 343 1718 347 1719
rect 343 1713 347 1714
rect 375 1718 379 1719
rect 375 1713 379 1714
rect 407 1718 411 1719
rect 407 1713 411 1714
rect 415 1718 419 1719
rect 415 1713 419 1714
rect 439 1718 443 1719
rect 439 1713 443 1714
rect 471 1718 475 1719
rect 471 1713 475 1714
rect 503 1718 507 1719
rect 503 1713 507 1714
rect 527 1718 531 1719
rect 527 1713 531 1714
rect 535 1718 539 1719
rect 535 1713 539 1714
rect 567 1718 571 1719
rect 567 1713 571 1714
rect 599 1718 603 1719
rect 599 1713 603 1714
rect 631 1718 635 1719
rect 631 1713 635 1714
rect 655 1718 659 1719
rect 655 1713 659 1714
rect 663 1718 667 1719
rect 663 1713 667 1714
rect 695 1718 699 1719
rect 695 1713 699 1714
rect 727 1718 731 1719
rect 727 1713 731 1714
rect 759 1718 763 1719
rect 759 1713 763 1714
rect 791 1718 795 1719
rect 791 1713 795 1714
rect 823 1718 827 1719
rect 823 1713 827 1714
rect 855 1718 859 1719
rect 855 1713 859 1714
rect 112 1705 114 1713
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 192 1703 194 1713
rect 206 1707 212 1708
rect 206 1703 207 1707
rect 211 1703 212 1707
rect 248 1703 250 1713
rect 320 1703 322 1713
rect 416 1703 418 1713
rect 528 1703 530 1713
rect 656 1703 658 1713
rect 792 1703 794 1713
rect 110 1699 116 1700
rect 190 1702 196 1703
rect 206 1702 212 1703
rect 246 1702 252 1703
rect 190 1698 191 1702
rect 195 1698 196 1702
rect 190 1697 196 1698
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 110 1682 116 1683
rect 190 1685 196 1686
rect 112 1671 114 1682
rect 190 1681 191 1685
rect 195 1681 196 1685
rect 190 1680 196 1681
rect 208 1680 210 1702
rect 246 1698 247 1702
rect 251 1698 252 1702
rect 246 1697 252 1698
rect 318 1702 324 1703
rect 318 1698 319 1702
rect 323 1698 324 1702
rect 318 1697 324 1698
rect 414 1702 420 1703
rect 414 1698 415 1702
rect 419 1698 420 1702
rect 414 1697 420 1698
rect 526 1702 532 1703
rect 526 1698 527 1702
rect 531 1698 532 1702
rect 526 1697 532 1698
rect 654 1702 660 1703
rect 654 1698 655 1702
rect 659 1698 660 1702
rect 654 1697 660 1698
rect 790 1702 796 1703
rect 790 1698 791 1702
rect 795 1698 796 1702
rect 790 1697 796 1698
rect 406 1691 412 1692
rect 406 1687 407 1691
rect 411 1687 412 1691
rect 406 1686 412 1687
rect 246 1685 252 1686
rect 246 1681 247 1685
rect 251 1681 252 1685
rect 246 1680 252 1681
rect 318 1685 324 1686
rect 318 1681 319 1685
rect 323 1681 324 1685
rect 318 1680 324 1681
rect 154 1671 160 1672
rect 192 1671 194 1680
rect 206 1679 212 1680
rect 206 1675 207 1679
rect 211 1675 212 1679
rect 206 1674 212 1675
rect 248 1671 250 1680
rect 320 1671 322 1680
rect 111 1670 115 1671
rect 111 1665 115 1666
rect 135 1670 139 1671
rect 154 1667 155 1671
rect 159 1667 160 1671
rect 154 1666 160 1667
rect 175 1670 179 1671
rect 112 1662 114 1665
rect 135 1664 139 1666
rect 134 1663 140 1664
rect 110 1661 116 1662
rect 110 1657 111 1661
rect 115 1657 116 1661
rect 134 1659 135 1663
rect 139 1659 140 1663
rect 134 1658 140 1659
rect 110 1656 116 1657
rect 134 1646 140 1647
rect 110 1644 116 1645
rect 110 1640 111 1644
rect 115 1640 116 1644
rect 134 1642 135 1646
rect 139 1642 140 1646
rect 134 1641 140 1642
rect 110 1639 116 1640
rect 112 1623 114 1639
rect 136 1623 138 1641
rect 156 1640 158 1666
rect 175 1664 179 1666
rect 191 1670 195 1671
rect 191 1665 195 1666
rect 247 1670 251 1671
rect 247 1665 251 1666
rect 263 1670 267 1671
rect 263 1664 267 1666
rect 319 1670 323 1671
rect 319 1665 323 1666
rect 391 1670 395 1671
rect 391 1664 395 1666
rect 174 1663 180 1664
rect 174 1659 175 1663
rect 179 1659 180 1663
rect 174 1658 180 1659
rect 262 1663 268 1664
rect 262 1659 263 1663
rect 267 1659 268 1663
rect 262 1658 268 1659
rect 390 1663 396 1664
rect 390 1659 391 1663
rect 395 1659 396 1663
rect 390 1658 396 1659
rect 342 1655 348 1656
rect 342 1651 343 1655
rect 347 1651 348 1655
rect 342 1650 348 1651
rect 174 1646 180 1647
rect 174 1642 175 1646
rect 179 1642 180 1646
rect 174 1641 180 1642
rect 262 1646 268 1647
rect 262 1642 263 1646
rect 267 1642 268 1646
rect 262 1641 268 1642
rect 154 1639 160 1640
rect 154 1635 155 1639
rect 159 1635 160 1639
rect 154 1634 160 1635
rect 176 1623 178 1641
rect 186 1631 192 1632
rect 186 1627 187 1631
rect 191 1627 192 1631
rect 186 1626 192 1627
rect 111 1622 115 1623
rect 111 1617 115 1618
rect 135 1622 139 1623
rect 135 1617 139 1618
rect 167 1622 171 1623
rect 167 1617 171 1618
rect 175 1622 179 1623
rect 175 1617 179 1618
rect 112 1609 114 1617
rect 110 1608 116 1609
rect 110 1604 111 1608
rect 115 1604 116 1608
rect 136 1607 138 1617
rect 168 1607 170 1617
rect 110 1603 116 1604
rect 134 1606 140 1607
rect 134 1602 135 1606
rect 139 1602 140 1606
rect 134 1601 140 1602
rect 166 1606 172 1607
rect 166 1602 167 1606
rect 171 1602 172 1606
rect 166 1601 172 1602
rect 150 1595 156 1596
rect 110 1591 116 1592
rect 110 1587 111 1591
rect 115 1587 116 1591
rect 150 1591 151 1595
rect 155 1591 156 1595
rect 150 1590 156 1591
rect 110 1586 116 1587
rect 134 1589 140 1590
rect 112 1583 114 1586
rect 134 1585 135 1589
rect 139 1585 140 1589
rect 134 1584 140 1585
rect 111 1582 115 1583
rect 111 1577 115 1578
rect 135 1582 139 1584
rect 112 1574 114 1577
rect 135 1576 139 1578
rect 134 1575 140 1576
rect 110 1573 116 1574
rect 110 1569 111 1573
rect 115 1569 116 1573
rect 134 1571 135 1575
rect 139 1571 140 1575
rect 134 1570 140 1571
rect 110 1568 116 1569
rect 134 1558 140 1559
rect 110 1556 116 1557
rect 110 1552 111 1556
rect 115 1552 116 1556
rect 134 1554 135 1558
rect 139 1554 140 1558
rect 134 1553 140 1554
rect 110 1551 116 1552
rect 112 1543 114 1551
rect 136 1543 138 1553
rect 152 1552 154 1590
rect 166 1589 172 1590
rect 166 1585 167 1589
rect 171 1585 172 1589
rect 166 1584 172 1585
rect 167 1582 171 1584
rect 167 1576 171 1578
rect 166 1575 172 1576
rect 166 1571 167 1575
rect 171 1571 172 1575
rect 166 1570 172 1571
rect 166 1558 172 1559
rect 166 1554 167 1558
rect 171 1554 172 1558
rect 166 1553 172 1554
rect 150 1551 156 1552
rect 150 1547 151 1551
rect 155 1547 156 1551
rect 150 1546 156 1547
rect 168 1543 170 1553
rect 111 1542 115 1543
rect 111 1537 115 1538
rect 135 1542 139 1543
rect 135 1537 139 1538
rect 167 1542 171 1543
rect 167 1537 171 1538
rect 175 1542 179 1543
rect 175 1537 179 1538
rect 112 1529 114 1537
rect 110 1528 116 1529
rect 110 1524 111 1528
rect 115 1524 116 1528
rect 136 1527 138 1537
rect 176 1527 178 1537
rect 110 1523 116 1524
rect 134 1526 140 1527
rect 134 1522 135 1526
rect 139 1522 140 1526
rect 134 1521 140 1522
rect 174 1526 180 1527
rect 174 1522 175 1526
rect 179 1522 180 1526
rect 174 1521 180 1522
rect 110 1511 116 1512
rect 102 1507 108 1508
rect 102 1503 103 1507
rect 107 1503 108 1507
rect 110 1507 111 1511
rect 115 1507 116 1511
rect 110 1506 116 1507
rect 134 1509 140 1510
rect 102 1502 108 1503
rect 104 1272 106 1502
rect 112 1499 114 1506
rect 134 1505 135 1509
rect 139 1505 140 1509
rect 134 1504 140 1505
rect 174 1509 180 1510
rect 174 1505 175 1509
rect 179 1505 180 1509
rect 174 1504 180 1505
rect 136 1499 138 1504
rect 176 1499 178 1504
rect 111 1498 115 1499
rect 111 1493 115 1494
rect 135 1498 139 1499
rect 135 1493 139 1494
rect 175 1498 179 1499
rect 175 1493 179 1494
rect 112 1474 114 1493
rect 176 1476 178 1493
rect 174 1475 180 1476
rect 110 1473 116 1474
rect 110 1469 111 1473
rect 115 1469 116 1473
rect 174 1471 175 1475
rect 179 1471 180 1475
rect 174 1470 180 1471
rect 110 1468 116 1469
rect 150 1467 156 1468
rect 150 1463 151 1467
rect 155 1463 156 1467
rect 150 1462 156 1463
rect 110 1456 116 1457
rect 110 1452 111 1456
rect 115 1452 116 1456
rect 110 1451 116 1452
rect 112 1431 114 1451
rect 111 1430 115 1431
rect 111 1425 115 1426
rect 135 1430 139 1431
rect 135 1425 139 1426
rect 112 1393 114 1425
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 136 1391 138 1425
rect 152 1396 154 1462
rect 174 1458 180 1459
rect 174 1454 175 1458
rect 179 1454 180 1458
rect 174 1453 180 1454
rect 176 1431 178 1453
rect 167 1430 171 1431
rect 167 1425 171 1426
rect 175 1430 179 1431
rect 175 1425 179 1426
rect 150 1395 156 1396
rect 150 1391 151 1395
rect 155 1391 156 1395
rect 168 1391 170 1425
rect 110 1387 116 1388
rect 134 1390 140 1391
rect 150 1390 156 1391
rect 166 1390 172 1391
rect 134 1386 135 1390
rect 139 1386 140 1390
rect 134 1385 140 1386
rect 166 1386 167 1390
rect 171 1386 172 1390
rect 166 1385 172 1386
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 110 1370 116 1371
rect 134 1373 140 1374
rect 112 1351 114 1370
rect 134 1369 135 1373
rect 139 1369 140 1373
rect 134 1368 140 1369
rect 166 1373 172 1374
rect 166 1369 167 1373
rect 171 1369 172 1373
rect 166 1368 172 1369
rect 136 1351 138 1368
rect 168 1351 170 1368
rect 111 1350 115 1351
rect 111 1345 115 1346
rect 135 1350 139 1351
rect 135 1345 139 1346
rect 167 1350 171 1351
rect 167 1345 171 1346
rect 112 1318 114 1345
rect 136 1320 138 1345
rect 168 1320 170 1345
rect 178 1335 184 1336
rect 178 1331 179 1335
rect 183 1331 184 1335
rect 178 1330 184 1331
rect 134 1319 140 1320
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1315 135 1319
rect 139 1315 140 1319
rect 134 1314 140 1315
rect 166 1319 172 1320
rect 166 1315 167 1319
rect 171 1315 172 1319
rect 166 1314 172 1315
rect 110 1312 116 1313
rect 150 1311 156 1312
rect 150 1307 151 1311
rect 155 1307 156 1311
rect 150 1306 156 1307
rect 134 1302 140 1303
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 134 1298 135 1302
rect 139 1298 140 1302
rect 134 1297 140 1298
rect 110 1295 116 1296
rect 102 1271 108 1272
rect 102 1267 103 1271
rect 107 1267 108 1271
rect 102 1266 108 1267
rect 112 1263 114 1295
rect 136 1263 138 1297
rect 111 1262 115 1263
rect 111 1257 115 1258
rect 135 1262 139 1263
rect 135 1257 139 1258
rect 112 1197 114 1257
rect 110 1196 116 1197
rect 110 1192 111 1196
rect 115 1192 116 1196
rect 136 1195 138 1257
rect 152 1200 154 1306
rect 166 1302 172 1303
rect 166 1298 167 1302
rect 171 1298 172 1302
rect 166 1297 172 1298
rect 168 1263 170 1297
rect 167 1262 171 1263
rect 167 1257 171 1258
rect 150 1199 156 1200
rect 150 1195 151 1199
rect 155 1195 156 1199
rect 168 1195 170 1257
rect 110 1191 116 1192
rect 134 1194 140 1195
rect 150 1194 156 1195
rect 166 1194 172 1195
rect 134 1190 135 1194
rect 139 1190 140 1194
rect 134 1189 140 1190
rect 166 1190 167 1194
rect 171 1190 172 1194
rect 166 1189 172 1190
rect 110 1179 116 1180
rect 110 1175 111 1179
rect 115 1175 116 1179
rect 110 1174 116 1175
rect 134 1177 140 1178
rect 112 1151 114 1174
rect 134 1173 135 1177
rect 139 1173 140 1177
rect 134 1172 140 1173
rect 166 1177 172 1178
rect 166 1173 167 1177
rect 171 1173 172 1177
rect 166 1172 172 1173
rect 136 1151 138 1172
rect 168 1151 170 1172
rect 111 1150 115 1151
rect 111 1145 115 1146
rect 135 1150 139 1151
rect 135 1145 139 1146
rect 167 1150 171 1151
rect 167 1145 171 1146
rect 112 1122 114 1145
rect 136 1124 138 1145
rect 168 1124 170 1145
rect 134 1123 140 1124
rect 110 1121 116 1122
rect 110 1117 111 1121
rect 115 1117 116 1121
rect 134 1119 135 1123
rect 139 1119 140 1123
rect 134 1118 140 1119
rect 166 1123 172 1124
rect 166 1119 167 1123
rect 171 1119 172 1123
rect 166 1118 172 1119
rect 110 1116 116 1117
rect 134 1106 140 1107
rect 110 1104 116 1105
rect 110 1100 111 1104
rect 115 1100 116 1104
rect 134 1102 135 1106
rect 139 1102 140 1106
rect 134 1101 140 1102
rect 166 1106 172 1107
rect 166 1102 167 1106
rect 171 1102 172 1106
rect 166 1101 172 1102
rect 110 1099 116 1100
rect 112 1035 114 1099
rect 136 1035 138 1101
rect 168 1035 170 1101
rect 180 1045 182 1330
rect 188 1280 190 1626
rect 264 1623 266 1641
rect 199 1622 203 1623
rect 199 1617 203 1618
rect 247 1622 251 1623
rect 247 1617 251 1618
rect 263 1622 267 1623
rect 263 1617 267 1618
rect 327 1622 331 1623
rect 327 1617 331 1618
rect 200 1607 202 1617
rect 248 1607 250 1617
rect 328 1607 330 1617
rect 344 1612 346 1650
rect 390 1646 396 1647
rect 390 1642 391 1646
rect 395 1642 396 1646
rect 390 1641 396 1642
rect 392 1623 394 1641
rect 408 1640 410 1686
rect 414 1685 420 1686
rect 414 1681 415 1685
rect 419 1681 420 1685
rect 414 1680 420 1681
rect 526 1685 532 1686
rect 526 1681 527 1685
rect 531 1681 532 1685
rect 526 1680 532 1681
rect 654 1685 660 1686
rect 654 1681 655 1685
rect 659 1681 660 1685
rect 654 1680 660 1681
rect 790 1685 796 1686
rect 790 1681 791 1685
rect 795 1681 796 1685
rect 790 1680 796 1681
rect 416 1671 418 1680
rect 528 1671 530 1680
rect 656 1671 658 1680
rect 792 1671 794 1680
rect 415 1670 419 1671
rect 415 1665 419 1666
rect 527 1670 531 1671
rect 527 1665 531 1666
rect 543 1670 547 1671
rect 543 1664 547 1666
rect 655 1670 659 1671
rect 655 1665 659 1666
rect 711 1670 715 1671
rect 711 1664 715 1666
rect 791 1670 795 1671
rect 791 1665 795 1666
rect 542 1663 548 1664
rect 542 1659 543 1663
rect 547 1659 548 1663
rect 542 1658 548 1659
rect 710 1663 716 1664
rect 710 1659 711 1663
rect 715 1659 716 1663
rect 710 1658 716 1659
rect 542 1646 548 1647
rect 542 1642 543 1646
rect 547 1642 548 1646
rect 542 1641 548 1642
rect 710 1646 716 1647
rect 710 1642 711 1646
rect 715 1642 716 1646
rect 710 1641 716 1642
rect 406 1639 412 1640
rect 406 1635 407 1639
rect 411 1635 412 1639
rect 406 1634 412 1635
rect 544 1623 546 1641
rect 582 1623 588 1624
rect 712 1623 714 1641
rect 391 1622 395 1623
rect 391 1617 395 1618
rect 439 1622 443 1623
rect 439 1617 443 1618
rect 543 1622 547 1623
rect 543 1617 547 1618
rect 567 1622 571 1623
rect 582 1619 583 1623
rect 587 1619 588 1623
rect 582 1618 588 1619
rect 711 1622 715 1623
rect 567 1617 571 1618
rect 342 1611 348 1612
rect 342 1607 343 1611
rect 347 1607 348 1611
rect 440 1607 442 1617
rect 568 1607 570 1617
rect 198 1606 204 1607
rect 198 1602 199 1606
rect 203 1602 204 1606
rect 198 1601 204 1602
rect 246 1606 252 1607
rect 246 1602 247 1606
rect 251 1602 252 1606
rect 246 1601 252 1602
rect 326 1606 332 1607
rect 342 1606 348 1607
rect 438 1606 444 1607
rect 326 1602 327 1606
rect 331 1602 332 1606
rect 326 1601 332 1602
rect 438 1602 439 1606
rect 443 1602 444 1606
rect 438 1601 444 1602
rect 566 1606 572 1607
rect 566 1602 567 1606
rect 571 1602 572 1606
rect 566 1601 572 1602
rect 584 1596 586 1618
rect 711 1617 715 1618
rect 855 1622 859 1623
rect 855 1617 859 1618
rect 712 1607 714 1617
rect 856 1607 858 1617
rect 872 1611 874 1758
rect 887 1756 891 1758
rect 919 1762 923 1763
rect 919 1756 923 1758
rect 951 1762 955 1763
rect 951 1756 955 1758
rect 983 1762 987 1763
rect 1695 1762 1699 1763
rect 983 1756 987 1758
rect 1190 1759 1196 1760
rect 886 1755 892 1756
rect 886 1751 887 1755
rect 891 1751 892 1755
rect 886 1750 892 1751
rect 918 1755 924 1756
rect 918 1751 919 1755
rect 923 1751 924 1755
rect 918 1750 924 1751
rect 950 1755 956 1756
rect 950 1751 951 1755
rect 955 1751 956 1755
rect 950 1750 956 1751
rect 982 1755 988 1756
rect 982 1751 983 1755
rect 987 1751 988 1755
rect 1190 1755 1191 1759
rect 1195 1755 1196 1759
rect 1695 1757 1699 1758
rect 1190 1754 1196 1755
rect 1696 1754 1698 1757
rect 982 1750 988 1751
rect 886 1738 892 1739
rect 886 1734 887 1738
rect 891 1734 892 1738
rect 886 1733 892 1734
rect 918 1738 924 1739
rect 918 1734 919 1738
rect 923 1734 924 1738
rect 918 1733 924 1734
rect 950 1738 956 1739
rect 950 1734 951 1738
rect 955 1734 956 1738
rect 950 1733 956 1734
rect 982 1738 988 1739
rect 982 1734 983 1738
rect 987 1734 988 1738
rect 982 1733 988 1734
rect 888 1719 890 1733
rect 920 1719 922 1733
rect 952 1719 954 1733
rect 984 1719 986 1733
rect 1062 1731 1068 1732
rect 1062 1727 1063 1731
rect 1067 1727 1068 1731
rect 1062 1726 1068 1727
rect 887 1718 891 1719
rect 887 1713 891 1714
rect 919 1718 923 1719
rect 919 1713 923 1714
rect 951 1718 955 1719
rect 951 1713 955 1714
rect 983 1718 987 1719
rect 983 1713 987 1714
rect 1047 1718 1051 1719
rect 1047 1713 1051 1714
rect 902 1711 908 1712
rect 894 1707 900 1708
rect 894 1703 895 1707
rect 899 1703 900 1707
rect 902 1707 903 1711
rect 907 1707 908 1711
rect 902 1706 908 1707
rect 894 1702 900 1703
rect 879 1670 883 1671
rect 879 1664 883 1666
rect 878 1663 884 1664
rect 878 1659 879 1663
rect 883 1659 884 1663
rect 878 1658 884 1659
rect 896 1656 898 1702
rect 904 1692 906 1706
rect 920 1703 922 1713
rect 1048 1703 1050 1713
rect 918 1702 924 1703
rect 918 1698 919 1702
rect 923 1698 924 1702
rect 918 1697 924 1698
rect 1046 1702 1052 1703
rect 1046 1698 1047 1702
rect 1051 1698 1052 1702
rect 1046 1697 1052 1698
rect 1064 1692 1066 1726
rect 1159 1718 1163 1719
rect 1159 1713 1163 1714
rect 1160 1703 1162 1713
rect 1158 1702 1164 1703
rect 1158 1698 1159 1702
rect 1163 1698 1164 1702
rect 1158 1697 1164 1698
rect 902 1691 908 1692
rect 902 1687 903 1691
rect 907 1687 908 1691
rect 902 1686 908 1687
rect 1062 1691 1068 1692
rect 1062 1687 1063 1691
rect 1067 1687 1068 1691
rect 1062 1686 1068 1687
rect 918 1685 924 1686
rect 918 1681 919 1685
rect 923 1681 924 1685
rect 918 1680 924 1681
rect 1046 1685 1052 1686
rect 1046 1681 1047 1685
rect 1051 1681 1052 1685
rect 1046 1680 1052 1681
rect 1158 1685 1164 1686
rect 1158 1681 1159 1685
rect 1163 1681 1164 1685
rect 1158 1680 1164 1681
rect 920 1671 922 1680
rect 1048 1671 1050 1680
rect 1160 1671 1162 1680
rect 919 1670 923 1671
rect 919 1665 923 1666
rect 1039 1670 1043 1671
rect 1039 1664 1043 1666
rect 1047 1670 1051 1671
rect 1047 1665 1051 1666
rect 1159 1670 1163 1671
rect 1159 1665 1163 1666
rect 1183 1670 1187 1671
rect 1183 1664 1187 1666
rect 1038 1663 1044 1664
rect 1038 1659 1039 1663
rect 1043 1659 1044 1663
rect 1038 1658 1044 1659
rect 1182 1663 1188 1664
rect 1182 1659 1183 1663
rect 1187 1659 1188 1663
rect 1182 1658 1188 1659
rect 894 1655 900 1656
rect 894 1651 895 1655
rect 899 1651 900 1655
rect 894 1650 900 1651
rect 878 1646 884 1647
rect 878 1642 879 1646
rect 883 1642 884 1646
rect 878 1641 884 1642
rect 1038 1646 1044 1647
rect 1038 1642 1039 1646
rect 1043 1642 1044 1646
rect 1038 1641 1044 1642
rect 1182 1646 1188 1647
rect 1182 1642 1183 1646
rect 1187 1642 1188 1646
rect 1182 1641 1188 1642
rect 880 1623 882 1641
rect 1018 1639 1024 1640
rect 1018 1635 1019 1639
rect 1023 1635 1024 1639
rect 1018 1634 1024 1635
rect 879 1622 883 1623
rect 879 1617 883 1618
rect 999 1622 1003 1623
rect 999 1617 1003 1618
rect 974 1611 980 1612
rect 872 1609 882 1611
rect 710 1606 716 1607
rect 710 1602 711 1606
rect 715 1602 716 1606
rect 710 1601 716 1602
rect 854 1606 860 1607
rect 854 1602 855 1606
rect 859 1602 860 1606
rect 854 1601 860 1602
rect 582 1595 588 1596
rect 582 1591 583 1595
rect 587 1591 588 1595
rect 582 1590 588 1591
rect 722 1595 728 1596
rect 722 1591 723 1595
rect 727 1591 728 1595
rect 722 1590 728 1591
rect 198 1589 204 1590
rect 198 1585 199 1589
rect 203 1585 204 1589
rect 198 1584 204 1585
rect 246 1589 252 1590
rect 246 1585 247 1589
rect 251 1585 252 1589
rect 246 1584 252 1585
rect 326 1589 332 1590
rect 326 1585 327 1589
rect 331 1585 332 1589
rect 326 1584 332 1585
rect 438 1589 444 1590
rect 438 1585 439 1589
rect 443 1585 444 1589
rect 438 1584 444 1585
rect 566 1589 572 1590
rect 566 1585 567 1589
rect 571 1585 572 1589
rect 566 1584 572 1585
rect 710 1589 716 1590
rect 710 1585 711 1589
rect 715 1585 716 1589
rect 710 1584 716 1585
rect 199 1582 203 1584
rect 199 1577 203 1578
rect 231 1582 235 1583
rect 231 1576 235 1578
rect 247 1582 251 1584
rect 247 1577 251 1578
rect 287 1582 291 1583
rect 287 1576 291 1578
rect 327 1582 331 1584
rect 327 1577 331 1578
rect 343 1582 347 1583
rect 343 1576 347 1578
rect 399 1582 403 1583
rect 399 1576 403 1578
rect 439 1582 443 1584
rect 439 1577 443 1578
rect 455 1582 459 1583
rect 455 1576 459 1578
rect 511 1582 515 1583
rect 511 1576 515 1578
rect 567 1582 571 1584
rect 567 1577 571 1578
rect 575 1582 579 1583
rect 575 1576 579 1578
rect 655 1582 659 1583
rect 655 1576 659 1578
rect 711 1582 715 1584
rect 711 1577 715 1578
rect 230 1575 236 1576
rect 230 1571 231 1575
rect 235 1571 236 1575
rect 230 1570 236 1571
rect 286 1575 292 1576
rect 286 1571 287 1575
rect 291 1571 292 1575
rect 286 1570 292 1571
rect 342 1575 348 1576
rect 342 1571 343 1575
rect 347 1571 348 1575
rect 342 1570 348 1571
rect 398 1575 404 1576
rect 398 1571 399 1575
rect 403 1571 404 1575
rect 398 1570 404 1571
rect 454 1575 460 1576
rect 454 1571 455 1575
rect 459 1571 460 1575
rect 454 1570 460 1571
rect 510 1575 516 1576
rect 510 1571 511 1575
rect 515 1571 516 1575
rect 510 1570 516 1571
rect 574 1575 580 1576
rect 574 1571 575 1575
rect 579 1571 580 1575
rect 574 1570 580 1571
rect 654 1575 660 1576
rect 654 1571 655 1575
rect 659 1571 660 1575
rect 654 1570 660 1571
rect 298 1567 304 1568
rect 298 1563 299 1567
rect 303 1563 304 1567
rect 298 1562 304 1563
rect 378 1567 384 1568
rect 378 1563 379 1567
rect 383 1563 384 1567
rect 378 1562 384 1563
rect 230 1558 236 1559
rect 230 1554 231 1558
rect 235 1554 236 1558
rect 230 1553 236 1554
rect 286 1558 292 1559
rect 286 1554 287 1558
rect 291 1554 292 1558
rect 286 1553 292 1554
rect 232 1543 234 1553
rect 288 1543 290 1553
rect 300 1544 302 1562
rect 342 1558 348 1559
rect 342 1554 343 1558
rect 347 1554 348 1558
rect 342 1553 348 1554
rect 298 1543 304 1544
rect 344 1543 346 1553
rect 380 1544 382 1562
rect 724 1560 726 1590
rect 854 1589 860 1590
rect 854 1585 855 1589
rect 859 1585 860 1589
rect 854 1584 860 1585
rect 751 1582 755 1583
rect 751 1576 755 1578
rect 855 1582 859 1584
rect 855 1576 859 1578
rect 750 1575 756 1576
rect 750 1571 751 1575
rect 755 1571 756 1575
rect 750 1570 756 1571
rect 854 1575 860 1576
rect 854 1571 855 1575
rect 859 1571 860 1575
rect 854 1570 860 1571
rect 730 1567 736 1568
rect 730 1563 731 1567
rect 735 1563 736 1567
rect 730 1562 736 1563
rect 722 1559 728 1560
rect 398 1558 404 1559
rect 398 1554 399 1558
rect 403 1554 404 1558
rect 398 1553 404 1554
rect 454 1558 460 1559
rect 454 1554 455 1558
rect 459 1554 460 1558
rect 454 1553 460 1554
rect 510 1558 516 1559
rect 510 1554 511 1558
rect 515 1554 516 1558
rect 510 1553 516 1554
rect 574 1558 580 1559
rect 574 1554 575 1558
rect 579 1554 580 1558
rect 574 1553 580 1554
rect 654 1558 660 1559
rect 654 1554 655 1558
rect 659 1554 660 1558
rect 722 1555 723 1559
rect 727 1555 728 1559
rect 722 1554 728 1555
rect 654 1553 660 1554
rect 378 1543 384 1544
rect 400 1543 402 1553
rect 456 1543 458 1553
rect 512 1543 514 1553
rect 554 1543 560 1544
rect 576 1543 578 1553
rect 656 1543 658 1553
rect 223 1542 227 1543
rect 223 1537 227 1538
rect 231 1542 235 1543
rect 231 1537 235 1538
rect 279 1542 283 1543
rect 279 1537 283 1538
rect 287 1542 291 1543
rect 298 1539 299 1543
rect 303 1539 304 1543
rect 298 1538 304 1539
rect 335 1542 339 1543
rect 287 1537 291 1538
rect 335 1537 339 1538
rect 343 1542 347 1543
rect 378 1539 379 1543
rect 383 1539 384 1543
rect 378 1538 384 1539
rect 399 1542 403 1543
rect 343 1537 347 1538
rect 399 1537 403 1538
rect 455 1542 459 1543
rect 455 1537 459 1538
rect 463 1542 467 1543
rect 463 1537 467 1538
rect 511 1542 515 1543
rect 511 1537 515 1538
rect 535 1542 539 1543
rect 554 1539 555 1543
rect 559 1539 560 1543
rect 554 1538 560 1539
rect 575 1542 579 1543
rect 535 1537 539 1538
rect 210 1535 216 1536
rect 210 1531 211 1535
rect 215 1531 216 1535
rect 210 1530 216 1531
rect 212 1516 214 1530
rect 224 1527 226 1537
rect 280 1527 282 1537
rect 336 1527 338 1537
rect 400 1527 402 1537
rect 464 1527 466 1537
rect 470 1531 476 1532
rect 470 1527 471 1531
rect 475 1527 476 1531
rect 536 1527 538 1537
rect 222 1526 228 1527
rect 222 1522 223 1526
rect 227 1522 228 1526
rect 222 1521 228 1522
rect 278 1526 284 1527
rect 278 1522 279 1526
rect 283 1522 284 1526
rect 278 1521 284 1522
rect 334 1526 340 1527
rect 334 1522 335 1526
rect 339 1522 340 1526
rect 334 1521 340 1522
rect 398 1526 404 1527
rect 398 1522 399 1526
rect 403 1522 404 1526
rect 398 1521 404 1522
rect 462 1526 468 1527
rect 470 1526 476 1527
rect 534 1526 540 1527
rect 462 1522 463 1526
rect 467 1522 468 1526
rect 462 1521 468 1522
rect 210 1515 216 1516
rect 210 1511 211 1515
rect 215 1511 216 1515
rect 210 1510 216 1511
rect 318 1515 324 1516
rect 318 1511 319 1515
rect 323 1511 324 1515
rect 318 1510 324 1511
rect 350 1515 356 1516
rect 350 1511 351 1515
rect 355 1511 356 1515
rect 350 1510 356 1511
rect 222 1509 228 1510
rect 222 1505 223 1509
rect 227 1505 228 1509
rect 222 1504 228 1505
rect 278 1509 284 1510
rect 278 1505 279 1509
rect 283 1505 284 1509
rect 278 1504 284 1505
rect 224 1499 226 1504
rect 280 1499 282 1504
rect 207 1498 211 1499
rect 207 1493 211 1494
rect 223 1498 227 1499
rect 223 1493 227 1494
rect 239 1498 243 1499
rect 239 1493 243 1494
rect 271 1498 275 1499
rect 271 1493 275 1494
rect 279 1498 283 1499
rect 279 1493 283 1494
rect 303 1498 307 1499
rect 303 1493 307 1494
rect 208 1476 210 1493
rect 240 1476 242 1493
rect 272 1476 274 1493
rect 304 1476 306 1493
rect 206 1475 212 1476
rect 206 1471 207 1475
rect 211 1471 212 1475
rect 206 1470 212 1471
rect 238 1475 244 1476
rect 238 1471 239 1475
rect 243 1471 244 1475
rect 238 1470 244 1471
rect 270 1475 276 1476
rect 270 1471 271 1475
rect 275 1471 276 1475
rect 270 1470 276 1471
rect 302 1475 308 1476
rect 302 1471 303 1475
rect 307 1471 308 1475
rect 302 1470 308 1471
rect 206 1458 212 1459
rect 206 1454 207 1458
rect 211 1454 212 1458
rect 206 1453 212 1454
rect 238 1458 244 1459
rect 238 1454 239 1458
rect 243 1454 244 1458
rect 238 1453 244 1454
rect 270 1458 276 1459
rect 270 1454 271 1458
rect 275 1454 276 1458
rect 270 1453 276 1454
rect 302 1458 308 1459
rect 302 1454 303 1458
rect 307 1454 308 1458
rect 302 1453 308 1454
rect 208 1431 210 1453
rect 240 1431 242 1453
rect 272 1431 274 1453
rect 304 1431 306 1453
rect 320 1452 322 1510
rect 334 1509 340 1510
rect 334 1505 335 1509
rect 339 1505 340 1509
rect 334 1504 340 1505
rect 336 1499 338 1504
rect 335 1498 339 1499
rect 335 1493 339 1494
rect 336 1476 338 1493
rect 334 1475 340 1476
rect 334 1471 335 1475
rect 339 1471 340 1475
rect 334 1470 340 1471
rect 334 1458 340 1459
rect 334 1454 335 1458
rect 339 1454 340 1458
rect 334 1453 340 1454
rect 318 1451 324 1452
rect 318 1447 319 1451
rect 323 1447 324 1451
rect 318 1446 324 1447
rect 336 1431 338 1453
rect 352 1452 354 1510
rect 398 1509 404 1510
rect 398 1505 399 1509
rect 403 1505 404 1509
rect 398 1504 404 1505
rect 462 1509 468 1510
rect 462 1505 463 1509
rect 467 1505 468 1509
rect 462 1504 468 1505
rect 400 1499 402 1504
rect 464 1499 466 1504
rect 367 1498 371 1499
rect 367 1493 371 1494
rect 399 1498 403 1499
rect 399 1493 403 1494
rect 431 1498 435 1499
rect 431 1493 435 1494
rect 463 1498 467 1499
rect 463 1493 467 1494
rect 368 1476 370 1493
rect 382 1483 388 1484
rect 382 1479 383 1483
rect 387 1479 388 1483
rect 382 1478 388 1479
rect 366 1475 372 1476
rect 366 1471 367 1475
rect 371 1471 372 1475
rect 366 1470 372 1471
rect 366 1458 372 1459
rect 366 1454 367 1458
rect 371 1454 372 1458
rect 366 1453 372 1454
rect 350 1451 356 1452
rect 350 1447 351 1451
rect 355 1447 356 1451
rect 350 1446 356 1447
rect 368 1431 370 1453
rect 384 1452 386 1478
rect 400 1476 402 1493
rect 432 1476 434 1493
rect 464 1476 466 1493
rect 472 1484 474 1526
rect 534 1522 535 1526
rect 539 1522 540 1526
rect 534 1521 540 1522
rect 556 1516 558 1538
rect 575 1537 579 1538
rect 607 1542 611 1543
rect 607 1537 611 1538
rect 655 1542 659 1543
rect 655 1537 659 1538
rect 687 1542 691 1543
rect 687 1537 691 1538
rect 608 1527 610 1537
rect 646 1535 652 1536
rect 638 1531 644 1532
rect 638 1527 639 1531
rect 643 1527 644 1531
rect 646 1531 647 1535
rect 651 1531 652 1535
rect 646 1530 652 1531
rect 606 1526 612 1527
rect 638 1526 644 1527
rect 606 1522 607 1526
rect 611 1522 612 1526
rect 606 1521 612 1522
rect 554 1515 560 1516
rect 554 1511 555 1515
rect 559 1511 560 1515
rect 554 1510 560 1511
rect 534 1509 540 1510
rect 534 1505 535 1509
rect 539 1505 540 1509
rect 534 1504 540 1505
rect 606 1509 612 1510
rect 606 1505 607 1509
rect 611 1505 612 1509
rect 606 1504 612 1505
rect 536 1499 538 1504
rect 608 1499 610 1504
rect 495 1498 499 1499
rect 495 1493 499 1494
rect 527 1498 531 1499
rect 527 1493 531 1494
rect 535 1498 539 1499
rect 535 1493 539 1494
rect 559 1498 563 1499
rect 559 1493 563 1494
rect 591 1498 595 1499
rect 591 1493 595 1494
rect 607 1498 611 1499
rect 607 1493 611 1494
rect 623 1498 627 1499
rect 623 1493 627 1494
rect 470 1483 476 1484
rect 470 1479 471 1483
rect 475 1479 476 1483
rect 470 1478 476 1479
rect 496 1476 498 1493
rect 528 1476 530 1493
rect 560 1476 562 1493
rect 592 1476 594 1493
rect 624 1476 626 1493
rect 398 1475 404 1476
rect 398 1471 399 1475
rect 403 1471 404 1475
rect 398 1470 404 1471
rect 430 1475 436 1476
rect 430 1471 431 1475
rect 435 1471 436 1475
rect 430 1470 436 1471
rect 462 1475 468 1476
rect 462 1471 463 1475
rect 467 1471 468 1475
rect 462 1470 468 1471
rect 494 1475 500 1476
rect 494 1471 495 1475
rect 499 1471 500 1475
rect 494 1470 500 1471
rect 526 1475 532 1476
rect 526 1471 527 1475
rect 531 1471 532 1475
rect 526 1470 532 1471
rect 558 1475 564 1476
rect 558 1471 559 1475
rect 563 1471 564 1475
rect 558 1470 564 1471
rect 590 1475 596 1476
rect 590 1471 591 1475
rect 595 1471 596 1475
rect 590 1470 596 1471
rect 622 1475 628 1476
rect 622 1471 623 1475
rect 627 1471 628 1475
rect 622 1470 628 1471
rect 640 1468 642 1526
rect 648 1516 650 1530
rect 688 1527 690 1537
rect 732 1536 734 1562
rect 750 1558 756 1559
rect 750 1554 751 1558
rect 755 1554 756 1558
rect 750 1553 756 1554
rect 854 1558 860 1559
rect 854 1554 855 1558
rect 859 1554 860 1558
rect 854 1553 860 1554
rect 752 1543 754 1553
rect 758 1551 764 1552
rect 758 1547 759 1551
rect 763 1547 764 1551
rect 758 1546 764 1547
rect 751 1542 755 1543
rect 751 1537 755 1538
rect 730 1535 736 1536
rect 730 1531 731 1535
rect 735 1531 736 1535
rect 730 1530 736 1531
rect 686 1526 692 1527
rect 686 1522 687 1526
rect 691 1522 692 1526
rect 686 1521 692 1522
rect 646 1515 652 1516
rect 646 1511 647 1515
rect 651 1511 652 1515
rect 646 1510 652 1511
rect 718 1515 724 1516
rect 718 1511 719 1515
rect 723 1511 724 1515
rect 718 1510 724 1511
rect 686 1509 692 1510
rect 686 1505 687 1509
rect 691 1505 692 1509
rect 686 1504 692 1505
rect 688 1499 690 1504
rect 663 1498 667 1499
rect 663 1493 667 1494
rect 687 1498 691 1499
rect 687 1493 691 1494
rect 703 1498 707 1499
rect 703 1493 707 1494
rect 664 1476 666 1493
rect 704 1476 706 1493
rect 662 1475 668 1476
rect 662 1471 663 1475
rect 667 1471 668 1475
rect 662 1470 668 1471
rect 702 1475 708 1476
rect 702 1471 703 1475
rect 707 1471 708 1475
rect 702 1470 708 1471
rect 446 1467 452 1468
rect 446 1463 447 1467
rect 451 1463 452 1467
rect 446 1462 452 1463
rect 542 1467 548 1468
rect 542 1463 543 1467
rect 547 1463 548 1467
rect 542 1462 548 1463
rect 638 1467 644 1468
rect 638 1463 639 1467
rect 643 1463 644 1467
rect 638 1462 644 1463
rect 682 1467 688 1468
rect 682 1463 683 1467
rect 687 1463 688 1467
rect 682 1462 688 1463
rect 398 1458 404 1459
rect 398 1454 399 1458
rect 403 1454 404 1458
rect 398 1453 404 1454
rect 430 1458 436 1459
rect 430 1454 431 1458
rect 435 1454 436 1458
rect 430 1453 436 1454
rect 382 1451 388 1452
rect 382 1447 383 1451
rect 387 1447 388 1451
rect 382 1446 388 1447
rect 400 1431 402 1453
rect 432 1431 434 1453
rect 199 1430 203 1431
rect 199 1425 203 1426
rect 207 1430 211 1431
rect 207 1425 211 1426
rect 231 1430 235 1431
rect 231 1425 235 1426
rect 239 1430 243 1431
rect 239 1425 243 1426
rect 263 1430 267 1431
rect 263 1425 267 1426
rect 271 1430 275 1431
rect 271 1425 275 1426
rect 295 1430 299 1431
rect 295 1425 299 1426
rect 303 1430 307 1431
rect 303 1425 307 1426
rect 327 1430 331 1431
rect 327 1425 331 1426
rect 335 1430 339 1431
rect 335 1425 339 1426
rect 359 1430 363 1431
rect 359 1425 363 1426
rect 367 1430 371 1431
rect 367 1425 371 1426
rect 391 1430 395 1431
rect 391 1425 395 1426
rect 399 1430 403 1431
rect 399 1425 403 1426
rect 423 1430 427 1431
rect 423 1425 427 1426
rect 431 1430 435 1431
rect 431 1425 435 1426
rect 200 1391 202 1425
rect 232 1391 234 1425
rect 264 1391 266 1425
rect 296 1391 298 1425
rect 328 1391 330 1425
rect 360 1391 362 1425
rect 378 1395 384 1396
rect 378 1391 379 1395
rect 383 1391 384 1395
rect 392 1391 394 1425
rect 424 1391 426 1425
rect 448 1404 450 1462
rect 462 1458 468 1459
rect 462 1454 463 1458
rect 467 1454 468 1458
rect 462 1453 468 1454
rect 494 1458 500 1459
rect 494 1454 495 1458
rect 499 1454 500 1458
rect 494 1453 500 1454
rect 526 1458 532 1459
rect 526 1454 527 1458
rect 531 1454 532 1458
rect 526 1453 532 1454
rect 464 1431 466 1453
rect 496 1431 498 1453
rect 528 1431 530 1453
rect 534 1451 540 1452
rect 534 1447 535 1451
rect 539 1447 540 1451
rect 534 1446 540 1447
rect 455 1430 459 1431
rect 455 1425 459 1426
rect 463 1430 467 1431
rect 463 1425 467 1426
rect 487 1430 491 1431
rect 487 1425 491 1426
rect 495 1430 499 1431
rect 495 1425 499 1426
rect 519 1430 523 1431
rect 519 1425 523 1426
rect 527 1430 531 1431
rect 536 1428 538 1446
rect 527 1425 531 1426
rect 534 1427 540 1428
rect 446 1403 452 1404
rect 446 1399 447 1403
rect 451 1399 452 1403
rect 446 1398 452 1399
rect 456 1391 458 1425
rect 488 1391 490 1425
rect 520 1391 522 1425
rect 534 1423 535 1427
rect 539 1423 540 1427
rect 534 1422 540 1423
rect 544 1404 546 1462
rect 558 1458 564 1459
rect 558 1454 559 1458
rect 563 1454 564 1458
rect 558 1453 564 1454
rect 590 1458 596 1459
rect 590 1454 591 1458
rect 595 1454 596 1458
rect 590 1453 596 1454
rect 622 1458 628 1459
rect 622 1454 623 1458
rect 627 1454 628 1458
rect 622 1453 628 1454
rect 662 1458 668 1459
rect 662 1454 663 1458
rect 667 1454 668 1458
rect 662 1453 668 1454
rect 684 1453 686 1462
rect 702 1458 708 1459
rect 702 1454 703 1458
rect 707 1454 708 1458
rect 702 1453 708 1454
rect 560 1431 562 1453
rect 592 1431 594 1453
rect 624 1431 626 1453
rect 664 1431 666 1453
rect 684 1451 690 1453
rect 551 1430 555 1431
rect 551 1425 555 1426
rect 559 1430 563 1431
rect 559 1425 563 1426
rect 583 1430 587 1431
rect 583 1425 587 1426
rect 591 1430 595 1431
rect 591 1425 595 1426
rect 615 1430 619 1431
rect 615 1425 619 1426
rect 623 1430 627 1431
rect 623 1425 627 1426
rect 647 1430 651 1431
rect 647 1425 651 1426
rect 663 1430 667 1431
rect 679 1430 683 1431
rect 663 1425 667 1426
rect 670 1427 676 1428
rect 542 1403 548 1404
rect 542 1399 543 1403
rect 547 1399 548 1403
rect 542 1398 548 1399
rect 552 1391 554 1425
rect 584 1391 586 1425
rect 616 1391 618 1425
rect 648 1391 650 1425
rect 670 1423 671 1427
rect 675 1423 676 1427
rect 679 1425 683 1426
rect 670 1422 676 1423
rect 198 1390 204 1391
rect 198 1386 199 1390
rect 203 1386 204 1390
rect 198 1385 204 1386
rect 230 1390 236 1391
rect 230 1386 231 1390
rect 235 1386 236 1390
rect 230 1385 236 1386
rect 262 1390 268 1391
rect 262 1386 263 1390
rect 267 1386 268 1390
rect 262 1385 268 1386
rect 294 1390 300 1391
rect 294 1386 295 1390
rect 299 1386 300 1390
rect 294 1385 300 1386
rect 326 1390 332 1391
rect 326 1386 327 1390
rect 331 1386 332 1390
rect 326 1385 332 1386
rect 358 1390 364 1391
rect 378 1390 384 1391
rect 390 1390 396 1391
rect 358 1386 359 1390
rect 363 1386 364 1390
rect 358 1385 364 1386
rect 346 1379 352 1380
rect 346 1375 347 1379
rect 351 1375 352 1379
rect 346 1374 352 1375
rect 198 1373 204 1374
rect 198 1369 199 1373
rect 203 1369 204 1373
rect 198 1368 204 1369
rect 230 1373 236 1374
rect 230 1369 231 1373
rect 235 1369 236 1373
rect 230 1368 236 1369
rect 262 1373 268 1374
rect 262 1369 263 1373
rect 267 1369 268 1373
rect 262 1368 268 1369
rect 294 1373 300 1374
rect 294 1369 295 1373
rect 299 1369 300 1373
rect 294 1368 300 1369
rect 326 1373 332 1374
rect 326 1369 327 1373
rect 331 1369 332 1373
rect 326 1368 332 1369
rect 200 1351 202 1368
rect 232 1351 234 1368
rect 264 1351 266 1368
rect 296 1351 298 1368
rect 328 1351 330 1368
rect 199 1350 203 1351
rect 199 1345 203 1346
rect 231 1350 235 1351
rect 231 1345 235 1346
rect 263 1350 267 1351
rect 263 1345 267 1346
rect 295 1350 299 1351
rect 295 1345 299 1346
rect 327 1350 331 1351
rect 327 1345 331 1346
rect 200 1320 202 1345
rect 232 1320 234 1345
rect 264 1320 266 1345
rect 296 1320 298 1345
rect 328 1320 330 1345
rect 198 1319 204 1320
rect 198 1315 199 1319
rect 203 1315 204 1319
rect 198 1314 204 1315
rect 230 1319 236 1320
rect 230 1315 231 1319
rect 235 1315 236 1319
rect 230 1314 236 1315
rect 262 1319 268 1320
rect 262 1315 263 1319
rect 267 1315 268 1319
rect 262 1314 268 1315
rect 294 1319 300 1320
rect 294 1315 295 1319
rect 299 1315 300 1319
rect 294 1314 300 1315
rect 326 1319 332 1320
rect 326 1315 327 1319
rect 331 1315 332 1319
rect 326 1314 332 1315
rect 348 1304 350 1374
rect 358 1373 364 1374
rect 358 1369 359 1373
rect 363 1369 364 1373
rect 358 1368 364 1369
rect 380 1368 382 1390
rect 390 1386 391 1390
rect 395 1386 396 1390
rect 390 1385 396 1386
rect 422 1390 428 1391
rect 422 1386 423 1390
rect 427 1386 428 1390
rect 422 1385 428 1386
rect 454 1390 460 1391
rect 454 1386 455 1390
rect 459 1386 460 1390
rect 454 1385 460 1386
rect 486 1390 492 1391
rect 486 1386 487 1390
rect 491 1386 492 1390
rect 486 1385 492 1386
rect 518 1390 524 1391
rect 518 1386 519 1390
rect 523 1386 524 1390
rect 518 1385 524 1386
rect 550 1390 556 1391
rect 550 1386 551 1390
rect 555 1386 556 1390
rect 550 1385 556 1386
rect 582 1390 588 1391
rect 582 1386 583 1390
rect 587 1386 588 1390
rect 582 1385 588 1386
rect 614 1390 620 1391
rect 614 1386 615 1390
rect 619 1386 620 1390
rect 614 1385 620 1386
rect 646 1390 652 1391
rect 646 1386 647 1390
rect 651 1386 652 1390
rect 646 1385 652 1386
rect 470 1379 476 1380
rect 470 1375 471 1379
rect 475 1375 476 1379
rect 470 1374 476 1375
rect 566 1379 572 1380
rect 566 1375 567 1379
rect 571 1375 572 1379
rect 566 1374 572 1375
rect 662 1379 668 1380
rect 662 1375 663 1379
rect 667 1375 668 1379
rect 662 1374 668 1375
rect 390 1373 396 1374
rect 390 1369 391 1373
rect 395 1369 396 1373
rect 390 1368 396 1369
rect 422 1373 428 1374
rect 422 1369 423 1373
rect 427 1369 428 1373
rect 422 1368 428 1369
rect 454 1373 460 1374
rect 454 1369 455 1373
rect 459 1369 460 1373
rect 454 1368 460 1369
rect 360 1351 362 1368
rect 378 1367 384 1368
rect 378 1363 379 1367
rect 383 1363 384 1367
rect 378 1362 384 1363
rect 392 1351 394 1368
rect 424 1351 426 1368
rect 456 1351 458 1368
rect 359 1350 363 1351
rect 359 1345 363 1346
rect 391 1350 395 1351
rect 391 1345 395 1346
rect 423 1350 427 1351
rect 423 1345 427 1346
rect 455 1350 459 1351
rect 455 1345 459 1346
rect 360 1320 362 1345
rect 392 1320 394 1345
rect 424 1320 426 1345
rect 456 1320 458 1345
rect 358 1319 364 1320
rect 358 1315 359 1319
rect 363 1315 364 1319
rect 358 1314 364 1315
rect 390 1319 396 1320
rect 390 1315 391 1319
rect 395 1315 396 1319
rect 390 1314 396 1315
rect 422 1319 428 1320
rect 422 1315 423 1319
rect 427 1315 428 1319
rect 422 1314 428 1315
rect 454 1319 460 1320
rect 454 1315 455 1319
rect 459 1315 460 1319
rect 454 1314 460 1315
rect 346 1303 352 1304
rect 198 1302 204 1303
rect 198 1298 199 1302
rect 203 1298 204 1302
rect 198 1297 204 1298
rect 230 1302 236 1303
rect 230 1298 231 1302
rect 235 1298 236 1302
rect 230 1297 236 1298
rect 262 1302 268 1303
rect 262 1298 263 1302
rect 267 1298 268 1302
rect 262 1297 268 1298
rect 294 1302 300 1303
rect 294 1298 295 1302
rect 299 1298 300 1302
rect 294 1297 300 1298
rect 326 1302 332 1303
rect 326 1298 327 1302
rect 331 1298 332 1302
rect 346 1299 347 1303
rect 351 1299 352 1303
rect 346 1298 352 1299
rect 358 1302 364 1303
rect 358 1298 359 1302
rect 363 1298 364 1302
rect 326 1297 332 1298
rect 358 1297 364 1298
rect 390 1302 396 1303
rect 390 1298 391 1302
rect 395 1298 396 1302
rect 390 1297 396 1298
rect 422 1302 428 1303
rect 422 1298 423 1302
rect 427 1298 428 1302
rect 422 1297 428 1298
rect 454 1302 460 1303
rect 454 1298 455 1302
rect 459 1298 460 1302
rect 454 1297 460 1298
rect 186 1279 192 1280
rect 186 1275 187 1279
rect 191 1275 192 1279
rect 186 1274 192 1275
rect 200 1263 202 1297
rect 232 1263 234 1297
rect 264 1263 266 1297
rect 296 1263 298 1297
rect 328 1263 330 1297
rect 360 1263 362 1297
rect 392 1263 394 1297
rect 424 1263 426 1297
rect 456 1263 458 1297
rect 472 1288 474 1374
rect 486 1373 492 1374
rect 486 1369 487 1373
rect 491 1369 492 1373
rect 486 1368 492 1369
rect 518 1373 524 1374
rect 518 1369 519 1373
rect 523 1369 524 1373
rect 518 1368 524 1369
rect 550 1373 556 1374
rect 550 1369 551 1373
rect 555 1369 556 1373
rect 550 1368 556 1369
rect 568 1368 570 1374
rect 582 1373 588 1374
rect 582 1369 583 1373
rect 587 1369 588 1373
rect 582 1368 588 1369
rect 614 1373 620 1374
rect 614 1369 615 1373
rect 619 1369 620 1373
rect 614 1368 620 1369
rect 646 1373 652 1374
rect 646 1369 647 1373
rect 651 1369 652 1373
rect 646 1368 652 1369
rect 488 1351 490 1368
rect 520 1351 522 1368
rect 552 1351 554 1368
rect 566 1367 572 1368
rect 566 1363 567 1367
rect 571 1363 572 1367
rect 566 1362 572 1363
rect 584 1351 586 1368
rect 616 1351 618 1368
rect 648 1351 650 1368
rect 487 1350 491 1351
rect 487 1345 491 1346
rect 519 1350 523 1351
rect 519 1345 523 1346
rect 551 1350 555 1351
rect 551 1345 555 1346
rect 583 1350 587 1351
rect 583 1345 587 1346
rect 615 1350 619 1351
rect 615 1345 619 1346
rect 647 1350 651 1351
rect 647 1345 651 1346
rect 488 1320 490 1345
rect 520 1320 522 1345
rect 552 1320 554 1345
rect 584 1320 586 1345
rect 616 1320 618 1345
rect 648 1320 650 1345
rect 486 1319 492 1320
rect 486 1315 487 1319
rect 491 1315 492 1319
rect 486 1314 492 1315
rect 518 1319 524 1320
rect 518 1315 519 1319
rect 523 1315 524 1319
rect 518 1314 524 1315
rect 550 1319 556 1320
rect 550 1315 551 1319
rect 555 1315 556 1319
rect 550 1314 556 1315
rect 582 1319 588 1320
rect 582 1315 583 1319
rect 587 1315 588 1319
rect 582 1314 588 1315
rect 614 1319 620 1320
rect 614 1315 615 1319
rect 619 1315 620 1319
rect 614 1314 620 1315
rect 646 1319 652 1320
rect 646 1315 647 1319
rect 651 1315 652 1319
rect 646 1314 652 1315
rect 626 1311 632 1312
rect 626 1307 627 1311
rect 631 1307 632 1311
rect 626 1306 632 1307
rect 486 1302 492 1303
rect 486 1298 487 1302
rect 491 1298 492 1302
rect 486 1297 492 1298
rect 518 1302 524 1303
rect 518 1298 519 1302
rect 523 1298 524 1302
rect 518 1297 524 1298
rect 550 1302 556 1303
rect 550 1298 551 1302
rect 555 1298 556 1302
rect 550 1297 556 1298
rect 582 1302 588 1303
rect 582 1298 583 1302
rect 587 1298 588 1302
rect 582 1297 588 1298
rect 614 1302 620 1303
rect 614 1298 615 1302
rect 619 1298 620 1302
rect 614 1297 620 1298
rect 470 1287 476 1288
rect 470 1283 471 1287
rect 475 1283 476 1287
rect 470 1282 476 1283
rect 488 1263 490 1297
rect 520 1263 522 1297
rect 552 1263 554 1297
rect 574 1271 580 1272
rect 574 1267 575 1271
rect 579 1267 580 1271
rect 574 1266 580 1267
rect 199 1262 203 1263
rect 199 1257 203 1258
rect 231 1262 235 1263
rect 231 1257 235 1258
rect 263 1262 267 1263
rect 263 1257 267 1258
rect 295 1262 299 1263
rect 295 1257 299 1258
rect 327 1262 331 1263
rect 327 1257 331 1258
rect 359 1262 363 1263
rect 359 1257 363 1258
rect 391 1262 395 1263
rect 391 1257 395 1258
rect 423 1262 427 1263
rect 423 1257 427 1258
rect 455 1262 459 1263
rect 455 1257 459 1258
rect 487 1262 491 1263
rect 487 1257 491 1258
rect 519 1262 523 1263
rect 519 1257 523 1258
rect 551 1262 555 1263
rect 551 1257 555 1258
rect 190 1235 196 1236
rect 190 1231 191 1235
rect 195 1231 196 1235
rect 190 1230 196 1231
rect 192 1076 194 1230
rect 200 1195 202 1257
rect 232 1195 234 1257
rect 264 1195 266 1257
rect 296 1195 298 1257
rect 328 1195 330 1257
rect 360 1195 362 1257
rect 392 1195 394 1257
rect 424 1195 426 1257
rect 456 1195 458 1257
rect 488 1195 490 1257
rect 520 1195 522 1257
rect 552 1195 554 1257
rect 198 1194 204 1195
rect 198 1190 199 1194
rect 203 1190 204 1194
rect 198 1189 204 1190
rect 230 1194 236 1195
rect 230 1190 231 1194
rect 235 1190 236 1194
rect 230 1189 236 1190
rect 262 1194 268 1195
rect 262 1190 263 1194
rect 267 1190 268 1194
rect 262 1189 268 1190
rect 294 1194 300 1195
rect 294 1190 295 1194
rect 299 1190 300 1194
rect 294 1189 300 1190
rect 326 1194 332 1195
rect 326 1190 327 1194
rect 331 1190 332 1194
rect 326 1189 332 1190
rect 358 1194 364 1195
rect 358 1190 359 1194
rect 363 1190 364 1194
rect 358 1189 364 1190
rect 390 1194 396 1195
rect 390 1190 391 1194
rect 395 1190 396 1194
rect 390 1189 396 1190
rect 422 1194 428 1195
rect 422 1190 423 1194
rect 427 1190 428 1194
rect 422 1189 428 1190
rect 454 1194 460 1195
rect 454 1190 455 1194
rect 459 1190 460 1194
rect 454 1189 460 1190
rect 486 1194 492 1195
rect 486 1190 487 1194
rect 491 1190 492 1194
rect 486 1189 492 1190
rect 518 1194 524 1195
rect 518 1190 519 1194
rect 523 1190 524 1194
rect 518 1189 524 1190
rect 550 1194 556 1195
rect 550 1190 551 1194
rect 555 1190 556 1194
rect 550 1189 556 1190
rect 566 1183 572 1184
rect 566 1179 567 1183
rect 571 1179 572 1183
rect 566 1178 572 1179
rect 198 1177 204 1178
rect 198 1173 199 1177
rect 203 1173 204 1177
rect 198 1172 204 1173
rect 230 1177 236 1178
rect 230 1173 231 1177
rect 235 1173 236 1177
rect 230 1172 236 1173
rect 262 1177 268 1178
rect 262 1173 263 1177
rect 267 1173 268 1177
rect 262 1172 268 1173
rect 294 1177 300 1178
rect 294 1173 295 1177
rect 299 1173 300 1177
rect 294 1172 300 1173
rect 326 1177 332 1178
rect 326 1173 327 1177
rect 331 1173 332 1177
rect 326 1172 332 1173
rect 358 1177 364 1178
rect 358 1173 359 1177
rect 363 1173 364 1177
rect 358 1172 364 1173
rect 390 1177 396 1178
rect 390 1173 391 1177
rect 395 1173 396 1177
rect 390 1172 396 1173
rect 422 1177 428 1178
rect 422 1173 423 1177
rect 427 1173 428 1177
rect 422 1172 428 1173
rect 454 1177 460 1178
rect 454 1173 455 1177
rect 459 1173 460 1177
rect 454 1172 460 1173
rect 486 1177 492 1178
rect 486 1173 487 1177
rect 491 1173 492 1177
rect 486 1172 492 1173
rect 518 1177 524 1178
rect 518 1173 519 1177
rect 523 1173 524 1177
rect 518 1172 524 1173
rect 550 1177 556 1178
rect 550 1173 551 1177
rect 555 1173 556 1177
rect 550 1172 556 1173
rect 200 1151 202 1172
rect 232 1151 234 1172
rect 264 1151 266 1172
rect 296 1151 298 1172
rect 328 1151 330 1172
rect 360 1151 362 1172
rect 392 1151 394 1172
rect 414 1151 420 1152
rect 424 1151 426 1172
rect 442 1171 448 1172
rect 442 1167 443 1171
rect 447 1167 448 1171
rect 442 1166 448 1167
rect 199 1150 203 1151
rect 199 1145 203 1146
rect 231 1150 235 1151
rect 231 1145 235 1146
rect 263 1150 267 1151
rect 263 1145 267 1146
rect 295 1150 299 1151
rect 295 1145 299 1146
rect 327 1150 331 1151
rect 327 1145 331 1146
rect 359 1150 363 1151
rect 359 1145 363 1146
rect 391 1150 395 1151
rect 414 1147 415 1151
rect 419 1147 420 1151
rect 414 1146 420 1147
rect 423 1150 427 1151
rect 391 1145 395 1146
rect 200 1124 202 1145
rect 232 1124 234 1145
rect 264 1124 266 1145
rect 282 1131 288 1132
rect 282 1127 283 1131
rect 287 1127 288 1131
rect 282 1126 288 1127
rect 198 1123 204 1124
rect 198 1119 199 1123
rect 203 1119 204 1123
rect 198 1118 204 1119
rect 230 1123 236 1124
rect 230 1119 231 1123
rect 235 1119 236 1123
rect 230 1118 236 1119
rect 262 1123 268 1124
rect 262 1119 263 1123
rect 267 1119 268 1123
rect 262 1118 268 1119
rect 246 1115 252 1116
rect 246 1111 247 1115
rect 251 1111 252 1115
rect 246 1110 252 1111
rect 198 1106 204 1107
rect 198 1102 199 1106
rect 203 1102 204 1106
rect 198 1101 204 1102
rect 230 1106 236 1107
rect 230 1102 231 1106
rect 235 1102 236 1106
rect 230 1101 236 1102
rect 190 1075 196 1076
rect 190 1071 191 1075
rect 195 1071 196 1075
rect 190 1070 196 1071
rect 187 1060 191 1061
rect 187 1055 191 1056
rect 179 1044 183 1045
rect 179 1039 183 1040
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 135 1034 139 1035
rect 135 1029 139 1030
rect 167 1034 171 1035
rect 167 1029 171 1030
rect 112 997 114 1029
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 136 995 138 1029
rect 168 995 170 1029
rect 110 991 116 992
rect 134 994 140 995
rect 134 990 135 994
rect 139 990 140 994
rect 134 989 140 990
rect 166 994 172 995
rect 166 990 167 994
rect 171 990 172 994
rect 166 989 172 990
rect 150 983 156 984
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 150 979 151 983
rect 155 979 156 983
rect 150 978 156 979
rect 110 974 116 975
rect 134 977 140 978
rect 112 955 114 974
rect 134 973 135 977
rect 139 973 140 977
rect 134 972 140 973
rect 136 955 138 972
rect 111 954 115 955
rect 111 949 115 950
rect 135 954 139 955
rect 135 949 139 950
rect 112 922 114 949
rect 136 924 138 949
rect 134 923 140 924
rect 110 921 116 922
rect 110 917 111 921
rect 115 917 116 921
rect 134 919 135 923
rect 139 919 140 923
rect 134 918 140 919
rect 110 916 116 917
rect 134 906 140 907
rect 110 904 116 905
rect 110 900 111 904
rect 115 900 116 904
rect 134 902 135 906
rect 139 902 140 906
rect 134 901 140 902
rect 110 899 116 900
rect 112 839 114 899
rect 136 839 138 901
rect 152 900 154 978
rect 166 977 172 978
rect 166 973 167 977
rect 171 973 172 977
rect 166 972 172 973
rect 168 955 170 972
rect 167 954 171 955
rect 167 949 171 950
rect 168 924 170 949
rect 166 923 172 924
rect 166 919 167 923
rect 171 919 172 923
rect 166 918 172 919
rect 188 916 190 1055
rect 200 1035 202 1101
rect 232 1035 234 1101
rect 199 1034 203 1035
rect 199 1029 203 1030
rect 231 1034 235 1035
rect 231 1029 235 1030
rect 200 995 202 1029
rect 232 995 234 1029
rect 248 1008 250 1110
rect 262 1106 268 1107
rect 262 1102 263 1106
rect 267 1102 268 1106
rect 262 1101 268 1102
rect 264 1035 266 1101
rect 284 1100 286 1126
rect 296 1124 298 1145
rect 328 1124 330 1145
rect 360 1124 362 1145
rect 392 1124 394 1145
rect 294 1123 300 1124
rect 294 1119 295 1123
rect 299 1119 300 1123
rect 294 1118 300 1119
rect 326 1123 332 1124
rect 326 1119 327 1123
rect 331 1119 332 1123
rect 326 1118 332 1119
rect 358 1123 364 1124
rect 358 1119 359 1123
rect 363 1119 364 1123
rect 358 1118 364 1119
rect 390 1123 396 1124
rect 390 1119 391 1123
rect 395 1119 396 1123
rect 390 1118 396 1119
rect 294 1106 300 1107
rect 294 1102 295 1106
rect 299 1102 300 1106
rect 294 1101 300 1102
rect 326 1106 332 1107
rect 326 1102 327 1106
rect 331 1102 332 1106
rect 326 1101 332 1102
rect 358 1106 364 1107
rect 358 1102 359 1106
rect 363 1102 364 1106
rect 358 1101 364 1102
rect 390 1106 396 1107
rect 390 1102 391 1106
rect 395 1102 396 1106
rect 390 1101 396 1102
rect 282 1099 288 1100
rect 282 1095 283 1099
rect 287 1095 288 1099
rect 282 1094 288 1095
rect 296 1035 298 1101
rect 306 1083 312 1084
rect 306 1079 307 1083
rect 311 1079 312 1083
rect 306 1078 312 1079
rect 263 1034 267 1035
rect 263 1029 267 1030
rect 295 1034 299 1035
rect 295 1029 299 1030
rect 246 1007 252 1008
rect 246 1003 247 1007
rect 251 1003 252 1007
rect 246 1002 252 1003
rect 264 995 266 1029
rect 198 994 204 995
rect 198 990 199 994
rect 203 990 204 994
rect 198 989 204 990
rect 230 994 236 995
rect 230 990 231 994
rect 235 990 236 994
rect 230 989 236 990
rect 262 994 268 995
rect 262 990 263 994
rect 267 990 268 994
rect 262 989 268 990
rect 198 977 204 978
rect 198 973 199 977
rect 203 973 204 977
rect 198 972 204 973
rect 230 977 236 978
rect 230 973 231 977
rect 235 973 236 977
rect 230 972 236 973
rect 262 977 268 978
rect 262 973 263 977
rect 267 973 268 977
rect 262 972 268 973
rect 200 955 202 972
rect 218 955 224 956
rect 232 955 234 972
rect 264 955 266 972
rect 199 954 203 955
rect 218 951 219 955
rect 223 951 224 955
rect 218 950 224 951
rect 231 954 235 955
rect 199 949 203 950
rect 200 925 202 949
rect 198 924 204 925
rect 198 920 199 924
rect 203 920 204 924
rect 198 919 204 920
rect 186 915 192 916
rect 186 911 187 915
rect 191 911 192 915
rect 186 910 192 911
rect 166 906 172 907
rect 166 902 167 906
rect 171 902 172 906
rect 166 901 172 902
rect 150 899 156 900
rect 150 895 151 899
rect 155 895 156 899
rect 150 894 156 895
rect 168 839 170 901
rect 182 899 188 900
rect 182 895 183 899
rect 187 895 188 899
rect 182 894 188 895
rect 111 838 115 839
rect 111 833 115 834
rect 135 838 139 839
rect 135 833 139 834
rect 167 838 171 839
rect 167 833 171 834
rect 112 805 114 833
rect 110 804 116 805
rect 110 800 111 804
rect 115 800 116 804
rect 136 803 138 833
rect 110 799 116 800
rect 134 802 140 803
rect 134 798 135 802
rect 139 798 140 802
rect 134 797 140 798
rect 150 791 156 792
rect 110 787 116 788
rect 110 783 111 787
rect 115 783 116 787
rect 150 787 151 791
rect 155 787 156 791
rect 150 786 156 787
rect 110 782 116 783
rect 134 785 140 786
rect 112 755 114 782
rect 134 781 135 785
rect 139 781 140 785
rect 134 780 140 781
rect 136 755 138 780
rect 111 754 115 755
rect 111 749 115 750
rect 135 754 139 755
rect 135 749 139 750
rect 112 726 114 749
rect 136 729 138 749
rect 134 728 140 729
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 134 724 135 728
rect 139 724 140 728
rect 134 723 140 724
rect 110 720 116 721
rect 110 708 116 709
rect 110 704 111 708
rect 115 704 116 708
rect 110 703 116 704
rect 112 643 114 703
rect 142 690 148 691
rect 142 686 143 690
rect 147 686 148 690
rect 142 685 148 686
rect 144 643 146 685
rect 111 642 115 643
rect 111 637 115 638
rect 135 642 139 643
rect 135 637 139 638
rect 143 642 147 643
rect 143 637 147 638
rect 112 605 114 637
rect 110 604 116 605
rect 110 600 111 604
rect 115 600 116 604
rect 136 603 138 637
rect 152 608 154 786
rect 167 642 171 643
rect 167 637 171 638
rect 150 607 156 608
rect 150 603 151 607
rect 155 603 156 607
rect 168 603 170 637
rect 110 599 116 600
rect 134 602 140 603
rect 150 602 156 603
rect 166 602 172 603
rect 134 598 135 602
rect 139 598 140 602
rect 134 597 140 598
rect 166 598 167 602
rect 171 598 172 602
rect 166 597 172 598
rect 184 592 186 894
rect 206 886 212 887
rect 206 882 207 886
rect 211 882 212 886
rect 206 881 212 882
rect 208 839 210 881
rect 220 876 222 950
rect 231 949 235 950
rect 263 954 267 955
rect 263 949 267 950
rect 279 954 283 955
rect 279 949 283 950
rect 280 929 282 949
rect 278 928 284 929
rect 278 924 279 928
rect 283 924 284 928
rect 278 923 284 924
rect 266 915 272 916
rect 266 911 267 915
rect 271 911 272 915
rect 266 910 272 911
rect 258 907 264 908
rect 258 903 259 907
rect 263 903 264 907
rect 258 902 264 903
rect 260 876 262 902
rect 218 875 224 876
rect 218 871 219 875
rect 223 871 224 875
rect 218 870 224 871
rect 258 875 264 876
rect 258 871 259 875
rect 263 871 264 875
rect 268 872 270 910
rect 278 881 284 882
rect 278 877 279 881
rect 283 877 284 881
rect 278 876 284 877
rect 308 876 310 1078
rect 328 1035 330 1101
rect 360 1035 362 1101
rect 383 1092 387 1093
rect 383 1087 387 1088
rect 327 1034 331 1035
rect 327 1029 331 1030
rect 359 1034 363 1035
rect 359 1029 363 1030
rect 328 998 330 1029
rect 384 1008 386 1087
rect 392 1035 394 1101
rect 399 1044 403 1045
rect 399 1039 403 1040
rect 391 1034 395 1035
rect 391 1029 395 1030
rect 400 1024 402 1039
rect 407 1034 411 1035
rect 407 1029 411 1030
rect 398 1023 404 1024
rect 398 1019 399 1023
rect 403 1019 404 1023
rect 398 1018 404 1019
rect 408 1015 410 1029
rect 416 1024 418 1146
rect 423 1145 427 1146
rect 424 1124 426 1145
rect 422 1123 428 1124
rect 422 1119 423 1123
rect 427 1119 428 1123
rect 422 1118 428 1119
rect 422 1106 428 1107
rect 422 1102 423 1106
rect 427 1102 428 1106
rect 422 1101 428 1102
rect 424 1035 426 1101
rect 444 1100 446 1166
rect 456 1151 458 1172
rect 488 1151 490 1172
rect 520 1151 522 1172
rect 542 1163 548 1164
rect 542 1159 543 1163
rect 547 1159 548 1163
rect 542 1158 548 1159
rect 455 1150 459 1151
rect 455 1145 459 1146
rect 487 1150 491 1151
rect 487 1145 491 1146
rect 519 1150 523 1151
rect 519 1145 523 1146
rect 456 1124 458 1145
rect 488 1124 490 1145
rect 520 1124 522 1145
rect 454 1123 460 1124
rect 454 1119 455 1123
rect 459 1119 460 1123
rect 454 1118 460 1119
rect 486 1123 492 1124
rect 486 1119 487 1123
rect 491 1119 492 1123
rect 486 1118 492 1119
rect 518 1123 524 1124
rect 518 1119 519 1123
rect 523 1119 524 1123
rect 518 1118 524 1119
rect 534 1115 540 1116
rect 534 1111 535 1115
rect 539 1111 540 1115
rect 534 1110 540 1111
rect 454 1106 460 1107
rect 454 1102 455 1106
rect 459 1102 460 1106
rect 454 1101 460 1102
rect 486 1106 492 1107
rect 486 1102 487 1106
rect 491 1102 492 1106
rect 486 1101 492 1102
rect 518 1106 524 1107
rect 518 1102 519 1106
rect 523 1102 524 1106
rect 518 1101 524 1102
rect 442 1099 448 1100
rect 442 1095 443 1099
rect 447 1095 448 1099
rect 442 1094 448 1095
rect 456 1035 458 1101
rect 488 1035 490 1101
rect 520 1035 522 1101
rect 536 1092 538 1110
rect 534 1091 540 1092
rect 534 1087 535 1091
rect 539 1087 540 1091
rect 534 1086 540 1087
rect 423 1034 427 1035
rect 423 1029 427 1030
rect 455 1034 459 1035
rect 455 1029 459 1030
rect 487 1034 491 1035
rect 487 1029 491 1030
rect 503 1034 507 1035
rect 503 1029 507 1030
rect 519 1034 523 1035
rect 519 1029 523 1030
rect 494 1027 500 1028
rect 414 1023 420 1024
rect 414 1019 415 1023
rect 419 1019 420 1023
rect 414 1018 420 1019
rect 458 1023 464 1024
rect 458 1019 459 1023
rect 463 1019 464 1023
rect 494 1023 495 1027
rect 499 1023 500 1027
rect 494 1022 500 1023
rect 458 1018 464 1019
rect 406 1014 412 1015
rect 406 1010 407 1014
rect 411 1010 412 1014
rect 406 1009 412 1010
rect 382 1007 388 1008
rect 382 1003 383 1007
rect 387 1003 388 1007
rect 382 1002 388 1003
rect 358 999 364 1000
rect 326 997 332 998
rect 326 993 327 997
rect 331 993 332 997
rect 358 995 359 999
rect 363 995 364 999
rect 358 994 364 995
rect 326 992 332 993
rect 318 983 324 984
rect 318 979 319 983
rect 323 979 324 983
rect 318 978 324 979
rect 320 964 322 978
rect 342 970 348 971
rect 342 966 343 970
rect 347 966 348 970
rect 342 965 348 966
rect 318 963 324 964
rect 318 959 319 963
rect 323 959 324 963
rect 318 958 324 959
rect 344 955 346 965
rect 319 954 323 955
rect 319 949 323 950
rect 343 954 347 955
rect 343 949 347 950
rect 320 925 322 949
rect 338 943 344 944
rect 338 939 339 943
rect 343 939 344 943
rect 338 938 344 939
rect 318 924 324 925
rect 318 920 319 924
rect 323 920 324 924
rect 318 919 324 920
rect 326 886 332 887
rect 326 882 327 886
rect 331 882 332 886
rect 326 881 332 882
rect 258 870 264 871
rect 266 871 272 872
rect 207 838 211 839
rect 207 833 211 834
rect 220 764 222 870
rect 260 864 262 870
rect 266 867 267 871
rect 271 867 272 871
rect 266 866 272 867
rect 258 863 264 864
rect 258 859 259 863
rect 263 859 264 863
rect 258 858 264 859
rect 280 839 282 876
rect 306 875 312 876
rect 306 871 307 875
rect 311 871 312 875
rect 306 870 312 871
rect 308 856 310 870
rect 306 855 312 856
rect 306 851 307 855
rect 311 851 312 855
rect 306 850 312 851
rect 302 839 308 840
rect 328 839 330 881
rect 340 876 342 938
rect 338 875 344 876
rect 338 871 339 875
rect 343 871 344 875
rect 338 870 344 871
rect 231 838 235 839
rect 231 833 235 834
rect 279 838 283 839
rect 302 835 303 839
rect 307 835 308 839
rect 302 834 308 835
rect 327 838 331 839
rect 279 833 283 834
rect 232 824 234 833
rect 230 823 236 824
rect 230 819 231 823
rect 235 819 236 823
rect 230 818 236 819
rect 230 782 236 783
rect 230 778 231 782
rect 235 778 236 782
rect 230 777 236 778
rect 218 763 224 764
rect 218 759 219 763
rect 223 759 224 763
rect 218 758 224 759
rect 232 755 234 777
rect 215 754 219 755
rect 215 749 219 750
rect 231 754 235 755
rect 231 749 235 750
rect 287 754 291 755
rect 287 749 291 750
rect 216 733 218 749
rect 214 732 220 733
rect 214 728 215 732
rect 219 728 220 732
rect 288 731 290 749
rect 214 727 220 728
rect 286 730 292 731
rect 286 726 287 730
rect 291 726 292 730
rect 286 725 292 726
rect 202 719 208 720
rect 202 715 203 719
rect 207 715 208 719
rect 202 714 208 715
rect 190 687 196 688
rect 190 683 191 687
rect 195 683 196 687
rect 190 682 196 683
rect 150 591 156 592
rect 110 587 116 588
rect 110 583 111 587
rect 115 583 116 587
rect 150 587 151 591
rect 155 587 156 591
rect 150 586 156 587
rect 182 591 188 592
rect 182 587 183 591
rect 187 587 188 591
rect 182 586 188 587
rect 110 582 116 583
rect 134 585 140 586
rect 112 563 114 582
rect 134 581 135 585
rect 139 581 140 585
rect 134 580 140 581
rect 136 563 138 580
rect 111 562 115 563
rect 111 557 115 558
rect 135 562 139 563
rect 135 557 139 558
rect 112 534 114 557
rect 136 536 138 557
rect 134 535 140 536
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 134 531 135 535
rect 139 531 140 535
rect 134 530 140 531
rect 110 528 116 529
rect 134 518 140 519
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 134 514 135 518
rect 139 514 140 518
rect 134 513 140 514
rect 110 511 116 512
rect 112 443 114 511
rect 136 443 138 513
rect 152 512 154 586
rect 166 585 172 586
rect 166 581 167 585
rect 171 581 172 585
rect 166 580 172 581
rect 168 563 170 580
rect 167 562 171 563
rect 167 557 171 558
rect 168 537 170 557
rect 166 536 172 537
rect 166 532 167 536
rect 171 532 172 536
rect 166 531 172 532
rect 150 511 156 512
rect 150 507 151 511
rect 155 507 156 511
rect 150 506 156 507
rect 174 498 180 499
rect 174 494 175 498
rect 179 494 180 498
rect 174 493 180 494
rect 176 443 178 493
rect 192 488 194 682
rect 204 676 206 714
rect 242 711 248 712
rect 242 707 243 711
rect 247 707 248 711
rect 242 706 248 707
rect 214 685 220 686
rect 214 681 215 685
rect 219 681 220 685
rect 214 680 220 681
rect 202 675 208 676
rect 202 671 203 675
rect 207 671 208 675
rect 202 670 208 671
rect 216 643 218 680
rect 234 679 240 680
rect 234 675 235 679
rect 239 675 240 679
rect 234 674 240 675
rect 236 648 238 674
rect 244 668 246 706
rect 278 699 284 700
rect 278 695 279 699
rect 283 695 284 699
rect 278 694 284 695
rect 242 667 248 668
rect 242 663 243 667
rect 247 663 248 667
rect 242 662 248 663
rect 244 660 246 662
rect 242 659 248 660
rect 242 655 243 659
rect 247 655 248 659
rect 242 654 248 655
rect 234 647 240 648
rect 234 643 235 647
rect 239 643 240 647
rect 207 642 211 643
rect 207 637 211 638
rect 215 642 219 643
rect 234 642 240 643
rect 215 637 219 638
rect 208 628 210 637
rect 236 632 238 642
rect 280 632 282 694
rect 286 689 292 690
rect 286 685 287 689
rect 291 685 292 689
rect 286 684 292 685
rect 288 643 290 684
rect 304 680 306 834
rect 327 833 331 834
rect 302 679 308 680
rect 302 675 303 679
rect 307 675 308 679
rect 302 674 308 675
rect 322 679 328 680
rect 322 675 323 679
rect 327 675 328 679
rect 322 674 328 675
rect 314 667 320 668
rect 314 663 315 667
rect 319 663 320 667
rect 314 662 320 663
rect 316 648 318 662
rect 314 647 320 648
rect 314 643 315 647
rect 319 643 320 647
rect 287 642 291 643
rect 314 642 320 643
rect 287 637 291 638
rect 294 639 300 640
rect 234 631 240 632
rect 206 627 212 628
rect 206 623 207 627
rect 211 623 212 627
rect 234 627 235 631
rect 239 627 240 631
rect 234 626 240 627
rect 278 631 284 632
rect 278 627 279 631
rect 283 627 284 631
rect 278 626 284 627
rect 288 623 290 637
rect 294 635 295 639
rect 299 635 300 639
rect 294 634 300 635
rect 206 622 212 623
rect 286 622 292 623
rect 286 618 287 622
rect 291 618 292 622
rect 286 617 292 618
rect 254 607 260 608
rect 254 603 255 607
rect 259 603 260 607
rect 254 602 260 603
rect 206 580 212 581
rect 206 576 207 580
rect 211 576 212 580
rect 206 575 212 576
rect 208 563 210 575
rect 207 562 211 563
rect 207 557 211 558
rect 247 562 251 563
rect 247 557 251 558
rect 248 541 250 557
rect 246 540 252 541
rect 246 536 247 540
rect 251 536 252 540
rect 246 535 252 536
rect 234 527 240 528
rect 234 523 235 527
rect 239 523 240 527
rect 234 522 240 523
rect 186 487 194 488
rect 186 483 187 487
rect 191 484 194 487
rect 236 484 238 522
rect 246 493 252 494
rect 246 489 247 493
rect 251 489 252 493
rect 246 488 252 489
rect 191 483 192 484
rect 186 482 192 483
rect 234 483 240 484
rect 188 460 190 482
rect 234 479 235 483
rect 239 479 240 483
rect 234 478 240 479
rect 186 459 192 460
rect 186 455 187 459
rect 191 455 192 459
rect 186 454 192 455
rect 248 443 250 488
rect 111 442 115 443
rect 111 437 115 438
rect 135 442 139 443
rect 135 437 139 438
rect 167 442 171 443
rect 167 437 171 438
rect 175 442 179 443
rect 175 437 179 438
rect 199 442 203 443
rect 199 437 203 438
rect 231 442 235 443
rect 231 437 235 438
rect 247 442 251 443
rect 247 437 251 438
rect 112 377 114 437
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 136 375 138 437
rect 168 375 170 437
rect 200 375 202 437
rect 232 375 234 437
rect 110 371 116 372
rect 134 374 140 375
rect 134 370 135 374
rect 139 370 140 374
rect 134 369 140 370
rect 166 374 172 375
rect 166 370 167 374
rect 171 370 172 374
rect 166 369 172 370
rect 198 374 204 375
rect 198 370 199 374
rect 203 370 204 374
rect 198 369 204 370
rect 230 374 236 375
rect 230 370 231 374
rect 235 370 236 374
rect 230 369 236 370
rect 247 363 253 364
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 247 359 248 363
rect 252 362 253 363
rect 256 362 258 602
rect 286 599 292 600
rect 286 595 287 599
rect 291 595 292 599
rect 296 596 298 634
rect 306 631 312 632
rect 306 627 307 631
rect 311 627 312 631
rect 306 626 312 627
rect 286 594 292 595
rect 294 595 300 596
rect 288 587 290 594
rect 294 591 295 595
rect 299 591 300 595
rect 294 590 300 591
rect 308 587 310 626
rect 288 585 310 587
rect 278 584 284 585
rect 278 580 279 584
rect 283 580 284 584
rect 278 579 284 580
rect 280 563 282 579
rect 279 562 283 563
rect 279 557 283 558
rect 303 562 307 563
rect 303 557 307 558
rect 304 539 306 557
rect 302 538 308 539
rect 302 534 303 538
rect 307 534 308 538
rect 302 533 308 534
rect 274 519 280 520
rect 274 515 275 519
rect 279 515 280 519
rect 274 514 280 515
rect 276 476 278 514
rect 294 507 300 508
rect 294 503 295 507
rect 299 503 300 507
rect 294 502 300 503
rect 274 475 280 476
rect 274 471 275 475
rect 279 471 280 475
rect 274 470 280 471
rect 276 468 278 470
rect 274 467 280 468
rect 274 463 275 467
rect 279 463 280 467
rect 274 462 280 463
rect 263 442 267 443
rect 263 437 267 438
rect 264 375 266 437
rect 296 404 298 502
rect 302 497 308 498
rect 302 493 303 497
rect 307 493 308 497
rect 302 492 308 493
rect 304 443 306 492
rect 316 480 318 642
rect 324 488 326 674
rect 340 640 342 870
rect 360 840 362 994
rect 398 976 404 977
rect 398 972 399 976
rect 403 972 404 976
rect 398 971 404 972
rect 400 955 402 971
rect 399 954 403 955
rect 399 949 403 950
rect 400 929 402 949
rect 416 944 418 1018
rect 460 996 462 1018
rect 458 995 464 996
rect 458 991 459 995
rect 463 991 464 995
rect 458 990 464 991
rect 496 988 498 1022
rect 504 1020 506 1029
rect 544 1024 546 1158
rect 552 1151 554 1172
rect 551 1150 555 1151
rect 551 1145 555 1146
rect 552 1124 554 1145
rect 550 1123 556 1124
rect 550 1119 551 1123
rect 555 1119 556 1123
rect 550 1118 556 1119
rect 550 1106 556 1107
rect 550 1102 551 1106
rect 555 1102 556 1106
rect 550 1101 556 1102
rect 552 1035 554 1101
rect 568 1100 570 1178
rect 566 1099 572 1100
rect 566 1095 567 1099
rect 571 1095 572 1099
rect 566 1094 572 1095
rect 551 1034 555 1035
rect 551 1029 555 1030
rect 542 1023 548 1024
rect 502 1019 508 1020
rect 502 1015 503 1019
rect 507 1015 508 1019
rect 542 1019 543 1023
rect 547 1019 548 1023
rect 542 1018 548 1019
rect 502 1014 508 1015
rect 530 991 536 992
rect 494 987 500 988
rect 494 983 495 987
rect 499 983 500 987
rect 530 987 531 991
rect 535 987 536 991
rect 530 986 536 987
rect 494 982 500 983
rect 502 972 508 973
rect 502 968 503 972
rect 507 968 508 972
rect 502 967 508 968
rect 504 955 506 967
rect 463 954 467 955
rect 463 949 467 950
rect 503 954 507 955
rect 503 949 507 950
rect 414 943 420 944
rect 414 939 415 943
rect 419 939 420 943
rect 414 938 420 939
rect 398 928 404 929
rect 398 924 399 928
rect 403 924 404 928
rect 398 923 404 924
rect 464 921 466 949
rect 462 920 468 921
rect 462 916 463 920
rect 467 916 468 920
rect 386 915 392 916
rect 462 915 468 916
rect 386 911 387 915
rect 391 911 392 915
rect 386 910 392 911
rect 388 872 390 910
rect 426 907 432 908
rect 426 903 427 907
rect 431 903 432 907
rect 426 902 432 903
rect 434 905 440 906
rect 398 881 404 882
rect 398 877 399 881
rect 403 877 404 881
rect 398 876 404 877
rect 386 871 392 872
rect 386 867 387 871
rect 391 867 392 871
rect 386 866 392 867
rect 358 839 364 840
rect 400 839 402 876
rect 414 875 420 876
rect 414 871 415 875
rect 419 871 420 875
rect 414 870 420 871
rect 416 856 418 870
rect 428 864 430 902
rect 434 901 435 905
rect 439 901 440 905
rect 434 900 440 901
rect 426 863 432 864
rect 426 859 427 863
rect 431 859 432 863
rect 426 858 432 859
rect 414 855 420 856
rect 414 851 415 855
rect 419 851 420 855
rect 414 850 420 851
rect 358 835 359 839
rect 363 835 364 839
rect 358 834 364 835
rect 399 838 403 839
rect 399 833 403 834
rect 407 838 411 839
rect 407 833 411 834
rect 408 824 410 833
rect 406 823 412 824
rect 406 819 407 823
rect 411 819 412 823
rect 406 818 412 819
rect 406 782 412 783
rect 406 778 407 782
rect 411 778 412 782
rect 406 777 412 778
rect 408 755 410 777
rect 391 754 395 755
rect 391 749 395 750
rect 407 754 411 755
rect 407 749 411 750
rect 392 733 394 749
rect 390 732 396 733
rect 390 728 391 732
rect 395 728 396 732
rect 390 727 396 728
rect 416 723 418 850
rect 436 839 438 900
rect 522 895 528 896
rect 522 891 523 895
rect 527 891 528 895
rect 522 890 528 891
rect 435 838 439 839
rect 435 833 439 834
rect 426 831 432 832
rect 426 827 427 831
rect 431 827 432 831
rect 426 826 432 827
rect 412 721 418 723
rect 390 685 396 686
rect 390 681 391 685
rect 395 681 396 685
rect 390 680 396 681
rect 412 680 414 721
rect 418 711 424 712
rect 418 707 419 711
rect 423 707 424 711
rect 418 706 424 707
rect 392 643 394 680
rect 410 679 416 680
rect 398 675 404 676
rect 398 671 399 675
rect 403 671 404 675
rect 410 675 411 679
rect 415 675 416 679
rect 410 674 416 675
rect 398 670 404 671
rect 391 642 395 643
rect 338 639 344 640
rect 338 635 339 639
rect 343 635 344 639
rect 391 637 395 638
rect 338 634 344 635
rect 400 596 402 670
rect 412 668 414 674
rect 420 668 422 706
rect 428 684 430 826
rect 471 754 475 755
rect 471 749 475 750
rect 472 725 474 749
rect 470 724 476 725
rect 470 720 471 724
rect 475 720 476 724
rect 470 719 476 720
rect 442 709 448 710
rect 442 705 443 709
rect 447 705 448 709
rect 442 704 448 705
rect 426 683 432 684
rect 426 679 427 683
rect 431 679 432 683
rect 426 678 432 679
rect 410 667 416 668
rect 410 663 411 667
rect 415 663 416 667
rect 410 662 416 663
rect 418 667 424 668
rect 418 663 419 667
rect 423 663 424 667
rect 418 662 424 663
rect 444 643 446 704
rect 524 676 526 890
rect 532 856 534 986
rect 544 880 546 1018
rect 576 1008 578 1266
rect 584 1263 586 1297
rect 616 1263 618 1297
rect 583 1262 587 1263
rect 583 1257 587 1258
rect 615 1262 619 1263
rect 615 1257 619 1258
rect 584 1195 586 1257
rect 606 1255 612 1256
rect 606 1251 607 1255
rect 611 1251 612 1255
rect 606 1250 612 1251
rect 590 1215 596 1216
rect 590 1211 591 1215
rect 595 1211 596 1215
rect 590 1210 596 1211
rect 592 1200 594 1210
rect 598 1207 604 1208
rect 598 1203 599 1207
rect 603 1203 604 1207
rect 598 1202 604 1203
rect 590 1199 596 1200
rect 590 1195 591 1199
rect 595 1195 596 1199
rect 582 1194 588 1195
rect 590 1194 596 1195
rect 582 1190 583 1194
rect 587 1190 588 1194
rect 582 1189 588 1190
rect 600 1184 602 1202
rect 598 1183 604 1184
rect 598 1179 599 1183
rect 603 1179 604 1183
rect 598 1178 604 1179
rect 582 1177 588 1178
rect 582 1173 583 1177
rect 587 1173 588 1177
rect 582 1172 588 1173
rect 584 1151 586 1172
rect 583 1150 587 1151
rect 583 1145 587 1146
rect 584 1125 586 1145
rect 582 1124 588 1125
rect 582 1120 583 1124
rect 587 1120 588 1124
rect 582 1119 588 1120
rect 590 1086 596 1087
rect 590 1082 591 1086
rect 595 1082 596 1086
rect 590 1081 596 1082
rect 592 1035 594 1081
rect 598 1075 604 1076
rect 598 1071 599 1075
rect 603 1074 604 1075
rect 608 1074 610 1250
rect 616 1195 618 1257
rect 628 1216 630 1306
rect 646 1302 652 1303
rect 646 1298 647 1302
rect 651 1298 652 1302
rect 646 1297 652 1298
rect 648 1263 650 1297
rect 664 1296 666 1374
rect 662 1295 668 1296
rect 662 1291 663 1295
rect 667 1291 668 1295
rect 662 1290 668 1291
rect 647 1262 651 1263
rect 647 1257 651 1258
rect 626 1215 632 1216
rect 626 1211 627 1215
rect 631 1211 632 1215
rect 626 1210 632 1211
rect 648 1195 650 1257
rect 654 1227 660 1228
rect 654 1223 655 1227
rect 659 1223 660 1227
rect 654 1222 660 1223
rect 614 1194 620 1195
rect 614 1190 615 1194
rect 619 1190 620 1194
rect 614 1189 620 1190
rect 646 1194 652 1195
rect 646 1190 647 1194
rect 651 1190 652 1194
rect 646 1189 652 1190
rect 614 1177 620 1178
rect 614 1173 615 1177
rect 619 1173 620 1177
rect 614 1172 620 1173
rect 646 1177 652 1178
rect 646 1173 647 1177
rect 651 1173 652 1177
rect 646 1172 652 1173
rect 616 1151 618 1172
rect 648 1151 650 1172
rect 615 1150 619 1151
rect 615 1145 619 1146
rect 647 1150 651 1151
rect 647 1145 651 1146
rect 656 1116 658 1222
rect 654 1115 660 1116
rect 654 1111 655 1115
rect 659 1111 660 1115
rect 654 1110 660 1111
rect 658 1105 664 1106
rect 658 1101 659 1105
rect 663 1101 664 1105
rect 658 1100 664 1101
rect 603 1072 610 1074
rect 603 1071 604 1072
rect 598 1070 604 1071
rect 583 1034 587 1035
rect 583 1029 587 1030
rect 591 1034 595 1035
rect 591 1029 595 1030
rect 584 1016 586 1029
rect 582 1015 588 1016
rect 582 1011 583 1015
rect 587 1011 588 1015
rect 582 1010 588 1011
rect 574 1007 580 1008
rect 574 1003 575 1007
rect 579 1003 580 1007
rect 574 1002 580 1003
rect 582 974 588 975
rect 582 970 583 974
rect 587 970 588 974
rect 582 969 588 970
rect 584 955 586 969
rect 600 956 602 1070
rect 606 1067 612 1068
rect 606 1063 607 1067
rect 611 1063 612 1067
rect 606 1062 612 1063
rect 598 955 604 956
rect 583 954 587 955
rect 583 949 587 950
rect 591 954 595 955
rect 598 951 599 955
rect 603 951 604 955
rect 598 950 604 951
rect 591 949 595 950
rect 592 927 594 949
rect 590 926 596 927
rect 590 922 591 926
rect 595 922 596 926
rect 590 921 596 922
rect 598 919 604 920
rect 598 915 599 919
rect 603 915 604 919
rect 598 914 604 915
rect 590 885 596 886
rect 590 881 591 885
rect 595 881 596 885
rect 590 880 596 881
rect 542 879 548 880
rect 542 875 543 879
rect 547 875 548 879
rect 542 874 548 875
rect 530 855 536 856
rect 530 851 531 855
rect 535 851 536 855
rect 530 850 536 851
rect 592 839 594 880
rect 600 860 602 914
rect 608 896 610 1062
rect 660 1035 662 1100
rect 672 1093 674 1422
rect 680 1391 682 1425
rect 678 1390 684 1391
rect 678 1386 679 1390
rect 683 1386 684 1390
rect 678 1385 684 1386
rect 678 1373 684 1374
rect 678 1369 679 1373
rect 683 1369 684 1373
rect 678 1368 684 1369
rect 680 1351 682 1368
rect 688 1360 690 1451
rect 704 1431 706 1453
rect 720 1452 722 1510
rect 743 1498 747 1499
rect 743 1493 747 1494
rect 744 1476 746 1493
rect 742 1475 748 1476
rect 742 1471 743 1475
rect 747 1471 748 1475
rect 742 1470 748 1471
rect 742 1458 748 1459
rect 742 1454 743 1458
rect 747 1454 748 1458
rect 742 1453 748 1454
rect 718 1451 724 1452
rect 718 1447 719 1451
rect 723 1447 724 1451
rect 718 1446 724 1447
rect 744 1431 746 1453
rect 703 1430 707 1431
rect 703 1425 707 1426
rect 719 1430 723 1431
rect 719 1425 723 1426
rect 743 1430 747 1431
rect 743 1425 747 1426
rect 694 1395 700 1396
rect 694 1391 695 1395
rect 699 1391 700 1395
rect 720 1394 722 1425
rect 750 1423 756 1424
rect 750 1419 751 1423
rect 755 1419 756 1423
rect 750 1418 756 1419
rect 694 1390 700 1391
rect 718 1393 724 1394
rect 686 1359 692 1360
rect 686 1355 687 1359
rect 691 1355 692 1359
rect 686 1354 692 1355
rect 679 1350 683 1351
rect 679 1345 683 1346
rect 680 1320 682 1345
rect 678 1319 684 1320
rect 678 1315 679 1319
rect 683 1315 684 1319
rect 678 1314 684 1315
rect 696 1312 698 1390
rect 718 1389 719 1393
rect 723 1389 724 1393
rect 718 1388 724 1389
rect 734 1366 740 1367
rect 734 1362 735 1366
rect 739 1362 740 1366
rect 734 1361 740 1362
rect 736 1351 738 1361
rect 711 1350 715 1351
rect 711 1345 715 1346
rect 735 1350 739 1351
rect 735 1345 739 1346
rect 743 1350 747 1351
rect 743 1345 747 1346
rect 712 1320 714 1345
rect 744 1321 746 1345
rect 742 1320 748 1321
rect 710 1319 716 1320
rect 710 1315 711 1319
rect 715 1315 716 1319
rect 742 1316 743 1320
rect 747 1316 748 1320
rect 742 1315 748 1316
rect 710 1314 716 1315
rect 694 1311 700 1312
rect 694 1307 695 1311
rect 699 1307 700 1311
rect 752 1308 754 1418
rect 760 1408 762 1546
rect 856 1543 858 1553
rect 775 1542 779 1543
rect 775 1537 779 1538
rect 855 1542 859 1543
rect 855 1537 859 1538
rect 871 1542 875 1543
rect 871 1537 875 1538
rect 776 1527 778 1537
rect 872 1527 874 1537
rect 774 1526 780 1527
rect 774 1522 775 1526
rect 779 1522 780 1526
rect 774 1521 780 1522
rect 870 1526 876 1527
rect 870 1522 871 1526
rect 875 1522 876 1526
rect 870 1521 876 1522
rect 774 1509 780 1510
rect 774 1505 775 1509
rect 779 1505 780 1509
rect 774 1504 780 1505
rect 870 1509 876 1510
rect 870 1505 871 1509
rect 875 1505 876 1509
rect 870 1504 876 1505
rect 776 1499 778 1504
rect 872 1499 874 1504
rect 775 1498 779 1499
rect 775 1493 779 1494
rect 807 1498 811 1499
rect 807 1493 811 1494
rect 871 1498 875 1499
rect 871 1493 875 1494
rect 776 1476 778 1493
rect 808 1477 810 1493
rect 806 1476 812 1477
rect 774 1475 780 1476
rect 774 1471 775 1475
rect 779 1471 780 1475
rect 806 1472 807 1476
rect 811 1472 812 1476
rect 806 1471 812 1472
rect 774 1470 780 1471
rect 774 1457 780 1458
rect 774 1453 775 1457
rect 779 1453 780 1457
rect 774 1452 780 1453
rect 806 1457 812 1458
rect 806 1453 807 1457
rect 811 1453 812 1457
rect 806 1452 812 1453
rect 776 1431 778 1452
rect 808 1431 810 1452
rect 814 1443 820 1444
rect 814 1439 815 1443
rect 819 1439 820 1443
rect 814 1438 820 1439
rect 767 1430 771 1431
rect 767 1425 771 1426
rect 775 1430 779 1431
rect 775 1425 779 1426
rect 807 1430 811 1431
rect 807 1425 811 1426
rect 768 1416 770 1425
rect 794 1423 800 1424
rect 794 1419 795 1423
rect 799 1419 800 1423
rect 794 1418 800 1419
rect 766 1415 772 1416
rect 766 1411 767 1415
rect 771 1411 772 1415
rect 766 1410 772 1411
rect 758 1407 764 1408
rect 758 1403 759 1407
rect 763 1403 764 1407
rect 758 1402 764 1403
rect 762 1395 768 1396
rect 762 1394 763 1395
rect 760 1391 763 1394
rect 767 1391 768 1395
rect 760 1390 768 1391
rect 694 1306 700 1307
rect 750 1307 756 1308
rect 750 1303 751 1307
rect 755 1303 756 1307
rect 678 1302 684 1303
rect 678 1298 679 1302
rect 683 1298 684 1302
rect 678 1297 684 1298
rect 710 1302 716 1303
rect 750 1302 756 1303
rect 710 1298 711 1302
rect 715 1298 716 1302
rect 710 1297 716 1298
rect 680 1263 682 1297
rect 712 1263 714 1297
rect 750 1282 756 1283
rect 734 1279 740 1280
rect 734 1275 735 1279
rect 739 1275 740 1279
rect 750 1278 751 1282
rect 755 1278 756 1282
rect 750 1277 756 1278
rect 734 1274 740 1275
rect 736 1264 738 1274
rect 734 1263 740 1264
rect 752 1263 754 1277
rect 760 1272 762 1390
rect 786 1387 792 1388
rect 786 1383 787 1387
rect 791 1383 792 1387
rect 786 1382 792 1383
rect 766 1368 772 1369
rect 766 1364 767 1368
rect 771 1364 772 1368
rect 766 1363 772 1364
rect 768 1351 770 1363
rect 767 1350 771 1351
rect 767 1345 771 1346
rect 788 1272 790 1382
rect 758 1271 764 1272
rect 758 1267 759 1271
rect 763 1267 764 1271
rect 758 1266 764 1267
rect 786 1271 792 1272
rect 786 1267 787 1271
rect 791 1267 792 1271
rect 786 1266 792 1267
rect 679 1262 683 1263
rect 679 1257 683 1258
rect 711 1262 715 1263
rect 734 1259 735 1263
rect 739 1259 740 1263
rect 734 1258 740 1259
rect 743 1262 747 1263
rect 711 1257 715 1258
rect 743 1257 747 1258
rect 751 1262 755 1263
rect 751 1257 755 1258
rect 680 1195 682 1257
rect 712 1195 714 1257
rect 744 1195 746 1257
rect 760 1256 762 1266
rect 775 1262 779 1263
rect 775 1257 779 1258
rect 758 1255 764 1256
rect 758 1251 759 1255
rect 763 1251 764 1255
rect 758 1250 764 1251
rect 776 1220 778 1257
rect 796 1224 798 1418
rect 808 1396 810 1425
rect 806 1395 812 1396
rect 806 1391 807 1395
rect 811 1391 812 1395
rect 806 1390 812 1391
rect 806 1372 812 1373
rect 806 1368 807 1372
rect 811 1368 812 1372
rect 806 1367 812 1368
rect 808 1351 810 1367
rect 816 1356 818 1438
rect 839 1430 843 1431
rect 839 1425 843 1426
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 814 1355 820 1356
rect 814 1351 815 1355
rect 819 1351 820 1355
rect 807 1350 811 1351
rect 814 1350 820 1351
rect 823 1350 827 1351
rect 807 1345 811 1346
rect 823 1345 827 1346
rect 824 1321 826 1345
rect 822 1320 828 1321
rect 822 1316 823 1320
rect 827 1316 828 1320
rect 822 1315 828 1316
rect 832 1308 834 1418
rect 840 1416 842 1425
rect 880 1420 882 1609
rect 974 1607 975 1611
rect 979 1607 980 1611
rect 1000 1607 1002 1617
rect 974 1606 980 1607
rect 998 1606 1004 1607
rect 959 1582 963 1583
rect 959 1576 963 1578
rect 958 1575 964 1576
rect 958 1571 959 1575
rect 963 1571 964 1575
rect 958 1570 964 1571
rect 976 1568 978 1606
rect 998 1602 999 1606
rect 1003 1602 1004 1606
rect 998 1601 1004 1602
rect 1020 1596 1022 1634
rect 1040 1623 1042 1641
rect 1184 1623 1186 1641
rect 1039 1622 1043 1623
rect 1039 1617 1043 1618
rect 1127 1622 1131 1623
rect 1127 1617 1131 1618
rect 1183 1622 1187 1623
rect 1183 1617 1187 1618
rect 1078 1611 1084 1612
rect 1078 1607 1079 1611
rect 1083 1607 1084 1611
rect 1128 1607 1130 1617
rect 1174 1611 1180 1612
rect 1174 1607 1175 1611
rect 1179 1607 1180 1611
rect 1078 1606 1084 1607
rect 1126 1606 1132 1607
rect 1174 1606 1180 1607
rect 1018 1595 1024 1596
rect 1018 1591 1019 1595
rect 1023 1591 1024 1595
rect 1018 1590 1024 1591
rect 998 1589 1004 1590
rect 998 1585 999 1589
rect 1003 1585 1004 1589
rect 998 1584 1004 1585
rect 999 1582 1003 1584
rect 999 1577 1003 1578
rect 1063 1582 1067 1583
rect 1063 1576 1067 1578
rect 1062 1575 1068 1576
rect 1062 1571 1063 1575
rect 1067 1571 1068 1575
rect 1062 1570 1068 1571
rect 1080 1568 1082 1606
rect 1126 1602 1127 1606
rect 1131 1602 1132 1606
rect 1126 1601 1132 1602
rect 1126 1589 1132 1590
rect 1126 1585 1127 1589
rect 1131 1585 1132 1589
rect 1126 1584 1132 1585
rect 1127 1582 1131 1584
rect 1127 1577 1131 1578
rect 1159 1582 1163 1583
rect 1159 1576 1163 1578
rect 1158 1575 1164 1576
rect 1158 1571 1159 1575
rect 1163 1571 1164 1575
rect 1158 1570 1164 1571
rect 1176 1568 1178 1606
rect 974 1567 980 1568
rect 974 1563 975 1567
rect 979 1563 980 1567
rect 974 1562 980 1563
rect 1078 1567 1084 1568
rect 1078 1563 1079 1567
rect 1083 1563 1084 1567
rect 1078 1562 1084 1563
rect 1174 1567 1180 1568
rect 1174 1563 1175 1567
rect 1179 1563 1180 1567
rect 1192 1563 1194 1754
rect 1694 1753 1700 1754
rect 1694 1749 1695 1753
rect 1699 1749 1700 1753
rect 1694 1748 1700 1749
rect 1694 1736 1700 1737
rect 1694 1732 1695 1736
rect 1699 1732 1700 1736
rect 1694 1731 1700 1732
rect 1696 1719 1698 1731
rect 1255 1718 1259 1719
rect 1255 1713 1259 1714
rect 1335 1718 1339 1719
rect 1335 1713 1339 1714
rect 1407 1718 1411 1719
rect 1407 1713 1411 1714
rect 1463 1718 1467 1719
rect 1463 1713 1467 1714
rect 1519 1718 1523 1719
rect 1519 1713 1523 1714
rect 1567 1718 1571 1719
rect 1567 1713 1571 1714
rect 1623 1718 1627 1719
rect 1623 1713 1627 1714
rect 1655 1718 1659 1719
rect 1655 1713 1659 1714
rect 1695 1718 1699 1719
rect 1695 1713 1699 1714
rect 1206 1711 1212 1712
rect 1198 1707 1204 1708
rect 1198 1703 1199 1707
rect 1203 1703 1204 1707
rect 1206 1707 1207 1711
rect 1211 1707 1212 1711
rect 1206 1706 1212 1707
rect 1198 1702 1204 1703
rect 1200 1656 1202 1702
rect 1208 1692 1210 1706
rect 1256 1703 1258 1713
rect 1336 1703 1338 1713
rect 1408 1703 1410 1713
rect 1464 1703 1466 1713
rect 1520 1703 1522 1713
rect 1568 1703 1570 1713
rect 1624 1703 1626 1713
rect 1656 1703 1658 1713
rect 1696 1705 1698 1713
rect 1694 1704 1700 1705
rect 1254 1702 1260 1703
rect 1254 1698 1255 1702
rect 1259 1698 1260 1702
rect 1254 1697 1260 1698
rect 1334 1702 1340 1703
rect 1334 1698 1335 1702
rect 1339 1698 1340 1702
rect 1334 1697 1340 1698
rect 1406 1702 1412 1703
rect 1406 1698 1407 1702
rect 1411 1698 1412 1702
rect 1406 1697 1412 1698
rect 1462 1702 1468 1703
rect 1462 1698 1463 1702
rect 1467 1698 1468 1702
rect 1462 1697 1468 1698
rect 1518 1702 1524 1703
rect 1518 1698 1519 1702
rect 1523 1698 1524 1702
rect 1518 1697 1524 1698
rect 1566 1702 1572 1703
rect 1566 1698 1567 1702
rect 1571 1698 1572 1702
rect 1566 1697 1572 1698
rect 1622 1702 1628 1703
rect 1622 1698 1623 1702
rect 1627 1698 1628 1702
rect 1622 1697 1628 1698
rect 1654 1702 1660 1703
rect 1654 1698 1655 1702
rect 1659 1698 1660 1702
rect 1694 1700 1695 1704
rect 1699 1700 1700 1704
rect 1694 1699 1700 1700
rect 1654 1697 1660 1698
rect 1206 1691 1212 1692
rect 1206 1687 1207 1691
rect 1211 1687 1212 1691
rect 1206 1686 1212 1687
rect 1694 1687 1700 1688
rect 1254 1685 1260 1686
rect 1254 1681 1255 1685
rect 1259 1681 1260 1685
rect 1254 1680 1260 1681
rect 1334 1685 1340 1686
rect 1334 1681 1335 1685
rect 1339 1681 1340 1685
rect 1334 1680 1340 1681
rect 1406 1685 1412 1686
rect 1406 1681 1407 1685
rect 1411 1681 1412 1685
rect 1406 1680 1412 1681
rect 1462 1685 1468 1686
rect 1462 1681 1463 1685
rect 1467 1681 1468 1685
rect 1462 1680 1468 1681
rect 1518 1685 1524 1686
rect 1518 1681 1519 1685
rect 1523 1681 1524 1685
rect 1518 1680 1524 1681
rect 1566 1685 1572 1686
rect 1566 1681 1567 1685
rect 1571 1681 1572 1685
rect 1566 1680 1572 1681
rect 1622 1685 1628 1686
rect 1622 1681 1623 1685
rect 1627 1681 1628 1685
rect 1622 1680 1628 1681
rect 1654 1685 1660 1686
rect 1654 1681 1655 1685
rect 1659 1681 1660 1685
rect 1694 1683 1695 1687
rect 1699 1683 1700 1687
rect 1694 1682 1700 1683
rect 1654 1680 1660 1681
rect 1256 1671 1258 1680
rect 1336 1671 1338 1680
rect 1408 1671 1410 1680
rect 1464 1671 1466 1680
rect 1470 1679 1476 1680
rect 1470 1675 1471 1679
rect 1475 1675 1476 1679
rect 1470 1674 1476 1675
rect 1255 1670 1259 1671
rect 1255 1665 1259 1666
rect 1319 1670 1323 1671
rect 1319 1664 1323 1666
rect 1335 1670 1339 1671
rect 1335 1665 1339 1666
rect 1407 1670 1411 1671
rect 1407 1665 1411 1666
rect 1439 1670 1443 1671
rect 1439 1664 1443 1666
rect 1463 1670 1467 1671
rect 1463 1665 1467 1666
rect 1318 1663 1324 1664
rect 1318 1659 1319 1663
rect 1323 1659 1324 1663
rect 1318 1658 1324 1659
rect 1438 1663 1444 1664
rect 1438 1659 1439 1663
rect 1443 1659 1444 1663
rect 1438 1658 1444 1659
rect 1198 1655 1204 1656
rect 1198 1651 1199 1655
rect 1203 1651 1204 1655
rect 1198 1650 1204 1651
rect 1318 1646 1324 1647
rect 1318 1642 1319 1646
rect 1323 1642 1324 1646
rect 1318 1641 1324 1642
rect 1438 1646 1444 1647
rect 1438 1642 1439 1646
rect 1443 1642 1444 1646
rect 1438 1641 1444 1642
rect 1320 1623 1322 1641
rect 1374 1639 1380 1640
rect 1374 1635 1375 1639
rect 1379 1635 1380 1639
rect 1374 1634 1380 1635
rect 1247 1622 1251 1623
rect 1247 1617 1251 1618
rect 1319 1622 1323 1623
rect 1319 1617 1323 1618
rect 1359 1622 1363 1623
rect 1359 1617 1363 1618
rect 1210 1615 1216 1616
rect 1210 1611 1211 1615
rect 1215 1611 1216 1615
rect 1210 1610 1216 1611
rect 1212 1596 1214 1610
rect 1248 1607 1250 1617
rect 1360 1607 1362 1617
rect 1246 1606 1252 1607
rect 1246 1602 1247 1606
rect 1251 1602 1252 1606
rect 1246 1601 1252 1602
rect 1358 1606 1364 1607
rect 1358 1602 1359 1606
rect 1363 1602 1364 1606
rect 1358 1601 1364 1602
rect 1376 1596 1378 1634
rect 1440 1623 1442 1641
rect 1472 1640 1474 1674
rect 1520 1671 1522 1680
rect 1568 1671 1570 1680
rect 1624 1671 1626 1680
rect 1656 1671 1658 1680
rect 1696 1671 1698 1682
rect 1519 1670 1523 1671
rect 1519 1665 1523 1666
rect 1559 1670 1563 1671
rect 1559 1664 1563 1666
rect 1567 1670 1571 1671
rect 1567 1665 1571 1666
rect 1623 1670 1627 1671
rect 1623 1665 1627 1666
rect 1655 1670 1659 1671
rect 1655 1664 1659 1666
rect 1695 1670 1699 1671
rect 1695 1665 1699 1666
rect 1558 1663 1564 1664
rect 1558 1659 1559 1663
rect 1563 1659 1564 1663
rect 1558 1658 1564 1659
rect 1654 1663 1660 1664
rect 1654 1659 1655 1663
rect 1659 1659 1660 1663
rect 1696 1662 1698 1665
rect 1654 1658 1660 1659
rect 1694 1661 1700 1662
rect 1694 1657 1695 1661
rect 1699 1657 1700 1661
rect 1694 1656 1700 1657
rect 1670 1655 1676 1656
rect 1670 1651 1671 1655
rect 1675 1651 1676 1655
rect 1670 1650 1676 1651
rect 1558 1646 1564 1647
rect 1558 1642 1559 1646
rect 1563 1642 1564 1646
rect 1558 1641 1564 1642
rect 1654 1646 1660 1647
rect 1654 1642 1655 1646
rect 1659 1642 1660 1646
rect 1654 1641 1660 1642
rect 1470 1639 1476 1640
rect 1470 1635 1471 1639
rect 1475 1635 1476 1639
rect 1470 1634 1476 1635
rect 1560 1623 1562 1641
rect 1656 1623 1658 1641
rect 1439 1622 1443 1623
rect 1439 1617 1443 1618
rect 1463 1622 1467 1623
rect 1463 1617 1467 1618
rect 1559 1622 1563 1623
rect 1559 1617 1563 1618
rect 1567 1622 1571 1623
rect 1567 1617 1571 1618
rect 1655 1622 1659 1623
rect 1655 1617 1659 1618
rect 1464 1607 1466 1617
rect 1478 1611 1484 1612
rect 1478 1607 1479 1611
rect 1483 1607 1484 1611
rect 1568 1607 1570 1617
rect 1656 1607 1658 1617
rect 1672 1612 1674 1650
rect 1694 1644 1700 1645
rect 1694 1640 1695 1644
rect 1699 1640 1700 1644
rect 1694 1639 1700 1640
rect 1696 1623 1698 1639
rect 1695 1622 1699 1623
rect 1695 1617 1699 1618
rect 1670 1611 1676 1612
rect 1670 1607 1671 1611
rect 1675 1607 1676 1611
rect 1696 1609 1698 1617
rect 1462 1606 1468 1607
rect 1478 1606 1484 1607
rect 1566 1606 1572 1607
rect 1462 1602 1463 1606
rect 1467 1602 1468 1606
rect 1462 1601 1468 1602
rect 1210 1595 1216 1596
rect 1210 1591 1211 1595
rect 1215 1591 1216 1595
rect 1210 1590 1216 1591
rect 1342 1595 1348 1596
rect 1342 1591 1343 1595
rect 1347 1591 1348 1595
rect 1342 1590 1348 1591
rect 1374 1595 1380 1596
rect 1374 1591 1375 1595
rect 1379 1591 1380 1595
rect 1374 1590 1380 1591
rect 1246 1589 1252 1590
rect 1246 1585 1247 1589
rect 1251 1585 1252 1589
rect 1246 1584 1252 1585
rect 1247 1582 1251 1584
rect 1247 1576 1251 1578
rect 1327 1582 1331 1583
rect 1327 1576 1331 1578
rect 1246 1575 1252 1576
rect 1246 1571 1247 1575
rect 1251 1571 1252 1575
rect 1246 1570 1252 1571
rect 1326 1575 1332 1576
rect 1326 1571 1327 1575
rect 1331 1571 1332 1575
rect 1326 1570 1332 1571
rect 1174 1562 1180 1563
rect 1188 1561 1194 1563
rect 958 1558 964 1559
rect 958 1554 959 1558
rect 963 1554 964 1558
rect 958 1553 964 1554
rect 1062 1558 1068 1559
rect 1062 1554 1063 1558
rect 1067 1554 1068 1558
rect 1062 1553 1068 1554
rect 1158 1558 1164 1559
rect 1158 1554 1159 1558
rect 1163 1554 1164 1558
rect 1158 1553 1164 1554
rect 960 1543 962 1553
rect 1030 1543 1036 1544
rect 1064 1543 1066 1553
rect 1102 1551 1108 1552
rect 1102 1547 1103 1551
rect 1107 1547 1108 1551
rect 1102 1546 1108 1547
rect 959 1542 963 1543
rect 959 1537 963 1538
rect 975 1542 979 1543
rect 1030 1539 1031 1543
rect 1035 1539 1036 1543
rect 1030 1538 1036 1539
rect 1063 1542 1067 1543
rect 975 1537 979 1538
rect 976 1527 978 1537
rect 974 1526 980 1527
rect 974 1522 975 1526
rect 979 1522 980 1526
rect 974 1521 980 1522
rect 990 1515 996 1516
rect 990 1511 991 1515
rect 995 1511 996 1515
rect 990 1510 996 1511
rect 974 1509 980 1510
rect 974 1505 975 1509
rect 979 1505 980 1509
rect 974 1504 980 1505
rect 976 1499 978 1504
rect 895 1498 899 1499
rect 895 1493 899 1494
rect 935 1498 939 1499
rect 935 1493 939 1494
rect 975 1498 979 1499
rect 975 1493 979 1494
rect 896 1477 898 1493
rect 918 1491 924 1492
rect 918 1487 919 1491
rect 923 1487 924 1491
rect 918 1486 924 1487
rect 894 1476 900 1477
rect 894 1472 895 1476
rect 899 1472 900 1476
rect 894 1471 900 1472
rect 886 1467 892 1468
rect 886 1463 887 1467
rect 891 1463 892 1467
rect 886 1462 892 1463
rect 888 1444 890 1462
rect 920 1460 922 1486
rect 936 1477 938 1493
rect 934 1476 940 1477
rect 934 1472 935 1476
rect 939 1472 940 1476
rect 934 1471 940 1472
rect 918 1459 924 1460
rect 918 1455 919 1459
rect 923 1455 924 1459
rect 918 1454 924 1455
rect 934 1457 940 1458
rect 934 1453 935 1457
rect 939 1453 940 1457
rect 934 1452 940 1453
rect 894 1448 900 1449
rect 894 1444 895 1448
rect 899 1444 900 1448
rect 886 1443 892 1444
rect 894 1443 900 1444
rect 886 1439 887 1443
rect 891 1439 892 1443
rect 886 1438 892 1439
rect 896 1431 898 1443
rect 910 1435 916 1436
rect 910 1431 911 1435
rect 915 1431 916 1435
rect 936 1431 938 1452
rect 992 1432 994 1510
rect 1023 1498 1027 1499
rect 1023 1493 1027 1494
rect 1024 1477 1026 1493
rect 1022 1476 1028 1477
rect 1022 1472 1023 1476
rect 1027 1472 1028 1476
rect 1022 1471 1028 1472
rect 1032 1436 1034 1538
rect 1063 1537 1067 1538
rect 1079 1542 1083 1543
rect 1079 1537 1083 1538
rect 1080 1527 1082 1537
rect 1094 1531 1100 1532
rect 1094 1527 1095 1531
rect 1099 1527 1100 1531
rect 1078 1526 1084 1527
rect 1094 1526 1100 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1078 1509 1084 1510
rect 1078 1505 1079 1509
rect 1083 1505 1084 1509
rect 1078 1504 1084 1505
rect 1080 1499 1082 1504
rect 1079 1498 1083 1499
rect 1079 1493 1083 1494
rect 1080 1476 1082 1493
rect 1078 1475 1084 1476
rect 1078 1471 1079 1475
rect 1083 1471 1084 1475
rect 1078 1470 1084 1471
rect 1096 1468 1098 1526
rect 1104 1524 1106 1546
rect 1160 1543 1162 1553
rect 1159 1542 1163 1543
rect 1159 1537 1163 1538
rect 1175 1542 1179 1543
rect 1175 1537 1179 1538
rect 1176 1527 1178 1537
rect 1188 1532 1190 1561
rect 1246 1558 1252 1559
rect 1246 1554 1247 1558
rect 1251 1554 1252 1558
rect 1246 1553 1252 1554
rect 1326 1558 1332 1559
rect 1326 1554 1327 1558
rect 1331 1554 1332 1558
rect 1326 1553 1332 1554
rect 1194 1551 1200 1552
rect 1194 1547 1195 1551
rect 1199 1547 1200 1551
rect 1194 1546 1200 1547
rect 1186 1531 1192 1532
rect 1186 1527 1187 1531
rect 1191 1527 1192 1531
rect 1174 1526 1180 1527
rect 1186 1526 1192 1527
rect 1102 1523 1108 1524
rect 1102 1519 1103 1523
rect 1107 1519 1108 1523
rect 1174 1522 1175 1526
rect 1179 1522 1180 1526
rect 1174 1521 1180 1522
rect 1102 1518 1108 1519
rect 1196 1516 1198 1546
rect 1248 1543 1250 1553
rect 1328 1543 1330 1553
rect 1344 1552 1346 1590
rect 1358 1589 1364 1590
rect 1358 1585 1359 1589
rect 1363 1585 1364 1589
rect 1358 1584 1364 1585
rect 1462 1589 1468 1590
rect 1462 1585 1463 1589
rect 1467 1585 1468 1589
rect 1462 1584 1468 1585
rect 1359 1582 1363 1584
rect 1359 1577 1363 1578
rect 1399 1582 1403 1583
rect 1399 1576 1403 1578
rect 1463 1582 1467 1584
rect 1463 1577 1467 1578
rect 1471 1582 1475 1583
rect 1471 1576 1475 1578
rect 1398 1575 1404 1576
rect 1398 1571 1399 1575
rect 1403 1571 1404 1575
rect 1398 1570 1404 1571
rect 1470 1575 1476 1576
rect 1470 1571 1471 1575
rect 1475 1571 1476 1575
rect 1470 1570 1476 1571
rect 1374 1567 1380 1568
rect 1374 1563 1375 1567
rect 1379 1563 1380 1567
rect 1374 1562 1380 1563
rect 1342 1551 1348 1552
rect 1342 1547 1343 1551
rect 1347 1547 1348 1551
rect 1342 1546 1348 1547
rect 1247 1542 1251 1543
rect 1247 1537 1251 1538
rect 1271 1542 1275 1543
rect 1271 1537 1275 1538
rect 1327 1542 1331 1543
rect 1327 1537 1331 1538
rect 1359 1542 1363 1543
rect 1359 1537 1363 1538
rect 1254 1535 1260 1536
rect 1214 1531 1220 1532
rect 1214 1527 1215 1531
rect 1219 1527 1220 1531
rect 1254 1531 1255 1535
rect 1259 1531 1260 1535
rect 1254 1530 1260 1531
rect 1214 1526 1220 1527
rect 1194 1515 1200 1516
rect 1194 1511 1195 1515
rect 1199 1511 1200 1515
rect 1194 1510 1200 1511
rect 1174 1509 1180 1510
rect 1174 1505 1175 1509
rect 1179 1505 1180 1509
rect 1174 1504 1180 1505
rect 1176 1499 1178 1504
rect 1111 1498 1115 1499
rect 1111 1493 1115 1494
rect 1167 1498 1171 1499
rect 1167 1493 1171 1494
rect 1175 1498 1179 1499
rect 1175 1493 1179 1494
rect 1199 1498 1203 1499
rect 1199 1493 1203 1494
rect 1112 1477 1114 1493
rect 1146 1491 1152 1492
rect 1146 1487 1147 1491
rect 1151 1487 1152 1491
rect 1146 1486 1152 1487
rect 1110 1476 1116 1477
rect 1110 1472 1111 1476
rect 1115 1472 1116 1476
rect 1110 1471 1116 1472
rect 1094 1467 1100 1468
rect 1094 1463 1095 1467
rect 1099 1463 1100 1467
rect 1094 1462 1100 1463
rect 1078 1458 1084 1459
rect 1038 1455 1044 1456
rect 1038 1451 1039 1455
rect 1043 1451 1044 1455
rect 1078 1454 1079 1458
rect 1083 1454 1084 1458
rect 1148 1456 1150 1486
rect 1168 1476 1170 1493
rect 1200 1476 1202 1493
rect 1166 1475 1172 1476
rect 1166 1471 1167 1475
rect 1171 1471 1172 1475
rect 1166 1470 1172 1471
rect 1198 1475 1204 1476
rect 1198 1471 1199 1475
rect 1203 1471 1204 1475
rect 1198 1470 1204 1471
rect 1166 1458 1172 1459
rect 1078 1453 1084 1454
rect 1126 1455 1132 1456
rect 1038 1450 1044 1451
rect 1030 1435 1036 1436
rect 990 1431 996 1432
rect 895 1430 899 1431
rect 910 1430 916 1431
rect 935 1430 939 1431
rect 895 1425 899 1426
rect 878 1419 884 1420
rect 838 1415 844 1416
rect 838 1411 839 1415
rect 843 1411 844 1415
rect 878 1415 879 1419
rect 883 1415 884 1419
rect 878 1414 884 1415
rect 896 1411 898 1425
rect 912 1421 914 1430
rect 935 1425 939 1426
rect 975 1430 979 1431
rect 990 1427 991 1431
rect 995 1427 996 1431
rect 990 1426 996 1427
rect 998 1431 1004 1432
rect 1030 1431 1031 1435
rect 1035 1431 1036 1435
rect 1040 1431 1042 1450
rect 1046 1439 1052 1440
rect 1046 1435 1047 1439
rect 1051 1435 1052 1439
rect 1046 1434 1052 1435
rect 998 1427 999 1431
rect 1003 1427 1004 1431
rect 998 1426 1004 1427
rect 1023 1430 1027 1431
rect 1030 1430 1036 1431
rect 1039 1430 1043 1431
rect 975 1425 979 1426
rect 946 1423 952 1424
rect 911 1420 915 1421
rect 902 1419 908 1420
rect 902 1415 903 1419
rect 907 1415 908 1419
rect 911 1415 915 1416
rect 918 1419 924 1420
rect 918 1415 919 1419
rect 923 1415 924 1419
rect 946 1419 947 1423
rect 951 1419 952 1423
rect 946 1418 952 1419
rect 902 1414 908 1415
rect 918 1414 924 1415
rect 838 1410 844 1411
rect 894 1410 900 1411
rect 894 1406 895 1410
rect 899 1406 900 1410
rect 894 1405 900 1406
rect 904 1403 906 1414
rect 896 1401 906 1403
rect 866 1387 872 1388
rect 866 1383 867 1387
rect 871 1383 872 1387
rect 866 1382 872 1383
rect 846 1379 852 1380
rect 846 1375 847 1379
rect 851 1375 852 1379
rect 846 1374 852 1375
rect 838 1368 844 1369
rect 838 1364 839 1368
rect 843 1364 844 1368
rect 838 1363 844 1364
rect 840 1351 842 1363
rect 839 1350 843 1351
rect 839 1345 843 1346
rect 830 1307 836 1308
rect 830 1303 831 1307
rect 835 1303 836 1307
rect 830 1302 836 1303
rect 830 1282 836 1283
rect 830 1278 831 1282
rect 835 1278 836 1282
rect 830 1277 836 1278
rect 832 1263 834 1277
rect 838 1271 844 1272
rect 838 1267 839 1271
rect 843 1267 844 1271
rect 838 1266 844 1267
rect 811 1262 815 1263
rect 811 1257 815 1258
rect 831 1262 835 1263
rect 831 1257 835 1258
rect 794 1223 800 1224
rect 774 1219 780 1220
rect 774 1215 775 1219
rect 779 1215 780 1219
rect 794 1219 795 1223
rect 799 1222 800 1223
rect 799 1219 802 1222
rect 794 1218 802 1219
rect 774 1214 780 1215
rect 790 1215 796 1216
rect 758 1211 764 1212
rect 758 1207 759 1211
rect 763 1207 764 1211
rect 790 1211 791 1215
rect 795 1211 796 1215
rect 790 1210 796 1211
rect 758 1206 764 1207
rect 678 1194 684 1195
rect 678 1190 679 1194
rect 683 1190 684 1194
rect 678 1189 684 1190
rect 710 1194 716 1195
rect 710 1190 711 1194
rect 715 1190 716 1194
rect 710 1189 716 1190
rect 742 1194 748 1195
rect 742 1190 743 1194
rect 747 1190 748 1194
rect 742 1189 748 1190
rect 760 1184 762 1206
rect 792 1192 794 1210
rect 790 1191 796 1192
rect 790 1187 791 1191
rect 795 1187 796 1191
rect 790 1186 796 1187
rect 758 1183 764 1184
rect 758 1179 759 1183
rect 763 1179 764 1183
rect 758 1178 764 1179
rect 678 1177 684 1178
rect 678 1173 679 1177
rect 683 1173 684 1177
rect 678 1172 684 1173
rect 710 1177 716 1178
rect 710 1173 711 1177
rect 715 1173 716 1177
rect 710 1172 716 1173
rect 742 1177 748 1178
rect 742 1173 743 1177
rect 747 1173 748 1177
rect 742 1172 748 1173
rect 774 1172 780 1173
rect 680 1151 682 1172
rect 712 1151 714 1172
rect 744 1151 746 1172
rect 774 1168 775 1172
rect 779 1168 780 1172
rect 774 1167 780 1168
rect 776 1151 778 1167
rect 679 1150 683 1151
rect 679 1145 683 1146
rect 687 1150 691 1151
rect 687 1145 691 1146
rect 711 1150 715 1151
rect 711 1145 715 1146
rect 743 1150 747 1151
rect 743 1145 747 1146
rect 775 1150 779 1151
rect 775 1145 779 1146
rect 688 1121 690 1145
rect 686 1120 692 1121
rect 686 1116 687 1120
rect 691 1116 692 1120
rect 686 1115 692 1116
rect 782 1119 788 1120
rect 782 1115 783 1119
rect 787 1115 788 1119
rect 782 1114 788 1115
rect 702 1095 708 1096
rect 671 1092 675 1093
rect 702 1091 703 1095
rect 707 1091 708 1095
rect 702 1090 708 1091
rect 671 1087 675 1088
rect 659 1034 663 1035
rect 659 1029 663 1030
rect 614 1023 620 1024
rect 614 1019 615 1023
rect 619 1019 620 1023
rect 614 1018 620 1019
rect 658 1023 664 1024
rect 658 1019 659 1023
rect 663 1019 664 1023
rect 658 1018 664 1019
rect 606 895 612 896
rect 606 891 607 895
rect 611 891 612 895
rect 606 890 612 891
rect 607 875 613 876
rect 607 871 608 875
rect 612 874 613 875
rect 616 874 618 1018
rect 660 956 662 1018
rect 658 955 664 956
rect 658 951 659 955
rect 663 951 664 955
rect 658 950 664 951
rect 679 954 683 955
rect 679 949 683 950
rect 680 925 682 949
rect 678 924 684 925
rect 678 920 679 924
rect 683 920 684 924
rect 678 919 684 920
rect 694 919 700 920
rect 694 915 695 919
rect 699 915 700 919
rect 694 914 700 915
rect 678 901 684 902
rect 678 897 679 901
rect 683 897 684 901
rect 678 896 684 897
rect 612 872 618 874
rect 612 871 613 872
rect 607 870 613 871
rect 598 859 604 860
rect 598 855 599 859
rect 603 855 604 859
rect 598 854 604 855
rect 608 840 610 870
rect 606 839 612 840
rect 680 839 682 896
rect 559 838 563 839
rect 559 833 563 834
rect 591 838 595 839
rect 606 835 607 839
rect 611 835 612 839
rect 606 834 612 835
rect 663 838 667 839
rect 591 833 595 834
rect 663 833 667 834
rect 679 838 683 839
rect 679 833 683 834
rect 560 803 562 833
rect 574 831 580 832
rect 574 827 575 831
rect 579 827 580 831
rect 574 826 580 827
rect 558 802 564 803
rect 558 798 559 802
rect 563 798 564 802
rect 558 797 564 798
rect 576 792 578 826
rect 664 818 666 833
rect 696 828 698 914
rect 704 868 706 1090
rect 711 1034 715 1035
rect 711 1029 715 1030
rect 712 1016 714 1029
rect 784 1024 786 1114
rect 792 1080 794 1186
rect 800 1164 802 1218
rect 812 1196 814 1257
rect 840 1256 842 1266
rect 838 1255 844 1256
rect 838 1251 839 1255
rect 843 1251 844 1255
rect 838 1250 844 1251
rect 848 1228 850 1374
rect 868 1272 870 1382
rect 886 1372 892 1373
rect 886 1368 887 1372
rect 891 1368 892 1372
rect 886 1367 892 1368
rect 888 1351 890 1367
rect 887 1350 891 1351
rect 887 1345 891 1346
rect 896 1339 898 1401
rect 903 1350 907 1351
rect 903 1345 907 1346
rect 888 1337 898 1339
rect 866 1271 872 1272
rect 866 1267 867 1271
rect 871 1267 872 1271
rect 866 1266 872 1267
rect 888 1256 890 1337
rect 904 1321 906 1345
rect 902 1320 908 1321
rect 902 1316 903 1320
rect 907 1316 908 1320
rect 902 1315 908 1316
rect 910 1282 916 1283
rect 910 1278 911 1282
rect 915 1278 916 1282
rect 910 1277 916 1278
rect 894 1271 900 1272
rect 894 1267 895 1271
rect 899 1270 900 1271
rect 899 1267 902 1270
rect 894 1266 902 1267
rect 886 1255 892 1256
rect 886 1251 887 1255
rect 891 1251 892 1255
rect 886 1250 892 1251
rect 900 1236 902 1266
rect 912 1263 914 1277
rect 911 1262 915 1263
rect 911 1257 915 1258
rect 920 1248 922 1414
rect 948 1384 950 1418
rect 976 1416 978 1425
rect 991 1420 995 1421
rect 966 1415 972 1416
rect 966 1411 967 1415
rect 971 1411 972 1415
rect 966 1410 972 1411
rect 974 1415 980 1416
rect 974 1411 975 1415
rect 979 1411 980 1415
rect 990 1415 991 1420
rect 995 1415 996 1420
rect 990 1414 996 1415
rect 974 1410 980 1411
rect 968 1388 970 1410
rect 1000 1396 1002 1426
rect 1023 1425 1027 1426
rect 1039 1425 1043 1426
rect 998 1395 1004 1396
rect 998 1391 999 1395
rect 1003 1391 1004 1395
rect 1024 1391 1026 1425
rect 1048 1416 1050 1434
rect 1080 1431 1082 1453
rect 1126 1451 1127 1455
rect 1131 1451 1132 1455
rect 1126 1450 1132 1451
rect 1146 1455 1152 1456
rect 1146 1451 1147 1455
rect 1151 1451 1152 1455
rect 1166 1454 1167 1458
rect 1171 1454 1172 1458
rect 1166 1453 1172 1454
rect 1198 1458 1204 1459
rect 1198 1454 1199 1458
rect 1203 1454 1204 1458
rect 1198 1453 1204 1454
rect 1146 1450 1152 1451
rect 1128 1431 1130 1450
rect 1138 1447 1144 1448
rect 1138 1443 1139 1447
rect 1143 1443 1144 1447
rect 1138 1442 1144 1443
rect 1063 1430 1067 1431
rect 1063 1425 1067 1426
rect 1079 1430 1083 1431
rect 1079 1425 1083 1426
rect 1111 1430 1115 1431
rect 1111 1425 1115 1426
rect 1127 1430 1131 1431
rect 1127 1425 1131 1426
rect 1046 1415 1052 1416
rect 1046 1411 1047 1415
rect 1051 1411 1052 1415
rect 1046 1410 1052 1411
rect 998 1390 1004 1391
rect 1022 1390 1028 1391
rect 966 1387 972 1388
rect 946 1383 952 1384
rect 946 1379 947 1383
rect 951 1379 952 1383
rect 966 1383 967 1387
rect 971 1383 972 1387
rect 1022 1386 1023 1390
rect 1027 1386 1028 1390
rect 1022 1385 1028 1386
rect 966 1382 972 1383
rect 946 1378 952 1379
rect 1022 1373 1028 1374
rect 1022 1369 1023 1373
rect 1027 1369 1028 1373
rect 974 1368 980 1369
rect 1022 1368 1028 1369
rect 974 1364 975 1368
rect 979 1364 980 1368
rect 974 1363 980 1364
rect 950 1355 956 1356
rect 950 1351 951 1355
rect 955 1351 956 1355
rect 976 1351 978 1363
rect 1024 1351 1026 1368
rect 950 1350 956 1351
rect 975 1350 979 1351
rect 930 1271 936 1272
rect 930 1267 931 1271
rect 935 1267 936 1271
rect 930 1266 936 1267
rect 918 1247 924 1248
rect 918 1243 919 1247
rect 923 1243 924 1247
rect 918 1242 924 1243
rect 898 1235 904 1236
rect 898 1231 899 1235
rect 903 1231 904 1235
rect 898 1230 904 1231
rect 846 1227 852 1228
rect 846 1223 847 1227
rect 851 1223 852 1227
rect 846 1222 852 1223
rect 932 1211 934 1266
rect 916 1209 934 1211
rect 822 1203 828 1204
rect 822 1199 823 1203
rect 827 1199 828 1203
rect 822 1198 828 1199
rect 810 1195 816 1196
rect 810 1191 811 1195
rect 815 1191 816 1195
rect 810 1190 816 1191
rect 798 1163 804 1164
rect 798 1159 799 1163
rect 803 1159 804 1163
rect 798 1158 804 1159
rect 814 1163 820 1164
rect 814 1159 815 1163
rect 819 1159 820 1163
rect 814 1158 820 1159
rect 799 1150 803 1151
rect 799 1145 803 1146
rect 800 1125 802 1145
rect 798 1124 804 1125
rect 798 1120 799 1124
rect 803 1120 804 1124
rect 798 1119 804 1120
rect 798 1101 804 1102
rect 798 1097 799 1101
rect 803 1097 804 1101
rect 798 1096 804 1097
rect 790 1079 796 1080
rect 790 1075 791 1079
rect 795 1075 796 1079
rect 790 1074 796 1075
rect 800 1035 802 1096
rect 816 1061 818 1158
rect 824 1072 826 1198
rect 838 1180 844 1181
rect 838 1176 839 1180
rect 843 1176 844 1180
rect 838 1175 844 1176
rect 840 1151 842 1175
rect 839 1150 843 1151
rect 839 1145 843 1146
rect 847 1150 851 1151
rect 847 1145 851 1146
rect 848 1127 850 1145
rect 846 1126 852 1127
rect 846 1122 847 1126
rect 851 1122 852 1126
rect 846 1121 852 1122
rect 854 1119 860 1120
rect 854 1115 855 1119
rect 859 1115 860 1119
rect 854 1114 860 1115
rect 846 1085 852 1086
rect 846 1081 847 1085
rect 851 1081 852 1085
rect 846 1080 852 1081
rect 822 1071 828 1072
rect 822 1067 823 1071
rect 827 1067 828 1071
rect 822 1066 828 1067
rect 815 1060 819 1061
rect 815 1055 819 1056
rect 848 1035 850 1080
rect 799 1034 803 1035
rect 799 1029 803 1030
rect 823 1034 827 1035
rect 847 1034 851 1035
rect 823 1029 827 1030
rect 830 1031 836 1032
rect 782 1023 788 1024
rect 782 1019 783 1023
rect 787 1019 788 1023
rect 782 1018 788 1019
rect 710 1015 716 1016
rect 710 1011 711 1015
rect 715 1011 716 1015
rect 710 1010 716 1011
rect 824 1010 826 1029
rect 830 1027 831 1031
rect 835 1027 836 1031
rect 847 1029 851 1030
rect 830 1026 836 1027
rect 822 1009 828 1010
rect 822 1005 823 1009
rect 827 1005 828 1009
rect 822 1004 828 1005
rect 822 979 828 980
rect 822 975 823 979
rect 827 975 828 979
rect 710 974 716 975
rect 822 974 828 975
rect 710 970 711 974
rect 715 970 716 974
rect 710 969 716 970
rect 814 969 820 970
rect 712 955 714 969
rect 814 965 815 969
rect 819 965 820 969
rect 814 964 820 965
rect 816 955 818 964
rect 711 954 715 955
rect 711 949 715 950
rect 727 954 731 955
rect 727 949 731 950
rect 815 954 819 955
rect 815 949 819 950
rect 728 927 730 949
rect 726 926 732 927
rect 726 922 727 926
rect 731 922 732 926
rect 816 924 818 949
rect 726 921 732 922
rect 814 923 820 924
rect 814 919 815 923
rect 819 919 820 923
rect 814 918 820 919
rect 802 915 808 916
rect 802 911 803 915
rect 807 911 808 915
rect 802 910 808 911
rect 726 885 732 886
rect 726 881 727 885
rect 731 881 732 885
rect 726 880 732 881
rect 702 867 708 868
rect 702 863 703 867
rect 707 863 708 867
rect 702 862 708 863
rect 728 839 730 880
rect 804 876 806 910
rect 814 906 820 907
rect 814 902 815 906
rect 819 902 820 906
rect 814 901 820 902
rect 802 875 808 876
rect 802 871 803 875
rect 807 871 808 875
rect 802 870 808 871
rect 746 867 752 868
rect 746 863 747 867
rect 751 863 752 867
rect 746 862 752 863
rect 727 838 731 839
rect 727 833 731 834
rect 694 827 700 828
rect 694 823 695 827
rect 699 823 700 827
rect 694 822 700 823
rect 662 817 668 818
rect 662 813 663 817
rect 667 813 668 817
rect 662 812 668 813
rect 574 791 580 792
rect 574 787 575 791
rect 579 787 580 791
rect 574 786 580 787
rect 558 785 564 786
rect 558 781 559 785
rect 563 781 564 785
rect 558 780 564 781
rect 560 755 562 780
rect 654 777 660 778
rect 654 773 655 777
rect 659 773 660 777
rect 654 772 660 773
rect 656 755 658 772
rect 559 754 563 755
rect 559 749 563 750
rect 615 754 619 755
rect 615 749 619 750
rect 655 754 659 755
rect 655 749 659 750
rect 719 754 723 755
rect 719 749 723 750
rect 616 731 618 749
rect 614 730 620 731
rect 614 726 615 730
rect 619 726 620 730
rect 720 729 722 749
rect 614 725 620 726
rect 718 728 724 729
rect 718 724 719 728
rect 723 724 724 728
rect 622 723 628 724
rect 718 723 724 724
rect 622 719 623 723
rect 627 719 628 723
rect 622 718 628 719
rect 566 699 572 700
rect 566 695 567 699
rect 571 695 572 699
rect 566 694 572 695
rect 554 679 560 680
rect 522 675 528 676
rect 522 671 523 675
rect 527 671 528 675
rect 554 675 555 679
rect 559 675 560 679
rect 554 674 560 675
rect 522 670 528 671
rect 458 667 464 668
rect 458 663 459 667
rect 463 663 464 667
rect 458 662 464 663
rect 407 642 411 643
rect 407 637 411 638
rect 443 642 447 643
rect 443 637 447 638
rect 408 623 410 637
rect 460 632 462 662
rect 535 642 539 643
rect 535 637 539 638
rect 414 631 420 632
rect 414 627 415 631
rect 419 627 420 631
rect 414 626 420 627
rect 458 631 464 632
rect 458 627 459 631
rect 463 627 464 631
rect 458 626 464 627
rect 518 631 524 632
rect 518 627 519 631
rect 523 627 524 631
rect 518 626 524 627
rect 406 622 412 623
rect 406 618 407 622
rect 411 618 412 622
rect 406 617 412 618
rect 398 595 404 596
rect 398 591 399 595
rect 403 591 404 595
rect 398 590 404 591
rect 398 584 404 585
rect 398 580 399 584
rect 403 580 404 584
rect 398 579 404 580
rect 378 563 384 564
rect 400 563 402 579
rect 378 559 379 563
rect 383 559 384 563
rect 378 558 384 559
rect 391 562 395 563
rect 380 488 382 558
rect 391 557 395 558
rect 399 562 403 563
rect 399 557 403 558
rect 392 537 394 557
rect 390 536 396 537
rect 390 532 391 536
rect 395 532 396 536
rect 390 531 396 532
rect 398 498 404 499
rect 398 494 399 498
rect 403 494 404 498
rect 398 493 404 494
rect 322 487 328 488
rect 322 483 323 487
rect 327 483 328 487
rect 322 482 328 483
rect 378 487 384 488
rect 378 483 379 487
rect 383 483 384 487
rect 378 482 384 483
rect 390 487 396 488
rect 390 483 391 487
rect 395 483 396 487
rect 390 482 396 483
rect 314 479 320 480
rect 314 475 315 479
rect 319 475 320 479
rect 314 474 320 475
rect 324 452 326 482
rect 382 479 388 480
rect 382 475 383 479
rect 387 475 388 479
rect 382 474 388 475
rect 322 451 328 452
rect 322 447 323 451
rect 327 447 328 451
rect 322 446 328 447
rect 303 442 307 443
rect 303 437 307 438
rect 375 442 379 443
rect 375 437 379 438
rect 294 403 300 404
rect 294 399 295 403
rect 299 399 300 403
rect 294 398 300 399
rect 304 395 306 437
rect 310 423 316 424
rect 310 419 311 423
rect 315 419 316 423
rect 310 418 316 419
rect 312 404 314 418
rect 354 407 360 408
rect 310 403 316 404
rect 310 399 311 403
rect 315 399 316 403
rect 354 403 355 407
rect 359 403 360 407
rect 354 402 360 403
rect 310 398 316 399
rect 302 394 308 395
rect 302 390 303 394
rect 307 390 308 394
rect 302 389 308 390
rect 262 374 268 375
rect 262 370 263 374
rect 267 370 268 374
rect 262 369 268 370
rect 356 368 358 402
rect 376 400 378 437
rect 384 408 386 474
rect 392 416 394 482
rect 400 443 402 493
rect 406 491 412 492
rect 406 487 407 491
rect 411 490 412 491
rect 416 490 418 626
rect 471 562 475 563
rect 471 557 475 558
rect 472 541 474 557
rect 470 540 476 541
rect 470 536 471 540
rect 475 536 476 540
rect 470 535 476 536
rect 458 527 464 528
rect 458 523 459 527
rect 463 523 464 527
rect 458 522 464 523
rect 411 488 418 490
rect 411 487 412 488
rect 406 486 412 487
rect 408 460 410 486
rect 460 484 462 522
rect 498 519 504 520
rect 498 515 499 519
rect 503 515 504 519
rect 498 514 504 515
rect 506 517 512 518
rect 470 493 476 494
rect 470 489 471 493
rect 475 489 476 493
rect 470 488 476 489
rect 458 483 464 484
rect 458 479 459 483
rect 463 479 464 483
rect 458 478 464 479
rect 406 459 412 460
rect 406 455 407 459
rect 411 455 412 459
rect 406 454 412 455
rect 472 443 474 488
rect 478 487 484 488
rect 478 483 479 487
rect 483 483 484 487
rect 478 482 484 483
rect 399 442 403 443
rect 399 437 403 438
rect 415 442 419 443
rect 415 437 419 438
rect 447 442 451 443
rect 447 437 451 438
rect 471 442 475 443
rect 471 437 475 438
rect 390 415 396 416
rect 390 411 391 415
rect 395 411 396 415
rect 390 410 396 411
rect 382 407 388 408
rect 382 403 383 407
rect 387 403 388 407
rect 382 402 388 403
rect 374 399 380 400
rect 374 395 375 399
rect 379 395 380 399
rect 374 394 380 395
rect 392 372 394 410
rect 416 375 418 437
rect 448 375 450 437
rect 480 408 482 482
rect 500 476 502 514
rect 506 513 507 517
rect 511 513 512 517
rect 506 512 512 513
rect 498 475 504 476
rect 498 471 499 475
rect 503 471 504 475
rect 498 470 504 471
rect 508 443 510 512
rect 487 442 491 443
rect 487 437 491 438
rect 507 442 511 443
rect 507 437 511 438
rect 478 407 484 408
rect 478 403 479 407
rect 483 403 484 407
rect 478 402 484 403
rect 488 378 490 437
rect 520 380 522 626
rect 536 624 538 637
rect 556 632 558 674
rect 554 631 560 632
rect 554 627 555 631
rect 559 627 560 631
rect 554 626 560 627
rect 534 623 540 624
rect 534 619 535 623
rect 539 619 540 623
rect 534 618 540 619
rect 526 611 532 612
rect 526 607 527 611
rect 531 607 532 611
rect 526 606 532 607
rect 528 564 530 606
rect 534 582 540 583
rect 534 578 535 582
rect 539 578 540 582
rect 534 577 540 578
rect 526 563 532 564
rect 536 563 538 577
rect 526 559 527 563
rect 531 559 532 563
rect 526 558 532 559
rect 535 562 539 563
rect 535 557 539 558
rect 536 533 538 557
rect 534 532 540 533
rect 534 528 535 532
rect 539 528 540 532
rect 534 527 540 528
rect 568 484 570 694
rect 614 689 620 690
rect 614 685 615 689
rect 619 685 620 689
rect 624 685 626 718
rect 730 711 736 712
rect 730 707 731 711
rect 735 707 736 711
rect 730 706 736 707
rect 718 705 724 706
rect 718 701 719 705
rect 723 701 724 705
rect 718 700 724 701
rect 614 684 620 685
rect 623 684 627 685
rect 616 643 618 684
rect 623 679 627 680
rect 720 643 722 700
rect 615 642 619 643
rect 671 642 675 643
rect 615 637 619 638
rect 634 639 640 640
rect 634 635 635 639
rect 639 635 640 639
rect 671 637 675 638
rect 719 642 723 643
rect 719 637 723 638
rect 634 634 640 635
rect 636 532 638 634
rect 672 603 674 637
rect 686 631 692 632
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 670 602 676 603
rect 670 598 671 602
rect 675 598 676 602
rect 670 597 676 598
rect 688 592 690 626
rect 732 608 734 706
rect 748 688 750 862
rect 816 839 818 901
rect 824 900 826 974
rect 822 899 828 900
rect 822 895 823 899
rect 827 895 828 899
rect 822 894 828 895
rect 815 838 819 839
rect 815 833 819 834
rect 816 824 818 833
rect 832 832 834 1026
rect 856 1020 858 1114
rect 862 1075 868 1076
rect 862 1071 863 1075
rect 867 1071 868 1075
rect 862 1070 868 1071
rect 864 1032 866 1070
rect 916 1056 918 1209
rect 952 1208 954 1350
rect 975 1345 979 1346
rect 983 1350 987 1351
rect 983 1345 987 1346
rect 1023 1350 1027 1351
rect 1023 1345 1027 1346
rect 984 1325 986 1345
rect 982 1324 988 1325
rect 982 1320 983 1324
rect 987 1320 988 1324
rect 1024 1321 1026 1345
rect 982 1319 988 1320
rect 1022 1320 1028 1321
rect 1022 1316 1023 1320
rect 1027 1316 1028 1320
rect 1022 1315 1028 1316
rect 970 1311 976 1312
rect 970 1307 971 1311
rect 975 1307 976 1311
rect 970 1306 976 1307
rect 962 1303 968 1304
rect 962 1299 963 1303
rect 967 1299 968 1303
rect 962 1298 968 1299
rect 964 1272 966 1298
rect 962 1271 968 1272
rect 962 1267 963 1271
rect 967 1267 968 1271
rect 972 1268 974 1306
rect 1022 1292 1028 1293
rect 1022 1288 1023 1292
rect 1027 1288 1028 1292
rect 1022 1287 1028 1288
rect 982 1277 988 1278
rect 982 1273 983 1277
rect 987 1273 988 1277
rect 982 1272 988 1273
rect 962 1266 968 1267
rect 970 1267 976 1268
rect 970 1263 971 1267
rect 975 1263 976 1267
rect 984 1263 986 1272
rect 1024 1263 1026 1287
rect 1038 1279 1044 1280
rect 1038 1275 1039 1279
rect 1043 1278 1044 1279
rect 1048 1278 1050 1410
rect 1064 1401 1066 1425
rect 1070 1407 1076 1408
rect 1070 1403 1071 1407
rect 1075 1403 1076 1407
rect 1070 1402 1076 1403
rect 1062 1400 1068 1401
rect 1062 1396 1063 1400
rect 1067 1396 1068 1400
rect 1054 1395 1060 1396
rect 1062 1395 1068 1396
rect 1054 1391 1055 1395
rect 1059 1391 1060 1395
rect 1054 1390 1060 1391
rect 1043 1276 1050 1278
rect 1043 1275 1044 1276
rect 1038 1274 1044 1275
rect 1056 1264 1058 1390
rect 1072 1384 1074 1402
rect 1112 1392 1114 1425
rect 1122 1419 1128 1420
rect 1122 1415 1123 1419
rect 1127 1415 1128 1419
rect 1122 1414 1128 1415
rect 1110 1391 1116 1392
rect 1102 1387 1108 1388
rect 1070 1383 1076 1384
rect 1070 1379 1071 1383
rect 1075 1379 1076 1383
rect 1102 1383 1103 1387
rect 1107 1383 1108 1387
rect 1110 1387 1111 1391
rect 1115 1387 1116 1391
rect 1110 1386 1116 1387
rect 1102 1382 1108 1383
rect 1070 1378 1076 1379
rect 1062 1372 1068 1373
rect 1062 1368 1063 1372
rect 1067 1368 1068 1372
rect 1062 1367 1068 1368
rect 1064 1351 1066 1367
rect 1063 1350 1067 1351
rect 1063 1345 1067 1346
rect 1064 1321 1066 1345
rect 1062 1320 1068 1321
rect 1062 1316 1063 1320
rect 1067 1316 1068 1320
rect 1062 1315 1068 1316
rect 1062 1301 1068 1302
rect 1062 1297 1063 1301
rect 1067 1297 1068 1301
rect 1062 1296 1068 1297
rect 1054 1263 1060 1264
rect 1064 1263 1066 1296
rect 1104 1278 1106 1382
rect 1124 1380 1126 1414
rect 1130 1395 1136 1396
rect 1130 1391 1131 1395
rect 1135 1391 1136 1395
rect 1130 1390 1136 1391
rect 1122 1379 1128 1380
rect 1122 1375 1123 1379
rect 1127 1375 1128 1379
rect 1122 1374 1128 1375
rect 1110 1373 1116 1374
rect 1110 1369 1111 1373
rect 1115 1369 1116 1373
rect 1110 1368 1116 1369
rect 1112 1351 1114 1368
rect 1124 1356 1126 1374
rect 1122 1355 1128 1356
rect 1122 1351 1123 1355
rect 1127 1351 1128 1355
rect 1111 1350 1115 1351
rect 1122 1350 1128 1351
rect 1111 1345 1115 1346
rect 1132 1312 1134 1390
rect 1130 1311 1136 1312
rect 1130 1307 1131 1311
rect 1135 1307 1136 1311
rect 1130 1306 1136 1307
rect 1140 1280 1142 1442
rect 1168 1431 1170 1453
rect 1182 1451 1188 1452
rect 1182 1447 1183 1451
rect 1187 1447 1188 1451
rect 1182 1446 1188 1447
rect 1151 1430 1155 1431
rect 1151 1425 1155 1426
rect 1167 1430 1171 1431
rect 1167 1425 1171 1426
rect 1152 1401 1154 1425
rect 1150 1400 1156 1401
rect 1150 1396 1151 1400
rect 1155 1396 1156 1400
rect 1150 1395 1156 1396
rect 1166 1387 1172 1388
rect 1166 1383 1167 1387
rect 1171 1383 1172 1387
rect 1166 1382 1172 1383
rect 1150 1372 1156 1373
rect 1150 1368 1151 1372
rect 1155 1368 1156 1372
rect 1150 1367 1156 1368
rect 1152 1351 1154 1367
rect 1151 1350 1155 1351
rect 1151 1345 1155 1346
rect 1159 1350 1163 1351
rect 1159 1345 1163 1346
rect 1160 1321 1162 1345
rect 1168 1344 1170 1382
rect 1166 1343 1172 1344
rect 1166 1339 1167 1343
rect 1171 1339 1172 1343
rect 1166 1338 1172 1339
rect 1158 1320 1164 1321
rect 1158 1316 1159 1320
rect 1163 1316 1164 1320
rect 1158 1315 1164 1316
rect 1174 1299 1180 1300
rect 1174 1295 1175 1299
rect 1179 1295 1180 1299
rect 1174 1294 1180 1295
rect 1110 1279 1116 1280
rect 1110 1278 1111 1279
rect 1104 1276 1111 1278
rect 1110 1275 1111 1276
rect 1115 1275 1116 1279
rect 1110 1274 1116 1275
rect 1138 1279 1144 1280
rect 1138 1275 1139 1279
rect 1143 1275 1144 1279
rect 1138 1274 1144 1275
rect 1154 1279 1160 1280
rect 1154 1274 1155 1279
rect 1159 1274 1160 1279
rect 1155 1271 1159 1272
rect 1176 1263 1178 1294
rect 959 1262 963 1263
rect 970 1262 976 1263
rect 983 1262 987 1263
rect 959 1257 963 1258
rect 983 1257 987 1258
rect 1015 1262 1019 1263
rect 1015 1257 1019 1258
rect 1023 1262 1027 1263
rect 1054 1259 1055 1263
rect 1059 1259 1060 1263
rect 1054 1258 1060 1259
rect 1063 1262 1067 1263
rect 1023 1257 1027 1258
rect 1063 1257 1067 1258
rect 1087 1262 1091 1263
rect 1087 1257 1091 1258
rect 1127 1262 1131 1263
rect 1127 1257 1131 1258
rect 1159 1262 1163 1263
rect 1159 1257 1163 1258
rect 1175 1262 1179 1263
rect 1175 1257 1179 1258
rect 950 1207 956 1208
rect 950 1203 951 1207
rect 955 1203 956 1207
rect 950 1202 956 1203
rect 960 1198 962 1257
rect 990 1255 996 1256
rect 990 1251 991 1255
rect 995 1251 996 1255
rect 990 1250 996 1251
rect 992 1232 994 1250
rect 990 1231 996 1232
rect 990 1227 991 1231
rect 995 1227 996 1231
rect 990 1226 996 1227
rect 992 1200 994 1226
rect 1016 1215 1018 1257
rect 1066 1227 1072 1228
rect 1038 1223 1044 1224
rect 1038 1219 1039 1223
rect 1043 1219 1044 1223
rect 1066 1223 1067 1227
rect 1071 1223 1072 1227
rect 1066 1222 1072 1223
rect 1038 1218 1044 1219
rect 1014 1214 1020 1215
rect 1014 1210 1015 1214
rect 1019 1210 1020 1214
rect 1014 1209 1020 1210
rect 990 1199 996 1200
rect 958 1197 964 1198
rect 958 1193 959 1197
rect 963 1193 964 1197
rect 990 1195 991 1199
rect 995 1195 996 1199
rect 990 1194 996 1195
rect 958 1192 964 1193
rect 930 1179 936 1180
rect 930 1178 931 1179
rect 924 1176 931 1178
rect 924 1080 926 1176
rect 930 1175 931 1176
rect 935 1175 936 1179
rect 930 1174 936 1175
rect 1006 1176 1012 1177
rect 1006 1172 1007 1176
rect 1011 1172 1012 1176
rect 1006 1171 1012 1172
rect 974 1170 980 1171
rect 974 1166 975 1170
rect 979 1166 980 1170
rect 974 1165 980 1166
rect 976 1151 978 1165
rect 1008 1151 1010 1171
rect 935 1150 939 1151
rect 935 1145 939 1146
rect 967 1150 971 1151
rect 967 1145 971 1146
rect 975 1150 979 1151
rect 975 1145 979 1146
rect 999 1150 1003 1151
rect 999 1145 1003 1146
rect 1007 1150 1011 1151
rect 1007 1145 1011 1146
rect 1031 1150 1035 1151
rect 1031 1145 1035 1146
rect 936 1124 938 1145
rect 954 1143 960 1144
rect 954 1139 955 1143
rect 959 1139 960 1143
rect 954 1138 960 1139
rect 934 1123 940 1124
rect 934 1119 935 1123
rect 939 1119 940 1123
rect 934 1118 940 1119
rect 934 1106 940 1107
rect 934 1102 935 1106
rect 939 1102 940 1106
rect 934 1101 940 1102
rect 922 1079 928 1080
rect 922 1075 923 1079
rect 927 1075 928 1079
rect 922 1074 928 1075
rect 914 1055 920 1056
rect 914 1051 915 1055
rect 919 1051 920 1055
rect 914 1050 920 1051
rect 936 1035 938 1101
rect 956 1100 958 1138
rect 968 1124 970 1145
rect 1000 1125 1002 1145
rect 998 1124 1004 1125
rect 1032 1124 1034 1145
rect 966 1123 972 1124
rect 966 1119 967 1123
rect 971 1119 972 1123
rect 998 1120 999 1124
rect 1003 1120 1004 1124
rect 1030 1123 1036 1124
rect 998 1119 1004 1120
rect 1014 1119 1020 1120
rect 966 1118 972 1119
rect 1014 1115 1015 1119
rect 1019 1115 1020 1119
rect 1030 1119 1031 1123
rect 1035 1119 1036 1123
rect 1030 1118 1036 1119
rect 1014 1114 1020 1115
rect 966 1106 972 1107
rect 966 1102 967 1106
rect 971 1102 972 1106
rect 966 1101 972 1102
rect 998 1101 1004 1102
rect 954 1099 960 1100
rect 954 1095 955 1099
rect 959 1095 960 1099
rect 954 1094 960 1095
rect 968 1035 970 1101
rect 998 1097 999 1101
rect 1003 1097 1004 1101
rect 998 1096 1004 1097
rect 1000 1035 1002 1096
rect 919 1034 923 1035
rect 862 1031 868 1032
rect 862 1027 863 1031
rect 867 1027 868 1031
rect 919 1029 923 1030
rect 935 1034 939 1035
rect 935 1029 939 1030
rect 967 1034 971 1035
rect 967 1029 971 1030
rect 975 1034 979 1035
rect 975 1029 979 1030
rect 999 1034 1003 1035
rect 999 1029 1003 1030
rect 862 1026 868 1027
rect 842 1019 848 1020
rect 842 1015 843 1019
rect 847 1015 848 1019
rect 842 1014 848 1015
rect 854 1019 860 1020
rect 854 1015 855 1019
rect 859 1015 860 1019
rect 854 1014 860 1015
rect 844 883 846 1014
rect 920 995 922 1029
rect 976 1010 978 1029
rect 1016 1024 1018 1114
rect 1030 1106 1036 1107
rect 1030 1102 1031 1106
rect 1035 1102 1036 1106
rect 1030 1101 1036 1102
rect 1032 1035 1034 1101
rect 1040 1064 1042 1218
rect 1068 1188 1070 1222
rect 1088 1220 1090 1257
rect 1102 1223 1108 1224
rect 1078 1219 1084 1220
rect 1078 1215 1079 1219
rect 1083 1215 1084 1219
rect 1078 1214 1084 1215
rect 1086 1219 1092 1220
rect 1086 1215 1087 1219
rect 1091 1215 1092 1219
rect 1102 1219 1103 1223
rect 1107 1219 1108 1223
rect 1102 1218 1108 1219
rect 1086 1214 1092 1215
rect 1080 1192 1082 1214
rect 1078 1191 1084 1192
rect 1066 1187 1072 1188
rect 1066 1183 1067 1187
rect 1071 1183 1072 1187
rect 1078 1187 1079 1191
rect 1083 1187 1084 1191
rect 1078 1186 1084 1187
rect 1066 1182 1072 1183
rect 1086 1172 1092 1173
rect 1086 1168 1087 1172
rect 1091 1168 1092 1172
rect 1086 1167 1092 1168
rect 1088 1151 1090 1167
rect 1063 1150 1067 1151
rect 1063 1145 1067 1146
rect 1087 1150 1091 1151
rect 1087 1145 1091 1146
rect 1095 1150 1099 1151
rect 1095 1145 1099 1146
rect 1064 1124 1066 1145
rect 1096 1125 1098 1145
rect 1094 1124 1100 1125
rect 1062 1123 1068 1124
rect 1062 1119 1063 1123
rect 1067 1119 1068 1123
rect 1094 1120 1095 1124
rect 1099 1120 1100 1124
rect 1094 1119 1100 1120
rect 1062 1118 1068 1119
rect 1082 1115 1088 1116
rect 1082 1111 1083 1115
rect 1087 1111 1088 1115
rect 1082 1110 1088 1111
rect 1062 1106 1068 1107
rect 1062 1102 1063 1106
rect 1067 1102 1068 1106
rect 1062 1101 1068 1102
rect 1038 1063 1044 1064
rect 1038 1059 1039 1063
rect 1043 1059 1044 1063
rect 1038 1058 1044 1059
rect 1064 1035 1066 1101
rect 1075 1092 1079 1093
rect 1075 1087 1079 1088
rect 1031 1034 1035 1035
rect 1031 1029 1035 1030
rect 1063 1034 1067 1035
rect 1063 1029 1067 1030
rect 1014 1023 1020 1024
rect 1014 1019 1015 1023
rect 1019 1019 1020 1023
rect 1014 1018 1020 1019
rect 1046 1019 1052 1020
rect 1046 1015 1047 1019
rect 1051 1015 1052 1019
rect 1046 1014 1052 1015
rect 974 1009 980 1010
rect 974 1005 975 1009
rect 979 1005 980 1009
rect 974 1004 980 1005
rect 918 994 924 995
rect 918 990 919 994
rect 923 990 924 994
rect 918 989 924 990
rect 934 983 940 984
rect 934 979 935 983
rect 939 979 940 983
rect 934 978 940 979
rect 918 977 924 978
rect 918 973 919 977
rect 923 973 924 977
rect 918 972 924 973
rect 854 955 860 956
rect 920 955 922 972
rect 854 951 855 955
rect 859 951 860 955
rect 854 950 860 951
rect 863 954 867 955
rect 856 896 858 950
rect 863 949 867 950
rect 919 954 923 955
rect 919 949 923 950
rect 864 927 866 949
rect 862 926 868 927
rect 862 922 863 926
rect 867 922 868 926
rect 862 921 868 922
rect 854 895 860 896
rect 854 891 855 895
rect 859 891 860 895
rect 854 890 860 891
rect 862 885 868 886
rect 844 881 854 883
rect 852 844 854 881
rect 862 881 863 885
rect 867 881 868 885
rect 862 880 868 881
rect 850 843 856 844
rect 850 839 851 843
rect 855 839 856 843
rect 864 839 866 880
rect 936 876 938 978
rect 966 969 972 970
rect 966 965 967 969
rect 971 965 972 969
rect 966 964 972 965
rect 968 955 970 964
rect 951 954 955 955
rect 951 949 955 950
rect 967 954 971 955
rect 967 949 971 950
rect 983 954 987 955
rect 983 949 987 950
rect 1039 954 1043 955
rect 1039 949 1043 950
rect 952 924 954 949
rect 984 925 986 949
rect 990 931 996 932
rect 990 927 991 931
rect 995 927 996 931
rect 990 926 996 927
rect 982 924 988 925
rect 950 923 956 924
rect 950 919 951 923
rect 955 919 956 923
rect 982 920 983 924
rect 987 920 988 924
rect 982 919 988 920
rect 950 918 956 919
rect 970 915 976 916
rect 970 911 971 915
rect 975 911 976 915
rect 970 910 976 911
rect 950 906 956 907
rect 950 902 951 906
rect 955 902 956 906
rect 950 901 956 902
rect 934 875 940 876
rect 934 871 935 875
rect 939 871 940 875
rect 934 870 940 871
rect 886 859 892 860
rect 886 855 887 859
rect 891 855 892 859
rect 886 854 892 855
rect 850 838 856 839
rect 863 838 867 839
rect 830 831 836 832
rect 830 827 831 831
rect 835 827 836 831
rect 830 826 836 827
rect 814 823 820 824
rect 814 819 815 823
rect 819 819 820 823
rect 814 818 820 819
rect 814 782 820 783
rect 814 778 815 782
rect 819 778 820 782
rect 814 777 820 778
rect 816 755 818 777
rect 767 754 771 755
rect 767 749 771 750
rect 815 754 819 755
rect 815 749 819 750
rect 768 736 770 749
rect 766 735 772 736
rect 766 731 767 735
rect 771 731 772 735
rect 766 730 772 731
rect 766 723 772 724
rect 766 719 767 723
rect 771 719 772 723
rect 766 718 772 719
rect 746 687 752 688
rect 746 683 747 687
rect 751 683 752 687
rect 746 682 752 683
rect 758 683 764 684
rect 758 679 759 683
rect 763 679 764 683
rect 758 678 764 679
rect 760 616 762 678
rect 768 676 770 718
rect 774 695 780 696
rect 774 691 775 695
rect 779 691 780 695
rect 774 690 780 691
rect 766 675 772 676
rect 766 671 767 675
rect 771 671 772 675
rect 766 670 772 671
rect 776 643 778 690
rect 832 680 834 826
rect 842 719 848 720
rect 842 715 843 719
rect 847 715 848 719
rect 842 714 848 715
rect 830 679 836 680
rect 830 675 831 679
rect 835 675 836 679
rect 830 674 836 675
rect 767 642 771 643
rect 767 637 771 638
rect 775 642 779 643
rect 775 637 779 638
rect 768 624 770 637
rect 832 624 834 674
rect 844 668 846 714
rect 852 692 854 838
rect 863 833 867 834
rect 888 832 890 854
rect 952 839 954 901
rect 972 884 974 910
rect 992 900 994 926
rect 1040 924 1042 949
rect 1038 923 1044 924
rect 1038 919 1039 923
rect 1043 919 1044 923
rect 1038 918 1044 919
rect 1038 906 1044 907
rect 998 903 1004 904
rect 990 899 996 900
rect 990 895 991 899
rect 995 895 996 899
rect 998 899 999 903
rect 1003 899 1004 903
rect 1038 902 1039 906
rect 1043 902 1044 906
rect 1038 901 1044 902
rect 998 898 1004 899
rect 990 894 996 895
rect 970 883 976 884
rect 970 879 971 883
rect 975 879 976 883
rect 970 878 976 879
rect 951 838 955 839
rect 951 833 955 834
rect 886 831 892 832
rect 886 827 887 831
rect 891 827 892 831
rect 886 826 892 827
rect 952 808 954 833
rect 992 824 994 894
rect 1000 839 1002 898
rect 1040 839 1042 901
rect 1048 888 1050 1014
rect 1064 1005 1066 1029
rect 1076 1012 1078 1087
rect 1074 1011 1080 1012
rect 1074 1007 1075 1011
rect 1079 1007 1080 1011
rect 1074 1006 1080 1007
rect 1062 1004 1068 1005
rect 1062 1000 1063 1004
rect 1067 1000 1068 1004
rect 1062 999 1068 1000
rect 1062 976 1068 977
rect 1062 972 1063 976
rect 1067 972 1068 976
rect 1062 971 1068 972
rect 1064 955 1066 971
rect 1084 964 1086 1110
rect 1094 1096 1100 1097
rect 1094 1092 1095 1096
rect 1099 1092 1100 1096
rect 1094 1091 1100 1092
rect 1096 1035 1098 1091
rect 1104 1084 1106 1218
rect 1128 1195 1130 1257
rect 1160 1195 1162 1257
rect 1126 1194 1132 1195
rect 1126 1190 1127 1194
rect 1131 1190 1132 1194
rect 1126 1189 1132 1190
rect 1158 1194 1164 1195
rect 1158 1190 1159 1194
rect 1163 1190 1164 1194
rect 1158 1189 1164 1190
rect 1142 1183 1148 1184
rect 1142 1179 1143 1183
rect 1147 1179 1148 1183
rect 1142 1178 1148 1179
rect 1126 1177 1132 1178
rect 1126 1173 1127 1177
rect 1131 1173 1132 1177
rect 1126 1172 1132 1173
rect 1128 1151 1130 1172
rect 1127 1150 1131 1151
rect 1127 1145 1131 1146
rect 1135 1150 1139 1151
rect 1135 1145 1139 1146
rect 1136 1124 1138 1145
rect 1144 1144 1146 1178
rect 1158 1177 1164 1178
rect 1158 1173 1159 1177
rect 1163 1173 1164 1177
rect 1158 1172 1164 1173
rect 1160 1151 1162 1172
rect 1159 1150 1163 1151
rect 1159 1145 1163 1146
rect 1167 1150 1171 1151
rect 1167 1145 1171 1146
rect 1142 1143 1148 1144
rect 1142 1139 1143 1143
rect 1147 1139 1148 1143
rect 1142 1138 1148 1139
rect 1168 1125 1170 1145
rect 1166 1124 1172 1125
rect 1134 1123 1140 1124
rect 1134 1119 1135 1123
rect 1139 1119 1140 1123
rect 1166 1120 1167 1124
rect 1171 1120 1172 1124
rect 1166 1119 1172 1120
rect 1134 1118 1140 1119
rect 1122 1115 1128 1116
rect 1122 1111 1123 1115
rect 1127 1111 1128 1115
rect 1122 1110 1128 1111
rect 1110 1107 1116 1108
rect 1110 1103 1111 1107
rect 1115 1103 1116 1107
rect 1110 1102 1116 1103
rect 1102 1083 1108 1084
rect 1102 1079 1103 1083
rect 1107 1079 1108 1083
rect 1102 1078 1108 1079
rect 1095 1034 1099 1035
rect 1095 1029 1099 1030
rect 1112 971 1114 1102
rect 1124 1088 1126 1110
rect 1134 1106 1140 1107
rect 1134 1102 1135 1106
rect 1139 1102 1140 1106
rect 1134 1101 1140 1102
rect 1122 1087 1128 1088
rect 1122 1083 1123 1087
rect 1127 1083 1128 1087
rect 1122 1082 1128 1083
rect 1136 1035 1138 1101
rect 1174 1086 1180 1087
rect 1174 1082 1175 1086
rect 1179 1082 1180 1086
rect 1174 1081 1180 1082
rect 1176 1035 1178 1081
rect 1119 1034 1123 1035
rect 1119 1029 1123 1030
rect 1135 1034 1139 1035
rect 1135 1029 1139 1030
rect 1167 1034 1171 1035
rect 1167 1029 1171 1030
rect 1175 1034 1179 1035
rect 1175 1029 1179 1030
rect 1120 998 1122 1029
rect 1118 997 1124 998
rect 1118 993 1119 997
rect 1123 993 1124 997
rect 1168 995 1170 1029
rect 1184 1016 1186 1446
rect 1190 1443 1196 1444
rect 1190 1439 1191 1443
rect 1195 1439 1196 1443
rect 1190 1438 1196 1439
rect 1192 1428 1194 1438
rect 1200 1431 1202 1453
rect 1216 1452 1218 1526
rect 1239 1498 1243 1499
rect 1239 1493 1243 1494
rect 1240 1476 1242 1493
rect 1238 1475 1244 1476
rect 1238 1471 1239 1475
rect 1243 1471 1244 1475
rect 1238 1470 1244 1471
rect 1256 1468 1258 1530
rect 1272 1527 1274 1537
rect 1360 1527 1362 1537
rect 1376 1532 1378 1562
rect 1398 1558 1404 1559
rect 1398 1554 1399 1558
rect 1403 1554 1404 1558
rect 1398 1553 1404 1554
rect 1470 1558 1476 1559
rect 1470 1554 1471 1558
rect 1475 1554 1476 1558
rect 1470 1553 1476 1554
rect 1400 1543 1402 1553
rect 1472 1543 1474 1553
rect 1399 1542 1403 1543
rect 1399 1537 1403 1538
rect 1439 1542 1443 1543
rect 1439 1537 1443 1538
rect 1471 1542 1475 1543
rect 1471 1537 1475 1538
rect 1374 1531 1380 1532
rect 1374 1527 1375 1531
rect 1379 1527 1380 1531
rect 1440 1527 1442 1537
rect 1446 1531 1452 1532
rect 1446 1527 1447 1531
rect 1451 1527 1452 1531
rect 1270 1526 1276 1527
rect 1270 1522 1271 1526
rect 1275 1522 1276 1526
rect 1270 1521 1276 1522
rect 1358 1526 1364 1527
rect 1374 1526 1380 1527
rect 1438 1526 1444 1527
rect 1446 1526 1452 1527
rect 1358 1522 1359 1526
rect 1363 1522 1364 1526
rect 1358 1521 1364 1522
rect 1438 1522 1439 1526
rect 1443 1522 1444 1526
rect 1438 1521 1444 1522
rect 1334 1515 1340 1516
rect 1334 1511 1335 1515
rect 1339 1511 1340 1515
rect 1334 1510 1340 1511
rect 1374 1515 1380 1516
rect 1374 1511 1375 1515
rect 1379 1511 1380 1515
rect 1374 1510 1380 1511
rect 1270 1509 1276 1510
rect 1270 1505 1271 1509
rect 1275 1505 1276 1509
rect 1270 1504 1276 1505
rect 1272 1499 1274 1504
rect 1271 1498 1275 1499
rect 1271 1493 1275 1494
rect 1279 1498 1283 1499
rect 1279 1493 1283 1494
rect 1319 1498 1323 1499
rect 1319 1493 1323 1494
rect 1280 1476 1282 1493
rect 1320 1476 1322 1493
rect 1278 1475 1284 1476
rect 1278 1471 1279 1475
rect 1283 1471 1284 1475
rect 1278 1470 1284 1471
rect 1318 1475 1324 1476
rect 1318 1471 1319 1475
rect 1323 1471 1324 1475
rect 1318 1470 1324 1471
rect 1230 1467 1236 1468
rect 1230 1463 1231 1467
rect 1235 1463 1236 1467
rect 1230 1462 1236 1463
rect 1254 1467 1260 1468
rect 1254 1463 1255 1467
rect 1259 1463 1260 1467
rect 1254 1462 1260 1463
rect 1214 1451 1220 1452
rect 1214 1447 1215 1451
rect 1219 1447 1220 1451
rect 1214 1446 1220 1447
rect 1199 1430 1203 1431
rect 1190 1427 1196 1428
rect 1190 1423 1191 1427
rect 1195 1423 1196 1427
rect 1199 1425 1203 1426
rect 1190 1422 1196 1423
rect 1192 1400 1194 1422
rect 1190 1399 1196 1400
rect 1190 1395 1191 1399
rect 1195 1395 1196 1399
rect 1190 1394 1196 1395
rect 1192 1284 1194 1394
rect 1200 1391 1202 1425
rect 1216 1420 1218 1446
rect 1214 1419 1220 1420
rect 1214 1415 1215 1419
rect 1219 1415 1220 1419
rect 1214 1414 1220 1415
rect 1232 1412 1234 1462
rect 1238 1458 1244 1459
rect 1318 1458 1324 1459
rect 1238 1454 1239 1458
rect 1243 1454 1244 1458
rect 1238 1453 1244 1454
rect 1278 1457 1284 1458
rect 1278 1453 1279 1457
rect 1283 1453 1284 1457
rect 1318 1454 1319 1458
rect 1323 1454 1324 1458
rect 1318 1453 1324 1454
rect 1240 1431 1242 1453
rect 1278 1452 1284 1453
rect 1280 1431 1282 1452
rect 1298 1451 1304 1452
rect 1298 1447 1299 1451
rect 1303 1447 1304 1451
rect 1298 1446 1304 1447
rect 1239 1430 1243 1431
rect 1239 1425 1243 1426
rect 1263 1430 1267 1431
rect 1263 1425 1267 1426
rect 1279 1430 1283 1431
rect 1279 1425 1283 1426
rect 1230 1411 1236 1412
rect 1214 1407 1220 1408
rect 1214 1403 1215 1407
rect 1219 1403 1220 1407
rect 1230 1407 1231 1411
rect 1235 1407 1236 1411
rect 1230 1406 1236 1407
rect 1214 1402 1220 1403
rect 1198 1390 1204 1391
rect 1198 1386 1199 1390
rect 1203 1386 1204 1390
rect 1198 1385 1204 1386
rect 1216 1380 1218 1402
rect 1264 1394 1266 1425
rect 1262 1393 1268 1394
rect 1262 1389 1263 1393
rect 1267 1389 1268 1393
rect 1262 1388 1268 1389
rect 1300 1384 1302 1446
rect 1320 1431 1322 1453
rect 1336 1452 1338 1510
rect 1358 1509 1364 1510
rect 1358 1505 1359 1509
rect 1363 1505 1364 1509
rect 1358 1504 1364 1505
rect 1360 1499 1362 1504
rect 1359 1498 1363 1499
rect 1359 1493 1363 1494
rect 1360 1476 1362 1493
rect 1358 1475 1364 1476
rect 1358 1471 1359 1475
rect 1363 1471 1364 1475
rect 1358 1470 1364 1471
rect 1358 1458 1364 1459
rect 1358 1454 1359 1458
rect 1363 1454 1364 1458
rect 1358 1453 1364 1454
rect 1334 1451 1340 1452
rect 1334 1447 1335 1451
rect 1339 1447 1340 1451
rect 1334 1446 1340 1447
rect 1360 1431 1362 1453
rect 1376 1452 1378 1510
rect 1438 1509 1444 1510
rect 1438 1505 1439 1509
rect 1443 1505 1444 1509
rect 1438 1504 1444 1505
rect 1440 1499 1442 1504
rect 1399 1498 1403 1499
rect 1399 1493 1403 1494
rect 1439 1498 1443 1499
rect 1439 1493 1443 1494
rect 1400 1476 1402 1493
rect 1440 1476 1442 1493
rect 1398 1475 1404 1476
rect 1398 1471 1399 1475
rect 1403 1471 1404 1475
rect 1398 1470 1404 1471
rect 1438 1475 1444 1476
rect 1438 1471 1439 1475
rect 1443 1471 1444 1475
rect 1438 1470 1444 1471
rect 1398 1458 1404 1459
rect 1398 1454 1399 1458
rect 1403 1454 1404 1458
rect 1398 1453 1404 1454
rect 1438 1458 1444 1459
rect 1438 1454 1439 1458
rect 1443 1454 1444 1458
rect 1438 1453 1444 1454
rect 1374 1451 1380 1452
rect 1374 1447 1375 1451
rect 1379 1447 1380 1451
rect 1374 1446 1380 1447
rect 1400 1431 1402 1453
rect 1440 1431 1442 1453
rect 1319 1430 1323 1431
rect 1319 1425 1323 1426
rect 1359 1430 1363 1431
rect 1359 1425 1363 1426
rect 1399 1430 1403 1431
rect 1399 1425 1403 1426
rect 1415 1430 1419 1431
rect 1415 1425 1419 1426
rect 1439 1430 1443 1431
rect 1439 1425 1443 1426
rect 1320 1392 1322 1425
rect 1406 1399 1412 1400
rect 1406 1395 1407 1399
rect 1411 1395 1412 1399
rect 1406 1394 1412 1395
rect 1318 1391 1324 1392
rect 1318 1387 1319 1391
rect 1323 1387 1324 1391
rect 1318 1386 1324 1387
rect 1298 1383 1304 1384
rect 1214 1379 1220 1380
rect 1214 1375 1215 1379
rect 1219 1375 1220 1379
rect 1298 1379 1299 1383
rect 1303 1379 1304 1383
rect 1298 1378 1304 1379
rect 1214 1374 1220 1375
rect 1198 1373 1204 1374
rect 1198 1369 1199 1373
rect 1203 1369 1204 1373
rect 1198 1368 1204 1369
rect 1246 1372 1252 1373
rect 1246 1368 1247 1372
rect 1251 1368 1252 1372
rect 1200 1351 1202 1368
rect 1246 1367 1252 1368
rect 1318 1372 1324 1373
rect 1318 1368 1319 1372
rect 1323 1368 1324 1372
rect 1318 1367 1324 1368
rect 1248 1351 1250 1367
rect 1320 1351 1322 1367
rect 1199 1350 1203 1351
rect 1199 1345 1203 1346
rect 1215 1350 1219 1351
rect 1215 1345 1219 1346
rect 1247 1350 1251 1351
rect 1247 1345 1251 1346
rect 1303 1350 1307 1351
rect 1303 1345 1307 1346
rect 1319 1350 1323 1351
rect 1319 1345 1323 1346
rect 1391 1350 1395 1351
rect 1391 1345 1395 1346
rect 1216 1321 1218 1345
rect 1238 1335 1244 1336
rect 1238 1331 1239 1335
rect 1243 1331 1244 1335
rect 1238 1330 1244 1331
rect 1214 1320 1220 1321
rect 1214 1316 1215 1320
rect 1219 1316 1220 1320
rect 1214 1315 1220 1316
rect 1214 1301 1220 1302
rect 1214 1297 1215 1301
rect 1219 1297 1220 1301
rect 1214 1296 1220 1297
rect 1190 1283 1196 1284
rect 1190 1279 1191 1283
rect 1195 1279 1196 1283
rect 1190 1278 1196 1279
rect 1192 1224 1194 1278
rect 1198 1271 1204 1272
rect 1198 1267 1199 1271
rect 1203 1267 1204 1271
rect 1198 1266 1204 1267
rect 1190 1223 1196 1224
rect 1190 1219 1191 1223
rect 1195 1219 1196 1223
rect 1190 1218 1196 1219
rect 1192 1208 1194 1218
rect 1200 1216 1202 1266
rect 1216 1263 1218 1296
rect 1215 1262 1219 1263
rect 1215 1257 1219 1258
rect 1198 1215 1204 1216
rect 1198 1210 1199 1215
rect 1203 1210 1204 1215
rect 1190 1207 1196 1208
rect 1199 1207 1203 1208
rect 1190 1203 1191 1207
rect 1195 1203 1196 1207
rect 1190 1202 1196 1203
rect 1200 1200 1202 1207
rect 1198 1199 1204 1200
rect 1198 1195 1199 1199
rect 1203 1195 1204 1199
rect 1216 1198 1218 1257
rect 1198 1194 1204 1195
rect 1214 1197 1220 1198
rect 1214 1193 1215 1197
rect 1219 1193 1220 1197
rect 1240 1196 1242 1330
rect 1304 1321 1306 1345
rect 1302 1320 1308 1321
rect 1392 1320 1394 1345
rect 1408 1342 1410 1394
rect 1416 1391 1418 1425
rect 1414 1390 1420 1391
rect 1414 1386 1415 1390
rect 1419 1386 1420 1390
rect 1414 1385 1420 1386
rect 1448 1380 1450 1526
rect 1480 1516 1482 1606
rect 1566 1602 1567 1606
rect 1571 1602 1572 1606
rect 1566 1601 1572 1602
rect 1654 1606 1660 1607
rect 1670 1606 1676 1607
rect 1694 1608 1700 1609
rect 1654 1602 1655 1606
rect 1659 1602 1660 1606
rect 1694 1604 1695 1608
rect 1699 1604 1700 1608
rect 1694 1603 1700 1604
rect 1654 1601 1660 1602
rect 1622 1595 1628 1596
rect 1622 1591 1623 1595
rect 1627 1591 1628 1595
rect 1622 1590 1628 1591
rect 1694 1591 1700 1592
rect 1566 1589 1572 1590
rect 1566 1585 1567 1589
rect 1571 1585 1572 1589
rect 1566 1584 1572 1585
rect 1535 1582 1539 1583
rect 1535 1576 1539 1578
rect 1567 1582 1571 1584
rect 1567 1577 1571 1578
rect 1607 1582 1611 1583
rect 1607 1576 1611 1578
rect 1534 1575 1540 1576
rect 1534 1571 1535 1575
rect 1539 1571 1540 1575
rect 1534 1570 1540 1571
rect 1606 1575 1612 1576
rect 1606 1571 1607 1575
rect 1611 1571 1612 1575
rect 1606 1570 1612 1571
rect 1546 1567 1552 1568
rect 1546 1563 1547 1567
rect 1551 1563 1552 1567
rect 1546 1562 1552 1563
rect 1534 1558 1540 1559
rect 1534 1554 1535 1558
rect 1539 1554 1540 1558
rect 1534 1553 1540 1554
rect 1536 1543 1538 1553
rect 1519 1542 1523 1543
rect 1519 1537 1523 1538
rect 1535 1542 1539 1543
rect 1535 1537 1539 1538
rect 1520 1527 1522 1537
rect 1548 1532 1550 1562
rect 1606 1558 1612 1559
rect 1606 1554 1607 1558
rect 1611 1554 1612 1558
rect 1606 1553 1612 1554
rect 1608 1543 1610 1553
rect 1624 1552 1626 1590
rect 1654 1589 1660 1590
rect 1654 1585 1655 1589
rect 1659 1585 1660 1589
rect 1694 1587 1695 1591
rect 1699 1587 1700 1591
rect 1694 1586 1700 1587
rect 1654 1584 1660 1585
rect 1655 1582 1659 1584
rect 1696 1583 1698 1586
rect 1655 1576 1659 1578
rect 1695 1582 1699 1583
rect 1695 1577 1699 1578
rect 1654 1575 1660 1576
rect 1654 1571 1655 1575
rect 1659 1571 1660 1575
rect 1696 1574 1698 1577
rect 1702 1575 1708 1576
rect 1654 1570 1660 1571
rect 1694 1573 1700 1574
rect 1694 1569 1695 1573
rect 1699 1569 1700 1573
rect 1702 1571 1703 1575
rect 1707 1571 1708 1575
rect 1702 1570 1708 1571
rect 1694 1568 1700 1569
rect 1670 1567 1676 1568
rect 1670 1563 1671 1567
rect 1675 1563 1676 1567
rect 1670 1562 1676 1563
rect 1654 1558 1660 1559
rect 1654 1554 1655 1558
rect 1659 1554 1660 1558
rect 1654 1553 1660 1554
rect 1622 1551 1628 1552
rect 1622 1547 1623 1551
rect 1627 1547 1628 1551
rect 1622 1546 1628 1547
rect 1656 1543 1658 1553
rect 1599 1542 1603 1543
rect 1599 1537 1603 1538
rect 1607 1542 1611 1543
rect 1607 1537 1611 1538
rect 1655 1542 1659 1543
rect 1655 1537 1659 1538
rect 1546 1531 1552 1532
rect 1546 1527 1547 1531
rect 1551 1527 1552 1531
rect 1600 1527 1602 1537
rect 1656 1527 1658 1537
rect 1672 1532 1674 1562
rect 1694 1556 1700 1557
rect 1694 1552 1695 1556
rect 1699 1552 1700 1556
rect 1694 1551 1700 1552
rect 1696 1543 1698 1551
rect 1695 1542 1699 1543
rect 1695 1537 1699 1538
rect 1670 1531 1676 1532
rect 1670 1527 1671 1531
rect 1675 1527 1676 1531
rect 1696 1529 1698 1537
rect 1518 1526 1524 1527
rect 1546 1526 1552 1527
rect 1598 1526 1604 1527
rect 1518 1522 1519 1526
rect 1523 1522 1524 1526
rect 1518 1521 1524 1522
rect 1598 1522 1599 1526
rect 1603 1522 1604 1526
rect 1598 1521 1604 1522
rect 1654 1526 1660 1527
rect 1670 1526 1676 1527
rect 1694 1528 1700 1529
rect 1654 1522 1655 1526
rect 1659 1522 1660 1526
rect 1694 1524 1695 1528
rect 1699 1524 1700 1528
rect 1694 1523 1700 1524
rect 1654 1521 1660 1522
rect 1478 1515 1484 1516
rect 1478 1511 1479 1515
rect 1483 1511 1484 1515
rect 1478 1510 1484 1511
rect 1638 1515 1644 1516
rect 1638 1511 1639 1515
rect 1643 1511 1644 1515
rect 1638 1510 1644 1511
rect 1694 1511 1700 1512
rect 1518 1509 1524 1510
rect 1518 1505 1519 1509
rect 1523 1505 1524 1509
rect 1518 1504 1524 1505
rect 1598 1509 1604 1510
rect 1598 1505 1599 1509
rect 1603 1505 1604 1509
rect 1598 1504 1604 1505
rect 1498 1503 1504 1504
rect 1498 1499 1499 1503
rect 1503 1499 1504 1503
rect 1520 1499 1522 1504
rect 1600 1499 1602 1504
rect 1479 1498 1483 1499
rect 1498 1498 1504 1499
rect 1519 1498 1523 1499
rect 1479 1493 1483 1494
rect 1480 1476 1482 1493
rect 1478 1475 1484 1476
rect 1478 1471 1479 1475
rect 1483 1471 1484 1475
rect 1478 1470 1484 1471
rect 1458 1467 1464 1468
rect 1458 1463 1459 1467
rect 1463 1463 1464 1467
rect 1458 1462 1464 1463
rect 1460 1416 1462 1462
rect 1478 1458 1484 1459
rect 1478 1454 1479 1458
rect 1483 1454 1484 1458
rect 1478 1453 1484 1454
rect 1480 1431 1482 1453
rect 1500 1452 1502 1498
rect 1519 1493 1523 1494
rect 1559 1498 1563 1499
rect 1559 1493 1563 1494
rect 1591 1498 1595 1499
rect 1591 1493 1595 1494
rect 1599 1498 1603 1499
rect 1599 1493 1603 1494
rect 1623 1498 1627 1499
rect 1623 1493 1627 1494
rect 1520 1476 1522 1493
rect 1560 1476 1562 1493
rect 1592 1476 1594 1493
rect 1624 1476 1626 1493
rect 1518 1475 1524 1476
rect 1518 1471 1519 1475
rect 1523 1471 1524 1475
rect 1518 1470 1524 1471
rect 1558 1475 1564 1476
rect 1558 1471 1559 1475
rect 1563 1471 1564 1475
rect 1558 1470 1564 1471
rect 1590 1475 1596 1476
rect 1590 1471 1591 1475
rect 1595 1471 1596 1475
rect 1590 1470 1596 1471
rect 1622 1475 1628 1476
rect 1622 1471 1623 1475
rect 1627 1471 1628 1475
rect 1622 1470 1628 1471
rect 1550 1467 1556 1468
rect 1550 1463 1551 1467
rect 1555 1463 1556 1467
rect 1550 1462 1556 1463
rect 1574 1467 1580 1468
rect 1574 1463 1575 1467
rect 1579 1463 1580 1467
rect 1574 1462 1580 1463
rect 1518 1458 1524 1459
rect 1518 1454 1519 1458
rect 1523 1454 1524 1458
rect 1518 1453 1524 1454
rect 1498 1451 1504 1452
rect 1498 1447 1499 1451
rect 1503 1447 1504 1451
rect 1498 1446 1504 1447
rect 1520 1431 1522 1453
rect 1479 1430 1483 1431
rect 1479 1425 1483 1426
rect 1519 1430 1523 1431
rect 1519 1425 1523 1426
rect 1535 1430 1539 1431
rect 1535 1425 1539 1426
rect 1470 1423 1476 1424
rect 1470 1419 1471 1423
rect 1475 1419 1476 1423
rect 1470 1418 1476 1419
rect 1458 1415 1464 1416
rect 1458 1411 1459 1415
rect 1463 1411 1464 1415
rect 1458 1410 1464 1411
rect 1472 1408 1474 1418
rect 1470 1407 1476 1408
rect 1470 1403 1471 1407
rect 1475 1403 1476 1407
rect 1470 1402 1476 1403
rect 1446 1379 1452 1380
rect 1446 1375 1447 1379
rect 1451 1375 1452 1379
rect 1446 1374 1452 1375
rect 1414 1373 1420 1374
rect 1414 1369 1415 1373
rect 1419 1369 1420 1373
rect 1414 1368 1420 1369
rect 1462 1372 1468 1373
rect 1462 1368 1463 1372
rect 1467 1368 1468 1372
rect 1416 1351 1418 1368
rect 1462 1367 1468 1368
rect 1464 1351 1466 1367
rect 1415 1350 1419 1351
rect 1415 1345 1419 1346
rect 1423 1350 1427 1351
rect 1423 1345 1427 1346
rect 1455 1350 1459 1351
rect 1455 1345 1459 1346
rect 1463 1350 1467 1351
rect 1463 1345 1467 1346
rect 1408 1340 1414 1342
rect 1302 1316 1303 1320
rect 1307 1316 1308 1320
rect 1302 1315 1308 1316
rect 1390 1319 1396 1320
rect 1390 1315 1391 1319
rect 1395 1315 1396 1319
rect 1390 1314 1396 1315
rect 1412 1312 1414 1340
rect 1424 1320 1426 1345
rect 1456 1321 1458 1345
rect 1454 1320 1460 1321
rect 1422 1319 1428 1320
rect 1422 1315 1423 1319
rect 1427 1315 1428 1319
rect 1454 1316 1455 1320
rect 1459 1316 1460 1320
rect 1454 1315 1460 1316
rect 1422 1314 1428 1315
rect 1286 1311 1292 1312
rect 1286 1307 1287 1311
rect 1291 1307 1292 1311
rect 1286 1306 1292 1307
rect 1410 1311 1416 1312
rect 1410 1307 1411 1311
rect 1415 1307 1416 1311
rect 1434 1311 1440 1312
rect 1434 1310 1435 1311
rect 1410 1306 1416 1307
rect 1432 1307 1435 1310
rect 1439 1307 1440 1311
rect 1432 1306 1440 1307
rect 1288 1284 1290 1306
rect 1302 1301 1308 1302
rect 1302 1297 1303 1301
rect 1307 1297 1308 1301
rect 1302 1296 1308 1297
rect 1390 1301 1396 1302
rect 1390 1297 1391 1301
rect 1395 1297 1396 1301
rect 1390 1296 1396 1297
rect 1286 1283 1292 1284
rect 1286 1279 1287 1283
rect 1291 1279 1292 1283
rect 1286 1278 1292 1279
rect 1304 1263 1306 1296
rect 1392 1263 1394 1296
rect 1412 1288 1414 1306
rect 1422 1302 1428 1303
rect 1422 1298 1423 1302
rect 1427 1298 1428 1302
rect 1422 1297 1428 1298
rect 1410 1287 1416 1288
rect 1410 1283 1411 1287
rect 1415 1283 1416 1287
rect 1410 1282 1416 1283
rect 1424 1263 1426 1297
rect 1255 1262 1259 1263
rect 1255 1257 1259 1258
rect 1295 1262 1299 1263
rect 1295 1257 1299 1258
rect 1303 1262 1307 1263
rect 1303 1257 1307 1258
rect 1343 1262 1347 1263
rect 1343 1257 1347 1258
rect 1375 1262 1379 1263
rect 1375 1257 1379 1258
rect 1391 1262 1395 1263
rect 1391 1257 1395 1258
rect 1407 1262 1411 1263
rect 1407 1257 1411 1258
rect 1423 1262 1427 1263
rect 1423 1257 1427 1258
rect 1214 1192 1220 1193
rect 1238 1195 1244 1196
rect 1256 1195 1258 1257
rect 1262 1207 1268 1208
rect 1262 1203 1263 1207
rect 1267 1203 1268 1207
rect 1262 1202 1268 1203
rect 1238 1191 1239 1195
rect 1243 1191 1244 1195
rect 1238 1190 1244 1191
rect 1254 1194 1260 1195
rect 1254 1190 1255 1194
rect 1259 1190 1260 1194
rect 1254 1189 1260 1190
rect 1254 1177 1260 1178
rect 1198 1176 1204 1177
rect 1198 1172 1199 1176
rect 1203 1172 1204 1176
rect 1254 1173 1255 1177
rect 1259 1173 1260 1177
rect 1254 1172 1260 1173
rect 1198 1171 1204 1172
rect 1200 1151 1202 1171
rect 1256 1151 1258 1172
rect 1199 1150 1203 1151
rect 1199 1145 1203 1146
rect 1247 1150 1251 1151
rect 1247 1145 1251 1146
rect 1255 1150 1259 1151
rect 1255 1145 1259 1146
rect 1248 1129 1250 1145
rect 1246 1128 1252 1129
rect 1246 1124 1247 1128
rect 1251 1124 1252 1128
rect 1246 1123 1252 1124
rect 1234 1115 1240 1116
rect 1234 1111 1235 1115
rect 1239 1111 1240 1115
rect 1234 1110 1240 1111
rect 1226 1107 1232 1108
rect 1226 1103 1227 1107
rect 1231 1103 1232 1107
rect 1226 1102 1232 1103
rect 1228 1076 1230 1102
rect 1194 1075 1200 1076
rect 1194 1071 1195 1075
rect 1199 1071 1200 1075
rect 1194 1070 1200 1071
rect 1226 1075 1232 1076
rect 1226 1071 1227 1075
rect 1231 1071 1232 1075
rect 1236 1072 1238 1110
rect 1246 1081 1252 1082
rect 1246 1077 1247 1081
rect 1251 1077 1252 1081
rect 1246 1076 1252 1077
rect 1264 1076 1266 1202
rect 1296 1198 1298 1257
rect 1294 1197 1300 1198
rect 1294 1193 1295 1197
rect 1299 1193 1300 1197
rect 1344 1195 1346 1257
rect 1350 1203 1356 1204
rect 1350 1199 1351 1203
rect 1355 1199 1356 1203
rect 1350 1198 1356 1199
rect 1294 1192 1300 1193
rect 1342 1194 1348 1195
rect 1342 1190 1343 1194
rect 1347 1190 1348 1194
rect 1342 1189 1348 1190
rect 1286 1183 1292 1184
rect 1286 1179 1287 1183
rect 1291 1179 1292 1183
rect 1286 1178 1292 1179
rect 1288 1164 1290 1178
rect 1342 1177 1348 1178
rect 1342 1173 1343 1177
rect 1347 1173 1348 1177
rect 1342 1172 1348 1173
rect 1310 1170 1316 1171
rect 1310 1166 1311 1170
rect 1315 1166 1316 1170
rect 1310 1165 1316 1166
rect 1286 1163 1292 1164
rect 1286 1159 1287 1163
rect 1291 1159 1292 1163
rect 1286 1158 1292 1159
rect 1312 1151 1314 1165
rect 1344 1151 1346 1172
rect 1287 1150 1291 1151
rect 1287 1145 1291 1146
rect 1311 1150 1315 1151
rect 1311 1145 1315 1146
rect 1335 1150 1339 1151
rect 1335 1145 1339 1146
rect 1343 1150 1347 1151
rect 1343 1145 1347 1146
rect 1288 1124 1290 1145
rect 1336 1127 1338 1145
rect 1334 1126 1340 1127
rect 1286 1123 1292 1124
rect 1286 1119 1287 1123
rect 1291 1119 1292 1123
rect 1334 1122 1335 1126
rect 1339 1122 1340 1126
rect 1334 1121 1340 1122
rect 1286 1118 1292 1119
rect 1278 1115 1284 1116
rect 1278 1111 1279 1115
rect 1283 1111 1284 1115
rect 1278 1110 1284 1111
rect 1226 1070 1232 1071
rect 1234 1071 1240 1072
rect 1196 1059 1198 1070
rect 1234 1067 1235 1071
rect 1239 1067 1240 1071
rect 1234 1066 1240 1067
rect 1192 1057 1198 1059
rect 1182 1015 1188 1016
rect 1182 1011 1183 1015
rect 1187 1011 1188 1015
rect 1182 1010 1188 1011
rect 1192 1008 1194 1057
rect 1248 1035 1250 1076
rect 1262 1075 1268 1076
rect 1262 1071 1263 1075
rect 1267 1071 1268 1075
rect 1262 1070 1268 1071
rect 1199 1034 1203 1035
rect 1199 1029 1203 1030
rect 1247 1034 1251 1035
rect 1247 1029 1251 1030
rect 1190 1007 1196 1008
rect 1190 1003 1191 1007
rect 1195 1003 1196 1007
rect 1200 1005 1202 1029
rect 1206 1011 1212 1012
rect 1206 1007 1207 1011
rect 1211 1007 1212 1011
rect 1206 1006 1212 1007
rect 1190 1002 1196 1003
rect 1198 1004 1204 1005
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1198 999 1204 1000
rect 1118 992 1124 993
rect 1166 994 1172 995
rect 1166 990 1167 994
rect 1171 990 1172 994
rect 1166 989 1172 990
rect 1208 988 1210 1006
rect 1248 998 1250 1029
rect 1264 1020 1266 1070
rect 1262 1019 1268 1020
rect 1262 1015 1263 1019
rect 1267 1015 1268 1019
rect 1262 1014 1268 1015
rect 1280 1008 1282 1110
rect 1286 1106 1292 1107
rect 1286 1102 1287 1106
rect 1291 1102 1292 1106
rect 1286 1101 1292 1102
rect 1288 1035 1290 1101
rect 1334 1085 1340 1086
rect 1334 1081 1335 1085
rect 1339 1081 1340 1085
rect 1334 1080 1340 1081
rect 1336 1035 1338 1080
rect 1352 1076 1354 1198
rect 1376 1195 1378 1257
rect 1408 1195 1410 1257
rect 1414 1207 1420 1208
rect 1414 1203 1415 1207
rect 1419 1203 1420 1207
rect 1414 1202 1420 1203
rect 1374 1194 1380 1195
rect 1374 1190 1375 1194
rect 1379 1190 1380 1194
rect 1374 1189 1380 1190
rect 1406 1194 1412 1195
rect 1406 1190 1407 1194
rect 1411 1190 1412 1194
rect 1406 1189 1412 1190
rect 1416 1184 1418 1202
rect 1423 1199 1429 1200
rect 1423 1195 1424 1199
rect 1428 1198 1429 1199
rect 1432 1198 1434 1306
rect 1438 1295 1444 1296
rect 1438 1291 1439 1295
rect 1443 1291 1444 1295
rect 1438 1290 1444 1291
rect 1454 1292 1460 1293
rect 1440 1288 1442 1290
rect 1454 1288 1455 1292
rect 1459 1288 1460 1292
rect 1438 1287 1444 1288
rect 1438 1283 1439 1287
rect 1443 1283 1444 1287
rect 1438 1282 1444 1283
rect 1446 1287 1452 1288
rect 1454 1287 1460 1288
rect 1446 1283 1447 1287
rect 1451 1283 1452 1287
rect 1446 1282 1452 1283
rect 1439 1262 1443 1263
rect 1439 1257 1443 1258
rect 1428 1196 1434 1198
rect 1428 1195 1429 1196
rect 1440 1195 1442 1257
rect 1448 1224 1450 1282
rect 1456 1263 1458 1287
rect 1472 1280 1474 1402
rect 1480 1394 1482 1425
rect 1478 1393 1484 1394
rect 1478 1389 1479 1393
rect 1483 1389 1484 1393
rect 1478 1388 1484 1389
rect 1486 1391 1492 1392
rect 1536 1391 1538 1425
rect 1552 1396 1554 1462
rect 1558 1458 1564 1459
rect 1558 1454 1559 1458
rect 1563 1454 1564 1458
rect 1558 1453 1564 1454
rect 1560 1431 1562 1453
rect 1559 1430 1563 1431
rect 1559 1425 1563 1426
rect 1576 1400 1578 1462
rect 1590 1458 1596 1459
rect 1590 1454 1591 1458
rect 1595 1454 1596 1458
rect 1590 1453 1596 1454
rect 1622 1458 1628 1459
rect 1622 1454 1623 1458
rect 1627 1454 1628 1458
rect 1622 1453 1628 1454
rect 1592 1431 1594 1453
rect 1624 1431 1626 1453
rect 1640 1452 1642 1510
rect 1654 1509 1660 1510
rect 1654 1505 1655 1509
rect 1659 1505 1660 1509
rect 1694 1507 1695 1511
rect 1699 1507 1700 1511
rect 1694 1506 1700 1507
rect 1654 1504 1660 1505
rect 1656 1499 1658 1504
rect 1696 1499 1698 1506
rect 1655 1498 1659 1499
rect 1655 1493 1659 1494
rect 1695 1498 1699 1499
rect 1695 1493 1699 1494
rect 1656 1476 1658 1493
rect 1654 1475 1660 1476
rect 1654 1471 1655 1475
rect 1659 1471 1660 1475
rect 1696 1474 1698 1493
rect 1654 1470 1660 1471
rect 1694 1473 1700 1474
rect 1694 1469 1695 1473
rect 1699 1469 1700 1473
rect 1694 1468 1700 1469
rect 1670 1467 1676 1468
rect 1670 1463 1671 1467
rect 1675 1463 1676 1467
rect 1670 1462 1676 1463
rect 1654 1458 1660 1459
rect 1654 1454 1655 1458
rect 1659 1454 1660 1458
rect 1654 1453 1660 1454
rect 1638 1451 1644 1452
rect 1638 1447 1639 1451
rect 1643 1447 1644 1451
rect 1638 1446 1644 1447
rect 1656 1431 1658 1453
rect 1672 1444 1674 1462
rect 1694 1456 1700 1457
rect 1694 1452 1695 1456
rect 1699 1452 1700 1456
rect 1694 1451 1700 1452
rect 1670 1443 1676 1444
rect 1670 1439 1671 1443
rect 1675 1439 1676 1443
rect 1670 1438 1676 1439
rect 1696 1431 1698 1451
rect 1704 1436 1706 1570
rect 1702 1435 1708 1436
rect 1702 1431 1703 1435
rect 1707 1431 1708 1435
rect 1583 1430 1587 1431
rect 1583 1425 1587 1426
rect 1591 1430 1595 1431
rect 1591 1425 1595 1426
rect 1623 1430 1627 1431
rect 1623 1425 1627 1426
rect 1655 1430 1659 1431
rect 1655 1425 1659 1426
rect 1695 1430 1699 1431
rect 1702 1430 1708 1431
rect 1695 1425 1699 1426
rect 1574 1399 1580 1400
rect 1550 1395 1556 1396
rect 1550 1391 1551 1395
rect 1555 1391 1556 1395
rect 1574 1395 1575 1399
rect 1579 1395 1580 1399
rect 1574 1394 1580 1395
rect 1584 1391 1586 1425
rect 1624 1391 1626 1425
rect 1656 1391 1658 1425
rect 1696 1393 1698 1425
rect 1694 1392 1700 1393
rect 1486 1387 1487 1391
rect 1491 1387 1492 1391
rect 1486 1386 1492 1387
rect 1534 1390 1540 1391
rect 1550 1390 1556 1391
rect 1582 1390 1588 1391
rect 1534 1386 1535 1390
rect 1539 1386 1540 1390
rect 1488 1356 1490 1386
rect 1534 1385 1540 1386
rect 1582 1386 1583 1390
rect 1587 1386 1588 1390
rect 1582 1385 1588 1386
rect 1622 1390 1628 1391
rect 1622 1386 1623 1390
rect 1627 1386 1628 1390
rect 1622 1385 1628 1386
rect 1654 1390 1660 1391
rect 1654 1386 1655 1390
rect 1659 1386 1660 1390
rect 1694 1388 1695 1392
rect 1699 1388 1700 1392
rect 1694 1387 1700 1388
rect 1654 1385 1660 1386
rect 1546 1379 1552 1380
rect 1546 1375 1547 1379
rect 1551 1375 1552 1379
rect 1546 1374 1552 1375
rect 1694 1375 1700 1376
rect 1534 1373 1540 1374
rect 1534 1369 1535 1373
rect 1539 1369 1540 1373
rect 1534 1368 1540 1369
rect 1486 1355 1492 1356
rect 1486 1351 1487 1355
rect 1491 1351 1492 1355
rect 1536 1351 1538 1368
rect 1486 1350 1492 1351
rect 1495 1350 1499 1351
rect 1495 1345 1499 1346
rect 1527 1350 1531 1351
rect 1527 1345 1531 1346
rect 1535 1350 1539 1351
rect 1535 1345 1539 1346
rect 1496 1320 1498 1345
rect 1528 1320 1530 1345
rect 1494 1319 1500 1320
rect 1494 1315 1495 1319
rect 1499 1315 1500 1319
rect 1494 1314 1500 1315
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1482 1311 1488 1312
rect 1482 1307 1483 1311
rect 1487 1307 1488 1311
rect 1482 1306 1488 1307
rect 1538 1311 1544 1312
rect 1538 1307 1539 1311
rect 1543 1307 1544 1311
rect 1538 1306 1544 1307
rect 1484 1284 1486 1306
rect 1494 1302 1500 1303
rect 1494 1298 1495 1302
rect 1499 1298 1500 1302
rect 1494 1297 1500 1298
rect 1526 1302 1532 1303
rect 1526 1298 1527 1302
rect 1531 1298 1532 1302
rect 1526 1297 1532 1298
rect 1482 1283 1488 1284
rect 1470 1279 1476 1280
rect 1470 1275 1471 1279
rect 1475 1275 1476 1279
rect 1482 1279 1483 1283
rect 1487 1279 1488 1283
rect 1482 1278 1488 1279
rect 1470 1274 1476 1275
rect 1496 1263 1498 1297
rect 1514 1295 1520 1296
rect 1514 1291 1515 1295
rect 1519 1291 1520 1295
rect 1514 1290 1520 1291
rect 1516 1277 1518 1290
rect 1515 1276 1519 1277
rect 1515 1271 1519 1272
rect 1528 1263 1530 1297
rect 1455 1262 1459 1263
rect 1455 1257 1459 1258
rect 1479 1262 1483 1263
rect 1479 1257 1483 1258
rect 1495 1262 1499 1263
rect 1495 1257 1499 1258
rect 1519 1262 1523 1263
rect 1519 1257 1523 1258
rect 1527 1262 1531 1263
rect 1527 1257 1531 1258
rect 1446 1223 1452 1224
rect 1446 1219 1447 1223
rect 1451 1219 1452 1223
rect 1446 1218 1452 1219
rect 1423 1194 1429 1195
rect 1438 1194 1444 1195
rect 1438 1190 1439 1194
rect 1443 1190 1444 1194
rect 1438 1189 1444 1190
rect 1416 1183 1424 1184
rect 1416 1180 1419 1183
rect 1418 1179 1419 1180
rect 1423 1179 1424 1183
rect 1418 1178 1424 1179
rect 1374 1177 1380 1178
rect 1374 1173 1375 1177
rect 1379 1173 1380 1177
rect 1374 1172 1380 1173
rect 1406 1177 1412 1178
rect 1406 1173 1407 1177
rect 1411 1173 1412 1177
rect 1406 1172 1412 1173
rect 1438 1177 1444 1178
rect 1438 1173 1439 1177
rect 1443 1173 1444 1177
rect 1438 1172 1444 1173
rect 1448 1172 1450 1218
rect 1454 1215 1460 1216
rect 1454 1211 1455 1215
rect 1459 1211 1460 1215
rect 1454 1210 1460 1211
rect 1456 1184 1458 1210
rect 1480 1195 1482 1257
rect 1498 1199 1504 1200
rect 1498 1195 1499 1199
rect 1503 1195 1504 1199
rect 1520 1195 1522 1257
rect 1540 1200 1542 1306
rect 1548 1296 1550 1374
rect 1582 1373 1588 1374
rect 1582 1369 1583 1373
rect 1587 1369 1588 1373
rect 1582 1368 1588 1369
rect 1622 1373 1628 1374
rect 1622 1369 1623 1373
rect 1627 1369 1628 1373
rect 1622 1368 1628 1369
rect 1654 1373 1660 1374
rect 1654 1369 1655 1373
rect 1659 1369 1660 1373
rect 1694 1371 1695 1375
rect 1699 1371 1700 1375
rect 1694 1370 1700 1371
rect 1654 1368 1660 1369
rect 1574 1367 1580 1368
rect 1574 1363 1575 1367
rect 1579 1363 1580 1367
rect 1574 1362 1580 1363
rect 1559 1350 1563 1351
rect 1559 1345 1563 1346
rect 1560 1320 1562 1345
rect 1558 1319 1564 1320
rect 1558 1315 1559 1319
rect 1563 1315 1564 1319
rect 1558 1314 1564 1315
rect 1558 1302 1564 1303
rect 1558 1298 1559 1302
rect 1563 1298 1564 1302
rect 1558 1297 1564 1298
rect 1546 1295 1552 1296
rect 1546 1291 1547 1295
rect 1551 1291 1552 1295
rect 1546 1290 1552 1291
rect 1560 1263 1562 1297
rect 1576 1296 1578 1362
rect 1584 1351 1586 1368
rect 1624 1351 1626 1368
rect 1656 1351 1658 1368
rect 1696 1351 1698 1370
rect 1583 1350 1587 1351
rect 1583 1345 1587 1346
rect 1591 1350 1595 1351
rect 1591 1345 1595 1346
rect 1623 1350 1627 1351
rect 1623 1345 1627 1346
rect 1655 1350 1659 1351
rect 1655 1345 1659 1346
rect 1695 1350 1699 1351
rect 1695 1345 1699 1346
rect 1592 1320 1594 1345
rect 1624 1320 1626 1345
rect 1656 1320 1658 1345
rect 1590 1319 1596 1320
rect 1590 1315 1591 1319
rect 1595 1315 1596 1319
rect 1590 1314 1596 1315
rect 1622 1319 1628 1320
rect 1622 1315 1623 1319
rect 1627 1315 1628 1319
rect 1622 1314 1628 1315
rect 1654 1319 1660 1320
rect 1654 1315 1655 1319
rect 1659 1315 1660 1319
rect 1696 1318 1698 1345
rect 1654 1314 1660 1315
rect 1694 1317 1700 1318
rect 1694 1313 1695 1317
rect 1699 1313 1700 1317
rect 1694 1312 1700 1313
rect 1670 1311 1676 1312
rect 1670 1307 1671 1311
rect 1675 1307 1676 1311
rect 1670 1306 1676 1307
rect 1590 1302 1596 1303
rect 1590 1298 1591 1302
rect 1595 1298 1596 1302
rect 1590 1297 1596 1298
rect 1622 1302 1628 1303
rect 1622 1298 1623 1302
rect 1627 1298 1628 1302
rect 1622 1297 1628 1298
rect 1654 1302 1660 1303
rect 1654 1298 1655 1302
rect 1659 1298 1660 1302
rect 1654 1297 1660 1298
rect 1574 1295 1580 1296
rect 1574 1291 1575 1295
rect 1579 1291 1580 1295
rect 1574 1290 1580 1291
rect 1592 1263 1594 1297
rect 1624 1263 1626 1297
rect 1656 1263 1658 1297
rect 1559 1262 1563 1263
rect 1559 1257 1563 1258
rect 1591 1262 1595 1263
rect 1591 1257 1595 1258
rect 1623 1262 1627 1263
rect 1623 1257 1627 1258
rect 1655 1262 1659 1263
rect 1655 1257 1659 1258
rect 1546 1203 1552 1204
rect 1538 1199 1544 1200
rect 1538 1195 1539 1199
rect 1543 1195 1544 1199
rect 1546 1199 1547 1203
rect 1551 1199 1552 1203
rect 1546 1198 1552 1199
rect 1478 1194 1484 1195
rect 1498 1194 1504 1195
rect 1518 1194 1524 1195
rect 1538 1194 1544 1195
rect 1478 1190 1479 1194
rect 1483 1190 1484 1194
rect 1478 1189 1484 1190
rect 1454 1183 1460 1184
rect 1454 1179 1455 1183
rect 1459 1179 1460 1183
rect 1454 1178 1460 1179
rect 1478 1177 1484 1178
rect 1478 1173 1479 1177
rect 1483 1173 1484 1177
rect 1478 1172 1484 1173
rect 1376 1151 1378 1172
rect 1408 1151 1410 1172
rect 1430 1171 1436 1172
rect 1430 1167 1431 1171
rect 1435 1167 1436 1171
rect 1430 1166 1436 1167
rect 1375 1150 1379 1151
rect 1375 1145 1379 1146
rect 1407 1150 1411 1151
rect 1407 1145 1411 1146
rect 1423 1150 1427 1151
rect 1423 1145 1427 1146
rect 1424 1124 1426 1145
rect 1422 1123 1428 1124
rect 1422 1119 1423 1123
rect 1427 1119 1428 1123
rect 1422 1118 1428 1119
rect 1422 1106 1428 1107
rect 1422 1102 1423 1106
rect 1427 1102 1428 1106
rect 1422 1101 1428 1102
rect 1350 1075 1356 1076
rect 1350 1071 1351 1075
rect 1355 1071 1356 1075
rect 1350 1070 1356 1071
rect 1424 1035 1426 1101
rect 1432 1100 1434 1166
rect 1440 1151 1442 1172
rect 1446 1171 1452 1172
rect 1446 1167 1447 1171
rect 1451 1167 1452 1171
rect 1446 1166 1452 1167
rect 1480 1151 1482 1172
rect 1439 1150 1443 1151
rect 1439 1145 1443 1146
rect 1455 1150 1459 1151
rect 1455 1145 1459 1146
rect 1479 1150 1483 1151
rect 1479 1145 1483 1146
rect 1487 1150 1491 1151
rect 1487 1145 1491 1146
rect 1456 1124 1458 1145
rect 1488 1124 1490 1145
rect 1454 1123 1460 1124
rect 1454 1119 1455 1123
rect 1459 1119 1460 1123
rect 1454 1118 1460 1119
rect 1486 1123 1492 1124
rect 1486 1119 1487 1123
rect 1491 1119 1492 1123
rect 1486 1118 1492 1119
rect 1500 1116 1502 1194
rect 1518 1190 1519 1194
rect 1523 1190 1524 1194
rect 1518 1189 1524 1190
rect 1548 1184 1550 1198
rect 1560 1195 1562 1257
rect 1592 1195 1594 1257
rect 1624 1195 1626 1257
rect 1656 1195 1658 1257
rect 1672 1200 1674 1306
rect 1694 1300 1700 1301
rect 1694 1296 1695 1300
rect 1699 1296 1700 1300
rect 1694 1295 1700 1296
rect 1696 1263 1698 1295
rect 1695 1262 1699 1263
rect 1695 1257 1699 1258
rect 1670 1199 1676 1200
rect 1670 1195 1671 1199
rect 1675 1195 1676 1199
rect 1696 1197 1698 1257
rect 1558 1194 1564 1195
rect 1558 1190 1559 1194
rect 1563 1190 1564 1194
rect 1558 1189 1564 1190
rect 1590 1194 1596 1195
rect 1590 1190 1591 1194
rect 1595 1190 1596 1194
rect 1590 1189 1596 1190
rect 1622 1194 1628 1195
rect 1622 1190 1623 1194
rect 1627 1190 1628 1194
rect 1622 1189 1628 1190
rect 1654 1194 1660 1195
rect 1670 1194 1676 1195
rect 1694 1196 1700 1197
rect 1654 1190 1655 1194
rect 1659 1190 1660 1194
rect 1694 1192 1695 1196
rect 1699 1192 1700 1196
rect 1694 1191 1700 1192
rect 1654 1189 1660 1190
rect 1546 1183 1552 1184
rect 1546 1179 1547 1183
rect 1551 1179 1552 1183
rect 1546 1178 1552 1179
rect 1574 1183 1580 1184
rect 1574 1179 1575 1183
rect 1579 1179 1580 1183
rect 1574 1178 1580 1179
rect 1610 1183 1616 1184
rect 1610 1179 1611 1183
rect 1615 1179 1616 1183
rect 1610 1178 1616 1179
rect 1694 1179 1700 1180
rect 1518 1177 1524 1178
rect 1518 1173 1519 1177
rect 1523 1173 1524 1177
rect 1518 1172 1524 1173
rect 1558 1177 1564 1178
rect 1558 1173 1559 1177
rect 1563 1173 1564 1177
rect 1558 1172 1564 1173
rect 1520 1151 1522 1172
rect 1560 1151 1562 1172
rect 1519 1150 1523 1151
rect 1519 1145 1523 1146
rect 1559 1150 1563 1151
rect 1559 1145 1563 1146
rect 1520 1124 1522 1145
rect 1560 1124 1562 1145
rect 1518 1123 1524 1124
rect 1518 1119 1519 1123
rect 1523 1119 1524 1123
rect 1518 1118 1524 1119
rect 1558 1123 1564 1124
rect 1558 1119 1559 1123
rect 1563 1119 1564 1123
rect 1558 1118 1564 1119
rect 1470 1115 1476 1116
rect 1470 1111 1471 1115
rect 1475 1111 1476 1115
rect 1470 1110 1476 1111
rect 1498 1115 1504 1116
rect 1498 1111 1499 1115
rect 1503 1111 1504 1115
rect 1498 1110 1504 1111
rect 1534 1115 1540 1116
rect 1534 1111 1535 1115
rect 1539 1111 1540 1115
rect 1534 1110 1540 1111
rect 1454 1106 1460 1107
rect 1454 1102 1455 1106
rect 1459 1102 1460 1106
rect 1454 1101 1460 1102
rect 1430 1099 1436 1100
rect 1430 1095 1431 1099
rect 1435 1095 1436 1099
rect 1430 1094 1436 1095
rect 1446 1075 1452 1076
rect 1446 1071 1447 1075
rect 1451 1071 1452 1075
rect 1446 1070 1452 1071
rect 1287 1034 1291 1035
rect 1287 1029 1291 1030
rect 1295 1034 1299 1035
rect 1295 1029 1299 1030
rect 1327 1034 1331 1035
rect 1327 1029 1331 1030
rect 1335 1034 1339 1035
rect 1335 1029 1339 1030
rect 1367 1034 1371 1035
rect 1367 1029 1371 1030
rect 1407 1034 1411 1035
rect 1407 1029 1411 1030
rect 1423 1034 1427 1035
rect 1423 1029 1427 1030
rect 1439 1034 1443 1035
rect 1439 1029 1443 1030
rect 1278 1007 1284 1008
rect 1278 1003 1279 1007
rect 1283 1003 1284 1007
rect 1278 1002 1284 1003
rect 1246 997 1252 998
rect 1246 993 1247 997
rect 1251 993 1252 997
rect 1296 995 1298 1029
rect 1328 1005 1330 1029
rect 1334 1011 1340 1012
rect 1334 1007 1335 1011
rect 1339 1007 1340 1011
rect 1334 1006 1340 1007
rect 1326 1004 1332 1005
rect 1326 1000 1327 1004
rect 1331 1000 1332 1004
rect 1326 999 1332 1000
rect 1246 992 1252 993
rect 1294 994 1300 995
rect 1294 990 1295 994
rect 1299 990 1300 994
rect 1294 989 1300 990
rect 1336 988 1338 1006
rect 1368 1005 1370 1029
rect 1366 1004 1372 1005
rect 1366 1000 1367 1004
rect 1371 1000 1372 1004
rect 1366 999 1372 1000
rect 1408 995 1410 1029
rect 1440 995 1442 1029
rect 1406 994 1412 995
rect 1382 991 1388 992
rect 1206 987 1212 988
rect 1206 983 1207 987
rect 1211 983 1212 987
rect 1206 982 1212 983
rect 1334 987 1340 988
rect 1334 983 1335 987
rect 1339 983 1340 987
rect 1382 987 1383 991
rect 1387 987 1388 991
rect 1406 990 1407 994
rect 1411 990 1412 994
rect 1406 989 1412 990
rect 1438 994 1444 995
rect 1438 990 1439 994
rect 1443 990 1444 994
rect 1438 989 1444 990
rect 1382 986 1388 987
rect 1334 982 1340 983
rect 1166 977 1172 978
rect 1294 977 1300 978
rect 1166 973 1167 977
rect 1171 973 1172 977
rect 1166 972 1172 973
rect 1198 976 1204 977
rect 1198 972 1199 976
rect 1203 972 1204 976
rect 1294 973 1295 977
rect 1299 973 1300 977
rect 1294 972 1300 973
rect 1326 976 1332 977
rect 1326 972 1327 976
rect 1331 972 1332 976
rect 1112 969 1126 971
rect 1082 963 1088 964
rect 1082 959 1083 963
rect 1087 959 1088 963
rect 1082 958 1088 959
rect 1063 954 1067 955
rect 1063 949 1067 950
rect 1071 954 1075 955
rect 1071 949 1075 950
rect 1111 954 1115 955
rect 1111 949 1115 950
rect 1072 925 1074 949
rect 1070 924 1076 925
rect 1112 924 1114 949
rect 1124 936 1126 969
rect 1134 970 1140 971
rect 1134 966 1135 970
rect 1139 966 1140 970
rect 1134 965 1140 966
rect 1136 955 1138 965
rect 1168 955 1170 972
rect 1198 971 1204 972
rect 1200 955 1202 971
rect 1262 970 1268 971
rect 1262 966 1263 970
rect 1267 966 1268 970
rect 1262 965 1268 966
rect 1264 955 1266 965
rect 1296 955 1298 972
rect 1326 971 1332 972
rect 1366 976 1372 977
rect 1366 972 1367 976
rect 1371 972 1372 976
rect 1366 971 1372 972
rect 1328 955 1330 971
rect 1368 955 1370 971
rect 1135 954 1139 955
rect 1135 949 1139 950
rect 1143 954 1147 955
rect 1143 949 1147 950
rect 1167 954 1171 955
rect 1167 949 1171 950
rect 1199 954 1203 955
rect 1199 949 1203 950
rect 1239 954 1243 955
rect 1239 949 1243 950
rect 1263 954 1267 955
rect 1263 949 1267 950
rect 1271 954 1275 955
rect 1271 949 1275 950
rect 1295 954 1299 955
rect 1295 949 1299 950
rect 1327 954 1331 955
rect 1327 949 1331 950
rect 1367 954 1371 955
rect 1367 949 1371 950
rect 1122 935 1128 936
rect 1122 931 1123 935
rect 1127 931 1128 935
rect 1122 930 1128 931
rect 1070 920 1071 924
rect 1075 920 1076 924
rect 1070 919 1076 920
rect 1110 923 1116 924
rect 1110 919 1111 923
rect 1115 919 1116 923
rect 1110 918 1116 919
rect 1094 915 1100 916
rect 1094 911 1095 915
rect 1099 911 1100 915
rect 1094 910 1100 911
rect 1070 896 1076 897
rect 1070 892 1071 896
rect 1075 892 1076 896
rect 1070 891 1076 892
rect 1046 887 1052 888
rect 1046 883 1047 887
rect 1051 883 1052 887
rect 1046 882 1052 883
rect 1072 839 1074 891
rect 1096 888 1098 910
rect 1110 905 1116 906
rect 1110 901 1111 905
rect 1115 901 1116 905
rect 1110 900 1116 901
rect 1078 887 1084 888
rect 1078 883 1079 887
rect 1083 883 1084 887
rect 1078 882 1084 883
rect 1094 887 1100 888
rect 1094 883 1095 887
rect 1099 883 1100 887
rect 1094 882 1100 883
rect 999 838 1003 839
rect 999 833 1003 834
rect 1031 838 1035 839
rect 1031 833 1035 834
rect 1039 838 1043 839
rect 1039 833 1043 834
rect 1071 838 1075 839
rect 1071 833 1075 834
rect 990 823 996 824
rect 990 819 991 823
rect 995 819 996 823
rect 990 818 996 819
rect 950 807 956 808
rect 950 803 951 807
rect 955 803 956 807
rect 1032 806 1034 833
rect 1055 812 1059 813
rect 1055 807 1059 808
rect 950 802 956 803
rect 1030 805 1036 806
rect 1030 801 1031 805
rect 1035 801 1036 805
rect 1056 804 1058 807
rect 1030 800 1036 801
rect 1042 803 1048 804
rect 1042 799 1043 803
rect 1047 799 1048 803
rect 1042 798 1048 799
rect 1054 803 1060 804
rect 1054 799 1055 803
rect 1059 799 1060 803
rect 1054 798 1060 799
rect 950 784 956 785
rect 950 780 951 784
rect 955 780 956 784
rect 950 779 956 780
rect 1014 784 1020 785
rect 1014 780 1015 784
rect 1019 780 1020 784
rect 1014 779 1020 780
rect 952 755 954 779
rect 1016 755 1018 779
rect 1034 775 1040 776
rect 1034 771 1035 775
rect 1039 771 1040 775
rect 1034 770 1040 771
rect 863 754 867 755
rect 863 749 867 750
rect 911 754 915 755
rect 911 749 915 750
rect 951 754 955 755
rect 951 749 955 750
rect 999 754 1003 755
rect 999 749 1003 750
rect 1015 754 1019 755
rect 1015 749 1019 750
rect 864 728 866 749
rect 912 731 914 749
rect 1000 736 1002 749
rect 998 735 1004 736
rect 998 731 999 735
rect 1003 731 1004 735
rect 910 730 916 731
rect 998 730 1004 731
rect 862 727 868 728
rect 862 723 863 727
rect 867 723 868 727
rect 910 726 911 730
rect 915 726 916 730
rect 910 725 916 726
rect 862 722 868 723
rect 862 710 868 711
rect 862 706 863 710
rect 867 706 868 710
rect 862 705 868 706
rect 850 691 856 692
rect 850 687 851 691
rect 855 687 856 691
rect 850 686 856 687
rect 842 667 848 668
rect 842 663 843 667
rect 847 663 848 667
rect 852 664 854 686
rect 842 662 848 663
rect 850 663 856 664
rect 850 659 851 663
rect 855 659 856 663
rect 850 658 856 659
rect 766 623 772 624
rect 766 619 767 623
rect 771 619 772 623
rect 766 618 772 619
rect 830 623 836 624
rect 830 619 831 623
rect 835 619 836 623
rect 830 618 836 619
rect 758 615 764 616
rect 758 611 759 615
rect 763 611 764 615
rect 758 610 764 611
rect 730 607 736 608
rect 730 603 731 607
rect 735 603 736 607
rect 730 602 736 603
rect 686 591 692 592
rect 686 587 687 591
rect 691 587 692 591
rect 686 586 692 587
rect 670 585 676 586
rect 670 581 671 585
rect 675 581 676 585
rect 670 580 676 581
rect 766 582 772 583
rect 672 563 674 580
rect 766 578 767 582
rect 771 578 772 582
rect 766 577 772 578
rect 768 563 770 577
rect 794 563 800 564
rect 647 562 651 563
rect 647 557 651 558
rect 671 562 675 563
rect 671 557 675 558
rect 727 562 731 563
rect 727 557 731 558
rect 767 562 771 563
rect 767 557 771 558
rect 775 562 779 563
rect 794 559 795 563
rect 799 559 800 563
rect 794 558 800 559
rect 775 557 779 558
rect 648 537 650 557
rect 728 541 730 557
rect 726 540 732 541
rect 646 536 652 537
rect 646 532 647 536
rect 651 532 652 536
rect 726 536 727 540
rect 731 536 732 540
rect 776 537 778 557
rect 726 535 732 536
rect 774 536 780 537
rect 634 531 640 532
rect 646 531 652 532
rect 774 532 775 536
rect 779 532 780 536
rect 774 531 780 532
rect 634 527 635 531
rect 639 527 640 531
rect 634 526 640 527
rect 714 527 720 528
rect 714 523 715 527
rect 719 523 720 527
rect 714 522 720 523
rect 610 503 616 504
rect 610 499 611 503
rect 615 499 616 503
rect 610 498 616 499
rect 654 498 660 499
rect 566 483 572 484
rect 566 479 567 483
rect 571 479 572 483
rect 566 478 572 479
rect 612 468 614 498
rect 654 494 655 498
rect 659 494 660 498
rect 654 493 660 494
rect 626 491 632 492
rect 626 487 627 491
rect 631 487 632 491
rect 626 486 632 487
rect 642 487 648 488
rect 610 467 616 468
rect 610 463 611 467
rect 615 463 616 467
rect 610 462 616 463
rect 534 459 540 460
rect 534 455 535 459
rect 539 455 540 459
rect 534 454 540 455
rect 526 403 532 404
rect 526 399 527 403
rect 531 399 532 403
rect 526 398 532 399
rect 518 379 524 380
rect 486 377 492 378
rect 414 374 420 375
rect 390 371 396 372
rect 354 367 360 368
rect 354 363 355 367
rect 359 363 360 367
rect 390 367 391 371
rect 395 367 396 371
rect 414 370 415 374
rect 419 370 420 374
rect 414 369 420 370
rect 446 374 452 375
rect 446 370 447 374
rect 451 370 452 374
rect 486 373 487 377
rect 491 373 492 377
rect 518 375 519 379
rect 523 375 524 379
rect 518 374 524 375
rect 486 372 492 373
rect 446 369 452 370
rect 390 366 396 367
rect 354 362 360 363
rect 430 363 436 364
rect 252 360 258 362
rect 252 359 253 360
rect 247 358 253 359
rect 430 359 431 363
rect 435 359 436 363
rect 430 358 436 359
rect 110 354 116 355
rect 134 357 140 358
rect 112 323 114 354
rect 134 353 135 357
rect 139 353 140 357
rect 134 352 140 353
rect 166 357 172 358
rect 166 353 167 357
rect 171 353 172 357
rect 166 352 172 353
rect 198 357 204 358
rect 198 353 199 357
rect 203 353 204 357
rect 198 352 204 353
rect 230 357 236 358
rect 230 353 231 357
rect 235 353 236 357
rect 230 352 236 353
rect 262 357 268 358
rect 414 357 420 358
rect 262 353 263 357
rect 267 353 268 357
rect 262 352 268 353
rect 294 356 300 357
rect 294 352 295 356
rect 299 352 300 356
rect 414 353 415 357
rect 419 353 420 357
rect 136 323 138 352
rect 154 351 160 352
rect 154 347 155 351
rect 159 347 160 351
rect 154 346 160 347
rect 111 322 115 323
rect 111 317 115 318
rect 135 322 139 323
rect 135 317 139 318
rect 83 308 87 309
rect 83 303 87 304
rect 84 284 86 303
rect 112 302 114 317
rect 136 304 138 317
rect 134 303 140 304
rect 110 301 116 302
rect 110 297 111 301
rect 115 297 116 301
rect 134 299 135 303
rect 139 299 140 303
rect 134 298 140 299
rect 110 296 116 297
rect 134 286 140 287
rect 110 284 116 285
rect 82 283 88 284
rect 82 279 83 283
rect 87 279 88 283
rect 110 280 111 284
rect 115 280 116 284
rect 134 282 135 286
rect 139 282 140 286
rect 134 281 140 282
rect 110 279 116 280
rect 82 278 88 279
rect 112 251 114 279
rect 136 251 138 281
rect 156 280 158 346
rect 168 323 170 352
rect 200 323 202 352
rect 232 323 234 352
rect 264 323 266 352
rect 294 351 300 352
rect 374 352 380 353
rect 414 352 420 353
rect 296 323 298 351
rect 374 348 375 352
rect 379 348 380 352
rect 374 347 380 348
rect 376 323 378 347
rect 416 323 418 352
rect 167 322 171 323
rect 167 317 171 318
rect 199 322 203 323
rect 199 317 203 318
rect 231 322 235 323
rect 231 317 235 318
rect 263 322 267 323
rect 263 317 267 318
rect 295 322 299 323
rect 295 317 299 318
rect 327 322 331 323
rect 327 317 331 318
rect 359 322 363 323
rect 359 317 363 318
rect 375 322 379 323
rect 375 317 379 318
rect 391 322 395 323
rect 391 317 395 318
rect 415 322 419 323
rect 415 317 419 318
rect 423 322 427 323
rect 423 317 427 318
rect 168 304 170 317
rect 200 304 202 317
rect 232 304 234 317
rect 264 304 266 317
rect 296 304 298 317
rect 328 304 330 317
rect 360 304 362 317
rect 392 304 394 317
rect 424 304 426 317
rect 166 303 172 304
rect 166 299 167 303
rect 171 299 172 303
rect 166 298 172 299
rect 198 303 204 304
rect 198 299 199 303
rect 203 299 204 303
rect 198 298 204 299
rect 230 303 236 304
rect 230 299 231 303
rect 235 299 236 303
rect 230 298 236 299
rect 262 303 268 304
rect 262 299 263 303
rect 267 299 268 303
rect 262 298 268 299
rect 294 303 300 304
rect 294 299 295 303
rect 299 299 300 303
rect 294 298 300 299
rect 326 303 332 304
rect 326 299 327 303
rect 331 299 332 303
rect 326 298 332 299
rect 358 303 364 304
rect 358 299 359 303
rect 363 299 364 303
rect 358 298 364 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 422 303 428 304
rect 422 299 423 303
rect 427 299 428 303
rect 422 298 428 299
rect 274 295 280 296
rect 274 291 275 295
rect 279 291 280 295
rect 274 290 280 291
rect 166 286 172 287
rect 166 282 167 286
rect 171 282 172 286
rect 166 281 172 282
rect 198 286 204 287
rect 198 282 199 286
rect 203 282 204 286
rect 198 281 204 282
rect 230 286 236 287
rect 230 282 231 286
rect 235 282 236 286
rect 230 281 236 282
rect 262 286 268 287
rect 262 282 263 286
rect 267 282 268 286
rect 262 281 268 282
rect 154 279 160 280
rect 154 275 155 279
rect 159 275 160 279
rect 154 274 160 275
rect 168 251 170 281
rect 200 251 202 281
rect 232 251 234 281
rect 264 251 266 281
rect 276 275 278 290
rect 294 286 300 287
rect 294 282 295 286
rect 299 282 300 286
rect 294 281 300 282
rect 326 286 332 287
rect 326 282 327 286
rect 331 282 332 286
rect 326 281 332 282
rect 358 286 364 287
rect 358 282 359 286
rect 363 282 364 286
rect 358 281 364 282
rect 390 286 396 287
rect 390 282 391 286
rect 395 282 396 286
rect 390 281 396 282
rect 422 286 428 287
rect 422 282 423 286
rect 427 282 428 286
rect 422 281 428 282
rect 272 273 278 275
rect 111 250 115 251
rect 111 245 115 246
rect 135 250 139 251
rect 135 245 139 246
rect 167 250 171 251
rect 167 245 171 246
rect 183 250 187 251
rect 183 245 187 246
rect 199 250 203 251
rect 199 245 203 246
rect 215 250 219 251
rect 215 245 219 246
rect 231 250 235 251
rect 231 245 235 246
rect 247 250 251 251
rect 247 245 251 246
rect 263 250 267 251
rect 263 245 267 246
rect 112 217 114 245
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 184 215 186 245
rect 216 215 218 245
rect 248 215 250 245
rect 272 228 274 273
rect 296 251 298 281
rect 328 251 330 281
rect 360 251 362 281
rect 366 279 372 280
rect 366 275 367 279
rect 371 275 372 279
rect 366 274 372 275
rect 279 250 283 251
rect 279 245 283 246
rect 295 250 299 251
rect 295 245 299 246
rect 311 250 315 251
rect 311 245 315 246
rect 327 250 331 251
rect 327 245 331 246
rect 343 250 347 251
rect 343 245 347 246
rect 359 250 363 251
rect 359 245 363 246
rect 270 227 276 228
rect 270 223 271 227
rect 275 223 276 227
rect 270 222 276 223
rect 280 215 282 245
rect 312 215 314 245
rect 330 227 336 228
rect 330 223 331 227
rect 335 223 336 227
rect 330 222 336 223
rect 110 211 116 212
rect 182 214 188 215
rect 182 210 183 214
rect 187 210 188 214
rect 182 209 188 210
rect 214 214 220 215
rect 214 210 215 214
rect 219 210 220 214
rect 214 209 220 210
rect 246 214 252 215
rect 246 210 247 214
rect 251 210 252 214
rect 246 209 252 210
rect 278 214 284 215
rect 278 210 279 214
rect 283 210 284 214
rect 278 209 284 210
rect 310 214 316 215
rect 310 210 311 214
rect 315 210 316 214
rect 310 209 316 210
rect 332 204 334 222
rect 344 215 346 245
rect 358 219 364 220
rect 358 215 359 219
rect 363 215 364 219
rect 342 214 348 215
rect 358 214 364 215
rect 342 210 343 214
rect 347 210 348 214
rect 342 209 348 210
rect 330 203 336 204
rect 110 199 116 200
rect 110 195 111 199
rect 115 195 116 199
rect 330 199 331 203
rect 335 199 336 203
rect 330 198 336 199
rect 110 194 116 195
rect 182 197 188 198
rect 112 175 114 194
rect 182 193 183 197
rect 187 193 188 197
rect 182 192 188 193
rect 214 197 220 198
rect 214 193 215 197
rect 219 193 220 197
rect 214 192 220 193
rect 246 197 252 198
rect 246 193 247 197
rect 251 193 252 197
rect 246 192 252 193
rect 278 197 284 198
rect 278 193 279 197
rect 283 193 284 197
rect 278 192 284 193
rect 310 197 316 198
rect 310 193 311 197
rect 315 193 316 197
rect 310 192 316 193
rect 342 197 348 198
rect 342 193 343 197
rect 347 193 348 197
rect 342 192 348 193
rect 360 192 362 214
rect 368 212 370 274
rect 392 251 394 281
rect 424 251 426 281
rect 432 280 434 358
rect 446 357 452 358
rect 446 353 447 357
rect 451 353 452 357
rect 446 352 452 353
rect 448 323 450 352
rect 502 350 508 351
rect 502 346 503 350
rect 507 346 508 350
rect 502 345 508 346
rect 504 323 506 345
rect 520 332 522 374
rect 528 372 530 398
rect 536 392 538 454
rect 606 451 612 452
rect 606 447 607 451
rect 611 447 612 451
rect 606 446 612 447
rect 550 443 556 444
rect 543 442 547 443
rect 550 439 551 443
rect 555 439 556 443
rect 550 438 556 439
rect 543 437 547 438
rect 544 395 546 437
rect 552 424 554 438
rect 550 423 556 424
rect 550 419 551 423
rect 555 419 556 423
rect 550 418 556 419
rect 552 404 554 418
rect 594 407 600 408
rect 550 403 556 404
rect 550 399 551 403
rect 555 399 556 403
rect 594 403 595 407
rect 599 403 600 407
rect 594 402 600 403
rect 550 398 556 399
rect 542 394 548 395
rect 534 391 540 392
rect 534 387 535 391
rect 539 387 540 391
rect 542 390 543 394
rect 547 390 548 394
rect 542 389 548 390
rect 534 386 540 387
rect 526 371 532 372
rect 526 367 527 371
rect 531 367 532 371
rect 596 368 598 402
rect 526 366 532 367
rect 594 367 600 368
rect 518 331 524 332
rect 518 327 519 331
rect 523 327 524 331
rect 518 326 524 327
rect 447 322 451 323
rect 447 317 451 318
rect 455 322 459 323
rect 455 317 459 318
rect 487 322 491 323
rect 487 317 491 318
rect 503 322 507 323
rect 503 317 507 318
rect 519 322 523 323
rect 519 317 523 318
rect 456 304 458 317
rect 488 304 490 317
rect 520 304 522 317
rect 528 309 530 366
rect 594 363 595 367
rect 599 363 600 367
rect 594 362 600 363
rect 534 356 540 357
rect 534 352 535 356
rect 539 352 540 356
rect 534 351 540 352
rect 536 323 538 351
rect 566 339 572 340
rect 566 335 567 339
rect 571 335 572 339
rect 566 334 572 335
rect 535 322 539 323
rect 535 317 539 318
rect 551 322 555 323
rect 551 317 555 318
rect 527 308 531 309
rect 552 304 554 317
rect 454 303 460 304
rect 454 299 455 303
rect 459 299 460 303
rect 454 298 460 299
rect 486 303 492 304
rect 486 299 487 303
rect 491 299 492 303
rect 486 298 492 299
rect 518 303 524 304
rect 527 303 531 304
rect 550 303 556 304
rect 518 299 519 303
rect 523 299 524 303
rect 518 298 524 299
rect 550 299 551 303
rect 555 299 556 303
rect 550 298 556 299
rect 568 296 570 334
rect 599 322 603 323
rect 599 317 603 318
rect 600 307 602 317
rect 598 306 604 307
rect 598 302 599 306
rect 603 302 604 306
rect 598 301 604 302
rect 530 295 536 296
rect 530 294 531 295
rect 528 291 531 294
rect 535 291 536 295
rect 528 290 536 291
rect 566 295 572 296
rect 566 291 567 295
rect 571 291 572 295
rect 566 290 572 291
rect 454 286 460 287
rect 454 282 455 286
rect 459 282 460 286
rect 454 281 460 282
rect 486 286 492 287
rect 486 282 487 286
rect 491 282 492 286
rect 486 281 492 282
rect 518 286 524 287
rect 518 282 519 286
rect 523 282 524 286
rect 518 281 524 282
rect 430 279 436 280
rect 430 275 431 279
rect 435 275 436 279
rect 430 274 436 275
rect 456 251 458 281
rect 488 251 490 281
rect 520 251 522 281
rect 375 250 379 251
rect 375 245 379 246
rect 391 250 395 251
rect 391 245 395 246
rect 407 250 411 251
rect 407 245 411 246
rect 423 250 427 251
rect 423 245 427 246
rect 439 250 443 251
rect 439 245 443 246
rect 455 250 459 251
rect 455 245 459 246
rect 471 250 475 251
rect 471 245 475 246
rect 487 250 491 251
rect 487 245 491 246
rect 503 250 507 251
rect 503 245 507 246
rect 519 250 523 251
rect 519 245 523 246
rect 376 215 378 245
rect 408 215 410 245
rect 440 215 442 245
rect 472 215 474 245
rect 504 215 506 245
rect 519 219 525 220
rect 519 215 520 219
rect 524 218 525 219
rect 528 218 530 290
rect 550 286 556 287
rect 550 282 551 286
rect 555 282 556 286
rect 550 281 556 282
rect 552 251 554 281
rect 582 279 588 280
rect 582 275 583 279
rect 587 275 588 279
rect 582 274 588 275
rect 535 250 539 251
rect 535 245 539 246
rect 551 250 555 251
rect 551 245 555 246
rect 567 250 571 251
rect 567 245 571 246
rect 524 216 530 218
rect 524 215 525 216
rect 536 215 538 245
rect 568 215 570 245
rect 584 232 586 274
rect 598 265 604 266
rect 598 261 599 265
rect 603 261 604 265
rect 608 261 610 446
rect 615 442 619 443
rect 615 437 619 438
rect 616 400 618 437
rect 628 404 630 486
rect 642 483 643 487
rect 647 483 648 487
rect 642 482 648 483
rect 644 416 646 482
rect 656 443 658 493
rect 666 487 672 488
rect 666 483 667 487
rect 671 483 672 487
rect 716 484 718 522
rect 746 519 752 520
rect 746 515 747 519
rect 751 515 752 519
rect 746 514 752 515
rect 726 493 732 494
rect 726 489 727 493
rect 731 489 732 493
rect 726 488 732 489
rect 666 482 672 483
rect 714 483 720 484
rect 668 468 670 482
rect 714 479 715 483
rect 719 479 720 483
rect 714 478 720 479
rect 666 467 672 468
rect 666 463 667 467
rect 671 463 672 467
rect 666 462 672 463
rect 686 451 692 452
rect 686 447 687 451
rect 691 447 692 451
rect 686 446 692 447
rect 655 442 659 443
rect 655 437 659 438
rect 671 442 675 443
rect 671 437 675 438
rect 642 415 648 416
rect 642 411 643 415
rect 647 411 648 415
rect 642 410 648 411
rect 626 403 632 404
rect 614 399 620 400
rect 614 395 615 399
rect 619 395 620 399
rect 626 399 627 403
rect 631 399 632 403
rect 626 398 632 399
rect 614 394 620 395
rect 644 372 646 410
rect 672 396 674 437
rect 678 435 684 436
rect 678 431 679 435
rect 683 431 684 435
rect 678 430 684 431
rect 670 395 676 396
rect 670 391 671 395
rect 675 391 676 395
rect 670 390 676 391
rect 642 371 648 372
rect 642 367 643 371
rect 647 367 648 371
rect 642 366 648 367
rect 670 354 676 355
rect 614 352 620 353
rect 614 348 615 352
rect 619 348 620 352
rect 670 350 671 354
rect 675 350 676 354
rect 670 349 676 350
rect 614 347 620 348
rect 616 323 618 347
rect 672 323 674 349
rect 615 322 619 323
rect 615 317 619 318
rect 671 322 675 323
rect 671 317 675 318
rect 622 275 628 276
rect 622 271 623 275
rect 627 271 628 275
rect 622 270 628 271
rect 598 260 604 261
rect 607 260 611 261
rect 600 251 602 260
rect 606 255 612 256
rect 606 251 607 255
rect 611 251 612 255
rect 599 250 603 251
rect 606 250 612 251
rect 624 248 626 270
rect 680 253 682 430
rect 688 404 690 446
rect 728 443 730 488
rect 734 487 740 488
rect 734 483 735 487
rect 739 483 740 487
rect 734 482 740 483
rect 727 442 731 443
rect 727 437 731 438
rect 736 412 738 482
rect 748 476 750 514
rect 766 507 772 508
rect 766 503 767 507
rect 771 503 772 507
rect 766 502 772 503
rect 746 475 752 476
rect 746 471 747 475
rect 751 471 752 475
rect 746 470 752 471
rect 748 416 750 470
rect 755 442 759 443
rect 755 437 759 438
rect 746 415 752 416
rect 734 411 740 412
rect 734 407 735 411
rect 739 407 740 411
rect 746 411 747 415
rect 751 411 752 415
rect 746 410 752 411
rect 734 406 740 407
rect 686 403 692 404
rect 686 399 687 403
rect 691 399 692 403
rect 686 398 692 399
rect 718 403 724 404
rect 718 399 719 403
rect 723 399 724 403
rect 718 398 724 399
rect 710 331 716 332
rect 710 327 711 331
rect 715 327 716 331
rect 710 326 716 327
rect 703 322 707 323
rect 703 317 707 318
rect 704 307 706 317
rect 702 306 708 307
rect 702 302 703 306
rect 707 302 708 306
rect 702 301 708 302
rect 702 265 708 266
rect 702 261 703 265
rect 707 261 708 265
rect 702 260 708 261
rect 672 251 682 253
rect 704 251 706 260
rect 712 256 714 326
rect 710 255 716 256
rect 710 251 711 255
rect 715 251 716 255
rect 639 250 643 251
rect 599 245 603 246
rect 622 247 628 248
rect 582 231 588 232
rect 582 227 583 231
rect 587 227 588 231
rect 582 226 588 227
rect 600 215 602 245
rect 622 243 623 247
rect 627 243 628 247
rect 672 248 674 251
rect 695 250 699 251
rect 639 245 643 246
rect 670 247 676 248
rect 622 242 628 243
rect 374 214 380 215
rect 366 211 372 212
rect 366 207 367 211
rect 371 207 372 211
rect 374 210 375 214
rect 379 210 380 214
rect 374 209 380 210
rect 406 214 412 215
rect 406 210 407 214
rect 411 210 412 214
rect 406 209 412 210
rect 438 214 444 215
rect 438 210 439 214
rect 443 210 444 214
rect 438 209 444 210
rect 470 214 476 215
rect 470 210 471 214
rect 475 210 476 214
rect 470 209 476 210
rect 502 214 508 215
rect 519 214 525 215
rect 534 214 540 215
rect 502 210 503 214
rect 507 210 508 214
rect 502 209 508 210
rect 534 210 535 214
rect 539 210 540 214
rect 534 209 540 210
rect 566 214 572 215
rect 566 210 567 214
rect 571 210 572 214
rect 566 209 572 210
rect 598 214 604 215
rect 598 210 599 214
rect 603 210 604 214
rect 598 209 604 210
rect 366 206 372 207
rect 486 203 492 204
rect 486 199 487 203
rect 491 199 492 203
rect 486 198 492 199
rect 614 203 620 204
rect 614 199 615 203
rect 619 199 620 203
rect 614 198 620 199
rect 374 197 380 198
rect 374 193 375 197
rect 379 193 380 197
rect 374 192 380 193
rect 406 197 412 198
rect 406 193 407 197
rect 411 193 412 197
rect 406 192 412 193
rect 438 197 444 198
rect 438 193 439 197
rect 443 193 444 197
rect 438 192 444 193
rect 470 197 476 198
rect 470 193 471 197
rect 475 193 476 197
rect 470 192 476 193
rect 488 192 490 198
rect 502 197 508 198
rect 502 193 503 197
rect 507 193 508 197
rect 502 192 508 193
rect 534 197 540 198
rect 534 193 535 197
rect 539 193 540 197
rect 534 192 540 193
rect 566 197 572 198
rect 566 193 567 197
rect 571 193 572 197
rect 566 192 572 193
rect 598 197 604 198
rect 598 193 599 197
rect 603 193 604 197
rect 598 192 604 193
rect 184 175 186 192
rect 216 175 218 192
rect 248 175 250 192
rect 280 175 282 192
rect 312 175 314 192
rect 344 175 346 192
rect 358 191 364 192
rect 358 187 359 191
rect 363 187 364 191
rect 358 186 364 187
rect 376 175 378 192
rect 408 175 410 192
rect 440 175 442 192
rect 472 175 474 192
rect 486 191 492 192
rect 486 187 487 191
rect 491 187 492 191
rect 486 186 492 187
rect 504 175 506 192
rect 536 175 538 192
rect 568 175 570 192
rect 600 175 602 192
rect 111 174 115 175
rect 111 169 115 170
rect 135 174 139 175
rect 112 166 114 169
rect 135 168 139 170
rect 167 174 171 175
rect 167 168 171 170
rect 183 174 187 175
rect 183 169 187 170
rect 215 174 219 175
rect 215 168 219 170
rect 247 174 251 175
rect 247 169 251 170
rect 263 174 267 175
rect 263 168 267 170
rect 279 174 283 175
rect 279 169 283 170
rect 311 174 315 175
rect 311 168 315 170
rect 343 174 347 175
rect 343 169 347 170
rect 367 174 371 175
rect 367 168 371 170
rect 375 174 379 175
rect 375 169 379 170
rect 407 174 411 175
rect 407 169 411 170
rect 415 174 419 175
rect 415 168 419 170
rect 439 174 443 175
rect 439 169 443 170
rect 471 174 475 175
rect 471 168 475 170
rect 503 174 507 175
rect 503 169 507 170
rect 535 174 539 175
rect 535 168 539 170
rect 567 174 571 175
rect 567 169 571 170
rect 599 174 603 175
rect 599 169 603 170
rect 607 174 611 175
rect 607 168 611 170
rect 134 167 140 168
rect 110 165 116 166
rect 110 161 111 165
rect 115 161 116 165
rect 134 163 135 167
rect 139 163 140 167
rect 134 162 140 163
rect 166 167 172 168
rect 166 163 167 167
rect 171 163 172 167
rect 166 162 172 163
rect 214 167 220 168
rect 214 163 215 167
rect 219 163 220 167
rect 214 162 220 163
rect 262 167 268 168
rect 262 163 263 167
rect 267 163 268 167
rect 262 162 268 163
rect 310 167 316 168
rect 310 163 311 167
rect 315 163 316 167
rect 310 162 316 163
rect 366 167 372 168
rect 366 163 367 167
rect 371 163 372 167
rect 366 162 372 163
rect 414 167 420 168
rect 414 163 415 167
rect 419 163 420 167
rect 414 162 420 163
rect 470 167 476 168
rect 470 163 471 167
rect 475 163 476 167
rect 470 162 476 163
rect 534 167 540 168
rect 534 163 535 167
rect 539 163 540 167
rect 534 162 540 163
rect 606 167 612 168
rect 606 163 607 167
rect 611 163 612 167
rect 606 162 612 163
rect 110 160 116 161
rect 150 159 156 160
rect 150 155 151 159
rect 155 155 156 159
rect 150 154 156 155
rect 134 150 140 151
rect 110 148 116 149
rect 110 144 111 148
rect 115 144 116 148
rect 134 146 135 150
rect 139 146 140 150
rect 134 145 140 146
rect 110 143 116 144
rect 112 123 114 143
rect 136 123 138 145
rect 111 122 115 123
rect 111 117 115 118
rect 135 122 139 123
rect 135 117 139 118
rect 112 109 114 117
rect 110 108 116 109
rect 110 104 111 108
rect 115 104 116 108
rect 136 107 138 117
rect 152 112 154 154
rect 166 150 172 151
rect 166 146 167 150
rect 171 146 172 150
rect 166 145 172 146
rect 214 150 220 151
rect 214 146 215 150
rect 219 146 220 150
rect 214 145 220 146
rect 262 150 268 151
rect 262 146 263 150
rect 267 146 268 150
rect 262 145 268 146
rect 310 150 316 151
rect 310 146 311 150
rect 315 146 316 150
rect 310 145 316 146
rect 366 150 372 151
rect 366 146 367 150
rect 371 146 372 150
rect 366 145 372 146
rect 414 150 420 151
rect 414 146 415 150
rect 419 146 420 150
rect 414 145 420 146
rect 470 150 476 151
rect 470 146 471 150
rect 475 146 476 150
rect 470 145 476 146
rect 534 150 540 151
rect 534 146 535 150
rect 539 146 540 150
rect 534 145 540 146
rect 606 150 612 151
rect 606 146 607 150
rect 611 146 612 150
rect 606 145 612 146
rect 168 123 170 145
rect 216 123 218 145
rect 264 123 266 145
rect 312 123 314 145
rect 368 123 370 145
rect 416 123 418 145
rect 472 123 474 145
rect 536 123 538 145
rect 608 123 610 145
rect 616 144 618 198
rect 614 143 620 144
rect 614 139 615 143
rect 619 139 620 143
rect 614 138 620 139
rect 167 122 171 123
rect 167 117 171 118
rect 199 122 203 123
rect 199 117 203 118
rect 215 122 219 123
rect 215 117 219 118
rect 231 122 235 123
rect 231 117 235 118
rect 263 122 267 123
rect 263 117 267 118
rect 295 122 299 123
rect 295 117 299 118
rect 311 122 315 123
rect 311 117 315 118
rect 327 122 331 123
rect 327 117 331 118
rect 359 122 363 123
rect 359 117 363 118
rect 367 122 371 123
rect 367 117 371 118
rect 391 122 395 123
rect 391 117 395 118
rect 415 122 419 123
rect 415 117 419 118
rect 423 122 427 123
rect 423 117 427 118
rect 455 122 459 123
rect 455 117 459 118
rect 471 122 475 123
rect 471 117 475 118
rect 487 122 491 123
rect 487 117 491 118
rect 519 122 523 123
rect 519 117 523 118
rect 535 122 539 123
rect 535 117 539 118
rect 551 122 555 123
rect 551 117 555 118
rect 607 122 611 123
rect 607 117 611 118
rect 150 111 156 112
rect 150 107 151 111
rect 155 107 156 111
rect 168 107 170 117
rect 200 107 202 117
rect 232 107 234 117
rect 264 107 266 117
rect 296 107 298 117
rect 328 107 330 117
rect 360 107 362 117
rect 392 107 394 117
rect 424 107 426 117
rect 456 107 458 117
rect 488 107 490 117
rect 520 107 522 117
rect 552 107 554 117
rect 608 107 610 117
rect 110 103 116 104
rect 134 106 140 107
rect 150 106 156 107
rect 166 106 172 107
rect 134 102 135 106
rect 139 102 140 106
rect 134 101 140 102
rect 166 102 167 106
rect 171 102 172 106
rect 166 101 172 102
rect 198 106 204 107
rect 198 102 199 106
rect 203 102 204 106
rect 198 101 204 102
rect 230 106 236 107
rect 230 102 231 106
rect 235 102 236 106
rect 230 101 236 102
rect 262 106 268 107
rect 262 102 263 106
rect 267 102 268 106
rect 262 101 268 102
rect 294 106 300 107
rect 294 102 295 106
rect 299 102 300 106
rect 294 101 300 102
rect 326 106 332 107
rect 326 102 327 106
rect 331 102 332 106
rect 326 101 332 102
rect 358 106 364 107
rect 358 102 359 106
rect 363 102 364 106
rect 358 101 364 102
rect 390 106 396 107
rect 390 102 391 106
rect 395 102 396 106
rect 390 101 396 102
rect 422 106 428 107
rect 422 102 423 106
rect 427 102 428 106
rect 422 101 428 102
rect 454 106 460 107
rect 454 102 455 106
rect 459 102 460 106
rect 454 101 460 102
rect 486 106 492 107
rect 486 102 487 106
rect 491 102 492 106
rect 486 101 492 102
rect 518 106 524 107
rect 518 102 519 106
rect 523 102 524 106
rect 518 101 524 102
rect 550 106 556 107
rect 550 102 551 106
rect 555 102 556 106
rect 550 101 556 102
rect 606 106 612 107
rect 606 102 607 106
rect 611 102 612 106
rect 606 101 612 102
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 110 86 116 87
rect 134 89 140 90
rect 112 83 114 86
rect 134 85 135 89
rect 139 85 140 89
rect 134 84 140 85
rect 166 89 172 90
rect 166 85 167 89
rect 171 85 172 89
rect 166 84 172 85
rect 198 89 204 90
rect 198 85 199 89
rect 203 85 204 89
rect 198 84 204 85
rect 230 89 236 90
rect 230 85 231 89
rect 235 85 236 89
rect 230 84 236 85
rect 262 89 268 90
rect 262 85 263 89
rect 267 85 268 89
rect 262 84 268 85
rect 294 89 300 90
rect 294 85 295 89
rect 299 85 300 89
rect 294 84 300 85
rect 326 89 332 90
rect 326 85 327 89
rect 331 85 332 89
rect 326 84 332 85
rect 358 89 364 90
rect 358 85 359 89
rect 363 85 364 89
rect 358 84 364 85
rect 390 89 396 90
rect 390 85 391 89
rect 395 85 396 89
rect 390 84 396 85
rect 422 89 428 90
rect 422 85 423 89
rect 427 85 428 89
rect 422 84 428 85
rect 454 89 460 90
rect 454 85 455 89
rect 459 85 460 89
rect 454 84 460 85
rect 486 89 492 90
rect 486 85 487 89
rect 491 85 492 89
rect 486 84 492 85
rect 518 89 524 90
rect 518 85 519 89
rect 523 85 524 89
rect 518 84 524 85
rect 550 89 556 90
rect 550 85 551 89
rect 555 85 556 89
rect 550 84 556 85
rect 606 89 612 90
rect 606 85 607 89
rect 611 85 612 89
rect 624 88 626 242
rect 640 215 642 245
rect 670 243 671 247
rect 675 243 676 247
rect 695 245 699 246
rect 703 250 707 251
rect 710 250 716 251
rect 703 245 707 246
rect 670 242 676 243
rect 696 236 698 245
rect 694 235 700 236
rect 654 231 660 232
rect 654 227 655 231
rect 659 227 660 231
rect 694 231 695 235
rect 699 231 700 235
rect 694 230 700 231
rect 654 226 660 227
rect 646 219 652 220
rect 646 215 647 219
rect 651 215 652 219
rect 638 214 644 215
rect 646 214 652 215
rect 638 210 639 214
rect 643 210 644 214
rect 638 209 644 210
rect 638 197 644 198
rect 638 193 639 197
rect 643 193 644 197
rect 638 192 644 193
rect 640 175 642 192
rect 639 174 643 175
rect 639 169 643 170
rect 648 160 650 214
rect 656 204 658 226
rect 720 224 722 398
rect 756 376 758 437
rect 768 408 770 502
rect 782 498 788 499
rect 782 494 783 498
rect 787 494 788 498
rect 782 493 788 494
rect 784 443 786 493
rect 796 488 798 558
rect 832 531 834 618
rect 824 529 834 531
rect 794 487 800 488
rect 794 483 795 487
rect 799 483 800 487
rect 794 482 800 483
rect 806 487 812 488
rect 806 483 807 487
rect 811 483 812 487
rect 806 482 812 483
rect 796 468 798 482
rect 794 467 800 468
rect 794 463 795 467
rect 799 463 800 467
rect 794 462 800 463
rect 783 442 787 443
rect 783 437 787 438
rect 808 428 810 482
rect 806 427 812 428
rect 806 423 807 427
rect 811 423 812 427
rect 806 422 812 423
rect 766 407 772 408
rect 766 403 767 407
rect 771 403 772 407
rect 766 402 772 403
rect 754 375 760 376
rect 754 371 755 375
rect 759 371 760 375
rect 754 370 760 371
rect 782 360 788 361
rect 782 356 783 360
rect 787 356 788 360
rect 782 355 788 356
rect 784 323 786 355
rect 783 322 787 323
rect 783 317 787 318
rect 807 322 811 323
rect 807 317 811 318
rect 808 307 810 317
rect 806 306 812 307
rect 806 302 807 306
rect 811 302 812 306
rect 806 301 812 302
rect 778 295 784 296
rect 778 291 779 295
rect 783 291 784 295
rect 778 290 784 291
rect 780 256 782 290
rect 806 265 812 266
rect 806 261 807 265
rect 811 261 812 265
rect 806 260 812 261
rect 778 255 784 256
rect 778 251 779 255
rect 783 251 784 255
rect 808 251 810 260
rect 824 256 826 529
rect 842 527 848 528
rect 842 523 843 527
rect 847 523 848 527
rect 842 522 848 523
rect 834 519 840 520
rect 834 515 835 519
rect 839 515 840 519
rect 834 514 840 515
rect 836 488 838 514
rect 834 487 840 488
rect 834 483 835 487
rect 839 483 840 487
rect 844 484 846 522
rect 834 482 840 483
rect 842 483 848 484
rect 842 479 843 483
rect 847 479 848 483
rect 842 478 848 479
rect 830 275 836 276
rect 830 271 831 275
rect 835 271 836 275
rect 830 270 836 271
rect 822 255 828 256
rect 822 251 823 255
rect 827 251 828 255
rect 778 250 784 251
rect 791 250 795 251
rect 791 245 795 246
rect 807 250 811 251
rect 822 250 828 251
rect 807 245 811 246
rect 718 223 724 224
rect 718 219 719 223
rect 723 219 724 223
rect 718 218 724 219
rect 792 215 794 245
rect 832 240 834 270
rect 839 250 843 251
rect 839 245 843 246
rect 806 239 812 240
rect 806 235 807 239
rect 811 235 812 239
rect 806 234 812 235
rect 830 239 836 240
rect 830 235 831 239
rect 835 235 836 239
rect 830 234 836 235
rect 790 214 796 215
rect 790 210 791 214
rect 795 210 796 214
rect 790 209 796 210
rect 808 204 810 234
rect 840 230 842 245
rect 852 240 854 658
rect 864 643 866 705
rect 1006 695 1012 696
rect 1006 691 1007 695
rect 1011 691 1012 695
rect 1006 690 1012 691
rect 910 689 916 690
rect 910 685 911 689
rect 915 685 916 689
rect 910 684 916 685
rect 983 684 987 685
rect 912 643 914 684
rect 982 679 988 680
rect 982 675 983 679
rect 987 675 988 679
rect 982 674 988 675
rect 1008 643 1010 690
rect 1036 684 1038 770
rect 1014 683 1020 684
rect 1014 679 1015 683
rect 1019 679 1020 683
rect 1014 678 1020 679
rect 1034 683 1040 684
rect 1034 679 1035 683
rect 1039 679 1040 683
rect 1034 678 1040 679
rect 1016 664 1018 678
rect 1014 663 1020 664
rect 1014 659 1015 663
rect 1019 659 1020 663
rect 1014 658 1020 659
rect 863 642 867 643
rect 863 637 867 638
rect 903 642 907 643
rect 903 637 907 638
rect 911 642 915 643
rect 911 637 915 638
rect 999 642 1003 643
rect 999 637 1003 638
rect 1007 642 1011 643
rect 1007 637 1011 638
rect 904 628 906 637
rect 918 635 924 636
rect 918 631 919 635
rect 923 631 924 635
rect 918 630 924 631
rect 950 631 956 632
rect 902 627 908 628
rect 902 623 903 627
rect 907 623 908 627
rect 902 622 908 623
rect 902 580 908 581
rect 902 576 903 580
rect 907 576 908 580
rect 902 575 908 576
rect 904 563 906 575
rect 871 562 875 563
rect 871 557 875 558
rect 903 562 907 563
rect 903 557 907 558
rect 872 541 874 557
rect 870 540 876 541
rect 870 536 871 540
rect 875 536 876 540
rect 870 535 876 536
rect 920 528 922 630
rect 950 627 951 631
rect 955 627 956 631
rect 950 626 956 627
rect 982 631 988 632
rect 982 627 983 631
rect 987 627 988 631
rect 982 626 988 627
rect 927 562 931 563
rect 927 557 931 558
rect 928 537 930 557
rect 926 536 932 537
rect 926 532 927 536
rect 931 532 932 536
rect 926 531 932 532
rect 918 527 924 528
rect 918 523 919 527
rect 923 523 924 527
rect 918 522 924 523
rect 934 498 940 499
rect 934 494 935 498
rect 939 494 940 498
rect 870 493 876 494
rect 934 493 940 494
rect 870 489 871 493
rect 875 489 876 493
rect 870 488 876 489
rect 872 443 874 488
rect 936 443 938 493
rect 942 487 948 488
rect 942 483 943 487
rect 947 483 948 487
rect 942 482 948 483
rect 944 444 946 482
rect 952 476 954 626
rect 958 599 964 600
rect 958 595 959 599
rect 963 595 964 599
rect 958 594 964 595
rect 960 488 962 594
rect 958 487 964 488
rect 958 483 959 487
rect 963 483 964 487
rect 958 482 964 483
rect 950 475 956 476
rect 950 471 951 475
rect 955 471 956 475
rect 950 470 956 471
rect 942 443 948 444
rect 958 443 964 444
rect 871 442 875 443
rect 871 437 875 438
rect 903 442 907 443
rect 903 437 907 438
rect 935 442 939 443
rect 942 439 943 443
rect 947 439 948 443
rect 942 438 948 439
rect 951 442 955 443
rect 958 439 959 443
rect 963 439 964 443
rect 958 438 964 439
rect 935 437 939 438
rect 951 437 955 438
rect 882 411 888 412
rect 882 407 883 411
rect 887 407 888 411
rect 882 406 888 407
rect 884 384 886 406
rect 882 383 888 384
rect 882 379 883 383
rect 887 379 888 383
rect 882 378 888 379
rect 904 375 906 437
rect 922 435 928 436
rect 922 431 923 435
rect 927 431 928 435
rect 922 430 928 431
rect 924 380 926 430
rect 952 395 954 437
rect 960 404 962 438
rect 958 403 964 404
rect 958 399 959 403
rect 963 399 964 403
rect 958 398 964 399
rect 950 394 956 395
rect 950 390 951 394
rect 955 390 956 394
rect 950 389 956 390
rect 922 379 928 380
rect 922 375 923 379
rect 927 375 928 379
rect 902 374 908 375
rect 922 374 928 375
rect 902 370 903 374
rect 907 370 908 374
rect 902 369 908 370
rect 984 365 986 626
rect 1000 623 1002 637
rect 1006 631 1012 632
rect 1006 627 1007 631
rect 1011 627 1012 631
rect 1006 626 1012 627
rect 998 622 1004 623
rect 998 618 999 622
rect 1003 618 1004 622
rect 998 617 1004 618
rect 990 584 996 585
rect 990 580 991 584
rect 995 580 996 584
rect 990 579 996 580
rect 992 563 994 579
rect 1008 564 1010 626
rect 1006 563 1012 564
rect 991 562 995 563
rect 1006 559 1007 563
rect 1011 559 1012 563
rect 1006 558 1012 559
rect 1031 562 1035 563
rect 991 557 995 558
rect 1031 557 1035 558
rect 1032 541 1034 557
rect 1030 540 1036 541
rect 1030 536 1031 540
rect 1035 536 1036 540
rect 1030 535 1036 536
rect 1030 493 1036 494
rect 1030 489 1031 493
rect 1035 489 1036 493
rect 1030 488 1036 489
rect 1002 483 1008 484
rect 1002 479 1003 483
rect 1007 479 1008 483
rect 1002 478 1008 479
rect 1004 368 1006 478
rect 1032 443 1034 488
rect 1044 460 1046 798
rect 1062 671 1068 672
rect 1062 667 1063 671
rect 1067 667 1068 671
rect 1062 666 1068 667
rect 1050 635 1056 636
rect 1050 631 1051 635
rect 1055 631 1056 635
rect 1050 630 1056 631
rect 1052 596 1054 630
rect 1050 595 1056 596
rect 1050 591 1051 595
rect 1055 591 1056 595
rect 1050 590 1056 591
rect 1054 519 1060 520
rect 1054 515 1055 519
rect 1059 515 1060 519
rect 1054 514 1060 515
rect 1056 480 1058 514
rect 1054 479 1060 480
rect 1054 475 1055 479
rect 1059 475 1060 479
rect 1054 474 1060 475
rect 1042 459 1048 460
rect 1042 455 1043 459
rect 1047 455 1048 459
rect 1042 454 1048 455
rect 1031 442 1035 443
rect 1031 437 1035 438
rect 1032 378 1034 437
rect 1056 404 1058 474
rect 1064 404 1066 666
rect 1080 644 1082 882
rect 1112 839 1114 900
rect 1103 838 1107 839
rect 1103 833 1107 834
rect 1111 838 1115 839
rect 1111 833 1115 834
rect 1104 803 1106 833
rect 1124 808 1126 930
rect 1144 925 1146 949
rect 1194 943 1200 944
rect 1194 939 1195 943
rect 1199 939 1200 943
rect 1194 938 1200 939
rect 1142 924 1148 925
rect 1142 920 1143 924
rect 1147 920 1148 924
rect 1142 919 1148 920
rect 1142 905 1148 906
rect 1142 901 1143 905
rect 1147 901 1148 905
rect 1142 900 1148 901
rect 1144 839 1146 900
rect 1143 838 1147 839
rect 1143 833 1147 834
rect 1167 838 1171 839
rect 1167 833 1171 834
rect 1110 807 1116 808
rect 1110 803 1111 807
rect 1115 803 1116 807
rect 1102 802 1108 803
rect 1110 802 1116 803
rect 1122 807 1128 808
rect 1122 803 1123 807
rect 1127 803 1128 807
rect 1168 806 1170 833
rect 1196 808 1198 938
rect 1240 924 1242 949
rect 1272 925 1274 949
rect 1270 924 1276 925
rect 1238 923 1244 924
rect 1238 919 1239 923
rect 1243 919 1244 923
rect 1270 920 1271 924
rect 1275 920 1276 924
rect 1270 919 1276 920
rect 1238 918 1244 919
rect 1230 915 1236 916
rect 1230 911 1231 915
rect 1235 911 1236 915
rect 1230 910 1236 911
rect 1354 911 1360 912
rect 1206 899 1212 900
rect 1206 895 1207 899
rect 1211 895 1212 899
rect 1206 894 1212 895
rect 1208 884 1210 894
rect 1206 883 1212 884
rect 1206 879 1207 883
rect 1211 879 1212 883
rect 1206 878 1212 879
rect 1232 824 1234 910
rect 1354 907 1355 911
rect 1359 907 1360 911
rect 1354 906 1360 907
rect 1238 905 1244 906
rect 1238 901 1239 905
rect 1243 901 1244 905
rect 1238 900 1244 901
rect 1270 905 1276 906
rect 1270 901 1271 905
rect 1275 901 1276 905
rect 1270 900 1276 901
rect 1240 839 1242 900
rect 1254 839 1260 840
rect 1272 839 1274 900
rect 1356 892 1358 906
rect 1374 903 1380 904
rect 1374 899 1375 903
rect 1379 899 1380 903
rect 1374 898 1380 899
rect 1354 891 1360 892
rect 1354 887 1355 891
rect 1359 887 1360 891
rect 1354 886 1360 887
rect 1239 838 1243 839
rect 1239 833 1243 834
rect 1247 838 1251 839
rect 1254 835 1255 839
rect 1259 835 1260 839
rect 1254 834 1260 835
rect 1271 838 1275 839
rect 1247 833 1251 834
rect 1230 823 1236 824
rect 1230 819 1231 823
rect 1235 819 1236 823
rect 1230 818 1236 819
rect 1194 807 1200 808
rect 1122 802 1128 803
rect 1166 805 1172 806
rect 1102 798 1103 802
rect 1107 798 1108 802
rect 1102 797 1108 798
rect 1102 785 1108 786
rect 1102 781 1103 785
rect 1107 781 1108 785
rect 1102 780 1108 781
rect 1104 755 1106 780
rect 1087 754 1091 755
rect 1087 749 1091 750
rect 1103 754 1107 755
rect 1103 749 1107 750
rect 1088 729 1090 749
rect 1086 728 1092 729
rect 1086 724 1087 728
rect 1091 724 1092 728
rect 1086 723 1092 724
rect 1094 690 1100 691
rect 1094 686 1095 690
rect 1099 686 1100 690
rect 1094 685 1100 686
rect 1086 679 1092 680
rect 1086 675 1087 679
rect 1091 675 1092 679
rect 1086 674 1092 675
rect 1078 643 1084 644
rect 1078 639 1079 643
rect 1083 639 1084 643
rect 1078 638 1084 639
rect 1088 452 1090 674
rect 1096 643 1098 685
rect 1102 679 1108 680
rect 1102 675 1103 679
rect 1107 675 1108 679
rect 1102 674 1108 675
rect 1104 656 1106 674
rect 1112 664 1114 802
rect 1166 801 1167 805
rect 1171 801 1172 805
rect 1194 803 1195 807
rect 1199 803 1200 807
rect 1248 806 1250 833
rect 1256 820 1258 834
rect 1271 833 1275 834
rect 1295 838 1299 839
rect 1295 833 1299 834
rect 1327 838 1331 839
rect 1327 833 1331 834
rect 1278 831 1284 832
rect 1278 827 1279 831
rect 1283 827 1284 831
rect 1278 826 1284 827
rect 1254 819 1260 820
rect 1254 815 1255 819
rect 1259 815 1260 819
rect 1254 814 1260 815
rect 1194 802 1200 803
rect 1246 805 1252 806
rect 1166 800 1172 801
rect 1246 801 1247 805
rect 1251 801 1252 805
rect 1246 800 1252 801
rect 1158 791 1164 792
rect 1158 787 1159 791
rect 1163 787 1164 791
rect 1158 786 1164 787
rect 1160 772 1162 786
rect 1230 784 1236 785
rect 1230 780 1231 784
rect 1235 780 1236 784
rect 1230 779 1236 780
rect 1182 778 1188 779
rect 1182 774 1183 778
rect 1187 774 1188 778
rect 1182 773 1188 774
rect 1158 771 1164 772
rect 1158 767 1159 771
rect 1163 767 1164 771
rect 1158 766 1164 767
rect 1184 755 1186 773
rect 1222 759 1228 760
rect 1222 755 1223 759
rect 1227 755 1228 759
rect 1232 755 1234 779
rect 1167 754 1171 755
rect 1167 749 1171 750
rect 1183 754 1187 755
rect 1183 749 1187 750
rect 1207 754 1211 755
rect 1222 754 1228 755
rect 1231 754 1235 755
rect 1207 749 1211 750
rect 1168 733 1170 749
rect 1166 732 1172 733
rect 1166 728 1167 732
rect 1171 728 1172 732
rect 1208 729 1210 749
rect 1166 727 1172 728
rect 1206 728 1212 729
rect 1206 724 1207 728
rect 1211 724 1212 728
rect 1206 723 1212 724
rect 1154 719 1160 720
rect 1154 715 1155 719
rect 1159 715 1160 719
rect 1154 714 1160 715
rect 1146 711 1152 712
rect 1146 707 1147 711
rect 1151 707 1152 711
rect 1146 706 1152 707
rect 1148 680 1150 706
rect 1146 679 1152 680
rect 1146 675 1147 679
rect 1151 675 1152 679
rect 1156 676 1158 714
rect 1224 712 1226 754
rect 1231 749 1235 750
rect 1247 754 1251 755
rect 1247 749 1251 750
rect 1248 728 1250 749
rect 1246 727 1252 728
rect 1246 723 1247 727
rect 1251 723 1252 727
rect 1246 722 1252 723
rect 1234 719 1240 720
rect 1234 715 1235 719
rect 1239 715 1240 719
rect 1234 714 1240 715
rect 1222 711 1228 712
rect 1222 707 1223 711
rect 1227 707 1228 711
rect 1222 706 1228 707
rect 1226 703 1232 704
rect 1206 700 1212 701
rect 1206 696 1207 700
rect 1211 696 1212 700
rect 1226 699 1227 703
rect 1231 699 1232 703
rect 1226 698 1232 699
rect 1206 695 1212 696
rect 1166 685 1172 686
rect 1166 681 1167 685
rect 1171 681 1172 685
rect 1166 680 1172 681
rect 1146 674 1152 675
rect 1154 675 1160 676
rect 1154 671 1155 675
rect 1159 671 1160 675
rect 1154 670 1160 671
rect 1110 663 1116 664
rect 1110 659 1111 663
rect 1115 659 1116 663
rect 1110 658 1116 659
rect 1102 655 1108 656
rect 1102 651 1103 655
rect 1107 651 1108 655
rect 1102 650 1108 651
rect 1095 642 1099 643
rect 1095 637 1099 638
rect 1104 568 1106 650
rect 1168 643 1170 680
rect 1182 679 1188 680
rect 1182 675 1183 679
rect 1187 675 1188 679
rect 1182 674 1188 675
rect 1174 659 1180 660
rect 1174 655 1175 659
rect 1179 655 1180 659
rect 1174 654 1180 655
rect 1119 642 1123 643
rect 1119 637 1123 638
rect 1167 642 1171 643
rect 1167 637 1171 638
rect 1120 628 1122 637
rect 1142 631 1148 632
rect 1110 627 1116 628
rect 1110 623 1111 627
rect 1115 623 1116 627
rect 1110 622 1116 623
rect 1118 627 1124 628
rect 1118 623 1119 627
rect 1123 623 1124 627
rect 1142 627 1143 631
rect 1147 627 1148 631
rect 1142 626 1148 627
rect 1118 622 1124 623
rect 1112 600 1114 622
rect 1110 599 1116 600
rect 1110 595 1111 599
rect 1115 595 1116 599
rect 1110 594 1116 595
rect 1118 580 1124 581
rect 1118 576 1119 580
rect 1123 576 1124 580
rect 1118 575 1124 576
rect 1102 567 1108 568
rect 1102 563 1103 567
rect 1107 563 1108 567
rect 1120 563 1122 575
rect 1095 562 1099 563
rect 1102 562 1108 563
rect 1119 562 1123 563
rect 1095 557 1099 558
rect 1096 537 1098 557
rect 1094 536 1100 537
rect 1094 532 1095 536
rect 1099 532 1100 536
rect 1094 531 1100 532
rect 1104 506 1106 562
rect 1119 557 1123 558
rect 1104 504 1114 506
rect 1144 504 1146 626
rect 1154 519 1160 520
rect 1154 515 1155 519
rect 1159 515 1160 519
rect 1154 514 1160 515
rect 1102 498 1108 499
rect 1102 494 1103 498
rect 1107 494 1108 498
rect 1102 493 1108 494
rect 1086 451 1092 452
rect 1086 447 1087 451
rect 1091 447 1092 451
rect 1086 446 1092 447
rect 1104 443 1106 493
rect 1112 488 1114 504
rect 1142 503 1148 504
rect 1142 499 1143 503
rect 1147 499 1148 503
rect 1142 498 1148 499
rect 1156 488 1158 514
rect 1110 487 1116 488
rect 1110 483 1111 487
rect 1115 483 1116 487
rect 1110 482 1116 483
rect 1154 487 1160 488
rect 1154 483 1155 487
rect 1159 483 1160 487
rect 1154 482 1160 483
rect 1156 475 1158 482
rect 1156 473 1170 475
rect 1075 442 1079 443
rect 1075 437 1079 438
rect 1103 442 1107 443
rect 1103 437 1107 438
rect 1054 403 1060 404
rect 1054 399 1055 403
rect 1059 399 1060 403
rect 1054 398 1060 399
rect 1062 403 1068 404
rect 1062 399 1063 403
rect 1067 399 1068 403
rect 1062 398 1068 399
rect 1064 380 1066 398
rect 1062 379 1068 380
rect 1030 377 1036 378
rect 1030 373 1031 377
rect 1035 373 1036 377
rect 1062 375 1063 379
rect 1067 375 1068 379
rect 1076 376 1078 437
rect 1168 416 1170 473
rect 1176 416 1178 654
rect 1184 640 1186 674
rect 1208 643 1210 695
rect 1228 683 1230 698
rect 1236 692 1238 714
rect 1246 710 1252 711
rect 1246 706 1247 710
rect 1251 706 1252 710
rect 1246 705 1252 706
rect 1234 691 1240 692
rect 1234 687 1235 691
rect 1239 687 1240 691
rect 1234 686 1240 687
rect 1228 681 1234 683
rect 1207 642 1211 643
rect 1182 639 1188 640
rect 1182 635 1183 639
rect 1187 635 1188 639
rect 1207 637 1211 638
rect 1215 642 1219 643
rect 1215 637 1219 638
rect 1182 634 1188 635
rect 1216 623 1218 637
rect 1222 631 1228 632
rect 1222 627 1223 631
rect 1227 627 1228 631
rect 1222 626 1228 627
rect 1214 622 1220 623
rect 1214 618 1215 622
rect 1219 618 1220 622
rect 1214 617 1220 618
rect 1206 584 1212 585
rect 1206 580 1207 584
rect 1211 580 1212 584
rect 1206 579 1212 580
rect 1208 563 1210 579
rect 1224 568 1226 626
rect 1222 567 1228 568
rect 1222 563 1223 567
rect 1227 563 1228 567
rect 1199 562 1203 563
rect 1199 557 1203 558
rect 1207 562 1211 563
rect 1222 562 1228 563
rect 1207 557 1211 558
rect 1200 541 1202 557
rect 1198 540 1204 541
rect 1198 536 1199 540
rect 1203 536 1204 540
rect 1198 535 1204 536
rect 1190 527 1196 528
rect 1190 523 1191 527
rect 1195 523 1196 527
rect 1190 522 1196 523
rect 1192 484 1194 522
rect 1222 507 1228 508
rect 1222 503 1223 507
rect 1227 503 1228 507
rect 1222 502 1228 503
rect 1198 493 1204 494
rect 1198 489 1199 493
rect 1203 489 1204 493
rect 1198 488 1204 489
rect 1224 488 1226 502
rect 1190 483 1196 484
rect 1190 479 1191 483
rect 1195 479 1196 483
rect 1190 478 1196 479
rect 1200 443 1202 488
rect 1222 487 1228 488
rect 1222 483 1223 487
rect 1227 483 1228 487
rect 1222 482 1228 483
rect 1214 479 1220 480
rect 1214 475 1215 479
rect 1219 475 1220 479
rect 1214 474 1220 475
rect 1199 442 1203 443
rect 1199 437 1203 438
rect 1190 423 1196 424
rect 1190 419 1191 423
rect 1195 419 1196 423
rect 1190 418 1196 419
rect 1162 415 1170 416
rect 1162 411 1163 415
rect 1167 411 1170 415
rect 1162 410 1170 411
rect 1174 415 1180 416
rect 1174 411 1175 415
rect 1179 411 1180 415
rect 1174 410 1180 411
rect 1164 409 1170 410
rect 1126 399 1132 400
rect 1126 395 1127 399
rect 1131 395 1132 399
rect 1126 394 1132 395
rect 1062 374 1068 375
rect 1074 375 1080 376
rect 1030 372 1036 373
rect 1074 371 1075 375
rect 1079 371 1080 375
rect 1074 370 1080 371
rect 1002 367 1008 368
rect 983 364 987 365
rect 918 363 924 364
rect 878 359 884 360
rect 878 355 879 359
rect 883 355 884 359
rect 918 359 919 363
rect 923 359 924 363
rect 1002 363 1003 367
rect 1007 363 1008 367
rect 1002 362 1008 363
rect 983 359 987 360
rect 1102 360 1108 361
rect 918 358 924 359
rect 878 354 884 355
rect 902 357 908 358
rect 880 256 882 354
rect 902 353 903 357
rect 907 353 908 357
rect 902 352 908 353
rect 904 323 906 352
rect 903 322 907 323
rect 903 317 907 318
rect 911 322 915 323
rect 911 317 915 318
rect 912 307 914 317
rect 910 306 916 307
rect 910 302 911 306
rect 915 302 916 306
rect 910 301 916 302
rect 920 296 922 358
rect 942 356 948 357
rect 942 352 943 356
rect 947 352 948 356
rect 1102 356 1103 360
rect 1107 356 1108 360
rect 1102 355 1108 356
rect 942 351 948 352
rect 944 323 946 351
rect 1046 350 1052 351
rect 1046 346 1047 350
rect 1051 346 1052 350
rect 1046 345 1052 346
rect 1038 343 1044 344
rect 1038 339 1039 343
rect 1043 339 1044 343
rect 1038 338 1044 339
rect 982 323 988 324
rect 943 322 947 323
rect 982 319 983 323
rect 987 319 988 323
rect 982 318 988 319
rect 999 322 1003 323
rect 943 317 947 318
rect 918 295 924 296
rect 918 291 919 295
rect 923 291 924 295
rect 918 290 924 291
rect 984 276 986 318
rect 999 317 1003 318
rect 1031 322 1035 323
rect 1031 317 1035 318
rect 1000 304 1002 317
rect 1032 304 1034 317
rect 1040 307 1042 338
rect 1048 323 1050 345
rect 1104 323 1106 355
rect 1047 322 1051 323
rect 1047 317 1051 318
rect 1063 322 1067 323
rect 1063 317 1067 318
rect 1103 322 1107 323
rect 1103 317 1107 318
rect 1111 322 1115 323
rect 1111 317 1115 318
rect 1040 305 1046 307
rect 998 303 1004 304
rect 998 299 999 303
rect 1003 299 1004 303
rect 998 298 1004 299
rect 1030 303 1036 304
rect 1030 299 1031 303
rect 1035 299 1036 303
rect 1030 298 1036 299
rect 1044 296 1046 305
rect 1064 304 1066 317
rect 1112 307 1114 317
rect 1110 306 1116 307
rect 1062 303 1068 304
rect 1062 299 1063 303
rect 1067 299 1068 303
rect 1110 302 1111 306
rect 1115 302 1116 306
rect 1110 301 1116 302
rect 1062 298 1068 299
rect 1042 295 1048 296
rect 1042 291 1043 295
rect 1047 291 1048 295
rect 1042 290 1048 291
rect 998 286 1004 287
rect 998 282 999 286
rect 1003 282 1004 286
rect 998 281 1004 282
rect 1030 286 1036 287
rect 1030 282 1031 286
rect 1035 282 1036 286
rect 1030 281 1036 282
rect 1062 286 1068 287
rect 1062 282 1063 286
rect 1067 282 1068 286
rect 1062 281 1068 282
rect 982 275 988 276
rect 982 271 983 275
rect 987 271 988 275
rect 982 270 988 271
rect 910 265 916 266
rect 910 261 911 265
rect 915 261 916 265
rect 910 260 916 261
rect 927 260 931 261
rect 878 255 884 256
rect 878 251 879 255
rect 883 251 884 255
rect 912 251 914 260
rect 926 255 932 256
rect 926 251 927 255
rect 931 251 932 255
rect 982 255 988 256
rect 982 251 983 255
rect 987 251 988 255
rect 1000 251 1002 281
rect 1006 275 1012 276
rect 1006 271 1007 275
rect 1011 271 1012 275
rect 1006 270 1012 271
rect 1008 252 1010 270
rect 1006 251 1012 252
rect 1032 251 1034 281
rect 1064 251 1066 281
rect 1082 271 1088 272
rect 1082 267 1083 271
rect 1087 267 1088 271
rect 1082 266 1088 267
rect 878 250 884 251
rect 911 250 915 251
rect 911 245 915 246
rect 919 250 923 251
rect 926 250 932 251
rect 967 250 971 251
rect 982 250 988 251
rect 999 250 1003 251
rect 919 245 923 246
rect 967 245 971 246
rect 850 239 856 240
rect 850 235 851 239
rect 855 235 856 239
rect 850 234 856 235
rect 838 229 844 230
rect 838 225 839 229
rect 843 225 844 229
rect 838 224 844 225
rect 920 220 922 245
rect 934 239 940 240
rect 934 235 935 239
rect 939 235 940 239
rect 968 236 970 245
rect 934 234 940 235
rect 966 235 972 236
rect 918 219 924 220
rect 918 215 919 219
rect 923 215 924 219
rect 918 214 924 215
rect 654 203 660 204
rect 654 199 655 203
rect 659 199 660 203
rect 654 198 660 199
rect 806 203 812 204
rect 806 199 807 203
rect 811 199 812 203
rect 936 200 938 234
rect 966 231 967 235
rect 971 231 972 235
rect 966 230 972 231
rect 984 224 986 250
rect 1006 247 1007 251
rect 1011 247 1012 251
rect 1006 246 1012 247
rect 1031 250 1035 251
rect 999 245 1003 246
rect 1031 245 1035 246
rect 1063 250 1067 251
rect 1063 245 1067 246
rect 982 223 988 224
rect 982 219 983 223
rect 987 219 988 223
rect 982 218 988 219
rect 1064 215 1066 245
rect 1074 219 1080 220
rect 1074 215 1075 219
rect 1079 215 1080 219
rect 1062 214 1068 215
rect 1074 214 1080 215
rect 1062 210 1063 214
rect 1067 210 1068 214
rect 1062 209 1068 210
rect 806 198 812 199
rect 934 199 940 200
rect 790 197 796 198
rect 694 194 700 195
rect 694 190 695 194
rect 699 190 700 194
rect 790 193 791 197
rect 795 193 796 197
rect 790 192 796 193
rect 918 196 924 197
rect 918 192 919 196
rect 923 192 924 196
rect 934 195 935 199
rect 939 195 940 199
rect 1062 197 1068 198
rect 934 194 940 195
rect 966 194 972 195
rect 694 189 700 190
rect 696 175 698 189
rect 792 175 794 192
rect 918 191 924 192
rect 830 189 836 190
rect 830 185 831 189
rect 835 185 836 189
rect 830 184 836 185
rect 832 175 834 184
rect 920 175 922 191
rect 966 190 967 194
rect 971 190 972 194
rect 1062 193 1063 197
rect 1067 193 1068 197
rect 1062 192 1068 193
rect 966 189 972 190
rect 968 175 970 189
rect 1064 175 1066 192
rect 687 174 691 175
rect 687 168 691 170
rect 695 174 699 175
rect 695 169 699 170
rect 775 174 779 175
rect 775 168 779 170
rect 791 174 795 175
rect 791 169 795 170
rect 831 174 835 175
rect 831 169 835 170
rect 863 174 867 175
rect 863 168 867 170
rect 919 174 923 175
rect 919 169 923 170
rect 959 174 963 175
rect 959 168 963 170
rect 967 174 971 175
rect 967 169 971 170
rect 1055 174 1059 175
rect 1055 168 1059 170
rect 1063 174 1067 175
rect 1063 169 1067 170
rect 686 167 692 168
rect 686 163 687 167
rect 691 163 692 167
rect 686 162 692 163
rect 774 167 780 168
rect 774 163 775 167
rect 779 163 780 167
rect 774 162 780 163
rect 862 167 868 168
rect 862 163 863 167
rect 867 163 868 167
rect 862 162 868 163
rect 958 167 964 168
rect 958 163 959 167
rect 963 163 964 167
rect 958 162 964 163
rect 1054 167 1060 168
rect 1054 163 1055 167
rect 1059 163 1060 167
rect 1054 162 1060 163
rect 1076 160 1078 214
rect 1084 204 1086 266
rect 1110 265 1116 266
rect 1110 261 1111 265
rect 1115 261 1116 265
rect 1110 260 1116 261
rect 1112 251 1114 260
rect 1128 256 1130 394
rect 1176 320 1178 410
rect 1192 388 1194 418
rect 1216 388 1218 474
rect 1232 468 1234 681
rect 1248 643 1250 705
rect 1256 680 1258 814
rect 1280 804 1282 826
rect 1296 804 1298 833
rect 1328 804 1330 833
rect 1356 816 1358 886
rect 1376 839 1378 898
rect 1384 884 1386 986
rect 1426 983 1432 984
rect 1426 979 1427 983
rect 1431 982 1432 983
rect 1431 979 1434 982
rect 1426 978 1434 979
rect 1406 977 1412 978
rect 1406 973 1407 977
rect 1411 973 1412 977
rect 1406 972 1412 973
rect 1408 955 1410 972
rect 1391 954 1395 955
rect 1391 949 1395 950
rect 1407 954 1411 955
rect 1407 949 1411 950
rect 1423 954 1427 955
rect 1423 949 1427 950
rect 1392 931 1394 949
rect 1398 947 1404 948
rect 1398 943 1399 947
rect 1403 943 1404 947
rect 1398 942 1404 943
rect 1390 930 1396 931
rect 1390 926 1391 930
rect 1395 926 1396 930
rect 1390 925 1396 926
rect 1400 900 1402 942
rect 1424 924 1426 949
rect 1422 923 1428 924
rect 1422 919 1423 923
rect 1427 919 1428 923
rect 1422 918 1428 919
rect 1422 906 1428 907
rect 1422 902 1423 906
rect 1427 902 1428 906
rect 1422 901 1428 902
rect 1398 899 1404 900
rect 1398 895 1399 899
rect 1403 895 1404 899
rect 1398 894 1404 895
rect 1414 891 1420 892
rect 1414 887 1415 891
rect 1419 887 1420 891
rect 1414 886 1420 887
rect 1382 883 1388 884
rect 1382 879 1383 883
rect 1387 879 1388 883
rect 1382 878 1388 879
rect 1375 838 1379 839
rect 1375 833 1379 834
rect 1416 824 1418 886
rect 1424 839 1426 901
rect 1432 900 1434 978
rect 1438 977 1444 978
rect 1438 973 1439 977
rect 1443 973 1444 977
rect 1438 972 1444 973
rect 1440 955 1442 972
rect 1439 954 1443 955
rect 1439 949 1443 950
rect 1430 899 1436 900
rect 1430 895 1431 899
rect 1435 895 1436 899
rect 1430 894 1436 895
rect 1423 838 1427 839
rect 1423 833 1427 834
rect 1414 823 1420 824
rect 1414 819 1415 823
rect 1419 819 1420 823
rect 1414 818 1420 819
rect 1354 815 1360 816
rect 1354 811 1355 815
rect 1359 811 1360 815
rect 1424 813 1426 833
rect 1354 810 1360 811
rect 1422 812 1428 813
rect 1422 808 1423 812
rect 1427 808 1428 812
rect 1422 807 1428 808
rect 1278 803 1284 804
rect 1278 799 1279 803
rect 1283 799 1284 803
rect 1278 798 1284 799
rect 1294 803 1300 804
rect 1294 799 1295 803
rect 1299 799 1300 803
rect 1294 798 1300 799
rect 1326 803 1332 804
rect 1326 799 1327 803
rect 1331 799 1332 803
rect 1326 798 1332 799
rect 1271 796 1275 797
rect 1270 791 1271 796
rect 1275 791 1276 796
rect 1270 790 1276 791
rect 1254 679 1260 680
rect 1254 675 1255 679
rect 1259 675 1260 679
rect 1254 674 1260 675
rect 1272 643 1274 790
rect 1294 785 1300 786
rect 1294 781 1295 785
rect 1299 781 1300 785
rect 1294 780 1300 781
rect 1326 784 1332 785
rect 1326 780 1327 784
rect 1331 780 1332 784
rect 1296 755 1298 780
rect 1326 779 1332 780
rect 1422 784 1428 785
rect 1422 780 1423 784
rect 1427 780 1428 784
rect 1422 779 1428 780
rect 1328 755 1330 779
rect 1424 755 1426 779
rect 1279 754 1283 755
rect 1279 749 1283 750
rect 1295 754 1299 755
rect 1295 749 1299 750
rect 1311 754 1315 755
rect 1311 749 1315 750
rect 1327 754 1331 755
rect 1327 749 1331 750
rect 1343 754 1347 755
rect 1343 749 1347 750
rect 1375 754 1379 755
rect 1375 749 1379 750
rect 1407 754 1411 755
rect 1407 749 1411 750
rect 1423 754 1427 755
rect 1423 749 1427 750
rect 1439 754 1443 755
rect 1439 749 1443 750
rect 1280 728 1282 749
rect 1312 728 1314 749
rect 1344 728 1346 749
rect 1376 728 1378 749
rect 1408 728 1410 749
rect 1440 728 1442 749
rect 1278 727 1284 728
rect 1278 723 1279 727
rect 1283 723 1284 727
rect 1278 722 1284 723
rect 1310 727 1316 728
rect 1310 723 1311 727
rect 1315 723 1316 727
rect 1310 722 1316 723
rect 1342 727 1348 728
rect 1342 723 1343 727
rect 1347 723 1348 727
rect 1342 722 1348 723
rect 1374 727 1380 728
rect 1374 723 1375 727
rect 1379 723 1380 727
rect 1374 722 1380 723
rect 1406 727 1412 728
rect 1406 723 1407 727
rect 1411 723 1412 727
rect 1406 722 1412 723
rect 1438 727 1444 728
rect 1438 723 1439 727
rect 1443 723 1444 727
rect 1438 722 1444 723
rect 1448 715 1450 1070
rect 1456 1035 1458 1101
rect 1455 1034 1459 1035
rect 1455 1029 1459 1030
rect 1454 1011 1460 1012
rect 1454 1007 1455 1011
rect 1459 1007 1460 1011
rect 1454 1006 1460 1007
rect 1456 984 1458 1006
rect 1472 1000 1474 1110
rect 1486 1106 1492 1107
rect 1486 1102 1487 1106
rect 1491 1102 1492 1106
rect 1486 1101 1492 1102
rect 1518 1106 1524 1107
rect 1518 1102 1519 1106
rect 1523 1102 1524 1106
rect 1518 1101 1524 1102
rect 1488 1035 1490 1101
rect 1520 1035 1522 1101
rect 1479 1034 1483 1035
rect 1479 1029 1483 1030
rect 1487 1034 1491 1035
rect 1487 1029 1491 1030
rect 1519 1034 1523 1035
rect 1519 1029 1523 1030
rect 1470 999 1476 1000
rect 1470 995 1471 999
rect 1475 995 1476 999
rect 1480 995 1482 1029
rect 1520 995 1522 1029
rect 1536 1000 1538 1110
rect 1558 1106 1564 1107
rect 1558 1102 1559 1106
rect 1563 1102 1564 1106
rect 1558 1101 1564 1102
rect 1560 1035 1562 1101
rect 1576 1100 1578 1178
rect 1590 1177 1596 1178
rect 1590 1173 1591 1177
rect 1595 1173 1596 1177
rect 1590 1172 1596 1173
rect 1592 1151 1594 1172
rect 1591 1150 1595 1151
rect 1591 1145 1595 1146
rect 1592 1124 1594 1145
rect 1590 1123 1596 1124
rect 1590 1119 1591 1123
rect 1595 1119 1596 1123
rect 1590 1118 1596 1119
rect 1612 1108 1614 1178
rect 1622 1177 1628 1178
rect 1622 1173 1623 1177
rect 1627 1173 1628 1177
rect 1622 1172 1628 1173
rect 1654 1177 1660 1178
rect 1654 1173 1655 1177
rect 1659 1173 1660 1177
rect 1694 1175 1695 1179
rect 1699 1175 1700 1179
rect 1694 1174 1700 1175
rect 1654 1172 1660 1173
rect 1624 1151 1626 1172
rect 1656 1151 1658 1172
rect 1696 1151 1698 1174
rect 1623 1150 1627 1151
rect 1623 1145 1627 1146
rect 1655 1150 1659 1151
rect 1655 1145 1659 1146
rect 1695 1150 1699 1151
rect 1695 1145 1699 1146
rect 1624 1124 1626 1145
rect 1656 1124 1658 1145
rect 1622 1123 1628 1124
rect 1622 1119 1623 1123
rect 1627 1119 1628 1123
rect 1622 1118 1628 1119
rect 1654 1123 1660 1124
rect 1654 1119 1655 1123
rect 1659 1119 1660 1123
rect 1696 1122 1698 1145
rect 1654 1118 1660 1119
rect 1694 1121 1700 1122
rect 1694 1117 1695 1121
rect 1699 1117 1700 1121
rect 1694 1116 1700 1117
rect 1670 1115 1676 1116
rect 1670 1111 1671 1115
rect 1675 1111 1676 1115
rect 1670 1110 1676 1111
rect 1610 1107 1616 1108
rect 1590 1106 1596 1107
rect 1590 1102 1591 1106
rect 1595 1102 1596 1106
rect 1610 1103 1611 1107
rect 1615 1103 1616 1107
rect 1610 1102 1616 1103
rect 1622 1106 1628 1107
rect 1622 1102 1623 1106
rect 1627 1102 1628 1106
rect 1590 1101 1596 1102
rect 1622 1101 1628 1102
rect 1654 1106 1660 1107
rect 1654 1102 1655 1106
rect 1659 1102 1660 1106
rect 1654 1101 1660 1102
rect 1574 1099 1580 1100
rect 1574 1095 1575 1099
rect 1579 1095 1580 1099
rect 1574 1094 1580 1095
rect 1592 1035 1594 1101
rect 1624 1035 1626 1101
rect 1656 1035 1658 1101
rect 1672 1092 1674 1110
rect 1694 1104 1700 1105
rect 1694 1100 1695 1104
rect 1699 1100 1700 1104
rect 1694 1099 1700 1100
rect 1670 1091 1676 1092
rect 1670 1087 1671 1091
rect 1675 1087 1676 1091
rect 1670 1086 1676 1087
rect 1696 1035 1698 1099
rect 1559 1034 1563 1035
rect 1559 1029 1563 1030
rect 1591 1034 1595 1035
rect 1591 1029 1595 1030
rect 1623 1034 1627 1035
rect 1623 1029 1627 1030
rect 1655 1034 1659 1035
rect 1655 1029 1659 1030
rect 1695 1034 1699 1035
rect 1695 1029 1699 1030
rect 1534 999 1540 1000
rect 1534 995 1535 999
rect 1539 995 1540 999
rect 1560 995 1562 1029
rect 1592 995 1594 1029
rect 1624 995 1626 1029
rect 1656 995 1658 1029
rect 1696 997 1698 1029
rect 1694 996 1700 997
rect 1470 994 1476 995
rect 1478 994 1484 995
rect 1478 990 1479 994
rect 1483 990 1484 994
rect 1478 989 1484 990
rect 1518 994 1524 995
rect 1534 994 1540 995
rect 1558 994 1564 995
rect 1518 990 1519 994
rect 1523 990 1524 994
rect 1518 989 1524 990
rect 1558 990 1559 994
rect 1563 990 1564 994
rect 1558 989 1564 990
rect 1590 994 1596 995
rect 1590 990 1591 994
rect 1595 990 1596 994
rect 1590 989 1596 990
rect 1622 994 1628 995
rect 1622 990 1623 994
rect 1627 990 1628 994
rect 1622 989 1628 990
rect 1654 994 1660 995
rect 1654 990 1655 994
rect 1659 990 1660 994
rect 1694 992 1695 996
rect 1699 992 1700 996
rect 1694 991 1700 992
rect 1654 989 1660 990
rect 1454 983 1460 984
rect 1454 979 1455 983
rect 1459 979 1460 983
rect 1454 978 1460 979
rect 1494 983 1500 984
rect 1494 979 1495 983
rect 1499 979 1500 983
rect 1494 978 1500 979
rect 1694 979 1700 980
rect 1478 977 1484 978
rect 1478 973 1479 977
rect 1483 973 1484 977
rect 1478 972 1484 973
rect 1480 955 1482 972
rect 1455 954 1459 955
rect 1455 949 1459 950
rect 1479 954 1483 955
rect 1479 949 1483 950
rect 1456 925 1458 949
rect 1454 924 1460 925
rect 1454 920 1455 924
rect 1459 920 1460 924
rect 1454 919 1460 920
rect 1470 903 1476 904
rect 1470 899 1471 903
rect 1475 899 1476 903
rect 1470 898 1476 899
rect 1472 839 1474 898
rect 1478 887 1484 888
rect 1478 883 1479 887
rect 1483 883 1484 887
rect 1478 882 1484 883
rect 1480 840 1482 882
rect 1478 839 1484 840
rect 1471 838 1475 839
rect 1478 835 1479 839
rect 1483 835 1484 839
rect 1478 834 1484 835
rect 1471 833 1475 834
rect 1472 813 1474 833
rect 1480 824 1482 834
rect 1478 823 1484 824
rect 1478 819 1479 823
rect 1483 819 1484 823
rect 1496 820 1498 978
rect 1518 977 1524 978
rect 1518 973 1519 977
rect 1523 973 1524 977
rect 1518 972 1524 973
rect 1558 977 1564 978
rect 1558 973 1559 977
rect 1563 973 1564 977
rect 1558 972 1564 973
rect 1590 977 1596 978
rect 1590 973 1591 977
rect 1595 973 1596 977
rect 1590 972 1596 973
rect 1622 977 1628 978
rect 1622 973 1623 977
rect 1627 973 1628 977
rect 1622 972 1628 973
rect 1654 977 1660 978
rect 1654 973 1655 977
rect 1659 973 1660 977
rect 1694 975 1695 979
rect 1699 975 1700 979
rect 1694 974 1700 975
rect 1654 972 1660 973
rect 1520 955 1522 972
rect 1538 971 1544 972
rect 1538 967 1539 971
rect 1543 967 1544 971
rect 1538 966 1544 967
rect 1519 954 1523 955
rect 1519 949 1523 950
rect 1520 924 1522 949
rect 1518 923 1524 924
rect 1518 919 1519 923
rect 1523 919 1524 923
rect 1518 918 1524 919
rect 1518 906 1524 907
rect 1518 902 1519 906
rect 1523 902 1524 906
rect 1518 901 1524 902
rect 1520 839 1522 901
rect 1540 900 1542 966
rect 1560 955 1562 972
rect 1592 955 1594 972
rect 1624 955 1626 972
rect 1656 955 1658 972
rect 1696 955 1698 974
rect 1559 954 1563 955
rect 1559 949 1563 950
rect 1591 954 1595 955
rect 1591 949 1595 950
rect 1623 954 1627 955
rect 1623 949 1627 950
rect 1655 954 1659 955
rect 1655 949 1659 950
rect 1695 954 1699 955
rect 1695 949 1699 950
rect 1560 924 1562 949
rect 1592 924 1594 949
rect 1624 924 1626 949
rect 1656 924 1658 949
rect 1558 923 1564 924
rect 1558 919 1559 923
rect 1563 919 1564 923
rect 1558 918 1564 919
rect 1590 923 1596 924
rect 1590 919 1591 923
rect 1595 919 1596 923
rect 1590 918 1596 919
rect 1622 923 1628 924
rect 1622 919 1623 923
rect 1627 919 1628 923
rect 1622 918 1628 919
rect 1654 923 1660 924
rect 1654 919 1655 923
rect 1659 919 1660 923
rect 1696 922 1698 949
rect 1654 918 1660 919
rect 1694 921 1700 922
rect 1694 917 1695 921
rect 1699 917 1700 921
rect 1694 916 1700 917
rect 1670 915 1676 916
rect 1670 911 1671 915
rect 1675 911 1676 915
rect 1670 910 1676 911
rect 1558 906 1564 907
rect 1558 902 1559 906
rect 1563 902 1564 906
rect 1558 901 1564 902
rect 1590 906 1596 907
rect 1590 902 1591 906
rect 1595 902 1596 906
rect 1590 901 1596 902
rect 1622 906 1628 907
rect 1622 902 1623 906
rect 1627 902 1628 906
rect 1622 901 1628 902
rect 1654 906 1660 907
rect 1654 902 1655 906
rect 1659 902 1660 906
rect 1654 901 1660 902
rect 1538 899 1544 900
rect 1538 895 1539 899
rect 1543 895 1544 899
rect 1538 894 1544 895
rect 1560 839 1562 901
rect 1592 839 1594 901
rect 1624 839 1626 901
rect 1656 839 1658 901
rect 1663 884 1667 885
rect 1662 879 1663 884
rect 1667 879 1668 884
rect 1662 878 1668 879
rect 1519 838 1523 839
rect 1519 833 1523 834
rect 1559 838 1563 839
rect 1559 833 1563 834
rect 1591 838 1595 839
rect 1591 833 1595 834
rect 1623 838 1627 839
rect 1623 833 1627 834
rect 1655 838 1659 839
rect 1655 833 1659 834
rect 1478 818 1484 819
rect 1494 819 1500 820
rect 1494 815 1495 819
rect 1499 815 1500 819
rect 1494 814 1500 815
rect 1470 812 1476 813
rect 1470 808 1471 812
rect 1475 808 1476 812
rect 1470 807 1476 808
rect 1520 803 1522 833
rect 1560 803 1562 833
rect 1592 803 1594 833
rect 1624 803 1626 833
rect 1656 803 1658 833
rect 1672 808 1674 910
rect 1694 904 1700 905
rect 1694 900 1695 904
rect 1699 900 1700 904
rect 1694 899 1700 900
rect 1696 839 1698 899
rect 1695 838 1699 839
rect 1695 833 1699 834
rect 1670 807 1676 808
rect 1670 803 1671 807
rect 1675 803 1676 807
rect 1696 805 1698 833
rect 1518 802 1524 803
rect 1518 798 1519 802
rect 1523 798 1524 802
rect 1518 797 1524 798
rect 1558 802 1564 803
rect 1558 798 1559 802
rect 1563 798 1564 802
rect 1558 797 1564 798
rect 1590 802 1596 803
rect 1590 798 1591 802
rect 1595 798 1596 802
rect 1590 797 1596 798
rect 1622 802 1628 803
rect 1622 798 1623 802
rect 1627 798 1628 802
rect 1622 797 1628 798
rect 1654 802 1660 803
rect 1670 802 1676 803
rect 1694 804 1700 805
rect 1654 798 1655 802
rect 1659 798 1660 802
rect 1694 800 1695 804
rect 1699 800 1700 804
rect 1694 799 1700 800
rect 1654 797 1660 798
rect 1694 787 1700 788
rect 1518 785 1524 786
rect 1470 784 1476 785
rect 1470 780 1471 784
rect 1475 780 1476 784
rect 1518 781 1519 785
rect 1523 781 1524 785
rect 1518 780 1524 781
rect 1558 785 1564 786
rect 1558 781 1559 785
rect 1563 781 1564 785
rect 1558 780 1564 781
rect 1590 785 1596 786
rect 1590 781 1591 785
rect 1595 781 1596 785
rect 1590 780 1596 781
rect 1622 785 1628 786
rect 1622 781 1623 785
rect 1627 781 1628 785
rect 1622 780 1628 781
rect 1654 785 1660 786
rect 1654 781 1655 785
rect 1659 781 1660 785
rect 1694 783 1695 787
rect 1699 783 1700 787
rect 1694 782 1700 783
rect 1654 780 1660 781
rect 1470 779 1476 780
rect 1498 779 1504 780
rect 1472 755 1474 779
rect 1498 775 1499 779
rect 1503 775 1504 779
rect 1498 774 1504 775
rect 1471 754 1475 755
rect 1471 749 1475 750
rect 1479 754 1483 755
rect 1479 749 1483 750
rect 1480 728 1482 749
rect 1478 727 1484 728
rect 1478 723 1479 727
rect 1483 723 1484 727
rect 1478 722 1484 723
rect 1448 713 1458 715
rect 1278 710 1284 711
rect 1278 706 1279 710
rect 1283 706 1284 710
rect 1278 705 1284 706
rect 1310 710 1316 711
rect 1310 706 1311 710
rect 1315 706 1316 710
rect 1310 705 1316 706
rect 1342 710 1348 711
rect 1342 706 1343 710
rect 1347 706 1348 710
rect 1342 705 1348 706
rect 1374 710 1380 711
rect 1374 706 1375 710
rect 1379 706 1380 710
rect 1374 705 1380 706
rect 1406 710 1412 711
rect 1406 706 1407 710
rect 1411 706 1412 710
rect 1406 705 1412 706
rect 1438 710 1444 711
rect 1438 706 1439 710
rect 1443 706 1444 710
rect 1438 705 1444 706
rect 1280 643 1282 705
rect 1312 643 1314 705
rect 1344 643 1346 705
rect 1358 679 1364 680
rect 1358 675 1359 679
rect 1363 675 1364 679
rect 1358 674 1364 675
rect 1247 642 1251 643
rect 1247 637 1251 638
rect 1260 641 1274 643
rect 1279 642 1283 643
rect 1260 523 1262 641
rect 1279 637 1283 638
rect 1311 642 1315 643
rect 1311 637 1315 638
rect 1335 642 1339 643
rect 1335 637 1339 638
rect 1343 642 1347 643
rect 1343 637 1347 638
rect 1266 635 1272 636
rect 1266 631 1267 635
rect 1271 631 1272 635
rect 1266 630 1272 631
rect 1268 596 1270 630
rect 1336 628 1338 637
rect 1360 632 1362 674
rect 1376 643 1378 705
rect 1408 643 1410 705
rect 1440 643 1442 705
rect 1446 703 1452 704
rect 1446 699 1447 703
rect 1451 699 1452 703
rect 1446 698 1452 699
rect 1375 642 1379 643
rect 1375 637 1379 638
rect 1407 642 1411 643
rect 1407 637 1411 638
rect 1415 642 1419 643
rect 1415 637 1419 638
rect 1439 642 1443 643
rect 1439 637 1443 638
rect 1358 631 1364 632
rect 1334 627 1340 628
rect 1334 623 1335 627
rect 1339 623 1340 627
rect 1358 627 1359 631
rect 1363 627 1364 631
rect 1358 626 1364 627
rect 1334 622 1340 623
rect 1346 619 1352 620
rect 1346 615 1347 619
rect 1351 615 1352 619
rect 1346 614 1352 615
rect 1348 600 1350 614
rect 1416 603 1418 637
rect 1434 607 1440 608
rect 1434 603 1435 607
rect 1439 603 1440 607
rect 1414 602 1420 603
rect 1434 602 1440 603
rect 1346 599 1352 600
rect 1266 595 1272 596
rect 1266 591 1267 595
rect 1271 591 1272 595
rect 1346 595 1347 599
rect 1351 595 1352 599
rect 1414 598 1415 602
rect 1419 598 1420 602
rect 1414 597 1420 598
rect 1346 594 1352 595
rect 1266 590 1272 591
rect 1334 580 1340 581
rect 1334 576 1335 580
rect 1339 576 1340 580
rect 1334 575 1340 576
rect 1336 563 1338 575
rect 1287 562 1291 563
rect 1287 557 1291 558
rect 1335 562 1339 563
rect 1335 557 1339 558
rect 1288 533 1290 557
rect 1286 532 1292 533
rect 1286 528 1287 532
rect 1291 528 1292 532
rect 1286 527 1292 528
rect 1260 521 1270 523
rect 1258 517 1264 518
rect 1258 513 1259 517
rect 1263 513 1264 517
rect 1258 512 1264 513
rect 1230 467 1236 468
rect 1230 463 1231 467
rect 1235 463 1236 467
rect 1230 462 1236 463
rect 1260 443 1262 512
rect 1231 442 1235 443
rect 1231 437 1235 438
rect 1259 442 1263 443
rect 1259 437 1263 438
rect 1232 396 1234 437
rect 1268 424 1270 521
rect 1348 476 1350 594
rect 1414 585 1420 586
rect 1414 581 1415 585
rect 1419 581 1420 585
rect 1414 580 1420 581
rect 1416 563 1418 580
rect 1415 562 1419 563
rect 1415 557 1419 558
rect 1423 562 1427 563
rect 1423 557 1427 558
rect 1424 536 1426 557
rect 1422 535 1428 536
rect 1378 531 1384 532
rect 1378 527 1379 531
rect 1383 527 1384 531
rect 1422 531 1423 535
rect 1427 531 1428 535
rect 1422 530 1428 531
rect 1436 528 1438 602
rect 1448 592 1450 698
rect 1456 692 1458 713
rect 1478 710 1484 711
rect 1478 706 1479 710
rect 1483 706 1484 710
rect 1478 705 1484 706
rect 1454 691 1460 692
rect 1454 687 1455 691
rect 1459 687 1460 691
rect 1454 686 1460 687
rect 1480 643 1482 705
rect 1500 704 1502 774
rect 1520 755 1522 780
rect 1560 755 1562 780
rect 1592 755 1594 780
rect 1624 755 1626 780
rect 1656 755 1658 780
rect 1696 755 1698 782
rect 1519 754 1523 755
rect 1519 749 1523 750
rect 1559 754 1563 755
rect 1559 749 1563 750
rect 1591 754 1595 755
rect 1591 749 1595 750
rect 1623 754 1627 755
rect 1623 749 1627 750
rect 1655 754 1659 755
rect 1655 749 1659 750
rect 1695 754 1699 755
rect 1695 749 1699 750
rect 1520 728 1522 749
rect 1560 728 1562 749
rect 1592 728 1594 749
rect 1624 728 1626 749
rect 1656 728 1658 749
rect 1518 727 1524 728
rect 1518 723 1519 727
rect 1523 723 1524 727
rect 1518 722 1524 723
rect 1558 727 1564 728
rect 1558 723 1559 727
rect 1563 723 1564 727
rect 1558 722 1564 723
rect 1590 727 1596 728
rect 1590 723 1591 727
rect 1595 723 1596 727
rect 1590 722 1596 723
rect 1622 727 1628 728
rect 1622 723 1623 727
rect 1627 723 1628 727
rect 1622 722 1628 723
rect 1654 727 1660 728
rect 1654 723 1655 727
rect 1659 723 1660 727
rect 1696 726 1698 749
rect 1654 722 1660 723
rect 1694 725 1700 726
rect 1694 721 1695 725
rect 1699 721 1700 725
rect 1694 720 1700 721
rect 1670 719 1676 720
rect 1670 715 1671 719
rect 1675 715 1676 719
rect 1670 714 1676 715
rect 1518 710 1524 711
rect 1518 706 1519 710
rect 1523 706 1524 710
rect 1518 705 1524 706
rect 1558 710 1564 711
rect 1558 706 1559 710
rect 1563 706 1564 710
rect 1558 705 1564 706
rect 1590 710 1596 711
rect 1590 706 1591 710
rect 1595 706 1596 710
rect 1590 705 1596 706
rect 1622 710 1628 711
rect 1622 706 1623 710
rect 1627 706 1628 710
rect 1622 705 1628 706
rect 1654 710 1660 711
rect 1654 706 1655 710
rect 1659 706 1660 710
rect 1654 705 1660 706
rect 1498 703 1504 704
rect 1498 699 1499 703
rect 1503 699 1504 703
rect 1498 698 1504 699
rect 1520 643 1522 705
rect 1560 643 1562 705
rect 1592 643 1594 705
rect 1624 643 1626 705
rect 1656 643 1658 705
rect 1479 642 1483 643
rect 1479 637 1483 638
rect 1519 642 1523 643
rect 1519 637 1523 638
rect 1543 642 1547 643
rect 1543 637 1547 638
rect 1559 642 1563 643
rect 1559 637 1563 638
rect 1591 642 1595 643
rect 1591 637 1595 638
rect 1607 642 1611 643
rect 1607 637 1611 638
rect 1623 642 1627 643
rect 1623 637 1627 638
rect 1655 642 1659 643
rect 1655 637 1659 638
rect 1480 603 1482 637
rect 1544 603 1546 637
rect 1608 603 1610 637
rect 1656 603 1658 637
rect 1672 620 1674 714
rect 1694 708 1700 709
rect 1694 704 1695 708
rect 1699 704 1700 708
rect 1694 703 1700 704
rect 1696 643 1698 703
rect 1695 642 1699 643
rect 1695 637 1699 638
rect 1670 619 1676 620
rect 1670 615 1671 619
rect 1675 615 1676 619
rect 1670 614 1676 615
rect 1696 605 1698 637
rect 1694 604 1700 605
rect 1478 602 1484 603
rect 1478 598 1479 602
rect 1483 598 1484 602
rect 1478 597 1484 598
rect 1542 602 1548 603
rect 1542 598 1543 602
rect 1547 598 1548 602
rect 1542 597 1548 598
rect 1606 602 1612 603
rect 1606 598 1607 602
rect 1611 598 1612 602
rect 1606 597 1612 598
rect 1654 602 1660 603
rect 1654 598 1655 602
rect 1659 598 1660 602
rect 1694 600 1695 604
rect 1699 600 1700 604
rect 1694 599 1700 600
rect 1654 597 1660 598
rect 1446 591 1452 592
rect 1446 587 1447 591
rect 1451 587 1452 591
rect 1446 586 1452 587
rect 1670 591 1676 592
rect 1670 587 1671 591
rect 1675 587 1676 591
rect 1670 586 1676 587
rect 1694 587 1700 588
rect 1478 585 1484 586
rect 1478 581 1479 585
rect 1483 581 1484 585
rect 1478 580 1484 581
rect 1542 585 1548 586
rect 1542 581 1543 585
rect 1547 581 1548 585
rect 1542 580 1548 581
rect 1606 585 1612 586
rect 1606 581 1607 585
rect 1611 581 1612 585
rect 1606 580 1612 581
rect 1654 585 1660 586
rect 1654 581 1655 585
rect 1659 581 1660 585
rect 1654 580 1660 581
rect 1480 563 1482 580
rect 1544 563 1546 580
rect 1608 563 1610 580
rect 1656 563 1658 580
rect 1479 562 1483 563
rect 1479 557 1483 558
rect 1527 562 1531 563
rect 1527 557 1531 558
rect 1543 562 1547 563
rect 1543 557 1547 558
rect 1575 562 1579 563
rect 1575 557 1579 558
rect 1607 562 1611 563
rect 1607 557 1611 558
rect 1623 562 1627 563
rect 1623 557 1627 558
rect 1655 562 1659 563
rect 1655 557 1659 558
rect 1480 536 1482 557
rect 1528 536 1530 557
rect 1576 536 1578 557
rect 1624 536 1626 557
rect 1656 536 1658 557
rect 1478 535 1484 536
rect 1478 531 1479 535
rect 1483 531 1484 535
rect 1478 530 1484 531
rect 1526 535 1532 536
rect 1526 531 1527 535
rect 1531 531 1532 535
rect 1526 530 1532 531
rect 1574 535 1580 536
rect 1574 531 1575 535
rect 1579 531 1580 535
rect 1574 530 1580 531
rect 1622 535 1628 536
rect 1622 531 1623 535
rect 1627 531 1628 535
rect 1622 530 1628 531
rect 1654 535 1660 536
rect 1654 531 1655 535
rect 1659 531 1660 535
rect 1654 530 1660 531
rect 1378 526 1384 527
rect 1434 527 1440 528
rect 1346 475 1352 476
rect 1346 471 1347 475
rect 1351 471 1352 475
rect 1346 470 1352 471
rect 1319 442 1323 443
rect 1319 437 1323 438
rect 1359 442 1363 443
rect 1359 437 1363 438
rect 1266 423 1272 424
rect 1266 419 1267 423
rect 1271 419 1272 423
rect 1266 418 1272 419
rect 1230 395 1236 396
rect 1230 391 1231 395
rect 1235 391 1236 395
rect 1230 390 1236 391
rect 1190 387 1196 388
rect 1190 383 1191 387
rect 1195 383 1196 387
rect 1190 382 1196 383
rect 1214 387 1220 388
rect 1214 383 1215 387
rect 1219 383 1220 387
rect 1214 382 1220 383
rect 1320 375 1322 437
rect 1330 435 1336 436
rect 1330 431 1331 435
rect 1335 431 1336 435
rect 1330 430 1336 431
rect 1318 374 1324 375
rect 1318 370 1319 374
rect 1323 370 1324 374
rect 1332 372 1334 430
rect 1338 423 1344 424
rect 1338 419 1339 423
rect 1343 419 1344 423
rect 1338 418 1344 419
rect 1340 380 1342 418
rect 1360 390 1362 437
rect 1366 415 1372 416
rect 1366 411 1367 415
rect 1371 411 1372 415
rect 1366 410 1372 411
rect 1368 400 1370 410
rect 1380 408 1382 526
rect 1434 523 1435 527
rect 1439 523 1440 527
rect 1434 522 1440 523
rect 1606 527 1612 528
rect 1606 523 1607 527
rect 1611 523 1612 527
rect 1606 522 1612 523
rect 1422 518 1428 519
rect 1422 514 1423 518
rect 1427 514 1428 518
rect 1422 513 1428 514
rect 1478 518 1484 519
rect 1478 514 1479 518
rect 1483 514 1484 518
rect 1478 513 1484 514
rect 1526 518 1532 519
rect 1526 514 1527 518
rect 1531 514 1532 518
rect 1526 513 1532 514
rect 1574 518 1580 519
rect 1574 514 1575 518
rect 1579 514 1580 518
rect 1574 513 1580 514
rect 1424 443 1426 513
rect 1480 443 1482 513
rect 1528 443 1530 513
rect 1576 443 1578 513
rect 1582 511 1588 512
rect 1582 507 1583 511
rect 1587 507 1588 511
rect 1582 506 1588 507
rect 1423 442 1427 443
rect 1423 437 1427 438
rect 1439 442 1443 443
rect 1439 437 1443 438
rect 1479 442 1483 443
rect 1479 437 1483 438
rect 1519 442 1523 443
rect 1519 437 1523 438
rect 1527 442 1531 443
rect 1527 437 1531 438
rect 1559 442 1563 443
rect 1559 437 1563 438
rect 1575 442 1579 443
rect 1575 437 1579 438
rect 1378 407 1384 408
rect 1378 403 1379 407
rect 1383 403 1384 407
rect 1378 402 1384 403
rect 1366 399 1372 400
rect 1366 395 1367 399
rect 1371 395 1372 399
rect 1366 394 1372 395
rect 1358 389 1364 390
rect 1358 385 1359 389
rect 1363 385 1364 389
rect 1358 384 1364 385
rect 1440 380 1442 437
rect 1454 399 1460 400
rect 1454 395 1455 399
rect 1459 395 1460 399
rect 1454 394 1460 395
rect 1338 379 1344 380
rect 1338 375 1339 379
rect 1343 375 1344 379
rect 1338 374 1344 375
rect 1438 379 1444 380
rect 1438 375 1439 379
rect 1443 375 1444 379
rect 1438 374 1444 375
rect 1318 369 1324 370
rect 1330 371 1336 372
rect 1330 367 1331 371
rect 1335 367 1336 371
rect 1330 366 1336 367
rect 1334 363 1340 364
rect 1194 359 1200 360
rect 1194 355 1195 359
rect 1199 355 1200 359
rect 1334 359 1335 363
rect 1339 359 1340 363
rect 1456 360 1458 394
rect 1480 375 1482 437
rect 1494 379 1500 380
rect 1494 375 1495 379
rect 1499 375 1500 379
rect 1520 375 1522 437
rect 1560 375 1562 437
rect 1478 374 1484 375
rect 1494 374 1500 375
rect 1518 374 1524 375
rect 1478 370 1479 374
rect 1483 370 1484 374
rect 1478 369 1484 370
rect 1334 358 1340 359
rect 1454 359 1460 360
rect 1318 357 1324 358
rect 1194 354 1200 355
rect 1230 354 1236 355
rect 1196 331 1198 354
rect 1230 350 1231 354
rect 1235 350 1236 354
rect 1318 353 1319 357
rect 1323 353 1324 357
rect 1318 352 1324 353
rect 1230 349 1236 350
rect 1184 329 1198 331
rect 1174 319 1180 320
rect 1174 315 1175 319
rect 1179 315 1180 319
rect 1174 314 1180 315
rect 1184 260 1186 329
rect 1232 323 1234 349
rect 1320 323 1322 352
rect 1199 322 1203 323
rect 1231 322 1235 323
rect 1199 317 1203 318
rect 1214 319 1220 320
rect 1200 312 1202 317
rect 1214 315 1215 319
rect 1219 315 1220 319
rect 1231 317 1235 318
rect 1287 322 1291 323
rect 1287 317 1291 318
rect 1319 322 1323 323
rect 1319 317 1323 318
rect 1214 314 1220 315
rect 1198 311 1204 312
rect 1198 307 1199 311
rect 1203 307 1204 311
rect 1198 306 1204 307
rect 1206 271 1212 272
rect 1206 267 1207 271
rect 1211 267 1212 271
rect 1206 266 1212 267
rect 1182 259 1188 260
rect 1126 255 1132 256
rect 1118 251 1124 252
rect 1103 250 1107 251
rect 1103 245 1107 246
rect 1111 250 1115 251
rect 1118 247 1119 251
rect 1123 247 1124 251
rect 1126 251 1127 255
rect 1131 251 1132 255
rect 1182 255 1183 259
rect 1187 255 1188 259
rect 1182 254 1188 255
rect 1208 251 1210 266
rect 1216 260 1218 314
rect 1288 305 1290 317
rect 1286 304 1292 305
rect 1320 304 1322 317
rect 1286 300 1287 304
rect 1291 300 1292 304
rect 1318 303 1324 304
rect 1286 299 1292 300
rect 1298 299 1304 300
rect 1298 295 1299 299
rect 1303 295 1304 299
rect 1318 299 1319 303
rect 1323 299 1324 303
rect 1318 298 1324 299
rect 1298 294 1304 295
rect 1286 281 1292 282
rect 1286 277 1287 281
rect 1291 277 1292 281
rect 1286 276 1292 277
rect 1214 259 1220 260
rect 1214 255 1215 259
rect 1219 255 1220 259
rect 1214 254 1220 255
rect 1288 251 1290 276
rect 1300 260 1302 294
rect 1318 286 1324 287
rect 1318 282 1319 286
rect 1323 282 1324 286
rect 1318 281 1324 282
rect 1298 259 1304 260
rect 1298 255 1299 259
rect 1303 255 1304 259
rect 1298 254 1304 255
rect 1320 251 1322 281
rect 1336 280 1338 358
rect 1438 356 1444 357
rect 1438 352 1439 356
rect 1443 352 1444 356
rect 1454 355 1455 359
rect 1459 355 1460 359
rect 1454 354 1460 355
rect 1478 357 1484 358
rect 1478 353 1479 357
rect 1483 353 1484 357
rect 1478 352 1484 353
rect 1438 351 1444 352
rect 1350 349 1356 350
rect 1350 345 1351 349
rect 1355 345 1356 349
rect 1350 344 1356 345
rect 1352 323 1354 344
rect 1440 323 1442 351
rect 1480 323 1482 352
rect 1351 322 1355 323
rect 1351 317 1355 318
rect 1383 322 1387 323
rect 1383 317 1387 318
rect 1415 322 1419 323
rect 1415 317 1419 318
rect 1439 322 1443 323
rect 1439 317 1443 318
rect 1447 322 1451 323
rect 1447 317 1451 318
rect 1479 322 1483 323
rect 1479 317 1483 318
rect 1352 304 1354 317
rect 1384 304 1386 317
rect 1416 304 1418 317
rect 1448 304 1450 317
rect 1480 304 1482 317
rect 1496 312 1498 374
rect 1518 370 1519 374
rect 1523 370 1524 374
rect 1518 369 1524 370
rect 1558 374 1564 375
rect 1558 370 1559 374
rect 1563 370 1564 374
rect 1558 369 1564 370
rect 1575 363 1581 364
rect 1575 359 1576 363
rect 1580 362 1581 363
rect 1584 362 1586 506
rect 1591 442 1595 443
rect 1591 437 1595 438
rect 1592 375 1594 437
rect 1608 380 1610 522
rect 1622 518 1628 519
rect 1622 514 1623 518
rect 1627 514 1628 518
rect 1622 513 1628 514
rect 1654 518 1660 519
rect 1654 514 1655 518
rect 1659 514 1660 518
rect 1654 513 1660 514
rect 1624 443 1626 513
rect 1656 443 1658 513
rect 1672 512 1674 586
rect 1694 583 1695 587
rect 1699 583 1700 587
rect 1694 582 1700 583
rect 1696 563 1698 582
rect 1695 562 1699 563
rect 1695 557 1699 558
rect 1696 534 1698 557
rect 1694 533 1700 534
rect 1694 529 1695 533
rect 1699 529 1700 533
rect 1694 528 1700 529
rect 1694 516 1700 517
rect 1694 512 1695 516
rect 1699 512 1700 516
rect 1670 511 1676 512
rect 1694 511 1700 512
rect 1670 507 1671 511
rect 1675 507 1676 511
rect 1670 506 1676 507
rect 1696 443 1698 511
rect 1623 442 1627 443
rect 1623 437 1627 438
rect 1655 442 1659 443
rect 1655 437 1659 438
rect 1695 442 1699 443
rect 1695 437 1699 438
rect 1606 379 1612 380
rect 1606 375 1607 379
rect 1611 375 1612 379
rect 1624 375 1626 437
rect 1656 375 1658 437
rect 1696 377 1698 437
rect 1694 376 1700 377
rect 1590 374 1596 375
rect 1606 374 1612 375
rect 1622 374 1628 375
rect 1590 370 1591 374
rect 1595 370 1596 374
rect 1590 369 1596 370
rect 1622 370 1623 374
rect 1627 370 1628 374
rect 1622 369 1628 370
rect 1654 374 1660 375
rect 1654 370 1655 374
rect 1659 370 1660 374
rect 1694 372 1695 376
rect 1699 372 1700 376
rect 1694 371 1700 372
rect 1654 369 1660 370
rect 1580 360 1586 362
rect 1723 364 1727 365
rect 1580 359 1581 360
rect 1575 358 1581 359
rect 1694 359 1700 360
rect 1723 359 1727 360
rect 1518 357 1524 358
rect 1518 353 1519 357
rect 1523 353 1524 357
rect 1518 352 1524 353
rect 1558 357 1564 358
rect 1558 353 1559 357
rect 1563 353 1564 357
rect 1558 352 1564 353
rect 1590 357 1596 358
rect 1590 353 1591 357
rect 1595 353 1596 357
rect 1590 352 1596 353
rect 1622 357 1628 358
rect 1622 353 1623 357
rect 1627 353 1628 357
rect 1622 352 1628 353
rect 1654 357 1660 358
rect 1654 353 1655 357
rect 1659 353 1660 357
rect 1694 355 1695 359
rect 1699 355 1700 359
rect 1694 354 1700 355
rect 1654 352 1660 353
rect 1520 323 1522 352
rect 1560 323 1562 352
rect 1592 323 1594 352
rect 1624 323 1626 352
rect 1642 351 1648 352
rect 1642 347 1643 351
rect 1647 347 1648 351
rect 1642 346 1648 347
rect 1519 322 1523 323
rect 1519 317 1523 318
rect 1559 322 1563 323
rect 1559 317 1563 318
rect 1591 322 1595 323
rect 1591 317 1595 318
rect 1623 322 1627 323
rect 1623 317 1627 318
rect 1494 311 1500 312
rect 1494 307 1495 311
rect 1499 307 1500 311
rect 1494 306 1500 307
rect 1520 304 1522 317
rect 1560 304 1562 317
rect 1592 304 1594 317
rect 1624 304 1626 317
rect 1350 303 1356 304
rect 1350 299 1351 303
rect 1355 299 1356 303
rect 1350 298 1356 299
rect 1382 303 1388 304
rect 1382 299 1383 303
rect 1387 299 1388 303
rect 1382 298 1388 299
rect 1414 303 1420 304
rect 1414 299 1415 303
rect 1419 299 1420 303
rect 1414 298 1420 299
rect 1446 303 1452 304
rect 1446 299 1447 303
rect 1451 299 1452 303
rect 1446 298 1452 299
rect 1478 303 1484 304
rect 1478 299 1479 303
rect 1483 299 1484 303
rect 1478 298 1484 299
rect 1518 303 1524 304
rect 1518 299 1519 303
rect 1523 299 1524 303
rect 1518 298 1524 299
rect 1558 303 1564 304
rect 1558 299 1559 303
rect 1563 299 1564 303
rect 1558 298 1564 299
rect 1590 303 1596 304
rect 1590 299 1591 303
rect 1595 299 1596 303
rect 1590 298 1596 299
rect 1622 303 1628 304
rect 1622 299 1623 303
rect 1627 299 1628 303
rect 1622 298 1628 299
rect 1530 295 1536 296
rect 1530 291 1531 295
rect 1535 291 1536 295
rect 1530 290 1536 291
rect 1350 286 1356 287
rect 1350 282 1351 286
rect 1355 282 1356 286
rect 1350 281 1356 282
rect 1382 286 1388 287
rect 1382 282 1383 286
rect 1387 282 1388 286
rect 1382 281 1388 282
rect 1414 286 1420 287
rect 1414 282 1415 286
rect 1419 282 1420 286
rect 1414 281 1420 282
rect 1446 286 1452 287
rect 1446 282 1447 286
rect 1451 282 1452 286
rect 1446 281 1452 282
rect 1478 286 1484 287
rect 1478 282 1479 286
rect 1483 282 1484 286
rect 1478 281 1484 282
rect 1518 286 1524 287
rect 1518 282 1519 286
rect 1523 282 1524 286
rect 1518 281 1524 282
rect 1334 279 1340 280
rect 1334 275 1335 279
rect 1339 275 1340 279
rect 1334 274 1340 275
rect 1352 251 1354 281
rect 1384 251 1386 281
rect 1416 251 1418 281
rect 1448 251 1450 281
rect 1480 251 1482 281
rect 1520 251 1522 281
rect 1126 250 1132 251
rect 1143 250 1147 251
rect 1118 246 1124 247
rect 1111 245 1115 246
rect 1104 215 1106 245
rect 1102 214 1108 215
rect 1102 210 1103 214
rect 1107 210 1108 214
rect 1102 209 1108 210
rect 1082 203 1088 204
rect 1082 199 1083 203
rect 1087 199 1088 203
rect 1082 198 1088 199
rect 1102 197 1108 198
rect 1102 193 1103 197
rect 1107 193 1108 197
rect 1102 192 1108 193
rect 1120 192 1122 246
rect 1143 245 1147 246
rect 1183 250 1187 251
rect 1183 245 1187 246
rect 1207 250 1211 251
rect 1207 245 1211 246
rect 1223 250 1227 251
rect 1223 245 1227 246
rect 1263 250 1267 251
rect 1263 245 1267 246
rect 1287 250 1291 251
rect 1287 245 1291 246
rect 1303 250 1307 251
rect 1303 245 1307 246
rect 1319 250 1323 251
rect 1319 245 1323 246
rect 1343 250 1347 251
rect 1343 245 1347 246
rect 1351 250 1355 251
rect 1351 245 1355 246
rect 1375 250 1379 251
rect 1375 245 1379 246
rect 1383 250 1387 251
rect 1383 245 1387 246
rect 1407 250 1411 251
rect 1407 245 1411 246
rect 1415 250 1419 251
rect 1415 245 1419 246
rect 1439 250 1443 251
rect 1439 245 1443 246
rect 1447 250 1451 251
rect 1447 245 1451 246
rect 1479 250 1483 251
rect 1479 245 1483 246
rect 1519 250 1523 251
rect 1519 245 1523 246
rect 1144 215 1146 245
rect 1184 215 1186 245
rect 1198 231 1204 232
rect 1198 227 1199 231
rect 1203 227 1204 231
rect 1198 226 1204 227
rect 1142 214 1148 215
rect 1142 210 1143 214
rect 1147 210 1148 214
rect 1142 209 1148 210
rect 1182 214 1188 215
rect 1182 210 1183 214
rect 1187 210 1188 214
rect 1182 209 1188 210
rect 1200 204 1202 226
rect 1224 215 1226 245
rect 1264 215 1266 245
rect 1304 215 1306 245
rect 1310 223 1316 224
rect 1310 219 1311 223
rect 1315 219 1316 223
rect 1310 218 1316 219
rect 1222 214 1228 215
rect 1222 210 1223 214
rect 1227 210 1228 214
rect 1222 209 1228 210
rect 1262 214 1268 215
rect 1262 210 1263 214
rect 1267 210 1268 214
rect 1262 209 1268 210
rect 1302 214 1308 215
rect 1302 210 1303 214
rect 1307 210 1308 214
rect 1302 209 1308 210
rect 1162 203 1168 204
rect 1162 199 1163 203
rect 1167 199 1168 203
rect 1162 198 1168 199
rect 1198 203 1204 204
rect 1198 199 1199 203
rect 1203 199 1204 203
rect 1198 198 1204 199
rect 1142 197 1148 198
rect 1142 193 1143 197
rect 1147 193 1148 197
rect 1142 192 1148 193
rect 1104 175 1106 192
rect 1118 191 1124 192
rect 1118 187 1119 191
rect 1123 187 1124 191
rect 1118 186 1124 187
rect 1144 175 1146 192
rect 1103 174 1107 175
rect 1103 169 1107 170
rect 1143 174 1147 175
rect 1143 169 1147 170
rect 1151 174 1155 175
rect 1151 168 1155 170
rect 1150 167 1156 168
rect 1150 163 1151 167
rect 1155 163 1156 167
rect 1150 162 1156 163
rect 646 159 652 160
rect 646 155 647 159
rect 651 155 652 159
rect 646 154 652 155
rect 998 159 1004 160
rect 998 155 999 159
rect 1003 155 1004 159
rect 998 154 1004 155
rect 1074 159 1080 160
rect 1074 155 1075 159
rect 1079 155 1080 159
rect 1074 154 1080 155
rect 686 150 692 151
rect 686 146 687 150
rect 691 146 692 150
rect 686 145 692 146
rect 774 150 780 151
rect 774 146 775 150
rect 779 146 780 150
rect 774 145 780 146
rect 862 150 868 151
rect 862 146 863 150
rect 867 146 868 150
rect 862 145 868 146
rect 958 150 964 151
rect 958 146 959 150
rect 963 146 964 150
rect 958 145 964 146
rect 688 123 690 145
rect 776 123 778 145
rect 864 123 866 145
rect 918 143 924 144
rect 918 139 919 143
rect 923 139 924 143
rect 918 138 924 139
rect 671 122 675 123
rect 671 117 675 118
rect 687 122 691 123
rect 687 117 691 118
rect 743 122 747 123
rect 743 117 747 118
rect 775 122 779 123
rect 775 117 779 118
rect 823 122 827 123
rect 823 117 827 118
rect 863 122 867 123
rect 863 117 867 118
rect 903 122 907 123
rect 903 117 907 118
rect 672 107 674 117
rect 744 107 746 117
rect 824 107 826 117
rect 904 107 906 117
rect 670 106 676 107
rect 670 102 671 106
rect 675 102 676 106
rect 670 101 676 102
rect 742 106 748 107
rect 742 102 743 106
rect 747 102 748 106
rect 742 101 748 102
rect 822 106 828 107
rect 822 102 823 106
rect 827 102 828 106
rect 822 101 828 102
rect 902 106 908 107
rect 902 102 903 106
rect 907 102 908 106
rect 902 101 908 102
rect 920 96 922 138
rect 960 123 962 145
rect 959 122 963 123
rect 959 117 963 118
rect 983 122 987 123
rect 983 117 987 118
rect 984 107 986 117
rect 1000 112 1002 154
rect 1054 150 1060 151
rect 1054 146 1055 150
rect 1059 146 1060 150
rect 1054 145 1060 146
rect 1150 150 1156 151
rect 1150 146 1151 150
rect 1155 146 1156 150
rect 1150 145 1156 146
rect 1026 135 1032 136
rect 1026 131 1027 135
rect 1031 131 1032 135
rect 1026 130 1032 131
rect 998 111 1004 112
rect 998 107 999 111
rect 1003 107 1004 111
rect 982 106 988 107
rect 998 106 1004 107
rect 982 102 983 106
rect 987 102 988 106
rect 982 101 988 102
rect 1028 96 1030 130
rect 1056 123 1058 145
rect 1152 123 1154 145
rect 1164 144 1166 198
rect 1182 197 1188 198
rect 1182 193 1183 197
rect 1187 193 1188 197
rect 1182 192 1188 193
rect 1222 197 1228 198
rect 1222 193 1223 197
rect 1227 193 1228 197
rect 1222 192 1228 193
rect 1262 197 1268 198
rect 1262 193 1263 197
rect 1267 193 1268 197
rect 1262 192 1268 193
rect 1302 197 1308 198
rect 1302 193 1303 197
rect 1307 193 1308 197
rect 1302 192 1308 193
rect 1184 175 1186 192
rect 1224 175 1226 192
rect 1264 175 1266 192
rect 1304 175 1306 192
rect 1183 174 1187 175
rect 1183 169 1187 170
rect 1223 174 1227 175
rect 1223 169 1227 170
rect 1239 174 1243 175
rect 1239 168 1243 170
rect 1263 174 1267 175
rect 1263 169 1267 170
rect 1303 174 1307 175
rect 1303 169 1307 170
rect 1238 167 1244 168
rect 1238 163 1239 167
rect 1243 163 1244 167
rect 1238 162 1244 163
rect 1312 160 1314 218
rect 1344 215 1346 245
rect 1376 215 1378 245
rect 1408 215 1410 245
rect 1440 215 1442 245
rect 1480 215 1482 245
rect 1520 215 1522 245
rect 1532 232 1534 290
rect 1558 286 1564 287
rect 1558 282 1559 286
rect 1563 282 1564 286
rect 1558 281 1564 282
rect 1590 286 1596 287
rect 1590 282 1591 286
rect 1595 282 1596 286
rect 1590 281 1596 282
rect 1622 286 1628 287
rect 1622 282 1623 286
rect 1627 282 1628 286
rect 1622 281 1628 282
rect 1560 251 1562 281
rect 1592 251 1594 281
rect 1606 279 1612 280
rect 1606 275 1607 279
rect 1611 275 1612 279
rect 1606 274 1612 275
rect 1559 250 1563 251
rect 1559 245 1563 246
rect 1591 250 1595 251
rect 1591 245 1595 246
rect 1530 231 1536 232
rect 1530 227 1531 231
rect 1535 227 1536 231
rect 1530 226 1536 227
rect 1560 215 1562 245
rect 1592 215 1594 245
rect 1598 219 1604 220
rect 1598 215 1599 219
rect 1603 215 1604 219
rect 1342 214 1348 215
rect 1342 210 1343 214
rect 1347 210 1348 214
rect 1342 209 1348 210
rect 1374 214 1380 215
rect 1374 210 1375 214
rect 1379 210 1380 214
rect 1374 209 1380 210
rect 1406 214 1412 215
rect 1406 210 1407 214
rect 1411 210 1412 214
rect 1406 209 1412 210
rect 1438 214 1444 215
rect 1438 210 1439 214
rect 1443 210 1444 214
rect 1438 209 1444 210
rect 1478 214 1484 215
rect 1478 210 1479 214
rect 1483 210 1484 214
rect 1478 209 1484 210
rect 1518 214 1524 215
rect 1518 210 1519 214
rect 1523 210 1524 214
rect 1518 209 1524 210
rect 1558 214 1564 215
rect 1558 210 1559 214
rect 1563 210 1564 214
rect 1558 209 1564 210
rect 1590 214 1596 215
rect 1598 214 1604 215
rect 1590 210 1591 214
rect 1595 210 1596 214
rect 1590 209 1596 210
rect 1578 203 1584 204
rect 1578 199 1579 203
rect 1583 199 1584 203
rect 1578 198 1584 199
rect 1342 197 1348 198
rect 1342 193 1343 197
rect 1347 193 1348 197
rect 1342 192 1348 193
rect 1374 197 1380 198
rect 1374 193 1375 197
rect 1379 193 1380 197
rect 1374 192 1380 193
rect 1406 197 1412 198
rect 1406 193 1407 197
rect 1411 193 1412 197
rect 1406 192 1412 193
rect 1438 197 1444 198
rect 1438 193 1439 197
rect 1443 193 1444 197
rect 1438 192 1444 193
rect 1478 197 1484 198
rect 1478 193 1479 197
rect 1483 193 1484 197
rect 1478 192 1484 193
rect 1518 197 1524 198
rect 1518 193 1519 197
rect 1523 193 1524 197
rect 1518 192 1524 193
rect 1558 197 1564 198
rect 1558 193 1559 197
rect 1563 193 1564 197
rect 1558 192 1564 193
rect 1344 175 1346 192
rect 1376 175 1378 192
rect 1408 175 1410 192
rect 1440 175 1442 192
rect 1480 175 1482 192
rect 1520 175 1522 192
rect 1560 175 1562 192
rect 1327 174 1331 175
rect 1327 168 1331 170
rect 1343 174 1347 175
rect 1343 169 1347 170
rect 1375 174 1379 175
rect 1375 169 1379 170
rect 1407 174 1411 175
rect 1407 169 1411 170
rect 1415 174 1419 175
rect 1415 168 1419 170
rect 1439 174 1443 175
rect 1439 169 1443 170
rect 1479 174 1483 175
rect 1479 169 1483 170
rect 1503 174 1507 175
rect 1503 168 1507 170
rect 1519 174 1523 175
rect 1519 169 1523 170
rect 1559 174 1563 175
rect 1559 169 1563 170
rect 1326 167 1332 168
rect 1326 163 1327 167
rect 1331 163 1332 167
rect 1326 162 1332 163
rect 1414 167 1420 168
rect 1414 163 1415 167
rect 1419 163 1420 167
rect 1414 162 1420 163
rect 1502 167 1508 168
rect 1502 163 1503 167
rect 1507 163 1508 167
rect 1502 162 1508 163
rect 1310 159 1316 160
rect 1310 155 1311 159
rect 1315 155 1316 159
rect 1310 154 1316 155
rect 1534 159 1540 160
rect 1534 155 1535 159
rect 1539 155 1540 159
rect 1534 154 1540 155
rect 1542 159 1548 160
rect 1542 155 1543 159
rect 1547 155 1548 159
rect 1542 154 1548 155
rect 1238 150 1244 151
rect 1238 146 1239 150
rect 1243 146 1244 150
rect 1238 145 1244 146
rect 1326 150 1332 151
rect 1326 146 1327 150
rect 1331 146 1332 150
rect 1326 145 1332 146
rect 1414 150 1420 151
rect 1414 146 1415 150
rect 1419 146 1420 150
rect 1414 145 1420 146
rect 1502 150 1508 151
rect 1502 146 1503 150
rect 1507 146 1508 150
rect 1502 145 1508 146
rect 1162 143 1168 144
rect 1162 139 1163 143
rect 1167 139 1168 143
rect 1162 138 1168 139
rect 1194 143 1200 144
rect 1194 139 1195 143
rect 1199 139 1200 143
rect 1194 138 1200 139
rect 1055 122 1059 123
rect 1055 117 1059 118
rect 1119 122 1123 123
rect 1119 117 1123 118
rect 1151 122 1155 123
rect 1151 117 1155 118
rect 1175 122 1179 123
rect 1175 117 1179 118
rect 1056 107 1058 117
rect 1070 111 1076 112
rect 1070 107 1071 111
rect 1075 107 1076 111
rect 1120 107 1122 117
rect 1176 107 1178 117
rect 1054 106 1060 107
rect 1070 106 1076 107
rect 1118 106 1124 107
rect 1054 102 1055 106
rect 1059 102 1060 106
rect 1054 101 1060 102
rect 918 95 924 96
rect 918 91 919 95
rect 923 91 924 95
rect 918 90 924 91
rect 1026 95 1032 96
rect 1026 91 1027 95
rect 1031 91 1032 95
rect 1026 90 1032 91
rect 670 89 676 90
rect 606 84 612 85
rect 622 87 628 88
rect 111 82 115 83
rect 111 77 115 78
rect 135 82 139 84
rect 135 77 139 78
rect 167 82 171 84
rect 167 77 171 78
rect 199 82 203 84
rect 199 77 203 78
rect 231 82 235 84
rect 231 77 235 78
rect 263 82 267 84
rect 263 77 267 78
rect 295 82 299 84
rect 295 77 299 78
rect 327 82 331 84
rect 327 77 331 78
rect 359 82 363 84
rect 359 77 363 78
rect 391 82 395 84
rect 391 77 395 78
rect 423 82 427 84
rect 423 77 427 78
rect 455 82 459 84
rect 455 77 459 78
rect 487 82 491 84
rect 487 77 491 78
rect 519 82 523 84
rect 519 77 523 78
rect 551 82 555 84
rect 551 77 555 78
rect 607 82 611 84
rect 622 83 623 87
rect 627 83 628 87
rect 670 85 671 89
rect 675 85 676 89
rect 670 84 676 85
rect 742 89 748 90
rect 742 85 743 89
rect 747 85 748 89
rect 742 84 748 85
rect 822 89 828 90
rect 822 85 823 89
rect 827 85 828 89
rect 822 84 828 85
rect 902 89 908 90
rect 902 85 903 89
rect 907 85 908 89
rect 902 84 908 85
rect 982 89 988 90
rect 982 85 983 89
rect 987 85 988 89
rect 982 84 988 85
rect 1054 89 1060 90
rect 1054 85 1055 89
rect 1059 85 1060 89
rect 1054 84 1060 85
rect 1072 84 1074 106
rect 1118 102 1119 106
rect 1123 102 1124 106
rect 1118 101 1124 102
rect 1174 106 1180 107
rect 1174 102 1175 106
rect 1179 102 1180 106
rect 1174 101 1180 102
rect 1196 96 1198 138
rect 1240 123 1242 145
rect 1328 123 1330 145
rect 1416 123 1418 145
rect 1504 123 1506 145
rect 1223 122 1227 123
rect 1223 117 1227 118
rect 1239 122 1243 123
rect 1239 117 1243 118
rect 1271 122 1275 123
rect 1271 117 1275 118
rect 1311 122 1315 123
rect 1311 117 1315 118
rect 1327 122 1331 123
rect 1327 117 1331 118
rect 1343 122 1347 123
rect 1343 117 1347 118
rect 1375 122 1379 123
rect 1375 117 1379 118
rect 1407 122 1411 123
rect 1407 117 1411 118
rect 1415 122 1419 123
rect 1415 117 1419 118
rect 1439 122 1443 123
rect 1439 117 1443 118
rect 1479 122 1483 123
rect 1479 117 1483 118
rect 1503 122 1507 123
rect 1503 117 1507 118
rect 1519 122 1523 123
rect 1519 117 1523 118
rect 1224 107 1226 117
rect 1272 107 1274 117
rect 1312 107 1314 117
rect 1344 107 1346 117
rect 1376 107 1378 117
rect 1408 107 1410 117
rect 1440 107 1442 117
rect 1480 107 1482 117
rect 1520 107 1522 117
rect 1536 112 1538 154
rect 1544 136 1546 154
rect 1580 144 1582 198
rect 1590 197 1596 198
rect 1590 193 1591 197
rect 1595 193 1596 197
rect 1590 192 1596 193
rect 1592 175 1594 192
rect 1591 174 1595 175
rect 1591 168 1595 170
rect 1590 167 1596 168
rect 1590 163 1591 167
rect 1595 163 1596 167
rect 1590 162 1596 163
rect 1590 150 1596 151
rect 1590 146 1591 150
rect 1595 146 1596 150
rect 1590 145 1596 146
rect 1578 143 1584 144
rect 1578 139 1579 143
rect 1583 139 1584 143
rect 1578 138 1584 139
rect 1542 135 1548 136
rect 1542 131 1543 135
rect 1547 131 1548 135
rect 1542 130 1548 131
rect 1592 123 1594 145
rect 1559 122 1563 123
rect 1559 117 1563 118
rect 1591 122 1595 123
rect 1591 117 1595 118
rect 1534 111 1540 112
rect 1534 107 1535 111
rect 1539 107 1540 111
rect 1560 107 1562 117
rect 1592 107 1594 117
rect 1222 106 1228 107
rect 1222 102 1223 106
rect 1227 102 1228 106
rect 1222 101 1228 102
rect 1270 106 1276 107
rect 1270 102 1271 106
rect 1275 102 1276 106
rect 1270 101 1276 102
rect 1310 106 1316 107
rect 1310 102 1311 106
rect 1315 102 1316 106
rect 1310 101 1316 102
rect 1342 106 1348 107
rect 1342 102 1343 106
rect 1347 102 1348 106
rect 1342 101 1348 102
rect 1374 106 1380 107
rect 1374 102 1375 106
rect 1379 102 1380 106
rect 1374 101 1380 102
rect 1406 106 1412 107
rect 1406 102 1407 106
rect 1411 102 1412 106
rect 1406 101 1412 102
rect 1438 106 1444 107
rect 1438 102 1439 106
rect 1443 102 1444 106
rect 1438 101 1444 102
rect 1478 106 1484 107
rect 1478 102 1479 106
rect 1483 102 1484 106
rect 1478 101 1484 102
rect 1518 106 1524 107
rect 1534 106 1540 107
rect 1558 106 1564 107
rect 1518 102 1519 106
rect 1523 102 1524 106
rect 1518 101 1524 102
rect 1558 102 1559 106
rect 1563 102 1564 106
rect 1558 101 1564 102
rect 1590 106 1596 107
rect 1590 102 1591 106
rect 1595 102 1596 106
rect 1590 101 1596 102
rect 1600 96 1602 214
rect 1608 204 1610 274
rect 1624 251 1626 281
rect 1644 280 1646 346
rect 1656 323 1658 352
rect 1696 323 1698 354
rect 1655 322 1659 323
rect 1655 317 1659 318
rect 1695 322 1699 323
rect 1695 317 1699 318
rect 1656 304 1658 317
rect 1654 303 1660 304
rect 1654 299 1655 303
rect 1659 299 1660 303
rect 1696 302 1698 317
rect 1654 298 1660 299
rect 1694 301 1700 302
rect 1694 297 1695 301
rect 1699 297 1700 301
rect 1694 296 1700 297
rect 1670 295 1676 296
rect 1670 291 1671 295
rect 1675 291 1676 295
rect 1724 292 1726 359
rect 1670 290 1676 291
rect 1722 291 1728 292
rect 1654 286 1660 287
rect 1654 282 1655 286
rect 1659 282 1660 286
rect 1654 281 1660 282
rect 1642 279 1648 280
rect 1642 275 1643 279
rect 1647 275 1648 279
rect 1642 274 1648 275
rect 1656 251 1658 281
rect 1623 250 1627 251
rect 1623 245 1627 246
rect 1655 250 1659 251
rect 1655 245 1659 246
rect 1624 215 1626 245
rect 1656 215 1658 245
rect 1672 220 1674 290
rect 1722 287 1723 291
rect 1727 287 1728 291
rect 1722 286 1728 287
rect 1694 284 1700 285
rect 1694 280 1695 284
rect 1699 280 1700 284
rect 1694 279 1700 280
rect 1696 251 1698 279
rect 1695 250 1699 251
rect 1695 245 1699 246
rect 1670 219 1676 220
rect 1670 215 1671 219
rect 1675 215 1676 219
rect 1696 217 1698 245
rect 1622 214 1628 215
rect 1622 210 1623 214
rect 1627 210 1628 214
rect 1622 209 1628 210
rect 1654 214 1660 215
rect 1670 214 1676 215
rect 1694 216 1700 217
rect 1654 210 1655 214
rect 1659 210 1660 214
rect 1694 212 1695 216
rect 1699 212 1700 216
rect 1694 211 1700 212
rect 1654 209 1660 210
rect 1606 203 1612 204
rect 1606 199 1607 203
rect 1611 199 1612 203
rect 1606 198 1612 199
rect 1642 203 1648 204
rect 1642 199 1643 203
rect 1647 199 1648 203
rect 1642 198 1648 199
rect 1694 199 1700 200
rect 1622 197 1628 198
rect 1622 193 1623 197
rect 1627 193 1628 197
rect 1622 192 1628 193
rect 1624 175 1626 192
rect 1623 174 1627 175
rect 1623 169 1627 170
rect 1644 144 1646 198
rect 1654 197 1660 198
rect 1654 193 1655 197
rect 1659 193 1660 197
rect 1694 195 1695 199
rect 1699 195 1700 199
rect 1694 194 1700 195
rect 1654 192 1660 193
rect 1656 175 1658 192
rect 1696 175 1698 194
rect 1655 174 1659 175
rect 1655 168 1659 170
rect 1695 174 1699 175
rect 1695 169 1699 170
rect 1654 167 1660 168
rect 1654 163 1655 167
rect 1659 163 1660 167
rect 1696 166 1698 169
rect 1654 162 1660 163
rect 1694 165 1700 166
rect 1694 161 1695 165
rect 1699 161 1700 165
rect 1694 160 1700 161
rect 1670 159 1676 160
rect 1670 155 1671 159
rect 1675 155 1676 159
rect 1670 154 1676 155
rect 1654 150 1660 151
rect 1654 146 1655 150
rect 1659 146 1660 150
rect 1654 145 1660 146
rect 1642 143 1648 144
rect 1642 139 1643 143
rect 1647 139 1648 143
rect 1642 138 1648 139
rect 1656 123 1658 145
rect 1623 122 1627 123
rect 1623 117 1627 118
rect 1655 122 1659 123
rect 1655 117 1659 118
rect 1624 107 1626 117
rect 1656 107 1658 117
rect 1672 112 1674 154
rect 1694 148 1700 149
rect 1694 144 1695 148
rect 1699 144 1700 148
rect 1694 143 1700 144
rect 1696 123 1698 143
rect 1695 122 1699 123
rect 1695 117 1699 118
rect 1670 111 1676 112
rect 1670 107 1671 111
rect 1675 107 1676 111
rect 1696 109 1698 117
rect 1622 106 1628 107
rect 1622 102 1623 106
rect 1627 102 1628 106
rect 1622 101 1628 102
rect 1654 106 1660 107
rect 1670 106 1676 107
rect 1694 108 1700 109
rect 1654 102 1655 106
rect 1659 102 1660 106
rect 1694 104 1695 108
rect 1699 104 1700 108
rect 1694 103 1700 104
rect 1654 101 1660 102
rect 1194 95 1200 96
rect 1194 91 1195 95
rect 1199 91 1200 95
rect 1600 95 1608 96
rect 1600 92 1603 95
rect 1194 90 1200 91
rect 1602 91 1603 92
rect 1607 91 1608 95
rect 1602 90 1608 91
rect 1694 91 1700 92
rect 1118 89 1124 90
rect 1118 85 1119 89
rect 1123 85 1124 89
rect 1118 84 1124 85
rect 1174 89 1180 90
rect 1174 85 1175 89
rect 1179 85 1180 89
rect 1174 84 1180 85
rect 1222 89 1228 90
rect 1222 85 1223 89
rect 1227 85 1228 89
rect 1222 84 1228 85
rect 1270 89 1276 90
rect 1270 85 1271 89
rect 1275 85 1276 89
rect 1270 84 1276 85
rect 1310 89 1316 90
rect 1310 85 1311 89
rect 1315 85 1316 89
rect 1310 84 1316 85
rect 1342 89 1348 90
rect 1342 85 1343 89
rect 1347 85 1348 89
rect 1342 84 1348 85
rect 1374 89 1380 90
rect 1374 85 1375 89
rect 1379 85 1380 89
rect 1374 84 1380 85
rect 1406 89 1412 90
rect 1406 85 1407 89
rect 1411 85 1412 89
rect 1406 84 1412 85
rect 1438 89 1444 90
rect 1438 85 1439 89
rect 1443 85 1444 89
rect 1438 84 1444 85
rect 1478 89 1484 90
rect 1478 85 1479 89
rect 1483 85 1484 89
rect 1478 84 1484 85
rect 1518 89 1524 90
rect 1518 85 1519 89
rect 1523 85 1524 89
rect 1518 84 1524 85
rect 1558 89 1564 90
rect 1558 85 1559 89
rect 1563 85 1564 89
rect 1558 84 1564 85
rect 1590 89 1596 90
rect 1590 85 1591 89
rect 1595 85 1596 89
rect 1590 84 1596 85
rect 1622 89 1628 90
rect 1622 85 1623 89
rect 1627 85 1628 89
rect 1622 84 1628 85
rect 1654 89 1660 90
rect 1654 85 1655 89
rect 1659 85 1660 89
rect 1694 87 1695 91
rect 1699 87 1700 91
rect 1694 86 1700 87
rect 1654 84 1660 85
rect 622 82 628 83
rect 671 82 675 84
rect 607 77 611 78
rect 671 77 675 78
rect 743 82 747 84
rect 743 77 747 78
rect 823 82 827 84
rect 823 77 827 78
rect 903 82 907 84
rect 903 77 907 78
rect 983 82 987 84
rect 983 77 987 78
rect 1055 82 1059 84
rect 1070 83 1076 84
rect 1070 79 1071 83
rect 1075 79 1076 83
rect 1070 78 1076 79
rect 1119 82 1123 84
rect 1055 77 1059 78
rect 1119 77 1123 78
rect 1175 82 1179 84
rect 1175 77 1179 78
rect 1223 82 1227 84
rect 1223 77 1227 78
rect 1271 82 1275 84
rect 1271 77 1275 78
rect 1311 82 1315 84
rect 1311 77 1315 78
rect 1343 82 1347 84
rect 1343 77 1347 78
rect 1375 82 1379 84
rect 1375 77 1379 78
rect 1407 82 1411 84
rect 1407 77 1411 78
rect 1439 82 1443 84
rect 1439 77 1443 78
rect 1479 82 1483 84
rect 1479 77 1483 78
rect 1519 82 1523 84
rect 1519 77 1523 78
rect 1559 82 1563 84
rect 1559 77 1563 78
rect 1591 82 1595 84
rect 1591 77 1595 78
rect 1623 82 1627 84
rect 1623 77 1627 78
rect 1655 82 1659 84
rect 1696 83 1698 86
rect 1655 77 1659 78
rect 1695 82 1699 83
rect 1695 77 1699 78
<< m4c >>
rect 111 1758 115 1762
rect 151 1758 155 1762
rect 183 1758 187 1762
rect 215 1758 219 1762
rect 247 1758 251 1762
rect 279 1758 283 1762
rect 311 1758 315 1762
rect 343 1758 347 1762
rect 375 1758 379 1762
rect 407 1758 411 1762
rect 439 1758 443 1762
rect 471 1758 475 1762
rect 503 1758 507 1762
rect 535 1758 539 1762
rect 567 1758 571 1762
rect 599 1758 603 1762
rect 631 1758 635 1762
rect 663 1758 667 1762
rect 695 1758 699 1762
rect 727 1758 731 1762
rect 759 1758 763 1762
rect 791 1758 795 1762
rect 823 1758 827 1762
rect 855 1758 859 1762
rect 887 1758 891 1762
rect 111 1714 115 1718
rect 151 1714 155 1718
rect 183 1714 187 1718
rect 191 1714 195 1718
rect 215 1714 219 1718
rect 247 1714 251 1718
rect 279 1714 283 1718
rect 311 1714 315 1718
rect 319 1714 323 1718
rect 343 1714 347 1718
rect 375 1714 379 1718
rect 407 1714 411 1718
rect 415 1714 419 1718
rect 439 1714 443 1718
rect 471 1714 475 1718
rect 503 1714 507 1718
rect 527 1714 531 1718
rect 535 1714 539 1718
rect 567 1714 571 1718
rect 599 1714 603 1718
rect 631 1714 635 1718
rect 655 1714 659 1718
rect 663 1714 667 1718
rect 695 1714 699 1718
rect 727 1714 731 1718
rect 759 1714 763 1718
rect 791 1714 795 1718
rect 823 1714 827 1718
rect 855 1714 859 1718
rect 111 1666 115 1670
rect 135 1666 139 1670
rect 175 1666 179 1670
rect 191 1666 195 1670
rect 247 1666 251 1670
rect 263 1666 267 1670
rect 319 1666 323 1670
rect 391 1666 395 1670
rect 111 1618 115 1622
rect 135 1618 139 1622
rect 167 1618 171 1622
rect 175 1618 179 1622
rect 111 1578 115 1582
rect 135 1578 139 1582
rect 167 1578 171 1582
rect 111 1538 115 1542
rect 135 1538 139 1542
rect 167 1538 171 1542
rect 175 1538 179 1542
rect 111 1494 115 1498
rect 135 1494 139 1498
rect 175 1494 179 1498
rect 111 1426 115 1430
rect 135 1426 139 1430
rect 167 1426 171 1430
rect 175 1426 179 1430
rect 111 1346 115 1350
rect 135 1346 139 1350
rect 167 1346 171 1350
rect 111 1258 115 1262
rect 135 1258 139 1262
rect 167 1258 171 1262
rect 111 1146 115 1150
rect 135 1146 139 1150
rect 167 1146 171 1150
rect 199 1618 203 1622
rect 247 1618 251 1622
rect 263 1618 267 1622
rect 327 1618 331 1622
rect 415 1666 419 1670
rect 527 1666 531 1670
rect 543 1666 547 1670
rect 655 1666 659 1670
rect 711 1666 715 1670
rect 791 1666 795 1670
rect 391 1618 395 1622
rect 439 1618 443 1622
rect 543 1618 547 1622
rect 567 1618 571 1622
rect 711 1618 715 1622
rect 855 1618 859 1622
rect 919 1758 923 1762
rect 951 1758 955 1762
rect 983 1758 987 1762
rect 1695 1758 1699 1762
rect 887 1714 891 1718
rect 919 1714 923 1718
rect 951 1714 955 1718
rect 983 1714 987 1718
rect 1047 1714 1051 1718
rect 879 1666 883 1670
rect 1159 1714 1163 1718
rect 919 1666 923 1670
rect 1039 1666 1043 1670
rect 1047 1666 1051 1670
rect 1159 1666 1163 1670
rect 1183 1666 1187 1670
rect 879 1618 883 1622
rect 999 1618 1003 1622
rect 199 1578 203 1582
rect 231 1578 235 1582
rect 247 1578 251 1582
rect 287 1578 291 1582
rect 327 1578 331 1582
rect 343 1578 347 1582
rect 399 1578 403 1582
rect 439 1578 443 1582
rect 455 1578 459 1582
rect 511 1578 515 1582
rect 567 1578 571 1582
rect 575 1578 579 1582
rect 655 1578 659 1582
rect 711 1578 715 1582
rect 751 1578 755 1582
rect 855 1578 859 1582
rect 223 1538 227 1542
rect 231 1538 235 1542
rect 279 1538 283 1542
rect 287 1538 291 1542
rect 335 1538 339 1542
rect 343 1538 347 1542
rect 399 1538 403 1542
rect 455 1538 459 1542
rect 463 1538 467 1542
rect 511 1538 515 1542
rect 535 1538 539 1542
rect 575 1538 579 1542
rect 207 1494 211 1498
rect 223 1494 227 1498
rect 239 1494 243 1498
rect 271 1494 275 1498
rect 279 1494 283 1498
rect 303 1494 307 1498
rect 335 1494 339 1498
rect 367 1494 371 1498
rect 399 1494 403 1498
rect 431 1494 435 1498
rect 463 1494 467 1498
rect 607 1538 611 1542
rect 655 1538 659 1542
rect 687 1538 691 1542
rect 495 1494 499 1498
rect 527 1494 531 1498
rect 535 1494 539 1498
rect 559 1494 563 1498
rect 591 1494 595 1498
rect 607 1494 611 1498
rect 623 1494 627 1498
rect 751 1538 755 1542
rect 663 1494 667 1498
rect 687 1494 691 1498
rect 703 1494 707 1498
rect 199 1426 203 1430
rect 207 1426 211 1430
rect 231 1426 235 1430
rect 239 1426 243 1430
rect 263 1426 267 1430
rect 271 1426 275 1430
rect 295 1426 299 1430
rect 303 1426 307 1430
rect 327 1426 331 1430
rect 335 1426 339 1430
rect 359 1426 363 1430
rect 367 1426 371 1430
rect 391 1426 395 1430
rect 399 1426 403 1430
rect 423 1426 427 1430
rect 431 1426 435 1430
rect 455 1426 459 1430
rect 463 1426 467 1430
rect 487 1426 491 1430
rect 495 1426 499 1430
rect 519 1426 523 1430
rect 527 1426 531 1430
rect 551 1426 555 1430
rect 559 1426 563 1430
rect 583 1426 587 1430
rect 591 1426 595 1430
rect 615 1426 619 1430
rect 623 1426 627 1430
rect 647 1426 651 1430
rect 663 1426 667 1430
rect 679 1426 683 1430
rect 199 1346 203 1350
rect 231 1346 235 1350
rect 263 1346 267 1350
rect 295 1346 299 1350
rect 327 1346 331 1350
rect 359 1346 363 1350
rect 391 1346 395 1350
rect 423 1346 427 1350
rect 455 1346 459 1350
rect 487 1346 491 1350
rect 519 1346 523 1350
rect 551 1346 555 1350
rect 583 1346 587 1350
rect 615 1346 619 1350
rect 647 1346 651 1350
rect 199 1258 203 1262
rect 231 1258 235 1262
rect 263 1258 267 1262
rect 295 1258 299 1262
rect 327 1258 331 1262
rect 359 1258 363 1262
rect 391 1258 395 1262
rect 423 1258 427 1262
rect 455 1258 459 1262
rect 487 1258 491 1262
rect 519 1258 523 1262
rect 551 1258 555 1262
rect 199 1146 203 1150
rect 231 1146 235 1150
rect 263 1146 267 1150
rect 295 1146 299 1150
rect 327 1146 331 1150
rect 359 1146 363 1150
rect 391 1146 395 1150
rect 423 1146 427 1150
rect 187 1056 191 1060
rect 179 1040 183 1044
rect 111 1030 115 1034
rect 135 1030 139 1034
rect 167 1030 171 1034
rect 111 950 115 954
rect 135 950 139 954
rect 167 950 171 954
rect 199 1030 203 1034
rect 231 1030 235 1034
rect 263 1030 267 1034
rect 295 1030 299 1034
rect 199 950 203 954
rect 231 950 235 954
rect 111 834 115 838
rect 135 834 139 838
rect 167 834 171 838
rect 111 750 115 754
rect 135 750 139 754
rect 111 638 115 642
rect 135 638 139 642
rect 143 638 147 642
rect 167 638 171 642
rect 263 950 267 954
rect 279 950 283 954
rect 383 1088 387 1092
rect 327 1030 331 1034
rect 359 1030 363 1034
rect 399 1040 403 1044
rect 391 1030 395 1034
rect 407 1030 411 1034
rect 455 1146 459 1150
rect 487 1146 491 1150
rect 519 1146 523 1150
rect 423 1030 427 1034
rect 455 1030 459 1034
rect 487 1030 491 1034
rect 503 1030 507 1034
rect 519 1030 523 1034
rect 319 950 323 954
rect 343 950 347 954
rect 207 834 211 838
rect 231 834 235 838
rect 279 834 283 838
rect 327 834 331 838
rect 215 750 219 754
rect 231 750 235 754
rect 287 750 291 754
rect 111 558 115 562
rect 135 558 139 562
rect 167 558 171 562
rect 207 638 211 642
rect 215 638 219 642
rect 287 638 291 642
rect 207 558 211 562
rect 247 558 251 562
rect 111 438 115 442
rect 135 438 139 442
rect 167 438 171 442
rect 175 438 179 442
rect 199 438 203 442
rect 231 438 235 442
rect 247 438 251 442
rect 279 558 283 562
rect 303 558 307 562
rect 263 438 267 442
rect 399 950 403 954
rect 551 1146 555 1150
rect 551 1030 555 1034
rect 463 950 467 954
rect 503 950 507 954
rect 399 834 403 838
rect 407 834 411 838
rect 391 750 395 754
rect 407 750 411 754
rect 435 834 439 838
rect 391 638 395 642
rect 471 750 475 754
rect 583 1258 587 1262
rect 615 1258 619 1262
rect 583 1146 587 1150
rect 647 1258 651 1262
rect 615 1146 619 1150
rect 647 1146 651 1150
rect 583 1030 587 1034
rect 591 1030 595 1034
rect 583 950 587 954
rect 591 950 595 954
rect 743 1494 747 1498
rect 703 1426 707 1430
rect 719 1426 723 1430
rect 743 1426 747 1430
rect 679 1346 683 1350
rect 711 1346 715 1350
rect 735 1346 739 1350
rect 743 1346 747 1350
rect 775 1538 779 1542
rect 855 1538 859 1542
rect 871 1538 875 1542
rect 775 1494 779 1498
rect 807 1494 811 1498
rect 871 1494 875 1498
rect 767 1426 771 1430
rect 775 1426 779 1430
rect 807 1426 811 1430
rect 767 1346 771 1350
rect 679 1258 683 1262
rect 711 1258 715 1262
rect 743 1258 747 1262
rect 751 1258 755 1262
rect 775 1258 779 1262
rect 839 1426 843 1430
rect 807 1346 811 1350
rect 823 1346 827 1350
rect 959 1578 963 1582
rect 1039 1618 1043 1622
rect 1127 1618 1131 1622
rect 1183 1618 1187 1622
rect 999 1578 1003 1582
rect 1063 1578 1067 1582
rect 1127 1578 1131 1582
rect 1159 1578 1163 1582
rect 1255 1714 1259 1718
rect 1335 1714 1339 1718
rect 1407 1714 1411 1718
rect 1463 1714 1467 1718
rect 1519 1714 1523 1718
rect 1567 1714 1571 1718
rect 1623 1714 1627 1718
rect 1655 1714 1659 1718
rect 1695 1714 1699 1718
rect 1255 1666 1259 1670
rect 1319 1666 1323 1670
rect 1335 1666 1339 1670
rect 1407 1666 1411 1670
rect 1439 1666 1443 1670
rect 1463 1666 1467 1670
rect 1247 1618 1251 1622
rect 1319 1618 1323 1622
rect 1359 1618 1363 1622
rect 1519 1666 1523 1670
rect 1559 1666 1563 1670
rect 1567 1666 1571 1670
rect 1623 1666 1627 1670
rect 1655 1666 1659 1670
rect 1695 1666 1699 1670
rect 1439 1618 1443 1622
rect 1463 1618 1467 1622
rect 1559 1618 1563 1622
rect 1567 1618 1571 1622
rect 1655 1618 1659 1622
rect 1695 1618 1699 1622
rect 1247 1578 1251 1582
rect 1327 1578 1331 1582
rect 959 1538 963 1542
rect 975 1538 979 1542
rect 1063 1538 1067 1542
rect 895 1494 899 1498
rect 935 1494 939 1498
rect 975 1494 979 1498
rect 1023 1494 1027 1498
rect 1079 1538 1083 1542
rect 1079 1494 1083 1498
rect 1159 1538 1163 1542
rect 1175 1538 1179 1542
rect 1359 1578 1363 1582
rect 1399 1578 1403 1582
rect 1463 1578 1467 1582
rect 1471 1578 1475 1582
rect 1247 1538 1251 1542
rect 1271 1538 1275 1542
rect 1327 1538 1331 1542
rect 1359 1538 1363 1542
rect 1111 1494 1115 1498
rect 1167 1494 1171 1498
rect 1175 1494 1179 1498
rect 1199 1494 1203 1498
rect 895 1426 899 1430
rect 935 1426 939 1430
rect 975 1426 979 1430
rect 1023 1426 1027 1430
rect 911 1416 915 1420
rect 839 1346 843 1350
rect 811 1258 815 1262
rect 831 1258 835 1262
rect 679 1146 683 1150
rect 687 1146 691 1150
rect 711 1146 715 1150
rect 743 1146 747 1150
rect 775 1146 779 1150
rect 671 1088 675 1092
rect 659 1030 663 1034
rect 679 950 683 954
rect 559 834 563 838
rect 591 834 595 838
rect 663 834 667 838
rect 679 834 683 838
rect 711 1030 715 1034
rect 887 1346 891 1350
rect 903 1346 907 1350
rect 911 1258 915 1262
rect 991 1419 995 1420
rect 991 1416 995 1419
rect 1039 1426 1043 1430
rect 1063 1426 1067 1430
rect 1079 1426 1083 1430
rect 1111 1426 1115 1430
rect 1127 1426 1131 1430
rect 799 1146 803 1150
rect 839 1146 843 1150
rect 847 1146 851 1150
rect 815 1056 819 1060
rect 799 1030 803 1034
rect 823 1030 827 1034
rect 847 1030 851 1034
rect 711 950 715 954
rect 727 950 731 954
rect 815 950 819 954
rect 727 834 731 838
rect 559 750 563 754
rect 615 750 619 754
rect 655 750 659 754
rect 719 750 723 754
rect 407 638 411 642
rect 443 638 447 642
rect 535 638 539 642
rect 391 558 395 562
rect 399 558 403 562
rect 303 438 307 442
rect 375 438 379 442
rect 471 558 475 562
rect 399 438 403 442
rect 415 438 419 442
rect 447 438 451 442
rect 471 438 475 442
rect 487 438 491 442
rect 507 438 511 442
rect 535 558 539 562
rect 623 680 627 684
rect 615 638 619 642
rect 671 638 675 642
rect 719 638 723 642
rect 815 834 819 838
rect 975 1346 979 1350
rect 983 1346 987 1350
rect 1023 1346 1027 1350
rect 1063 1346 1067 1350
rect 1111 1346 1115 1350
rect 1151 1426 1155 1430
rect 1167 1426 1171 1430
rect 1151 1346 1155 1350
rect 1159 1346 1163 1350
rect 1155 1275 1159 1276
rect 1155 1272 1159 1275
rect 959 1258 963 1262
rect 983 1258 987 1262
rect 1015 1258 1019 1262
rect 1023 1258 1027 1262
rect 1063 1258 1067 1262
rect 1087 1258 1091 1262
rect 1127 1258 1131 1262
rect 1159 1258 1163 1262
rect 1175 1258 1179 1262
rect 935 1146 939 1150
rect 967 1146 971 1150
rect 975 1146 979 1150
rect 999 1146 1003 1150
rect 1007 1146 1011 1150
rect 1031 1146 1035 1150
rect 919 1030 923 1034
rect 935 1030 939 1034
rect 967 1030 971 1034
rect 975 1030 979 1034
rect 999 1030 1003 1034
rect 1063 1146 1067 1150
rect 1087 1146 1091 1150
rect 1095 1146 1099 1150
rect 1075 1088 1079 1092
rect 1031 1030 1035 1034
rect 1063 1030 1067 1034
rect 863 950 867 954
rect 919 950 923 954
rect 951 950 955 954
rect 967 950 971 954
rect 983 950 987 954
rect 1039 950 1043 954
rect 767 750 771 754
rect 815 750 819 754
rect 767 638 771 642
rect 775 638 779 642
rect 863 834 867 838
rect 951 834 955 838
rect 1127 1146 1131 1150
rect 1135 1146 1139 1150
rect 1159 1146 1163 1150
rect 1167 1146 1171 1150
rect 1095 1030 1099 1034
rect 1119 1030 1123 1034
rect 1135 1030 1139 1034
rect 1167 1030 1171 1034
rect 1175 1030 1179 1034
rect 1239 1494 1243 1498
rect 1399 1538 1403 1542
rect 1439 1538 1443 1542
rect 1471 1538 1475 1542
rect 1271 1494 1275 1498
rect 1279 1494 1283 1498
rect 1319 1494 1323 1498
rect 1199 1426 1203 1430
rect 1239 1426 1243 1430
rect 1263 1426 1267 1430
rect 1279 1426 1283 1430
rect 1359 1494 1363 1498
rect 1399 1494 1403 1498
rect 1439 1494 1443 1498
rect 1319 1426 1323 1430
rect 1359 1426 1363 1430
rect 1399 1426 1403 1430
rect 1415 1426 1419 1430
rect 1439 1426 1443 1430
rect 1199 1346 1203 1350
rect 1215 1346 1219 1350
rect 1247 1346 1251 1350
rect 1303 1346 1307 1350
rect 1319 1346 1323 1350
rect 1391 1346 1395 1350
rect 1215 1258 1219 1262
rect 1199 1211 1203 1212
rect 1199 1208 1203 1211
rect 1535 1578 1539 1582
rect 1567 1578 1571 1582
rect 1607 1578 1611 1582
rect 1519 1538 1523 1542
rect 1535 1538 1539 1542
rect 1655 1578 1659 1582
rect 1695 1578 1699 1582
rect 1599 1538 1603 1542
rect 1607 1538 1611 1542
rect 1655 1538 1659 1542
rect 1695 1538 1699 1542
rect 1479 1494 1483 1498
rect 1519 1494 1523 1498
rect 1559 1494 1563 1498
rect 1591 1494 1595 1498
rect 1599 1494 1603 1498
rect 1623 1494 1627 1498
rect 1479 1426 1483 1430
rect 1519 1426 1523 1430
rect 1535 1426 1539 1430
rect 1415 1346 1419 1350
rect 1423 1346 1427 1350
rect 1455 1346 1459 1350
rect 1463 1346 1467 1350
rect 1255 1258 1259 1262
rect 1295 1258 1299 1262
rect 1303 1258 1307 1262
rect 1343 1258 1347 1262
rect 1375 1258 1379 1262
rect 1391 1258 1395 1262
rect 1407 1258 1411 1262
rect 1423 1258 1427 1262
rect 1199 1146 1203 1150
rect 1247 1146 1251 1150
rect 1255 1146 1259 1150
rect 1287 1146 1291 1150
rect 1311 1146 1315 1150
rect 1335 1146 1339 1150
rect 1343 1146 1347 1150
rect 1199 1030 1203 1034
rect 1247 1030 1251 1034
rect 1439 1258 1443 1262
rect 1559 1426 1563 1430
rect 1655 1494 1659 1498
rect 1695 1494 1699 1498
rect 1583 1426 1587 1430
rect 1591 1426 1595 1430
rect 1623 1426 1627 1430
rect 1655 1426 1659 1430
rect 1695 1426 1699 1430
rect 1495 1346 1499 1350
rect 1527 1346 1531 1350
rect 1535 1346 1539 1350
rect 1515 1272 1519 1276
rect 1455 1258 1459 1262
rect 1479 1258 1483 1262
rect 1495 1258 1499 1262
rect 1519 1258 1523 1262
rect 1527 1258 1531 1262
rect 1559 1346 1563 1350
rect 1583 1346 1587 1350
rect 1591 1346 1595 1350
rect 1623 1346 1627 1350
rect 1655 1346 1659 1350
rect 1695 1346 1699 1350
rect 1559 1258 1563 1262
rect 1591 1258 1595 1262
rect 1623 1258 1627 1262
rect 1655 1258 1659 1262
rect 1375 1146 1379 1150
rect 1407 1146 1411 1150
rect 1423 1146 1427 1150
rect 1439 1146 1443 1150
rect 1455 1146 1459 1150
rect 1479 1146 1483 1150
rect 1487 1146 1491 1150
rect 1695 1258 1699 1262
rect 1519 1146 1523 1150
rect 1559 1146 1563 1150
rect 1287 1030 1291 1034
rect 1295 1030 1299 1034
rect 1327 1030 1331 1034
rect 1335 1030 1339 1034
rect 1367 1030 1371 1034
rect 1407 1030 1411 1034
rect 1423 1030 1427 1034
rect 1439 1030 1443 1034
rect 1063 950 1067 954
rect 1071 950 1075 954
rect 1111 950 1115 954
rect 1135 950 1139 954
rect 1143 950 1147 954
rect 1167 950 1171 954
rect 1199 950 1203 954
rect 1239 950 1243 954
rect 1263 950 1267 954
rect 1271 950 1275 954
rect 1295 950 1299 954
rect 1327 950 1331 954
rect 1367 950 1371 954
rect 999 834 1003 838
rect 1031 834 1035 838
rect 1039 834 1043 838
rect 1071 834 1075 838
rect 1055 808 1059 812
rect 863 750 867 754
rect 911 750 915 754
rect 951 750 955 754
rect 999 750 1003 754
rect 1015 750 1019 754
rect 647 558 651 562
rect 671 558 675 562
rect 727 558 731 562
rect 767 558 771 562
rect 775 558 779 562
rect 111 318 115 322
rect 135 318 139 322
rect 83 304 87 308
rect 167 318 171 322
rect 199 318 203 322
rect 231 318 235 322
rect 263 318 267 322
rect 295 318 299 322
rect 327 318 331 322
rect 359 318 363 322
rect 375 318 379 322
rect 391 318 395 322
rect 415 318 419 322
rect 423 318 427 322
rect 111 246 115 250
rect 135 246 139 250
rect 167 246 171 250
rect 183 246 187 250
rect 199 246 203 250
rect 215 246 219 250
rect 231 246 235 250
rect 247 246 251 250
rect 263 246 267 250
rect 279 246 283 250
rect 295 246 299 250
rect 311 246 315 250
rect 327 246 331 250
rect 343 246 347 250
rect 359 246 363 250
rect 543 438 547 442
rect 447 318 451 322
rect 455 318 459 322
rect 487 318 491 322
rect 503 318 507 322
rect 519 318 523 322
rect 535 318 539 322
rect 551 318 555 322
rect 527 304 531 308
rect 599 318 603 322
rect 375 246 379 250
rect 391 246 395 250
rect 407 246 411 250
rect 423 246 427 250
rect 439 246 443 250
rect 455 246 459 250
rect 471 246 475 250
rect 487 246 491 250
rect 503 246 507 250
rect 519 246 523 250
rect 535 246 539 250
rect 551 246 555 250
rect 567 246 571 250
rect 615 438 619 442
rect 655 438 659 442
rect 671 438 675 442
rect 615 318 619 322
rect 671 318 675 322
rect 607 256 611 260
rect 599 246 603 250
rect 727 438 731 442
rect 755 438 759 442
rect 703 318 707 322
rect 639 246 643 250
rect 111 170 115 174
rect 135 170 139 174
rect 167 170 171 174
rect 183 170 187 174
rect 215 170 219 174
rect 247 170 251 174
rect 263 170 267 174
rect 279 170 283 174
rect 311 170 315 174
rect 343 170 347 174
rect 367 170 371 174
rect 375 170 379 174
rect 407 170 411 174
rect 415 170 419 174
rect 439 170 443 174
rect 471 170 475 174
rect 503 170 507 174
rect 535 170 539 174
rect 567 170 571 174
rect 599 170 603 174
rect 607 170 611 174
rect 111 118 115 122
rect 135 118 139 122
rect 167 118 171 122
rect 199 118 203 122
rect 215 118 219 122
rect 231 118 235 122
rect 263 118 267 122
rect 295 118 299 122
rect 311 118 315 122
rect 327 118 331 122
rect 359 118 363 122
rect 367 118 371 122
rect 391 118 395 122
rect 415 118 419 122
rect 423 118 427 122
rect 455 118 459 122
rect 471 118 475 122
rect 487 118 491 122
rect 519 118 523 122
rect 535 118 539 122
rect 551 118 555 122
rect 607 118 611 122
rect 695 246 699 250
rect 703 246 707 250
rect 639 170 643 174
rect 783 438 787 442
rect 783 318 787 322
rect 807 318 811 322
rect 791 246 795 250
rect 807 246 811 250
rect 839 246 843 250
rect 983 680 987 684
rect 863 638 867 642
rect 903 638 907 642
rect 911 638 915 642
rect 999 638 1003 642
rect 1007 638 1011 642
rect 871 558 875 562
rect 903 558 907 562
rect 927 558 931 562
rect 871 438 875 442
rect 903 438 907 442
rect 935 438 939 442
rect 951 438 955 442
rect 991 558 995 562
rect 1031 558 1035 562
rect 1031 438 1035 442
rect 1103 834 1107 838
rect 1111 834 1115 838
rect 1143 834 1147 838
rect 1167 834 1171 838
rect 1239 834 1243 838
rect 1247 834 1251 838
rect 1271 834 1275 838
rect 1087 750 1091 754
rect 1103 750 1107 754
rect 1295 834 1299 838
rect 1327 834 1331 838
rect 1167 750 1171 754
rect 1183 750 1187 754
rect 1207 750 1211 754
rect 1231 750 1235 754
rect 1247 750 1251 754
rect 1095 638 1099 642
rect 1119 638 1123 642
rect 1167 638 1171 642
rect 1095 558 1099 562
rect 1119 558 1123 562
rect 1075 438 1079 442
rect 1103 438 1107 442
rect 1207 638 1211 642
rect 1215 638 1219 642
rect 1199 558 1203 562
rect 1207 558 1211 562
rect 1199 438 1203 442
rect 983 360 987 364
rect 903 318 907 322
rect 911 318 915 322
rect 943 318 947 322
rect 999 318 1003 322
rect 1031 318 1035 322
rect 1047 318 1051 322
rect 1063 318 1067 322
rect 1103 318 1107 322
rect 1111 318 1115 322
rect 927 256 931 260
rect 911 246 915 250
rect 919 246 923 250
rect 967 246 971 250
rect 999 246 1003 250
rect 1031 246 1035 250
rect 1063 246 1067 250
rect 687 170 691 174
rect 695 170 699 174
rect 775 170 779 174
rect 791 170 795 174
rect 831 170 835 174
rect 863 170 867 174
rect 919 170 923 174
rect 959 170 963 174
rect 967 170 971 174
rect 1055 170 1059 174
rect 1063 170 1067 174
rect 1391 950 1395 954
rect 1407 950 1411 954
rect 1423 950 1427 954
rect 1375 834 1379 838
rect 1439 950 1443 954
rect 1423 834 1427 838
rect 1271 795 1275 796
rect 1271 792 1275 795
rect 1279 750 1283 754
rect 1295 750 1299 754
rect 1311 750 1315 754
rect 1327 750 1331 754
rect 1343 750 1347 754
rect 1375 750 1379 754
rect 1407 750 1411 754
rect 1423 750 1427 754
rect 1439 750 1443 754
rect 1455 1030 1459 1034
rect 1479 1030 1483 1034
rect 1487 1030 1491 1034
rect 1519 1030 1523 1034
rect 1591 1146 1595 1150
rect 1623 1146 1627 1150
rect 1655 1146 1659 1150
rect 1695 1146 1699 1150
rect 1559 1030 1563 1034
rect 1591 1030 1595 1034
rect 1623 1030 1627 1034
rect 1655 1030 1659 1034
rect 1695 1030 1699 1034
rect 1455 950 1459 954
rect 1479 950 1483 954
rect 1471 834 1475 838
rect 1519 950 1523 954
rect 1559 950 1563 954
rect 1591 950 1595 954
rect 1623 950 1627 954
rect 1655 950 1659 954
rect 1695 950 1699 954
rect 1663 883 1667 884
rect 1663 880 1667 883
rect 1519 834 1523 838
rect 1559 834 1563 838
rect 1591 834 1595 838
rect 1623 834 1627 838
rect 1655 834 1659 838
rect 1695 834 1699 838
rect 1471 750 1475 754
rect 1479 750 1483 754
rect 1247 638 1251 642
rect 1279 638 1283 642
rect 1311 638 1315 642
rect 1335 638 1339 642
rect 1343 638 1347 642
rect 1375 638 1379 642
rect 1407 638 1411 642
rect 1415 638 1419 642
rect 1439 638 1443 642
rect 1287 558 1291 562
rect 1335 558 1339 562
rect 1231 438 1235 442
rect 1259 438 1263 442
rect 1415 558 1419 562
rect 1423 558 1427 562
rect 1519 750 1523 754
rect 1559 750 1563 754
rect 1591 750 1595 754
rect 1623 750 1627 754
rect 1655 750 1659 754
rect 1695 750 1699 754
rect 1479 638 1483 642
rect 1519 638 1523 642
rect 1543 638 1547 642
rect 1559 638 1563 642
rect 1591 638 1595 642
rect 1607 638 1611 642
rect 1623 638 1627 642
rect 1655 638 1659 642
rect 1695 638 1699 642
rect 1479 558 1483 562
rect 1527 558 1531 562
rect 1543 558 1547 562
rect 1575 558 1579 562
rect 1607 558 1611 562
rect 1623 558 1627 562
rect 1655 558 1659 562
rect 1319 438 1323 442
rect 1359 438 1363 442
rect 1423 438 1427 442
rect 1439 438 1443 442
rect 1479 438 1483 442
rect 1519 438 1523 442
rect 1527 438 1531 442
rect 1559 438 1563 442
rect 1575 438 1579 442
rect 1199 318 1203 322
rect 1231 318 1235 322
rect 1287 318 1291 322
rect 1319 318 1323 322
rect 1103 246 1107 250
rect 1111 246 1115 250
rect 1351 318 1355 322
rect 1383 318 1387 322
rect 1415 318 1419 322
rect 1439 318 1443 322
rect 1447 318 1451 322
rect 1479 318 1483 322
rect 1591 438 1595 442
rect 1695 558 1699 562
rect 1623 438 1627 442
rect 1655 438 1659 442
rect 1695 438 1699 442
rect 1723 360 1727 364
rect 1519 318 1523 322
rect 1559 318 1563 322
rect 1591 318 1595 322
rect 1623 318 1627 322
rect 1143 246 1147 250
rect 1183 246 1187 250
rect 1207 246 1211 250
rect 1223 246 1227 250
rect 1263 246 1267 250
rect 1287 246 1291 250
rect 1303 246 1307 250
rect 1319 246 1323 250
rect 1343 246 1347 250
rect 1351 246 1355 250
rect 1375 246 1379 250
rect 1383 246 1387 250
rect 1407 246 1411 250
rect 1415 246 1419 250
rect 1439 246 1443 250
rect 1447 246 1451 250
rect 1479 246 1483 250
rect 1519 246 1523 250
rect 1103 170 1107 174
rect 1143 170 1147 174
rect 1151 170 1155 174
rect 671 118 675 122
rect 687 118 691 122
rect 743 118 747 122
rect 775 118 779 122
rect 823 118 827 122
rect 863 118 867 122
rect 903 118 907 122
rect 959 118 963 122
rect 983 118 987 122
rect 1183 170 1187 174
rect 1223 170 1227 174
rect 1239 170 1243 174
rect 1263 170 1267 174
rect 1303 170 1307 174
rect 1559 246 1563 250
rect 1591 246 1595 250
rect 1327 170 1331 174
rect 1343 170 1347 174
rect 1375 170 1379 174
rect 1407 170 1411 174
rect 1415 170 1419 174
rect 1439 170 1443 174
rect 1479 170 1483 174
rect 1503 170 1507 174
rect 1519 170 1523 174
rect 1559 170 1563 174
rect 1055 118 1059 122
rect 1119 118 1123 122
rect 1151 118 1155 122
rect 1175 118 1179 122
rect 111 78 115 82
rect 135 78 139 82
rect 167 78 171 82
rect 199 78 203 82
rect 231 78 235 82
rect 263 78 267 82
rect 295 78 299 82
rect 327 78 331 82
rect 359 78 363 82
rect 391 78 395 82
rect 423 78 427 82
rect 455 78 459 82
rect 487 78 491 82
rect 519 78 523 82
rect 551 78 555 82
rect 1223 118 1227 122
rect 1239 118 1243 122
rect 1271 118 1275 122
rect 1311 118 1315 122
rect 1327 118 1331 122
rect 1343 118 1347 122
rect 1375 118 1379 122
rect 1407 118 1411 122
rect 1415 118 1419 122
rect 1439 118 1443 122
rect 1479 118 1483 122
rect 1503 118 1507 122
rect 1519 118 1523 122
rect 1591 170 1595 174
rect 1559 118 1563 122
rect 1591 118 1595 122
rect 1655 318 1659 322
rect 1695 318 1699 322
rect 1623 246 1627 250
rect 1655 246 1659 250
rect 1695 246 1699 250
rect 1623 170 1627 174
rect 1655 170 1659 174
rect 1695 170 1699 174
rect 1623 118 1627 122
rect 1655 118 1659 122
rect 1695 118 1699 122
rect 607 78 611 82
rect 671 78 675 82
rect 743 78 747 82
rect 823 78 827 82
rect 903 78 907 82
rect 983 78 987 82
rect 1055 78 1059 82
rect 1119 78 1123 82
rect 1175 78 1179 82
rect 1223 78 1227 82
rect 1271 78 1275 82
rect 1311 78 1315 82
rect 1343 78 1347 82
rect 1375 78 1379 82
rect 1407 78 1411 82
rect 1439 78 1443 82
rect 1479 78 1483 82
rect 1519 78 1523 82
rect 1559 78 1563 82
rect 1591 78 1595 82
rect 1623 78 1627 82
rect 1655 78 1659 82
rect 1695 78 1699 82
<< m4 >>
rect 84 1757 85 1763
rect 91 1762 1719 1763
rect 91 1758 111 1762
rect 115 1758 151 1762
rect 155 1758 183 1762
rect 187 1758 215 1762
rect 219 1758 247 1762
rect 251 1758 279 1762
rect 283 1758 311 1762
rect 315 1758 343 1762
rect 347 1758 375 1762
rect 379 1758 407 1762
rect 411 1758 439 1762
rect 443 1758 471 1762
rect 475 1758 503 1762
rect 507 1758 535 1762
rect 539 1758 567 1762
rect 571 1758 599 1762
rect 603 1758 631 1762
rect 635 1758 663 1762
rect 667 1758 695 1762
rect 699 1758 727 1762
rect 731 1758 759 1762
rect 763 1758 791 1762
rect 795 1758 823 1762
rect 827 1758 855 1762
rect 859 1758 887 1762
rect 891 1758 919 1762
rect 923 1758 951 1762
rect 955 1758 983 1762
rect 987 1758 1695 1762
rect 1699 1758 1719 1762
rect 91 1757 1719 1758
rect 1725 1757 1726 1763
rect 96 1713 97 1719
rect 103 1718 1731 1719
rect 103 1714 111 1718
rect 115 1714 151 1718
rect 155 1714 183 1718
rect 187 1714 191 1718
rect 195 1714 215 1718
rect 219 1714 247 1718
rect 251 1714 279 1718
rect 283 1714 311 1718
rect 315 1714 319 1718
rect 323 1714 343 1718
rect 347 1714 375 1718
rect 379 1714 407 1718
rect 411 1714 415 1718
rect 419 1714 439 1718
rect 443 1714 471 1718
rect 475 1714 503 1718
rect 507 1714 527 1718
rect 531 1714 535 1718
rect 539 1714 567 1718
rect 571 1714 599 1718
rect 603 1714 631 1718
rect 635 1714 655 1718
rect 659 1714 663 1718
rect 667 1714 695 1718
rect 699 1714 727 1718
rect 731 1714 759 1718
rect 763 1714 791 1718
rect 795 1714 823 1718
rect 827 1714 855 1718
rect 859 1714 887 1718
rect 891 1714 919 1718
rect 923 1714 951 1718
rect 955 1714 983 1718
rect 987 1714 1047 1718
rect 1051 1714 1159 1718
rect 1163 1714 1255 1718
rect 1259 1714 1335 1718
rect 1339 1714 1407 1718
rect 1411 1714 1463 1718
rect 1467 1714 1519 1718
rect 1523 1714 1567 1718
rect 1571 1714 1623 1718
rect 1627 1714 1655 1718
rect 1659 1714 1695 1718
rect 1699 1714 1731 1718
rect 103 1713 1731 1714
rect 1737 1713 1738 1719
rect 84 1665 85 1671
rect 91 1670 1719 1671
rect 91 1666 111 1670
rect 115 1666 135 1670
rect 139 1666 175 1670
rect 179 1666 191 1670
rect 195 1666 247 1670
rect 251 1666 263 1670
rect 267 1666 319 1670
rect 323 1666 391 1670
rect 395 1666 415 1670
rect 419 1666 527 1670
rect 531 1666 543 1670
rect 547 1666 655 1670
rect 659 1666 711 1670
rect 715 1666 791 1670
rect 795 1666 879 1670
rect 883 1666 919 1670
rect 923 1666 1039 1670
rect 1043 1666 1047 1670
rect 1051 1666 1159 1670
rect 1163 1666 1183 1670
rect 1187 1666 1255 1670
rect 1259 1666 1319 1670
rect 1323 1666 1335 1670
rect 1339 1666 1407 1670
rect 1411 1666 1439 1670
rect 1443 1666 1463 1670
rect 1467 1666 1519 1670
rect 1523 1666 1559 1670
rect 1563 1666 1567 1670
rect 1571 1666 1623 1670
rect 1627 1666 1655 1670
rect 1659 1666 1695 1670
rect 1699 1666 1719 1670
rect 91 1665 1719 1666
rect 1725 1665 1726 1671
rect 96 1617 97 1623
rect 103 1622 1731 1623
rect 103 1618 111 1622
rect 115 1618 135 1622
rect 139 1618 167 1622
rect 171 1618 175 1622
rect 179 1618 199 1622
rect 203 1618 247 1622
rect 251 1618 263 1622
rect 267 1618 327 1622
rect 331 1618 391 1622
rect 395 1618 439 1622
rect 443 1618 543 1622
rect 547 1618 567 1622
rect 571 1618 711 1622
rect 715 1618 855 1622
rect 859 1618 879 1622
rect 883 1618 999 1622
rect 1003 1618 1039 1622
rect 1043 1618 1127 1622
rect 1131 1618 1183 1622
rect 1187 1618 1247 1622
rect 1251 1618 1319 1622
rect 1323 1618 1359 1622
rect 1363 1618 1439 1622
rect 1443 1618 1463 1622
rect 1467 1618 1559 1622
rect 1563 1618 1567 1622
rect 1571 1618 1655 1622
rect 1659 1618 1695 1622
rect 1699 1618 1731 1622
rect 103 1617 1731 1618
rect 1737 1617 1738 1623
rect 84 1577 85 1583
rect 91 1582 1719 1583
rect 91 1578 111 1582
rect 115 1578 135 1582
rect 139 1578 167 1582
rect 171 1578 199 1582
rect 203 1578 231 1582
rect 235 1578 247 1582
rect 251 1578 287 1582
rect 291 1578 327 1582
rect 331 1578 343 1582
rect 347 1578 399 1582
rect 403 1578 439 1582
rect 443 1578 455 1582
rect 459 1578 511 1582
rect 515 1578 567 1582
rect 571 1578 575 1582
rect 579 1578 655 1582
rect 659 1578 711 1582
rect 715 1578 751 1582
rect 755 1578 855 1582
rect 859 1578 959 1582
rect 963 1578 999 1582
rect 1003 1578 1063 1582
rect 1067 1578 1127 1582
rect 1131 1578 1159 1582
rect 1163 1578 1247 1582
rect 1251 1578 1327 1582
rect 1331 1578 1359 1582
rect 1363 1578 1399 1582
rect 1403 1578 1463 1582
rect 1467 1578 1471 1582
rect 1475 1578 1535 1582
rect 1539 1578 1567 1582
rect 1571 1578 1607 1582
rect 1611 1578 1655 1582
rect 1659 1578 1695 1582
rect 1699 1578 1719 1582
rect 91 1577 1719 1578
rect 1725 1577 1726 1583
rect 96 1537 97 1543
rect 103 1542 1731 1543
rect 103 1538 111 1542
rect 115 1538 135 1542
rect 139 1538 167 1542
rect 171 1538 175 1542
rect 179 1538 223 1542
rect 227 1538 231 1542
rect 235 1538 279 1542
rect 283 1538 287 1542
rect 291 1538 335 1542
rect 339 1538 343 1542
rect 347 1538 399 1542
rect 403 1538 455 1542
rect 459 1538 463 1542
rect 467 1538 511 1542
rect 515 1538 535 1542
rect 539 1538 575 1542
rect 579 1538 607 1542
rect 611 1538 655 1542
rect 659 1538 687 1542
rect 691 1538 751 1542
rect 755 1538 775 1542
rect 779 1538 855 1542
rect 859 1538 871 1542
rect 875 1538 959 1542
rect 963 1538 975 1542
rect 979 1538 1063 1542
rect 1067 1538 1079 1542
rect 1083 1538 1159 1542
rect 1163 1538 1175 1542
rect 1179 1538 1247 1542
rect 1251 1538 1271 1542
rect 1275 1538 1327 1542
rect 1331 1538 1359 1542
rect 1363 1538 1399 1542
rect 1403 1538 1439 1542
rect 1443 1538 1471 1542
rect 1475 1538 1519 1542
rect 1523 1538 1535 1542
rect 1539 1538 1599 1542
rect 1603 1538 1607 1542
rect 1611 1538 1655 1542
rect 1659 1538 1695 1542
rect 1699 1538 1731 1542
rect 103 1537 1731 1538
rect 1737 1537 1738 1543
rect 84 1493 85 1499
rect 91 1498 1719 1499
rect 91 1494 111 1498
rect 115 1494 135 1498
rect 139 1494 175 1498
rect 179 1494 207 1498
rect 211 1494 223 1498
rect 227 1494 239 1498
rect 243 1494 271 1498
rect 275 1494 279 1498
rect 283 1494 303 1498
rect 307 1494 335 1498
rect 339 1494 367 1498
rect 371 1494 399 1498
rect 403 1494 431 1498
rect 435 1494 463 1498
rect 467 1494 495 1498
rect 499 1494 527 1498
rect 531 1494 535 1498
rect 539 1494 559 1498
rect 563 1494 591 1498
rect 595 1494 607 1498
rect 611 1494 623 1498
rect 627 1494 663 1498
rect 667 1494 687 1498
rect 691 1494 703 1498
rect 707 1494 743 1498
rect 747 1494 775 1498
rect 779 1494 807 1498
rect 811 1494 871 1498
rect 875 1494 895 1498
rect 899 1494 935 1498
rect 939 1494 975 1498
rect 979 1494 1023 1498
rect 1027 1494 1079 1498
rect 1083 1494 1111 1498
rect 1115 1494 1167 1498
rect 1171 1494 1175 1498
rect 1179 1494 1199 1498
rect 1203 1494 1239 1498
rect 1243 1494 1271 1498
rect 1275 1494 1279 1498
rect 1283 1494 1319 1498
rect 1323 1494 1359 1498
rect 1363 1494 1399 1498
rect 1403 1494 1439 1498
rect 1443 1494 1479 1498
rect 1483 1494 1519 1498
rect 1523 1494 1559 1498
rect 1563 1494 1591 1498
rect 1595 1494 1599 1498
rect 1603 1494 1623 1498
rect 1627 1494 1655 1498
rect 1659 1494 1695 1498
rect 1699 1494 1719 1498
rect 91 1493 1719 1494
rect 1725 1493 1726 1499
rect 96 1425 97 1431
rect 103 1430 1731 1431
rect 103 1426 111 1430
rect 115 1426 135 1430
rect 139 1426 167 1430
rect 171 1426 175 1430
rect 179 1426 199 1430
rect 203 1426 207 1430
rect 211 1426 231 1430
rect 235 1426 239 1430
rect 243 1426 263 1430
rect 267 1426 271 1430
rect 275 1426 295 1430
rect 299 1426 303 1430
rect 307 1426 327 1430
rect 331 1426 335 1430
rect 339 1426 359 1430
rect 363 1426 367 1430
rect 371 1426 391 1430
rect 395 1426 399 1430
rect 403 1426 423 1430
rect 427 1426 431 1430
rect 435 1426 455 1430
rect 459 1426 463 1430
rect 467 1426 487 1430
rect 491 1426 495 1430
rect 499 1426 519 1430
rect 523 1426 527 1430
rect 531 1426 551 1430
rect 555 1426 559 1430
rect 563 1426 583 1430
rect 587 1426 591 1430
rect 595 1426 615 1430
rect 619 1426 623 1430
rect 627 1426 647 1430
rect 651 1426 663 1430
rect 667 1426 679 1430
rect 683 1426 703 1430
rect 707 1426 719 1430
rect 723 1426 743 1430
rect 747 1426 767 1430
rect 771 1426 775 1430
rect 779 1426 807 1430
rect 811 1426 839 1430
rect 843 1426 895 1430
rect 899 1426 935 1430
rect 939 1426 975 1430
rect 979 1426 1023 1430
rect 1027 1426 1039 1430
rect 1043 1426 1063 1430
rect 1067 1426 1079 1430
rect 1083 1426 1111 1430
rect 1115 1426 1127 1430
rect 1131 1426 1151 1430
rect 1155 1426 1167 1430
rect 1171 1426 1199 1430
rect 1203 1426 1239 1430
rect 1243 1426 1263 1430
rect 1267 1426 1279 1430
rect 1283 1426 1319 1430
rect 1323 1426 1359 1430
rect 1363 1426 1399 1430
rect 1403 1426 1415 1430
rect 1419 1426 1439 1430
rect 1443 1426 1479 1430
rect 1483 1426 1519 1430
rect 1523 1426 1535 1430
rect 1539 1426 1559 1430
rect 1563 1426 1583 1430
rect 1587 1426 1591 1430
rect 1595 1426 1623 1430
rect 1627 1426 1655 1430
rect 1659 1426 1695 1430
rect 1699 1426 1731 1430
rect 103 1425 1731 1426
rect 1737 1425 1738 1431
rect 910 1420 916 1421
rect 990 1420 996 1421
rect 910 1416 911 1420
rect 915 1416 991 1420
rect 995 1416 996 1420
rect 910 1415 916 1416
rect 990 1415 996 1416
rect 84 1345 85 1351
rect 91 1350 1719 1351
rect 91 1346 111 1350
rect 115 1346 135 1350
rect 139 1346 167 1350
rect 171 1346 199 1350
rect 203 1346 231 1350
rect 235 1346 263 1350
rect 267 1346 295 1350
rect 299 1346 327 1350
rect 331 1346 359 1350
rect 363 1346 391 1350
rect 395 1346 423 1350
rect 427 1346 455 1350
rect 459 1346 487 1350
rect 491 1346 519 1350
rect 523 1346 551 1350
rect 555 1346 583 1350
rect 587 1346 615 1350
rect 619 1346 647 1350
rect 651 1346 679 1350
rect 683 1346 711 1350
rect 715 1346 735 1350
rect 739 1346 743 1350
rect 747 1346 767 1350
rect 771 1346 807 1350
rect 811 1346 823 1350
rect 827 1346 839 1350
rect 843 1346 887 1350
rect 891 1346 903 1350
rect 907 1346 975 1350
rect 979 1346 983 1350
rect 987 1346 1023 1350
rect 1027 1346 1063 1350
rect 1067 1346 1111 1350
rect 1115 1346 1151 1350
rect 1155 1346 1159 1350
rect 1163 1346 1199 1350
rect 1203 1346 1215 1350
rect 1219 1346 1247 1350
rect 1251 1346 1303 1350
rect 1307 1346 1319 1350
rect 1323 1346 1391 1350
rect 1395 1346 1415 1350
rect 1419 1346 1423 1350
rect 1427 1346 1455 1350
rect 1459 1346 1463 1350
rect 1467 1346 1495 1350
rect 1499 1346 1527 1350
rect 1531 1346 1535 1350
rect 1539 1346 1559 1350
rect 1563 1346 1583 1350
rect 1587 1346 1591 1350
rect 1595 1346 1623 1350
rect 1627 1346 1655 1350
rect 1659 1346 1695 1350
rect 1699 1346 1719 1350
rect 91 1345 1719 1346
rect 1725 1345 1726 1351
rect 1150 1271 1151 1277
rect 1157 1276 1160 1277
rect 1159 1272 1160 1276
rect 1157 1271 1160 1272
rect 1514 1276 1520 1277
rect 1574 1276 1575 1277
rect 1514 1272 1515 1276
rect 1519 1272 1575 1276
rect 1514 1271 1520 1272
rect 1574 1271 1575 1272
rect 1581 1271 1582 1277
rect 96 1257 97 1263
rect 103 1262 1731 1263
rect 103 1258 111 1262
rect 115 1258 135 1262
rect 139 1258 167 1262
rect 171 1258 199 1262
rect 203 1258 231 1262
rect 235 1258 263 1262
rect 267 1258 295 1262
rect 299 1258 327 1262
rect 331 1258 359 1262
rect 363 1258 391 1262
rect 395 1258 423 1262
rect 427 1258 455 1262
rect 459 1258 487 1262
rect 491 1258 519 1262
rect 523 1258 551 1262
rect 555 1258 583 1262
rect 587 1258 615 1262
rect 619 1258 647 1262
rect 651 1258 679 1262
rect 683 1258 711 1262
rect 715 1258 743 1262
rect 747 1258 751 1262
rect 755 1258 775 1262
rect 779 1258 811 1262
rect 815 1258 831 1262
rect 835 1258 911 1262
rect 915 1258 959 1262
rect 963 1258 983 1262
rect 987 1258 1015 1262
rect 1019 1258 1023 1262
rect 1027 1258 1063 1262
rect 1067 1258 1087 1262
rect 1091 1258 1127 1262
rect 1131 1258 1159 1262
rect 1163 1258 1175 1262
rect 1179 1258 1215 1262
rect 1219 1258 1255 1262
rect 1259 1258 1295 1262
rect 1299 1258 1303 1262
rect 1307 1258 1343 1262
rect 1347 1258 1375 1262
rect 1379 1258 1391 1262
rect 1395 1258 1407 1262
rect 1411 1258 1423 1262
rect 1427 1258 1439 1262
rect 1443 1258 1455 1262
rect 1459 1258 1479 1262
rect 1483 1258 1495 1262
rect 1499 1258 1519 1262
rect 1523 1258 1527 1262
rect 1531 1258 1559 1262
rect 1563 1258 1591 1262
rect 1595 1258 1623 1262
rect 1627 1258 1655 1262
rect 1659 1258 1695 1262
rect 1699 1258 1731 1262
rect 103 1257 1731 1258
rect 1737 1257 1738 1263
rect 1198 1207 1199 1213
rect 1205 1207 1206 1213
rect 84 1145 85 1151
rect 91 1150 1719 1151
rect 91 1146 111 1150
rect 115 1146 135 1150
rect 139 1146 167 1150
rect 171 1146 199 1150
rect 203 1146 231 1150
rect 235 1146 263 1150
rect 267 1146 295 1150
rect 299 1146 327 1150
rect 331 1146 359 1150
rect 363 1146 391 1150
rect 395 1146 423 1150
rect 427 1146 455 1150
rect 459 1146 487 1150
rect 491 1146 519 1150
rect 523 1146 551 1150
rect 555 1146 583 1150
rect 587 1146 615 1150
rect 619 1146 647 1150
rect 651 1146 679 1150
rect 683 1146 687 1150
rect 691 1146 711 1150
rect 715 1146 743 1150
rect 747 1146 775 1150
rect 779 1146 799 1150
rect 803 1146 839 1150
rect 843 1146 847 1150
rect 851 1146 935 1150
rect 939 1146 967 1150
rect 971 1146 975 1150
rect 979 1146 999 1150
rect 1003 1146 1007 1150
rect 1011 1146 1031 1150
rect 1035 1146 1063 1150
rect 1067 1146 1087 1150
rect 1091 1146 1095 1150
rect 1099 1146 1127 1150
rect 1131 1146 1135 1150
rect 1139 1146 1159 1150
rect 1163 1146 1167 1150
rect 1171 1146 1199 1150
rect 1203 1146 1247 1150
rect 1251 1146 1255 1150
rect 1259 1146 1287 1150
rect 1291 1146 1311 1150
rect 1315 1146 1335 1150
rect 1339 1146 1343 1150
rect 1347 1146 1375 1150
rect 1379 1146 1407 1150
rect 1411 1146 1423 1150
rect 1427 1146 1439 1150
rect 1443 1146 1455 1150
rect 1459 1146 1479 1150
rect 1483 1146 1487 1150
rect 1491 1146 1519 1150
rect 1523 1146 1559 1150
rect 1563 1146 1591 1150
rect 1595 1146 1623 1150
rect 1627 1146 1655 1150
rect 1659 1146 1695 1150
rect 1699 1146 1719 1150
rect 91 1145 1719 1146
rect 1725 1145 1726 1151
rect 382 1092 388 1093
rect 670 1092 676 1093
rect 1074 1092 1080 1093
rect 382 1088 383 1092
rect 387 1088 671 1092
rect 675 1088 1075 1092
rect 1079 1088 1080 1092
rect 382 1087 388 1088
rect 670 1087 676 1088
rect 1074 1087 1080 1088
rect 186 1060 192 1061
rect 814 1060 820 1061
rect 186 1056 187 1060
rect 191 1056 815 1060
rect 819 1056 820 1060
rect 186 1055 192 1056
rect 814 1055 820 1056
rect 178 1044 184 1045
rect 398 1044 404 1045
rect 178 1040 179 1044
rect 183 1040 399 1044
rect 403 1040 404 1044
rect 178 1039 184 1040
rect 398 1039 404 1040
rect 96 1029 97 1035
rect 103 1034 1731 1035
rect 103 1030 111 1034
rect 115 1030 135 1034
rect 139 1030 167 1034
rect 171 1030 199 1034
rect 203 1030 231 1034
rect 235 1030 263 1034
rect 267 1030 295 1034
rect 299 1030 327 1034
rect 331 1030 359 1034
rect 363 1030 391 1034
rect 395 1030 407 1034
rect 411 1030 423 1034
rect 427 1030 455 1034
rect 459 1030 487 1034
rect 491 1030 503 1034
rect 507 1030 519 1034
rect 523 1030 551 1034
rect 555 1030 583 1034
rect 587 1030 591 1034
rect 595 1030 659 1034
rect 663 1030 711 1034
rect 715 1030 799 1034
rect 803 1030 823 1034
rect 827 1030 847 1034
rect 851 1030 919 1034
rect 923 1030 935 1034
rect 939 1030 967 1034
rect 971 1030 975 1034
rect 979 1030 999 1034
rect 1003 1030 1031 1034
rect 1035 1030 1063 1034
rect 1067 1030 1095 1034
rect 1099 1030 1119 1034
rect 1123 1030 1135 1034
rect 1139 1030 1167 1034
rect 1171 1030 1175 1034
rect 1179 1030 1199 1034
rect 1203 1030 1247 1034
rect 1251 1030 1287 1034
rect 1291 1030 1295 1034
rect 1299 1030 1327 1034
rect 1331 1030 1335 1034
rect 1339 1030 1367 1034
rect 1371 1030 1407 1034
rect 1411 1030 1423 1034
rect 1427 1030 1439 1034
rect 1443 1030 1455 1034
rect 1459 1030 1479 1034
rect 1483 1030 1487 1034
rect 1491 1030 1519 1034
rect 1523 1030 1559 1034
rect 1563 1030 1591 1034
rect 1595 1030 1623 1034
rect 1627 1030 1655 1034
rect 1659 1030 1695 1034
rect 1699 1030 1731 1034
rect 103 1029 1731 1030
rect 1737 1029 1738 1035
rect 84 949 85 955
rect 91 954 1719 955
rect 91 950 111 954
rect 115 950 135 954
rect 139 950 167 954
rect 171 950 199 954
rect 203 950 231 954
rect 235 950 263 954
rect 267 950 279 954
rect 283 950 319 954
rect 323 950 343 954
rect 347 950 399 954
rect 403 950 463 954
rect 467 950 503 954
rect 507 950 583 954
rect 587 950 591 954
rect 595 950 679 954
rect 683 950 711 954
rect 715 950 727 954
rect 731 950 815 954
rect 819 950 863 954
rect 867 950 919 954
rect 923 950 951 954
rect 955 950 967 954
rect 971 950 983 954
rect 987 950 1039 954
rect 1043 950 1063 954
rect 1067 950 1071 954
rect 1075 950 1111 954
rect 1115 950 1135 954
rect 1139 950 1143 954
rect 1147 950 1167 954
rect 1171 950 1199 954
rect 1203 950 1239 954
rect 1243 950 1263 954
rect 1267 950 1271 954
rect 1275 950 1295 954
rect 1299 950 1327 954
rect 1331 950 1367 954
rect 1371 950 1391 954
rect 1395 950 1407 954
rect 1411 950 1423 954
rect 1427 950 1439 954
rect 1443 950 1455 954
rect 1459 950 1479 954
rect 1483 950 1519 954
rect 1523 950 1559 954
rect 1563 950 1591 954
rect 1595 950 1623 954
rect 1627 950 1655 954
rect 1659 950 1695 954
rect 1699 950 1719 954
rect 91 949 1719 950
rect 1725 949 1726 955
rect 1574 879 1575 885
rect 1581 884 1582 885
rect 1662 884 1668 885
rect 1581 880 1663 884
rect 1667 880 1668 884
rect 1581 879 1582 880
rect 1662 879 1668 880
rect 96 833 97 839
rect 103 838 1731 839
rect 103 834 111 838
rect 115 834 135 838
rect 139 834 167 838
rect 171 834 207 838
rect 211 834 231 838
rect 235 834 279 838
rect 283 834 327 838
rect 331 834 399 838
rect 403 834 407 838
rect 411 834 435 838
rect 439 834 559 838
rect 563 834 591 838
rect 595 834 663 838
rect 667 834 679 838
rect 683 834 727 838
rect 731 834 815 838
rect 819 834 863 838
rect 867 834 951 838
rect 955 834 999 838
rect 1003 834 1031 838
rect 1035 834 1039 838
rect 1043 834 1071 838
rect 1075 834 1103 838
rect 1107 834 1111 838
rect 1115 834 1143 838
rect 1147 834 1167 838
rect 1171 834 1239 838
rect 1243 834 1247 838
rect 1251 834 1271 838
rect 1275 834 1295 838
rect 1299 834 1327 838
rect 1331 834 1375 838
rect 1379 834 1423 838
rect 1427 834 1471 838
rect 1475 834 1519 838
rect 1523 834 1559 838
rect 1563 834 1591 838
rect 1595 834 1623 838
rect 1627 834 1655 838
rect 1659 834 1695 838
rect 1699 834 1731 838
rect 103 833 1731 834
rect 1737 833 1738 839
rect 1054 812 1060 813
rect 1150 812 1151 813
rect 1054 808 1055 812
rect 1059 808 1151 812
rect 1054 807 1060 808
rect 1150 807 1151 808
rect 1157 807 1158 813
rect 1198 791 1199 797
rect 1205 796 1206 797
rect 1270 796 1276 797
rect 1205 792 1271 796
rect 1275 792 1276 796
rect 1205 791 1206 792
rect 1270 791 1276 792
rect 84 749 85 755
rect 91 754 1719 755
rect 91 750 111 754
rect 115 750 135 754
rect 139 750 215 754
rect 219 750 231 754
rect 235 750 287 754
rect 291 750 391 754
rect 395 750 407 754
rect 411 750 471 754
rect 475 750 559 754
rect 563 750 615 754
rect 619 750 655 754
rect 659 750 719 754
rect 723 750 767 754
rect 771 750 815 754
rect 819 750 863 754
rect 867 750 911 754
rect 915 750 951 754
rect 955 750 999 754
rect 1003 750 1015 754
rect 1019 750 1087 754
rect 1091 750 1103 754
rect 1107 750 1167 754
rect 1171 750 1183 754
rect 1187 750 1207 754
rect 1211 750 1231 754
rect 1235 750 1247 754
rect 1251 750 1279 754
rect 1283 750 1295 754
rect 1299 750 1311 754
rect 1315 750 1327 754
rect 1331 750 1343 754
rect 1347 750 1375 754
rect 1379 750 1407 754
rect 1411 750 1423 754
rect 1427 750 1439 754
rect 1443 750 1471 754
rect 1475 750 1479 754
rect 1483 750 1519 754
rect 1523 750 1559 754
rect 1563 750 1591 754
rect 1595 750 1623 754
rect 1627 750 1655 754
rect 1659 750 1695 754
rect 1699 750 1719 754
rect 91 749 1719 750
rect 1725 749 1726 755
rect 622 684 628 685
rect 982 684 988 685
rect 622 680 623 684
rect 627 680 983 684
rect 987 680 988 684
rect 622 679 628 680
rect 982 679 988 680
rect 96 637 97 643
rect 103 642 1731 643
rect 103 638 111 642
rect 115 638 135 642
rect 139 638 143 642
rect 147 638 167 642
rect 171 638 207 642
rect 211 638 215 642
rect 219 638 287 642
rect 291 638 391 642
rect 395 638 407 642
rect 411 638 443 642
rect 447 638 535 642
rect 539 638 615 642
rect 619 638 671 642
rect 675 638 719 642
rect 723 638 767 642
rect 771 638 775 642
rect 779 638 863 642
rect 867 638 903 642
rect 907 638 911 642
rect 915 638 999 642
rect 1003 638 1007 642
rect 1011 638 1095 642
rect 1099 638 1119 642
rect 1123 638 1167 642
rect 1171 638 1207 642
rect 1211 638 1215 642
rect 1219 638 1247 642
rect 1251 638 1279 642
rect 1283 638 1311 642
rect 1315 638 1335 642
rect 1339 638 1343 642
rect 1347 638 1375 642
rect 1379 638 1407 642
rect 1411 638 1415 642
rect 1419 638 1439 642
rect 1443 638 1479 642
rect 1483 638 1519 642
rect 1523 638 1543 642
rect 1547 638 1559 642
rect 1563 638 1591 642
rect 1595 638 1607 642
rect 1611 638 1623 642
rect 1627 638 1655 642
rect 1659 638 1695 642
rect 1699 638 1731 642
rect 103 637 1731 638
rect 1737 637 1738 643
rect 84 557 85 563
rect 91 562 1719 563
rect 91 558 111 562
rect 115 558 135 562
rect 139 558 167 562
rect 171 558 207 562
rect 211 558 247 562
rect 251 558 279 562
rect 283 558 303 562
rect 307 558 391 562
rect 395 558 399 562
rect 403 558 471 562
rect 475 558 535 562
rect 539 558 647 562
rect 651 558 671 562
rect 675 558 727 562
rect 731 558 767 562
rect 771 558 775 562
rect 779 558 871 562
rect 875 558 903 562
rect 907 558 927 562
rect 931 558 991 562
rect 995 558 1031 562
rect 1035 558 1095 562
rect 1099 558 1119 562
rect 1123 558 1199 562
rect 1203 558 1207 562
rect 1211 558 1287 562
rect 1291 558 1335 562
rect 1339 558 1415 562
rect 1419 558 1423 562
rect 1427 558 1479 562
rect 1483 558 1527 562
rect 1531 558 1543 562
rect 1547 558 1575 562
rect 1579 558 1607 562
rect 1611 558 1623 562
rect 1627 558 1655 562
rect 1659 558 1695 562
rect 1699 558 1719 562
rect 91 557 1719 558
rect 1725 557 1726 563
rect 96 437 97 443
rect 103 442 1731 443
rect 103 438 111 442
rect 115 438 135 442
rect 139 438 167 442
rect 171 438 175 442
rect 179 438 199 442
rect 203 438 231 442
rect 235 438 247 442
rect 251 438 263 442
rect 267 438 303 442
rect 307 438 375 442
rect 379 438 399 442
rect 403 438 415 442
rect 419 438 447 442
rect 451 438 471 442
rect 475 438 487 442
rect 491 438 507 442
rect 511 438 543 442
rect 547 438 615 442
rect 619 438 655 442
rect 659 438 671 442
rect 675 438 727 442
rect 731 438 755 442
rect 759 438 783 442
rect 787 438 871 442
rect 875 438 903 442
rect 907 438 935 442
rect 939 438 951 442
rect 955 438 1031 442
rect 1035 438 1075 442
rect 1079 438 1103 442
rect 1107 438 1199 442
rect 1203 438 1231 442
rect 1235 438 1259 442
rect 1263 438 1319 442
rect 1323 438 1359 442
rect 1363 438 1423 442
rect 1427 438 1439 442
rect 1443 438 1479 442
rect 1483 438 1519 442
rect 1523 438 1527 442
rect 1531 438 1559 442
rect 1563 438 1575 442
rect 1579 438 1591 442
rect 1595 438 1623 442
rect 1627 438 1655 442
rect 1659 438 1695 442
rect 1699 438 1731 442
rect 103 437 1731 438
rect 1737 437 1738 443
rect 982 364 988 365
rect 1722 364 1728 365
rect 982 360 983 364
rect 987 360 1723 364
rect 1727 360 1728 364
rect 982 359 988 360
rect 1722 359 1728 360
rect 84 317 85 323
rect 91 322 1719 323
rect 91 318 111 322
rect 115 318 135 322
rect 139 318 167 322
rect 171 318 199 322
rect 203 318 231 322
rect 235 318 263 322
rect 267 318 295 322
rect 299 318 327 322
rect 331 318 359 322
rect 363 318 375 322
rect 379 318 391 322
rect 395 318 415 322
rect 419 318 423 322
rect 427 318 447 322
rect 451 318 455 322
rect 459 318 487 322
rect 491 318 503 322
rect 507 318 519 322
rect 523 318 535 322
rect 539 318 551 322
rect 555 318 599 322
rect 603 318 615 322
rect 619 318 671 322
rect 675 318 703 322
rect 707 318 783 322
rect 787 318 807 322
rect 811 318 903 322
rect 907 318 911 322
rect 915 318 943 322
rect 947 318 999 322
rect 1003 318 1031 322
rect 1035 318 1047 322
rect 1051 318 1063 322
rect 1067 318 1103 322
rect 1107 318 1111 322
rect 1115 318 1199 322
rect 1203 318 1231 322
rect 1235 318 1287 322
rect 1291 318 1319 322
rect 1323 318 1351 322
rect 1355 318 1383 322
rect 1387 318 1415 322
rect 1419 318 1439 322
rect 1443 318 1447 322
rect 1451 318 1479 322
rect 1483 318 1519 322
rect 1523 318 1559 322
rect 1563 318 1591 322
rect 1595 318 1623 322
rect 1627 318 1655 322
rect 1659 318 1695 322
rect 1699 318 1719 322
rect 91 317 1719 318
rect 1725 317 1726 323
rect 82 308 88 309
rect 526 308 532 309
rect 82 304 83 308
rect 87 304 527 308
rect 531 304 532 308
rect 82 303 88 304
rect 526 303 532 304
rect 606 260 612 261
rect 926 260 932 261
rect 606 256 607 260
rect 611 256 927 260
rect 931 256 932 260
rect 606 255 612 256
rect 926 255 932 256
rect 96 245 97 251
rect 103 250 1731 251
rect 103 246 111 250
rect 115 246 135 250
rect 139 246 167 250
rect 171 246 183 250
rect 187 246 199 250
rect 203 246 215 250
rect 219 246 231 250
rect 235 246 247 250
rect 251 246 263 250
rect 267 246 279 250
rect 283 246 295 250
rect 299 246 311 250
rect 315 246 327 250
rect 331 246 343 250
rect 347 246 359 250
rect 363 246 375 250
rect 379 246 391 250
rect 395 246 407 250
rect 411 246 423 250
rect 427 246 439 250
rect 443 246 455 250
rect 459 246 471 250
rect 475 246 487 250
rect 491 246 503 250
rect 507 246 519 250
rect 523 246 535 250
rect 539 246 551 250
rect 555 246 567 250
rect 571 246 599 250
rect 603 246 639 250
rect 643 246 695 250
rect 699 246 703 250
rect 707 246 791 250
rect 795 246 807 250
rect 811 246 839 250
rect 843 246 911 250
rect 915 246 919 250
rect 923 246 967 250
rect 971 246 999 250
rect 1003 246 1031 250
rect 1035 246 1063 250
rect 1067 246 1103 250
rect 1107 246 1111 250
rect 1115 246 1143 250
rect 1147 246 1183 250
rect 1187 246 1207 250
rect 1211 246 1223 250
rect 1227 246 1263 250
rect 1267 246 1287 250
rect 1291 246 1303 250
rect 1307 246 1319 250
rect 1323 246 1343 250
rect 1347 246 1351 250
rect 1355 246 1375 250
rect 1379 246 1383 250
rect 1387 246 1407 250
rect 1411 246 1415 250
rect 1419 246 1439 250
rect 1443 246 1447 250
rect 1451 246 1479 250
rect 1483 246 1519 250
rect 1523 246 1559 250
rect 1563 246 1591 250
rect 1595 246 1623 250
rect 1627 246 1655 250
rect 1659 246 1695 250
rect 1699 246 1731 250
rect 103 245 1731 246
rect 1737 245 1738 251
rect 84 169 85 175
rect 91 174 1719 175
rect 91 170 111 174
rect 115 170 135 174
rect 139 170 167 174
rect 171 170 183 174
rect 187 170 215 174
rect 219 170 247 174
rect 251 170 263 174
rect 267 170 279 174
rect 283 170 311 174
rect 315 170 343 174
rect 347 170 367 174
rect 371 170 375 174
rect 379 170 407 174
rect 411 170 415 174
rect 419 170 439 174
rect 443 170 471 174
rect 475 170 503 174
rect 507 170 535 174
rect 539 170 567 174
rect 571 170 599 174
rect 603 170 607 174
rect 611 170 639 174
rect 643 170 687 174
rect 691 170 695 174
rect 699 170 775 174
rect 779 170 791 174
rect 795 170 831 174
rect 835 170 863 174
rect 867 170 919 174
rect 923 170 959 174
rect 963 170 967 174
rect 971 170 1055 174
rect 1059 170 1063 174
rect 1067 170 1103 174
rect 1107 170 1143 174
rect 1147 170 1151 174
rect 1155 170 1183 174
rect 1187 170 1223 174
rect 1227 170 1239 174
rect 1243 170 1263 174
rect 1267 170 1303 174
rect 1307 170 1327 174
rect 1331 170 1343 174
rect 1347 170 1375 174
rect 1379 170 1407 174
rect 1411 170 1415 174
rect 1419 170 1439 174
rect 1443 170 1479 174
rect 1483 170 1503 174
rect 1507 170 1519 174
rect 1523 170 1559 174
rect 1563 170 1591 174
rect 1595 170 1623 174
rect 1627 170 1655 174
rect 1659 170 1695 174
rect 1699 170 1719 174
rect 91 169 1719 170
rect 1725 169 1726 175
rect 96 117 97 123
rect 103 122 1731 123
rect 103 118 111 122
rect 115 118 135 122
rect 139 118 167 122
rect 171 118 199 122
rect 203 118 215 122
rect 219 118 231 122
rect 235 118 263 122
rect 267 118 295 122
rect 299 118 311 122
rect 315 118 327 122
rect 331 118 359 122
rect 363 118 367 122
rect 371 118 391 122
rect 395 118 415 122
rect 419 118 423 122
rect 427 118 455 122
rect 459 118 471 122
rect 475 118 487 122
rect 491 118 519 122
rect 523 118 535 122
rect 539 118 551 122
rect 555 118 607 122
rect 611 118 671 122
rect 675 118 687 122
rect 691 118 743 122
rect 747 118 775 122
rect 779 118 823 122
rect 827 118 863 122
rect 867 118 903 122
rect 907 118 959 122
rect 963 118 983 122
rect 987 118 1055 122
rect 1059 118 1119 122
rect 1123 118 1151 122
rect 1155 118 1175 122
rect 1179 118 1223 122
rect 1227 118 1239 122
rect 1243 118 1271 122
rect 1275 118 1311 122
rect 1315 118 1327 122
rect 1331 118 1343 122
rect 1347 118 1375 122
rect 1379 118 1407 122
rect 1411 118 1415 122
rect 1419 118 1439 122
rect 1443 118 1479 122
rect 1483 118 1503 122
rect 1507 118 1519 122
rect 1523 118 1559 122
rect 1563 118 1591 122
rect 1595 118 1623 122
rect 1627 118 1655 122
rect 1659 118 1695 122
rect 1699 118 1731 122
rect 103 117 1731 118
rect 1737 117 1738 123
rect 84 77 85 83
rect 91 82 1719 83
rect 91 78 111 82
rect 115 78 135 82
rect 139 78 167 82
rect 171 78 199 82
rect 203 78 231 82
rect 235 78 263 82
rect 267 78 295 82
rect 299 78 327 82
rect 331 78 359 82
rect 363 78 391 82
rect 395 78 423 82
rect 427 78 455 82
rect 459 78 487 82
rect 491 78 519 82
rect 523 78 551 82
rect 555 78 607 82
rect 611 78 671 82
rect 675 78 743 82
rect 747 78 823 82
rect 827 78 903 82
rect 907 78 983 82
rect 987 78 1055 82
rect 1059 78 1119 82
rect 1123 78 1175 82
rect 1179 78 1223 82
rect 1227 78 1271 82
rect 1275 78 1311 82
rect 1315 78 1343 82
rect 1347 78 1375 82
rect 1379 78 1407 82
rect 1411 78 1439 82
rect 1443 78 1479 82
rect 1483 78 1519 82
rect 1523 78 1559 82
rect 1563 78 1591 82
rect 1595 78 1623 82
rect 1627 78 1655 82
rect 1659 78 1695 82
rect 1699 78 1719 82
rect 91 77 1719 78
rect 1725 77 1726 83
<< m5c >>
rect 85 1757 91 1763
rect 1719 1757 1725 1763
rect 97 1713 103 1719
rect 1731 1713 1737 1719
rect 85 1665 91 1671
rect 1719 1665 1725 1671
rect 97 1617 103 1623
rect 1731 1617 1737 1623
rect 85 1577 91 1583
rect 1719 1577 1725 1583
rect 97 1537 103 1543
rect 1731 1537 1737 1543
rect 85 1493 91 1499
rect 1719 1493 1725 1499
rect 97 1425 103 1431
rect 1731 1425 1737 1431
rect 85 1345 91 1351
rect 1719 1345 1725 1351
rect 1151 1276 1157 1277
rect 1151 1272 1155 1276
rect 1155 1272 1157 1276
rect 1151 1271 1157 1272
rect 1575 1271 1581 1277
rect 97 1257 103 1263
rect 1731 1257 1737 1263
rect 1199 1212 1205 1213
rect 1199 1208 1203 1212
rect 1203 1208 1205 1212
rect 1199 1207 1205 1208
rect 85 1145 91 1151
rect 1719 1145 1725 1151
rect 97 1029 103 1035
rect 1731 1029 1737 1035
rect 85 949 91 955
rect 1719 949 1725 955
rect 1575 879 1581 885
rect 97 833 103 839
rect 1731 833 1737 839
rect 1151 807 1157 813
rect 1199 791 1205 797
rect 85 749 91 755
rect 1719 749 1725 755
rect 97 637 103 643
rect 1731 637 1737 643
rect 85 557 91 563
rect 1719 557 1725 563
rect 97 437 103 443
rect 1731 437 1737 443
rect 85 317 91 323
rect 1719 317 1725 323
rect 97 245 103 251
rect 1731 245 1737 251
rect 85 169 91 175
rect 1719 169 1725 175
rect 97 117 103 123
rect 1731 117 1737 123
rect 85 77 91 83
rect 1719 77 1725 83
<< m5 >>
rect 84 1763 92 1800
rect 84 1757 85 1763
rect 91 1757 92 1763
rect 84 1671 92 1757
rect 84 1665 85 1671
rect 91 1665 92 1671
rect 84 1583 92 1665
rect 84 1577 85 1583
rect 91 1577 92 1583
rect 84 1499 92 1577
rect 84 1493 85 1499
rect 91 1493 92 1499
rect 84 1351 92 1493
rect 84 1345 85 1351
rect 91 1345 92 1351
rect 84 1151 92 1345
rect 84 1145 85 1151
rect 91 1145 92 1151
rect 84 955 92 1145
rect 84 949 85 955
rect 91 949 92 955
rect 84 755 92 949
rect 84 749 85 755
rect 91 749 92 755
rect 84 563 92 749
rect 84 557 85 563
rect 91 557 92 563
rect 84 323 92 557
rect 84 317 85 323
rect 91 317 92 323
rect 84 175 92 317
rect 84 169 85 175
rect 91 169 92 175
rect 84 83 92 169
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 1719 104 1800
rect 96 1713 97 1719
rect 103 1713 104 1719
rect 96 1623 104 1713
rect 96 1617 97 1623
rect 103 1617 104 1623
rect 96 1543 104 1617
rect 96 1537 97 1543
rect 103 1537 104 1543
rect 96 1431 104 1537
rect 96 1425 97 1431
rect 103 1425 104 1431
rect 96 1263 104 1425
rect 1718 1763 1726 1800
rect 1718 1757 1719 1763
rect 1725 1757 1726 1763
rect 1718 1671 1726 1757
rect 1718 1665 1719 1671
rect 1725 1665 1726 1671
rect 1718 1583 1726 1665
rect 1718 1577 1719 1583
rect 1725 1577 1726 1583
rect 1718 1499 1726 1577
rect 1718 1493 1719 1499
rect 1725 1493 1726 1499
rect 1718 1351 1726 1493
rect 1718 1345 1719 1351
rect 1725 1345 1726 1351
rect 1150 1277 1158 1278
rect 1150 1271 1151 1277
rect 1157 1271 1158 1277
rect 1150 1270 1158 1271
rect 1574 1277 1582 1278
rect 1574 1271 1575 1277
rect 1581 1271 1582 1277
rect 1574 1270 1582 1271
rect 96 1257 97 1263
rect 103 1257 104 1263
rect 96 1035 104 1257
rect 96 1029 97 1035
rect 103 1029 104 1035
rect 96 839 104 1029
rect 96 833 97 839
rect 103 833 104 839
rect 96 643 104 833
rect 1152 814 1156 1270
rect 1198 1213 1206 1214
rect 1198 1207 1199 1213
rect 1205 1207 1206 1213
rect 1198 1206 1206 1207
rect 1150 813 1158 814
rect 1150 807 1151 813
rect 1157 807 1158 813
rect 1150 806 1158 807
rect 1200 798 1204 1206
rect 1576 886 1580 1270
rect 1718 1151 1726 1345
rect 1718 1145 1719 1151
rect 1725 1145 1726 1151
rect 1718 955 1726 1145
rect 1718 949 1719 955
rect 1725 949 1726 955
rect 1574 885 1582 886
rect 1574 879 1575 885
rect 1581 879 1582 885
rect 1574 878 1582 879
rect 1198 797 1206 798
rect 1198 791 1199 797
rect 1205 791 1206 797
rect 1198 790 1206 791
rect 96 637 97 643
rect 103 637 104 643
rect 96 443 104 637
rect 96 437 97 443
rect 103 437 104 443
rect 96 251 104 437
rect 96 245 97 251
rect 103 245 104 251
rect 96 123 104 245
rect 96 117 97 123
rect 103 117 104 123
rect 96 72 104 117
rect 1718 755 1726 949
rect 1718 749 1719 755
rect 1725 749 1726 755
rect 1718 563 1726 749
rect 1718 557 1719 563
rect 1725 557 1726 563
rect 1718 323 1726 557
rect 1718 317 1719 323
rect 1725 317 1726 323
rect 1718 175 1726 317
rect 1718 169 1719 175
rect 1725 169 1726 175
rect 1718 83 1726 169
rect 1718 77 1719 83
rect 1725 77 1726 83
rect 1718 72 1726 77
rect 1730 1719 1738 1800
rect 1730 1713 1731 1719
rect 1737 1713 1738 1719
rect 1730 1623 1738 1713
rect 1730 1617 1731 1623
rect 1737 1617 1738 1623
rect 1730 1543 1738 1617
rect 1730 1537 1731 1543
rect 1737 1537 1738 1543
rect 1730 1431 1738 1537
rect 1730 1425 1731 1431
rect 1737 1425 1738 1431
rect 1730 1263 1738 1425
rect 1730 1257 1731 1263
rect 1737 1257 1738 1263
rect 1730 1035 1738 1257
rect 1730 1029 1731 1035
rect 1737 1029 1738 1035
rect 1730 839 1738 1029
rect 1730 833 1731 839
rect 1737 833 1738 839
rect 1730 643 1738 833
rect 1730 637 1731 643
rect 1737 637 1738 643
rect 1730 443 1738 637
rect 1730 437 1731 443
rect 1737 437 1738 443
rect 1730 251 1738 437
rect 1730 245 1731 251
rect 1737 245 1738 251
rect 1730 123 1738 245
rect 1730 117 1731 123
rect 1737 117 1738 123
rect 1730 72 1738 117
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__43
timestamp 1731220320
transform 1 0 1688 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220320
transform 1 0 104 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220320
transform 1 0 1688 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220320
transform 1 0 104 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220320
transform 1 0 1688 0 -1 1664
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220320
transform 1 0 104 0 -1 1664
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220320
transform 1 0 1688 0 1 1584
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220320
transform 1 0 104 0 1 1584
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220320
transform 1 0 1688 0 -1 1576
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220320
transform 1 0 104 0 -1 1576
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220320
transform 1 0 1688 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220320
transform 1 0 104 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220320
transform 1 0 1688 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220320
transform 1 0 104 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220320
transform 1 0 1688 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220320
transform 1 0 104 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220320
transform 1 0 1688 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220320
transform 1 0 104 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220320
transform 1 0 1688 0 1 1172
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220320
transform 1 0 104 0 1 1172
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220320
transform 1 0 1688 0 -1 1124
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220320
transform 1 0 104 0 -1 1124
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220320
transform 1 0 1688 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220320
transform 1 0 104 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220320
transform 1 0 1688 0 -1 924
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220320
transform 1 0 104 0 -1 924
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220320
transform 1 0 1688 0 1 780
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220320
transform 1 0 104 0 1 780
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220320
transform 1 0 1688 0 -1 728
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220320
transform 1 0 104 0 -1 728
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220320
transform 1 0 1688 0 1 580
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220320
transform 1 0 104 0 1 580
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220320
transform 1 0 1688 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220320
transform 1 0 104 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220320
transform 1 0 1688 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220320
transform 1 0 104 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220320
transform 1 0 1688 0 -1 304
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220320
transform 1 0 104 0 -1 304
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220320
transform 1 0 1688 0 1 192
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220320
transform 1 0 104 0 1 192
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220320
transform 1 0 1688 0 -1 168
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220320
transform 1 0 104 0 -1 168
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220320
transform 1 0 1688 0 1 84
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220320
transform 1 0 104 0 1 84
box 7 3 12 24
use _0_0std_0_0cells_0_0INVX1  splt_ar0_ai
timestamp 1731220320
transform 1 0 1472 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  splt_ar0_an
timestamp 1731220320
transform 1 0 1464 0 1 776
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_55_6
timestamp 1731220320
transform 1 0 1056 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_54_6
timestamp 1731220320
transform 1 0 1024 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_53_6
timestamp 1731220320
transform 1 0 960 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_52_6
timestamp 1731220320
transform 1 0 928 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_51_6
timestamp 1731220320
transform 1 0 1120 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_50_6
timestamp 1731220320
transform 1 0 1152 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ac__latch__inv
timestamp 1731220320
transform 1 0 1280 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0OR2X1  splt_ar2_an
timestamp 1731220320
transform 1 0 1448 0 -1 928
box 4 4 48 48
use _0_0std_0_0cells_0_0INVX1  splt_ar1_ai
timestamp 1731220320
transform 1 0 1240 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  splt_ar1_an
timestamp 1731220320
transform 1 0 1200 0 -1 732
box 4 6 36 48
use _0_0cell_0_0ginvx0  splt_ac_acx1
timestamp 1731220320
transform 1 0 1288 0 1 776
box 8 6 28 32
use _0_0cell_0_0gcelem3x0  splt_ac_acx0
timestamp 1731220320
transform 1 0 1320 0 1 752
box 8 5 92 72
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_544_6
timestamp 1731220320
transform 1 0 1024 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_543_6
timestamp 1731220320
transform 1 0 992 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_542_6
timestamp 1731220320
transform 1 0 1056 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_541_6
timestamp 1731220320
transform 1 0 1048 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_540_6
timestamp 1731220320
transform 1 0 976 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_539_6
timestamp 1731220320
transform 1 0 952 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_538_6
timestamp 1731220320
transform 1 0 1144 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_537_6
timestamp 1731220320
transform 1 0 1136 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_536_6
timestamp 1731220320
transform 1 0 1096 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_535_6
timestamp 1731220320
transform 1 0 1176 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_534_6
timestamp 1731220320
transform 1 0 1216 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_533_6
timestamp 1731220320
transform 1 0 1256 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_532_6
timestamp 1731220320
transform 1 0 1320 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_531_6
timestamp 1731220320
transform 1 0 1232 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_530_6
timestamp 1731220320
transform 1 0 1168 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_529_6
timestamp 1731220320
transform 1 0 1112 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_528_6
timestamp 1731220320
transform 1 0 1048 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_527_6
timestamp 1731220320
transform 1 0 1216 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_526_6
timestamp 1731220320
transform 1 0 1264 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_525_6
timestamp 1731220320
transform 1 0 1304 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_524_6
timestamp 1731220320
transform 1 0 1336 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_523_6
timestamp 1731220320
transform 1 0 1368 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_522_6
timestamp 1731220320
transform 1 0 1400 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_521_6
timestamp 1731220320
transform 1 0 1432 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_520_6
timestamp 1731220320
transform 1 0 1472 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_519_6
timestamp 1731220320
transform 1 0 1512 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_518_6
timestamp 1731220320
transform 1 0 1496 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_517_6
timestamp 1731220320
transform 1 0 1408 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_516_6
timestamp 1731220320
transform 1 0 1584 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_515_6
timestamp 1731220320
transform 1 0 1552 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_514_6
timestamp 1731220320
transform 1 0 1512 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_513_6
timestamp 1731220320
transform 1 0 1472 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_512_6
timestamp 1731220320
transform 1 0 1432 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_511_6
timestamp 1731220320
transform 1 0 1400 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_510_6
timestamp 1731220320
transform 1 0 1368 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_59_6
timestamp 1731220320
transform 1 0 1336 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_58_6
timestamp 1731220320
transform 1 0 1296 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_57_6
timestamp 1731220320
transform 1 0 1512 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_56_6
timestamp 1731220320
transform 1 0 1472 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_55_6
timestamp 1731220320
transform 1 0 1440 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_54_6
timestamp 1731220320
transform 1 0 1408 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_53_6
timestamp 1731220320
transform 1 0 1376 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_52_6
timestamp 1731220320
transform 1 0 1344 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_51_6
timestamp 1731220320
transform 1 0 1312 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_50_6
timestamp 1731220320
transform 1 0 1312 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  splt_ap_aand
timestamp 1731220320
transform 1 0 1016 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0OR2X1  splt_ar3_an
timestamp 1731220320
transform 1 0 1224 0 1 776
box 4 4 48 48
use _0_0std_0_0cells_0_0AND2X1  splt_ar1__r
timestamp 1731220320
transform 1 0 1232 0 1 956
box 8 4 52 52
use _0_0std_0_0cells_0_0LATCHINV  splt_ac__latch_al
timestamp 1731220320
transform 1 0 1160 0 -1 1144
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  splt_ac__latch_anx
timestamp 1731220320
transform 1 0 1240 0 -1 1132
box 4 6 36 64
use _0_0std_0_0cells_0_0AND2X1  splt_ar2__r
timestamp 1731220320
transform 1 0 1104 0 1 956
box 8 4 52 52
use _0_0std_0_0cells_0_0NOR2X1  splt_anor__ra
timestamp 1731220320
transform 1 0 1416 0 1 776
box 4 6 36 48
use _0_0std_0_0cells_0_0LATCH  splt_alatch_57_6
timestamp 1731220320
transform 1 0 1208 0 1 336
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_56_6
timestamp 1731220320
transform 1 0 1088 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_55_6
timestamp 1731220320
transform 1 0 784 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_54_6
timestamp 1731220320
transform 1 0 744 0 1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_53_6
timestamp 1731220320
transform 1 0 888 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_52_6
timestamp 1731220320
transform 1 0 792 0 1 764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_51_6
timestamp 1731220320
transform 1 0 688 0 1 956
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_50_6
timestamp 1731220320
transform 1 0 824 0 -1 1140
box 8 5 100 68
use _0_0std_0_0cells_0_0INVX1  snk_ar_ai
timestamp 1731220320
transform 1 0 1288 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  snk_ar_an
timestamp 1731220320
transform 1 0 1320 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_569_6
timestamp 1731220320
transform 1 0 864 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_568_6
timestamp 1731220320
transform 1 0 768 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_567_6
timestamp 1731220320
transform 1 0 648 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_566_6
timestamp 1731220320
transform 1 0 528 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_565_6
timestamp 1731220320
transform 1 0 456 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_564_6
timestamp 1731220320
transform 1 0 360 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_563_6
timestamp 1731220320
transform 1 0 296 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_562_6
timestamp 1731220320
transform 1 0 272 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_561_6
timestamp 1731220320
transform 1 0 216 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_560_6
timestamp 1731220320
transform 1 0 168 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_559_6
timestamp 1731220320
transform 1 0 128 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_558_6
timestamp 1731220320
transform 1 0 280 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_557_6
timestamp 1731220320
transform 1 0 224 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_556_6
timestamp 1731220320
transform 1 0 160 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_555_6
timestamp 1731220320
transform 1 0 128 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_554_6
timestamp 1731220320
transform 1 0 128 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_553_6
timestamp 1731220320
transform 1 0 160 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_552_6
timestamp 1731220320
transform 1 0 192 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_551_6
timestamp 1731220320
transform 1 0 240 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_550_6
timestamp 1731220320
transform 1 0 560 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_549_6
timestamp 1731220320
transform 1 0 432 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_548_6
timestamp 1731220320
transform 1 0 320 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_547_6
timestamp 1731220320
transform 1 0 256 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_546_6
timestamp 1731220320
transform 1 0 168 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_545_6
timestamp 1731220320
transform 1 0 128 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_544_6
timestamp 1731220320
transform 1 0 704 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_543_6
timestamp 1731220320
transform 1 0 536 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_542_6
timestamp 1731220320
transform 1 0 384 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_541_6
timestamp 1731220320
transform 1 0 312 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_540_6
timestamp 1731220320
transform 1 0 240 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_539_6
timestamp 1731220320
transform 1 0 184 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_538_6
timestamp 1731220320
transform 1 0 648 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_537_6
timestamp 1731220320
transform 1 0 520 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_536_6
timestamp 1731220320
transform 1 0 408 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_535_6
timestamp 1731220320
transform 1 0 208 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_534_6
timestamp 1731220320
transform 1 0 176 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_533_6
timestamp 1731220320
transform 1 0 144 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_532_6
timestamp 1731220320
transform 1 0 240 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_531_6
timestamp 1731220320
transform 1 0 272 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_530_6
timestamp 1731220320
transform 1 0 304 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_529_6
timestamp 1731220320
transform 1 0 336 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_528_6
timestamp 1731220320
transform 1 0 368 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_527_6
timestamp 1731220320
transform 1 0 400 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_526_6
timestamp 1731220320
transform 1 0 432 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_525_6
timestamp 1731220320
transform 1 0 464 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_524_6
timestamp 1731220320
transform 1 0 496 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_523_6
timestamp 1731220320
transform 1 0 528 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_522_6
timestamp 1731220320
transform 1 0 560 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_521_6
timestamp 1731220320
transform 1 0 592 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_520_6
timestamp 1731220320
transform 1 0 624 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_519_6
timestamp 1731220320
transform 1 0 656 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_518_6
timestamp 1731220320
transform 1 0 688 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_517_6
timestamp 1731220320
transform 1 0 720 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_516_6
timestamp 1731220320
transform 1 0 752 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_515_6
timestamp 1731220320
transform 1 0 784 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_514_6
timestamp 1731220320
transform 1 0 816 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_513_6
timestamp 1731220320
transform 1 0 848 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_512_6
timestamp 1731220320
transform 1 0 880 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_511_6
timestamp 1731220320
transform 1 0 912 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_510_6
timestamp 1731220320
transform 1 0 944 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_59_6
timestamp 1731220320
transform 1 0 976 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_58_6
timestamp 1731220320
transform 1 0 1040 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_57_6
timestamp 1731220320
transform 1 0 912 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_56_6
timestamp 1731220320
transform 1 0 784 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_55_6
timestamp 1731220320
transform 1 0 872 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_54_6
timestamp 1731220320
transform 1 0 1032 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_53_6
timestamp 1731220320
transform 1 0 992 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_52_6
timestamp 1731220320
transform 1 0 1056 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_51_6
timestamp 1731220320
transform 1 0 1072 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_50_6
timestamp 1731220320
transform 1 0 1072 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_57_6
timestamp 1731220320
transform 1 0 896 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_56_6
timestamp 1731220320
transform 1 0 1056 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_55_6
timestamp 1731220320
transform 1 0 784 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_54_6
timestamp 1731220320
transform 1 0 664 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_53_6
timestamp 1731220320
transform 1 0 856 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_52_6
timestamp 1731220320
transform 1 0 552 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_51_6
timestamp 1731220320
transform 1 0 808 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_50_6
timestamp 1731220320
transform 1 0 912 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar2_an
timestamp 1731220320
transform 1 0 1056 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  m_ar1_ai
timestamp 1731220320
transform 1 0 1032 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar1_an
timestamp 1731220320
transform 1 0 1064 0 -1 928
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  m_ar3_ai
timestamp 1731220320
transform 1 0 1432 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar3_an
timestamp 1731220320
transform 1 0 1360 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0AND2X1  m_aand__ct
timestamp 1731220320
transform 1 0 1360 0 -1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0OR2X1  m_aor__ca
timestamp 1731220320
transform 1 0 1008 0 1 776
box 4 4 48 48
use _0_0std_0_0cells_0_0INVX1  m_ar0_ai
timestamp 1731220320
transform 1 0 1160 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar0_an
timestamp 1731220320
transform 1 0 1192 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  m_ar4_ai
timestamp 1731220320
transform 1 0 1128 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar4_an
timestamp 1731220320
transform 1 0 1088 0 -1 1128
box 4 6 36 48
use _0_0cell_0_0ginvx0  m_ac1_acx1
timestamp 1731220320
transform 1 0 1104 0 -1 928
box 8 6 28 32
use _0_0cell_0_0gcelem3x0  m_ac1_acx0
timestamp 1731220320
transform 1 0 1136 0 -1 952
box 8 5 92 72
use _0_0cell_0_0ginvx0  m_ac0_acx1
timestamp 1731220320
transform 1 0 1232 0 -1 928
box 8 6 28 32
use _0_0cell_0_0gcelem3x0  m_ac0_acx0
timestamp 1731220320
transform 1 0 1264 0 -1 952
box 8 5 92 72
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_544_6
timestamp 1731220320
transform 1 0 544 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_543_6
timestamp 1731220320
transform 1 0 632 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_542_6
timestamp 1731220320
transform 1 0 600 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_541_6
timestamp 1731220320
transform 1 0 680 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_540_6
timestamp 1731220320
transform 1 0 768 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_539_6
timestamp 1731220320
transform 1 0 856 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_538_6
timestamp 1731220320
transform 1 0 896 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_537_6
timestamp 1731220320
transform 1 0 816 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_536_6
timestamp 1731220320
transform 1 0 736 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_535_6
timestamp 1731220320
transform 1 0 664 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_534_6
timestamp 1731220320
transform 1 0 600 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_533_6
timestamp 1731220320
transform 1 0 544 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_532_6
timestamp 1731220320
transform 1 0 512 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_531_6
timestamp 1731220320
transform 1 0 480 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_530_6
timestamp 1731220320
transform 1 0 448 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_529_6
timestamp 1731220320
transform 1 0 416 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_528_6
timestamp 1731220320
transform 1 0 384 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_527_6
timestamp 1731220320
transform 1 0 352 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_526_6
timestamp 1731220320
transform 1 0 320 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_525_6
timestamp 1731220320
transform 1 0 288 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_524_6
timestamp 1731220320
transform 1 0 256 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_523_6
timestamp 1731220320
transform 1 0 224 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_522_6
timestamp 1731220320
transform 1 0 192 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_521_6
timestamp 1731220320
transform 1 0 160 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_520_6
timestamp 1731220320
transform 1 0 128 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_519_6
timestamp 1731220320
transform 1 0 128 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_518_6
timestamp 1731220320
transform 1 0 160 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_517_6
timestamp 1731220320
transform 1 0 208 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_516_6
timestamp 1731220320
transform 1 0 256 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_515_6
timestamp 1731220320
transform 1 0 304 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_514_6
timestamp 1731220320
transform 1 0 360 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_513_6
timestamp 1731220320
transform 1 0 408 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_512_6
timestamp 1731220320
transform 1 0 464 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_511_6
timestamp 1731220320
transform 1 0 528 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_510_6
timestamp 1731220320
transform 1 0 592 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_59_6
timestamp 1731220320
transform 1 0 560 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_58_6
timestamp 1731220320
transform 1 0 528 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_57_6
timestamp 1731220320
transform 1 0 496 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_56_6
timestamp 1731220320
transform 1 0 512 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_55_6
timestamp 1731220320
transform 1 0 480 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_54_6
timestamp 1731220320
transform 1 0 448 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_53_6
timestamp 1731220320
transform 1 0 416 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_52_6
timestamp 1731220320
transform 1 0 384 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_51_6
timestamp 1731220320
transform 1 0 408 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_50_6
timestamp 1731220320
transform 1 0 440 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  m_ap_aand
timestamp 1731220320
transform 1 0 472 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  m_aand__cf
timestamp 1731220320
transform 1 0 1152 0 1 764
box 8 4 52 52
use _0_0std_0_0cells_0_0INVX1  m_ainv__cd
timestamp 1731220320
transform 1 0 1096 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad__cd_ainvs_51_6
timestamp 1731220320
transform 1 0 1416 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad__cd_ainvs_50_6
timestamp 1731220320
transform 1 0 1400 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0LATCH  m_alatch_57_6
timestamp 1731220320
transform 1 0 680 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_56_6
timestamp 1731220320
transform 1 0 944 0 1 176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_55_6
timestamp 1731220320
transform 1 0 672 0 1 176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_54_6
timestamp 1731220320
transform 1 0 512 0 1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_53_6
timestamp 1731220320
transform 1 0 592 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_52_6
timestamp 1731220320
transform 1 0 384 0 1 764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_51_6
timestamp 1731220320
transform 1 0 704 0 -1 940
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_50_6
timestamp 1731220320
transform 1 0 840 0 -1 940
box 8 5 100 68
use _0_0std_0_0cells_0_0MUX2X1  m_amux_57_6
timestamp 1731220320
transform 1 0 1344 0 1 336
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_56_6
timestamp 1731220320
transform 1 0 1192 0 -1 320
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_55_6
timestamp 1731220320
transform 1 0 824 0 1 176
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_54_6
timestamp 1731220320
transform 1 0 760 0 -1 744
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_53_6
timestamp 1731220320
transform 1 0 992 0 -1 744
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_52_6
timestamp 1731220320
transform 1 0 648 0 1 764
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_51_6
timestamp 1731220320
transform 1 0 808 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_50_6
timestamp 1731220320
transform 1 0 960 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_55_6
timestamp 1731220320
transform 1 0 1432 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_54_6
timestamp 1731220320
transform 1 0 1392 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_53_6
timestamp 1731220320
transform 1 0 1312 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_52_6
timestamp 1731220320
transform 1 0 1264 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_51_6
timestamp 1731220320
transform 1 0 1232 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_50_6
timestamp 1731220320
transform 1 0 1160 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ar0_ai
timestamp 1731220320
transform 1 0 968 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  c_ar0_an
timestamp 1731220320
transform 1 0 888 0 -1 1480
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_544_6
timestamp 1731220320
transform 1 0 256 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_543_6
timestamp 1731220320
transform 1 0 224 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_542_6
timestamp 1731220320
transform 1 0 192 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_541_6
timestamp 1731220320
transform 1 0 224 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_540_6
timestamp 1731220320
transform 1 0 192 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_539_6
timestamp 1731220320
transform 1 0 160 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_538_6
timestamp 1731220320
transform 1 0 128 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_537_6
timestamp 1731220320
transform 1 0 288 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_536_6
timestamp 1731220320
transform 1 0 320 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_535_6
timestamp 1731220320
transform 1 0 352 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_534_6
timestamp 1731220320
transform 1 0 384 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_533_6
timestamp 1731220320
transform 1 0 512 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_532_6
timestamp 1731220320
transform 1 0 480 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_531_6
timestamp 1731220320
transform 1 0 448 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_530_6
timestamp 1731220320
transform 1 0 416 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_529_6
timestamp 1731220320
transform 1 0 480 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_528_6
timestamp 1731220320
transform 1 0 448 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_527_6
timestamp 1731220320
transform 1 0 416 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_526_6
timestamp 1731220320
transform 1 0 384 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_525_6
timestamp 1731220320
transform 1 0 352 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_524_6
timestamp 1731220320
transform 1 0 320 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_523_6
timestamp 1731220320
transform 1 0 288 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_522_6
timestamp 1731220320
transform 1 0 256 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_521_6
timestamp 1731220320
transform 1 0 224 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_520_6
timestamp 1731220320
transform 1 0 192 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_519_6
timestamp 1731220320
transform 1 0 160 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_518_6
timestamp 1731220320
transform 1 0 128 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_517_6
timestamp 1731220320
transform 1 0 128 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_516_6
timestamp 1731220320
transform 1 0 160 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_515_6
timestamp 1731220320
transform 1 0 192 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_514_6
timestamp 1731220320
transform 1 0 224 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_513_6
timestamp 1731220320
transform 1 0 256 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_512_6
timestamp 1731220320
transform 1 0 288 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_511_6
timestamp 1731220320
transform 1 0 320 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_510_6
timestamp 1731220320
transform 1 0 448 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_59_6
timestamp 1731220320
transform 1 0 416 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_58_6
timestamp 1731220320
transform 1 0 384 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_57_6
timestamp 1731220320
transform 1 0 352 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_56_6
timestamp 1731220320
transform 1 0 544 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_55_6
timestamp 1731220320
transform 1 0 512 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_54_6
timestamp 1731220320
transform 1 0 480 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_53_6
timestamp 1731220320
transform 1 0 424 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_52_6
timestamp 1731220320
transform 1 0 392 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_51_6
timestamp 1731220320
transform 1 0 456 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_50_6
timestamp 1731220320
transform 1 0 488 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  c_ap_aand
timestamp 1731220320
transform 1 0 312 0 1 956
box 8 4 52 52
use _0_0cell_0_0ginvx0  c_ac_acx1
timestamp 1731220320
transform 1 0 768 0 -1 1480
box 8 6 28 32
use _0_0cell_0_0gcelem2x0  c_ac_acx0
timestamp 1731220320
transform 1 0 800 0 -1 1496
box 8 4 84 60
use _0_0std_0_0cells_0_0OR2X1  c_ar2_an
timestamp 1731220320
transform 1 0 1016 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  c_ar1_an
timestamp 1731220320
transform 1 0 1104 0 -1 1480
box 4 4 48 48
use _0_0cell_0_0gcelem2x0  c_ac__ra_acx0
timestamp 1731220320
transform 1 0 928 0 -1 1496
box 8 4 84 60
use _0_0std_0_0cells_0_0LATCH  c_alatch_57_6
timestamp 1731220320
transform 1 0 576 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_56_6
timestamp 1731220320
transform 1 0 888 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_55_6
timestamp 1731220320
transform 1 0 648 0 1 336
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_54_6
timestamp 1731220320
transform 1 0 280 0 -1 552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_53_6
timestamp 1731220320
transform 1 0 264 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_52_6
timestamp 1731220320
transform 1 0 208 0 1 764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_51_6
timestamp 1731220320
transform 1 0 568 0 -1 940
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_50_6
timestamp 1731220320
transform 1 0 560 0 1 956
box 8 5 100 68
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_569_6
timestamp 1731220320
transform 1 0 1272 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_568_6
timestamp 1731220320
transform 1 0 1304 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_567_6
timestamp 1731220320
transform 1 0 1336 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_566_6
timestamp 1731220320
transform 1 0 1368 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_565_6
timestamp 1731220320
transform 1 0 1400 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_564_6
timestamp 1731220320
transform 1 0 1432 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_563_6
timestamp 1731220320
transform 1 0 1408 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_562_6
timestamp 1731220320
transform 1 0 1416 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_561_6
timestamp 1731220320
transform 1 0 1472 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_560_6
timestamp 1731220320
transform 1 0 1520 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_559_6
timestamp 1731220320
transform 1 0 1568 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_558_6
timestamp 1731220320
transform 1 0 1552 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_557_6
timestamp 1731220320
transform 1 0 1512 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_556_6
timestamp 1731220320
transform 1 0 1472 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_555_6
timestamp 1731220320
transform 1 0 1552 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_554_6
timestamp 1731220320
transform 1 0 1584 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_553_6
timestamp 1731220320
transform 1 0 1584 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_552_6
timestamp 1731220320
transform 1 0 1584 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_551_6
timestamp 1731220320
transform 1 0 1552 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_550_6
timestamp 1731220320
transform 1 0 1616 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_549_6
timestamp 1731220320
transform 1 0 1648 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_548_6
timestamp 1731220320
transform 1 0 1648 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_547_6
timestamp 1731220320
transform 1 0 1616 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_546_6
timestamp 1731220320
transform 1 0 1648 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_545_6
timestamp 1731220320
transform 1 0 1648 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_544_6
timestamp 1731220320
transform 1 0 1616 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_543_6
timestamp 1731220320
transform 1 0 1648 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_542_6
timestamp 1731220320
transform 1 0 1616 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_541_6
timestamp 1731220320
transform 1 0 1584 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_540_6
timestamp 1731220320
transform 1 0 1616 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_539_6
timestamp 1731220320
transform 1 0 1648 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_538_6
timestamp 1731220320
transform 1 0 1648 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_537_6
timestamp 1731220320
transform 1 0 1600 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_536_6
timestamp 1731220320
transform 1 0 1536 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_535_6
timestamp 1731220320
transform 1 0 1472 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_534_6
timestamp 1731220320
transform 1 0 1648 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_533_6
timestamp 1731220320
transform 1 0 1616 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_532_6
timestamp 1731220320
transform 1 0 1584 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_531_6
timestamp 1731220320
transform 1 0 1552 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_530_6
timestamp 1731220320
transform 1 0 1512 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_529_6
timestamp 1731220320
transform 1 0 1472 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_528_6
timestamp 1731220320
transform 1 0 1512 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_527_6
timestamp 1731220320
transform 1 0 1552 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_526_6
timestamp 1731220320
transform 1 0 1584 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_525_6
timestamp 1731220320
transform 1 0 1616 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_524_6
timestamp 1731220320
transform 1 0 1648 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_523_6
timestamp 1731220320
transform 1 0 1648 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_522_6
timestamp 1731220320
transform 1 0 1616 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_521_6
timestamp 1731220320
transform 1 0 1584 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_520_6
timestamp 1731220320
transform 1 0 1552 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_519_6
timestamp 1731220320
transform 1 0 1512 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_518_6
timestamp 1731220320
transform 1 0 1648 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_517_6
timestamp 1731220320
transform 1 0 1616 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_516_6
timestamp 1731220320
transform 1 0 1584 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_515_6
timestamp 1731220320
transform 1 0 1552 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_514_6
timestamp 1731220320
transform 1 0 1512 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_513_6
timestamp 1731220320
transform 1 0 1512 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_512_6
timestamp 1731220320
transform 1 0 1552 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_511_6
timestamp 1731220320
transform 1 0 1552 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_510_6
timestamp 1731220320
transform 1 0 1512 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_59_6
timestamp 1731220320
transform 1 0 1520 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_58_6
timestamp 1731220320
transform 1 0 1528 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_57_6
timestamp 1731220320
transform 1 0 1512 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_56_6
timestamp 1731220320
transform 1 0 1472 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_55_6
timestamp 1731220320
transform 1 0 1512 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_54_6
timestamp 1731220320
transform 1 0 1528 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_53_6
timestamp 1731220320
transform 1 0 1464 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_52_6
timestamp 1731220320
transform 1 0 1392 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_51_6
timestamp 1731220320
transform 1 0 1240 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_50_6
timestamp 1731220320
transform 1 0 1168 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ar0_ai
timestamp 1731220320
transform 1 0 1016 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  a_ar0_an
timestamp 1731220320
transform 1 0 1056 0 1 1364
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_544_6
timestamp 1731220320
transform 1 0 160 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_543_6
timestamp 1731220320
transform 1 0 160 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_542_6
timestamp 1731220320
transform 1 0 224 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_541_6
timestamp 1731220320
transform 1 0 256 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_540_6
timestamp 1731220320
transform 1 0 288 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_539_6
timestamp 1731220320
transform 1 0 320 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_538_6
timestamp 1731220320
transform 1 0 352 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_537_6
timestamp 1731220320
transform 1 0 336 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_536_6
timestamp 1731220320
transform 1 0 464 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_535_6
timestamp 1731220320
transform 1 0 432 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_534_6
timestamp 1731220320
transform 1 0 400 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_533_6
timestamp 1731220320
transform 1 0 368 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_532_6
timestamp 1731220320
transform 1 0 304 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_531_6
timestamp 1731220320
transform 1 0 272 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_530_6
timestamp 1731220320
transform 1 0 240 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_529_6
timestamp 1731220320
transform 1 0 208 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_528_6
timestamp 1731220320
transform 1 0 176 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_527_6
timestamp 1731220320
transform 1 0 256 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_526_6
timestamp 1731220320
transform 1 0 224 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_525_6
timestamp 1731220320
transform 1 0 192 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_524_6
timestamp 1731220320
transform 1 0 160 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_523_6
timestamp 1731220320
transform 1 0 128 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_522_6
timestamp 1731220320
transform 1 0 192 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_521_6
timestamp 1731220320
transform 1 0 160 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_520_6
timestamp 1731220320
transform 1 0 128 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_519_6
timestamp 1731220320
transform 1 0 128 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_518_6
timestamp 1731220320
transform 1 0 128 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_517_6
timestamp 1731220320
transform 1 0 128 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_516_6
timestamp 1731220320
transform 1 0 128 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_515_6
timestamp 1731220320
transform 1 0 128 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_514_6
timestamp 1731220320
transform 1 0 160 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_513_6
timestamp 1731220320
transform 1 0 256 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_512_6
timestamp 1731220320
transform 1 0 544 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_511_6
timestamp 1731220320
transform 1 0 544 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_510_6
timestamp 1731220320
transform 1 0 512 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_59_6
timestamp 1731220320
transform 1 0 576 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_58_6
timestamp 1731220320
transform 1 0 608 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_57_6
timestamp 1731220320
transform 1 0 640 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_56_6
timestamp 1731220320
transform 1 0 640 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_55_6
timestamp 1731220320
transform 1 0 608 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_54_6
timestamp 1731220320
transform 1 0 576 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_53_6
timestamp 1731220320
transform 1 0 520 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_52_6
timestamp 1731220320
transform 1 0 552 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_51_6
timestamp 1731220320
transform 1 0 584 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_50_6
timestamp 1731220320
transform 1 0 736 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  a_ap_aand
timestamp 1731220320
transform 1 0 944 0 1 1156
box 8 4 52 52
use _0_0cell_0_0ginvx0  a_ac_acx1
timestamp 1731220320
transform 1 0 1104 0 1 1364
box 8 6 28 32
use _0_0cell_0_0gcelem3x0  a_ac_acx0
timestamp 1731220320
transform 1 0 1056 0 -1 1348
box 8 5 92 72
use _0_0std_0_0cells_0_0NOR2X1  a_ar2_an
timestamp 1731220320
transform 1 0 1016 0 -1 1324
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  a_ar1_ai
timestamp 1731220320
transform 1 0 1192 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  a_ar1_an
timestamp 1731220320
transform 1 0 1144 0 1 1364
box 4 6 36 48
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_57_6_al
timestamp 1731220320
transform 1 0 1200 0 1 560
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_57_6_anx
timestamp 1731220320
transform 1 0 1328 0 1 572
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_56_6_al
timestamp 1731220320
transform 1 0 1088 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_56_6_anx
timestamp 1731220320
transform 1 0 1192 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_55_6_al
timestamp 1731220320
transform 1 0 640 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_55_6_anx
timestamp 1731220320
transform 1 0 720 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_54_6_al
timestamp 1731220320
transform 1 0 384 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_54_6_anx
timestamp 1731220320
transform 1 0 464 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_53_6_al
timestamp 1731220320
transform 1 0 392 0 1 560
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_53_6_anx
timestamp 1731220320
transform 1 0 384 0 -1 736
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_52_6_al
timestamp 1731220320
transform 1 0 312 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_52_6_anx
timestamp 1731220320
transform 1 0 392 0 -1 932
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_51_6_al
timestamp 1731220320
transform 1 0 1000 0 1 1152
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_51_6_anx
timestamp 1731220320
transform 1 0 1080 0 1 1164
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_50_6_al
timestamp 1731220320
transform 1 0 816 0 -1 1340
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_50_6_anx
timestamp 1731220320
transform 1 0 832 0 1 1360
box 4 6 36 64
use _0_0std_0_0cells_0_0FAX1  a_aadder_57_6
timestamp 1731220320
transform 1 0 1256 0 -1 560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_56_6
timestamp 1731220320
transform 1 0 1072 0 1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_55_6
timestamp 1731220320
transform 1 0 752 0 1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_54_6
timestamp 1731220320
transform 1 0 504 0 -1 560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_53_6
timestamp 1731220320
transform 1 0 440 0 -1 752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_52_6
timestamp 1731220320
transform 1 0 432 0 -1 948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_51_6
timestamp 1731220320
transform 1 0 656 0 -1 1148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_50_6
timestamp 1731220320
transform 1 0 808 0 1 1148
box 3 5 132 108
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_57_6_al
timestamp 1731220320
transform 1 0 1080 0 -1 748
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_57_6_anx
timestamp 1731220320
transform 1 0 1160 0 -1 736
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_56_6_al
timestamp 1731220320
transform 1 0 984 0 1 560
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_56_6_anx
timestamp 1731220320
transform 1 0 1112 0 1 572
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_55_6_al
timestamp 1731220320
transform 1 0 768 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_55_6_anx
timestamp 1731220320
transform 1 0 864 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_54_6_al
timestamp 1731220320
transform 1 0 160 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_54_6_anx
timestamp 1731220320
transform 1 0 240 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_53_6_al
timestamp 1731220320
transform 1 0 128 0 -1 748
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_53_6_anx
timestamp 1731220320
transform 1 0 208 0 -1 736
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_52_6_al
timestamp 1731220320
transform 1 0 392 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_52_6_anx
timestamp 1731220320
transform 1 0 496 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_51_6_al
timestamp 1731220320
transform 1 0 896 0 -1 1340
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_51_6_anx
timestamp 1731220320
transform 1 0 976 0 -1 1328
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_50_6_al
timestamp 1731220320
transform 1 0 880 0 1 1348
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_50_6_anx
timestamp 1731220320
transform 1 0 968 0 1 1360
box 4 6 36 64
use _0_0std_0_0cells_0_0TIELOX1  a_atlo
timestamp 1731220320
transform 1 0 800 0 1 1364
box 8 6 28 37
use _0_0std_0_0cells_0_0OR2X1  i_ar0_an
timestamp 1731220320
transform 1 0 1456 0 1 1364
box 4 4 48 48
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_55_6
timestamp 1731220320
transform 1 0 1352 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_54_6
timestamp 1731220320
transform 1 0 1352 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_53_6
timestamp 1731220320
transform 1 0 1320 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_52_6
timestamp 1731220320
transform 1 0 1240 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_51_6
timestamp 1731220320
transform 1 0 1120 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_50_6
timestamp 1731220320
transform 1 0 1152 0 -1 1580
box 8 7 28 34
use _0_0cell_0_0ginvx0  i_ac_acx1
timestamp 1731220320
transform 1 0 1272 0 -1 1480
box 8 6 28 32
use _0_0cell_0_0gcelem2x0  i_ac_acx0
timestamp 1731220320
transform 1 0 1312 0 1 1348
box 8 4 84 60
use _0_0std_0_0cells_0_0INVX1  i_ar1_ai
timestamp 1731220320
transform 1 0 1192 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0OR2X1  i_ar1_an
timestamp 1731220320
transform 1 0 1240 0 1 1364
box 4 4 48 48
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_544_6
timestamp 1731220320
transform 1 0 656 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_543_6
timestamp 1731220320
transform 1 0 696 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_542_6
timestamp 1731220320
transform 1 0 680 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_541_6
timestamp 1731220320
transform 1 0 600 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_540_6
timestamp 1731220320
transform 1 0 616 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_539_6
timestamp 1731220320
transform 1 0 672 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_538_6
timestamp 1731220320
transform 1 0 672 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_537_6
timestamp 1731220320
transform 1 0 704 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_536_6
timestamp 1731220320
transform 1 0 736 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_535_6
timestamp 1731220320
transform 1 0 704 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_534_6
timestamp 1731220320
transform 1 0 672 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_533_6
timestamp 1731220320
transform 1 0 640 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_532_6
timestamp 1731220320
transform 1 0 608 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_531_6
timestamp 1731220320
transform 1 0 576 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_530_6
timestamp 1731220320
transform 1 0 544 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_529_6
timestamp 1731220320
transform 1 0 512 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_528_6
timestamp 1731220320
transform 1 0 480 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_527_6
timestamp 1731220320
transform 1 0 448 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_526_6
timestamp 1731220320
transform 1 0 416 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_525_6
timestamp 1731220320
transform 1 0 384 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_524_6
timestamp 1731220320
transform 1 0 352 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_523_6
timestamp 1731220320
transform 1 0 320 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_522_6
timestamp 1731220320
transform 1 0 288 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_521_6
timestamp 1731220320
transform 1 0 256 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_520_6
timestamp 1731220320
transform 1 0 224 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_519_6
timestamp 1731220320
transform 1 0 192 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_518_6
timestamp 1731220320
transform 1 0 160 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_517_6
timestamp 1731220320
transform 1 0 128 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_516_6
timestamp 1731220320
transform 1 0 168 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_515_6
timestamp 1731220320
transform 1 0 200 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_514_6
timestamp 1731220320
transform 1 0 232 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_513_6
timestamp 1731220320
transform 1 0 264 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_512_6
timestamp 1731220320
transform 1 0 328 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_511_6
timestamp 1731220320
transform 1 0 328 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_510_6
timestamp 1731220320
transform 1 0 392 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_59_6
timestamp 1731220320
transform 1 0 336 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_58_6
timestamp 1731220320
transform 1 0 392 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_57_6
timestamp 1731220320
transform 1 0 448 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_56_6
timestamp 1731220320
transform 1 0 504 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_55_6
timestamp 1731220320
transform 1 0 568 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_54_6
timestamp 1731220320
transform 1 0 704 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_53_6
timestamp 1731220320
transform 1 0 848 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_52_6
timestamp 1731220320
transform 1 0 952 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_51_6
timestamp 1731220320
transform 1 0 848 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_50_6
timestamp 1731220320
transform 1 0 744 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  i_ap_aand
timestamp 1731220320
transform 1 0 704 0 1 1352
box 8 4 52 52
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_57_6_al
timestamp 1731220320
transform 1 0 920 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_57_6_anx
timestamp 1731220320
transform 1 0 896 0 1 572
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_56_6_al
timestamp 1731220320
transform 1 0 936 0 1 332
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_56_6_anx
timestamp 1731220320
transform 1 0 1024 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_55_6_al
timestamp 1731220320
transform 1 0 528 0 1 332
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_55_6_anx
timestamp 1731220320
transform 1 0 608 0 1 344
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_54_6_al
timestamp 1731220320
transform 1 0 288 0 1 332
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_54_6_anx
timestamp 1731220320
transform 1 0 368 0 1 344
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_53_6_al
timestamp 1731220320
transform 1 0 272 0 1 560
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_53_6_anx
timestamp 1731220320
transform 1 0 200 0 1 572
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_52_6_al
timestamp 1731220320
transform 1 0 192 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_52_6_anx
timestamp 1731220320
transform 1 0 272 0 -1 932
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_51_6_al
timestamp 1731220320
transform 1 0 576 0 -1 1144
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_51_6_anx
timestamp 1731220320
transform 1 0 768 0 1 1164
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_50_6_al
timestamp 1731220320
transform 1 0 736 0 -1 1340
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_50_6_anx
timestamp 1731220320
transform 1 0 760 0 1 1360
box 4 6 36 64
use _0_0std_0_0cells_0_0INVX1  src_ar_ai
timestamp 1731220320
transform 1 0 944 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0OR2X1  src_ar_an
timestamp 1731220320
transform 1 0 976 0 -1 928
box 4 4 48 48
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_57_6
timestamp 1731220320
transform 1 0 1432 0 1 348
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_56_6
timestamp 1731220320
transform 1 0 1280 0 -1 308
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_55_6
timestamp 1731220320
transform 1 0 912 0 1 188
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_54_6
timestamp 1731220320
transform 1 0 712 0 -1 732
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_53_6
timestamp 1731220320
transform 1 0 944 0 1 776
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_52_6
timestamp 1731220320
transform 1 0 672 0 -1 928
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_51_6
timestamp 1731220320
transform 1 0 792 0 -1 1128
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_50_6
timestamp 1731220320
transform 1 0 992 0 -1 1128
box 8 6 28 37
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_55_6
timestamp 1731220320
transform 1 0 1448 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_54_6
timestamp 1731220320
transform 1 0 1416 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_53_6
timestamp 1731220320
transform 1 0 1368 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_52_6
timestamp 1731220320
transform 1 0 1336 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_51_6
timestamp 1731220320
transform 1 0 1400 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_50_6
timestamp 1731220320
transform 1 0 1416 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ar0_ai
timestamp 1731220320
transform 1 0 1488 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  c__copy_ar0_an
timestamp 1731220320
transform 1 0 1448 0 -1 1324
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_544_6
timestamp 1731220320
transform 1 0 1248 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_543_6
timestamp 1731220320
transform 1 0 1432 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_542_6
timestamp 1731220320
transform 1 0 1472 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_541_6
timestamp 1731220320
transform 1 0 1480 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_540_6
timestamp 1731220320
transform 1 0 1584 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_539_6
timestamp 1731220320
transform 1 0 1648 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_538_6
timestamp 1731220320
transform 1 0 1616 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_537_6
timestamp 1731220320
transform 1 0 1584 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_536_6
timestamp 1731220320
transform 1 0 1616 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_535_6
timestamp 1731220320
transform 1 0 1648 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_534_6
timestamp 1731220320
transform 1 0 1648 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_533_6
timestamp 1731220320
transform 1 0 1616 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_532_6
timestamp 1731220320
transform 1 0 1584 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_531_6
timestamp 1731220320
transform 1 0 1552 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_530_6
timestamp 1731220320
transform 1 0 1648 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_529_6
timestamp 1731220320
transform 1 0 1616 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_528_6
timestamp 1731220320
transform 1 0 1576 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_527_6
timestamp 1731220320
transform 1 0 1552 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_526_6
timestamp 1731220320
transform 1 0 1584 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_525_6
timestamp 1731220320
transform 1 0 1648 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_524_6
timestamp 1731220320
transform 1 0 1616 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_523_6
timestamp 1731220320
transform 1 0 1592 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_522_6
timestamp 1731220320
transform 1 0 1648 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_521_6
timestamp 1731220320
transform 1 0 1648 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_520_6
timestamp 1731220320
transform 1 0 1600 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_519_6
timestamp 1731220320
transform 1 0 1560 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_518_6
timestamp 1731220320
transform 1 0 1648 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_517_6
timestamp 1731220320
transform 1 0 1648 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_516_6
timestamp 1731220320
transform 1 0 1552 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_515_6
timestamp 1731220320
transform 1 0 1432 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_514_6
timestamp 1731220320
transform 1 0 1648 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_513_6
timestamp 1731220320
transform 1 0 1616 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_512_6
timestamp 1731220320
transform 1 0 1560 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_511_6
timestamp 1731220320
transform 1 0 1512 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_510_6
timestamp 1731220320
transform 1 0 1456 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_59_6
timestamp 1731220320
transform 1 0 1400 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_58_6
timestamp 1731220320
transform 1 0 1328 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_57_6
timestamp 1731220320
transform 1 0 1248 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_56_6
timestamp 1731220320
transform 1 0 1152 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_55_6
timestamp 1731220320
transform 1 0 1176 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_54_6
timestamp 1731220320
transform 1 0 1312 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_53_6
timestamp 1731220320
transform 1 0 1352 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_52_6
timestamp 1731220320
transform 1 0 1456 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_51_6
timestamp 1731220320
transform 1 0 1432 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_50_6
timestamp 1731220320
transform 1 0 1408 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  c__copy_ap_aand
timestamp 1731220320
transform 1 0 1280 0 1 1156
box 8 4 52 52
use _0_0cell_0_0ginvx0  c__copy_ac_acx1
timestamp 1731220320
transform 1 0 1384 0 -1 1324
box 8 6 28 32
use _0_0cell_0_0gcelem2x0  c__copy_ac_acx0
timestamp 1731220320
transform 1 0 1296 0 -1 1340
box 8 4 84 60
use _0_0std_0_0cells_0_0OR2X1  c__copy_ar2_an
timestamp 1731220320
transform 1 0 1152 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  c__copy_ar1_an
timestamp 1731220320
transform 1 0 1192 0 1 1168
box 4 4 48 48
use _0_0cell_0_0gcelem2x0  c__copy_ac__ra_acx0
timestamp 1731220320
transform 1 0 1208 0 -1 1340
box 8 4 84 60
use _0_0std_0_0cells_0_0LATCH  c__copy_alatch_50_6
timestamp 1731220320
transform 1 0 1312 0 -1 1140
box 8 5 100 68
<< labels >>
rlabel m1 s 638 1796 642 1800 6 L.d[0]
port 0 nsew signal input
rlabel m1 s 80 1666 84 1670 6 L.d[1]
port 1 nsew signal input
rlabel m1 s 80 1398 84 1402 6 L.d[2]
port 2 nsew signal input
rlabel m1 s 80 866 84 870 6 L.d[3]
port 3 nsew signal input
rlabel m1 s 80 470 84 474 6 L.d[4]
port 4 nsew signal input
rlabel m1 s 80 602 84 606 6 L.d[5]
port 5 nsew signal input
rlabel m1 s 1748 262 1752 266 6 L.d[6]
port 6 nsew signal input
rlabel m1 s 1748 454 1752 458 6 L.d[7]
port 7 nsew signal input
rlabel m1 s 1748 1222 1752 1226 6 L.r
port 8 nsew signal input
rlabel m1 s 1190 1796 1194 1800 6 L.a
port 9 nsew signal tristate
rlabel m1 s 1748 646 1752 650 6 C.d[0]
port 10 nsew signal input
rlabel m1 s 1748 838 1752 842 6 C.r
port 11 nsew signal input
rlabel m1 s 1748 1030 1752 1034 6 C.a
port 12 nsew signal tristate
rlabel m1 s 80 1534 84 1538 6 R.d[0]
port 13 nsew signal tristate
rlabel m1 s 80 1266 84 1270 6 R.d[1]
port 14 nsew signal tristate
rlabel m1 s 80 1002 84 1006 6 R.d[2]
port 15 nsew signal tristate
rlabel m1 s 80 734 84 738 6 R.d[3]
port 16 nsew signal tristate
rlabel m1 s 80 334 84 338 6 R.d[4]
port 17 nsew signal tristate
rlabel m1 s 80 202 84 206 6 R.d[5]
port 18 nsew signal tristate
rlabel m1 s 1190 72 1194 76 6 R.d[6]
port 19 nsew signal tristate
rlabel m1 s 638 72 642 76 6 R.d[7]
port 20 nsew signal tristate
rlabel m1 s 1748 1414 1752 1418 6 R.r
port 21 nsew signal tristate
rlabel m1 s 1748 1606 1752 1610 6 R.a
port 22 nsew signal input
rlabel m1 s 80 1134 84 1138 6 Reset
port 23 nsew signal input
<< end >>
