magic
tech sky130l
timestamp 1731001196
<< m1 >>
rect 208 1139 212 1167
rect 384 1139 388 1167
rect 472 1139 476 1167
rect 480 1131 484 1167
rect 648 1139 652 1167
rect 736 1139 740 1167
rect 232 1099 236 1127
rect 320 1099 324 1127
rect 744 1131 748 1167
rect 408 1099 412 1127
rect 384 863 388 887
rect 480 831 484 859
rect 776 595 780 615
rect 912 559 916 591
rect 480 451 484 479
rect 568 451 572 539
rect 368 419 372 447
rect 728 419 732 447
rect 960 415 964 443
rect 224 315 228 339
rect 264 179 268 203
<< m2c >>
rect 111 1181 115 1185
rect 1111 1181 1115 1185
rect 208 1167 212 1171
rect 111 1163 115 1167
rect 208 1135 212 1139
rect 384 1167 388 1171
rect 384 1135 388 1139
rect 472 1167 476 1171
rect 472 1135 476 1139
rect 480 1167 484 1171
rect 648 1167 652 1171
rect 648 1135 652 1139
rect 736 1167 740 1171
rect 736 1135 740 1139
rect 744 1167 748 1171
rect 232 1127 236 1131
rect 111 1101 115 1105
rect 232 1095 236 1099
rect 320 1127 324 1131
rect 320 1095 324 1099
rect 408 1127 412 1131
rect 480 1127 484 1131
rect 1111 1163 1115 1167
rect 744 1127 748 1131
rect 1111 1101 1115 1105
rect 408 1095 412 1099
rect 111 1083 115 1087
rect 1111 1083 1115 1087
rect 111 1037 115 1041
rect 1111 1037 1115 1041
rect 111 1019 115 1023
rect 1111 1019 1115 1023
rect 111 965 115 969
rect 1111 965 1115 969
rect 111 947 115 951
rect 1111 947 1115 951
rect 111 901 115 905
rect 1111 901 1115 905
rect 384 887 388 891
rect 111 883 115 887
rect 1111 883 1115 887
rect 384 859 388 863
rect 480 859 484 863
rect 111 829 115 833
rect 480 827 484 831
rect 1111 829 1115 833
rect 111 811 115 815
rect 1111 811 1115 815
rect 111 765 115 769
rect 1111 765 1115 769
rect 111 747 115 751
rect 1111 747 1115 751
rect 111 697 115 701
rect 1111 697 1115 701
rect 111 679 115 683
rect 1111 679 1115 683
rect 111 629 115 633
rect 1111 629 1115 633
rect 776 615 780 619
rect 111 611 115 615
rect 1111 611 1115 615
rect 776 591 780 595
rect 912 591 916 595
rect 111 557 115 561
rect 912 555 916 559
rect 1111 557 1115 561
rect 111 539 115 543
rect 568 539 572 543
rect 1111 539 1115 543
rect 111 493 115 497
rect 480 479 484 483
rect 111 475 115 479
rect 368 447 372 451
rect 480 447 484 451
rect 1111 493 1115 497
rect 1111 475 1115 479
rect 568 447 572 451
rect 728 447 732 451
rect 111 417 115 421
rect 368 415 372 419
rect 728 415 732 419
rect 960 443 964 447
rect 1111 417 1115 421
rect 960 411 964 415
rect 111 399 115 403
rect 1111 399 1115 403
rect 111 353 115 357
rect 1111 353 1115 357
rect 224 339 228 343
rect 111 335 115 339
rect 1111 335 1115 339
rect 224 311 228 315
rect 111 281 115 285
rect 1111 281 1115 285
rect 111 263 115 267
rect 1111 263 1115 267
rect 111 217 115 221
rect 1111 217 1115 221
rect 264 203 268 207
rect 111 199 115 203
rect 1111 199 1115 203
rect 264 175 268 179
rect 111 133 115 137
rect 1111 133 1115 137
rect 111 115 115 119
rect 1111 115 1115 119
<< m2 >>
rect 134 1200 140 1201
rect 134 1196 135 1200
rect 139 1196 140 1200
rect 134 1195 140 1196
rect 222 1200 228 1201
rect 222 1196 223 1200
rect 227 1196 228 1200
rect 222 1195 228 1196
rect 310 1200 316 1201
rect 310 1196 311 1200
rect 315 1196 316 1200
rect 310 1195 316 1196
rect 398 1200 404 1201
rect 398 1196 399 1200
rect 403 1196 404 1200
rect 398 1195 404 1196
rect 486 1200 492 1201
rect 486 1196 487 1200
rect 491 1196 492 1200
rect 486 1195 492 1196
rect 574 1200 580 1201
rect 574 1196 575 1200
rect 579 1196 580 1200
rect 574 1195 580 1196
rect 662 1200 668 1201
rect 662 1196 663 1200
rect 667 1196 668 1200
rect 662 1195 668 1196
rect 750 1200 756 1201
rect 750 1196 751 1200
rect 755 1196 756 1200
rect 750 1195 756 1196
rect 110 1185 116 1186
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 110 1180 116 1181
rect 1110 1185 1116 1186
rect 1110 1181 1111 1185
rect 1115 1181 1116 1185
rect 1110 1180 1116 1181
rect 207 1171 213 1172
rect 207 1170 208 1171
rect 197 1168 208 1170
rect 110 1167 116 1168
rect 110 1163 111 1167
rect 115 1163 116 1167
rect 207 1167 208 1168
rect 212 1167 213 1171
rect 290 1171 296 1172
rect 290 1170 291 1171
rect 285 1168 291 1170
rect 207 1166 213 1167
rect 290 1167 291 1168
rect 295 1167 296 1171
rect 383 1171 389 1172
rect 383 1170 384 1171
rect 373 1168 384 1170
rect 290 1166 296 1167
rect 383 1167 384 1168
rect 388 1167 389 1171
rect 471 1171 477 1172
rect 471 1170 472 1171
rect 461 1168 472 1170
rect 383 1166 389 1167
rect 471 1167 472 1168
rect 476 1167 477 1171
rect 471 1166 477 1167
rect 479 1171 485 1172
rect 479 1167 480 1171
rect 484 1170 485 1171
rect 647 1171 653 1172
rect 647 1170 648 1171
rect 484 1168 513 1170
rect 637 1168 648 1170
rect 484 1167 485 1168
rect 479 1166 485 1167
rect 647 1167 648 1168
rect 652 1167 653 1171
rect 735 1171 741 1172
rect 735 1170 736 1171
rect 725 1168 736 1170
rect 647 1166 653 1167
rect 735 1167 736 1168
rect 740 1167 741 1171
rect 735 1166 741 1167
rect 743 1171 749 1172
rect 743 1167 744 1171
rect 748 1170 749 1171
rect 748 1168 777 1170
rect 748 1167 749 1168
rect 743 1166 749 1167
rect 1110 1167 1116 1168
rect 110 1162 116 1163
rect 1110 1163 1111 1167
rect 1115 1163 1116 1167
rect 1110 1162 1116 1163
rect 142 1155 148 1156
rect 142 1151 143 1155
rect 147 1151 148 1155
rect 142 1150 148 1151
rect 230 1155 236 1156
rect 230 1151 231 1155
rect 235 1151 236 1155
rect 230 1150 236 1151
rect 318 1155 324 1156
rect 318 1151 319 1155
rect 323 1151 324 1155
rect 318 1150 324 1151
rect 406 1155 412 1156
rect 406 1151 407 1155
rect 411 1151 412 1155
rect 406 1150 412 1151
rect 494 1155 500 1156
rect 494 1151 495 1155
rect 499 1151 500 1155
rect 494 1150 500 1151
rect 582 1155 588 1156
rect 582 1151 583 1155
rect 587 1151 588 1155
rect 582 1150 588 1151
rect 670 1155 676 1156
rect 670 1151 671 1155
rect 675 1151 676 1155
rect 670 1150 676 1151
rect 758 1155 764 1156
rect 758 1151 759 1155
rect 763 1151 764 1155
rect 758 1150 764 1151
rect 522 1147 528 1148
rect 522 1143 523 1147
rect 527 1143 528 1147
rect 522 1142 528 1143
rect 207 1139 213 1140
rect 207 1135 208 1139
rect 212 1138 213 1139
rect 260 1138 262 1141
rect 212 1136 262 1138
rect 290 1139 296 1140
rect 212 1135 213 1136
rect 207 1134 213 1135
rect 290 1135 291 1139
rect 295 1138 296 1139
rect 348 1138 350 1141
rect 295 1136 350 1138
rect 383 1139 389 1140
rect 295 1135 296 1136
rect 290 1134 296 1135
rect 383 1135 384 1139
rect 388 1138 389 1139
rect 436 1138 438 1141
rect 388 1136 438 1138
rect 471 1139 477 1140
rect 388 1135 389 1136
rect 383 1134 389 1135
rect 471 1135 472 1139
rect 476 1138 477 1139
rect 612 1138 614 1141
rect 476 1136 614 1138
rect 647 1139 653 1140
rect 476 1135 477 1136
rect 471 1134 477 1135
rect 647 1135 648 1139
rect 652 1138 653 1139
rect 700 1138 702 1141
rect 652 1136 702 1138
rect 735 1139 741 1140
rect 652 1135 653 1136
rect 647 1134 653 1135
rect 735 1135 736 1139
rect 740 1138 741 1139
rect 788 1138 790 1141
rect 740 1136 790 1138
rect 740 1135 741 1136
rect 735 1134 741 1135
rect 231 1131 237 1132
rect 231 1130 232 1131
rect 196 1128 232 1130
rect 192 1126 198 1128
rect 231 1127 232 1128
rect 236 1127 237 1131
rect 319 1131 325 1132
rect 319 1130 320 1131
rect 284 1128 320 1130
rect 231 1126 237 1127
rect 280 1126 286 1128
rect 319 1127 320 1128
rect 324 1127 325 1131
rect 407 1131 413 1132
rect 407 1130 408 1131
rect 372 1128 408 1130
rect 319 1126 325 1127
rect 368 1126 374 1128
rect 407 1127 408 1128
rect 412 1127 413 1131
rect 479 1131 485 1132
rect 479 1130 480 1131
rect 460 1128 480 1130
rect 407 1126 413 1127
rect 456 1126 462 1128
rect 479 1127 480 1128
rect 484 1127 485 1131
rect 479 1126 485 1127
rect 522 1131 528 1132
rect 522 1127 523 1131
rect 527 1130 528 1131
rect 743 1131 749 1132
rect 743 1130 744 1131
rect 527 1128 744 1130
rect 527 1127 528 1128
rect 522 1126 528 1127
rect 743 1127 744 1128
rect 748 1127 749 1131
rect 743 1126 749 1127
rect 189 1124 194 1126
rect 277 1124 282 1126
rect 365 1124 370 1126
rect 453 1124 458 1126
rect 158 1117 164 1118
rect 158 1113 159 1117
rect 163 1113 164 1117
rect 158 1112 164 1113
rect 246 1117 252 1118
rect 246 1113 247 1117
rect 251 1113 252 1117
rect 246 1112 252 1113
rect 334 1117 340 1118
rect 334 1113 335 1117
rect 339 1113 340 1117
rect 334 1112 340 1113
rect 422 1117 428 1118
rect 422 1113 423 1117
rect 427 1113 428 1117
rect 422 1112 428 1113
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 110 1100 116 1101
rect 1110 1105 1116 1106
rect 1110 1101 1111 1105
rect 1115 1101 1116 1105
rect 1110 1100 1116 1101
rect 231 1099 237 1100
rect 231 1095 232 1099
rect 236 1098 237 1099
rect 319 1099 325 1100
rect 236 1096 265 1098
rect 236 1095 237 1096
rect 231 1094 237 1095
rect 319 1095 320 1099
rect 324 1098 325 1099
rect 407 1099 413 1100
rect 324 1096 353 1098
rect 324 1095 325 1096
rect 319 1094 325 1095
rect 407 1095 408 1099
rect 412 1098 413 1099
rect 412 1096 441 1098
rect 412 1095 413 1096
rect 407 1094 413 1095
rect 110 1087 116 1088
rect 110 1083 111 1087
rect 115 1083 116 1087
rect 246 1087 252 1088
rect 246 1086 247 1087
rect 209 1084 247 1086
rect 110 1082 116 1083
rect 246 1083 247 1084
rect 251 1083 252 1087
rect 246 1082 252 1083
rect 1110 1087 1116 1088
rect 1110 1083 1111 1087
rect 1115 1083 1116 1087
rect 1110 1082 1116 1083
rect 150 1072 156 1073
rect 150 1068 151 1072
rect 155 1068 156 1072
rect 150 1067 156 1068
rect 238 1072 244 1073
rect 238 1068 239 1072
rect 243 1068 244 1072
rect 238 1067 244 1068
rect 326 1072 332 1073
rect 326 1068 327 1072
rect 331 1068 332 1072
rect 326 1067 332 1068
rect 414 1072 420 1073
rect 414 1068 415 1072
rect 419 1068 420 1072
rect 414 1067 420 1068
rect 134 1056 140 1057
rect 134 1052 135 1056
rect 139 1052 140 1056
rect 134 1051 140 1052
rect 222 1056 228 1057
rect 222 1052 223 1056
rect 227 1052 228 1056
rect 222 1051 228 1052
rect 310 1056 316 1057
rect 310 1052 311 1056
rect 315 1052 316 1056
rect 310 1051 316 1052
rect 398 1056 404 1057
rect 398 1052 399 1056
rect 403 1052 404 1056
rect 398 1051 404 1052
rect 378 1043 384 1044
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 378 1039 379 1043
rect 383 1042 384 1043
rect 383 1040 417 1042
rect 1110 1041 1116 1042
rect 383 1039 384 1040
rect 378 1038 384 1039
rect 110 1036 116 1037
rect 1110 1037 1111 1041
rect 1115 1037 1116 1041
rect 1110 1036 1116 1037
rect 318 1031 324 1032
rect 202 1027 208 1028
rect 202 1026 203 1027
rect 197 1024 203 1026
rect 110 1023 116 1024
rect 110 1019 111 1023
rect 115 1019 116 1023
rect 202 1023 203 1024
rect 207 1023 208 1027
rect 318 1027 319 1031
rect 323 1027 324 1031
rect 318 1026 324 1027
rect 406 1031 412 1032
rect 406 1027 407 1031
rect 411 1027 412 1031
rect 406 1026 412 1027
rect 285 1024 321 1026
rect 373 1024 410 1026
rect 202 1022 208 1023
rect 1110 1023 1116 1024
rect 110 1018 116 1019
rect 1110 1019 1111 1023
rect 1115 1019 1116 1023
rect 1110 1018 1116 1019
rect 142 1011 148 1012
rect 142 1007 143 1011
rect 147 1007 148 1011
rect 142 1006 148 1007
rect 230 1011 236 1012
rect 230 1007 231 1011
rect 235 1007 236 1011
rect 230 1006 236 1007
rect 318 1011 324 1012
rect 318 1007 319 1011
rect 323 1007 324 1011
rect 318 1006 324 1007
rect 406 1011 412 1012
rect 406 1007 407 1011
rect 411 1007 412 1011
rect 406 1006 412 1007
rect 328 1004 350 1006
rect 416 1004 438 1006
rect 170 1003 176 1004
rect 170 999 171 1003
rect 175 999 176 1003
rect 170 998 176 999
rect 258 1003 264 1004
rect 258 999 259 1003
rect 263 999 264 1003
rect 258 998 264 999
rect 326 1003 332 1004
rect 326 999 327 1003
rect 331 999 332 1003
rect 348 1001 350 1004
rect 414 1003 420 1004
rect 326 998 332 999
rect 414 999 415 1003
rect 419 999 420 1003
rect 436 1001 438 1004
rect 414 998 420 999
rect 202 995 208 996
rect 202 994 203 995
rect 180 992 203 994
rect 176 990 182 992
rect 202 991 203 992
rect 207 991 208 995
rect 202 990 208 991
rect 258 991 264 992
rect 173 988 178 990
rect 258 987 259 991
rect 263 987 264 991
rect 258 986 264 987
rect 346 991 352 992
rect 346 987 347 991
rect 351 987 352 991
rect 346 986 352 987
rect 434 991 440 992
rect 434 987 435 991
rect 439 987 440 991
rect 434 986 440 987
rect 142 981 148 982
rect 142 977 143 981
rect 147 977 148 981
rect 142 976 148 977
rect 230 981 236 982
rect 230 977 231 981
rect 235 977 236 981
rect 230 976 236 977
rect 318 981 324 982
rect 318 977 319 981
rect 323 977 324 981
rect 318 976 324 977
rect 406 981 412 982
rect 406 977 407 981
rect 411 977 412 981
rect 406 976 412 977
rect 110 969 116 970
rect 110 965 111 969
rect 115 965 116 969
rect 110 964 116 965
rect 1110 969 1116 970
rect 1110 965 1111 969
rect 1115 965 1116 969
rect 1110 964 1116 965
rect 230 963 236 964
rect 230 962 231 963
rect 197 960 231 962
rect 230 959 231 960
rect 235 959 236 963
rect 318 963 324 964
rect 318 962 319 963
rect 285 960 319 962
rect 230 958 236 959
rect 318 959 319 960
rect 323 959 324 963
rect 406 963 412 964
rect 406 962 407 963
rect 373 960 407 962
rect 318 958 324 959
rect 406 959 407 960
rect 411 959 412 963
rect 406 958 412 959
rect 110 951 116 952
rect 110 947 111 951
rect 115 947 116 951
rect 1110 951 1116 952
rect 457 948 470 950
rect 110 946 116 947
rect 466 947 472 948
rect 466 943 467 947
rect 471 943 472 947
rect 1110 947 1111 951
rect 1115 947 1116 951
rect 1110 946 1116 947
rect 466 942 472 943
rect 134 936 140 937
rect 134 932 135 936
rect 139 932 140 936
rect 134 931 140 932
rect 222 936 228 937
rect 222 932 223 936
rect 227 932 228 936
rect 222 931 228 932
rect 310 936 316 937
rect 310 932 311 936
rect 315 932 316 936
rect 310 931 316 932
rect 398 936 404 937
rect 398 932 399 936
rect 403 932 404 936
rect 398 931 404 932
rect 134 920 140 921
rect 134 916 135 920
rect 139 916 140 920
rect 134 915 140 916
rect 222 920 228 921
rect 222 916 223 920
rect 227 916 228 920
rect 222 915 228 916
rect 310 920 316 921
rect 310 916 311 920
rect 315 916 316 920
rect 310 915 316 916
rect 398 920 404 921
rect 398 916 399 920
rect 403 916 404 920
rect 398 915 404 916
rect 110 905 116 906
rect 110 901 111 905
rect 115 901 116 905
rect 110 900 116 901
rect 1110 905 1116 906
rect 1110 901 1111 905
rect 1115 901 1116 905
rect 1110 900 1116 901
rect 206 891 212 892
rect 110 887 116 888
rect 110 883 111 887
rect 115 883 116 887
rect 110 882 116 883
rect 196 884 198 889
rect 206 887 207 891
rect 211 890 212 891
rect 290 891 296 892
rect 211 888 249 890
rect 211 887 212 888
rect 206 886 212 887
rect 290 887 291 891
rect 295 890 296 891
rect 383 891 389 892
rect 295 888 337 890
rect 295 887 296 888
rect 290 886 296 887
rect 383 887 384 891
rect 388 890 389 891
rect 388 888 425 890
rect 388 887 389 888
rect 383 886 389 887
rect 1110 887 1116 888
rect 196 883 204 884
rect 196 880 199 883
rect 198 879 199 880
rect 203 879 204 883
rect 1110 883 1111 887
rect 1115 883 1116 887
rect 1110 882 1116 883
rect 198 878 204 879
rect 142 875 148 876
rect 142 871 143 875
rect 147 871 148 875
rect 142 870 148 871
rect 230 875 236 876
rect 230 871 231 875
rect 235 871 236 875
rect 230 870 236 871
rect 318 875 324 876
rect 318 871 319 875
rect 323 871 324 875
rect 318 870 324 871
rect 406 875 412 876
rect 406 871 407 875
rect 411 871 412 875
rect 406 870 412 871
rect 206 863 212 864
rect 206 862 207 863
rect 173 860 207 862
rect 206 859 207 860
rect 211 859 212 863
rect 290 863 296 864
rect 290 862 291 863
rect 261 860 291 862
rect 206 858 212 859
rect 290 859 291 860
rect 295 859 296 863
rect 383 863 389 864
rect 383 862 384 863
rect 349 860 384 862
rect 290 858 296 859
rect 383 859 384 860
rect 388 859 389 863
rect 466 863 472 864
rect 466 862 467 863
rect 437 860 467 862
rect 383 858 389 859
rect 466 859 467 860
rect 471 859 472 863
rect 466 858 472 859
rect 479 863 485 864
rect 479 859 480 863
rect 484 862 485 863
rect 484 860 526 862
rect 484 859 485 860
rect 479 858 485 859
rect 180 856 202 858
rect 176 854 182 856
rect 198 855 204 856
rect 173 852 178 854
rect 198 851 199 855
rect 203 851 204 855
rect 198 850 204 851
rect 258 855 264 856
rect 258 851 259 855
rect 263 851 264 855
rect 258 850 264 851
rect 346 855 352 856
rect 346 851 347 855
rect 351 851 352 855
rect 346 850 352 851
rect 434 855 440 856
rect 524 855 526 860
rect 434 851 435 855
rect 439 851 440 855
rect 434 850 440 851
rect 142 845 148 846
rect 142 841 143 845
rect 147 841 148 845
rect 142 840 148 841
rect 230 845 236 846
rect 230 841 231 845
rect 235 841 236 845
rect 230 840 236 841
rect 318 845 324 846
rect 318 841 319 845
rect 323 841 324 845
rect 318 840 324 841
rect 406 845 412 846
rect 406 841 407 845
rect 411 841 412 845
rect 406 840 412 841
rect 494 845 500 846
rect 494 841 495 845
rect 499 841 500 845
rect 494 840 500 841
rect 110 833 116 834
rect 110 829 111 833
rect 115 829 116 833
rect 1110 833 1116 834
rect 479 831 485 832
rect 479 830 480 831
rect 110 828 116 829
rect 461 828 480 830
rect 230 827 236 828
rect 230 826 231 827
rect 197 824 231 826
rect 230 823 231 824
rect 235 823 236 827
rect 318 827 324 828
rect 318 826 319 827
rect 285 824 319 826
rect 230 822 236 823
rect 318 823 319 824
rect 323 823 324 827
rect 406 827 412 828
rect 406 826 407 827
rect 373 824 407 826
rect 318 822 324 823
rect 406 823 407 824
rect 411 823 412 827
rect 479 827 480 828
rect 484 827 485 831
rect 1110 829 1111 833
rect 1115 829 1116 833
rect 1110 828 1116 829
rect 479 826 485 827
rect 406 822 412 823
rect 110 815 116 816
rect 110 811 111 815
rect 115 811 116 815
rect 110 810 116 811
rect 474 815 480 816
rect 474 811 475 815
rect 479 814 480 815
rect 1110 815 1116 816
rect 479 812 505 814
rect 479 811 480 812
rect 474 810 480 811
rect 1110 811 1111 815
rect 1115 811 1116 815
rect 1110 810 1116 811
rect 134 800 140 801
rect 134 796 135 800
rect 139 796 140 800
rect 134 795 140 796
rect 222 800 228 801
rect 222 796 223 800
rect 227 796 228 800
rect 222 795 228 796
rect 310 800 316 801
rect 310 796 311 800
rect 315 796 316 800
rect 310 795 316 796
rect 398 800 404 801
rect 398 796 399 800
rect 403 796 404 800
rect 398 795 404 796
rect 486 800 492 801
rect 486 796 487 800
rect 491 796 492 800
rect 486 795 492 796
rect 134 784 140 785
rect 134 780 135 784
rect 139 780 140 784
rect 134 779 140 780
rect 230 784 236 785
rect 230 780 231 784
rect 235 780 236 784
rect 230 779 236 780
rect 358 784 364 785
rect 358 780 359 784
rect 363 780 364 784
rect 358 779 364 780
rect 502 784 508 785
rect 502 780 503 784
rect 507 780 508 784
rect 502 779 508 780
rect 646 784 652 785
rect 646 780 647 784
rect 651 780 652 784
rect 646 779 652 780
rect 798 784 804 785
rect 798 780 799 784
rect 803 780 804 784
rect 798 779 804 780
rect 958 784 964 785
rect 958 780 959 784
rect 963 780 964 784
rect 958 779 964 780
rect 110 769 116 770
rect 110 765 111 769
rect 115 765 116 769
rect 561 768 658 770
rect 1110 769 1116 770
rect 110 764 116 765
rect 654 767 660 768
rect 654 763 655 767
rect 659 763 660 767
rect 1110 765 1111 769
rect 1115 765 1116 769
rect 1110 764 1116 765
rect 654 762 660 763
rect 366 759 372 760
rect 366 758 367 759
rect 319 756 367 758
rect 214 755 220 756
rect 214 754 215 755
rect 197 752 215 754
rect 110 751 116 752
rect 110 747 111 751
rect 115 747 116 751
rect 214 751 215 752
rect 219 751 220 755
rect 319 754 321 756
rect 366 755 367 756
rect 371 755 372 759
rect 510 759 516 760
rect 510 758 511 759
rect 366 754 372 755
rect 439 756 511 758
rect 439 754 441 756
rect 510 755 511 756
rect 515 755 516 759
rect 510 754 516 755
rect 570 755 576 756
rect 293 752 321 754
rect 421 752 441 754
rect 214 750 220 751
rect 570 751 571 755
rect 575 754 576 755
rect 938 755 944 756
rect 938 754 939 755
rect 575 752 673 754
rect 861 752 939 754
rect 575 751 576 752
rect 570 750 576 751
rect 938 751 939 752
rect 943 751 944 755
rect 938 750 944 751
rect 946 755 952 756
rect 946 751 947 755
rect 951 754 952 755
rect 951 752 985 754
rect 951 751 952 752
rect 946 750 952 751
rect 1110 751 1116 752
rect 110 746 116 747
rect 1110 747 1111 751
rect 1115 747 1116 751
rect 1110 746 1116 747
rect 142 739 148 740
rect 142 735 143 739
rect 147 735 148 739
rect 142 734 148 735
rect 238 739 244 740
rect 238 735 239 739
rect 243 735 244 739
rect 238 734 244 735
rect 366 739 372 740
rect 366 735 367 739
rect 371 735 372 739
rect 366 734 372 735
rect 510 739 516 740
rect 510 735 511 739
rect 515 735 516 739
rect 510 734 516 735
rect 654 739 660 740
rect 654 735 655 739
rect 659 735 660 739
rect 654 734 660 735
rect 806 739 812 740
rect 806 735 807 739
rect 811 735 812 739
rect 806 734 812 735
rect 966 739 972 740
rect 966 735 967 739
rect 971 735 972 739
rect 966 734 972 735
rect 252 732 270 734
rect 376 732 398 734
rect 664 732 686 734
rect 170 731 176 732
rect 170 727 171 731
rect 175 727 176 731
rect 170 726 176 727
rect 214 723 220 724
rect 214 719 215 723
rect 219 722 220 723
rect 252 722 254 732
rect 268 729 270 732
rect 374 731 380 732
rect 374 727 375 731
rect 379 727 380 731
rect 396 729 398 732
rect 426 731 432 732
rect 374 726 380 727
rect 426 727 427 731
rect 431 730 432 731
rect 558 731 564 732
rect 431 728 494 730
rect 431 727 432 728
rect 426 726 432 727
rect 219 720 254 722
rect 290 723 296 724
rect 492 723 494 728
rect 558 727 559 731
rect 563 730 564 731
rect 662 731 668 732
rect 563 728 606 730
rect 563 727 564 728
rect 558 726 564 727
rect 518 723 524 724
rect 219 719 220 720
rect 214 718 220 719
rect 290 719 291 723
rect 295 719 296 723
rect 290 718 296 719
rect 386 721 392 722
rect 386 717 387 721
rect 391 717 392 721
rect 518 719 519 723
rect 523 722 524 723
rect 540 722 542 725
rect 604 723 606 728
rect 662 727 663 731
rect 667 727 668 731
rect 684 729 686 732
rect 994 731 1000 732
rect 662 726 668 727
rect 858 727 864 728
rect 858 726 859 727
rect 837 724 859 726
rect 714 723 720 724
rect 523 720 542 722
rect 523 719 524 720
rect 518 718 524 719
rect 714 719 715 723
rect 719 719 720 723
rect 858 723 859 724
rect 863 723 864 727
rect 994 727 995 731
rect 999 727 1000 731
rect 994 726 1000 727
rect 1014 731 1020 732
rect 1014 727 1015 731
rect 1019 730 1020 731
rect 1019 728 1054 730
rect 1019 727 1020 728
rect 1014 726 1020 727
rect 858 722 864 723
rect 946 723 952 724
rect 1052 723 1054 728
rect 714 718 720 719
rect 826 721 832 722
rect 386 716 392 717
rect 826 717 827 721
rect 831 717 832 721
rect 946 719 947 723
rect 951 719 952 723
rect 946 718 952 719
rect 826 716 832 717
rect 262 713 268 714
rect 262 709 263 713
rect 267 709 268 713
rect 262 708 268 709
rect 358 713 364 714
rect 358 709 359 713
rect 363 709 364 713
rect 358 708 364 709
rect 462 713 468 714
rect 462 709 463 713
rect 467 709 468 713
rect 462 708 468 709
rect 574 713 580 714
rect 574 709 575 713
rect 579 709 580 713
rect 574 708 580 709
rect 686 713 692 714
rect 686 709 687 713
rect 691 709 692 713
rect 686 708 692 709
rect 798 713 804 714
rect 798 709 799 713
rect 803 709 804 713
rect 798 708 804 709
rect 918 713 924 714
rect 918 709 919 713
rect 923 709 924 713
rect 918 708 924 709
rect 1022 713 1028 714
rect 1022 709 1023 713
rect 1027 709 1028 713
rect 1022 708 1028 709
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 1110 701 1116 702
rect 326 699 332 700
rect 326 698 327 699
rect 110 696 116 697
rect 317 696 327 698
rect 326 695 327 696
rect 331 695 332 699
rect 426 699 432 700
rect 426 698 427 699
rect 413 696 427 698
rect 326 694 332 695
rect 426 695 427 696
rect 431 695 432 699
rect 558 699 564 700
rect 558 698 559 699
rect 517 696 559 698
rect 426 694 432 695
rect 558 695 559 696
rect 563 695 564 699
rect 858 699 864 700
rect 858 698 859 699
rect 853 696 859 698
rect 558 694 564 695
rect 682 695 688 696
rect 682 694 683 695
rect 629 692 683 694
rect 682 691 683 692
rect 687 691 688 695
rect 858 695 859 696
rect 863 695 864 699
rect 1110 697 1111 701
rect 1115 697 1116 701
rect 1110 696 1116 697
rect 858 694 864 695
rect 1014 695 1020 696
rect 1014 694 1015 695
rect 973 692 1015 694
rect 682 690 688 691
rect 1014 691 1015 692
rect 1019 691 1020 695
rect 1014 690 1020 691
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 110 678 116 679
rect 642 683 648 684
rect 642 679 643 683
rect 647 682 648 683
rect 1022 683 1028 684
rect 647 680 697 682
rect 647 679 648 680
rect 642 678 648 679
rect 1022 679 1023 683
rect 1027 682 1028 683
rect 1110 683 1116 684
rect 1027 680 1033 682
rect 1027 679 1028 680
rect 1022 678 1028 679
rect 1110 679 1111 683
rect 1115 679 1116 683
rect 1110 678 1116 679
rect 254 668 260 669
rect 254 664 255 668
rect 259 664 260 668
rect 254 663 260 664
rect 350 668 356 669
rect 350 664 351 668
rect 355 664 356 668
rect 350 663 356 664
rect 454 668 460 669
rect 454 664 455 668
rect 459 664 460 668
rect 454 663 460 664
rect 566 668 572 669
rect 566 664 567 668
rect 571 664 572 668
rect 566 663 572 664
rect 678 668 684 669
rect 678 664 679 668
rect 683 664 684 668
rect 678 663 684 664
rect 790 668 796 669
rect 790 664 791 668
rect 795 664 796 668
rect 790 663 796 664
rect 910 668 916 669
rect 910 664 911 668
rect 915 664 916 668
rect 910 663 916 664
rect 1014 668 1020 669
rect 1014 664 1015 668
rect 1019 664 1020 668
rect 1014 663 1020 664
rect 1022 659 1028 660
rect 506 655 512 656
rect 506 651 507 655
rect 511 654 512 655
rect 642 655 648 656
rect 642 654 643 655
rect 511 652 643 654
rect 511 651 512 652
rect 506 650 512 651
rect 642 651 643 652
rect 647 651 648 655
rect 1022 655 1023 659
rect 1027 658 1028 659
rect 1050 659 1056 660
rect 1050 658 1051 659
rect 1027 656 1051 658
rect 1027 655 1028 656
rect 1022 654 1028 655
rect 1050 655 1051 656
rect 1055 655 1056 659
rect 1050 654 1056 655
rect 642 650 648 651
rect 826 651 832 652
rect 470 648 476 649
rect 470 644 471 648
rect 475 644 476 648
rect 470 643 476 644
rect 566 648 572 649
rect 566 644 567 648
rect 571 644 572 648
rect 566 643 572 644
rect 670 648 676 649
rect 670 644 671 648
rect 675 644 676 648
rect 670 643 676 644
rect 782 648 788 649
rect 782 644 783 648
rect 787 644 788 648
rect 826 647 827 651
rect 831 650 832 651
rect 831 648 878 650
rect 831 647 832 648
rect 826 646 832 647
rect 782 643 788 644
rect 876 634 878 648
rect 902 648 908 649
rect 902 644 903 648
rect 907 644 908 648
rect 902 643 908 644
rect 1014 648 1020 649
rect 1014 644 1015 648
rect 1019 644 1020 648
rect 1014 643 1020 644
rect 110 633 116 634
rect 110 629 111 633
rect 115 629 116 633
rect 729 632 794 634
rect 876 632 921 634
rect 1110 633 1116 634
rect 110 628 116 629
rect 790 631 796 632
rect 790 627 791 631
rect 795 627 796 631
rect 1110 629 1111 633
rect 1115 629 1116 633
rect 1110 628 1116 629
rect 790 626 796 627
rect 574 623 580 624
rect 574 619 575 623
rect 579 619 580 623
rect 574 618 580 619
rect 678 623 684 624
rect 678 619 679 623
rect 683 619 684 623
rect 678 618 684 619
rect 775 619 781 620
rect 533 616 578 618
rect 629 616 681 618
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 775 615 776 619
rect 780 618 781 619
rect 1082 619 1088 620
rect 1082 618 1083 619
rect 780 616 809 618
rect 1077 616 1083 618
rect 780 615 781 616
rect 775 614 781 615
rect 1082 615 1083 616
rect 1087 615 1088 619
rect 1082 614 1088 615
rect 1110 615 1116 616
rect 110 610 116 611
rect 1110 611 1111 615
rect 1115 611 1116 615
rect 1110 610 1116 611
rect 478 603 484 604
rect 478 599 479 603
rect 483 599 484 603
rect 478 598 484 599
rect 574 603 580 604
rect 574 599 575 603
rect 579 599 580 603
rect 574 598 580 599
rect 678 603 684 604
rect 678 599 679 603
rect 683 599 684 603
rect 678 598 684 599
rect 790 603 796 604
rect 790 599 791 603
rect 795 599 796 603
rect 790 598 796 599
rect 910 603 916 604
rect 910 599 911 603
rect 915 599 916 603
rect 910 598 916 599
rect 1022 603 1028 604
rect 1022 599 1023 603
rect 1027 599 1028 603
rect 1022 598 1028 599
rect 584 596 606 598
rect 688 596 710 598
rect 920 596 942 598
rect 506 595 512 596
rect 506 591 507 595
rect 511 591 512 595
rect 506 590 512 591
rect 582 595 588 596
rect 582 591 583 595
rect 587 591 588 595
rect 604 593 606 596
rect 686 595 692 596
rect 582 590 588 591
rect 686 591 687 595
rect 691 591 692 595
rect 708 593 710 596
rect 775 595 781 596
rect 686 590 692 591
rect 775 591 776 595
rect 780 594 781 595
rect 911 595 917 596
rect 780 592 794 594
rect 780 591 781 592
rect 775 590 781 591
rect 554 587 560 588
rect 554 586 555 587
rect 532 584 555 586
rect 528 582 534 584
rect 554 583 555 584
rect 559 583 560 587
rect 650 587 656 588
rect 650 586 651 587
rect 620 584 651 586
rect 554 582 560 583
rect 616 582 622 584
rect 650 583 651 584
rect 655 583 656 587
rect 738 587 744 588
rect 738 586 739 587
rect 708 584 739 586
rect 650 582 656 583
rect 704 582 710 584
rect 738 583 739 584
rect 743 583 744 587
rect 738 582 744 583
rect 792 582 794 592
rect 911 591 912 595
rect 916 594 917 595
rect 920 594 922 596
rect 916 592 922 594
rect 940 593 942 596
rect 1050 595 1056 596
rect 916 591 917 592
rect 911 590 917 591
rect 1050 591 1051 595
rect 1055 591 1056 595
rect 1050 590 1056 591
rect 798 587 804 588
rect 798 583 799 587
rect 803 586 804 587
rect 820 586 822 589
rect 1002 587 1008 588
rect 1002 586 1003 587
rect 803 584 822 586
rect 972 584 1003 586
rect 803 583 804 584
rect 798 582 804 583
rect 874 583 880 584
rect 525 580 530 582
rect 613 580 618 582
rect 701 580 706 582
rect 789 580 794 582
rect 874 579 875 583
rect 879 579 880 583
rect 968 582 974 584
rect 1002 583 1003 584
rect 1007 583 1008 587
rect 1082 587 1088 588
rect 1082 586 1083 587
rect 1060 584 1083 586
rect 1002 582 1008 583
rect 1056 582 1062 584
rect 1082 583 1083 584
rect 1087 583 1088 587
rect 1082 582 1088 583
rect 965 580 970 582
rect 1053 580 1058 582
rect 874 578 880 579
rect 494 573 500 574
rect 494 569 495 573
rect 499 569 500 573
rect 494 568 500 569
rect 582 573 588 574
rect 582 569 583 573
rect 587 569 588 573
rect 582 568 588 569
rect 670 573 676 574
rect 670 569 671 573
rect 675 569 676 573
rect 670 568 676 569
rect 758 573 764 574
rect 758 569 759 573
rect 763 569 764 573
rect 758 568 764 569
rect 846 573 852 574
rect 846 569 847 573
rect 851 569 852 573
rect 846 568 852 569
rect 934 573 940 574
rect 934 569 935 573
rect 939 569 940 573
rect 934 568 940 569
rect 1022 573 1028 574
rect 1022 569 1023 573
rect 1027 569 1028 573
rect 1022 568 1028 569
rect 110 561 116 562
rect 110 557 111 561
rect 115 557 116 561
rect 1110 561 1116 562
rect 110 556 116 557
rect 554 559 560 560
rect 554 555 555 559
rect 559 555 560 559
rect 911 559 917 560
rect 911 558 912 559
rect 901 556 912 558
rect 554 554 560 555
rect 650 555 656 556
rect 556 552 601 554
rect 650 551 651 555
rect 655 554 656 555
rect 738 555 744 556
rect 655 552 689 554
rect 655 551 656 552
rect 650 550 656 551
rect 738 551 739 555
rect 743 554 744 555
rect 911 555 912 556
rect 916 555 917 559
rect 1110 557 1111 561
rect 1115 557 1116 561
rect 1110 556 1116 557
rect 911 554 917 555
rect 1002 555 1008 556
rect 743 552 777 554
rect 743 551 744 552
rect 738 550 744 551
rect 1002 551 1003 555
rect 1007 554 1008 555
rect 1007 552 1041 554
rect 1007 551 1008 552
rect 1002 550 1008 551
rect 110 543 116 544
rect 110 539 111 543
rect 115 539 116 543
rect 567 543 573 544
rect 567 542 568 543
rect 545 540 568 542
rect 110 538 116 539
rect 567 539 568 540
rect 572 539 573 543
rect 1022 543 1028 544
rect 1022 542 1023 543
rect 985 540 1023 542
rect 567 538 573 539
rect 1022 539 1023 540
rect 1027 539 1028 543
rect 1022 538 1028 539
rect 1110 543 1116 544
rect 1110 539 1111 543
rect 1115 539 1116 543
rect 1110 538 1116 539
rect 486 528 492 529
rect 486 524 487 528
rect 491 524 492 528
rect 486 523 492 524
rect 574 528 580 529
rect 574 524 575 528
rect 579 524 580 528
rect 574 523 580 524
rect 662 528 668 529
rect 662 524 663 528
rect 667 524 668 528
rect 662 523 668 524
rect 750 528 756 529
rect 750 524 751 528
rect 755 524 756 528
rect 750 523 756 524
rect 838 528 844 529
rect 926 528 932 529
rect 838 524 839 528
rect 843 524 844 528
rect 838 523 844 524
rect 854 527 860 528
rect 854 523 855 527
rect 859 526 860 527
rect 874 527 880 528
rect 874 526 875 527
rect 859 524 875 526
rect 859 523 860 524
rect 854 522 860 523
rect 874 523 875 524
rect 879 523 880 527
rect 926 524 927 528
rect 931 524 932 528
rect 926 523 932 524
rect 1014 528 1020 529
rect 1014 524 1015 528
rect 1019 524 1020 528
rect 1014 523 1020 524
rect 874 522 880 523
rect 374 512 380 513
rect 374 508 375 512
rect 379 508 380 512
rect 374 507 380 508
rect 486 512 492 513
rect 486 508 487 512
rect 491 508 492 512
rect 486 507 492 508
rect 598 512 604 513
rect 598 508 599 512
rect 603 508 604 512
rect 598 507 604 508
rect 718 512 724 513
rect 718 508 719 512
rect 723 508 724 512
rect 718 507 724 508
rect 846 512 852 513
rect 846 508 847 512
rect 851 508 852 512
rect 846 507 852 508
rect 982 512 988 513
rect 982 508 983 512
rect 987 508 988 512
rect 982 507 988 508
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 856 496 865 498
rect 1110 497 1116 498
rect 110 492 116 493
rect 854 495 860 496
rect 726 491 732 492
rect 726 490 727 491
rect 679 488 727 490
rect 479 483 485 484
rect 479 482 480 483
rect 437 480 480 482
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 479 479 480 480
rect 484 479 485 483
rect 554 483 560 484
rect 554 482 555 483
rect 549 480 555 482
rect 479 478 485 479
rect 554 479 555 480
rect 559 479 560 483
rect 679 482 681 488
rect 726 487 727 488
rect 731 487 732 491
rect 854 491 855 495
rect 859 491 860 495
rect 1110 493 1111 497
rect 1115 493 1116 497
rect 1110 492 1116 493
rect 854 490 860 491
rect 726 486 732 487
rect 661 480 681 482
rect 710 483 716 484
rect 554 478 560 479
rect 710 479 711 483
rect 715 482 716 483
rect 1050 483 1056 484
rect 1050 482 1051 483
rect 715 480 745 482
rect 1045 480 1051 482
rect 715 479 716 480
rect 710 478 716 479
rect 1050 479 1051 480
rect 1055 479 1056 483
rect 1050 478 1056 479
rect 1110 479 1116 480
rect 110 474 116 475
rect 1110 475 1111 479
rect 1115 475 1116 479
rect 1110 474 1116 475
rect 382 467 388 468
rect 382 463 383 467
rect 387 463 388 467
rect 382 462 388 463
rect 494 467 500 468
rect 494 463 495 467
rect 499 463 500 467
rect 494 462 500 463
rect 606 467 612 468
rect 606 463 607 467
rect 611 463 612 467
rect 606 462 612 463
rect 726 467 732 468
rect 726 463 727 467
rect 731 463 732 467
rect 726 462 732 463
rect 854 467 860 468
rect 854 463 855 467
rect 859 463 860 467
rect 854 462 860 463
rect 990 467 996 468
rect 990 463 991 467
rect 995 463 996 467
rect 990 462 996 463
rect 736 460 758 462
rect 410 459 416 460
rect 410 455 411 459
rect 415 455 416 459
rect 410 454 416 455
rect 734 459 740 460
rect 734 455 735 459
rect 739 455 740 459
rect 756 457 758 460
rect 1018 459 1024 460
rect 734 454 740 455
rect 1018 455 1019 459
rect 1023 455 1024 459
rect 1018 454 1024 455
rect 367 451 373 452
rect 358 447 364 448
rect 358 446 359 447
rect 300 444 359 446
rect 296 442 302 444
rect 358 443 359 444
rect 363 443 364 447
rect 367 447 368 451
rect 372 450 373 451
rect 479 451 485 452
rect 372 448 422 450
rect 372 447 373 448
rect 367 446 373 447
rect 420 443 422 448
rect 479 447 480 451
rect 484 450 485 451
rect 524 450 526 453
rect 484 448 526 450
rect 567 451 573 452
rect 484 447 485 448
rect 479 446 485 447
rect 554 447 560 448
rect 554 446 555 447
rect 548 444 555 446
rect 358 442 364 443
rect 544 442 550 444
rect 554 443 555 444
rect 559 443 560 447
rect 567 447 568 451
rect 572 450 573 451
rect 636 450 638 453
rect 572 448 638 450
rect 727 451 733 452
rect 572 447 573 448
rect 567 446 573 447
rect 727 447 728 451
rect 732 450 733 451
rect 818 451 824 452
rect 732 448 782 450
rect 732 447 733 448
rect 727 446 733 447
rect 554 442 560 443
rect 658 443 664 444
rect 780 443 782 448
rect 818 447 819 451
rect 823 450 824 451
rect 884 450 886 453
rect 823 448 886 450
rect 823 447 824 448
rect 818 446 824 447
rect 959 447 965 448
rect 959 446 960 447
rect 916 444 960 446
rect 293 440 298 442
rect 541 440 546 442
rect 658 439 659 443
rect 663 439 664 443
rect 912 442 918 444
rect 959 443 960 444
rect 964 443 965 447
rect 1050 447 1056 448
rect 1050 446 1051 447
rect 1044 444 1051 446
rect 959 442 965 443
rect 1040 442 1046 444
rect 1050 443 1051 444
rect 1055 443 1056 447
rect 1050 442 1056 443
rect 909 440 914 442
rect 1037 440 1042 442
rect 658 438 664 439
rect 262 433 268 434
rect 262 429 263 433
rect 267 429 268 433
rect 262 428 268 429
rect 390 433 396 434
rect 390 429 391 433
rect 395 429 396 433
rect 390 428 396 429
rect 510 433 516 434
rect 510 429 511 433
rect 515 429 516 433
rect 510 428 516 429
rect 630 433 636 434
rect 630 429 631 433
rect 635 429 636 433
rect 630 428 636 429
rect 750 433 756 434
rect 750 429 751 433
rect 755 429 756 433
rect 750 428 756 429
rect 878 433 884 434
rect 878 429 879 433
rect 883 429 884 433
rect 878 428 884 429
rect 1006 433 1012 434
rect 1006 429 1007 433
rect 1011 429 1012 433
rect 1006 428 1012 429
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 1110 421 1116 422
rect 367 419 373 420
rect 367 418 368 419
rect 110 416 116 417
rect 317 416 368 418
rect 367 415 368 416
rect 372 415 373 419
rect 727 419 733 420
rect 727 418 728 419
rect 685 416 728 418
rect 367 414 373 415
rect 458 415 464 416
rect 458 411 459 415
rect 463 414 464 415
rect 727 415 728 416
rect 732 415 733 419
rect 818 419 824 420
rect 818 418 819 419
rect 805 416 819 418
rect 727 414 733 415
rect 818 415 819 416
rect 823 415 824 419
rect 1110 417 1111 421
rect 1115 417 1116 421
rect 1110 416 1116 417
rect 818 414 824 415
rect 959 415 965 416
rect 463 412 529 414
rect 463 411 464 412
rect 458 410 464 411
rect 959 411 960 415
rect 964 414 965 415
rect 964 412 1025 414
rect 964 411 965 412
rect 959 410 965 411
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 970 403 976 404
rect 970 402 971 403
rect 441 400 454 402
rect 929 400 971 402
rect 110 398 116 399
rect 450 399 456 400
rect 450 395 451 399
rect 455 395 456 399
rect 970 399 971 400
rect 975 399 976 403
rect 970 398 976 399
rect 1110 403 1116 404
rect 1110 399 1111 403
rect 1115 399 1116 403
rect 1110 398 1116 399
rect 450 394 456 395
rect 254 388 260 389
rect 254 384 255 388
rect 259 384 260 388
rect 254 383 260 384
rect 382 388 388 389
rect 382 384 383 388
rect 387 384 388 388
rect 382 383 388 384
rect 502 388 508 389
rect 502 384 503 388
rect 507 384 508 388
rect 502 383 508 384
rect 622 388 628 389
rect 622 384 623 388
rect 627 384 628 388
rect 622 383 628 384
rect 742 388 748 389
rect 742 384 743 388
rect 747 384 748 388
rect 742 383 748 384
rect 870 388 876 389
rect 870 384 871 388
rect 875 384 876 388
rect 870 383 876 384
rect 998 388 1004 389
rect 998 384 999 388
rect 1003 384 1004 388
rect 998 383 1004 384
rect 134 372 140 373
rect 134 368 135 372
rect 139 368 140 372
rect 134 367 140 368
rect 254 372 260 373
rect 254 368 255 372
rect 259 368 260 372
rect 254 367 260 368
rect 414 372 420 373
rect 414 368 415 372
rect 419 368 420 372
rect 414 367 420 368
rect 582 372 588 373
rect 582 368 583 372
rect 587 368 588 372
rect 582 367 588 368
rect 758 372 764 373
rect 758 368 759 372
rect 763 368 764 372
rect 758 367 764 368
rect 934 372 940 373
rect 934 368 935 372
rect 939 368 940 372
rect 934 367 940 368
rect 658 359 664 360
rect 110 357 116 358
rect 110 353 111 357
rect 115 353 116 357
rect 658 355 659 359
rect 663 358 664 359
rect 663 356 777 358
rect 1110 357 1116 358
rect 663 355 664 356
rect 658 354 664 355
rect 110 352 116 353
rect 1110 353 1111 357
rect 1115 353 1116 357
rect 1110 352 1116 353
rect 202 343 208 344
rect 202 342 203 343
rect 197 340 203 342
rect 110 339 116 340
rect 110 335 111 339
rect 115 335 116 339
rect 202 339 203 340
rect 207 339 208 343
rect 202 338 208 339
rect 223 343 229 344
rect 223 339 224 343
rect 228 342 229 343
rect 490 343 496 344
rect 490 342 491 343
rect 228 340 281 342
rect 477 340 491 342
rect 228 339 229 340
rect 223 338 229 339
rect 490 339 491 340
rect 495 339 496 343
rect 490 338 496 339
rect 498 343 504 344
rect 498 339 499 343
rect 503 342 504 343
rect 898 343 904 344
rect 503 340 609 342
rect 503 339 504 340
rect 498 338 504 339
rect 898 339 899 343
rect 903 342 904 343
rect 903 340 961 342
rect 903 339 904 340
rect 898 338 904 339
rect 1110 339 1116 340
rect 110 334 116 335
rect 1110 335 1111 339
rect 1115 335 1116 339
rect 1110 334 1116 335
rect 142 327 148 328
rect 142 323 143 327
rect 147 323 148 327
rect 142 322 148 323
rect 262 327 268 328
rect 262 323 263 327
rect 267 323 268 327
rect 262 322 268 323
rect 422 327 428 328
rect 422 323 423 327
rect 427 323 428 327
rect 422 322 428 323
rect 590 327 596 328
rect 590 323 591 327
rect 595 323 596 327
rect 590 322 596 323
rect 766 327 772 328
rect 766 323 767 327
rect 771 323 772 327
rect 766 322 772 323
rect 942 327 948 328
rect 942 323 943 327
rect 947 323 948 327
rect 942 322 948 323
rect 290 319 296 320
rect 223 315 229 316
rect 223 314 224 315
rect 173 312 224 314
rect 223 311 224 312
rect 228 311 229 315
rect 290 315 291 319
rect 295 315 296 319
rect 290 314 296 315
rect 450 319 456 320
rect 450 315 451 319
rect 455 315 456 319
rect 450 314 456 315
rect 618 319 624 320
rect 618 315 619 319
rect 623 315 624 319
rect 794 319 800 320
rect 618 314 624 315
rect 638 315 644 316
rect 223 310 229 311
rect 638 311 639 315
rect 643 314 644 315
rect 794 315 795 319
rect 799 315 800 319
rect 794 314 800 315
rect 970 319 976 320
rect 970 315 971 319
rect 975 315 976 319
rect 970 314 976 315
rect 990 315 996 316
rect 643 312 750 314
rect 643 311 644 312
rect 638 310 644 311
rect 180 308 206 310
rect 176 306 182 308
rect 202 307 208 308
rect 173 304 178 306
rect 202 303 203 307
rect 207 303 208 307
rect 202 302 208 303
rect 298 307 304 308
rect 298 303 299 307
rect 303 303 304 307
rect 298 302 304 303
rect 450 307 456 308
rect 450 303 451 307
rect 455 303 456 307
rect 450 302 456 303
rect 602 307 608 308
rect 748 307 750 312
rect 990 311 991 315
rect 995 314 996 315
rect 995 312 1054 314
rect 995 311 996 312
rect 990 310 996 311
rect 898 307 904 308
rect 1052 307 1054 312
rect 602 303 603 307
rect 607 303 608 307
rect 602 302 608 303
rect 898 303 899 307
rect 903 303 904 307
rect 898 302 904 303
rect 142 297 148 298
rect 142 293 143 297
rect 147 293 148 297
rect 142 292 148 293
rect 270 297 276 298
rect 270 293 271 297
rect 275 293 276 297
rect 270 292 276 293
rect 422 297 428 298
rect 422 293 423 297
rect 427 293 428 297
rect 422 292 428 293
rect 574 297 580 298
rect 574 293 575 297
rect 579 293 580 297
rect 574 292 580 293
rect 718 297 724 298
rect 718 293 719 297
rect 723 293 724 297
rect 718 292 724 293
rect 870 297 876 298
rect 870 293 871 297
rect 875 293 876 297
rect 870 292 876 293
rect 1022 297 1028 298
rect 1022 293 1023 297
rect 1027 293 1028 297
rect 1022 292 1028 293
rect 110 285 116 286
rect 110 281 111 285
rect 115 281 116 285
rect 1110 285 1116 286
rect 222 283 228 284
rect 222 282 223 283
rect 110 280 116 281
rect 197 280 223 282
rect 222 279 223 280
rect 227 279 228 283
rect 382 283 388 284
rect 382 282 383 283
rect 325 280 383 282
rect 222 278 228 279
rect 382 279 383 280
rect 387 279 388 283
rect 638 283 644 284
rect 638 282 639 283
rect 629 280 639 282
rect 382 278 388 279
rect 638 279 639 280
rect 643 279 644 283
rect 794 283 800 284
rect 794 282 795 283
rect 773 280 795 282
rect 638 278 644 279
rect 794 279 795 280
rect 799 279 800 283
rect 990 283 996 284
rect 990 282 991 283
rect 925 280 991 282
rect 794 278 800 279
rect 990 279 991 280
rect 995 279 996 283
rect 1110 281 1111 285
rect 1115 281 1116 285
rect 1110 280 1116 281
rect 990 278 996 279
rect 110 267 116 268
rect 110 263 111 267
rect 115 263 116 267
rect 522 267 528 268
rect 522 266 523 267
rect 473 264 523 266
rect 110 262 116 263
rect 522 263 523 264
rect 527 263 528 267
rect 522 262 528 263
rect 1022 267 1028 268
rect 1022 263 1023 267
rect 1027 266 1028 267
rect 1110 267 1116 268
rect 1027 264 1033 266
rect 1027 263 1028 264
rect 1022 262 1028 263
rect 1110 263 1111 267
rect 1115 263 1116 267
rect 1110 262 1116 263
rect 134 252 140 253
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 262 252 268 253
rect 262 248 263 252
rect 267 248 268 252
rect 262 247 268 248
rect 414 252 420 253
rect 414 248 415 252
rect 419 248 420 252
rect 414 247 420 248
rect 566 252 572 253
rect 566 248 567 252
rect 571 248 572 252
rect 566 247 572 248
rect 710 252 716 253
rect 710 248 711 252
rect 715 248 716 252
rect 710 247 716 248
rect 862 252 868 253
rect 862 248 863 252
rect 867 248 868 252
rect 862 247 868 248
rect 1014 252 1020 253
rect 1014 248 1015 252
rect 1019 248 1020 252
rect 1014 247 1020 248
rect 174 236 180 237
rect 174 232 175 236
rect 179 232 180 236
rect 174 231 180 232
rect 326 236 332 237
rect 326 232 327 236
rect 331 232 332 236
rect 326 231 332 232
rect 486 236 492 237
rect 486 232 487 236
rect 491 232 492 236
rect 486 231 492 232
rect 654 236 660 237
rect 654 232 655 236
rect 659 232 660 236
rect 654 231 660 232
rect 830 236 836 237
rect 830 232 831 236
rect 835 232 836 236
rect 830 231 836 232
rect 1006 236 1012 237
rect 1006 232 1007 236
rect 1011 232 1012 236
rect 1006 231 1012 232
rect 602 223 608 224
rect 110 221 116 222
rect 110 217 111 221
rect 115 217 116 221
rect 602 219 603 223
rect 607 222 608 223
rect 607 220 673 222
rect 1110 221 1116 222
rect 607 219 608 220
rect 602 218 608 219
rect 110 216 116 217
rect 1110 217 1111 221
rect 1115 217 1116 221
rect 1110 216 1116 217
rect 170 211 176 212
rect 170 207 171 211
rect 175 207 176 211
rect 170 206 176 207
rect 263 207 269 208
rect 172 204 201 206
rect 110 203 116 204
rect 110 199 111 203
rect 115 199 116 203
rect 263 203 264 207
rect 268 206 269 207
rect 434 207 440 208
rect 268 204 353 206
rect 268 203 269 204
rect 263 202 269 203
rect 434 203 435 207
rect 439 206 440 207
rect 770 207 776 208
rect 439 204 513 206
rect 439 203 440 204
rect 434 202 440 203
rect 770 203 771 207
rect 775 206 776 207
rect 1074 207 1080 208
rect 1074 206 1075 207
rect 775 204 857 206
rect 1069 204 1075 206
rect 775 203 776 204
rect 770 202 776 203
rect 1074 203 1075 204
rect 1079 203 1080 207
rect 1074 202 1080 203
rect 1110 203 1116 204
rect 110 198 116 199
rect 1110 199 1111 203
rect 1115 199 1116 203
rect 1110 198 1116 199
rect 182 191 188 192
rect 182 187 183 191
rect 187 187 188 191
rect 182 186 188 187
rect 334 191 340 192
rect 334 187 335 191
rect 339 187 340 191
rect 334 186 340 187
rect 494 191 500 192
rect 494 187 495 191
rect 499 187 500 191
rect 494 186 500 187
rect 662 191 668 192
rect 662 187 663 191
rect 667 187 668 191
rect 662 186 668 187
rect 838 191 844 192
rect 838 187 839 191
rect 843 187 844 191
rect 838 186 844 187
rect 1014 191 1020 192
rect 1014 187 1015 191
rect 1019 187 1020 191
rect 1014 186 1020 187
rect 522 183 528 184
rect 263 179 269 180
rect 263 178 264 179
rect 213 176 264 178
rect 263 175 264 176
rect 268 175 269 179
rect 434 179 440 180
rect 434 178 435 179
rect 365 176 435 178
rect 263 174 269 175
rect 434 175 435 176
rect 439 175 440 179
rect 522 179 523 183
rect 527 179 528 183
rect 522 178 528 179
rect 770 179 776 180
rect 770 178 771 179
rect 693 176 771 178
rect 434 174 440 175
rect 770 175 771 176
rect 775 175 776 179
rect 770 174 776 175
rect 818 175 824 176
rect 818 171 819 175
rect 823 174 824 175
rect 868 174 870 177
rect 823 172 870 174
rect 1022 175 1028 176
rect 823 171 824 172
rect 818 170 824 171
rect 1022 171 1023 175
rect 1027 174 1028 175
rect 1044 174 1046 177
rect 1027 172 1046 174
rect 1027 171 1028 172
rect 1022 170 1028 171
rect 202 167 208 168
rect 202 163 203 167
rect 207 166 208 167
rect 290 167 296 168
rect 207 164 262 166
rect 207 163 208 164
rect 202 162 208 163
rect 170 159 176 160
rect 260 159 262 164
rect 290 163 291 167
rect 295 166 296 167
rect 378 167 384 168
rect 295 164 350 166
rect 295 163 296 164
rect 290 162 296 163
rect 348 159 350 164
rect 378 163 379 167
rect 383 166 384 167
rect 466 167 472 168
rect 383 164 438 166
rect 383 163 384 164
rect 378 162 384 163
rect 436 159 438 164
rect 466 163 467 167
rect 471 166 472 167
rect 554 167 560 168
rect 471 164 526 166
rect 471 163 472 164
rect 466 162 472 163
rect 524 159 526 164
rect 554 163 555 167
rect 559 166 560 167
rect 642 167 648 168
rect 559 164 614 166
rect 559 163 560 164
rect 554 162 560 163
rect 612 159 614 164
rect 642 163 643 167
rect 647 166 648 167
rect 730 167 736 168
rect 647 164 702 166
rect 647 163 648 164
rect 642 162 648 163
rect 700 159 702 164
rect 730 163 731 167
rect 735 166 736 167
rect 735 164 790 166
rect 735 163 736 164
rect 730 162 736 163
rect 788 159 790 164
rect 914 163 920 164
rect 914 162 915 163
rect 884 160 915 162
rect 170 155 171 159
rect 175 155 176 159
rect 880 158 886 160
rect 914 159 915 160
rect 919 159 920 163
rect 1002 163 1008 164
rect 1002 162 1003 163
rect 972 160 1003 162
rect 914 158 920 159
rect 968 158 974 160
rect 1002 159 1003 160
rect 1007 159 1008 163
rect 1074 163 1080 164
rect 1074 162 1075 163
rect 1060 160 1075 162
rect 1002 158 1008 159
rect 1056 158 1062 160
rect 1074 159 1075 160
rect 1079 159 1080 163
rect 1074 158 1080 159
rect 877 156 882 158
rect 965 156 970 158
rect 1053 156 1058 158
rect 170 154 176 155
rect 142 149 148 150
rect 142 145 143 149
rect 147 145 148 149
rect 142 144 148 145
rect 230 149 236 150
rect 230 145 231 149
rect 235 145 236 149
rect 230 144 236 145
rect 318 149 324 150
rect 318 145 319 149
rect 323 145 324 149
rect 318 144 324 145
rect 406 149 412 150
rect 406 145 407 149
rect 411 145 412 149
rect 406 144 412 145
rect 494 149 500 150
rect 494 145 495 149
rect 499 145 500 149
rect 494 144 500 145
rect 582 149 588 150
rect 582 145 583 149
rect 587 145 588 149
rect 582 144 588 145
rect 670 149 676 150
rect 670 145 671 149
rect 675 145 676 149
rect 670 144 676 145
rect 758 149 764 150
rect 758 145 759 149
rect 763 145 764 149
rect 758 144 764 145
rect 846 149 852 150
rect 846 145 847 149
rect 851 145 852 149
rect 846 144 852 145
rect 934 149 940 150
rect 934 145 935 149
rect 939 145 940 149
rect 934 144 940 145
rect 1022 149 1028 150
rect 1022 145 1023 149
rect 1027 145 1028 149
rect 1022 144 1028 145
rect 110 137 116 138
rect 110 133 111 137
rect 115 133 116 137
rect 1110 137 1116 138
rect 202 135 208 136
rect 202 134 203 135
rect 110 132 116 133
rect 197 132 203 134
rect 202 131 203 132
rect 207 131 208 135
rect 290 135 296 136
rect 290 134 291 135
rect 285 132 291 134
rect 202 130 208 131
rect 290 131 291 132
rect 295 131 296 135
rect 378 135 384 136
rect 378 134 379 135
rect 373 132 379 134
rect 290 130 296 131
rect 378 131 379 132
rect 383 131 384 135
rect 466 135 472 136
rect 466 134 467 135
rect 461 132 467 134
rect 378 130 384 131
rect 466 131 467 132
rect 471 131 472 135
rect 554 135 560 136
rect 554 134 555 135
rect 549 132 555 134
rect 466 130 472 131
rect 554 131 555 132
rect 559 131 560 135
rect 642 135 648 136
rect 642 134 643 135
rect 637 132 643 134
rect 554 130 560 131
rect 642 131 643 132
rect 647 131 648 135
rect 730 135 736 136
rect 730 134 731 135
rect 725 132 731 134
rect 642 130 648 131
rect 730 131 731 132
rect 735 131 736 135
rect 818 135 824 136
rect 818 134 819 135
rect 813 132 819 134
rect 730 130 736 131
rect 818 131 819 132
rect 823 131 824 135
rect 1110 133 1111 137
rect 1115 133 1116 137
rect 1110 132 1116 133
rect 818 130 824 131
rect 914 131 920 132
rect 914 127 915 131
rect 919 130 920 131
rect 1002 131 1008 132
rect 919 128 953 130
rect 919 127 920 128
rect 914 126 920 127
rect 1002 127 1003 131
rect 1007 130 1008 131
rect 1007 128 1041 130
rect 1007 127 1008 128
rect 1002 126 1008 127
rect 110 119 116 120
rect 110 115 111 119
rect 115 115 116 119
rect 110 114 116 115
rect 1110 119 1116 120
rect 1110 115 1111 119
rect 1115 115 1116 119
rect 1110 114 1116 115
rect 134 104 140 105
rect 134 100 135 104
rect 139 100 140 104
rect 134 99 140 100
rect 222 104 228 105
rect 222 100 223 104
rect 227 100 228 104
rect 222 99 228 100
rect 310 104 316 105
rect 310 100 311 104
rect 315 100 316 104
rect 310 99 316 100
rect 398 104 404 105
rect 398 100 399 104
rect 403 100 404 104
rect 398 99 404 100
rect 486 104 492 105
rect 486 100 487 104
rect 491 100 492 104
rect 486 99 492 100
rect 574 104 580 105
rect 574 100 575 104
rect 579 100 580 104
rect 574 99 580 100
rect 662 104 668 105
rect 662 100 663 104
rect 667 100 668 104
rect 662 99 668 100
rect 750 104 756 105
rect 750 100 751 104
rect 755 100 756 104
rect 750 99 756 100
rect 838 104 844 105
rect 838 100 839 104
rect 843 100 844 104
rect 838 99 844 100
rect 926 104 932 105
rect 926 100 927 104
rect 931 100 932 104
rect 926 99 932 100
rect 1014 104 1020 105
rect 1014 100 1015 104
rect 1019 100 1020 104
rect 1014 99 1020 100
<< m3c >>
rect 135 1196 139 1200
rect 223 1196 227 1200
rect 311 1196 315 1200
rect 399 1196 403 1200
rect 487 1196 491 1200
rect 575 1196 579 1200
rect 663 1196 667 1200
rect 751 1196 755 1200
rect 111 1181 115 1185
rect 1111 1181 1115 1185
rect 111 1163 115 1167
rect 291 1167 295 1171
rect 1111 1163 1115 1167
rect 143 1151 147 1155
rect 231 1151 235 1155
rect 319 1151 323 1155
rect 407 1151 411 1155
rect 495 1151 499 1155
rect 583 1151 587 1155
rect 671 1151 675 1155
rect 759 1151 763 1155
rect 523 1143 527 1147
rect 291 1135 295 1139
rect 523 1127 527 1131
rect 159 1113 163 1117
rect 247 1113 251 1117
rect 335 1113 339 1117
rect 423 1113 427 1117
rect 111 1101 115 1105
rect 1111 1101 1115 1105
rect 111 1083 115 1087
rect 247 1083 251 1087
rect 1111 1083 1115 1087
rect 151 1068 155 1072
rect 239 1068 243 1072
rect 327 1068 331 1072
rect 415 1068 419 1072
rect 135 1052 139 1056
rect 223 1052 227 1056
rect 311 1052 315 1056
rect 399 1052 403 1056
rect 111 1037 115 1041
rect 379 1039 383 1043
rect 1111 1037 1115 1041
rect 111 1019 115 1023
rect 203 1023 207 1027
rect 319 1027 323 1031
rect 407 1027 411 1031
rect 1111 1019 1115 1023
rect 143 1007 147 1011
rect 231 1007 235 1011
rect 319 1007 323 1011
rect 407 1007 411 1011
rect 171 999 175 1003
rect 259 999 263 1003
rect 327 999 331 1003
rect 415 999 419 1003
rect 203 991 207 995
rect 259 987 263 991
rect 347 987 351 991
rect 435 987 439 991
rect 143 977 147 981
rect 231 977 235 981
rect 319 977 323 981
rect 407 977 411 981
rect 111 965 115 969
rect 1111 965 1115 969
rect 231 959 235 963
rect 319 959 323 963
rect 407 959 411 963
rect 111 947 115 951
rect 467 943 471 947
rect 1111 947 1115 951
rect 135 932 139 936
rect 223 932 227 936
rect 311 932 315 936
rect 399 932 403 936
rect 135 916 139 920
rect 223 916 227 920
rect 311 916 315 920
rect 399 916 403 920
rect 111 901 115 905
rect 1111 901 1115 905
rect 111 883 115 887
rect 207 887 211 891
rect 291 887 295 891
rect 199 879 203 883
rect 1111 883 1115 887
rect 143 871 147 875
rect 231 871 235 875
rect 319 871 323 875
rect 407 871 411 875
rect 207 859 211 863
rect 291 859 295 863
rect 467 859 471 863
rect 199 851 203 855
rect 259 851 263 855
rect 347 851 351 855
rect 435 851 439 855
rect 143 841 147 845
rect 231 841 235 845
rect 319 841 323 845
rect 407 841 411 845
rect 495 841 499 845
rect 111 829 115 833
rect 231 823 235 827
rect 319 823 323 827
rect 407 823 411 827
rect 1111 829 1115 833
rect 111 811 115 815
rect 475 811 479 815
rect 1111 811 1115 815
rect 135 796 139 800
rect 223 796 227 800
rect 311 796 315 800
rect 399 796 403 800
rect 487 796 491 800
rect 135 780 139 784
rect 231 780 235 784
rect 359 780 363 784
rect 503 780 507 784
rect 647 780 651 784
rect 799 780 803 784
rect 959 780 963 784
rect 111 765 115 769
rect 655 763 659 767
rect 1111 765 1115 769
rect 111 747 115 751
rect 215 751 219 755
rect 367 755 371 759
rect 511 755 515 759
rect 571 751 575 755
rect 939 751 943 755
rect 947 751 951 755
rect 1111 747 1115 751
rect 143 735 147 739
rect 239 735 243 739
rect 367 735 371 739
rect 511 735 515 739
rect 655 735 659 739
rect 807 735 811 739
rect 967 735 971 739
rect 171 727 175 731
rect 215 719 219 723
rect 375 727 379 731
rect 427 727 431 731
rect 559 727 563 731
rect 291 719 295 723
rect 387 717 391 721
rect 519 719 523 723
rect 663 727 667 731
rect 715 719 719 723
rect 859 723 863 727
rect 995 727 999 731
rect 1015 727 1019 731
rect 827 717 831 721
rect 947 719 951 723
rect 263 709 267 713
rect 359 709 363 713
rect 463 709 467 713
rect 575 709 579 713
rect 687 709 691 713
rect 799 709 803 713
rect 919 709 923 713
rect 1023 709 1027 713
rect 111 697 115 701
rect 327 695 331 699
rect 427 695 431 699
rect 559 695 563 699
rect 683 691 687 695
rect 859 695 863 699
rect 1111 697 1115 701
rect 1015 691 1019 695
rect 111 679 115 683
rect 643 679 647 683
rect 1023 679 1027 683
rect 1111 679 1115 683
rect 255 664 259 668
rect 351 664 355 668
rect 455 664 459 668
rect 567 664 571 668
rect 679 664 683 668
rect 791 664 795 668
rect 911 664 915 668
rect 1015 664 1019 668
rect 507 651 511 655
rect 643 651 647 655
rect 1023 655 1027 659
rect 1051 655 1055 659
rect 471 644 475 648
rect 567 644 571 648
rect 671 644 675 648
rect 783 644 787 648
rect 827 647 831 651
rect 903 644 907 648
rect 1015 644 1019 648
rect 111 629 115 633
rect 791 627 795 631
rect 1111 629 1115 633
rect 575 619 579 623
rect 679 619 683 623
rect 111 611 115 615
rect 1083 615 1087 619
rect 1111 611 1115 615
rect 479 599 483 603
rect 575 599 579 603
rect 679 599 683 603
rect 791 599 795 603
rect 911 599 915 603
rect 1023 599 1027 603
rect 507 591 511 595
rect 583 591 587 595
rect 687 591 691 595
rect 555 583 559 587
rect 651 583 655 587
rect 739 583 743 587
rect 1051 591 1055 595
rect 799 583 803 587
rect 875 579 879 583
rect 1003 583 1007 587
rect 1083 583 1087 587
rect 495 569 499 573
rect 583 569 587 573
rect 671 569 675 573
rect 759 569 763 573
rect 847 569 851 573
rect 935 569 939 573
rect 1023 569 1027 573
rect 111 557 115 561
rect 555 555 559 559
rect 651 551 655 555
rect 739 551 743 555
rect 1111 557 1115 561
rect 1003 551 1007 555
rect 111 539 115 543
rect 1023 539 1027 543
rect 1111 539 1115 543
rect 487 524 491 528
rect 575 524 579 528
rect 663 524 667 528
rect 751 524 755 528
rect 839 524 843 528
rect 855 523 859 527
rect 875 523 879 527
rect 927 524 931 528
rect 1015 524 1019 528
rect 375 508 379 512
rect 487 508 491 512
rect 599 508 603 512
rect 719 508 723 512
rect 847 508 851 512
rect 983 508 987 512
rect 111 493 115 497
rect 111 475 115 479
rect 555 479 559 483
rect 727 487 731 491
rect 855 491 859 495
rect 1111 493 1115 497
rect 711 479 715 483
rect 1051 479 1055 483
rect 1111 475 1115 479
rect 383 463 387 467
rect 495 463 499 467
rect 607 463 611 467
rect 727 463 731 467
rect 855 463 859 467
rect 991 463 995 467
rect 411 455 415 459
rect 735 455 739 459
rect 1019 455 1023 459
rect 359 443 363 447
rect 555 443 559 447
rect 819 447 823 451
rect 659 439 663 443
rect 1051 443 1055 447
rect 263 429 267 433
rect 391 429 395 433
rect 511 429 515 433
rect 631 429 635 433
rect 751 429 755 433
rect 879 429 883 433
rect 1007 429 1011 433
rect 111 417 115 421
rect 459 411 463 415
rect 819 415 823 419
rect 1111 417 1115 421
rect 111 399 115 403
rect 451 395 455 399
rect 971 399 975 403
rect 1111 399 1115 403
rect 255 384 259 388
rect 383 384 387 388
rect 503 384 507 388
rect 623 384 627 388
rect 743 384 747 388
rect 871 384 875 388
rect 999 384 1003 388
rect 135 368 139 372
rect 255 368 259 372
rect 415 368 419 372
rect 583 368 587 372
rect 759 368 763 372
rect 935 368 939 372
rect 111 353 115 357
rect 659 355 663 359
rect 1111 353 1115 357
rect 111 335 115 339
rect 203 339 207 343
rect 491 339 495 343
rect 499 339 503 343
rect 899 339 903 343
rect 1111 335 1115 339
rect 143 323 147 327
rect 263 323 267 327
rect 423 323 427 327
rect 591 323 595 327
rect 767 323 771 327
rect 943 323 947 327
rect 291 315 295 319
rect 451 315 455 319
rect 619 315 623 319
rect 639 311 643 315
rect 795 315 799 319
rect 971 315 975 319
rect 203 303 207 307
rect 299 303 303 307
rect 451 303 455 307
rect 991 311 995 315
rect 603 303 607 307
rect 899 303 903 307
rect 143 293 147 297
rect 271 293 275 297
rect 423 293 427 297
rect 575 293 579 297
rect 719 293 723 297
rect 871 293 875 297
rect 1023 293 1027 297
rect 111 281 115 285
rect 223 279 227 283
rect 383 279 387 283
rect 639 279 643 283
rect 795 279 799 283
rect 991 279 995 283
rect 1111 281 1115 285
rect 111 263 115 267
rect 523 263 527 267
rect 1023 263 1027 267
rect 1111 263 1115 267
rect 135 248 139 252
rect 263 248 267 252
rect 415 248 419 252
rect 567 248 571 252
rect 711 248 715 252
rect 863 248 867 252
rect 1015 248 1019 252
rect 175 232 179 236
rect 327 232 331 236
rect 487 232 491 236
rect 655 232 659 236
rect 831 232 835 236
rect 1007 232 1011 236
rect 111 217 115 221
rect 603 219 607 223
rect 1111 217 1115 221
rect 171 207 175 211
rect 111 199 115 203
rect 435 203 439 207
rect 771 203 775 207
rect 1075 203 1079 207
rect 1111 199 1115 203
rect 183 187 187 191
rect 335 187 339 191
rect 495 187 499 191
rect 663 187 667 191
rect 839 187 843 191
rect 1015 187 1019 191
rect 435 175 439 179
rect 523 179 527 183
rect 771 175 775 179
rect 819 171 823 175
rect 1023 171 1027 175
rect 203 163 207 167
rect 291 163 295 167
rect 379 163 383 167
rect 467 163 471 167
rect 555 163 559 167
rect 643 163 647 167
rect 731 163 735 167
rect 171 155 175 159
rect 915 159 919 163
rect 1003 159 1007 163
rect 1075 159 1079 163
rect 143 145 147 149
rect 231 145 235 149
rect 319 145 323 149
rect 407 145 411 149
rect 495 145 499 149
rect 583 145 587 149
rect 671 145 675 149
rect 759 145 763 149
rect 847 145 851 149
rect 935 145 939 149
rect 1023 145 1027 149
rect 111 133 115 137
rect 203 131 207 135
rect 291 131 295 135
rect 379 131 383 135
rect 467 131 471 135
rect 555 131 559 135
rect 643 131 647 135
rect 731 131 735 135
rect 819 131 823 135
rect 1111 133 1115 137
rect 915 127 919 131
rect 1003 127 1007 131
rect 111 115 115 119
rect 1111 115 1115 119
rect 135 100 139 104
rect 223 100 227 104
rect 311 100 315 104
rect 399 100 403 104
rect 487 100 491 104
rect 575 100 579 104
rect 663 100 667 104
rect 751 100 755 104
rect 839 100 843 104
rect 927 100 931 104
rect 1015 100 1019 104
<< m3 >>
rect 111 1206 115 1207
rect 111 1201 115 1202
rect 135 1206 139 1207
rect 135 1201 139 1202
rect 223 1206 227 1207
rect 223 1201 227 1202
rect 311 1206 315 1207
rect 311 1201 315 1202
rect 399 1206 403 1207
rect 399 1201 403 1202
rect 487 1206 491 1207
rect 487 1201 491 1202
rect 575 1206 579 1207
rect 575 1201 579 1202
rect 663 1206 667 1207
rect 663 1201 667 1202
rect 751 1206 755 1207
rect 751 1201 755 1202
rect 1111 1206 1115 1207
rect 1111 1201 1115 1202
rect 112 1186 114 1201
rect 134 1200 140 1201
rect 134 1196 135 1200
rect 139 1196 140 1200
rect 134 1195 140 1196
rect 222 1200 228 1201
rect 222 1196 223 1200
rect 227 1196 228 1200
rect 222 1195 228 1196
rect 310 1200 316 1201
rect 310 1196 311 1200
rect 315 1196 316 1200
rect 310 1195 316 1196
rect 398 1200 404 1201
rect 398 1196 399 1200
rect 403 1196 404 1200
rect 398 1195 404 1196
rect 486 1200 492 1201
rect 486 1196 487 1200
rect 491 1196 492 1200
rect 486 1195 492 1196
rect 574 1200 580 1201
rect 574 1196 575 1200
rect 579 1196 580 1200
rect 574 1195 580 1196
rect 662 1200 668 1201
rect 662 1196 663 1200
rect 667 1196 668 1200
rect 662 1195 668 1196
rect 750 1200 756 1201
rect 750 1196 751 1200
rect 755 1196 756 1200
rect 750 1195 756 1196
rect 1112 1186 1114 1201
rect 110 1185 116 1186
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 110 1180 116 1181
rect 1110 1185 1116 1186
rect 1110 1181 1111 1185
rect 1115 1181 1116 1185
rect 1110 1180 1116 1181
rect 290 1171 296 1172
rect 110 1167 116 1168
rect 110 1163 111 1167
rect 115 1163 116 1167
rect 290 1167 291 1171
rect 295 1167 296 1171
rect 290 1166 296 1167
rect 1110 1167 1116 1168
rect 110 1162 116 1163
rect 112 1131 114 1162
rect 142 1155 148 1156
rect 142 1151 143 1155
rect 147 1151 148 1155
rect 142 1150 148 1151
rect 230 1155 236 1156
rect 230 1151 231 1155
rect 235 1151 236 1155
rect 230 1150 236 1151
rect 144 1131 146 1150
rect 232 1131 234 1150
rect 292 1140 294 1166
rect 1110 1163 1111 1167
rect 1115 1163 1116 1167
rect 1110 1162 1116 1163
rect 318 1155 324 1156
rect 318 1151 319 1155
rect 323 1151 324 1155
rect 318 1150 324 1151
rect 406 1155 412 1156
rect 406 1151 407 1155
rect 411 1151 412 1155
rect 406 1150 412 1151
rect 494 1155 500 1156
rect 494 1151 495 1155
rect 499 1151 500 1155
rect 494 1150 500 1151
rect 582 1155 588 1156
rect 582 1151 583 1155
rect 587 1151 588 1155
rect 582 1150 588 1151
rect 670 1155 676 1156
rect 670 1151 671 1155
rect 675 1151 676 1155
rect 670 1150 676 1151
rect 758 1155 764 1156
rect 758 1151 759 1155
rect 763 1151 764 1155
rect 758 1150 764 1151
rect 290 1139 296 1140
rect 290 1135 291 1139
rect 295 1135 296 1139
rect 290 1134 296 1135
rect 320 1131 322 1150
rect 408 1131 410 1150
rect 496 1131 498 1150
rect 522 1147 528 1148
rect 522 1143 523 1147
rect 527 1143 528 1147
rect 522 1142 528 1143
rect 524 1132 526 1142
rect 522 1131 528 1132
rect 584 1131 586 1150
rect 672 1131 674 1150
rect 760 1131 762 1150
rect 1112 1131 1114 1162
rect 111 1130 115 1131
rect 111 1125 115 1126
rect 143 1130 147 1131
rect 143 1125 147 1126
rect 159 1130 163 1131
rect 159 1125 163 1126
rect 231 1130 235 1131
rect 231 1125 235 1126
rect 247 1130 251 1131
rect 247 1125 251 1126
rect 319 1130 323 1131
rect 319 1125 323 1126
rect 335 1130 339 1131
rect 335 1125 339 1126
rect 407 1130 411 1131
rect 407 1125 411 1126
rect 423 1130 427 1131
rect 423 1125 427 1126
rect 495 1130 499 1131
rect 522 1127 523 1131
rect 527 1127 528 1131
rect 522 1126 528 1127
rect 583 1130 587 1131
rect 495 1125 499 1126
rect 583 1125 587 1126
rect 671 1130 675 1131
rect 671 1125 675 1126
rect 759 1130 763 1131
rect 759 1125 763 1126
rect 1111 1130 1115 1131
rect 1111 1125 1115 1126
rect 112 1106 114 1125
rect 160 1118 162 1125
rect 248 1118 250 1125
rect 336 1118 338 1125
rect 424 1118 426 1125
rect 158 1117 164 1118
rect 158 1113 159 1117
rect 163 1113 164 1117
rect 158 1112 164 1113
rect 246 1117 252 1118
rect 246 1113 247 1117
rect 251 1113 252 1117
rect 246 1112 252 1113
rect 334 1117 340 1118
rect 334 1113 335 1117
rect 339 1113 340 1117
rect 334 1112 340 1113
rect 422 1117 428 1118
rect 422 1113 423 1117
rect 427 1113 428 1117
rect 422 1112 428 1113
rect 1112 1106 1114 1125
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 110 1100 116 1101
rect 1110 1105 1116 1106
rect 1110 1101 1111 1105
rect 1115 1101 1116 1105
rect 1110 1100 1116 1101
rect 110 1087 116 1088
rect 110 1083 111 1087
rect 115 1083 116 1087
rect 110 1082 116 1083
rect 246 1087 252 1088
rect 246 1083 247 1087
rect 251 1083 252 1087
rect 246 1082 252 1083
rect 1110 1087 1116 1088
rect 1110 1083 1111 1087
rect 1115 1083 1116 1087
rect 1110 1082 1116 1083
rect 112 1063 114 1082
rect 150 1072 156 1073
rect 150 1068 151 1072
rect 155 1068 156 1072
rect 150 1067 156 1068
rect 238 1072 244 1073
rect 238 1068 239 1072
rect 243 1068 244 1072
rect 238 1067 244 1068
rect 152 1063 154 1067
rect 240 1063 242 1067
rect 111 1062 115 1063
rect 111 1057 115 1058
rect 135 1062 139 1063
rect 135 1057 139 1058
rect 151 1062 155 1063
rect 151 1057 155 1058
rect 223 1062 227 1063
rect 223 1057 227 1058
rect 239 1062 243 1063
rect 239 1057 243 1058
rect 112 1042 114 1057
rect 134 1056 140 1057
rect 134 1052 135 1056
rect 139 1052 140 1056
rect 134 1051 140 1052
rect 222 1056 228 1057
rect 222 1052 223 1056
rect 227 1052 228 1056
rect 222 1051 228 1052
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 110 1036 116 1037
rect 202 1027 208 1028
rect 110 1023 116 1024
rect 110 1019 111 1023
rect 115 1019 116 1023
rect 202 1023 203 1027
rect 207 1023 208 1027
rect 202 1022 208 1023
rect 110 1018 116 1019
rect 112 995 114 1018
rect 142 1011 148 1012
rect 142 1007 143 1011
rect 147 1007 148 1011
rect 142 1006 148 1007
rect 144 995 146 1006
rect 171 1004 175 1005
rect 170 999 171 1004
rect 175 999 176 1004
rect 170 998 176 999
rect 204 996 206 1022
rect 230 1011 236 1012
rect 230 1007 231 1011
rect 235 1007 236 1011
rect 230 1006 236 1007
rect 202 995 208 996
rect 232 995 234 1006
rect 248 1002 250 1082
rect 326 1072 332 1073
rect 326 1068 327 1072
rect 331 1068 332 1072
rect 326 1067 332 1068
rect 414 1072 420 1073
rect 414 1068 415 1072
rect 419 1068 420 1072
rect 414 1067 420 1068
rect 328 1063 330 1067
rect 416 1063 418 1067
rect 1112 1063 1114 1082
rect 311 1062 315 1063
rect 311 1057 315 1058
rect 327 1062 331 1063
rect 327 1057 331 1058
rect 399 1062 403 1063
rect 399 1057 403 1058
rect 415 1062 419 1063
rect 415 1057 419 1058
rect 1111 1062 1115 1063
rect 1111 1057 1115 1058
rect 310 1056 316 1057
rect 310 1052 311 1056
rect 315 1052 316 1056
rect 310 1051 316 1052
rect 398 1056 404 1057
rect 398 1052 399 1056
rect 403 1052 404 1056
rect 398 1051 404 1052
rect 378 1043 384 1044
rect 378 1039 379 1043
rect 383 1039 384 1043
rect 1112 1042 1114 1057
rect 378 1038 384 1039
rect 1110 1041 1116 1042
rect 318 1031 324 1032
rect 318 1027 319 1031
rect 323 1027 324 1031
rect 318 1026 330 1027
rect 320 1025 330 1026
rect 318 1011 324 1012
rect 318 1007 319 1011
rect 323 1007 324 1011
rect 318 1006 324 1007
rect 258 1003 264 1004
rect 258 1002 259 1003
rect 248 1000 259 1002
rect 258 999 259 1000
rect 263 999 264 1003
rect 258 998 264 999
rect 320 995 322 1006
rect 328 1004 330 1025
rect 380 1005 382 1038
rect 1110 1037 1111 1041
rect 1115 1037 1116 1041
rect 1110 1036 1116 1037
rect 406 1031 412 1032
rect 406 1027 407 1031
rect 411 1027 412 1031
rect 406 1026 412 1027
rect 408 1019 410 1026
rect 1110 1023 1116 1024
rect 1110 1019 1111 1023
rect 1115 1019 1116 1023
rect 408 1017 418 1019
rect 1110 1018 1116 1019
rect 406 1011 412 1012
rect 406 1007 407 1011
rect 411 1007 412 1011
rect 406 1006 412 1007
rect 379 1004 383 1005
rect 326 1003 332 1004
rect 326 999 327 1003
rect 331 999 332 1003
rect 379 999 383 1000
rect 326 998 332 999
rect 408 995 410 1006
rect 416 1004 418 1017
rect 414 1003 420 1004
rect 414 999 415 1003
rect 419 999 420 1003
rect 414 998 420 999
rect 1112 995 1114 1018
rect 111 994 115 995
rect 111 989 115 990
rect 143 994 147 995
rect 202 991 203 995
rect 207 991 208 995
rect 202 990 208 991
rect 231 994 235 995
rect 319 994 323 995
rect 143 989 147 990
rect 231 989 235 990
rect 258 991 264 992
rect 112 970 114 989
rect 144 982 146 989
rect 232 982 234 989
rect 258 987 259 991
rect 263 987 264 991
rect 407 994 411 995
rect 319 989 323 990
rect 346 991 352 992
rect 258 986 264 987
rect 142 981 148 982
rect 142 977 143 981
rect 147 977 148 981
rect 142 976 148 977
rect 230 981 236 982
rect 230 977 231 981
rect 235 977 236 981
rect 230 976 236 977
rect 260 971 262 986
rect 320 982 322 989
rect 346 987 347 991
rect 351 987 352 991
rect 1111 994 1115 995
rect 407 989 411 990
rect 434 991 440 992
rect 346 986 352 987
rect 318 981 324 982
rect 318 977 319 981
rect 323 977 324 981
rect 318 976 324 977
rect 110 969 116 970
rect 110 965 111 969
rect 115 965 116 969
rect 110 964 116 965
rect 232 969 262 971
rect 232 964 234 969
rect 230 963 236 964
rect 230 959 231 963
rect 235 959 236 963
rect 230 958 236 959
rect 318 963 324 964
rect 348 963 350 986
rect 408 982 410 989
rect 434 987 435 991
rect 439 987 440 991
rect 1111 989 1115 990
rect 434 986 440 987
rect 406 981 412 982
rect 406 977 407 981
rect 411 977 412 981
rect 406 976 412 977
rect 436 971 438 986
rect 408 969 438 971
rect 1112 970 1114 989
rect 1110 969 1116 970
rect 408 964 410 969
rect 1110 965 1111 969
rect 1115 965 1116 969
rect 1110 964 1116 965
rect 318 959 319 963
rect 323 961 350 963
rect 406 963 412 964
rect 323 959 324 961
rect 318 958 324 959
rect 406 959 407 963
rect 411 959 412 963
rect 406 958 412 959
rect 110 951 116 952
rect 110 947 111 951
rect 115 947 116 951
rect 1110 951 1116 952
rect 110 946 116 947
rect 466 947 472 948
rect 112 927 114 946
rect 466 943 467 947
rect 471 943 472 947
rect 1110 947 1111 951
rect 1115 947 1116 951
rect 1110 946 1116 947
rect 466 942 472 943
rect 134 936 140 937
rect 134 932 135 936
rect 139 932 140 936
rect 134 931 140 932
rect 222 936 228 937
rect 222 932 223 936
rect 227 932 228 936
rect 222 931 228 932
rect 310 936 316 937
rect 310 932 311 936
rect 315 932 316 936
rect 310 931 316 932
rect 398 936 404 937
rect 398 932 399 936
rect 403 932 404 936
rect 398 931 404 932
rect 136 927 138 931
rect 224 927 226 931
rect 312 927 314 931
rect 400 927 402 931
rect 111 926 115 927
rect 111 921 115 922
rect 135 926 139 927
rect 135 921 139 922
rect 223 926 227 927
rect 223 921 227 922
rect 311 926 315 927
rect 311 921 315 922
rect 399 926 403 927
rect 399 921 403 922
rect 112 906 114 921
rect 134 920 140 921
rect 134 916 135 920
rect 139 916 140 920
rect 134 915 140 916
rect 222 920 228 921
rect 222 916 223 920
rect 227 916 228 920
rect 222 915 228 916
rect 310 920 316 921
rect 310 916 311 920
rect 315 916 316 920
rect 310 915 316 916
rect 398 920 404 921
rect 398 916 399 920
rect 403 916 404 920
rect 398 915 404 916
rect 110 905 116 906
rect 110 901 111 905
rect 115 901 116 905
rect 110 900 116 901
rect 206 891 212 892
rect 110 887 116 888
rect 110 883 111 887
rect 115 883 116 887
rect 206 887 207 891
rect 211 887 212 891
rect 206 886 212 887
rect 290 891 296 892
rect 290 887 291 891
rect 295 887 296 891
rect 290 886 296 887
rect 110 882 116 883
rect 198 883 204 884
rect 112 859 114 882
rect 198 879 199 883
rect 203 879 204 883
rect 198 878 204 879
rect 142 875 148 876
rect 142 871 143 875
rect 147 871 148 875
rect 142 870 148 871
rect 144 859 146 870
rect 111 858 115 859
rect 111 853 115 854
rect 143 858 147 859
rect 200 856 202 878
rect 208 864 210 886
rect 230 875 236 876
rect 230 871 231 875
rect 235 871 236 875
rect 230 870 236 871
rect 206 863 212 864
rect 206 859 207 863
rect 211 859 212 863
rect 232 859 234 870
rect 292 864 294 886
rect 318 875 324 876
rect 318 871 319 875
rect 323 871 324 875
rect 318 870 324 871
rect 406 875 412 876
rect 406 871 407 875
rect 411 871 412 875
rect 406 870 412 871
rect 290 863 296 864
rect 290 859 291 863
rect 295 859 296 863
rect 320 859 322 870
rect 408 859 410 870
rect 468 864 470 942
rect 1112 927 1114 946
rect 1111 926 1115 927
rect 1111 921 1115 922
rect 1112 906 1114 921
rect 1110 905 1116 906
rect 1110 901 1111 905
rect 1115 901 1116 905
rect 1110 900 1116 901
rect 1110 887 1116 888
rect 1110 883 1111 887
rect 1115 883 1116 887
rect 1110 882 1116 883
rect 466 863 472 864
rect 466 859 467 863
rect 471 859 472 863
rect 1112 859 1114 882
rect 206 858 212 859
rect 231 858 235 859
rect 290 858 296 859
rect 319 858 323 859
rect 143 853 147 854
rect 198 855 204 856
rect 112 834 114 853
rect 144 846 146 853
rect 198 851 199 855
rect 203 851 204 855
rect 231 853 235 854
rect 258 855 264 856
rect 198 850 204 851
rect 232 846 234 853
rect 258 851 259 855
rect 263 851 264 855
rect 407 858 411 859
rect 466 858 472 859
rect 495 858 499 859
rect 319 853 323 854
rect 346 855 352 856
rect 258 850 264 851
rect 142 845 148 846
rect 142 841 143 845
rect 147 841 148 845
rect 142 840 148 841
rect 230 845 236 846
rect 230 841 231 845
rect 235 841 236 845
rect 230 840 236 841
rect 260 835 262 850
rect 320 846 322 853
rect 346 851 347 855
rect 351 851 352 855
rect 407 853 411 854
rect 434 855 440 856
rect 346 850 352 851
rect 318 845 324 846
rect 318 841 319 845
rect 323 841 324 845
rect 318 840 324 841
rect 110 833 116 834
rect 110 829 111 833
rect 115 829 116 833
rect 110 828 116 829
rect 232 833 262 835
rect 232 828 234 833
rect 230 827 236 828
rect 230 823 231 827
rect 235 823 236 827
rect 230 822 236 823
rect 318 827 324 828
rect 348 827 350 850
rect 408 846 410 853
rect 434 851 435 855
rect 439 851 440 855
rect 495 853 499 854
rect 1111 858 1115 859
rect 1111 853 1115 854
rect 434 850 440 851
rect 406 845 412 846
rect 406 841 407 845
rect 411 841 412 845
rect 406 840 412 841
rect 436 835 438 850
rect 496 846 498 853
rect 494 845 500 846
rect 494 841 495 845
rect 499 841 500 845
rect 494 840 500 841
rect 408 833 438 835
rect 1112 834 1114 853
rect 1110 833 1116 834
rect 408 828 410 833
rect 1110 829 1111 833
rect 1115 829 1116 833
rect 1110 828 1116 829
rect 318 823 319 827
rect 323 825 350 827
rect 406 827 412 828
rect 323 823 324 825
rect 318 822 324 823
rect 406 823 407 827
rect 411 823 412 827
rect 406 822 412 823
rect 110 815 116 816
rect 110 811 111 815
rect 115 811 116 815
rect 110 810 116 811
rect 474 815 480 816
rect 474 811 475 815
rect 479 811 480 815
rect 474 810 480 811
rect 1110 815 1116 816
rect 1110 811 1111 815
rect 1115 811 1116 815
rect 1110 810 1116 811
rect 112 791 114 810
rect 134 800 140 801
rect 134 796 135 800
rect 139 796 140 800
rect 134 795 140 796
rect 222 800 228 801
rect 222 796 223 800
rect 227 796 228 800
rect 222 795 228 796
rect 310 800 316 801
rect 310 796 311 800
rect 315 796 316 800
rect 310 795 316 796
rect 398 800 404 801
rect 398 796 399 800
rect 403 796 404 800
rect 398 795 404 796
rect 136 791 138 795
rect 224 791 226 795
rect 312 791 314 795
rect 400 791 402 795
rect 111 790 115 791
rect 111 785 115 786
rect 135 790 139 791
rect 135 785 139 786
rect 223 790 227 791
rect 223 785 227 786
rect 231 790 235 791
rect 231 785 235 786
rect 311 790 315 791
rect 311 785 315 786
rect 359 790 363 791
rect 359 785 363 786
rect 399 790 403 791
rect 399 785 403 786
rect 112 770 114 785
rect 134 784 140 785
rect 134 780 135 784
rect 139 780 140 784
rect 134 779 140 780
rect 230 784 236 785
rect 230 780 231 784
rect 235 780 236 784
rect 230 779 236 780
rect 358 784 364 785
rect 358 780 359 784
rect 363 780 364 784
rect 358 779 364 780
rect 110 769 116 770
rect 110 765 111 769
rect 115 765 116 769
rect 110 764 116 765
rect 366 759 372 760
rect 171 756 175 757
rect 110 751 116 752
rect 171 751 175 752
rect 214 755 220 756
rect 214 751 215 755
rect 219 751 220 755
rect 366 755 367 759
rect 371 755 372 759
rect 476 757 478 810
rect 486 800 492 801
rect 486 796 487 800
rect 491 796 492 800
rect 486 795 492 796
rect 488 791 490 795
rect 1112 791 1114 810
rect 487 790 491 791
rect 487 785 491 786
rect 503 790 507 791
rect 503 785 507 786
rect 647 790 651 791
rect 647 785 651 786
rect 799 790 803 791
rect 799 785 803 786
rect 959 790 963 791
rect 959 785 963 786
rect 1111 790 1115 791
rect 1111 785 1115 786
rect 502 784 508 785
rect 502 780 503 784
rect 507 780 508 784
rect 502 779 508 780
rect 646 784 652 785
rect 646 780 647 784
rect 651 780 652 784
rect 646 779 652 780
rect 798 784 804 785
rect 798 780 799 784
rect 803 780 804 784
rect 798 779 804 780
rect 958 784 964 785
rect 958 780 959 784
rect 963 780 964 784
rect 958 779 964 780
rect 1112 770 1114 785
rect 1110 769 1116 770
rect 654 767 660 768
rect 654 763 655 767
rect 659 763 660 767
rect 1110 765 1111 769
rect 1115 765 1116 769
rect 1110 764 1116 765
rect 654 762 660 763
rect 510 759 516 760
rect 475 756 479 757
rect 366 754 378 755
rect 368 753 378 754
rect 110 747 111 751
rect 115 747 116 751
rect 110 746 116 747
rect 112 727 114 746
rect 142 739 148 740
rect 142 735 143 739
rect 147 735 148 739
rect 142 734 148 735
rect 144 727 146 734
rect 172 732 174 751
rect 214 750 220 751
rect 170 731 176 732
rect 170 727 171 731
rect 175 727 176 731
rect 111 726 115 727
rect 111 721 115 722
rect 143 726 147 727
rect 170 726 176 727
rect 216 724 218 750
rect 291 740 295 741
rect 238 739 244 740
rect 238 735 239 739
rect 243 735 244 739
rect 291 735 295 736
rect 366 739 372 740
rect 366 735 367 739
rect 371 735 372 739
rect 238 734 244 735
rect 240 727 242 734
rect 239 726 243 727
rect 143 721 147 722
rect 214 723 220 724
rect 112 702 114 721
rect 214 719 215 723
rect 219 719 220 723
rect 239 721 243 722
rect 263 726 267 727
rect 292 724 294 735
rect 366 734 372 735
rect 368 727 370 734
rect 376 732 378 753
rect 510 755 511 759
rect 515 755 516 759
rect 570 755 576 756
rect 510 754 522 755
rect 512 753 522 754
rect 475 751 479 752
rect 510 739 516 740
rect 510 735 511 739
rect 515 735 516 739
rect 510 734 516 735
rect 374 731 380 732
rect 374 727 375 731
rect 379 727 380 731
rect 359 726 363 727
rect 263 721 267 722
rect 290 723 296 724
rect 214 718 220 719
rect 264 714 266 721
rect 290 719 291 723
rect 295 719 296 723
rect 359 721 363 722
rect 367 726 371 727
rect 374 726 380 727
rect 426 731 432 732
rect 426 727 427 731
rect 431 727 432 731
rect 512 727 514 734
rect 426 726 432 727
rect 463 726 467 727
rect 367 721 371 722
rect 386 721 392 722
rect 290 718 296 719
rect 360 714 362 721
rect 386 717 387 721
rect 391 717 392 721
rect 386 716 392 717
rect 262 713 268 714
rect 262 709 263 713
rect 267 709 268 713
rect 262 708 268 709
rect 358 713 364 714
rect 358 709 359 713
rect 363 709 364 713
rect 358 708 364 709
rect 110 701 116 702
rect 388 701 390 716
rect 110 697 111 701
rect 115 697 116 701
rect 327 700 331 701
rect 387 700 391 701
rect 428 700 430 726
rect 463 721 467 722
rect 511 726 515 727
rect 520 724 522 753
rect 570 751 571 755
rect 575 751 576 755
rect 570 750 576 751
rect 572 741 574 750
rect 656 747 658 762
rect 938 755 944 756
rect 938 751 939 755
rect 943 751 944 755
rect 938 750 944 751
rect 946 755 952 756
rect 946 751 947 755
rect 951 751 952 755
rect 946 750 952 751
rect 1110 751 1116 752
rect 656 745 666 747
rect 571 740 575 741
rect 571 735 575 736
rect 654 739 660 740
rect 654 735 655 739
rect 659 735 660 739
rect 654 734 660 735
rect 558 731 564 732
rect 558 727 559 731
rect 563 727 564 731
rect 656 727 658 734
rect 664 732 666 745
rect 940 741 942 750
rect 939 740 943 741
rect 806 739 812 740
rect 806 735 807 739
rect 811 735 812 739
rect 939 735 943 736
rect 806 734 812 735
rect 662 731 668 732
rect 662 727 663 731
rect 667 727 668 731
rect 808 727 810 734
rect 858 727 864 728
rect 558 726 564 727
rect 575 726 579 727
rect 511 721 515 722
rect 518 723 524 724
rect 464 714 466 721
rect 518 719 519 723
rect 523 719 524 723
rect 518 718 524 719
rect 462 713 468 714
rect 462 709 463 713
rect 467 709 468 713
rect 462 708 468 709
rect 560 700 562 726
rect 575 721 579 722
rect 655 726 659 727
rect 662 726 668 727
rect 687 726 691 727
rect 655 721 659 722
rect 799 726 803 727
rect 687 721 691 722
rect 714 723 720 724
rect 576 714 578 721
rect 688 714 690 721
rect 714 719 715 723
rect 719 719 720 723
rect 799 721 803 722
rect 807 726 811 727
rect 858 723 859 727
rect 863 723 864 727
rect 858 722 864 723
rect 919 726 923 727
rect 948 724 950 750
rect 1110 747 1111 751
rect 1115 747 1116 751
rect 1110 746 1116 747
rect 995 740 999 741
rect 966 739 972 740
rect 966 735 967 739
rect 971 735 972 739
rect 995 735 999 736
rect 966 734 972 735
rect 968 727 970 734
rect 996 732 998 735
rect 994 731 1000 732
rect 994 727 995 731
rect 999 727 1000 731
rect 967 726 971 727
rect 994 726 1000 727
rect 1014 731 1020 732
rect 1014 727 1015 731
rect 1019 727 1020 731
rect 1112 727 1114 746
rect 1014 726 1020 727
rect 1023 726 1027 727
rect 807 721 811 722
rect 826 721 832 722
rect 714 718 720 719
rect 574 713 580 714
rect 574 709 575 713
rect 579 709 580 713
rect 574 708 580 709
rect 686 713 692 714
rect 686 709 687 713
rect 691 709 692 713
rect 686 708 692 709
rect 110 696 116 697
rect 326 695 327 700
rect 331 695 332 700
rect 387 695 391 696
rect 426 699 432 700
rect 426 695 427 699
rect 431 695 432 699
rect 326 694 332 695
rect 426 694 432 695
rect 558 699 564 700
rect 716 699 718 718
rect 800 714 802 721
rect 826 717 827 721
rect 831 717 832 721
rect 826 716 832 717
rect 798 713 804 714
rect 798 709 799 713
rect 803 709 804 713
rect 798 708 804 709
rect 558 695 559 699
rect 563 695 564 699
rect 696 698 718 699
rect 692 697 718 698
rect 692 696 698 697
rect 558 694 564 695
rect 682 695 688 696
rect 682 691 683 695
rect 687 691 688 695
rect 692 691 694 696
rect 682 690 694 691
rect 684 689 694 690
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 110 678 116 679
rect 642 683 648 684
rect 642 679 643 683
rect 647 679 648 683
rect 642 678 648 679
rect 112 655 114 678
rect 254 668 260 669
rect 254 664 255 668
rect 259 664 260 668
rect 254 663 260 664
rect 350 668 356 669
rect 350 664 351 668
rect 355 664 356 668
rect 350 663 356 664
rect 454 668 460 669
rect 454 664 455 668
rect 459 664 460 668
rect 454 663 460 664
rect 566 668 572 669
rect 566 664 567 668
rect 571 664 572 668
rect 566 663 572 664
rect 256 655 258 663
rect 352 655 354 663
rect 456 655 458 663
rect 506 655 512 656
rect 568 655 570 663
rect 644 656 646 678
rect 678 668 684 669
rect 678 664 679 668
rect 683 664 684 668
rect 678 663 684 664
rect 790 668 796 669
rect 790 664 791 668
rect 795 664 796 668
rect 790 663 796 664
rect 642 655 648 656
rect 680 655 682 663
rect 792 655 794 663
rect 111 654 115 655
rect 111 649 115 650
rect 255 654 259 655
rect 255 649 259 650
rect 351 654 355 655
rect 351 649 355 650
rect 455 654 459 655
rect 455 649 459 650
rect 471 654 475 655
rect 506 651 507 655
rect 511 651 512 655
rect 506 650 512 651
rect 567 654 571 655
rect 642 651 643 655
rect 647 651 648 655
rect 642 650 648 651
rect 671 654 675 655
rect 471 649 475 650
rect 112 634 114 649
rect 470 648 476 649
rect 470 644 471 648
rect 475 644 476 648
rect 470 643 476 644
rect 110 633 116 634
rect 110 629 111 633
rect 115 629 116 633
rect 110 628 116 629
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 110 610 116 611
rect 112 587 114 610
rect 478 603 484 604
rect 478 599 479 603
rect 483 599 484 603
rect 478 598 484 599
rect 480 587 482 598
rect 508 596 510 650
rect 567 649 571 650
rect 671 649 675 650
rect 679 654 683 655
rect 679 649 683 650
rect 783 654 787 655
rect 783 649 787 650
rect 791 654 795 655
rect 828 652 830 716
rect 860 700 862 722
rect 919 721 923 722
rect 946 723 952 724
rect 920 714 922 721
rect 946 719 947 723
rect 951 719 952 723
rect 967 721 971 722
rect 946 718 952 719
rect 918 713 924 714
rect 918 709 919 713
rect 923 709 924 713
rect 918 708 924 709
rect 858 699 864 700
rect 858 695 859 699
rect 863 695 864 699
rect 1016 696 1018 726
rect 1023 721 1027 722
rect 1111 726 1115 727
rect 1111 721 1115 722
rect 1024 714 1026 721
rect 1022 713 1028 714
rect 1022 709 1023 713
rect 1027 709 1028 713
rect 1022 708 1028 709
rect 1112 702 1114 721
rect 1110 701 1116 702
rect 1110 697 1111 701
rect 1115 697 1116 701
rect 1110 696 1116 697
rect 858 694 864 695
rect 1014 695 1020 696
rect 1014 691 1015 695
rect 1019 691 1020 695
rect 1014 690 1020 691
rect 1022 683 1028 684
rect 1022 679 1023 683
rect 1027 679 1028 683
rect 1022 678 1028 679
rect 1110 683 1116 684
rect 1110 679 1111 683
rect 1115 679 1116 683
rect 1110 678 1116 679
rect 910 668 916 669
rect 910 664 911 668
rect 915 664 916 668
rect 910 663 916 664
rect 1014 668 1020 669
rect 1014 664 1015 668
rect 1019 664 1020 668
rect 1014 663 1020 664
rect 912 655 914 663
rect 1016 655 1018 663
rect 1024 660 1026 678
rect 1022 659 1028 660
rect 1022 655 1023 659
rect 1027 655 1028 659
rect 903 654 907 655
rect 791 649 795 650
rect 826 651 832 652
rect 566 648 572 649
rect 566 644 567 648
rect 571 644 572 648
rect 566 643 572 644
rect 670 648 676 649
rect 670 644 671 648
rect 675 644 676 648
rect 670 643 676 644
rect 782 648 788 649
rect 782 644 783 648
rect 787 644 788 648
rect 826 647 827 651
rect 831 647 832 651
rect 903 649 907 650
rect 911 654 915 655
rect 911 649 915 650
rect 1015 654 1019 655
rect 1022 654 1028 655
rect 1050 659 1056 660
rect 1050 655 1051 659
rect 1055 655 1056 659
rect 1112 655 1114 678
rect 1050 654 1056 655
rect 1111 654 1115 655
rect 1015 649 1019 650
rect 826 646 832 647
rect 902 648 908 649
rect 782 643 788 644
rect 902 644 903 648
rect 907 644 908 648
rect 902 643 908 644
rect 1014 648 1020 649
rect 1014 644 1015 648
rect 1019 644 1020 648
rect 1014 643 1020 644
rect 790 631 796 632
rect 790 627 791 631
rect 795 627 796 631
rect 790 626 796 627
rect 574 623 580 624
rect 574 619 575 623
rect 579 619 580 623
rect 574 618 580 619
rect 678 623 684 624
rect 678 619 679 623
rect 683 619 684 623
rect 678 618 690 619
rect 576 611 578 618
rect 680 617 690 618
rect 576 609 586 611
rect 574 603 580 604
rect 574 599 575 603
rect 579 599 580 603
rect 574 598 580 599
rect 506 595 512 596
rect 506 591 507 595
rect 511 591 512 595
rect 506 590 512 591
rect 554 587 560 588
rect 576 587 578 598
rect 584 596 586 609
rect 678 603 684 604
rect 678 599 679 603
rect 683 599 684 603
rect 678 598 684 599
rect 582 595 588 596
rect 582 591 583 595
rect 587 591 588 595
rect 582 590 588 591
rect 650 587 656 588
rect 680 587 682 598
rect 688 596 690 617
rect 792 611 794 626
rect 792 609 802 611
rect 790 603 796 604
rect 790 599 791 603
rect 795 599 796 603
rect 790 598 796 599
rect 686 595 692 596
rect 686 591 687 595
rect 691 591 692 595
rect 686 590 692 591
rect 738 587 744 588
rect 792 587 794 598
rect 800 588 802 609
rect 910 603 916 604
rect 910 599 911 603
rect 915 599 916 603
rect 910 598 916 599
rect 1022 603 1028 604
rect 1022 599 1023 603
rect 1027 599 1028 603
rect 1022 598 1028 599
rect 798 587 804 588
rect 912 587 914 598
rect 1002 587 1008 588
rect 1024 587 1026 598
rect 1052 596 1054 654
rect 1111 649 1115 650
rect 1112 634 1114 649
rect 1110 633 1116 634
rect 1110 629 1111 633
rect 1115 629 1116 633
rect 1110 628 1116 629
rect 1082 619 1088 620
rect 1082 615 1083 619
rect 1087 615 1088 619
rect 1082 614 1088 615
rect 1110 615 1116 616
rect 1050 595 1056 596
rect 1050 591 1051 595
rect 1055 591 1056 595
rect 1050 590 1056 591
rect 1084 588 1086 614
rect 1110 611 1111 615
rect 1115 611 1116 615
rect 1110 610 1116 611
rect 1082 587 1088 588
rect 1112 587 1114 610
rect 111 586 115 587
rect 111 581 115 582
rect 479 586 483 587
rect 479 581 483 582
rect 495 586 499 587
rect 554 583 555 587
rect 559 583 560 587
rect 554 582 560 583
rect 575 586 579 587
rect 495 581 499 582
rect 112 562 114 581
rect 496 574 498 581
rect 494 573 500 574
rect 494 569 495 573
rect 499 569 500 573
rect 494 568 500 569
rect 110 561 116 562
rect 110 557 111 561
rect 115 557 116 561
rect 556 560 558 582
rect 575 581 579 582
rect 583 586 587 587
rect 650 583 651 587
rect 655 583 656 587
rect 650 582 656 583
rect 671 586 675 587
rect 583 581 587 582
rect 584 574 586 581
rect 582 573 588 574
rect 582 569 583 573
rect 587 569 588 573
rect 582 568 588 569
rect 110 556 116 557
rect 554 559 560 560
rect 554 555 555 559
rect 559 555 560 559
rect 652 556 654 582
rect 671 581 675 582
rect 679 586 683 587
rect 738 583 739 587
rect 743 583 744 587
rect 738 582 744 583
rect 759 586 763 587
rect 679 581 683 582
rect 672 574 674 581
rect 670 573 676 574
rect 670 569 671 573
rect 675 569 676 573
rect 670 568 676 569
rect 740 556 742 582
rect 759 581 763 582
rect 791 586 795 587
rect 798 583 799 587
rect 803 583 804 587
rect 798 582 804 583
rect 847 586 851 587
rect 911 586 915 587
rect 791 581 795 582
rect 847 581 851 582
rect 874 583 880 584
rect 760 574 762 581
rect 848 574 850 581
rect 874 579 875 583
rect 879 579 880 583
rect 911 581 915 582
rect 935 586 939 587
rect 1002 583 1003 587
rect 1007 583 1008 587
rect 1002 582 1008 583
rect 1023 586 1027 587
rect 1082 583 1083 587
rect 1087 583 1088 587
rect 1082 582 1088 583
rect 1111 586 1115 587
rect 935 581 939 582
rect 874 578 880 579
rect 758 573 764 574
rect 758 569 759 573
rect 763 569 764 573
rect 758 568 764 569
rect 846 573 852 574
rect 846 569 847 573
rect 851 569 852 573
rect 846 568 852 569
rect 554 554 560 555
rect 650 555 656 556
rect 650 551 651 555
rect 655 551 656 555
rect 650 550 656 551
rect 738 555 744 556
rect 738 551 739 555
rect 743 551 744 555
rect 738 550 744 551
rect 110 543 116 544
rect 110 539 111 543
rect 115 539 116 543
rect 110 538 116 539
rect 112 519 114 538
rect 486 528 492 529
rect 486 524 487 528
rect 491 524 492 528
rect 486 523 492 524
rect 574 528 580 529
rect 574 524 575 528
rect 579 524 580 528
rect 574 523 580 524
rect 662 528 668 529
rect 662 524 663 528
rect 667 524 668 528
rect 662 523 668 524
rect 750 528 756 529
rect 750 524 751 528
rect 755 524 756 528
rect 750 523 756 524
rect 838 528 844 529
rect 876 528 878 578
rect 936 574 938 581
rect 934 573 940 574
rect 934 569 935 573
rect 939 569 940 573
rect 934 568 940 569
rect 1004 556 1006 582
rect 1023 581 1027 582
rect 1111 581 1115 582
rect 1024 574 1026 581
rect 1022 573 1028 574
rect 1022 569 1023 573
rect 1027 569 1028 573
rect 1022 568 1028 569
rect 1112 562 1114 581
rect 1110 561 1116 562
rect 1110 557 1111 561
rect 1115 557 1116 561
rect 1110 556 1116 557
rect 1002 555 1008 556
rect 1002 551 1003 555
rect 1007 551 1008 555
rect 1002 550 1008 551
rect 1022 543 1028 544
rect 1022 539 1023 543
rect 1027 539 1028 543
rect 1022 538 1028 539
rect 1110 543 1116 544
rect 1110 539 1111 543
rect 1115 539 1116 543
rect 1110 538 1116 539
rect 926 528 932 529
rect 838 524 839 528
rect 843 524 844 528
rect 838 523 844 524
rect 854 527 860 528
rect 854 523 855 527
rect 859 523 860 527
rect 488 519 490 523
rect 576 519 578 523
rect 664 519 666 523
rect 752 519 754 523
rect 840 519 842 523
rect 854 522 860 523
rect 874 527 880 528
rect 874 523 875 527
rect 879 523 880 527
rect 926 524 927 528
rect 931 524 932 528
rect 926 523 932 524
rect 1014 528 1020 529
rect 1014 524 1015 528
rect 1019 524 1020 528
rect 1014 523 1020 524
rect 874 522 880 523
rect 111 518 115 519
rect 111 513 115 514
rect 375 518 379 519
rect 375 513 379 514
rect 487 518 491 519
rect 487 513 491 514
rect 575 518 579 519
rect 575 513 579 514
rect 599 518 603 519
rect 599 513 603 514
rect 663 518 667 519
rect 663 513 667 514
rect 719 518 723 519
rect 719 513 723 514
rect 751 518 755 519
rect 751 513 755 514
rect 839 518 843 519
rect 839 513 843 514
rect 847 518 851 519
rect 847 513 851 514
rect 112 498 114 513
rect 374 512 380 513
rect 374 508 375 512
rect 379 508 380 512
rect 374 507 380 508
rect 486 512 492 513
rect 486 508 487 512
rect 491 508 492 512
rect 486 507 492 508
rect 598 512 604 513
rect 598 508 599 512
rect 603 508 604 512
rect 598 507 604 508
rect 718 512 724 513
rect 718 508 719 512
rect 723 508 724 512
rect 718 507 724 508
rect 846 512 852 513
rect 846 508 847 512
rect 851 508 852 512
rect 846 507 852 508
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 856 496 858 522
rect 928 519 930 523
rect 1016 519 1018 523
rect 927 518 931 519
rect 927 513 931 514
rect 983 518 987 519
rect 983 513 987 514
rect 1015 518 1019 519
rect 1015 513 1019 514
rect 982 512 988 513
rect 982 508 983 512
rect 987 508 988 512
rect 982 507 988 508
rect 1024 499 1026 538
rect 1112 519 1114 538
rect 1111 518 1115 519
rect 1111 513 1115 514
rect 1020 497 1026 499
rect 1112 498 1114 513
rect 1110 497 1116 498
rect 110 492 116 493
rect 854 495 860 496
rect 726 491 732 492
rect 726 487 727 491
rect 731 487 732 491
rect 854 491 855 495
rect 859 491 860 495
rect 854 490 860 491
rect 726 486 732 487
rect 554 483 560 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 554 479 555 483
rect 559 479 560 483
rect 554 478 560 479
rect 710 483 716 484
rect 710 479 711 483
rect 715 479 716 483
rect 728 483 730 486
rect 728 481 738 483
rect 710 478 716 479
rect 110 474 116 475
rect 112 447 114 474
rect 382 467 388 468
rect 382 463 383 467
rect 387 463 388 467
rect 382 462 388 463
rect 494 467 500 468
rect 494 463 495 467
rect 499 463 500 467
rect 494 462 500 463
rect 358 447 364 448
rect 384 447 386 462
rect 411 460 415 461
rect 410 455 411 460
rect 415 455 416 460
rect 410 454 416 455
rect 496 447 498 462
rect 556 448 558 478
rect 606 467 612 468
rect 606 463 607 467
rect 611 463 612 467
rect 606 462 612 463
rect 554 447 560 448
rect 608 447 610 462
rect 712 461 714 478
rect 726 467 732 468
rect 726 463 727 467
rect 731 463 732 467
rect 726 462 732 463
rect 711 460 715 461
rect 711 455 715 456
rect 728 447 730 462
rect 736 460 738 481
rect 854 467 860 468
rect 854 463 855 467
rect 859 463 860 467
rect 854 462 860 463
rect 990 467 996 468
rect 990 463 991 467
rect 995 463 996 467
rect 990 462 996 463
rect 734 459 740 460
rect 734 455 735 459
rect 739 455 740 459
rect 734 454 740 455
rect 818 451 824 452
rect 818 447 819 451
rect 823 447 824 451
rect 856 447 858 462
rect 992 447 994 462
rect 1020 460 1022 497
rect 1110 493 1111 497
rect 1115 493 1116 497
rect 1110 492 1116 493
rect 1050 483 1056 484
rect 1050 479 1051 483
rect 1055 479 1056 483
rect 1050 478 1056 479
rect 1110 479 1116 480
rect 1018 459 1024 460
rect 1018 455 1019 459
rect 1023 455 1024 459
rect 1018 454 1024 455
rect 1052 448 1054 478
rect 1110 475 1111 479
rect 1115 475 1116 479
rect 1110 474 1116 475
rect 1050 447 1056 448
rect 1112 447 1114 474
rect 111 446 115 447
rect 111 441 115 442
rect 263 446 267 447
rect 358 443 359 447
rect 363 443 364 447
rect 358 442 364 443
rect 383 446 387 447
rect 263 441 267 442
rect 112 422 114 441
rect 264 434 266 441
rect 262 433 268 434
rect 262 429 263 433
rect 267 429 268 433
rect 262 428 268 429
rect 110 421 116 422
rect 360 421 362 442
rect 383 441 387 442
rect 391 446 395 447
rect 391 441 395 442
rect 495 446 499 447
rect 495 441 499 442
rect 511 446 515 447
rect 554 443 555 447
rect 559 443 560 447
rect 554 442 560 443
rect 607 446 611 447
rect 511 441 515 442
rect 607 441 611 442
rect 631 446 635 447
rect 727 446 731 447
rect 631 441 635 442
rect 658 443 664 444
rect 392 434 394 441
rect 512 434 514 441
rect 632 434 634 441
rect 658 439 659 443
rect 663 439 664 443
rect 727 441 731 442
rect 751 446 755 447
rect 818 446 824 447
rect 855 446 859 447
rect 751 441 755 442
rect 658 438 664 439
rect 390 433 396 434
rect 390 429 391 433
rect 395 429 396 433
rect 390 428 396 429
rect 510 433 516 434
rect 510 429 511 433
rect 515 429 516 433
rect 510 428 516 429
rect 630 433 636 434
rect 630 429 631 433
rect 635 429 636 433
rect 630 428 636 429
rect 110 417 111 421
rect 115 417 116 421
rect 110 416 116 417
rect 359 420 363 421
rect 459 420 463 421
rect 359 415 363 416
rect 458 415 464 416
rect 458 411 459 415
rect 463 411 464 415
rect 458 410 464 411
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 110 398 116 399
rect 450 399 456 400
rect 112 379 114 398
rect 450 395 451 399
rect 455 395 456 399
rect 450 394 456 395
rect 254 388 260 389
rect 254 384 255 388
rect 259 384 260 388
rect 254 383 260 384
rect 382 388 388 389
rect 382 384 383 388
rect 387 384 388 388
rect 382 383 388 384
rect 256 379 258 383
rect 384 379 386 383
rect 111 378 115 379
rect 111 373 115 374
rect 135 378 139 379
rect 135 373 139 374
rect 255 378 259 379
rect 255 373 259 374
rect 383 378 387 379
rect 383 373 387 374
rect 415 378 419 379
rect 415 373 419 374
rect 112 358 114 373
rect 134 372 140 373
rect 134 368 135 372
rect 139 368 140 372
rect 134 367 140 368
rect 254 372 260 373
rect 254 368 255 372
rect 259 368 260 372
rect 254 367 260 368
rect 414 372 420 373
rect 414 368 415 372
rect 419 368 420 372
rect 414 367 420 368
rect 110 357 116 358
rect 110 353 111 357
rect 115 353 116 357
rect 110 352 116 353
rect 202 343 208 344
rect 110 339 116 340
rect 110 335 111 339
rect 115 335 116 339
rect 202 339 203 343
rect 207 339 208 343
rect 202 338 208 339
rect 110 334 116 335
rect 112 311 114 334
rect 142 327 148 328
rect 142 323 143 327
rect 147 323 148 327
rect 142 322 148 323
rect 144 311 146 322
rect 111 310 115 311
rect 111 305 115 306
rect 143 310 147 311
rect 204 308 206 338
rect 262 327 268 328
rect 262 323 263 327
rect 267 323 268 327
rect 422 327 428 328
rect 262 322 268 323
rect 291 324 295 325
rect 264 311 266 322
rect 422 323 423 327
rect 427 323 428 327
rect 422 322 428 323
rect 290 319 296 320
rect 290 315 291 319
rect 295 315 296 319
rect 290 314 296 315
rect 424 311 426 322
rect 452 320 454 394
rect 502 388 508 389
rect 502 384 503 388
rect 507 384 508 388
rect 502 383 508 384
rect 622 388 628 389
rect 622 384 623 388
rect 627 384 628 388
rect 622 383 628 384
rect 504 379 506 383
rect 624 379 626 383
rect 503 378 507 379
rect 503 373 507 374
rect 583 378 587 379
rect 583 373 587 374
rect 623 378 627 379
rect 623 373 627 374
rect 582 372 588 373
rect 582 368 583 372
rect 587 368 588 372
rect 582 367 588 368
rect 660 360 662 438
rect 752 434 754 441
rect 750 433 756 434
rect 750 429 751 433
rect 755 429 756 433
rect 750 428 756 429
rect 820 420 822 446
rect 855 441 859 442
rect 879 446 883 447
rect 879 441 883 442
rect 991 446 995 447
rect 991 441 995 442
rect 1007 446 1011 447
rect 1050 443 1051 447
rect 1055 443 1056 447
rect 1050 442 1056 443
rect 1111 446 1115 447
rect 1007 441 1011 442
rect 1111 441 1115 442
rect 880 434 882 441
rect 1008 434 1010 441
rect 878 433 884 434
rect 878 429 879 433
rect 883 429 884 433
rect 878 428 884 429
rect 1006 433 1012 434
rect 1006 429 1007 433
rect 1011 429 1012 433
rect 1006 428 1012 429
rect 1112 422 1114 441
rect 1110 421 1116 422
rect 818 419 824 420
rect 818 415 819 419
rect 823 415 824 419
rect 1110 417 1111 421
rect 1115 417 1116 421
rect 1110 416 1116 417
rect 818 414 824 415
rect 970 403 976 404
rect 970 399 971 403
rect 975 399 976 403
rect 970 398 976 399
rect 1110 403 1116 404
rect 1110 399 1111 403
rect 1115 399 1116 403
rect 1110 398 1116 399
rect 742 388 748 389
rect 742 384 743 388
rect 747 384 748 388
rect 742 383 748 384
rect 870 388 876 389
rect 870 384 871 388
rect 875 384 876 388
rect 870 383 876 384
rect 744 379 746 383
rect 872 379 874 383
rect 743 378 747 379
rect 743 373 747 374
rect 759 378 763 379
rect 759 373 763 374
rect 871 378 875 379
rect 871 373 875 374
rect 935 378 939 379
rect 935 373 939 374
rect 758 372 764 373
rect 758 368 759 372
rect 763 368 764 372
rect 758 367 764 368
rect 934 372 940 373
rect 934 368 935 372
rect 939 368 940 372
rect 934 367 940 368
rect 658 359 664 360
rect 658 355 659 359
rect 663 355 664 359
rect 658 354 664 355
rect 490 343 496 344
rect 490 338 491 343
rect 495 338 496 343
rect 498 343 504 344
rect 498 339 499 343
rect 503 339 504 343
rect 898 343 904 344
rect 498 338 504 339
rect 619 340 623 341
rect 491 335 495 336
rect 500 325 502 338
rect 898 339 899 343
rect 903 339 904 343
rect 898 338 904 339
rect 619 335 623 336
rect 590 327 596 328
rect 499 324 503 325
rect 590 323 591 327
rect 595 323 596 327
rect 590 322 596 323
rect 450 319 456 320
rect 499 319 503 320
rect 450 315 451 319
rect 455 315 456 319
rect 450 314 456 315
rect 592 311 594 322
rect 620 320 622 335
rect 766 327 772 328
rect 766 323 767 327
rect 771 323 772 327
rect 766 322 772 323
rect 618 319 624 320
rect 618 315 619 319
rect 623 315 624 319
rect 618 314 624 315
rect 638 315 644 316
rect 638 311 639 315
rect 643 311 644 315
rect 768 311 770 322
rect 794 319 800 320
rect 794 315 795 319
rect 799 315 800 319
rect 794 314 800 315
rect 263 310 267 311
rect 143 305 147 306
rect 202 307 208 308
rect 112 286 114 305
rect 144 298 146 305
rect 202 303 203 307
rect 207 303 208 307
rect 263 305 267 306
rect 271 310 275 311
rect 423 310 427 311
rect 271 305 275 306
rect 298 307 304 308
rect 202 302 208 303
rect 272 298 274 305
rect 298 303 299 307
rect 303 303 304 307
rect 575 310 579 311
rect 423 305 427 306
rect 450 307 456 308
rect 298 302 304 303
rect 142 297 148 298
rect 142 293 143 297
rect 147 293 148 297
rect 142 292 148 293
rect 270 297 276 298
rect 270 293 271 297
rect 275 293 276 297
rect 270 292 276 293
rect 110 285 116 286
rect 300 285 302 302
rect 424 298 426 305
rect 450 303 451 307
rect 455 303 456 307
rect 575 305 579 306
rect 591 310 595 311
rect 638 310 644 311
rect 719 310 723 311
rect 591 305 595 306
rect 602 307 608 308
rect 450 302 456 303
rect 422 297 428 298
rect 422 293 423 297
rect 427 293 428 297
rect 422 292 428 293
rect 452 285 454 302
rect 576 298 578 305
rect 602 303 603 307
rect 607 303 608 307
rect 602 302 608 303
rect 574 297 580 298
rect 574 293 575 297
rect 579 293 580 297
rect 574 292 580 293
rect 110 281 111 285
rect 115 281 116 285
rect 223 284 227 285
rect 299 284 303 285
rect 383 284 387 285
rect 451 284 455 285
rect 110 280 116 281
rect 222 279 223 284
rect 227 279 228 284
rect 299 279 303 280
rect 382 279 383 284
rect 387 279 388 284
rect 451 279 455 280
rect 222 278 228 279
rect 382 278 388 279
rect 110 267 116 268
rect 110 263 111 267
rect 115 263 116 267
rect 110 262 116 263
rect 522 267 528 268
rect 522 263 523 267
rect 527 263 528 267
rect 522 262 528 263
rect 112 243 114 262
rect 134 252 140 253
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 262 252 268 253
rect 262 248 263 252
rect 267 248 268 252
rect 262 247 268 248
rect 414 252 420 253
rect 414 248 415 252
rect 419 248 420 252
rect 414 247 420 248
rect 136 243 138 247
rect 264 243 266 247
rect 416 243 418 247
rect 111 242 115 243
rect 111 237 115 238
rect 135 242 139 243
rect 135 237 139 238
rect 175 242 179 243
rect 175 237 179 238
rect 263 242 267 243
rect 263 237 267 238
rect 327 242 331 243
rect 327 237 331 238
rect 415 242 419 243
rect 415 237 419 238
rect 487 242 491 243
rect 487 237 491 238
rect 112 222 114 237
rect 174 236 180 237
rect 174 232 175 236
rect 179 232 180 236
rect 174 231 180 232
rect 326 236 332 237
rect 326 232 327 236
rect 331 232 332 236
rect 326 231 332 232
rect 486 236 492 237
rect 486 232 487 236
rect 491 232 492 236
rect 486 231 492 232
rect 110 221 116 222
rect 110 217 111 221
rect 115 217 116 221
rect 110 216 116 217
rect 170 211 176 212
rect 170 207 171 211
rect 175 207 176 211
rect 170 206 176 207
rect 434 207 440 208
rect 110 203 116 204
rect 110 199 111 203
rect 115 199 116 203
rect 110 198 116 199
rect 112 163 114 198
rect 111 162 115 163
rect 111 157 115 158
rect 143 162 147 163
rect 172 160 174 206
rect 434 203 435 207
rect 439 203 440 207
rect 434 202 440 203
rect 182 191 188 192
rect 182 187 183 191
rect 187 187 188 191
rect 182 186 188 187
rect 334 191 340 192
rect 334 187 335 191
rect 339 187 340 191
rect 334 186 340 187
rect 184 163 186 186
rect 202 167 208 168
rect 202 163 203 167
rect 207 163 208 167
rect 290 167 296 168
rect 290 163 291 167
rect 295 163 296 167
rect 336 163 338 186
rect 436 180 438 202
rect 494 191 500 192
rect 494 187 495 191
rect 499 187 500 191
rect 494 186 500 187
rect 434 179 440 180
rect 434 175 435 179
rect 439 175 440 179
rect 434 174 440 175
rect 378 167 384 168
rect 378 163 379 167
rect 383 163 384 167
rect 466 167 472 168
rect 466 163 467 167
rect 471 163 472 167
rect 496 163 498 186
rect 524 184 526 262
rect 566 252 572 253
rect 566 248 567 252
rect 571 248 572 252
rect 566 247 572 248
rect 568 243 570 247
rect 567 242 571 243
rect 567 237 571 238
rect 604 224 606 302
rect 640 284 642 310
rect 719 305 723 306
rect 767 310 771 311
rect 767 305 771 306
rect 720 298 722 305
rect 718 297 724 298
rect 718 293 719 297
rect 723 293 724 297
rect 718 292 724 293
rect 796 284 798 314
rect 871 310 875 311
rect 900 308 902 338
rect 942 327 948 328
rect 942 323 943 327
rect 947 323 948 327
rect 942 322 948 323
rect 944 311 946 322
rect 972 320 974 398
rect 998 388 1004 389
rect 998 384 999 388
rect 1003 384 1004 388
rect 998 383 1004 384
rect 1000 379 1002 383
rect 1112 379 1114 398
rect 999 378 1003 379
rect 999 373 1003 374
rect 1111 378 1115 379
rect 1111 373 1115 374
rect 1112 358 1114 373
rect 1110 357 1116 358
rect 1110 353 1111 357
rect 1115 353 1116 357
rect 1110 352 1116 353
rect 1110 339 1116 340
rect 1110 335 1111 339
rect 1115 335 1116 339
rect 1110 334 1116 335
rect 970 319 976 320
rect 970 315 971 319
rect 975 315 976 319
rect 970 314 976 315
rect 990 315 996 316
rect 990 311 991 315
rect 995 311 996 315
rect 1112 311 1114 334
rect 943 310 947 311
rect 990 310 996 311
rect 1023 310 1027 311
rect 871 305 875 306
rect 898 307 904 308
rect 872 298 874 305
rect 898 303 899 307
rect 903 303 904 307
rect 943 305 947 306
rect 898 302 904 303
rect 870 297 876 298
rect 870 293 871 297
rect 875 293 876 297
rect 870 292 876 293
rect 992 284 994 310
rect 1023 305 1027 306
rect 1111 310 1115 311
rect 1111 305 1115 306
rect 1024 298 1026 305
rect 1022 297 1028 298
rect 1022 293 1023 297
rect 1027 293 1028 297
rect 1022 292 1028 293
rect 1112 286 1114 305
rect 1110 285 1116 286
rect 638 283 644 284
rect 638 279 639 283
rect 643 279 644 283
rect 638 278 644 279
rect 794 283 800 284
rect 794 279 795 283
rect 799 279 800 283
rect 794 278 800 279
rect 990 283 996 284
rect 990 279 991 283
rect 995 279 996 283
rect 1110 281 1111 285
rect 1115 281 1116 285
rect 1110 280 1116 281
rect 990 278 996 279
rect 1022 267 1028 268
rect 1022 263 1023 267
rect 1027 263 1028 267
rect 1022 262 1028 263
rect 1110 267 1116 268
rect 1110 263 1111 267
rect 1115 263 1116 267
rect 1110 262 1116 263
rect 710 252 716 253
rect 710 248 711 252
rect 715 248 716 252
rect 710 247 716 248
rect 862 252 868 253
rect 862 248 863 252
rect 867 248 868 252
rect 862 247 868 248
rect 1014 252 1020 253
rect 1014 248 1015 252
rect 1019 248 1020 252
rect 1014 247 1020 248
rect 712 243 714 247
rect 864 243 866 247
rect 1016 243 1018 247
rect 655 242 659 243
rect 655 237 659 238
rect 711 242 715 243
rect 711 237 715 238
rect 831 242 835 243
rect 831 237 835 238
rect 863 242 867 243
rect 863 237 867 238
rect 1007 242 1011 243
rect 1007 237 1011 238
rect 1015 242 1019 243
rect 1015 237 1019 238
rect 654 236 660 237
rect 654 232 655 236
rect 659 232 660 236
rect 654 231 660 232
rect 830 236 836 237
rect 830 232 831 236
rect 835 232 836 236
rect 830 231 836 232
rect 1006 236 1012 237
rect 1006 232 1007 236
rect 1011 232 1012 236
rect 1006 231 1012 232
rect 602 223 608 224
rect 602 219 603 223
rect 607 219 608 223
rect 602 218 608 219
rect 770 207 776 208
rect 770 203 771 207
rect 775 203 776 207
rect 770 202 776 203
rect 662 191 668 192
rect 662 187 663 191
rect 667 187 668 191
rect 662 186 668 187
rect 522 183 528 184
rect 522 179 523 183
rect 527 179 528 183
rect 522 178 528 179
rect 554 167 560 168
rect 554 163 555 167
rect 559 163 560 167
rect 642 167 648 168
rect 642 163 643 167
rect 647 163 648 167
rect 664 163 666 186
rect 772 180 774 202
rect 838 191 844 192
rect 838 187 839 191
rect 843 187 844 191
rect 838 186 844 187
rect 1014 191 1020 192
rect 1014 187 1015 191
rect 1019 187 1020 191
rect 1014 186 1020 187
rect 770 179 776 180
rect 770 175 771 179
rect 775 175 776 179
rect 770 174 776 175
rect 818 175 824 176
rect 818 171 819 175
rect 823 171 824 175
rect 818 170 824 171
rect 730 167 736 168
rect 730 163 731 167
rect 735 163 736 167
rect 183 162 187 163
rect 202 162 208 163
rect 231 162 235 163
rect 290 162 296 163
rect 319 162 323 163
rect 143 157 147 158
rect 170 159 176 160
rect 112 138 114 157
rect 144 150 146 157
rect 170 155 171 159
rect 175 155 176 159
rect 183 157 187 158
rect 170 154 176 155
rect 142 149 148 150
rect 142 145 143 149
rect 147 145 148 149
rect 142 144 148 145
rect 110 137 116 138
rect 110 133 111 137
rect 115 133 116 137
rect 204 136 206 162
rect 231 157 235 158
rect 232 150 234 157
rect 230 149 236 150
rect 230 145 231 149
rect 235 145 236 149
rect 230 144 236 145
rect 292 136 294 162
rect 319 157 323 158
rect 335 162 339 163
rect 378 162 384 163
rect 407 162 411 163
rect 466 162 472 163
rect 495 162 499 163
rect 554 162 560 163
rect 583 162 587 163
rect 642 162 648 163
rect 663 162 667 163
rect 335 157 339 158
rect 320 150 322 157
rect 318 149 324 150
rect 318 145 319 149
rect 323 145 324 149
rect 318 144 324 145
rect 380 136 382 162
rect 407 157 411 158
rect 408 150 410 157
rect 406 149 412 150
rect 406 145 407 149
rect 411 145 412 149
rect 406 144 412 145
rect 468 136 470 162
rect 495 157 499 158
rect 496 150 498 157
rect 494 149 500 150
rect 494 145 495 149
rect 499 145 500 149
rect 494 144 500 145
rect 556 136 558 162
rect 583 157 587 158
rect 584 150 586 157
rect 582 149 588 150
rect 582 145 583 149
rect 587 145 588 149
rect 582 144 588 145
rect 644 136 646 162
rect 663 157 667 158
rect 671 162 675 163
rect 730 162 736 163
rect 759 162 763 163
rect 671 157 675 158
rect 672 150 674 157
rect 670 149 676 150
rect 670 145 671 149
rect 675 145 676 149
rect 670 144 676 145
rect 732 136 734 162
rect 759 157 763 158
rect 760 150 762 157
rect 758 149 764 150
rect 758 145 759 149
rect 763 145 764 149
rect 758 144 764 145
rect 820 136 822 170
rect 840 163 842 186
rect 914 163 920 164
rect 1002 163 1008 164
rect 1016 163 1018 186
rect 1024 176 1026 262
rect 1112 243 1114 262
rect 1111 242 1115 243
rect 1111 237 1115 238
rect 1112 222 1114 237
rect 1110 221 1116 222
rect 1110 217 1111 221
rect 1115 217 1116 221
rect 1110 216 1116 217
rect 1074 207 1080 208
rect 1074 203 1075 207
rect 1079 203 1080 207
rect 1074 202 1080 203
rect 1110 203 1116 204
rect 1022 175 1028 176
rect 1022 171 1023 175
rect 1027 171 1028 175
rect 1022 170 1028 171
rect 1076 164 1078 202
rect 1110 199 1111 203
rect 1115 199 1116 203
rect 1110 198 1116 199
rect 1074 163 1080 164
rect 1112 163 1114 198
rect 839 162 843 163
rect 839 157 843 158
rect 847 162 851 163
rect 914 159 915 163
rect 919 159 920 163
rect 914 158 920 159
rect 935 162 939 163
rect 1002 159 1003 163
rect 1007 159 1008 163
rect 1002 158 1008 159
rect 1015 162 1019 163
rect 847 157 851 158
rect 848 150 850 157
rect 846 149 852 150
rect 846 145 847 149
rect 851 145 852 149
rect 846 144 852 145
rect 110 132 116 133
rect 202 135 208 136
rect 202 131 203 135
rect 207 131 208 135
rect 202 130 208 131
rect 290 135 296 136
rect 290 131 291 135
rect 295 131 296 135
rect 290 130 296 131
rect 378 135 384 136
rect 378 131 379 135
rect 383 131 384 135
rect 378 130 384 131
rect 466 135 472 136
rect 466 131 467 135
rect 471 131 472 135
rect 466 130 472 131
rect 554 135 560 136
rect 554 131 555 135
rect 559 131 560 135
rect 554 130 560 131
rect 642 135 648 136
rect 642 131 643 135
rect 647 131 648 135
rect 642 130 648 131
rect 730 135 736 136
rect 730 131 731 135
rect 735 131 736 135
rect 730 130 736 131
rect 818 135 824 136
rect 818 131 819 135
rect 823 131 824 135
rect 916 132 918 158
rect 935 157 939 158
rect 936 150 938 157
rect 934 149 940 150
rect 934 145 935 149
rect 939 145 940 149
rect 934 144 940 145
rect 1004 132 1006 158
rect 1015 157 1019 158
rect 1023 162 1027 163
rect 1074 159 1075 163
rect 1079 159 1080 163
rect 1074 158 1080 159
rect 1111 162 1115 163
rect 1023 157 1027 158
rect 1111 157 1115 158
rect 1024 150 1026 157
rect 1022 149 1028 150
rect 1022 145 1023 149
rect 1027 145 1028 149
rect 1022 144 1028 145
rect 1112 138 1114 157
rect 1110 137 1116 138
rect 1110 133 1111 137
rect 1115 133 1116 137
rect 1110 132 1116 133
rect 818 130 824 131
rect 914 131 920 132
rect 914 127 915 131
rect 919 127 920 131
rect 914 126 920 127
rect 1002 131 1008 132
rect 1002 127 1003 131
rect 1007 127 1008 131
rect 1002 126 1008 127
rect 110 119 116 120
rect 110 115 111 119
rect 115 115 116 119
rect 110 114 116 115
rect 1110 119 1116 120
rect 1110 115 1111 119
rect 1115 115 1116 119
rect 1110 114 1116 115
rect 112 99 114 114
rect 134 104 140 105
rect 134 100 135 104
rect 139 100 140 104
rect 134 99 140 100
rect 222 104 228 105
rect 222 100 223 104
rect 227 100 228 104
rect 222 99 228 100
rect 310 104 316 105
rect 310 100 311 104
rect 315 100 316 104
rect 310 99 316 100
rect 398 104 404 105
rect 398 100 399 104
rect 403 100 404 104
rect 398 99 404 100
rect 486 104 492 105
rect 486 100 487 104
rect 491 100 492 104
rect 486 99 492 100
rect 574 104 580 105
rect 574 100 575 104
rect 579 100 580 104
rect 574 99 580 100
rect 662 104 668 105
rect 662 100 663 104
rect 667 100 668 104
rect 662 99 668 100
rect 750 104 756 105
rect 750 100 751 104
rect 755 100 756 104
rect 750 99 756 100
rect 838 104 844 105
rect 838 100 839 104
rect 843 100 844 104
rect 838 99 844 100
rect 926 104 932 105
rect 926 100 927 104
rect 931 100 932 104
rect 926 99 932 100
rect 1014 104 1020 105
rect 1014 100 1015 104
rect 1019 100 1020 104
rect 1014 99 1020 100
rect 1112 99 1114 114
rect 111 98 115 99
rect 111 93 115 94
rect 135 98 139 99
rect 135 93 139 94
rect 223 98 227 99
rect 223 93 227 94
rect 311 98 315 99
rect 311 93 315 94
rect 399 98 403 99
rect 399 93 403 94
rect 487 98 491 99
rect 487 93 491 94
rect 575 98 579 99
rect 575 93 579 94
rect 663 98 667 99
rect 663 93 667 94
rect 751 98 755 99
rect 751 93 755 94
rect 839 98 843 99
rect 839 93 843 94
rect 927 98 931 99
rect 927 93 931 94
rect 1015 98 1019 99
rect 1015 93 1019 94
rect 1111 98 1115 99
rect 1111 93 1115 94
<< m4c >>
rect 111 1202 115 1206
rect 135 1202 139 1206
rect 223 1202 227 1206
rect 311 1202 315 1206
rect 399 1202 403 1206
rect 487 1202 491 1206
rect 575 1202 579 1206
rect 663 1202 667 1206
rect 751 1202 755 1206
rect 1111 1202 1115 1206
rect 111 1126 115 1130
rect 143 1126 147 1130
rect 159 1126 163 1130
rect 231 1126 235 1130
rect 247 1126 251 1130
rect 319 1126 323 1130
rect 335 1126 339 1130
rect 407 1126 411 1130
rect 423 1126 427 1130
rect 495 1126 499 1130
rect 583 1126 587 1130
rect 671 1126 675 1130
rect 759 1126 763 1130
rect 1111 1126 1115 1130
rect 111 1058 115 1062
rect 135 1058 139 1062
rect 151 1058 155 1062
rect 223 1058 227 1062
rect 239 1058 243 1062
rect 171 1003 175 1004
rect 171 1000 175 1003
rect 311 1058 315 1062
rect 327 1058 331 1062
rect 399 1058 403 1062
rect 415 1058 419 1062
rect 1111 1058 1115 1062
rect 379 1000 383 1004
rect 111 990 115 994
rect 143 990 147 994
rect 231 990 235 994
rect 319 990 323 994
rect 407 990 411 994
rect 1111 990 1115 994
rect 111 922 115 926
rect 135 922 139 926
rect 223 922 227 926
rect 311 922 315 926
rect 399 922 403 926
rect 111 854 115 858
rect 143 854 147 858
rect 1111 922 1115 926
rect 231 854 235 858
rect 319 854 323 858
rect 407 854 411 858
rect 495 854 499 858
rect 1111 854 1115 858
rect 111 786 115 790
rect 135 786 139 790
rect 223 786 227 790
rect 231 786 235 790
rect 311 786 315 790
rect 359 786 363 790
rect 399 786 403 790
rect 171 752 175 756
rect 487 786 491 790
rect 503 786 507 790
rect 647 786 651 790
rect 799 786 803 790
rect 959 786 963 790
rect 1111 786 1115 790
rect 111 722 115 726
rect 143 722 147 726
rect 291 736 295 740
rect 239 722 243 726
rect 263 722 267 726
rect 475 752 479 756
rect 359 722 363 726
rect 367 722 371 726
rect 463 722 467 726
rect 511 722 515 726
rect 571 736 575 740
rect 939 736 943 740
rect 575 722 579 726
rect 655 722 659 726
rect 687 722 691 726
rect 799 722 803 726
rect 807 722 811 726
rect 919 722 923 726
rect 995 736 999 740
rect 327 699 331 700
rect 327 696 331 699
rect 387 696 391 700
rect 111 650 115 654
rect 255 650 259 654
rect 351 650 355 654
rect 455 650 459 654
rect 471 650 475 654
rect 567 650 571 654
rect 671 650 675 654
rect 679 650 683 654
rect 783 650 787 654
rect 791 650 795 654
rect 967 722 971 726
rect 1023 722 1027 726
rect 1111 722 1115 726
rect 903 650 907 654
rect 911 650 915 654
rect 1015 650 1019 654
rect 1111 650 1115 654
rect 111 582 115 586
rect 479 582 483 586
rect 495 582 499 586
rect 575 582 579 586
rect 583 582 587 586
rect 671 582 675 586
rect 679 582 683 586
rect 759 582 763 586
rect 791 582 795 586
rect 847 582 851 586
rect 911 582 915 586
rect 935 582 939 586
rect 1023 582 1027 586
rect 1111 582 1115 586
rect 111 514 115 518
rect 375 514 379 518
rect 487 514 491 518
rect 575 514 579 518
rect 599 514 603 518
rect 663 514 667 518
rect 719 514 723 518
rect 751 514 755 518
rect 839 514 843 518
rect 847 514 851 518
rect 927 514 931 518
rect 983 514 987 518
rect 1015 514 1019 518
rect 1111 514 1115 518
rect 411 459 415 460
rect 411 456 415 459
rect 711 456 715 460
rect 111 442 115 446
rect 263 442 267 446
rect 383 442 387 446
rect 391 442 395 446
rect 495 442 499 446
rect 511 442 515 446
rect 607 442 611 446
rect 631 442 635 446
rect 727 442 731 446
rect 751 442 755 446
rect 359 416 363 420
rect 459 416 463 420
rect 111 374 115 378
rect 135 374 139 378
rect 255 374 259 378
rect 383 374 387 378
rect 415 374 419 378
rect 111 306 115 310
rect 143 306 147 310
rect 291 320 295 324
rect 503 374 507 378
rect 583 374 587 378
rect 623 374 627 378
rect 855 442 859 446
rect 879 442 883 446
rect 991 442 995 446
rect 1007 442 1011 446
rect 1111 442 1115 446
rect 743 374 747 378
rect 759 374 763 378
rect 871 374 875 378
rect 935 374 939 378
rect 491 339 495 340
rect 491 336 495 339
rect 619 336 623 340
rect 499 320 503 324
rect 263 306 267 310
rect 271 306 275 310
rect 423 306 427 310
rect 575 306 579 310
rect 591 306 595 310
rect 223 283 227 284
rect 223 280 227 283
rect 299 280 303 284
rect 383 283 387 284
rect 383 280 387 283
rect 451 280 455 284
rect 111 238 115 242
rect 135 238 139 242
rect 175 238 179 242
rect 263 238 267 242
rect 327 238 331 242
rect 415 238 419 242
rect 487 238 491 242
rect 111 158 115 162
rect 143 158 147 162
rect 567 238 571 242
rect 719 306 723 310
rect 767 306 771 310
rect 871 306 875 310
rect 999 374 1003 378
rect 1111 374 1115 378
rect 943 306 947 310
rect 1023 306 1027 310
rect 1111 306 1115 310
rect 655 238 659 242
rect 711 238 715 242
rect 831 238 835 242
rect 863 238 867 242
rect 1007 238 1011 242
rect 1015 238 1019 242
rect 183 158 187 162
rect 231 158 235 162
rect 319 158 323 162
rect 335 158 339 162
rect 407 158 411 162
rect 495 158 499 162
rect 583 158 587 162
rect 663 158 667 162
rect 671 158 675 162
rect 759 158 763 162
rect 1111 238 1115 242
rect 839 158 843 162
rect 847 158 851 162
rect 935 158 939 162
rect 1015 158 1019 162
rect 1023 158 1027 162
rect 1111 158 1115 162
rect 111 94 115 98
rect 135 94 139 98
rect 223 94 227 98
rect 311 94 315 98
rect 399 94 403 98
rect 487 94 491 98
rect 575 94 579 98
rect 663 94 667 98
rect 751 94 755 98
rect 839 94 843 98
rect 927 94 931 98
rect 1015 94 1019 98
rect 1111 94 1115 98
<< m4 >>
rect 84 1201 85 1207
rect 91 1206 1135 1207
rect 91 1202 111 1206
rect 115 1202 135 1206
rect 139 1202 223 1206
rect 227 1202 311 1206
rect 315 1202 399 1206
rect 403 1202 487 1206
rect 491 1202 575 1206
rect 579 1202 663 1206
rect 667 1202 751 1206
rect 755 1202 1111 1206
rect 1115 1202 1135 1206
rect 91 1201 1135 1202
rect 1141 1201 1142 1207
rect 96 1125 97 1131
rect 103 1130 1147 1131
rect 103 1126 111 1130
rect 115 1126 143 1130
rect 147 1126 159 1130
rect 163 1126 231 1130
rect 235 1126 247 1130
rect 251 1126 319 1130
rect 323 1126 335 1130
rect 339 1126 407 1130
rect 411 1126 423 1130
rect 427 1126 495 1130
rect 499 1126 583 1130
rect 587 1126 671 1130
rect 675 1126 759 1130
rect 763 1126 1111 1130
rect 1115 1126 1147 1130
rect 103 1125 1147 1126
rect 1153 1125 1154 1131
rect 84 1057 85 1063
rect 91 1062 1135 1063
rect 91 1058 111 1062
rect 115 1058 135 1062
rect 139 1058 151 1062
rect 155 1058 223 1062
rect 227 1058 239 1062
rect 243 1058 311 1062
rect 315 1058 327 1062
rect 331 1058 399 1062
rect 403 1058 415 1062
rect 419 1058 1111 1062
rect 1115 1058 1135 1062
rect 91 1057 1135 1058
rect 1141 1057 1142 1063
rect 170 1004 176 1005
rect 378 1004 384 1005
rect 170 1000 171 1004
rect 175 1000 379 1004
rect 383 1000 384 1004
rect 170 999 176 1000
rect 378 999 384 1000
rect 96 989 97 995
rect 103 994 1147 995
rect 103 990 111 994
rect 115 990 143 994
rect 147 990 231 994
rect 235 990 319 994
rect 323 990 407 994
rect 411 990 1111 994
rect 1115 990 1147 994
rect 103 989 1147 990
rect 1153 989 1154 995
rect 84 921 85 927
rect 91 926 1135 927
rect 91 922 111 926
rect 115 922 135 926
rect 139 922 223 926
rect 227 922 311 926
rect 315 922 399 926
rect 403 922 1111 926
rect 1115 922 1135 926
rect 91 921 1135 922
rect 1141 921 1142 927
rect 96 853 97 859
rect 103 858 1147 859
rect 103 854 111 858
rect 115 854 143 858
rect 147 854 231 858
rect 235 854 319 858
rect 323 854 407 858
rect 411 854 495 858
rect 499 854 1111 858
rect 1115 854 1147 858
rect 103 853 1147 854
rect 1153 853 1154 859
rect 84 785 85 791
rect 91 790 1135 791
rect 91 786 111 790
rect 115 786 135 790
rect 139 786 223 790
rect 227 786 231 790
rect 235 786 311 790
rect 315 786 359 790
rect 363 786 399 790
rect 403 786 487 790
rect 491 786 503 790
rect 507 786 647 790
rect 651 786 799 790
rect 803 786 959 790
rect 963 786 1111 790
rect 1115 786 1135 790
rect 91 785 1135 786
rect 1141 785 1142 791
rect 170 756 176 757
rect 474 756 480 757
rect 170 752 171 756
rect 175 752 475 756
rect 479 752 480 756
rect 170 751 176 752
rect 474 751 480 752
rect 290 740 296 741
rect 570 740 576 741
rect 290 736 291 740
rect 295 736 571 740
rect 575 736 576 740
rect 290 735 296 736
rect 570 735 576 736
rect 938 740 944 741
rect 994 740 1000 741
rect 938 736 939 740
rect 943 736 995 740
rect 999 736 1000 740
rect 938 735 944 736
rect 994 735 1000 736
rect 96 721 97 727
rect 103 726 1147 727
rect 103 722 111 726
rect 115 722 143 726
rect 147 722 239 726
rect 243 722 263 726
rect 267 722 359 726
rect 363 722 367 726
rect 371 722 463 726
rect 467 722 511 726
rect 515 722 575 726
rect 579 722 655 726
rect 659 722 687 726
rect 691 722 799 726
rect 803 722 807 726
rect 811 722 919 726
rect 923 722 967 726
rect 971 722 1023 726
rect 1027 722 1111 726
rect 1115 722 1147 726
rect 103 721 1147 722
rect 1153 721 1154 727
rect 326 700 332 701
rect 386 700 392 701
rect 326 696 327 700
rect 331 696 387 700
rect 391 696 392 700
rect 326 695 332 696
rect 386 695 392 696
rect 84 649 85 655
rect 91 654 1135 655
rect 91 650 111 654
rect 115 650 255 654
rect 259 650 351 654
rect 355 650 455 654
rect 459 650 471 654
rect 475 650 567 654
rect 571 650 671 654
rect 675 650 679 654
rect 683 650 783 654
rect 787 650 791 654
rect 795 650 903 654
rect 907 650 911 654
rect 915 650 1015 654
rect 1019 650 1111 654
rect 1115 650 1135 654
rect 91 649 1135 650
rect 1141 649 1142 655
rect 96 581 97 587
rect 103 586 1147 587
rect 103 582 111 586
rect 115 582 479 586
rect 483 582 495 586
rect 499 582 575 586
rect 579 582 583 586
rect 587 582 671 586
rect 675 582 679 586
rect 683 582 759 586
rect 763 582 791 586
rect 795 582 847 586
rect 851 582 911 586
rect 915 582 935 586
rect 939 582 1023 586
rect 1027 582 1111 586
rect 1115 582 1147 586
rect 103 581 1147 582
rect 1153 581 1154 587
rect 84 513 85 519
rect 91 518 1135 519
rect 91 514 111 518
rect 115 514 375 518
rect 379 514 487 518
rect 491 514 575 518
rect 579 514 599 518
rect 603 514 663 518
rect 667 514 719 518
rect 723 514 751 518
rect 755 514 839 518
rect 843 514 847 518
rect 851 514 927 518
rect 931 514 983 518
rect 987 514 1015 518
rect 1019 514 1111 518
rect 1115 514 1135 518
rect 91 513 1135 514
rect 1141 513 1142 519
rect 410 460 416 461
rect 710 460 716 461
rect 410 456 411 460
rect 415 456 711 460
rect 715 456 716 460
rect 410 455 416 456
rect 710 455 716 456
rect 96 441 97 447
rect 103 446 1147 447
rect 103 442 111 446
rect 115 442 263 446
rect 267 442 383 446
rect 387 442 391 446
rect 395 442 495 446
rect 499 442 511 446
rect 515 442 607 446
rect 611 442 631 446
rect 635 442 727 446
rect 731 442 751 446
rect 755 442 855 446
rect 859 442 879 446
rect 883 442 991 446
rect 995 442 1007 446
rect 1011 442 1111 446
rect 1115 442 1147 446
rect 103 441 1147 442
rect 1153 441 1154 447
rect 358 420 364 421
rect 458 420 464 421
rect 358 416 359 420
rect 363 416 459 420
rect 463 416 464 420
rect 358 415 364 416
rect 458 415 464 416
rect 84 373 85 379
rect 91 378 1135 379
rect 91 374 111 378
rect 115 374 135 378
rect 139 374 255 378
rect 259 374 383 378
rect 387 374 415 378
rect 419 374 503 378
rect 507 374 583 378
rect 587 374 623 378
rect 627 374 743 378
rect 747 374 759 378
rect 763 374 871 378
rect 875 374 935 378
rect 939 374 999 378
rect 1003 374 1111 378
rect 1115 374 1135 378
rect 91 373 1135 374
rect 1141 373 1142 379
rect 490 340 496 341
rect 618 340 624 341
rect 490 336 491 340
rect 495 336 619 340
rect 623 336 624 340
rect 490 335 496 336
rect 618 335 624 336
rect 290 324 296 325
rect 498 324 504 325
rect 290 320 291 324
rect 295 320 499 324
rect 503 320 504 324
rect 290 319 296 320
rect 498 319 504 320
rect 96 305 97 311
rect 103 310 1147 311
rect 103 306 111 310
rect 115 306 143 310
rect 147 306 263 310
rect 267 306 271 310
rect 275 306 423 310
rect 427 306 575 310
rect 579 306 591 310
rect 595 306 719 310
rect 723 306 767 310
rect 771 306 871 310
rect 875 306 943 310
rect 947 306 1023 310
rect 1027 306 1111 310
rect 1115 306 1147 310
rect 103 305 1147 306
rect 1153 305 1154 311
rect 222 284 228 285
rect 298 284 304 285
rect 222 280 223 284
rect 227 280 299 284
rect 303 280 304 284
rect 222 279 228 280
rect 298 279 304 280
rect 382 284 388 285
rect 450 284 456 285
rect 382 280 383 284
rect 387 280 451 284
rect 455 280 456 284
rect 382 279 388 280
rect 450 279 456 280
rect 84 237 85 243
rect 91 242 1135 243
rect 91 238 111 242
rect 115 238 135 242
rect 139 238 175 242
rect 179 238 263 242
rect 267 238 327 242
rect 331 238 415 242
rect 419 238 487 242
rect 491 238 567 242
rect 571 238 655 242
rect 659 238 711 242
rect 715 238 831 242
rect 835 238 863 242
rect 867 238 1007 242
rect 1011 238 1015 242
rect 1019 238 1111 242
rect 1115 238 1135 242
rect 91 237 1135 238
rect 1141 237 1142 243
rect 96 157 97 163
rect 103 162 1147 163
rect 103 158 111 162
rect 115 158 143 162
rect 147 158 183 162
rect 187 158 231 162
rect 235 158 319 162
rect 323 158 335 162
rect 339 158 407 162
rect 411 158 495 162
rect 499 158 583 162
rect 587 158 663 162
rect 667 158 671 162
rect 675 158 759 162
rect 763 158 839 162
rect 843 158 847 162
rect 851 158 935 162
rect 939 158 1015 162
rect 1019 158 1023 162
rect 1027 158 1111 162
rect 1115 158 1147 162
rect 103 157 1147 158
rect 1153 157 1154 163
rect 84 93 85 99
rect 91 98 1135 99
rect 91 94 111 98
rect 115 94 135 98
rect 139 94 223 98
rect 227 94 311 98
rect 315 94 399 98
rect 403 94 487 98
rect 491 94 575 98
rect 579 94 663 98
rect 667 94 751 98
rect 755 94 839 98
rect 843 94 927 98
rect 931 94 1015 98
rect 1019 94 1111 98
rect 1115 94 1135 98
rect 91 93 1135 94
rect 1141 93 1142 99
<< m5c >>
rect 85 1201 91 1207
rect 1135 1201 1141 1207
rect 97 1125 103 1131
rect 1147 1125 1153 1131
rect 85 1057 91 1063
rect 1135 1057 1141 1063
rect 97 989 103 995
rect 1147 989 1153 995
rect 85 921 91 927
rect 1135 921 1141 927
rect 97 853 103 859
rect 1147 853 1153 859
rect 85 785 91 791
rect 1135 785 1141 791
rect 97 721 103 727
rect 1147 721 1153 727
rect 85 649 91 655
rect 1135 649 1141 655
rect 97 581 103 587
rect 1147 581 1153 587
rect 85 513 91 519
rect 1135 513 1141 519
rect 97 441 103 447
rect 1147 441 1153 447
rect 85 373 91 379
rect 1135 373 1141 379
rect 97 305 103 311
rect 1147 305 1153 311
rect 85 237 91 243
rect 1135 237 1141 243
rect 97 157 103 163
rect 1147 157 1153 163
rect 85 93 91 99
rect 1135 93 1141 99
<< m5 >>
rect 84 1207 92 1224
rect 84 1201 85 1207
rect 91 1201 92 1207
rect 84 1063 92 1201
rect 84 1057 85 1063
rect 91 1057 92 1063
rect 84 927 92 1057
rect 84 921 85 927
rect 91 921 92 927
rect 84 791 92 921
rect 84 785 85 791
rect 91 785 92 791
rect 84 655 92 785
rect 84 649 85 655
rect 91 649 92 655
rect 84 519 92 649
rect 84 513 85 519
rect 91 513 92 519
rect 84 379 92 513
rect 84 373 85 379
rect 91 373 92 379
rect 84 243 92 373
rect 84 237 85 243
rect 91 237 92 243
rect 84 99 92 237
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 1131 104 1224
rect 96 1125 97 1131
rect 103 1125 104 1131
rect 96 995 104 1125
rect 96 989 97 995
rect 103 989 104 995
rect 96 859 104 989
rect 96 853 97 859
rect 103 853 104 859
rect 96 727 104 853
rect 96 721 97 727
rect 103 721 104 727
rect 96 587 104 721
rect 96 581 97 587
rect 103 581 104 587
rect 96 447 104 581
rect 96 441 97 447
rect 103 441 104 447
rect 96 311 104 441
rect 96 305 97 311
rect 103 305 104 311
rect 96 163 104 305
rect 96 157 97 163
rect 103 157 104 163
rect 96 72 104 157
rect 1134 1207 1142 1224
rect 1134 1201 1135 1207
rect 1141 1201 1142 1207
rect 1134 1063 1142 1201
rect 1134 1057 1135 1063
rect 1141 1057 1142 1063
rect 1134 927 1142 1057
rect 1134 921 1135 927
rect 1141 921 1142 927
rect 1134 791 1142 921
rect 1134 785 1135 791
rect 1141 785 1142 791
rect 1134 655 1142 785
rect 1134 649 1135 655
rect 1141 649 1142 655
rect 1134 519 1142 649
rect 1134 513 1135 519
rect 1141 513 1142 519
rect 1134 379 1142 513
rect 1134 373 1135 379
rect 1141 373 1142 379
rect 1134 243 1142 373
rect 1134 237 1135 243
rect 1141 237 1142 243
rect 1134 99 1142 237
rect 1134 93 1135 99
rect 1141 93 1142 99
rect 1134 72 1142 93
rect 1146 1131 1154 1224
rect 1146 1125 1147 1131
rect 1153 1125 1154 1131
rect 1146 995 1154 1125
rect 1146 989 1147 995
rect 1153 989 1154 995
rect 1146 859 1154 989
rect 1146 853 1147 859
rect 1153 853 1154 859
rect 1146 727 1154 853
rect 1146 721 1147 727
rect 1153 721 1154 727
rect 1146 587 1154 721
rect 1146 581 1147 587
rect 1153 581 1154 587
rect 1146 447 1154 581
rect 1146 441 1147 447
rect 1153 441 1154 447
rect 1146 311 1154 441
rect 1146 305 1147 311
rect 1153 305 1154 311
rect 1146 163 1154 305
rect 1146 157 1147 163
rect 1153 157 1154 163
rect 1146 72 1154 157
use _0_0std_0_0cells_0_0MUX2X1  mux_564_6
timestamp 1731001196
transform 1 0 128 0 1 96
box 8 2 80 63
use welltap_svt  __well_tap__0
timestamp 1731001196
transform 1 0 104 0 1 112
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0MUX2X1  mux_564_6
timestamp 1731001196
transform 1 0 128 0 1 96
box 8 2 80 63
use welltap_svt  __well_tap__0
timestamp 1731001196
transform 1 0 104 0 1 112
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0MUX2X1  mux_565_6
timestamp 1731001196
transform 1 0 216 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_565_6
timestamp 1731001196
transform 1 0 216 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_566_6
timestamp 1731001196
transform 1 0 304 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_566_6
timestamp 1731001196
transform 1 0 304 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_567_6
timestamp 1731001196
transform 1 0 392 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_567_6
timestamp 1731001196
transform 1 0 392 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_568_6
timestamp 1731001196
transform 1 0 480 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_568_6
timestamp 1731001196
transform 1 0 480 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_569_6
timestamp 1731001196
transform 1 0 568 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_569_6
timestamp 1731001196
transform 1 0 568 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_570_6
timestamp 1731001196
transform 1 0 656 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_570_6
timestamp 1731001196
transform 1 0 656 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_571_6
timestamp 1731001196
transform 1 0 744 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_571_6
timestamp 1731001196
transform 1 0 744 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_599_6
timestamp 1731001196
transform 1 0 832 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_599_6
timestamp 1731001196
transform 1 0 832 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_598_6
timestamp 1731001196
transform 1 0 920 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_598_6
timestamp 1731001196
transform 1 0 920 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_597_6
timestamp 1731001196
transform 1 0 1008 0 1 96
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_597_6
timestamp 1731001196
transform 1 0 1008 0 1 96
box 8 2 80 63
use welltap_svt  __well_tap__1
timestamp 1731001196
transform 1 0 1104 0 1 112
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1731001196
transform 1 0 1104 0 1 112
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1731001196
transform 1 0 104 0 -1 224
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1731001196
transform 1 0 104 0 -1 224
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_563_6
timestamp 1731001196
transform 1 0 168 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_563_6
timestamp 1731001196
transform 1 0 168 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_562_6
timestamp 1731001196
transform 1 0 320 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_562_6
timestamp 1731001196
transform 1 0 320 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_561_6
timestamp 1731001196
transform 1 0 480 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_561_6
timestamp 1731001196
transform 1 0 480 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_573_6
timestamp 1731001196
transform 1 0 648 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_573_6
timestamp 1731001196
transform 1 0 648 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_572_6
timestamp 1731001196
transform 1 0 824 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_572_6
timestamp 1731001196
transform 1 0 824 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_596_6
timestamp 1731001196
transform 1 0 1000 0 -1 240
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_596_6
timestamp 1731001196
transform 1 0 1000 0 -1 240
box 8 2 80 63
use welltap_svt  __well_tap__3
timestamp 1731001196
transform 1 0 1104 0 -1 224
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1731001196
transform 1 0 1104 0 -1 224
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_558_6
timestamp 1731001196
transform 1 0 128 0 1 244
box 8 2 80 63
use welltap_svt  __well_tap__4
timestamp 1731001196
transform 1 0 104 0 1 260
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_558_6
timestamp 1731001196
transform 1 0 128 0 1 244
box 8 2 80 63
use welltap_svt  __well_tap__4
timestamp 1731001196
transform 1 0 104 0 1 260
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_559_6
timestamp 1731001196
transform 1 0 256 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_559_6
timestamp 1731001196
transform 1 0 256 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_560_6
timestamp 1731001196
transform 1 0 408 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_560_6
timestamp 1731001196
transform 1 0 408 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_574_6
timestamp 1731001196
transform 1 0 560 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_574_6
timestamp 1731001196
transform 1 0 560 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_575_6
timestamp 1731001196
transform 1 0 704 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_575_6
timestamp 1731001196
transform 1 0 704 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_594_6
timestamp 1731001196
transform 1 0 856 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_594_6
timestamp 1731001196
transform 1 0 856 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_595_6
timestamp 1731001196
transform 1 0 1008 0 1 244
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_595_6
timestamp 1731001196
transform 1 0 1008 0 1 244
box 8 2 80 63
use welltap_svt  __well_tap__5
timestamp 1731001196
transform 1 0 1104 0 1 260
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1731001196
transform 1 0 1104 0 1 260
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_557_6
timestamp 1731001196
transform 1 0 128 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_557_6
timestamp 1731001196
transform 1 0 128 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_556_6
timestamp 1731001196
transform 1 0 248 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_556_6
timestamp 1731001196
transform 1 0 248 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_554_6
timestamp 1731001196
transform 1 0 408 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_554_6
timestamp 1731001196
transform 1 0 408 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_555_6
timestamp 1731001196
transform 1 0 576 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_555_6
timestamp 1731001196
transform 1 0 576 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_576_6
timestamp 1731001196
transform 1 0 752 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_576_6
timestamp 1731001196
transform 1 0 752 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_593_6
timestamp 1731001196
transform 1 0 928 0 -1 376
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_593_6
timestamp 1731001196
transform 1 0 928 0 -1 376
box 8 2 80 63
use welltap_svt  __well_tap__6
timestamp 1731001196
transform 1 0 104 0 -1 360
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1731001196
transform 1 0 104 0 1 396
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1731001196
transform 1 0 104 0 -1 360
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1731001196
transform 1 0 104 0 1 396
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_552_6
timestamp 1731001196
transform 1 0 248 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_552_6
timestamp 1731001196
transform 1 0 248 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_553_6
timestamp 1731001196
transform 1 0 376 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_553_6
timestamp 1731001196
transform 1 0 376 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_551_6
timestamp 1731001196
transform 1 0 496 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_551_6
timestamp 1731001196
transform 1 0 496 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_577_6
timestamp 1731001196
transform 1 0 616 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_577_6
timestamp 1731001196
transform 1 0 616 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_578_6
timestamp 1731001196
transform 1 0 736 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_578_6
timestamp 1731001196
transform 1 0 736 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_592_6
timestamp 1731001196
transform 1 0 864 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_592_6
timestamp 1731001196
transform 1 0 864 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_591_6
timestamp 1731001196
transform 1 0 992 0 1 380
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_591_6
timestamp 1731001196
transform 1 0 992 0 1 380
box 8 2 80 63
use welltap_svt  __well_tap__7
timestamp 1731001196
transform 1 0 1104 0 -1 360
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1731001196
transform 1 0 1104 0 1 396
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1731001196
transform 1 0 1104 0 -1 360
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1731001196
transform 1 0 1104 0 1 396
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_549_6
timestamp 1731001196
transform 1 0 368 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_549_6
timestamp 1731001196
transform 1 0 368 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_550_6
timestamp 1731001196
transform 1 0 480 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_550_6
timestamp 1731001196
transform 1 0 480 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_547_6
timestamp 1731001196
transform 1 0 592 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_547_6
timestamp 1731001196
transform 1 0 592 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_548_6
timestamp 1731001196
transform 1 0 712 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_548_6
timestamp 1731001196
transform 1 0 712 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_579_6
timestamp 1731001196
transform 1 0 840 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_579_6
timestamp 1731001196
transform 1 0 840 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_590_6
timestamp 1731001196
transform 1 0 976 0 -1 516
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_590_6
timestamp 1731001196
transform 1 0 976 0 -1 516
box 8 2 80 63
use welltap_svt  __well_tap__10
timestamp 1731001196
transform 1 0 104 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1731001196
transform 1 0 104 0 -1 500
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_546_6
timestamp 1731001196
transform 1 0 480 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_546_6
timestamp 1731001196
transform 1 0 480 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_545_6
timestamp 1731001196
transform 1 0 568 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_545_6
timestamp 1731001196
transform 1 0 568 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_544_6
timestamp 1731001196
transform 1 0 656 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_544_6
timestamp 1731001196
transform 1 0 656 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_543_6
timestamp 1731001196
transform 1 0 744 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_543_6
timestamp 1731001196
transform 1 0 744 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_580_6
timestamp 1731001196
transform 1 0 832 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_580_6
timestamp 1731001196
transform 1 0 832 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_589_6
timestamp 1731001196
transform 1 0 920 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_589_6
timestamp 1731001196
transform 1 0 920 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_588_6
timestamp 1731001196
transform 1 0 1008 0 1 520
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_588_6
timestamp 1731001196
transform 1 0 1008 0 1 520
box 8 2 80 63
use welltap_svt  __well_tap__11
timestamp 1731001196
transform 1 0 1104 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1731001196
transform 1 0 1104 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1731001196
transform 1 0 104 0 1 536
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1731001196
transform 1 0 104 0 1 536
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_539_6
timestamp 1731001196
transform 1 0 464 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_539_6
timestamp 1731001196
transform 1 0 464 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_540_6
timestamp 1731001196
transform 1 0 560 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_540_6
timestamp 1731001196
transform 1 0 560 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_541_6
timestamp 1731001196
transform 1 0 664 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_541_6
timestamp 1731001196
transform 1 0 664 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_542_6
timestamp 1731001196
transform 1 0 776 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_542_6
timestamp 1731001196
transform 1 0 776 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_581_6
timestamp 1731001196
transform 1 0 896 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_581_6
timestamp 1731001196
transform 1 0 896 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_587_6
timestamp 1731001196
transform 1 0 1008 0 -1 652
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_587_6
timestamp 1731001196
transform 1 0 1008 0 -1 652
box 8 2 80 63
use welltap_svt  __well_tap__13
timestamp 1731001196
transform 1 0 1104 0 1 536
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1731001196
transform 1 0 1104 0 1 536
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1731001196
transform 1 0 104 0 -1 636
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1731001196
transform 1 0 104 0 -1 636
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_534_6
timestamp 1731001196
transform 1 0 248 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_534_6
timestamp 1731001196
transform 1 0 248 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_535_6
timestamp 1731001196
transform 1 0 344 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_535_6
timestamp 1731001196
transform 1 0 344 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_536_6
timestamp 1731001196
transform 1 0 448 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_536_6
timestamp 1731001196
transform 1 0 448 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_537_6
timestamp 1731001196
transform 1 0 560 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_537_6
timestamp 1731001196
transform 1 0 560 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_538_6
timestamp 1731001196
transform 1 0 672 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_538_6
timestamp 1731001196
transform 1 0 672 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_582_6
timestamp 1731001196
transform 1 0 784 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_582_6
timestamp 1731001196
transform 1 0 784 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_585_6
timestamp 1731001196
transform 1 0 904 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_585_6
timestamp 1731001196
transform 1 0 904 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_586_6
timestamp 1731001196
transform 1 0 1008 0 1 660
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_586_6
timestamp 1731001196
transform 1 0 1008 0 1 660
box 8 2 80 63
use welltap_svt  __well_tap__15
timestamp 1731001196
transform 1 0 1104 0 -1 636
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1731001196
transform 1 0 1104 0 -1 636
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_529_6
timestamp 1731001196
transform 1 0 128 0 -1 788
box 8 2 80 63
use welltap_svt  __well_tap__16
timestamp 1731001196
transform 1 0 104 0 1 676
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_529_6
timestamp 1731001196
transform 1 0 128 0 -1 788
box 8 2 80 63
use welltap_svt  __well_tap__16
timestamp 1731001196
transform 1 0 104 0 1 676
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_530_6
timestamp 1731001196
transform 1 0 224 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_530_6
timestamp 1731001196
transform 1 0 224 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_531_6
timestamp 1731001196
transform 1 0 352 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_531_6
timestamp 1731001196
transform 1 0 352 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_532_6
timestamp 1731001196
transform 1 0 496 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_532_6
timestamp 1731001196
transform 1 0 496 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_533_6
timestamp 1731001196
transform 1 0 640 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_533_6
timestamp 1731001196
transform 1 0 640 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_583_6
timestamp 1731001196
transform 1 0 792 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_583_6
timestamp 1731001196
transform 1 0 792 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_584_6
timestamp 1731001196
transform 1 0 952 0 -1 788
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_584_6
timestamp 1731001196
transform 1 0 952 0 -1 788
box 8 2 80 63
use welltap_svt  __well_tap__17
timestamp 1731001196
transform 1 0 1104 0 1 676
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1731001196
transform 1 0 1104 0 1 676
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_524_6
timestamp 1731001196
transform 1 0 128 0 1 792
box 8 2 80 63
use welltap_svt  __well_tap__18
timestamp 1731001196
transform 1 0 104 0 -1 772
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_524_6
timestamp 1731001196
transform 1 0 128 0 1 792
box 8 2 80 63
use welltap_svt  __well_tap__18
timestamp 1731001196
transform 1 0 104 0 -1 772
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_525_6
timestamp 1731001196
transform 1 0 216 0 1 792
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_525_6
timestamp 1731001196
transform 1 0 216 0 1 792
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_526_6
timestamp 1731001196
transform 1 0 304 0 1 792
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_526_6
timestamp 1731001196
transform 1 0 304 0 1 792
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_527_6
timestamp 1731001196
transform 1 0 392 0 1 792
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_527_6
timestamp 1731001196
transform 1 0 392 0 1 792
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_528_6
timestamp 1731001196
transform 1 0 480 0 1 792
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_528_6
timestamp 1731001196
transform 1 0 480 0 1 792
box 8 2 80 63
use welltap_svt  __well_tap__19
timestamp 1731001196
transform 1 0 1104 0 -1 772
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1731001196
transform 1 0 1104 0 -1 772
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_523_6
timestamp 1731001196
transform 1 0 128 0 -1 924
box 8 2 80 63
use welltap_svt  __well_tap__20
timestamp 1731001196
transform 1 0 104 0 1 808
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_523_6
timestamp 1731001196
transform 1 0 128 0 -1 924
box 8 2 80 63
use welltap_svt  __well_tap__20
timestamp 1731001196
transform 1 0 104 0 1 808
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_522_6
timestamp 1731001196
transform 1 0 216 0 -1 924
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_522_6
timestamp 1731001196
transform 1 0 216 0 -1 924
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_521_6
timestamp 1731001196
transform 1 0 304 0 -1 924
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_521_6
timestamp 1731001196
transform 1 0 304 0 -1 924
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_520_6
timestamp 1731001196
transform 1 0 392 0 -1 924
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_520_6
timestamp 1731001196
transform 1 0 392 0 -1 924
box 8 2 80 63
use welltap_svt  __well_tap__21
timestamp 1731001196
transform 1 0 1104 0 1 808
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1731001196
transform 1 0 1104 0 1 808
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1731001196
transform 1 0 104 0 -1 908
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1731001196
transform 1 0 104 0 -1 908
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1731001196
transform 1 0 1104 0 -1 908
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1731001196
transform 1 0 1104 0 -1 908
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_516_6
timestamp 1731001196
transform 1 0 128 0 1 928
box 8 2 80 63
use welltap_svt  __well_tap__24
timestamp 1731001196
transform 1 0 104 0 1 944
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_516_6
timestamp 1731001196
transform 1 0 128 0 1 928
box 8 2 80 63
use welltap_svt  __well_tap__24
timestamp 1731001196
transform 1 0 104 0 1 944
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_517_6
timestamp 1731001196
transform 1 0 216 0 1 928
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_517_6
timestamp 1731001196
transform 1 0 216 0 1 928
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_518_6
timestamp 1731001196
transform 1 0 304 0 1 928
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_518_6
timestamp 1731001196
transform 1 0 304 0 1 928
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_519_6
timestamp 1731001196
transform 1 0 392 0 1 928
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_519_6
timestamp 1731001196
transform 1 0 392 0 1 928
box 8 2 80 63
use welltap_svt  __well_tap__25
timestamp 1731001196
transform 1 0 1104 0 1 944
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1731001196
transform 1 0 1104 0 1 944
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_515_6
timestamp 1731001196
transform 1 0 128 0 -1 1060
box 8 2 80 63
use welltap_svt  __well_tap__26
timestamp 1731001196
transform 1 0 104 0 -1 1044
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_515_6
timestamp 1731001196
transform 1 0 128 0 -1 1060
box 8 2 80 63
use welltap_svt  __well_tap__26
timestamp 1731001196
transform 1 0 104 0 -1 1044
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_512_6
timestamp 1731001196
transform 1 0 216 0 -1 1060
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_512_6
timestamp 1731001196
transform 1 0 216 0 -1 1060
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_513_6
timestamp 1731001196
transform 1 0 304 0 -1 1060
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_513_6
timestamp 1731001196
transform 1 0 304 0 -1 1060
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_514_6
timestamp 1731001196
transform 1 0 392 0 -1 1060
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_514_6
timestamp 1731001196
transform 1 0 392 0 -1 1060
box 8 2 80 63
use welltap_svt  __well_tap__27
timestamp 1731001196
transform 1 0 1104 0 -1 1044
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1731001196
transform 1 0 1104 0 -1 1044
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_511_6
timestamp 1731001196
transform 1 0 144 0 1 1064
box 8 2 80 63
use welltap_svt  __well_tap__28
timestamp 1731001196
transform 1 0 104 0 1 1080
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_511_6
timestamp 1731001196
transform 1 0 144 0 1 1064
box 8 2 80 63
use welltap_svt  __well_tap__28
timestamp 1731001196
transform 1 0 104 0 1 1080
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_510_6
timestamp 1731001196
transform 1 0 232 0 1 1064
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_510_6
timestamp 1731001196
transform 1 0 232 0 1 1064
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_59_6
timestamp 1731001196
transform 1 0 320 0 1 1064
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_59_6
timestamp 1731001196
transform 1 0 320 0 1 1064
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_58_6
timestamp 1731001196
transform 1 0 408 0 1 1064
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_58_6
timestamp 1731001196
transform 1 0 408 0 1 1064
box 8 2 80 63
use welltap_svt  __well_tap__29
timestamp 1731001196
transform 1 0 1104 0 1 1080
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1731001196
transform 1 0 1104 0 1 1080
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_50_6
timestamp 1731001196
transform 1 0 128 0 -1 1204
box 8 2 80 63
use welltap_svt  __well_tap__30
timestamp 1731001196
transform 1 0 104 0 -1 1188
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_50_6
timestamp 1731001196
transform 1 0 128 0 -1 1204
box 8 2 80 63
use welltap_svt  __well_tap__30
timestamp 1731001196
transform 1 0 104 0 -1 1188
box 8 4 12 24
use _0_0std_0_0cells_0_0MUX2X1  mux_51_6
timestamp 1731001196
transform 1 0 216 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_51_6
timestamp 1731001196
transform 1 0 216 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_52_6
timestamp 1731001196
transform 1 0 304 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_52_6
timestamp 1731001196
transform 1 0 304 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_53_6
timestamp 1731001196
transform 1 0 392 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_53_6
timestamp 1731001196
transform 1 0 392 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_57_6
timestamp 1731001196
transform 1 0 480 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_57_6
timestamp 1731001196
transform 1 0 480 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_54_6
timestamp 1731001196
transform 1 0 568 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_54_6
timestamp 1731001196
transform 1 0 568 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_55_6
timestamp 1731001196
transform 1 0 656 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_55_6
timestamp 1731001196
transform 1 0 656 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_56_6
timestamp 1731001196
transform 1 0 744 0 -1 1204
box 8 2 80 63
use _0_0std_0_0cells_0_0MUX2X1  mux_56_6
timestamp 1731001196
transform 1 0 744 0 -1 1204
box 8 2 80 63
use welltap_svt  __well_tap__31
timestamp 1731001196
transform 1 0 1104 0 -1 1188
box 8 4 12 24
use welltap_svt  __well_tap__31
timestamp 1731001196
transform 1 0 1104 0 -1 1188
box 8 4 12 24
<< end >>
