magic
tech sky130l
timestamp 1731220307
<< m1 >>
rect 638 1796 642 1800
rect 1190 1796 1194 1800
rect 80 1666 84 1670
rect 1748 1606 1752 1610
rect 80 1534 84 1538
rect 1748 1414 1752 1418
rect 80 1398 84 1402
rect 80 1266 84 1270
rect 1748 1222 1752 1226
rect 80 1134 84 1138
rect 1748 1030 1752 1034
rect 80 1002 84 1006
rect 80 866 84 870
rect 1748 838 1752 842
rect 80 734 84 738
rect 1748 646 1752 650
rect 80 602 84 606
rect 80 470 84 474
rect 1748 454 1752 458
rect 80 334 84 338
rect 1748 262 1752 266
rect 80 202 84 206
rect 638 72 642 76
rect 1190 72 1194 76
<< m2 >>
rect 150 1755 156 1756
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 150 1751 151 1755
rect 155 1751 156 1755
rect 150 1750 156 1751
rect 182 1755 188 1756
rect 182 1751 183 1755
rect 187 1751 188 1755
rect 182 1750 188 1751
rect 214 1755 220 1756
rect 214 1751 215 1755
rect 219 1751 220 1755
rect 214 1750 220 1751
rect 246 1755 252 1756
rect 246 1751 247 1755
rect 251 1751 252 1755
rect 246 1750 252 1751
rect 278 1755 284 1756
rect 278 1751 279 1755
rect 283 1751 284 1755
rect 278 1750 284 1751
rect 310 1755 316 1756
rect 310 1751 311 1755
rect 315 1751 316 1755
rect 310 1750 316 1751
rect 342 1755 348 1756
rect 342 1751 343 1755
rect 347 1751 348 1755
rect 342 1750 348 1751
rect 374 1755 380 1756
rect 374 1751 375 1755
rect 379 1751 380 1755
rect 374 1750 380 1751
rect 406 1755 412 1756
rect 406 1751 407 1755
rect 411 1751 412 1755
rect 406 1750 412 1751
rect 438 1755 444 1756
rect 438 1751 439 1755
rect 443 1751 444 1755
rect 438 1750 444 1751
rect 470 1755 476 1756
rect 470 1751 471 1755
rect 475 1751 476 1755
rect 470 1750 476 1751
rect 502 1755 508 1756
rect 502 1751 503 1755
rect 507 1751 508 1755
rect 502 1750 508 1751
rect 534 1755 540 1756
rect 534 1751 535 1755
rect 539 1751 540 1755
rect 534 1750 540 1751
rect 566 1755 572 1756
rect 566 1751 567 1755
rect 571 1751 572 1755
rect 566 1750 572 1751
rect 598 1755 604 1756
rect 598 1751 599 1755
rect 603 1751 604 1755
rect 598 1750 604 1751
rect 630 1755 636 1756
rect 630 1751 631 1755
rect 635 1751 636 1755
rect 630 1750 636 1751
rect 662 1755 668 1756
rect 662 1751 663 1755
rect 667 1751 668 1755
rect 662 1750 668 1751
rect 694 1755 700 1756
rect 694 1751 695 1755
rect 699 1751 700 1755
rect 694 1750 700 1751
rect 726 1755 732 1756
rect 726 1751 727 1755
rect 731 1751 732 1755
rect 726 1750 732 1751
rect 758 1755 764 1756
rect 758 1751 759 1755
rect 763 1751 764 1755
rect 758 1750 764 1751
rect 790 1755 796 1756
rect 790 1751 791 1755
rect 795 1751 796 1755
rect 790 1750 796 1751
rect 822 1755 828 1756
rect 822 1751 823 1755
rect 827 1751 828 1755
rect 822 1750 828 1751
rect 854 1755 860 1756
rect 854 1751 855 1755
rect 859 1751 860 1755
rect 854 1750 860 1751
rect 886 1755 892 1756
rect 886 1751 887 1755
rect 891 1751 892 1755
rect 886 1750 892 1751
rect 918 1755 924 1756
rect 918 1751 919 1755
rect 923 1751 924 1755
rect 918 1750 924 1751
rect 950 1755 956 1756
rect 950 1751 951 1755
rect 955 1751 956 1755
rect 950 1750 956 1751
rect 982 1755 988 1756
rect 982 1751 983 1755
rect 987 1751 988 1755
rect 982 1750 988 1751
rect 1694 1753 1700 1754
rect 110 1748 116 1749
rect 1694 1749 1695 1753
rect 1699 1749 1700 1753
rect 1694 1748 1700 1749
rect 150 1738 156 1739
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 150 1734 151 1738
rect 155 1734 156 1738
rect 150 1733 156 1734
rect 182 1738 188 1739
rect 182 1734 183 1738
rect 187 1734 188 1738
rect 182 1733 188 1734
rect 214 1738 220 1739
rect 214 1734 215 1738
rect 219 1734 220 1738
rect 214 1733 220 1734
rect 246 1738 252 1739
rect 246 1734 247 1738
rect 251 1734 252 1738
rect 246 1733 252 1734
rect 278 1738 284 1739
rect 278 1734 279 1738
rect 283 1734 284 1738
rect 278 1733 284 1734
rect 310 1738 316 1739
rect 310 1734 311 1738
rect 315 1734 316 1738
rect 310 1733 316 1734
rect 342 1738 348 1739
rect 342 1734 343 1738
rect 347 1734 348 1738
rect 342 1733 348 1734
rect 374 1738 380 1739
rect 374 1734 375 1738
rect 379 1734 380 1738
rect 374 1733 380 1734
rect 406 1738 412 1739
rect 406 1734 407 1738
rect 411 1734 412 1738
rect 406 1733 412 1734
rect 438 1738 444 1739
rect 438 1734 439 1738
rect 443 1734 444 1738
rect 438 1733 444 1734
rect 470 1738 476 1739
rect 470 1734 471 1738
rect 475 1734 476 1738
rect 470 1733 476 1734
rect 502 1738 508 1739
rect 502 1734 503 1738
rect 507 1734 508 1738
rect 502 1733 508 1734
rect 534 1738 540 1739
rect 534 1734 535 1738
rect 539 1734 540 1738
rect 534 1733 540 1734
rect 566 1738 572 1739
rect 566 1734 567 1738
rect 571 1734 572 1738
rect 566 1733 572 1734
rect 598 1738 604 1739
rect 598 1734 599 1738
rect 603 1734 604 1738
rect 598 1733 604 1734
rect 630 1738 636 1739
rect 630 1734 631 1738
rect 635 1734 636 1738
rect 630 1733 636 1734
rect 662 1738 668 1739
rect 662 1734 663 1738
rect 667 1734 668 1738
rect 662 1733 668 1734
rect 694 1738 700 1739
rect 694 1734 695 1738
rect 699 1734 700 1738
rect 694 1733 700 1734
rect 726 1738 732 1739
rect 726 1734 727 1738
rect 731 1734 732 1738
rect 726 1733 732 1734
rect 758 1738 764 1739
rect 758 1734 759 1738
rect 763 1734 764 1738
rect 758 1733 764 1734
rect 790 1738 796 1739
rect 790 1734 791 1738
rect 795 1734 796 1738
rect 790 1733 796 1734
rect 822 1738 828 1739
rect 822 1734 823 1738
rect 827 1734 828 1738
rect 822 1733 828 1734
rect 854 1738 860 1739
rect 854 1734 855 1738
rect 859 1734 860 1738
rect 854 1733 860 1734
rect 886 1738 892 1739
rect 886 1734 887 1738
rect 891 1734 892 1738
rect 886 1733 892 1734
rect 918 1738 924 1739
rect 918 1734 919 1738
rect 923 1734 924 1738
rect 918 1733 924 1734
rect 950 1738 956 1739
rect 950 1734 951 1738
rect 955 1734 956 1738
rect 950 1733 956 1734
rect 982 1738 988 1739
rect 982 1734 983 1738
rect 987 1734 988 1738
rect 982 1733 988 1734
rect 1694 1736 1700 1737
rect 110 1731 116 1732
rect 1694 1732 1695 1736
rect 1699 1732 1700 1736
rect 1694 1731 1700 1732
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 1694 1704 1700 1705
rect 110 1699 116 1700
rect 190 1702 196 1703
rect 190 1698 191 1702
rect 195 1698 196 1702
rect 190 1697 196 1698
rect 246 1702 252 1703
rect 246 1698 247 1702
rect 251 1698 252 1702
rect 246 1697 252 1698
rect 318 1702 324 1703
rect 318 1698 319 1702
rect 323 1698 324 1702
rect 318 1697 324 1698
rect 414 1702 420 1703
rect 414 1698 415 1702
rect 419 1698 420 1702
rect 414 1697 420 1698
rect 526 1702 532 1703
rect 526 1698 527 1702
rect 531 1698 532 1702
rect 526 1697 532 1698
rect 654 1702 660 1703
rect 654 1698 655 1702
rect 659 1698 660 1702
rect 654 1697 660 1698
rect 790 1702 796 1703
rect 790 1698 791 1702
rect 795 1698 796 1702
rect 790 1697 796 1698
rect 918 1702 924 1703
rect 918 1698 919 1702
rect 923 1698 924 1702
rect 918 1697 924 1698
rect 1046 1702 1052 1703
rect 1046 1698 1047 1702
rect 1051 1698 1052 1702
rect 1046 1697 1052 1698
rect 1158 1702 1164 1703
rect 1158 1698 1159 1702
rect 1163 1698 1164 1702
rect 1158 1697 1164 1698
rect 1254 1702 1260 1703
rect 1254 1698 1255 1702
rect 1259 1698 1260 1702
rect 1254 1697 1260 1698
rect 1334 1702 1340 1703
rect 1334 1698 1335 1702
rect 1339 1698 1340 1702
rect 1334 1697 1340 1698
rect 1406 1702 1412 1703
rect 1406 1698 1407 1702
rect 1411 1698 1412 1702
rect 1406 1697 1412 1698
rect 1462 1702 1468 1703
rect 1462 1698 1463 1702
rect 1467 1698 1468 1702
rect 1462 1697 1468 1698
rect 1518 1702 1524 1703
rect 1518 1698 1519 1702
rect 1523 1698 1524 1702
rect 1518 1697 1524 1698
rect 1566 1702 1572 1703
rect 1566 1698 1567 1702
rect 1571 1698 1572 1702
rect 1566 1697 1572 1698
rect 1622 1702 1628 1703
rect 1622 1698 1623 1702
rect 1627 1698 1628 1702
rect 1622 1697 1628 1698
rect 1654 1702 1660 1703
rect 1654 1698 1655 1702
rect 1659 1698 1660 1702
rect 1694 1700 1695 1704
rect 1699 1700 1700 1704
rect 1694 1699 1700 1700
rect 1654 1697 1660 1698
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 1694 1687 1700 1688
rect 110 1682 116 1683
rect 190 1685 196 1686
rect 190 1681 191 1685
rect 195 1681 196 1685
rect 190 1680 196 1681
rect 246 1685 252 1686
rect 246 1681 247 1685
rect 251 1681 252 1685
rect 246 1680 252 1681
rect 318 1685 324 1686
rect 318 1681 319 1685
rect 323 1681 324 1685
rect 318 1680 324 1681
rect 414 1685 420 1686
rect 414 1681 415 1685
rect 419 1681 420 1685
rect 414 1680 420 1681
rect 526 1685 532 1686
rect 526 1681 527 1685
rect 531 1681 532 1685
rect 526 1680 532 1681
rect 654 1685 660 1686
rect 654 1681 655 1685
rect 659 1681 660 1685
rect 654 1680 660 1681
rect 790 1685 796 1686
rect 790 1681 791 1685
rect 795 1681 796 1685
rect 790 1680 796 1681
rect 918 1685 924 1686
rect 918 1681 919 1685
rect 923 1681 924 1685
rect 918 1680 924 1681
rect 1046 1685 1052 1686
rect 1046 1681 1047 1685
rect 1051 1681 1052 1685
rect 1046 1680 1052 1681
rect 1158 1685 1164 1686
rect 1158 1681 1159 1685
rect 1163 1681 1164 1685
rect 1158 1680 1164 1681
rect 1254 1685 1260 1686
rect 1254 1681 1255 1685
rect 1259 1681 1260 1685
rect 1254 1680 1260 1681
rect 1334 1685 1340 1686
rect 1334 1681 1335 1685
rect 1339 1681 1340 1685
rect 1334 1680 1340 1681
rect 1406 1685 1412 1686
rect 1406 1681 1407 1685
rect 1411 1681 1412 1685
rect 1406 1680 1412 1681
rect 1462 1685 1468 1686
rect 1462 1681 1463 1685
rect 1467 1681 1468 1685
rect 1462 1680 1468 1681
rect 1518 1685 1524 1686
rect 1518 1681 1519 1685
rect 1523 1681 1524 1685
rect 1518 1680 1524 1681
rect 1566 1685 1572 1686
rect 1566 1681 1567 1685
rect 1571 1681 1572 1685
rect 1566 1680 1572 1681
rect 1622 1685 1628 1686
rect 1622 1681 1623 1685
rect 1627 1681 1628 1685
rect 1622 1680 1628 1681
rect 1654 1685 1660 1686
rect 1654 1681 1655 1685
rect 1659 1681 1660 1685
rect 1694 1683 1695 1687
rect 1699 1683 1700 1687
rect 1694 1682 1700 1683
rect 1654 1680 1660 1681
rect 134 1663 140 1664
rect 110 1661 116 1662
rect 110 1657 111 1661
rect 115 1657 116 1661
rect 134 1659 135 1663
rect 139 1659 140 1663
rect 134 1658 140 1659
rect 174 1663 180 1664
rect 174 1659 175 1663
rect 179 1659 180 1663
rect 174 1658 180 1659
rect 262 1663 268 1664
rect 262 1659 263 1663
rect 267 1659 268 1663
rect 262 1658 268 1659
rect 390 1663 396 1664
rect 390 1659 391 1663
rect 395 1659 396 1663
rect 390 1658 396 1659
rect 542 1663 548 1664
rect 542 1659 543 1663
rect 547 1659 548 1663
rect 542 1658 548 1659
rect 710 1663 716 1664
rect 710 1659 711 1663
rect 715 1659 716 1663
rect 710 1658 716 1659
rect 878 1663 884 1664
rect 878 1659 879 1663
rect 883 1659 884 1663
rect 878 1658 884 1659
rect 1038 1663 1044 1664
rect 1038 1659 1039 1663
rect 1043 1659 1044 1663
rect 1038 1658 1044 1659
rect 1182 1663 1188 1664
rect 1182 1659 1183 1663
rect 1187 1659 1188 1663
rect 1182 1658 1188 1659
rect 1318 1663 1324 1664
rect 1318 1659 1319 1663
rect 1323 1659 1324 1663
rect 1318 1658 1324 1659
rect 1438 1663 1444 1664
rect 1438 1659 1439 1663
rect 1443 1659 1444 1663
rect 1438 1658 1444 1659
rect 1558 1663 1564 1664
rect 1558 1659 1559 1663
rect 1563 1659 1564 1663
rect 1558 1658 1564 1659
rect 1654 1663 1660 1664
rect 1654 1659 1655 1663
rect 1659 1659 1660 1663
rect 1654 1658 1660 1659
rect 1694 1661 1700 1662
rect 110 1656 116 1657
rect 1694 1657 1695 1661
rect 1699 1657 1700 1661
rect 1694 1656 1700 1657
rect 134 1646 140 1647
rect 110 1644 116 1645
rect 110 1640 111 1644
rect 115 1640 116 1644
rect 134 1642 135 1646
rect 139 1642 140 1646
rect 134 1641 140 1642
rect 174 1646 180 1647
rect 174 1642 175 1646
rect 179 1642 180 1646
rect 174 1641 180 1642
rect 262 1646 268 1647
rect 262 1642 263 1646
rect 267 1642 268 1646
rect 262 1641 268 1642
rect 390 1646 396 1647
rect 390 1642 391 1646
rect 395 1642 396 1646
rect 390 1641 396 1642
rect 542 1646 548 1647
rect 542 1642 543 1646
rect 547 1642 548 1646
rect 542 1641 548 1642
rect 710 1646 716 1647
rect 710 1642 711 1646
rect 715 1642 716 1646
rect 710 1641 716 1642
rect 878 1646 884 1647
rect 878 1642 879 1646
rect 883 1642 884 1646
rect 878 1641 884 1642
rect 1038 1646 1044 1647
rect 1038 1642 1039 1646
rect 1043 1642 1044 1646
rect 1038 1641 1044 1642
rect 1182 1646 1188 1647
rect 1182 1642 1183 1646
rect 1187 1642 1188 1646
rect 1182 1641 1188 1642
rect 1318 1646 1324 1647
rect 1318 1642 1319 1646
rect 1323 1642 1324 1646
rect 1318 1641 1324 1642
rect 1438 1646 1444 1647
rect 1438 1642 1439 1646
rect 1443 1642 1444 1646
rect 1438 1641 1444 1642
rect 1558 1646 1564 1647
rect 1558 1642 1559 1646
rect 1563 1642 1564 1646
rect 1558 1641 1564 1642
rect 1654 1646 1660 1647
rect 1654 1642 1655 1646
rect 1659 1642 1660 1646
rect 1654 1641 1660 1642
rect 1694 1644 1700 1645
rect 110 1639 116 1640
rect 1694 1640 1695 1644
rect 1699 1640 1700 1644
rect 1694 1639 1700 1640
rect 110 1608 116 1609
rect 110 1604 111 1608
rect 115 1604 116 1608
rect 1694 1608 1700 1609
rect 110 1603 116 1604
rect 134 1606 140 1607
rect 134 1602 135 1606
rect 139 1602 140 1606
rect 134 1601 140 1602
rect 166 1606 172 1607
rect 166 1602 167 1606
rect 171 1602 172 1606
rect 166 1601 172 1602
rect 198 1606 204 1607
rect 198 1602 199 1606
rect 203 1602 204 1606
rect 198 1601 204 1602
rect 246 1606 252 1607
rect 246 1602 247 1606
rect 251 1602 252 1606
rect 246 1601 252 1602
rect 326 1606 332 1607
rect 326 1602 327 1606
rect 331 1602 332 1606
rect 326 1601 332 1602
rect 438 1606 444 1607
rect 438 1602 439 1606
rect 443 1602 444 1606
rect 438 1601 444 1602
rect 566 1606 572 1607
rect 566 1602 567 1606
rect 571 1602 572 1606
rect 566 1601 572 1602
rect 710 1606 716 1607
rect 710 1602 711 1606
rect 715 1602 716 1606
rect 710 1601 716 1602
rect 854 1606 860 1607
rect 854 1602 855 1606
rect 859 1602 860 1606
rect 854 1601 860 1602
rect 998 1606 1004 1607
rect 998 1602 999 1606
rect 1003 1602 1004 1606
rect 998 1601 1004 1602
rect 1126 1606 1132 1607
rect 1126 1602 1127 1606
rect 1131 1602 1132 1606
rect 1126 1601 1132 1602
rect 1246 1606 1252 1607
rect 1246 1602 1247 1606
rect 1251 1602 1252 1606
rect 1246 1601 1252 1602
rect 1358 1606 1364 1607
rect 1358 1602 1359 1606
rect 1363 1602 1364 1606
rect 1358 1601 1364 1602
rect 1462 1606 1468 1607
rect 1462 1602 1463 1606
rect 1467 1602 1468 1606
rect 1462 1601 1468 1602
rect 1566 1606 1572 1607
rect 1566 1602 1567 1606
rect 1571 1602 1572 1606
rect 1566 1601 1572 1602
rect 1654 1606 1660 1607
rect 1654 1602 1655 1606
rect 1659 1602 1660 1606
rect 1694 1604 1695 1608
rect 1699 1604 1700 1608
rect 1694 1603 1700 1604
rect 1654 1601 1660 1602
rect 110 1591 116 1592
rect 110 1587 111 1591
rect 115 1587 116 1591
rect 1694 1591 1700 1592
rect 110 1586 116 1587
rect 134 1589 140 1590
rect 134 1585 135 1589
rect 139 1585 140 1589
rect 134 1584 140 1585
rect 166 1589 172 1590
rect 166 1585 167 1589
rect 171 1585 172 1589
rect 166 1584 172 1585
rect 198 1589 204 1590
rect 198 1585 199 1589
rect 203 1585 204 1589
rect 198 1584 204 1585
rect 246 1589 252 1590
rect 246 1585 247 1589
rect 251 1585 252 1589
rect 246 1584 252 1585
rect 326 1589 332 1590
rect 326 1585 327 1589
rect 331 1585 332 1589
rect 326 1584 332 1585
rect 438 1589 444 1590
rect 438 1585 439 1589
rect 443 1585 444 1589
rect 438 1584 444 1585
rect 566 1589 572 1590
rect 566 1585 567 1589
rect 571 1585 572 1589
rect 566 1584 572 1585
rect 710 1589 716 1590
rect 710 1585 711 1589
rect 715 1585 716 1589
rect 710 1584 716 1585
rect 854 1589 860 1590
rect 854 1585 855 1589
rect 859 1585 860 1589
rect 854 1584 860 1585
rect 998 1589 1004 1590
rect 998 1585 999 1589
rect 1003 1585 1004 1589
rect 998 1584 1004 1585
rect 1126 1589 1132 1590
rect 1126 1585 1127 1589
rect 1131 1585 1132 1589
rect 1126 1584 1132 1585
rect 1246 1589 1252 1590
rect 1246 1585 1247 1589
rect 1251 1585 1252 1589
rect 1246 1584 1252 1585
rect 1358 1589 1364 1590
rect 1358 1585 1359 1589
rect 1363 1585 1364 1589
rect 1358 1584 1364 1585
rect 1462 1589 1468 1590
rect 1462 1585 1463 1589
rect 1467 1585 1468 1589
rect 1462 1584 1468 1585
rect 1566 1589 1572 1590
rect 1566 1585 1567 1589
rect 1571 1585 1572 1589
rect 1566 1584 1572 1585
rect 1654 1589 1660 1590
rect 1654 1585 1655 1589
rect 1659 1585 1660 1589
rect 1694 1587 1695 1591
rect 1699 1587 1700 1591
rect 1694 1586 1700 1587
rect 1654 1584 1660 1585
rect 134 1575 140 1576
rect 110 1573 116 1574
rect 110 1569 111 1573
rect 115 1569 116 1573
rect 134 1571 135 1575
rect 139 1571 140 1575
rect 134 1570 140 1571
rect 166 1575 172 1576
rect 166 1571 167 1575
rect 171 1571 172 1575
rect 166 1570 172 1571
rect 230 1575 236 1576
rect 230 1571 231 1575
rect 235 1571 236 1575
rect 230 1570 236 1571
rect 286 1575 292 1576
rect 286 1571 287 1575
rect 291 1571 292 1575
rect 286 1570 292 1571
rect 342 1575 348 1576
rect 342 1571 343 1575
rect 347 1571 348 1575
rect 342 1570 348 1571
rect 398 1575 404 1576
rect 398 1571 399 1575
rect 403 1571 404 1575
rect 398 1570 404 1571
rect 454 1575 460 1576
rect 454 1571 455 1575
rect 459 1571 460 1575
rect 454 1570 460 1571
rect 510 1575 516 1576
rect 510 1571 511 1575
rect 515 1571 516 1575
rect 510 1570 516 1571
rect 574 1575 580 1576
rect 574 1571 575 1575
rect 579 1571 580 1575
rect 574 1570 580 1571
rect 654 1575 660 1576
rect 654 1571 655 1575
rect 659 1571 660 1575
rect 654 1570 660 1571
rect 750 1575 756 1576
rect 750 1571 751 1575
rect 755 1571 756 1575
rect 750 1570 756 1571
rect 854 1575 860 1576
rect 854 1571 855 1575
rect 859 1571 860 1575
rect 854 1570 860 1571
rect 958 1575 964 1576
rect 958 1571 959 1575
rect 963 1571 964 1575
rect 958 1570 964 1571
rect 1062 1575 1068 1576
rect 1062 1571 1063 1575
rect 1067 1571 1068 1575
rect 1062 1570 1068 1571
rect 1158 1575 1164 1576
rect 1158 1571 1159 1575
rect 1163 1571 1164 1575
rect 1158 1570 1164 1571
rect 1246 1575 1252 1576
rect 1246 1571 1247 1575
rect 1251 1571 1252 1575
rect 1246 1570 1252 1571
rect 1326 1575 1332 1576
rect 1326 1571 1327 1575
rect 1331 1571 1332 1575
rect 1326 1570 1332 1571
rect 1398 1575 1404 1576
rect 1398 1571 1399 1575
rect 1403 1571 1404 1575
rect 1398 1570 1404 1571
rect 1470 1575 1476 1576
rect 1470 1571 1471 1575
rect 1475 1571 1476 1575
rect 1470 1570 1476 1571
rect 1534 1575 1540 1576
rect 1534 1571 1535 1575
rect 1539 1571 1540 1575
rect 1534 1570 1540 1571
rect 1606 1575 1612 1576
rect 1606 1571 1607 1575
rect 1611 1571 1612 1575
rect 1606 1570 1612 1571
rect 1654 1575 1660 1576
rect 1654 1571 1655 1575
rect 1659 1571 1660 1575
rect 1654 1570 1660 1571
rect 1694 1573 1700 1574
rect 110 1568 116 1569
rect 1694 1569 1695 1573
rect 1699 1569 1700 1573
rect 1694 1568 1700 1569
rect 134 1558 140 1559
rect 110 1556 116 1557
rect 110 1552 111 1556
rect 115 1552 116 1556
rect 134 1554 135 1558
rect 139 1554 140 1558
rect 134 1553 140 1554
rect 166 1558 172 1559
rect 166 1554 167 1558
rect 171 1554 172 1558
rect 166 1553 172 1554
rect 230 1558 236 1559
rect 230 1554 231 1558
rect 235 1554 236 1558
rect 230 1553 236 1554
rect 286 1558 292 1559
rect 286 1554 287 1558
rect 291 1554 292 1558
rect 286 1553 292 1554
rect 342 1558 348 1559
rect 342 1554 343 1558
rect 347 1554 348 1558
rect 342 1553 348 1554
rect 398 1558 404 1559
rect 398 1554 399 1558
rect 403 1554 404 1558
rect 398 1553 404 1554
rect 454 1558 460 1559
rect 454 1554 455 1558
rect 459 1554 460 1558
rect 454 1553 460 1554
rect 510 1558 516 1559
rect 510 1554 511 1558
rect 515 1554 516 1558
rect 510 1553 516 1554
rect 574 1558 580 1559
rect 574 1554 575 1558
rect 579 1554 580 1558
rect 574 1553 580 1554
rect 654 1558 660 1559
rect 654 1554 655 1558
rect 659 1554 660 1558
rect 654 1553 660 1554
rect 750 1558 756 1559
rect 750 1554 751 1558
rect 755 1554 756 1558
rect 750 1553 756 1554
rect 854 1558 860 1559
rect 854 1554 855 1558
rect 859 1554 860 1558
rect 854 1553 860 1554
rect 958 1558 964 1559
rect 958 1554 959 1558
rect 963 1554 964 1558
rect 958 1553 964 1554
rect 1062 1558 1068 1559
rect 1062 1554 1063 1558
rect 1067 1554 1068 1558
rect 1062 1553 1068 1554
rect 1158 1558 1164 1559
rect 1158 1554 1159 1558
rect 1163 1554 1164 1558
rect 1158 1553 1164 1554
rect 1246 1558 1252 1559
rect 1246 1554 1247 1558
rect 1251 1554 1252 1558
rect 1246 1553 1252 1554
rect 1326 1558 1332 1559
rect 1326 1554 1327 1558
rect 1331 1554 1332 1558
rect 1326 1553 1332 1554
rect 1398 1558 1404 1559
rect 1398 1554 1399 1558
rect 1403 1554 1404 1558
rect 1398 1553 1404 1554
rect 1470 1558 1476 1559
rect 1470 1554 1471 1558
rect 1475 1554 1476 1558
rect 1470 1553 1476 1554
rect 1534 1558 1540 1559
rect 1534 1554 1535 1558
rect 1539 1554 1540 1558
rect 1534 1553 1540 1554
rect 1606 1558 1612 1559
rect 1606 1554 1607 1558
rect 1611 1554 1612 1558
rect 1606 1553 1612 1554
rect 1654 1558 1660 1559
rect 1654 1554 1655 1558
rect 1659 1554 1660 1558
rect 1654 1553 1660 1554
rect 1694 1556 1700 1557
rect 110 1551 116 1552
rect 1694 1552 1695 1556
rect 1699 1552 1700 1556
rect 1694 1551 1700 1552
rect 110 1528 116 1529
rect 110 1524 111 1528
rect 115 1524 116 1528
rect 1694 1528 1700 1529
rect 110 1523 116 1524
rect 134 1526 140 1527
rect 134 1522 135 1526
rect 139 1522 140 1526
rect 134 1521 140 1522
rect 174 1526 180 1527
rect 174 1522 175 1526
rect 179 1522 180 1526
rect 174 1521 180 1522
rect 222 1526 228 1527
rect 222 1522 223 1526
rect 227 1522 228 1526
rect 222 1521 228 1522
rect 278 1526 284 1527
rect 278 1522 279 1526
rect 283 1522 284 1526
rect 278 1521 284 1522
rect 334 1526 340 1527
rect 334 1522 335 1526
rect 339 1522 340 1526
rect 334 1521 340 1522
rect 398 1526 404 1527
rect 398 1522 399 1526
rect 403 1522 404 1526
rect 398 1521 404 1522
rect 462 1526 468 1527
rect 462 1522 463 1526
rect 467 1522 468 1526
rect 462 1521 468 1522
rect 534 1526 540 1527
rect 534 1522 535 1526
rect 539 1522 540 1526
rect 534 1521 540 1522
rect 606 1526 612 1527
rect 606 1522 607 1526
rect 611 1522 612 1526
rect 606 1521 612 1522
rect 686 1526 692 1527
rect 686 1522 687 1526
rect 691 1522 692 1526
rect 686 1521 692 1522
rect 774 1526 780 1527
rect 774 1522 775 1526
rect 779 1522 780 1526
rect 774 1521 780 1522
rect 870 1526 876 1527
rect 870 1522 871 1526
rect 875 1522 876 1526
rect 870 1521 876 1522
rect 974 1526 980 1527
rect 974 1522 975 1526
rect 979 1522 980 1526
rect 974 1521 980 1522
rect 1078 1526 1084 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1174 1526 1180 1527
rect 1174 1522 1175 1526
rect 1179 1522 1180 1526
rect 1174 1521 1180 1522
rect 1270 1526 1276 1527
rect 1270 1522 1271 1526
rect 1275 1522 1276 1526
rect 1270 1521 1276 1522
rect 1358 1526 1364 1527
rect 1358 1522 1359 1526
rect 1363 1522 1364 1526
rect 1358 1521 1364 1522
rect 1438 1526 1444 1527
rect 1438 1522 1439 1526
rect 1443 1522 1444 1526
rect 1438 1521 1444 1522
rect 1518 1526 1524 1527
rect 1518 1522 1519 1526
rect 1523 1522 1524 1526
rect 1518 1521 1524 1522
rect 1598 1526 1604 1527
rect 1598 1522 1599 1526
rect 1603 1522 1604 1526
rect 1598 1521 1604 1522
rect 1654 1526 1660 1527
rect 1654 1522 1655 1526
rect 1659 1522 1660 1526
rect 1694 1524 1695 1528
rect 1699 1524 1700 1528
rect 1694 1523 1700 1524
rect 1654 1521 1660 1522
rect 110 1511 116 1512
rect 110 1507 111 1511
rect 115 1507 116 1511
rect 1694 1511 1700 1512
rect 110 1506 116 1507
rect 134 1509 140 1510
rect 134 1505 135 1509
rect 139 1505 140 1509
rect 134 1504 140 1505
rect 174 1509 180 1510
rect 174 1505 175 1509
rect 179 1505 180 1509
rect 174 1504 180 1505
rect 222 1509 228 1510
rect 222 1505 223 1509
rect 227 1505 228 1509
rect 222 1504 228 1505
rect 278 1509 284 1510
rect 278 1505 279 1509
rect 283 1505 284 1509
rect 278 1504 284 1505
rect 334 1509 340 1510
rect 334 1505 335 1509
rect 339 1505 340 1509
rect 334 1504 340 1505
rect 398 1509 404 1510
rect 398 1505 399 1509
rect 403 1505 404 1509
rect 398 1504 404 1505
rect 462 1509 468 1510
rect 462 1505 463 1509
rect 467 1505 468 1509
rect 462 1504 468 1505
rect 534 1509 540 1510
rect 534 1505 535 1509
rect 539 1505 540 1509
rect 534 1504 540 1505
rect 606 1509 612 1510
rect 606 1505 607 1509
rect 611 1505 612 1509
rect 606 1504 612 1505
rect 686 1509 692 1510
rect 686 1505 687 1509
rect 691 1505 692 1509
rect 686 1504 692 1505
rect 774 1509 780 1510
rect 774 1505 775 1509
rect 779 1505 780 1509
rect 774 1504 780 1505
rect 870 1509 876 1510
rect 870 1505 871 1509
rect 875 1505 876 1509
rect 870 1504 876 1505
rect 974 1509 980 1510
rect 974 1505 975 1509
rect 979 1505 980 1509
rect 974 1504 980 1505
rect 1078 1509 1084 1510
rect 1078 1505 1079 1509
rect 1083 1505 1084 1509
rect 1078 1504 1084 1505
rect 1174 1509 1180 1510
rect 1174 1505 1175 1509
rect 1179 1505 1180 1509
rect 1174 1504 1180 1505
rect 1270 1509 1276 1510
rect 1270 1505 1271 1509
rect 1275 1505 1276 1509
rect 1270 1504 1276 1505
rect 1358 1509 1364 1510
rect 1358 1505 1359 1509
rect 1363 1505 1364 1509
rect 1358 1504 1364 1505
rect 1438 1509 1444 1510
rect 1438 1505 1439 1509
rect 1443 1505 1444 1509
rect 1438 1504 1444 1505
rect 1518 1509 1524 1510
rect 1518 1505 1519 1509
rect 1523 1505 1524 1509
rect 1518 1504 1524 1505
rect 1598 1509 1604 1510
rect 1598 1505 1599 1509
rect 1603 1505 1604 1509
rect 1598 1504 1604 1505
rect 1654 1509 1660 1510
rect 1654 1505 1655 1509
rect 1659 1505 1660 1509
rect 1694 1507 1695 1511
rect 1699 1507 1700 1511
rect 1694 1506 1700 1507
rect 1654 1504 1660 1505
rect 806 1476 812 1477
rect 174 1475 180 1476
rect 110 1473 116 1474
rect 110 1469 111 1473
rect 115 1469 116 1473
rect 174 1471 175 1475
rect 179 1471 180 1475
rect 174 1470 180 1471
rect 206 1475 212 1476
rect 206 1471 207 1475
rect 211 1471 212 1475
rect 206 1470 212 1471
rect 238 1475 244 1476
rect 238 1471 239 1475
rect 243 1471 244 1475
rect 238 1470 244 1471
rect 270 1475 276 1476
rect 270 1471 271 1475
rect 275 1471 276 1475
rect 270 1470 276 1471
rect 302 1475 308 1476
rect 302 1471 303 1475
rect 307 1471 308 1475
rect 302 1470 308 1471
rect 334 1475 340 1476
rect 334 1471 335 1475
rect 339 1471 340 1475
rect 334 1470 340 1471
rect 366 1475 372 1476
rect 366 1471 367 1475
rect 371 1471 372 1475
rect 366 1470 372 1471
rect 398 1475 404 1476
rect 398 1471 399 1475
rect 403 1471 404 1475
rect 398 1470 404 1471
rect 430 1475 436 1476
rect 430 1471 431 1475
rect 435 1471 436 1475
rect 430 1470 436 1471
rect 462 1475 468 1476
rect 462 1471 463 1475
rect 467 1471 468 1475
rect 462 1470 468 1471
rect 494 1475 500 1476
rect 494 1471 495 1475
rect 499 1471 500 1475
rect 494 1470 500 1471
rect 526 1475 532 1476
rect 526 1471 527 1475
rect 531 1471 532 1475
rect 526 1470 532 1471
rect 558 1475 564 1476
rect 558 1471 559 1475
rect 563 1471 564 1475
rect 558 1470 564 1471
rect 590 1475 596 1476
rect 590 1471 591 1475
rect 595 1471 596 1475
rect 590 1470 596 1471
rect 622 1475 628 1476
rect 622 1471 623 1475
rect 627 1471 628 1475
rect 622 1470 628 1471
rect 662 1475 668 1476
rect 662 1471 663 1475
rect 667 1471 668 1475
rect 662 1470 668 1471
rect 702 1475 708 1476
rect 702 1471 703 1475
rect 707 1471 708 1475
rect 702 1470 708 1471
rect 742 1475 748 1476
rect 742 1471 743 1475
rect 747 1471 748 1475
rect 742 1470 748 1471
rect 774 1475 780 1476
rect 774 1471 775 1475
rect 779 1471 780 1475
rect 806 1472 807 1476
rect 811 1472 812 1476
rect 806 1471 812 1472
rect 894 1476 900 1477
rect 894 1472 895 1476
rect 899 1472 900 1476
rect 894 1471 900 1472
rect 934 1476 940 1477
rect 934 1472 935 1476
rect 939 1472 940 1476
rect 934 1471 940 1472
rect 1022 1476 1028 1477
rect 1110 1476 1116 1477
rect 1022 1472 1023 1476
rect 1027 1472 1028 1476
rect 1022 1471 1028 1472
rect 1078 1475 1084 1476
rect 1078 1471 1079 1475
rect 1083 1471 1084 1475
rect 1110 1472 1111 1476
rect 1115 1472 1116 1476
rect 1110 1471 1116 1472
rect 1166 1475 1172 1476
rect 1166 1471 1167 1475
rect 1171 1471 1172 1475
rect 774 1470 780 1471
rect 1078 1470 1084 1471
rect 1166 1470 1172 1471
rect 1198 1475 1204 1476
rect 1198 1471 1199 1475
rect 1203 1471 1204 1475
rect 1198 1470 1204 1471
rect 1238 1475 1244 1476
rect 1238 1471 1239 1475
rect 1243 1471 1244 1475
rect 1238 1470 1244 1471
rect 1278 1475 1284 1476
rect 1278 1471 1279 1475
rect 1283 1471 1284 1475
rect 1278 1470 1284 1471
rect 1318 1475 1324 1476
rect 1318 1471 1319 1475
rect 1323 1471 1324 1475
rect 1318 1470 1324 1471
rect 1358 1475 1364 1476
rect 1358 1471 1359 1475
rect 1363 1471 1364 1475
rect 1358 1470 1364 1471
rect 1398 1475 1404 1476
rect 1398 1471 1399 1475
rect 1403 1471 1404 1475
rect 1398 1470 1404 1471
rect 1438 1475 1444 1476
rect 1438 1471 1439 1475
rect 1443 1471 1444 1475
rect 1438 1470 1444 1471
rect 1478 1475 1484 1476
rect 1478 1471 1479 1475
rect 1483 1471 1484 1475
rect 1478 1470 1484 1471
rect 1518 1475 1524 1476
rect 1518 1471 1519 1475
rect 1523 1471 1524 1475
rect 1518 1470 1524 1471
rect 1558 1475 1564 1476
rect 1558 1471 1559 1475
rect 1563 1471 1564 1475
rect 1558 1470 1564 1471
rect 1590 1475 1596 1476
rect 1590 1471 1591 1475
rect 1595 1471 1596 1475
rect 1590 1470 1596 1471
rect 1622 1475 1628 1476
rect 1622 1471 1623 1475
rect 1627 1471 1628 1475
rect 1622 1470 1628 1471
rect 1654 1475 1660 1476
rect 1654 1471 1655 1475
rect 1659 1471 1660 1475
rect 1654 1470 1660 1471
rect 1694 1473 1700 1474
rect 110 1468 116 1469
rect 1694 1469 1695 1473
rect 1699 1469 1700 1473
rect 1694 1468 1700 1469
rect 174 1458 180 1459
rect 110 1456 116 1457
rect 110 1452 111 1456
rect 115 1452 116 1456
rect 174 1454 175 1458
rect 179 1454 180 1458
rect 174 1453 180 1454
rect 206 1458 212 1459
rect 206 1454 207 1458
rect 211 1454 212 1458
rect 206 1453 212 1454
rect 238 1458 244 1459
rect 238 1454 239 1458
rect 243 1454 244 1458
rect 238 1453 244 1454
rect 270 1458 276 1459
rect 270 1454 271 1458
rect 275 1454 276 1458
rect 270 1453 276 1454
rect 302 1458 308 1459
rect 302 1454 303 1458
rect 307 1454 308 1458
rect 302 1453 308 1454
rect 334 1458 340 1459
rect 334 1454 335 1458
rect 339 1454 340 1458
rect 334 1453 340 1454
rect 366 1458 372 1459
rect 366 1454 367 1458
rect 371 1454 372 1458
rect 366 1453 372 1454
rect 398 1458 404 1459
rect 398 1454 399 1458
rect 403 1454 404 1458
rect 398 1453 404 1454
rect 430 1458 436 1459
rect 430 1454 431 1458
rect 435 1454 436 1458
rect 430 1453 436 1454
rect 462 1458 468 1459
rect 462 1454 463 1458
rect 467 1454 468 1458
rect 462 1453 468 1454
rect 494 1458 500 1459
rect 494 1454 495 1458
rect 499 1454 500 1458
rect 494 1453 500 1454
rect 526 1458 532 1459
rect 526 1454 527 1458
rect 531 1454 532 1458
rect 526 1453 532 1454
rect 558 1458 564 1459
rect 558 1454 559 1458
rect 563 1454 564 1458
rect 558 1453 564 1454
rect 590 1458 596 1459
rect 590 1454 591 1458
rect 595 1454 596 1458
rect 590 1453 596 1454
rect 622 1458 628 1459
rect 622 1454 623 1458
rect 627 1454 628 1458
rect 622 1453 628 1454
rect 662 1458 668 1459
rect 662 1454 663 1458
rect 667 1454 668 1458
rect 662 1453 668 1454
rect 702 1458 708 1459
rect 702 1454 703 1458
rect 707 1454 708 1458
rect 702 1453 708 1454
rect 742 1458 748 1459
rect 1078 1458 1084 1459
rect 742 1454 743 1458
rect 747 1454 748 1458
rect 742 1453 748 1454
rect 774 1457 780 1458
rect 774 1453 775 1457
rect 779 1453 780 1457
rect 774 1452 780 1453
rect 806 1457 812 1458
rect 806 1453 807 1457
rect 811 1453 812 1457
rect 806 1452 812 1453
rect 934 1457 940 1458
rect 934 1453 935 1457
rect 939 1453 940 1457
rect 934 1452 940 1453
rect 1038 1455 1044 1456
rect 110 1451 116 1452
rect 1038 1451 1039 1455
rect 1043 1451 1044 1455
rect 1078 1454 1079 1458
rect 1083 1454 1084 1458
rect 1166 1458 1172 1459
rect 1078 1453 1084 1454
rect 1126 1455 1132 1456
rect 1038 1450 1044 1451
rect 1126 1451 1127 1455
rect 1131 1451 1132 1455
rect 1166 1454 1167 1458
rect 1171 1454 1172 1458
rect 1166 1453 1172 1454
rect 1198 1458 1204 1459
rect 1198 1454 1199 1458
rect 1203 1454 1204 1458
rect 1198 1453 1204 1454
rect 1238 1458 1244 1459
rect 1318 1458 1324 1459
rect 1238 1454 1239 1458
rect 1243 1454 1244 1458
rect 1238 1453 1244 1454
rect 1278 1457 1284 1458
rect 1278 1453 1279 1457
rect 1283 1453 1284 1457
rect 1318 1454 1319 1458
rect 1323 1454 1324 1458
rect 1318 1453 1324 1454
rect 1358 1458 1364 1459
rect 1358 1454 1359 1458
rect 1363 1454 1364 1458
rect 1358 1453 1364 1454
rect 1398 1458 1404 1459
rect 1398 1454 1399 1458
rect 1403 1454 1404 1458
rect 1398 1453 1404 1454
rect 1438 1458 1444 1459
rect 1438 1454 1439 1458
rect 1443 1454 1444 1458
rect 1438 1453 1444 1454
rect 1478 1458 1484 1459
rect 1478 1454 1479 1458
rect 1483 1454 1484 1458
rect 1478 1453 1484 1454
rect 1518 1458 1524 1459
rect 1518 1454 1519 1458
rect 1523 1454 1524 1458
rect 1518 1453 1524 1454
rect 1558 1458 1564 1459
rect 1558 1454 1559 1458
rect 1563 1454 1564 1458
rect 1558 1453 1564 1454
rect 1590 1458 1596 1459
rect 1590 1454 1591 1458
rect 1595 1454 1596 1458
rect 1590 1453 1596 1454
rect 1622 1458 1628 1459
rect 1622 1454 1623 1458
rect 1627 1454 1628 1458
rect 1622 1453 1628 1454
rect 1654 1458 1660 1459
rect 1654 1454 1655 1458
rect 1659 1454 1660 1458
rect 1654 1453 1660 1454
rect 1694 1456 1700 1457
rect 1278 1452 1284 1453
rect 1694 1452 1695 1456
rect 1699 1452 1700 1456
rect 1694 1451 1700 1452
rect 1126 1450 1132 1451
rect 894 1448 900 1449
rect 894 1444 895 1448
rect 899 1444 900 1448
rect 894 1443 900 1444
rect 766 1415 772 1416
rect 766 1411 767 1415
rect 771 1411 772 1415
rect 766 1410 772 1411
rect 838 1415 844 1416
rect 838 1411 839 1415
rect 843 1411 844 1415
rect 974 1415 980 1416
rect 974 1411 975 1415
rect 979 1411 980 1415
rect 838 1410 844 1411
rect 894 1410 900 1411
rect 974 1410 980 1411
rect 894 1406 895 1410
rect 899 1406 900 1410
rect 894 1405 900 1406
rect 1062 1400 1068 1401
rect 1062 1396 1063 1400
rect 1067 1396 1068 1400
rect 806 1395 812 1396
rect 1062 1395 1068 1396
rect 1150 1400 1156 1401
rect 1150 1396 1151 1400
rect 1155 1396 1156 1400
rect 1150 1395 1156 1396
rect 718 1393 724 1394
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 134 1390 140 1391
rect 134 1386 135 1390
rect 139 1386 140 1390
rect 134 1385 140 1386
rect 166 1390 172 1391
rect 166 1386 167 1390
rect 171 1386 172 1390
rect 166 1385 172 1386
rect 198 1390 204 1391
rect 198 1386 199 1390
rect 203 1386 204 1390
rect 198 1385 204 1386
rect 230 1390 236 1391
rect 230 1386 231 1390
rect 235 1386 236 1390
rect 230 1385 236 1386
rect 262 1390 268 1391
rect 262 1386 263 1390
rect 267 1386 268 1390
rect 262 1385 268 1386
rect 294 1390 300 1391
rect 294 1386 295 1390
rect 299 1386 300 1390
rect 294 1385 300 1386
rect 326 1390 332 1391
rect 326 1386 327 1390
rect 331 1386 332 1390
rect 326 1385 332 1386
rect 358 1390 364 1391
rect 358 1386 359 1390
rect 363 1386 364 1390
rect 358 1385 364 1386
rect 390 1390 396 1391
rect 390 1386 391 1390
rect 395 1386 396 1390
rect 390 1385 396 1386
rect 422 1390 428 1391
rect 422 1386 423 1390
rect 427 1386 428 1390
rect 422 1385 428 1386
rect 454 1390 460 1391
rect 454 1386 455 1390
rect 459 1386 460 1390
rect 454 1385 460 1386
rect 486 1390 492 1391
rect 486 1386 487 1390
rect 491 1386 492 1390
rect 486 1385 492 1386
rect 518 1390 524 1391
rect 518 1386 519 1390
rect 523 1386 524 1390
rect 518 1385 524 1386
rect 550 1390 556 1391
rect 550 1386 551 1390
rect 555 1386 556 1390
rect 550 1385 556 1386
rect 582 1390 588 1391
rect 582 1386 583 1390
rect 587 1386 588 1390
rect 582 1385 588 1386
rect 614 1390 620 1391
rect 614 1386 615 1390
rect 619 1386 620 1390
rect 614 1385 620 1386
rect 646 1390 652 1391
rect 646 1386 647 1390
rect 651 1386 652 1390
rect 646 1385 652 1386
rect 678 1390 684 1391
rect 678 1386 679 1390
rect 683 1386 684 1390
rect 718 1389 719 1393
rect 723 1389 724 1393
rect 806 1391 807 1395
rect 811 1391 812 1395
rect 1262 1393 1268 1394
rect 1110 1391 1116 1392
rect 806 1390 812 1391
rect 1022 1390 1028 1391
rect 718 1388 724 1389
rect 678 1385 684 1386
rect 1022 1386 1023 1390
rect 1027 1386 1028 1390
rect 1110 1387 1111 1391
rect 1115 1387 1116 1391
rect 1110 1386 1116 1387
rect 1198 1390 1204 1391
rect 1198 1386 1199 1390
rect 1203 1386 1204 1390
rect 1262 1389 1263 1393
rect 1267 1389 1268 1393
rect 1478 1393 1484 1394
rect 1262 1388 1268 1389
rect 1318 1391 1324 1392
rect 1318 1387 1319 1391
rect 1323 1387 1324 1391
rect 1318 1386 1324 1387
rect 1414 1390 1420 1391
rect 1414 1386 1415 1390
rect 1419 1386 1420 1390
rect 1478 1389 1479 1393
rect 1483 1389 1484 1393
rect 1694 1392 1700 1393
rect 1478 1388 1484 1389
rect 1534 1390 1540 1391
rect 1022 1385 1028 1386
rect 1198 1385 1204 1386
rect 1414 1385 1420 1386
rect 1534 1386 1535 1390
rect 1539 1386 1540 1390
rect 1534 1385 1540 1386
rect 1582 1390 1588 1391
rect 1582 1386 1583 1390
rect 1587 1386 1588 1390
rect 1582 1385 1588 1386
rect 1622 1390 1628 1391
rect 1622 1386 1623 1390
rect 1627 1386 1628 1390
rect 1622 1385 1628 1386
rect 1654 1390 1660 1391
rect 1654 1386 1655 1390
rect 1659 1386 1660 1390
rect 1694 1388 1695 1392
rect 1699 1388 1700 1392
rect 1694 1387 1700 1388
rect 1654 1385 1660 1386
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 1694 1375 1700 1376
rect 110 1370 116 1371
rect 134 1373 140 1374
rect 134 1369 135 1373
rect 139 1369 140 1373
rect 134 1368 140 1369
rect 166 1373 172 1374
rect 166 1369 167 1373
rect 171 1369 172 1373
rect 166 1368 172 1369
rect 198 1373 204 1374
rect 198 1369 199 1373
rect 203 1369 204 1373
rect 198 1368 204 1369
rect 230 1373 236 1374
rect 230 1369 231 1373
rect 235 1369 236 1373
rect 230 1368 236 1369
rect 262 1373 268 1374
rect 262 1369 263 1373
rect 267 1369 268 1373
rect 262 1368 268 1369
rect 294 1373 300 1374
rect 294 1369 295 1373
rect 299 1369 300 1373
rect 294 1368 300 1369
rect 326 1373 332 1374
rect 326 1369 327 1373
rect 331 1369 332 1373
rect 326 1368 332 1369
rect 358 1373 364 1374
rect 358 1369 359 1373
rect 363 1369 364 1373
rect 358 1368 364 1369
rect 390 1373 396 1374
rect 390 1369 391 1373
rect 395 1369 396 1373
rect 390 1368 396 1369
rect 422 1373 428 1374
rect 422 1369 423 1373
rect 427 1369 428 1373
rect 422 1368 428 1369
rect 454 1373 460 1374
rect 454 1369 455 1373
rect 459 1369 460 1373
rect 454 1368 460 1369
rect 486 1373 492 1374
rect 486 1369 487 1373
rect 491 1369 492 1373
rect 486 1368 492 1369
rect 518 1373 524 1374
rect 518 1369 519 1373
rect 523 1369 524 1373
rect 518 1368 524 1369
rect 550 1373 556 1374
rect 550 1369 551 1373
rect 555 1369 556 1373
rect 550 1368 556 1369
rect 582 1373 588 1374
rect 582 1369 583 1373
rect 587 1369 588 1373
rect 582 1368 588 1369
rect 614 1373 620 1374
rect 614 1369 615 1373
rect 619 1369 620 1373
rect 614 1368 620 1369
rect 646 1373 652 1374
rect 646 1369 647 1373
rect 651 1369 652 1373
rect 646 1368 652 1369
rect 678 1373 684 1374
rect 1022 1373 1028 1374
rect 1110 1373 1116 1374
rect 1198 1373 1204 1374
rect 1414 1373 1420 1374
rect 1534 1373 1540 1374
rect 678 1369 679 1373
rect 683 1369 684 1373
rect 806 1372 812 1373
rect 678 1368 684 1369
rect 766 1368 772 1369
rect 734 1366 740 1367
rect 734 1362 735 1366
rect 739 1362 740 1366
rect 766 1364 767 1368
rect 771 1364 772 1368
rect 806 1368 807 1372
rect 811 1368 812 1372
rect 886 1372 892 1373
rect 806 1367 812 1368
rect 838 1368 844 1369
rect 766 1363 772 1364
rect 838 1364 839 1368
rect 843 1364 844 1368
rect 886 1368 887 1372
rect 891 1368 892 1372
rect 1022 1369 1023 1373
rect 1027 1369 1028 1373
rect 886 1367 892 1368
rect 974 1368 980 1369
rect 1022 1368 1028 1369
rect 1062 1372 1068 1373
rect 1062 1368 1063 1372
rect 1067 1368 1068 1372
rect 1110 1369 1111 1373
rect 1115 1369 1116 1373
rect 1110 1368 1116 1369
rect 1150 1372 1156 1373
rect 1150 1368 1151 1372
rect 1155 1368 1156 1372
rect 1198 1369 1199 1373
rect 1203 1369 1204 1373
rect 1198 1368 1204 1369
rect 1246 1372 1252 1373
rect 1246 1368 1247 1372
rect 1251 1368 1252 1372
rect 838 1363 844 1364
rect 974 1364 975 1368
rect 979 1364 980 1368
rect 1062 1367 1068 1368
rect 1150 1367 1156 1368
rect 1246 1367 1252 1368
rect 1318 1372 1324 1373
rect 1318 1368 1319 1372
rect 1323 1368 1324 1372
rect 1414 1369 1415 1373
rect 1419 1369 1420 1373
rect 1414 1368 1420 1369
rect 1462 1372 1468 1373
rect 1462 1368 1463 1372
rect 1467 1368 1468 1372
rect 1534 1369 1535 1373
rect 1539 1369 1540 1373
rect 1534 1368 1540 1369
rect 1582 1373 1588 1374
rect 1582 1369 1583 1373
rect 1587 1369 1588 1373
rect 1582 1368 1588 1369
rect 1622 1373 1628 1374
rect 1622 1369 1623 1373
rect 1627 1369 1628 1373
rect 1622 1368 1628 1369
rect 1654 1373 1660 1374
rect 1654 1369 1655 1373
rect 1659 1369 1660 1373
rect 1694 1371 1695 1375
rect 1699 1371 1700 1375
rect 1694 1370 1700 1371
rect 1654 1368 1660 1369
rect 1318 1367 1324 1368
rect 1462 1367 1468 1368
rect 974 1363 980 1364
rect 734 1361 740 1362
rect 982 1324 988 1325
rect 742 1320 748 1321
rect 134 1319 140 1320
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1315 135 1319
rect 139 1315 140 1319
rect 134 1314 140 1315
rect 166 1319 172 1320
rect 166 1315 167 1319
rect 171 1315 172 1319
rect 166 1314 172 1315
rect 198 1319 204 1320
rect 198 1315 199 1319
rect 203 1315 204 1319
rect 198 1314 204 1315
rect 230 1319 236 1320
rect 230 1315 231 1319
rect 235 1315 236 1319
rect 230 1314 236 1315
rect 262 1319 268 1320
rect 262 1315 263 1319
rect 267 1315 268 1319
rect 262 1314 268 1315
rect 294 1319 300 1320
rect 294 1315 295 1319
rect 299 1315 300 1319
rect 294 1314 300 1315
rect 326 1319 332 1320
rect 326 1315 327 1319
rect 331 1315 332 1319
rect 326 1314 332 1315
rect 358 1319 364 1320
rect 358 1315 359 1319
rect 363 1315 364 1319
rect 358 1314 364 1315
rect 390 1319 396 1320
rect 390 1315 391 1319
rect 395 1315 396 1319
rect 390 1314 396 1315
rect 422 1319 428 1320
rect 422 1315 423 1319
rect 427 1315 428 1319
rect 422 1314 428 1315
rect 454 1319 460 1320
rect 454 1315 455 1319
rect 459 1315 460 1319
rect 454 1314 460 1315
rect 486 1319 492 1320
rect 486 1315 487 1319
rect 491 1315 492 1319
rect 486 1314 492 1315
rect 518 1319 524 1320
rect 518 1315 519 1319
rect 523 1315 524 1319
rect 518 1314 524 1315
rect 550 1319 556 1320
rect 550 1315 551 1319
rect 555 1315 556 1319
rect 550 1314 556 1315
rect 582 1319 588 1320
rect 582 1315 583 1319
rect 587 1315 588 1319
rect 582 1314 588 1315
rect 614 1319 620 1320
rect 614 1315 615 1319
rect 619 1315 620 1319
rect 614 1314 620 1315
rect 646 1319 652 1320
rect 646 1315 647 1319
rect 651 1315 652 1319
rect 646 1314 652 1315
rect 678 1319 684 1320
rect 678 1315 679 1319
rect 683 1315 684 1319
rect 678 1314 684 1315
rect 710 1319 716 1320
rect 710 1315 711 1319
rect 715 1315 716 1319
rect 742 1316 743 1320
rect 747 1316 748 1320
rect 742 1315 748 1316
rect 822 1320 828 1321
rect 822 1316 823 1320
rect 827 1316 828 1320
rect 822 1315 828 1316
rect 902 1320 908 1321
rect 902 1316 903 1320
rect 907 1316 908 1320
rect 982 1320 983 1324
rect 987 1320 988 1324
rect 982 1319 988 1320
rect 1022 1320 1028 1321
rect 902 1315 908 1316
rect 1022 1316 1023 1320
rect 1027 1316 1028 1320
rect 1022 1315 1028 1316
rect 1062 1320 1068 1321
rect 1062 1316 1063 1320
rect 1067 1316 1068 1320
rect 1062 1315 1068 1316
rect 1158 1320 1164 1321
rect 1158 1316 1159 1320
rect 1163 1316 1164 1320
rect 1158 1315 1164 1316
rect 1214 1320 1220 1321
rect 1214 1316 1215 1320
rect 1219 1316 1220 1320
rect 1214 1315 1220 1316
rect 1302 1320 1308 1321
rect 1454 1320 1460 1321
rect 1302 1316 1303 1320
rect 1307 1316 1308 1320
rect 1302 1315 1308 1316
rect 1390 1319 1396 1320
rect 1390 1315 1391 1319
rect 1395 1315 1396 1319
rect 710 1314 716 1315
rect 1390 1314 1396 1315
rect 1422 1319 1428 1320
rect 1422 1315 1423 1319
rect 1427 1315 1428 1319
rect 1454 1316 1455 1320
rect 1459 1316 1460 1320
rect 1454 1315 1460 1316
rect 1494 1319 1500 1320
rect 1494 1315 1495 1319
rect 1499 1315 1500 1319
rect 1422 1314 1428 1315
rect 1494 1314 1500 1315
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1558 1319 1564 1320
rect 1558 1315 1559 1319
rect 1563 1315 1564 1319
rect 1558 1314 1564 1315
rect 1590 1319 1596 1320
rect 1590 1315 1591 1319
rect 1595 1315 1596 1319
rect 1590 1314 1596 1315
rect 1622 1319 1628 1320
rect 1622 1315 1623 1319
rect 1627 1315 1628 1319
rect 1622 1314 1628 1315
rect 1654 1319 1660 1320
rect 1654 1315 1655 1319
rect 1659 1315 1660 1319
rect 1654 1314 1660 1315
rect 1694 1317 1700 1318
rect 110 1312 116 1313
rect 1694 1313 1695 1317
rect 1699 1313 1700 1317
rect 1694 1312 1700 1313
rect 134 1302 140 1303
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 134 1298 135 1302
rect 139 1298 140 1302
rect 134 1297 140 1298
rect 166 1302 172 1303
rect 166 1298 167 1302
rect 171 1298 172 1302
rect 166 1297 172 1298
rect 198 1302 204 1303
rect 198 1298 199 1302
rect 203 1298 204 1302
rect 198 1297 204 1298
rect 230 1302 236 1303
rect 230 1298 231 1302
rect 235 1298 236 1302
rect 230 1297 236 1298
rect 262 1302 268 1303
rect 262 1298 263 1302
rect 267 1298 268 1302
rect 262 1297 268 1298
rect 294 1302 300 1303
rect 294 1298 295 1302
rect 299 1298 300 1302
rect 294 1297 300 1298
rect 326 1302 332 1303
rect 326 1298 327 1302
rect 331 1298 332 1302
rect 326 1297 332 1298
rect 358 1302 364 1303
rect 358 1298 359 1302
rect 363 1298 364 1302
rect 358 1297 364 1298
rect 390 1302 396 1303
rect 390 1298 391 1302
rect 395 1298 396 1302
rect 390 1297 396 1298
rect 422 1302 428 1303
rect 422 1298 423 1302
rect 427 1298 428 1302
rect 422 1297 428 1298
rect 454 1302 460 1303
rect 454 1298 455 1302
rect 459 1298 460 1302
rect 454 1297 460 1298
rect 486 1302 492 1303
rect 486 1298 487 1302
rect 491 1298 492 1302
rect 486 1297 492 1298
rect 518 1302 524 1303
rect 518 1298 519 1302
rect 523 1298 524 1302
rect 518 1297 524 1298
rect 550 1302 556 1303
rect 550 1298 551 1302
rect 555 1298 556 1302
rect 550 1297 556 1298
rect 582 1302 588 1303
rect 582 1298 583 1302
rect 587 1298 588 1302
rect 582 1297 588 1298
rect 614 1302 620 1303
rect 614 1298 615 1302
rect 619 1298 620 1302
rect 614 1297 620 1298
rect 646 1302 652 1303
rect 646 1298 647 1302
rect 651 1298 652 1302
rect 646 1297 652 1298
rect 678 1302 684 1303
rect 678 1298 679 1302
rect 683 1298 684 1302
rect 678 1297 684 1298
rect 710 1302 716 1303
rect 1422 1302 1428 1303
rect 710 1298 711 1302
rect 715 1298 716 1302
rect 710 1297 716 1298
rect 1062 1301 1068 1302
rect 1062 1297 1063 1301
rect 1067 1297 1068 1301
rect 1214 1301 1220 1302
rect 1062 1296 1068 1297
rect 1174 1299 1180 1300
rect 110 1295 116 1296
rect 1174 1295 1175 1299
rect 1179 1295 1180 1299
rect 1214 1297 1215 1301
rect 1219 1297 1220 1301
rect 1214 1296 1220 1297
rect 1302 1301 1308 1302
rect 1302 1297 1303 1301
rect 1307 1297 1308 1301
rect 1302 1296 1308 1297
rect 1390 1301 1396 1302
rect 1390 1297 1391 1301
rect 1395 1297 1396 1301
rect 1422 1298 1423 1302
rect 1427 1298 1428 1302
rect 1422 1297 1428 1298
rect 1494 1302 1500 1303
rect 1494 1298 1495 1302
rect 1499 1298 1500 1302
rect 1494 1297 1500 1298
rect 1526 1302 1532 1303
rect 1526 1298 1527 1302
rect 1531 1298 1532 1302
rect 1526 1297 1532 1298
rect 1558 1302 1564 1303
rect 1558 1298 1559 1302
rect 1563 1298 1564 1302
rect 1558 1297 1564 1298
rect 1590 1302 1596 1303
rect 1590 1298 1591 1302
rect 1595 1298 1596 1302
rect 1590 1297 1596 1298
rect 1622 1302 1628 1303
rect 1622 1298 1623 1302
rect 1627 1298 1628 1302
rect 1622 1297 1628 1298
rect 1654 1302 1660 1303
rect 1654 1298 1655 1302
rect 1659 1298 1660 1302
rect 1654 1297 1660 1298
rect 1694 1300 1700 1301
rect 1390 1296 1396 1297
rect 1694 1296 1695 1300
rect 1699 1296 1700 1300
rect 1694 1295 1700 1296
rect 1174 1294 1180 1295
rect 1022 1292 1028 1293
rect 1022 1288 1023 1292
rect 1027 1288 1028 1292
rect 1022 1287 1028 1288
rect 1454 1292 1460 1293
rect 1454 1288 1455 1292
rect 1459 1288 1460 1292
rect 1454 1287 1460 1288
rect 750 1282 756 1283
rect 750 1278 751 1282
rect 755 1278 756 1282
rect 750 1277 756 1278
rect 830 1282 836 1283
rect 830 1278 831 1282
rect 835 1278 836 1282
rect 830 1277 836 1278
rect 910 1282 916 1283
rect 910 1278 911 1282
rect 915 1278 916 1282
rect 910 1277 916 1278
rect 982 1277 988 1278
rect 982 1273 983 1277
rect 987 1273 988 1277
rect 982 1272 988 1273
rect 774 1219 780 1220
rect 774 1215 775 1219
rect 779 1215 780 1219
rect 1086 1219 1092 1220
rect 1086 1215 1087 1219
rect 1091 1215 1092 1219
rect 774 1214 780 1215
rect 1014 1214 1020 1215
rect 1086 1214 1092 1215
rect 1014 1210 1015 1214
rect 1019 1210 1020 1214
rect 1014 1209 1020 1210
rect 958 1197 964 1198
rect 110 1196 116 1197
rect 110 1192 111 1196
rect 115 1192 116 1196
rect 810 1195 816 1196
rect 110 1191 116 1192
rect 134 1194 140 1195
rect 134 1190 135 1194
rect 139 1190 140 1194
rect 134 1189 140 1190
rect 166 1194 172 1195
rect 166 1190 167 1194
rect 171 1190 172 1194
rect 166 1189 172 1190
rect 198 1194 204 1195
rect 198 1190 199 1194
rect 203 1190 204 1194
rect 198 1189 204 1190
rect 230 1194 236 1195
rect 230 1190 231 1194
rect 235 1190 236 1194
rect 230 1189 236 1190
rect 262 1194 268 1195
rect 262 1190 263 1194
rect 267 1190 268 1194
rect 262 1189 268 1190
rect 294 1194 300 1195
rect 294 1190 295 1194
rect 299 1190 300 1194
rect 294 1189 300 1190
rect 326 1194 332 1195
rect 326 1190 327 1194
rect 331 1190 332 1194
rect 326 1189 332 1190
rect 358 1194 364 1195
rect 358 1190 359 1194
rect 363 1190 364 1194
rect 358 1189 364 1190
rect 390 1194 396 1195
rect 390 1190 391 1194
rect 395 1190 396 1194
rect 390 1189 396 1190
rect 422 1194 428 1195
rect 422 1190 423 1194
rect 427 1190 428 1194
rect 422 1189 428 1190
rect 454 1194 460 1195
rect 454 1190 455 1194
rect 459 1190 460 1194
rect 454 1189 460 1190
rect 486 1194 492 1195
rect 486 1190 487 1194
rect 491 1190 492 1194
rect 486 1189 492 1190
rect 518 1194 524 1195
rect 518 1190 519 1194
rect 523 1190 524 1194
rect 518 1189 524 1190
rect 550 1194 556 1195
rect 550 1190 551 1194
rect 555 1190 556 1194
rect 550 1189 556 1190
rect 582 1194 588 1195
rect 582 1190 583 1194
rect 587 1190 588 1194
rect 582 1189 588 1190
rect 614 1194 620 1195
rect 614 1190 615 1194
rect 619 1190 620 1194
rect 614 1189 620 1190
rect 646 1194 652 1195
rect 646 1190 647 1194
rect 651 1190 652 1194
rect 646 1189 652 1190
rect 678 1194 684 1195
rect 678 1190 679 1194
rect 683 1190 684 1194
rect 678 1189 684 1190
rect 710 1194 716 1195
rect 710 1190 711 1194
rect 715 1190 716 1194
rect 710 1189 716 1190
rect 742 1194 748 1195
rect 742 1190 743 1194
rect 747 1190 748 1194
rect 810 1191 811 1195
rect 815 1191 816 1195
rect 958 1193 959 1197
rect 963 1193 964 1197
rect 1214 1197 1220 1198
rect 958 1192 964 1193
rect 1126 1194 1132 1195
rect 810 1190 816 1191
rect 1126 1190 1127 1194
rect 1131 1190 1132 1194
rect 742 1189 748 1190
rect 1126 1189 1132 1190
rect 1158 1194 1164 1195
rect 1158 1190 1159 1194
rect 1163 1190 1164 1194
rect 1214 1193 1215 1197
rect 1219 1193 1220 1197
rect 1294 1197 1300 1198
rect 1214 1192 1220 1193
rect 1254 1194 1260 1195
rect 1158 1189 1164 1190
rect 1254 1190 1255 1194
rect 1259 1190 1260 1194
rect 1294 1193 1295 1197
rect 1299 1193 1300 1197
rect 1694 1196 1700 1197
rect 1294 1192 1300 1193
rect 1342 1194 1348 1195
rect 1254 1189 1260 1190
rect 1342 1190 1343 1194
rect 1347 1190 1348 1194
rect 1342 1189 1348 1190
rect 1374 1194 1380 1195
rect 1374 1190 1375 1194
rect 1379 1190 1380 1194
rect 1374 1189 1380 1190
rect 1406 1194 1412 1195
rect 1406 1190 1407 1194
rect 1411 1190 1412 1194
rect 1406 1189 1412 1190
rect 1438 1194 1444 1195
rect 1438 1190 1439 1194
rect 1443 1190 1444 1194
rect 1438 1189 1444 1190
rect 1478 1194 1484 1195
rect 1478 1190 1479 1194
rect 1483 1190 1484 1194
rect 1478 1189 1484 1190
rect 1518 1194 1524 1195
rect 1518 1190 1519 1194
rect 1523 1190 1524 1194
rect 1518 1189 1524 1190
rect 1558 1194 1564 1195
rect 1558 1190 1559 1194
rect 1563 1190 1564 1194
rect 1558 1189 1564 1190
rect 1590 1194 1596 1195
rect 1590 1190 1591 1194
rect 1595 1190 1596 1194
rect 1590 1189 1596 1190
rect 1622 1194 1628 1195
rect 1622 1190 1623 1194
rect 1627 1190 1628 1194
rect 1622 1189 1628 1190
rect 1654 1194 1660 1195
rect 1654 1190 1655 1194
rect 1659 1190 1660 1194
rect 1694 1192 1695 1196
rect 1699 1192 1700 1196
rect 1694 1191 1700 1192
rect 1654 1189 1660 1190
rect 838 1180 844 1181
rect 110 1179 116 1180
rect 110 1175 111 1179
rect 115 1175 116 1179
rect 110 1174 116 1175
rect 134 1177 140 1178
rect 134 1173 135 1177
rect 139 1173 140 1177
rect 134 1172 140 1173
rect 166 1177 172 1178
rect 166 1173 167 1177
rect 171 1173 172 1177
rect 166 1172 172 1173
rect 198 1177 204 1178
rect 198 1173 199 1177
rect 203 1173 204 1177
rect 198 1172 204 1173
rect 230 1177 236 1178
rect 230 1173 231 1177
rect 235 1173 236 1177
rect 230 1172 236 1173
rect 262 1177 268 1178
rect 262 1173 263 1177
rect 267 1173 268 1177
rect 262 1172 268 1173
rect 294 1177 300 1178
rect 294 1173 295 1177
rect 299 1173 300 1177
rect 294 1172 300 1173
rect 326 1177 332 1178
rect 326 1173 327 1177
rect 331 1173 332 1177
rect 326 1172 332 1173
rect 358 1177 364 1178
rect 358 1173 359 1177
rect 363 1173 364 1177
rect 358 1172 364 1173
rect 390 1177 396 1178
rect 390 1173 391 1177
rect 395 1173 396 1177
rect 390 1172 396 1173
rect 422 1177 428 1178
rect 422 1173 423 1177
rect 427 1173 428 1177
rect 422 1172 428 1173
rect 454 1177 460 1178
rect 454 1173 455 1177
rect 459 1173 460 1177
rect 454 1172 460 1173
rect 486 1177 492 1178
rect 486 1173 487 1177
rect 491 1173 492 1177
rect 486 1172 492 1173
rect 518 1177 524 1178
rect 518 1173 519 1177
rect 523 1173 524 1177
rect 518 1172 524 1173
rect 550 1177 556 1178
rect 550 1173 551 1177
rect 555 1173 556 1177
rect 550 1172 556 1173
rect 582 1177 588 1178
rect 582 1173 583 1177
rect 587 1173 588 1177
rect 582 1172 588 1173
rect 614 1177 620 1178
rect 614 1173 615 1177
rect 619 1173 620 1177
rect 614 1172 620 1173
rect 646 1177 652 1178
rect 646 1173 647 1177
rect 651 1173 652 1177
rect 646 1172 652 1173
rect 678 1177 684 1178
rect 678 1173 679 1177
rect 683 1173 684 1177
rect 678 1172 684 1173
rect 710 1177 716 1178
rect 710 1173 711 1177
rect 715 1173 716 1177
rect 710 1172 716 1173
rect 742 1177 748 1178
rect 742 1173 743 1177
rect 747 1173 748 1177
rect 838 1176 839 1180
rect 843 1176 844 1180
rect 1694 1179 1700 1180
rect 1126 1177 1132 1178
rect 838 1175 844 1176
rect 1006 1176 1012 1177
rect 742 1172 748 1173
rect 774 1172 780 1173
rect 774 1168 775 1172
rect 779 1168 780 1172
rect 1006 1172 1007 1176
rect 1011 1172 1012 1176
rect 1126 1173 1127 1177
rect 1131 1173 1132 1177
rect 1006 1171 1012 1172
rect 1086 1172 1092 1173
rect 1126 1172 1132 1173
rect 1158 1177 1164 1178
rect 1254 1177 1260 1178
rect 1158 1173 1159 1177
rect 1163 1173 1164 1177
rect 1158 1172 1164 1173
rect 1198 1176 1204 1177
rect 1198 1172 1199 1176
rect 1203 1172 1204 1176
rect 1254 1173 1255 1177
rect 1259 1173 1260 1177
rect 1254 1172 1260 1173
rect 1342 1177 1348 1178
rect 1342 1173 1343 1177
rect 1347 1173 1348 1177
rect 1342 1172 1348 1173
rect 1374 1177 1380 1178
rect 1374 1173 1375 1177
rect 1379 1173 1380 1177
rect 1374 1172 1380 1173
rect 1406 1177 1412 1178
rect 1406 1173 1407 1177
rect 1411 1173 1412 1177
rect 1406 1172 1412 1173
rect 1438 1177 1444 1178
rect 1438 1173 1439 1177
rect 1443 1173 1444 1177
rect 1438 1172 1444 1173
rect 1478 1177 1484 1178
rect 1478 1173 1479 1177
rect 1483 1173 1484 1177
rect 1478 1172 1484 1173
rect 1518 1177 1524 1178
rect 1518 1173 1519 1177
rect 1523 1173 1524 1177
rect 1518 1172 1524 1173
rect 1558 1177 1564 1178
rect 1558 1173 1559 1177
rect 1563 1173 1564 1177
rect 1558 1172 1564 1173
rect 1590 1177 1596 1178
rect 1590 1173 1591 1177
rect 1595 1173 1596 1177
rect 1590 1172 1596 1173
rect 1622 1177 1628 1178
rect 1622 1173 1623 1177
rect 1627 1173 1628 1177
rect 1622 1172 1628 1173
rect 1654 1177 1660 1178
rect 1654 1173 1655 1177
rect 1659 1173 1660 1177
rect 1694 1175 1695 1179
rect 1699 1175 1700 1179
rect 1694 1174 1700 1175
rect 1654 1172 1660 1173
rect 774 1167 780 1168
rect 974 1170 980 1171
rect 974 1166 975 1170
rect 979 1166 980 1170
rect 1086 1168 1087 1172
rect 1091 1168 1092 1172
rect 1198 1171 1204 1172
rect 1086 1167 1092 1168
rect 1310 1170 1316 1171
rect 974 1165 980 1166
rect 1310 1166 1311 1170
rect 1315 1166 1316 1170
rect 1310 1165 1316 1166
rect 1246 1128 1252 1129
rect 846 1126 852 1127
rect 582 1124 588 1125
rect 134 1123 140 1124
rect 110 1121 116 1122
rect 110 1117 111 1121
rect 115 1117 116 1121
rect 134 1119 135 1123
rect 139 1119 140 1123
rect 134 1118 140 1119
rect 166 1123 172 1124
rect 166 1119 167 1123
rect 171 1119 172 1123
rect 166 1118 172 1119
rect 198 1123 204 1124
rect 198 1119 199 1123
rect 203 1119 204 1123
rect 198 1118 204 1119
rect 230 1123 236 1124
rect 230 1119 231 1123
rect 235 1119 236 1123
rect 230 1118 236 1119
rect 262 1123 268 1124
rect 262 1119 263 1123
rect 267 1119 268 1123
rect 262 1118 268 1119
rect 294 1123 300 1124
rect 294 1119 295 1123
rect 299 1119 300 1123
rect 294 1118 300 1119
rect 326 1123 332 1124
rect 326 1119 327 1123
rect 331 1119 332 1123
rect 326 1118 332 1119
rect 358 1123 364 1124
rect 358 1119 359 1123
rect 363 1119 364 1123
rect 358 1118 364 1119
rect 390 1123 396 1124
rect 390 1119 391 1123
rect 395 1119 396 1123
rect 390 1118 396 1119
rect 422 1123 428 1124
rect 422 1119 423 1123
rect 427 1119 428 1123
rect 422 1118 428 1119
rect 454 1123 460 1124
rect 454 1119 455 1123
rect 459 1119 460 1123
rect 454 1118 460 1119
rect 486 1123 492 1124
rect 486 1119 487 1123
rect 491 1119 492 1123
rect 486 1118 492 1119
rect 518 1123 524 1124
rect 518 1119 519 1123
rect 523 1119 524 1123
rect 518 1118 524 1119
rect 550 1123 556 1124
rect 550 1119 551 1123
rect 555 1119 556 1123
rect 582 1120 583 1124
rect 587 1120 588 1124
rect 798 1124 804 1125
rect 582 1119 588 1120
rect 686 1120 692 1121
rect 550 1118 556 1119
rect 110 1116 116 1117
rect 686 1116 687 1120
rect 691 1116 692 1120
rect 798 1120 799 1124
rect 803 1120 804 1124
rect 846 1122 847 1126
rect 851 1122 852 1126
rect 998 1124 1004 1125
rect 1094 1124 1100 1125
rect 1166 1124 1172 1125
rect 846 1121 852 1122
rect 934 1123 940 1124
rect 798 1119 804 1120
rect 934 1119 935 1123
rect 939 1119 940 1123
rect 934 1118 940 1119
rect 966 1123 972 1124
rect 966 1119 967 1123
rect 971 1119 972 1123
rect 998 1120 999 1124
rect 1003 1120 1004 1124
rect 998 1119 1004 1120
rect 1030 1123 1036 1124
rect 1030 1119 1031 1123
rect 1035 1119 1036 1123
rect 966 1118 972 1119
rect 1030 1118 1036 1119
rect 1062 1123 1068 1124
rect 1062 1119 1063 1123
rect 1067 1119 1068 1123
rect 1094 1120 1095 1124
rect 1099 1120 1100 1124
rect 1094 1119 1100 1120
rect 1134 1123 1140 1124
rect 1134 1119 1135 1123
rect 1139 1119 1140 1123
rect 1166 1120 1167 1124
rect 1171 1120 1172 1124
rect 1246 1124 1247 1128
rect 1251 1124 1252 1128
rect 1334 1126 1340 1127
rect 1246 1123 1252 1124
rect 1286 1123 1292 1124
rect 1166 1119 1172 1120
rect 1286 1119 1287 1123
rect 1291 1119 1292 1123
rect 1334 1122 1335 1126
rect 1339 1122 1340 1126
rect 1334 1121 1340 1122
rect 1422 1123 1428 1124
rect 1062 1118 1068 1119
rect 1134 1118 1140 1119
rect 1286 1118 1292 1119
rect 1422 1119 1423 1123
rect 1427 1119 1428 1123
rect 1422 1118 1428 1119
rect 1454 1123 1460 1124
rect 1454 1119 1455 1123
rect 1459 1119 1460 1123
rect 1454 1118 1460 1119
rect 1486 1123 1492 1124
rect 1486 1119 1487 1123
rect 1491 1119 1492 1123
rect 1486 1118 1492 1119
rect 1518 1123 1524 1124
rect 1518 1119 1519 1123
rect 1523 1119 1524 1123
rect 1518 1118 1524 1119
rect 1558 1123 1564 1124
rect 1558 1119 1559 1123
rect 1563 1119 1564 1123
rect 1558 1118 1564 1119
rect 1590 1123 1596 1124
rect 1590 1119 1591 1123
rect 1595 1119 1596 1123
rect 1590 1118 1596 1119
rect 1622 1123 1628 1124
rect 1622 1119 1623 1123
rect 1627 1119 1628 1123
rect 1622 1118 1628 1119
rect 1654 1123 1660 1124
rect 1654 1119 1655 1123
rect 1659 1119 1660 1123
rect 1654 1118 1660 1119
rect 1694 1121 1700 1122
rect 1694 1117 1695 1121
rect 1699 1117 1700 1121
rect 1694 1116 1700 1117
rect 686 1115 692 1116
rect 134 1106 140 1107
rect 110 1104 116 1105
rect 110 1100 111 1104
rect 115 1100 116 1104
rect 134 1102 135 1106
rect 139 1102 140 1106
rect 134 1101 140 1102
rect 166 1106 172 1107
rect 166 1102 167 1106
rect 171 1102 172 1106
rect 166 1101 172 1102
rect 198 1106 204 1107
rect 198 1102 199 1106
rect 203 1102 204 1106
rect 198 1101 204 1102
rect 230 1106 236 1107
rect 230 1102 231 1106
rect 235 1102 236 1106
rect 230 1101 236 1102
rect 262 1106 268 1107
rect 262 1102 263 1106
rect 267 1102 268 1106
rect 262 1101 268 1102
rect 294 1106 300 1107
rect 294 1102 295 1106
rect 299 1102 300 1106
rect 294 1101 300 1102
rect 326 1106 332 1107
rect 326 1102 327 1106
rect 331 1102 332 1106
rect 326 1101 332 1102
rect 358 1106 364 1107
rect 358 1102 359 1106
rect 363 1102 364 1106
rect 358 1101 364 1102
rect 390 1106 396 1107
rect 390 1102 391 1106
rect 395 1102 396 1106
rect 390 1101 396 1102
rect 422 1106 428 1107
rect 422 1102 423 1106
rect 427 1102 428 1106
rect 422 1101 428 1102
rect 454 1106 460 1107
rect 454 1102 455 1106
rect 459 1102 460 1106
rect 454 1101 460 1102
rect 486 1106 492 1107
rect 486 1102 487 1106
rect 491 1102 492 1106
rect 486 1101 492 1102
rect 518 1106 524 1107
rect 518 1102 519 1106
rect 523 1102 524 1106
rect 518 1101 524 1102
rect 550 1106 556 1107
rect 934 1106 940 1107
rect 550 1102 551 1106
rect 555 1102 556 1106
rect 550 1101 556 1102
rect 658 1105 664 1106
rect 658 1101 659 1105
rect 663 1101 664 1105
rect 934 1102 935 1106
rect 939 1102 940 1106
rect 658 1100 664 1101
rect 798 1101 804 1102
rect 934 1101 940 1102
rect 966 1106 972 1107
rect 966 1102 967 1106
rect 971 1102 972 1106
rect 1030 1106 1036 1107
rect 1030 1102 1031 1106
rect 1035 1102 1036 1106
rect 966 1101 972 1102
rect 998 1101 1004 1102
rect 1030 1101 1036 1102
rect 1062 1106 1068 1107
rect 1062 1102 1063 1106
rect 1067 1102 1068 1106
rect 1062 1101 1068 1102
rect 1134 1106 1140 1107
rect 1134 1102 1135 1106
rect 1139 1102 1140 1106
rect 1134 1101 1140 1102
rect 1286 1106 1292 1107
rect 1286 1102 1287 1106
rect 1291 1102 1292 1106
rect 1286 1101 1292 1102
rect 1422 1106 1428 1107
rect 1422 1102 1423 1106
rect 1427 1102 1428 1106
rect 1422 1101 1428 1102
rect 1454 1106 1460 1107
rect 1454 1102 1455 1106
rect 1459 1102 1460 1106
rect 1454 1101 1460 1102
rect 1486 1106 1492 1107
rect 1486 1102 1487 1106
rect 1491 1102 1492 1106
rect 1486 1101 1492 1102
rect 1518 1106 1524 1107
rect 1518 1102 1519 1106
rect 1523 1102 1524 1106
rect 1518 1101 1524 1102
rect 1558 1106 1564 1107
rect 1558 1102 1559 1106
rect 1563 1102 1564 1106
rect 1558 1101 1564 1102
rect 1590 1106 1596 1107
rect 1590 1102 1591 1106
rect 1595 1102 1596 1106
rect 1590 1101 1596 1102
rect 1622 1106 1628 1107
rect 1622 1102 1623 1106
rect 1627 1102 1628 1106
rect 1622 1101 1628 1102
rect 1654 1106 1660 1107
rect 1654 1102 1655 1106
rect 1659 1102 1660 1106
rect 1654 1101 1660 1102
rect 1694 1104 1700 1105
rect 110 1099 116 1100
rect 798 1097 799 1101
rect 803 1097 804 1101
rect 798 1096 804 1097
rect 998 1097 999 1101
rect 1003 1097 1004 1101
rect 1694 1100 1695 1104
rect 1699 1100 1700 1104
rect 1694 1099 1700 1100
rect 998 1096 1004 1097
rect 1094 1096 1100 1097
rect 1094 1092 1095 1096
rect 1099 1092 1100 1096
rect 1094 1091 1100 1092
rect 590 1086 596 1087
rect 1174 1086 1180 1087
rect 590 1082 591 1086
rect 595 1082 596 1086
rect 590 1081 596 1082
rect 846 1085 852 1086
rect 846 1081 847 1085
rect 851 1081 852 1085
rect 1174 1082 1175 1086
rect 1179 1082 1180 1086
rect 1334 1085 1340 1086
rect 1174 1081 1180 1082
rect 1246 1081 1252 1082
rect 846 1080 852 1081
rect 1246 1077 1247 1081
rect 1251 1077 1252 1081
rect 1334 1081 1335 1085
rect 1339 1081 1340 1085
rect 1334 1080 1340 1081
rect 1246 1076 1252 1077
rect 502 1019 508 1020
rect 502 1015 503 1019
rect 507 1015 508 1019
rect 406 1014 412 1015
rect 502 1014 508 1015
rect 582 1015 588 1016
rect 406 1010 407 1014
rect 411 1010 412 1014
rect 582 1011 583 1015
rect 587 1011 588 1015
rect 582 1010 588 1011
rect 710 1015 716 1016
rect 710 1011 711 1015
rect 715 1011 716 1015
rect 710 1010 716 1011
rect 406 1009 412 1010
rect 822 1009 828 1010
rect 822 1005 823 1009
rect 827 1005 828 1009
rect 822 1004 828 1005
rect 974 1009 980 1010
rect 974 1005 975 1009
rect 979 1005 980 1009
rect 974 1004 980 1005
rect 1062 1004 1068 1005
rect 1062 1000 1063 1004
rect 1067 1000 1068 1004
rect 1062 999 1068 1000
rect 1198 1004 1204 1005
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1198 999 1204 1000
rect 1326 1004 1332 1005
rect 1326 1000 1327 1004
rect 1331 1000 1332 1004
rect 1326 999 1332 1000
rect 1366 1004 1372 1005
rect 1366 1000 1367 1004
rect 1371 1000 1372 1004
rect 1366 999 1372 1000
rect 326 997 332 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 134 994 140 995
rect 134 990 135 994
rect 139 990 140 994
rect 134 989 140 990
rect 166 994 172 995
rect 166 990 167 994
rect 171 990 172 994
rect 166 989 172 990
rect 198 994 204 995
rect 198 990 199 994
rect 203 990 204 994
rect 198 989 204 990
rect 230 994 236 995
rect 230 990 231 994
rect 235 990 236 994
rect 230 989 236 990
rect 262 994 268 995
rect 262 990 263 994
rect 267 990 268 994
rect 326 993 327 997
rect 331 993 332 997
rect 1118 997 1124 998
rect 326 992 332 993
rect 918 994 924 995
rect 262 989 268 990
rect 918 990 919 994
rect 923 990 924 994
rect 1118 993 1119 997
rect 1123 993 1124 997
rect 1246 997 1252 998
rect 1118 992 1124 993
rect 1166 994 1172 995
rect 918 989 924 990
rect 1166 990 1167 994
rect 1171 990 1172 994
rect 1246 993 1247 997
rect 1251 993 1252 997
rect 1694 996 1700 997
rect 1246 992 1252 993
rect 1294 994 1300 995
rect 1166 989 1172 990
rect 1294 990 1295 994
rect 1299 990 1300 994
rect 1294 989 1300 990
rect 1406 994 1412 995
rect 1406 990 1407 994
rect 1411 990 1412 994
rect 1406 989 1412 990
rect 1438 994 1444 995
rect 1438 990 1439 994
rect 1443 990 1444 994
rect 1438 989 1444 990
rect 1478 994 1484 995
rect 1478 990 1479 994
rect 1483 990 1484 994
rect 1478 989 1484 990
rect 1518 994 1524 995
rect 1518 990 1519 994
rect 1523 990 1524 994
rect 1518 989 1524 990
rect 1558 994 1564 995
rect 1558 990 1559 994
rect 1563 990 1564 994
rect 1558 989 1564 990
rect 1590 994 1596 995
rect 1590 990 1591 994
rect 1595 990 1596 994
rect 1590 989 1596 990
rect 1622 994 1628 995
rect 1622 990 1623 994
rect 1627 990 1628 994
rect 1622 989 1628 990
rect 1654 994 1660 995
rect 1654 990 1655 994
rect 1659 990 1660 994
rect 1694 992 1695 996
rect 1699 992 1700 996
rect 1694 991 1700 992
rect 1654 989 1660 990
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 1694 979 1700 980
rect 110 974 116 975
rect 134 977 140 978
rect 134 973 135 977
rect 139 973 140 977
rect 134 972 140 973
rect 166 977 172 978
rect 166 973 167 977
rect 171 973 172 977
rect 166 972 172 973
rect 198 977 204 978
rect 198 973 199 977
rect 203 973 204 977
rect 198 972 204 973
rect 230 977 236 978
rect 230 973 231 977
rect 235 973 236 977
rect 230 972 236 973
rect 262 977 268 978
rect 918 977 924 978
rect 1166 977 1172 978
rect 1294 977 1300 978
rect 1406 977 1412 978
rect 262 973 263 977
rect 267 973 268 977
rect 262 972 268 973
rect 398 976 404 977
rect 398 972 399 976
rect 403 972 404 976
rect 582 974 588 975
rect 398 971 404 972
rect 502 972 508 973
rect 342 970 348 971
rect 342 966 343 970
rect 347 966 348 970
rect 502 968 503 972
rect 507 968 508 972
rect 582 970 583 974
rect 587 970 588 974
rect 582 969 588 970
rect 710 974 716 975
rect 710 970 711 974
rect 715 970 716 974
rect 918 973 919 977
rect 923 973 924 977
rect 918 972 924 973
rect 1062 976 1068 977
rect 1062 972 1063 976
rect 1067 972 1068 976
rect 1166 973 1167 977
rect 1171 973 1172 977
rect 1166 972 1172 973
rect 1198 976 1204 977
rect 1198 972 1199 976
rect 1203 972 1204 976
rect 1294 973 1295 977
rect 1299 973 1300 977
rect 1294 972 1300 973
rect 1326 976 1332 977
rect 1326 972 1327 976
rect 1331 972 1332 976
rect 1062 971 1068 972
rect 1198 971 1204 972
rect 1326 971 1332 972
rect 1366 976 1372 977
rect 1366 972 1367 976
rect 1371 972 1372 976
rect 1406 973 1407 977
rect 1411 973 1412 977
rect 1406 972 1412 973
rect 1438 977 1444 978
rect 1438 973 1439 977
rect 1443 973 1444 977
rect 1438 972 1444 973
rect 1478 977 1484 978
rect 1478 973 1479 977
rect 1483 973 1484 977
rect 1478 972 1484 973
rect 1518 977 1524 978
rect 1518 973 1519 977
rect 1523 973 1524 977
rect 1518 972 1524 973
rect 1558 977 1564 978
rect 1558 973 1559 977
rect 1563 973 1564 977
rect 1558 972 1564 973
rect 1590 977 1596 978
rect 1590 973 1591 977
rect 1595 973 1596 977
rect 1590 972 1596 973
rect 1622 977 1628 978
rect 1622 973 1623 977
rect 1627 973 1628 977
rect 1622 972 1628 973
rect 1654 977 1660 978
rect 1654 973 1655 977
rect 1659 973 1660 977
rect 1694 975 1695 979
rect 1699 975 1700 979
rect 1694 974 1700 975
rect 1654 972 1660 973
rect 1366 971 1372 972
rect 1134 970 1140 971
rect 710 969 716 970
rect 814 969 820 970
rect 502 967 508 968
rect 342 965 348 966
rect 814 965 815 969
rect 819 965 820 969
rect 814 964 820 965
rect 966 969 972 970
rect 966 965 967 969
rect 971 965 972 969
rect 1134 966 1135 970
rect 1139 966 1140 970
rect 1134 965 1140 966
rect 1262 970 1268 971
rect 1262 966 1263 970
rect 1267 966 1268 970
rect 1262 965 1268 966
rect 966 964 972 965
rect 1390 930 1396 931
rect 278 928 284 929
rect 198 924 204 925
rect 134 923 140 924
rect 110 921 116 922
rect 110 917 111 921
rect 115 917 116 921
rect 134 919 135 923
rect 139 919 140 923
rect 134 918 140 919
rect 166 923 172 924
rect 166 919 167 923
rect 171 919 172 923
rect 198 920 199 924
rect 203 920 204 924
rect 278 924 279 928
rect 283 924 284 928
rect 398 928 404 929
rect 278 923 284 924
rect 318 924 324 925
rect 198 919 204 920
rect 318 920 319 924
rect 323 920 324 924
rect 398 924 399 928
rect 403 924 404 928
rect 398 923 404 924
rect 590 926 596 927
rect 590 922 591 926
rect 595 922 596 926
rect 726 926 732 927
rect 590 921 596 922
rect 678 924 684 925
rect 318 919 324 920
rect 462 920 468 921
rect 166 918 172 919
rect 110 916 116 917
rect 462 916 463 920
rect 467 916 468 920
rect 678 920 679 924
rect 683 920 684 924
rect 726 922 727 926
rect 731 922 732 926
rect 862 926 868 927
rect 726 921 732 922
rect 814 923 820 924
rect 678 919 684 920
rect 814 919 815 923
rect 819 919 820 923
rect 862 922 863 926
rect 867 922 868 926
rect 1390 926 1391 930
rect 1395 926 1396 930
rect 1390 925 1396 926
rect 982 924 988 925
rect 1070 924 1076 925
rect 1142 924 1148 925
rect 1270 924 1276 925
rect 1454 924 1460 925
rect 862 921 868 922
rect 950 923 956 924
rect 814 918 820 919
rect 950 919 951 923
rect 955 919 956 923
rect 982 920 983 924
rect 987 920 988 924
rect 982 919 988 920
rect 1038 923 1044 924
rect 1038 919 1039 923
rect 1043 919 1044 923
rect 1070 920 1071 924
rect 1075 920 1076 924
rect 1070 919 1076 920
rect 1110 923 1116 924
rect 1110 919 1111 923
rect 1115 919 1116 923
rect 1142 920 1143 924
rect 1147 920 1148 924
rect 1142 919 1148 920
rect 1238 923 1244 924
rect 1238 919 1239 923
rect 1243 919 1244 923
rect 1270 920 1271 924
rect 1275 920 1276 924
rect 1270 919 1276 920
rect 1422 923 1428 924
rect 1422 919 1423 923
rect 1427 919 1428 923
rect 1454 920 1455 924
rect 1459 920 1460 924
rect 1454 919 1460 920
rect 1518 923 1524 924
rect 1518 919 1519 923
rect 1523 919 1524 923
rect 950 918 956 919
rect 1038 918 1044 919
rect 1110 918 1116 919
rect 1238 918 1244 919
rect 1422 918 1428 919
rect 1518 918 1524 919
rect 1558 923 1564 924
rect 1558 919 1559 923
rect 1563 919 1564 923
rect 1558 918 1564 919
rect 1590 923 1596 924
rect 1590 919 1591 923
rect 1595 919 1596 923
rect 1590 918 1596 919
rect 1622 923 1628 924
rect 1622 919 1623 923
rect 1627 919 1628 923
rect 1622 918 1628 919
rect 1654 923 1660 924
rect 1654 919 1655 923
rect 1659 919 1660 923
rect 1654 918 1660 919
rect 1694 921 1700 922
rect 1694 917 1695 921
rect 1699 917 1700 921
rect 1694 916 1700 917
rect 462 915 468 916
rect 134 906 140 907
rect 110 904 116 905
rect 110 900 111 904
rect 115 900 116 904
rect 134 902 135 906
rect 139 902 140 906
rect 134 901 140 902
rect 166 906 172 907
rect 814 906 820 907
rect 166 902 167 906
rect 171 902 172 906
rect 166 901 172 902
rect 434 905 440 906
rect 434 901 435 905
rect 439 901 440 905
rect 814 902 815 906
rect 819 902 820 906
rect 434 900 440 901
rect 678 901 684 902
rect 814 901 820 902
rect 950 906 956 907
rect 950 902 951 906
rect 955 902 956 906
rect 1038 906 1044 907
rect 1422 906 1428 907
rect 950 901 956 902
rect 998 903 1004 904
rect 110 899 116 900
rect 678 897 679 901
rect 683 897 684 901
rect 998 899 999 903
rect 1003 899 1004 903
rect 1038 902 1039 906
rect 1043 902 1044 906
rect 1038 901 1044 902
rect 1110 905 1116 906
rect 1110 901 1111 905
rect 1115 901 1116 905
rect 1110 900 1116 901
rect 1142 905 1148 906
rect 1142 901 1143 905
rect 1147 901 1148 905
rect 1142 900 1148 901
rect 1238 905 1244 906
rect 1238 901 1239 905
rect 1243 901 1244 905
rect 1238 900 1244 901
rect 1270 905 1276 906
rect 1270 901 1271 905
rect 1275 901 1276 905
rect 1270 900 1276 901
rect 1374 903 1380 904
rect 998 898 1004 899
rect 1374 899 1375 903
rect 1379 899 1380 903
rect 1422 902 1423 906
rect 1427 902 1428 906
rect 1518 906 1524 907
rect 1422 901 1428 902
rect 1470 903 1476 904
rect 1374 898 1380 899
rect 1470 899 1471 903
rect 1475 899 1476 903
rect 1518 902 1519 906
rect 1523 902 1524 906
rect 1518 901 1524 902
rect 1558 906 1564 907
rect 1558 902 1559 906
rect 1563 902 1564 906
rect 1558 901 1564 902
rect 1590 906 1596 907
rect 1590 902 1591 906
rect 1595 902 1596 906
rect 1590 901 1596 902
rect 1622 906 1628 907
rect 1622 902 1623 906
rect 1627 902 1628 906
rect 1622 901 1628 902
rect 1654 906 1660 907
rect 1654 902 1655 906
rect 1659 902 1660 906
rect 1654 901 1660 902
rect 1694 904 1700 905
rect 1694 900 1695 904
rect 1699 900 1700 904
rect 1694 899 1700 900
rect 1470 898 1476 899
rect 678 896 684 897
rect 1070 896 1076 897
rect 1070 892 1071 896
rect 1075 892 1076 896
rect 1070 891 1076 892
rect 206 886 212 887
rect 206 882 207 886
rect 211 882 212 886
rect 326 886 332 887
rect 326 882 327 886
rect 331 882 332 886
rect 590 885 596 886
rect 206 881 212 882
rect 278 881 284 882
rect 326 881 332 882
rect 398 881 404 882
rect 278 877 279 881
rect 283 877 284 881
rect 278 876 284 877
rect 398 877 399 881
rect 403 877 404 881
rect 590 881 591 885
rect 595 881 596 885
rect 590 880 596 881
rect 726 885 732 886
rect 726 881 727 885
rect 731 881 732 885
rect 726 880 732 881
rect 862 885 868 886
rect 862 881 863 885
rect 867 881 868 885
rect 862 880 868 881
rect 398 876 404 877
rect 230 823 236 824
rect 230 819 231 823
rect 235 819 236 823
rect 230 818 236 819
rect 406 823 412 824
rect 406 819 407 823
rect 411 819 412 823
rect 406 818 412 819
rect 814 823 820 824
rect 814 819 815 823
rect 819 819 820 823
rect 814 818 820 819
rect 662 817 668 818
rect 662 813 663 817
rect 667 813 668 817
rect 662 812 668 813
rect 1422 812 1428 813
rect 1422 808 1423 812
rect 1427 808 1428 812
rect 950 807 956 808
rect 1422 807 1428 808
rect 1470 812 1476 813
rect 1470 808 1471 812
rect 1475 808 1476 812
rect 1470 807 1476 808
rect 110 804 116 805
rect 110 800 111 804
rect 115 800 116 804
rect 950 803 951 807
rect 955 803 956 807
rect 110 799 116 800
rect 134 802 140 803
rect 134 798 135 802
rect 139 798 140 802
rect 134 797 140 798
rect 558 802 564 803
rect 950 802 956 803
rect 1030 805 1036 806
rect 558 798 559 802
rect 563 798 564 802
rect 1030 801 1031 805
rect 1035 801 1036 805
rect 1166 805 1172 806
rect 1030 800 1036 801
rect 1102 802 1108 803
rect 558 797 564 798
rect 1102 798 1103 802
rect 1107 798 1108 802
rect 1166 801 1167 805
rect 1171 801 1172 805
rect 1166 800 1172 801
rect 1246 805 1252 806
rect 1246 801 1247 805
rect 1251 801 1252 805
rect 1694 804 1700 805
rect 1246 800 1252 801
rect 1294 803 1300 804
rect 1294 799 1295 803
rect 1299 799 1300 803
rect 1294 798 1300 799
rect 1326 803 1332 804
rect 1326 799 1327 803
rect 1331 799 1332 803
rect 1326 798 1332 799
rect 1518 802 1524 803
rect 1518 798 1519 802
rect 1523 798 1524 802
rect 1102 797 1108 798
rect 1518 797 1524 798
rect 1558 802 1564 803
rect 1558 798 1559 802
rect 1563 798 1564 802
rect 1558 797 1564 798
rect 1590 802 1596 803
rect 1590 798 1591 802
rect 1595 798 1596 802
rect 1590 797 1596 798
rect 1622 802 1628 803
rect 1622 798 1623 802
rect 1627 798 1628 802
rect 1622 797 1628 798
rect 1654 802 1660 803
rect 1654 798 1655 802
rect 1659 798 1660 802
rect 1694 800 1695 804
rect 1699 800 1700 804
rect 1694 799 1700 800
rect 1654 797 1660 798
rect 110 787 116 788
rect 110 783 111 787
rect 115 783 116 787
rect 1694 787 1700 788
rect 110 782 116 783
rect 134 785 140 786
rect 134 781 135 785
rect 139 781 140 785
rect 558 785 564 786
rect 1102 785 1108 786
rect 1294 785 1300 786
rect 1518 785 1524 786
rect 134 780 140 781
rect 230 782 236 783
rect 230 778 231 782
rect 235 778 236 782
rect 230 777 236 778
rect 406 782 412 783
rect 406 778 407 782
rect 411 778 412 782
rect 558 781 559 785
rect 563 781 564 785
rect 950 784 956 785
rect 558 780 564 781
rect 814 782 820 783
rect 814 778 815 782
rect 819 778 820 782
rect 950 780 951 784
rect 955 780 956 784
rect 950 779 956 780
rect 1014 784 1020 785
rect 1014 780 1015 784
rect 1019 780 1020 784
rect 1102 781 1103 785
rect 1107 781 1108 785
rect 1102 780 1108 781
rect 1230 784 1236 785
rect 1230 780 1231 784
rect 1235 780 1236 784
rect 1294 781 1295 785
rect 1299 781 1300 785
rect 1294 780 1300 781
rect 1326 784 1332 785
rect 1326 780 1327 784
rect 1331 780 1332 784
rect 1014 779 1020 780
rect 1230 779 1236 780
rect 1326 779 1332 780
rect 1422 784 1428 785
rect 1422 780 1423 784
rect 1427 780 1428 784
rect 1422 779 1428 780
rect 1470 784 1476 785
rect 1470 780 1471 784
rect 1475 780 1476 784
rect 1518 781 1519 785
rect 1523 781 1524 785
rect 1518 780 1524 781
rect 1558 785 1564 786
rect 1558 781 1559 785
rect 1563 781 1564 785
rect 1558 780 1564 781
rect 1590 785 1596 786
rect 1590 781 1591 785
rect 1595 781 1596 785
rect 1590 780 1596 781
rect 1622 785 1628 786
rect 1622 781 1623 785
rect 1627 781 1628 785
rect 1622 780 1628 781
rect 1654 785 1660 786
rect 1654 781 1655 785
rect 1659 781 1660 785
rect 1694 783 1695 787
rect 1699 783 1700 787
rect 1694 782 1700 783
rect 1654 780 1660 781
rect 1470 779 1476 780
rect 406 777 412 778
rect 654 777 660 778
rect 814 777 820 778
rect 1182 778 1188 779
rect 654 773 655 777
rect 659 773 660 777
rect 1182 774 1183 778
rect 1187 774 1188 778
rect 1182 773 1188 774
rect 654 772 660 773
rect 766 735 772 736
rect 214 732 220 733
rect 134 728 140 729
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 134 724 135 728
rect 139 724 140 728
rect 214 728 215 732
rect 219 728 220 732
rect 390 732 396 733
rect 214 727 220 728
rect 286 730 292 731
rect 286 726 287 730
rect 291 726 292 730
rect 390 728 391 732
rect 395 728 396 732
rect 766 731 767 735
rect 771 731 772 735
rect 998 735 1004 736
rect 998 731 999 735
rect 1003 731 1004 735
rect 390 727 396 728
rect 614 730 620 731
rect 766 730 772 731
rect 910 730 916 731
rect 998 730 1004 731
rect 1166 732 1172 733
rect 286 725 292 726
rect 614 726 615 730
rect 619 726 620 730
rect 614 725 620 726
rect 718 728 724 729
rect 134 723 140 724
rect 470 724 476 725
rect 110 720 116 721
rect 470 720 471 724
rect 475 720 476 724
rect 718 724 719 728
rect 723 724 724 728
rect 718 723 724 724
rect 862 727 868 728
rect 862 723 863 727
rect 867 723 868 727
rect 910 726 911 730
rect 915 726 916 730
rect 910 725 916 726
rect 1086 728 1092 729
rect 1086 724 1087 728
rect 1091 724 1092 728
rect 1166 728 1167 732
rect 1171 728 1172 732
rect 1166 727 1172 728
rect 1206 728 1212 729
rect 1086 723 1092 724
rect 1206 724 1207 728
rect 1211 724 1212 728
rect 1206 723 1212 724
rect 1246 727 1252 728
rect 1246 723 1247 727
rect 1251 723 1252 727
rect 862 722 868 723
rect 1246 722 1252 723
rect 1278 727 1284 728
rect 1278 723 1279 727
rect 1283 723 1284 727
rect 1278 722 1284 723
rect 1310 727 1316 728
rect 1310 723 1311 727
rect 1315 723 1316 727
rect 1310 722 1316 723
rect 1342 727 1348 728
rect 1342 723 1343 727
rect 1347 723 1348 727
rect 1342 722 1348 723
rect 1374 727 1380 728
rect 1374 723 1375 727
rect 1379 723 1380 727
rect 1374 722 1380 723
rect 1406 727 1412 728
rect 1406 723 1407 727
rect 1411 723 1412 727
rect 1406 722 1412 723
rect 1438 727 1444 728
rect 1438 723 1439 727
rect 1443 723 1444 727
rect 1438 722 1444 723
rect 1478 727 1484 728
rect 1478 723 1479 727
rect 1483 723 1484 727
rect 1478 722 1484 723
rect 1518 727 1524 728
rect 1518 723 1519 727
rect 1523 723 1524 727
rect 1518 722 1524 723
rect 1558 727 1564 728
rect 1558 723 1559 727
rect 1563 723 1564 727
rect 1558 722 1564 723
rect 1590 727 1596 728
rect 1590 723 1591 727
rect 1595 723 1596 727
rect 1590 722 1596 723
rect 1622 727 1628 728
rect 1622 723 1623 727
rect 1627 723 1628 727
rect 1622 722 1628 723
rect 1654 727 1660 728
rect 1654 723 1655 727
rect 1659 723 1660 727
rect 1654 722 1660 723
rect 1694 725 1700 726
rect 1694 721 1695 725
rect 1699 721 1700 725
rect 1694 720 1700 721
rect 470 719 476 720
rect 862 710 868 711
rect 442 709 448 710
rect 110 708 116 709
rect 110 704 111 708
rect 115 704 116 708
rect 442 705 443 709
rect 447 705 448 709
rect 862 706 863 710
rect 867 706 868 710
rect 442 704 448 705
rect 718 705 724 706
rect 862 705 868 706
rect 1246 710 1252 711
rect 1246 706 1247 710
rect 1251 706 1252 710
rect 1246 705 1252 706
rect 1278 710 1284 711
rect 1278 706 1279 710
rect 1283 706 1284 710
rect 1278 705 1284 706
rect 1310 710 1316 711
rect 1310 706 1311 710
rect 1315 706 1316 710
rect 1310 705 1316 706
rect 1342 710 1348 711
rect 1342 706 1343 710
rect 1347 706 1348 710
rect 1342 705 1348 706
rect 1374 710 1380 711
rect 1374 706 1375 710
rect 1379 706 1380 710
rect 1374 705 1380 706
rect 1406 710 1412 711
rect 1406 706 1407 710
rect 1411 706 1412 710
rect 1406 705 1412 706
rect 1438 710 1444 711
rect 1438 706 1439 710
rect 1443 706 1444 710
rect 1438 705 1444 706
rect 1478 710 1484 711
rect 1478 706 1479 710
rect 1483 706 1484 710
rect 1478 705 1484 706
rect 1518 710 1524 711
rect 1518 706 1519 710
rect 1523 706 1524 710
rect 1518 705 1524 706
rect 1558 710 1564 711
rect 1558 706 1559 710
rect 1563 706 1564 710
rect 1558 705 1564 706
rect 1590 710 1596 711
rect 1590 706 1591 710
rect 1595 706 1596 710
rect 1590 705 1596 706
rect 1622 710 1628 711
rect 1622 706 1623 710
rect 1627 706 1628 710
rect 1622 705 1628 706
rect 1654 710 1660 711
rect 1654 706 1655 710
rect 1659 706 1660 710
rect 1654 705 1660 706
rect 1694 708 1700 709
rect 110 703 116 704
rect 718 701 719 705
rect 723 701 724 705
rect 1694 704 1695 708
rect 1699 704 1700 708
rect 1694 703 1700 704
rect 718 700 724 701
rect 1206 700 1212 701
rect 1206 696 1207 700
rect 1211 696 1212 700
rect 774 695 780 696
rect 774 691 775 695
rect 779 691 780 695
rect 142 690 148 691
rect 774 690 780 691
rect 1006 695 1012 696
rect 1206 695 1212 696
rect 1006 691 1007 695
rect 1011 691 1012 695
rect 1006 690 1012 691
rect 1094 690 1100 691
rect 142 686 143 690
rect 147 686 148 690
rect 286 689 292 690
rect 142 685 148 686
rect 214 685 220 686
rect 214 681 215 685
rect 219 681 220 685
rect 286 685 287 689
rect 291 685 292 689
rect 614 689 620 690
rect 286 684 292 685
rect 390 685 396 686
rect 214 680 220 681
rect 390 681 391 685
rect 395 681 396 685
rect 614 685 615 689
rect 619 685 620 689
rect 614 684 620 685
rect 910 689 916 690
rect 910 685 911 689
rect 915 685 916 689
rect 1094 686 1095 690
rect 1099 686 1100 690
rect 1094 685 1100 686
rect 1166 685 1172 686
rect 910 684 916 685
rect 390 680 396 681
rect 1166 681 1167 685
rect 1171 681 1172 685
rect 1166 680 1172 681
rect 206 627 212 628
rect 206 623 207 627
rect 211 623 212 627
rect 902 627 908 628
rect 534 623 540 624
rect 206 622 212 623
rect 286 622 292 623
rect 286 618 287 622
rect 291 618 292 622
rect 286 617 292 618
rect 406 622 412 623
rect 406 618 407 622
rect 411 618 412 622
rect 534 619 535 623
rect 539 619 540 623
rect 534 618 540 619
rect 766 623 772 624
rect 766 619 767 623
rect 771 619 772 623
rect 902 623 903 627
rect 907 623 908 627
rect 1118 627 1124 628
rect 1118 623 1119 627
rect 1123 623 1124 627
rect 1334 627 1340 628
rect 1334 623 1335 627
rect 1339 623 1340 627
rect 902 622 908 623
rect 998 622 1004 623
rect 1118 622 1124 623
rect 1214 622 1220 623
rect 1334 622 1340 623
rect 766 618 772 619
rect 998 618 999 622
rect 1003 618 1004 622
rect 406 617 412 618
rect 998 617 1004 618
rect 1214 618 1215 622
rect 1219 618 1220 622
rect 1214 617 1220 618
rect 110 604 116 605
rect 110 600 111 604
rect 115 600 116 604
rect 1694 604 1700 605
rect 110 599 116 600
rect 134 602 140 603
rect 134 598 135 602
rect 139 598 140 602
rect 134 597 140 598
rect 166 602 172 603
rect 166 598 167 602
rect 171 598 172 602
rect 166 597 172 598
rect 670 602 676 603
rect 670 598 671 602
rect 675 598 676 602
rect 670 597 676 598
rect 1414 602 1420 603
rect 1414 598 1415 602
rect 1419 598 1420 602
rect 1414 597 1420 598
rect 1478 602 1484 603
rect 1478 598 1479 602
rect 1483 598 1484 602
rect 1478 597 1484 598
rect 1542 602 1548 603
rect 1542 598 1543 602
rect 1547 598 1548 602
rect 1542 597 1548 598
rect 1606 602 1612 603
rect 1606 598 1607 602
rect 1611 598 1612 602
rect 1606 597 1612 598
rect 1654 602 1660 603
rect 1654 598 1655 602
rect 1659 598 1660 602
rect 1694 600 1695 604
rect 1699 600 1700 604
rect 1694 599 1700 600
rect 1654 597 1660 598
rect 110 587 116 588
rect 110 583 111 587
rect 115 583 116 587
rect 1694 587 1700 588
rect 110 582 116 583
rect 134 585 140 586
rect 134 581 135 585
rect 139 581 140 585
rect 134 580 140 581
rect 166 585 172 586
rect 670 585 676 586
rect 1414 585 1420 586
rect 166 581 167 585
rect 171 581 172 585
rect 278 584 284 585
rect 166 580 172 581
rect 206 580 212 581
rect 206 576 207 580
rect 211 576 212 580
rect 278 580 279 584
rect 283 580 284 584
rect 278 579 284 580
rect 398 584 404 585
rect 398 580 399 584
rect 403 580 404 584
rect 398 579 404 580
rect 534 582 540 583
rect 534 578 535 582
rect 539 578 540 582
rect 670 581 671 585
rect 675 581 676 585
rect 990 584 996 585
rect 670 580 676 581
rect 766 582 772 583
rect 534 577 540 578
rect 766 578 767 582
rect 771 578 772 582
rect 766 577 772 578
rect 902 580 908 581
rect 206 575 212 576
rect 902 576 903 580
rect 907 576 908 580
rect 990 580 991 584
rect 995 580 996 584
rect 1206 584 1212 585
rect 990 579 996 580
rect 1118 580 1124 581
rect 902 575 908 576
rect 1118 576 1119 580
rect 1123 576 1124 580
rect 1206 580 1207 584
rect 1211 580 1212 584
rect 1414 581 1415 585
rect 1419 581 1420 585
rect 1206 579 1212 580
rect 1334 580 1340 581
rect 1414 580 1420 581
rect 1478 585 1484 586
rect 1478 581 1479 585
rect 1483 581 1484 585
rect 1478 580 1484 581
rect 1542 585 1548 586
rect 1542 581 1543 585
rect 1547 581 1548 585
rect 1542 580 1548 581
rect 1606 585 1612 586
rect 1606 581 1607 585
rect 1611 581 1612 585
rect 1606 580 1612 581
rect 1654 585 1660 586
rect 1654 581 1655 585
rect 1659 581 1660 585
rect 1694 583 1695 587
rect 1699 583 1700 587
rect 1694 582 1700 583
rect 1654 580 1660 581
rect 1118 575 1124 576
rect 1334 576 1335 580
rect 1339 576 1340 580
rect 1334 575 1340 576
rect 246 540 252 541
rect 166 536 172 537
rect 134 535 140 536
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 134 531 135 535
rect 139 531 140 535
rect 166 532 167 536
rect 171 532 172 536
rect 246 536 247 540
rect 251 536 252 540
rect 470 540 476 541
rect 246 535 252 536
rect 302 538 308 539
rect 302 534 303 538
rect 307 534 308 538
rect 302 533 308 534
rect 390 536 396 537
rect 166 531 172 532
rect 390 532 391 536
rect 395 532 396 536
rect 470 536 471 540
rect 475 536 476 540
rect 726 540 732 541
rect 470 535 476 536
rect 646 536 652 537
rect 390 531 396 532
rect 534 532 540 533
rect 134 530 140 531
rect 110 528 116 529
rect 534 528 535 532
rect 539 528 540 532
rect 646 532 647 536
rect 651 532 652 536
rect 726 536 727 540
rect 731 536 732 540
rect 870 540 876 541
rect 726 535 732 536
rect 774 536 780 537
rect 646 531 652 532
rect 774 532 775 536
rect 779 532 780 536
rect 870 536 871 540
rect 875 536 876 540
rect 1030 540 1036 541
rect 870 535 876 536
rect 926 536 932 537
rect 774 531 780 532
rect 926 532 927 536
rect 931 532 932 536
rect 1030 536 1031 540
rect 1035 536 1036 540
rect 1198 540 1204 541
rect 1030 535 1036 536
rect 1094 536 1100 537
rect 926 531 932 532
rect 1094 532 1095 536
rect 1099 532 1100 536
rect 1198 536 1199 540
rect 1203 536 1204 540
rect 1198 535 1204 536
rect 1422 535 1428 536
rect 1094 531 1100 532
rect 1286 532 1292 533
rect 534 527 540 528
rect 1286 528 1287 532
rect 1291 528 1292 532
rect 1422 531 1423 535
rect 1427 531 1428 535
rect 1422 530 1428 531
rect 1478 535 1484 536
rect 1478 531 1479 535
rect 1483 531 1484 535
rect 1478 530 1484 531
rect 1526 535 1532 536
rect 1526 531 1527 535
rect 1531 531 1532 535
rect 1526 530 1532 531
rect 1574 535 1580 536
rect 1574 531 1575 535
rect 1579 531 1580 535
rect 1574 530 1580 531
rect 1622 535 1628 536
rect 1622 531 1623 535
rect 1627 531 1628 535
rect 1622 530 1628 531
rect 1654 535 1660 536
rect 1654 531 1655 535
rect 1659 531 1660 535
rect 1654 530 1660 531
rect 1694 533 1700 534
rect 1694 529 1695 533
rect 1699 529 1700 533
rect 1694 528 1700 529
rect 1286 527 1292 528
rect 134 518 140 519
rect 1422 518 1428 519
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 134 514 135 518
rect 139 514 140 518
rect 134 513 140 514
rect 506 517 512 518
rect 506 513 507 517
rect 511 513 512 517
rect 506 512 512 513
rect 1258 517 1264 518
rect 1258 513 1259 517
rect 1263 513 1264 517
rect 1422 514 1423 518
rect 1427 514 1428 518
rect 1422 513 1428 514
rect 1478 518 1484 519
rect 1478 514 1479 518
rect 1483 514 1484 518
rect 1478 513 1484 514
rect 1526 518 1532 519
rect 1526 514 1527 518
rect 1531 514 1532 518
rect 1526 513 1532 514
rect 1574 518 1580 519
rect 1574 514 1575 518
rect 1579 514 1580 518
rect 1574 513 1580 514
rect 1622 518 1628 519
rect 1622 514 1623 518
rect 1627 514 1628 518
rect 1622 513 1628 514
rect 1654 518 1660 519
rect 1654 514 1655 518
rect 1659 514 1660 518
rect 1654 513 1660 514
rect 1694 516 1700 517
rect 1258 512 1264 513
rect 1694 512 1695 516
rect 1699 512 1700 516
rect 110 511 116 512
rect 1694 511 1700 512
rect 174 498 180 499
rect 398 498 404 499
rect 174 494 175 498
rect 179 494 180 498
rect 302 497 308 498
rect 174 493 180 494
rect 246 493 252 494
rect 246 489 247 493
rect 251 489 252 493
rect 302 493 303 497
rect 307 493 308 497
rect 398 494 399 498
rect 403 494 404 498
rect 654 498 660 499
rect 654 494 655 498
rect 659 494 660 498
rect 782 498 788 499
rect 782 494 783 498
rect 787 494 788 498
rect 934 498 940 499
rect 934 494 935 498
rect 939 494 940 498
rect 1102 498 1108 499
rect 1102 494 1103 498
rect 1107 494 1108 498
rect 398 493 404 494
rect 470 493 476 494
rect 654 493 660 494
rect 726 493 732 494
rect 782 493 788 494
rect 870 493 876 494
rect 934 493 940 494
rect 1030 493 1036 494
rect 1102 493 1108 494
rect 1198 493 1204 494
rect 302 492 308 493
rect 246 488 252 489
rect 470 489 471 493
rect 475 489 476 493
rect 470 488 476 489
rect 726 489 727 493
rect 731 489 732 493
rect 726 488 732 489
rect 870 489 871 493
rect 875 489 876 493
rect 870 488 876 489
rect 1030 489 1031 493
rect 1035 489 1036 493
rect 1030 488 1036 489
rect 1198 489 1199 493
rect 1203 489 1204 493
rect 1198 488 1204 489
rect 374 399 380 400
rect 374 395 375 399
rect 379 395 380 399
rect 614 399 620 400
rect 614 395 615 399
rect 619 395 620 399
rect 302 394 308 395
rect 374 394 380 395
rect 542 394 548 395
rect 614 394 620 395
rect 670 395 676 396
rect 1230 395 1236 396
rect 302 390 303 394
rect 307 390 308 394
rect 302 389 308 390
rect 542 390 543 394
rect 547 390 548 394
rect 670 391 671 395
rect 675 391 676 395
rect 670 390 676 391
rect 950 394 956 395
rect 950 390 951 394
rect 955 390 956 394
rect 1230 391 1231 395
rect 1235 391 1236 395
rect 1230 390 1236 391
rect 542 389 548 390
rect 950 389 956 390
rect 1358 389 1364 390
rect 1358 385 1359 389
rect 1363 385 1364 389
rect 1358 384 1364 385
rect 1438 379 1444 380
rect 486 377 492 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 110 371 116 372
rect 134 374 140 375
rect 134 370 135 374
rect 139 370 140 374
rect 134 369 140 370
rect 166 374 172 375
rect 166 370 167 374
rect 171 370 172 374
rect 166 369 172 370
rect 198 374 204 375
rect 198 370 199 374
rect 203 370 204 374
rect 198 369 204 370
rect 230 374 236 375
rect 230 370 231 374
rect 235 370 236 374
rect 230 369 236 370
rect 262 374 268 375
rect 262 370 263 374
rect 267 370 268 374
rect 262 369 268 370
rect 414 374 420 375
rect 414 370 415 374
rect 419 370 420 374
rect 414 369 420 370
rect 446 374 452 375
rect 446 370 447 374
rect 451 370 452 374
rect 486 373 487 377
rect 491 373 492 377
rect 1030 377 1036 378
rect 486 372 492 373
rect 754 375 760 376
rect 754 371 755 375
rect 759 371 760 375
rect 754 370 760 371
rect 902 374 908 375
rect 902 370 903 374
rect 907 370 908 374
rect 1030 373 1031 377
rect 1035 373 1036 377
rect 1030 372 1036 373
rect 1074 375 1080 376
rect 1438 375 1439 379
rect 1443 375 1444 379
rect 1694 376 1700 377
rect 1074 371 1075 375
rect 1079 371 1080 375
rect 1074 370 1080 371
rect 1318 374 1324 375
rect 1438 374 1444 375
rect 1478 374 1484 375
rect 1318 370 1319 374
rect 1323 370 1324 374
rect 446 369 452 370
rect 902 369 908 370
rect 1318 369 1324 370
rect 1478 370 1479 374
rect 1483 370 1484 374
rect 1478 369 1484 370
rect 1518 374 1524 375
rect 1518 370 1519 374
rect 1523 370 1524 374
rect 1518 369 1524 370
rect 1558 374 1564 375
rect 1558 370 1559 374
rect 1563 370 1564 374
rect 1558 369 1564 370
rect 1590 374 1596 375
rect 1590 370 1591 374
rect 1595 370 1596 374
rect 1590 369 1596 370
rect 1622 374 1628 375
rect 1622 370 1623 374
rect 1627 370 1628 374
rect 1622 369 1628 370
rect 1654 374 1660 375
rect 1654 370 1655 374
rect 1659 370 1660 374
rect 1694 372 1695 376
rect 1699 372 1700 376
rect 1694 371 1700 372
rect 1654 369 1660 370
rect 782 360 788 361
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 134 357 140 358
rect 134 353 135 357
rect 139 353 140 357
rect 134 352 140 353
rect 166 357 172 358
rect 166 353 167 357
rect 171 353 172 357
rect 166 352 172 353
rect 198 357 204 358
rect 198 353 199 357
rect 203 353 204 357
rect 198 352 204 353
rect 230 357 236 358
rect 230 353 231 357
rect 235 353 236 357
rect 230 352 236 353
rect 262 357 268 358
rect 414 357 420 358
rect 262 353 263 357
rect 267 353 268 357
rect 262 352 268 353
rect 294 356 300 357
rect 294 352 295 356
rect 299 352 300 356
rect 414 353 415 357
rect 419 353 420 357
rect 294 351 300 352
rect 374 352 380 353
rect 414 352 420 353
rect 446 357 452 358
rect 446 353 447 357
rect 451 353 452 357
rect 446 352 452 353
rect 534 356 540 357
rect 534 352 535 356
rect 539 352 540 356
rect 782 356 783 360
rect 787 356 788 360
rect 1102 360 1108 361
rect 782 355 788 356
rect 902 357 908 358
rect 670 354 676 355
rect 374 348 375 352
rect 379 348 380 352
rect 534 351 540 352
rect 614 352 620 353
rect 374 347 380 348
rect 502 350 508 351
rect 502 346 503 350
rect 507 346 508 350
rect 614 348 615 352
rect 619 348 620 352
rect 670 350 671 354
rect 675 350 676 354
rect 902 353 903 357
rect 907 353 908 357
rect 902 352 908 353
rect 942 356 948 357
rect 942 352 943 356
rect 947 352 948 356
rect 1102 356 1103 360
rect 1107 356 1108 360
rect 1694 359 1700 360
rect 1102 355 1108 356
rect 1318 357 1324 358
rect 1478 357 1484 358
rect 942 351 948 352
rect 1230 354 1236 355
rect 670 349 676 350
rect 1046 350 1052 351
rect 614 347 620 348
rect 502 345 508 346
rect 1046 346 1047 350
rect 1051 346 1052 350
rect 1230 350 1231 354
rect 1235 350 1236 354
rect 1318 353 1319 357
rect 1323 353 1324 357
rect 1318 352 1324 353
rect 1438 356 1444 357
rect 1438 352 1439 356
rect 1443 352 1444 356
rect 1478 353 1479 357
rect 1483 353 1484 357
rect 1478 352 1484 353
rect 1518 357 1524 358
rect 1518 353 1519 357
rect 1523 353 1524 357
rect 1518 352 1524 353
rect 1558 357 1564 358
rect 1558 353 1559 357
rect 1563 353 1564 357
rect 1558 352 1564 353
rect 1590 357 1596 358
rect 1590 353 1591 357
rect 1595 353 1596 357
rect 1590 352 1596 353
rect 1622 357 1628 358
rect 1622 353 1623 357
rect 1627 353 1628 357
rect 1622 352 1628 353
rect 1654 357 1660 358
rect 1654 353 1655 357
rect 1659 353 1660 357
rect 1694 355 1695 359
rect 1699 355 1700 359
rect 1694 354 1700 355
rect 1654 352 1660 353
rect 1438 351 1444 352
rect 1230 349 1236 350
rect 1350 349 1356 350
rect 1046 345 1052 346
rect 1350 345 1351 349
rect 1355 345 1356 349
rect 1350 344 1356 345
rect 1198 311 1204 312
rect 1198 307 1199 311
rect 1203 307 1204 311
rect 598 306 604 307
rect 134 303 140 304
rect 110 301 116 302
rect 110 297 111 301
rect 115 297 116 301
rect 134 299 135 303
rect 139 299 140 303
rect 134 298 140 299
rect 166 303 172 304
rect 166 299 167 303
rect 171 299 172 303
rect 166 298 172 299
rect 198 303 204 304
rect 198 299 199 303
rect 203 299 204 303
rect 198 298 204 299
rect 230 303 236 304
rect 230 299 231 303
rect 235 299 236 303
rect 230 298 236 299
rect 262 303 268 304
rect 262 299 263 303
rect 267 299 268 303
rect 262 298 268 299
rect 294 303 300 304
rect 294 299 295 303
rect 299 299 300 303
rect 294 298 300 299
rect 326 303 332 304
rect 326 299 327 303
rect 331 299 332 303
rect 326 298 332 299
rect 358 303 364 304
rect 358 299 359 303
rect 363 299 364 303
rect 358 298 364 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 422 303 428 304
rect 422 299 423 303
rect 427 299 428 303
rect 422 298 428 299
rect 454 303 460 304
rect 454 299 455 303
rect 459 299 460 303
rect 454 298 460 299
rect 486 303 492 304
rect 486 299 487 303
rect 491 299 492 303
rect 486 298 492 299
rect 518 303 524 304
rect 518 299 519 303
rect 523 299 524 303
rect 518 298 524 299
rect 550 303 556 304
rect 550 299 551 303
rect 555 299 556 303
rect 598 302 599 306
rect 603 302 604 306
rect 598 301 604 302
rect 702 306 708 307
rect 702 302 703 306
rect 707 302 708 306
rect 702 301 708 302
rect 806 306 812 307
rect 806 302 807 306
rect 811 302 812 306
rect 806 301 812 302
rect 910 306 916 307
rect 910 302 911 306
rect 915 302 916 306
rect 1110 306 1116 307
rect 1198 306 1204 307
rect 910 301 916 302
rect 998 303 1004 304
rect 550 298 556 299
rect 998 299 999 303
rect 1003 299 1004 303
rect 998 298 1004 299
rect 1030 303 1036 304
rect 1030 299 1031 303
rect 1035 299 1036 303
rect 1030 298 1036 299
rect 1062 303 1068 304
rect 1062 299 1063 303
rect 1067 299 1068 303
rect 1110 302 1111 306
rect 1115 302 1116 306
rect 1110 301 1116 302
rect 1286 304 1292 305
rect 1286 300 1287 304
rect 1291 300 1292 304
rect 1286 299 1292 300
rect 1318 303 1324 304
rect 1318 299 1319 303
rect 1323 299 1324 303
rect 1062 298 1068 299
rect 1318 298 1324 299
rect 1350 303 1356 304
rect 1350 299 1351 303
rect 1355 299 1356 303
rect 1350 298 1356 299
rect 1382 303 1388 304
rect 1382 299 1383 303
rect 1387 299 1388 303
rect 1382 298 1388 299
rect 1414 303 1420 304
rect 1414 299 1415 303
rect 1419 299 1420 303
rect 1414 298 1420 299
rect 1446 303 1452 304
rect 1446 299 1447 303
rect 1451 299 1452 303
rect 1446 298 1452 299
rect 1478 303 1484 304
rect 1478 299 1479 303
rect 1483 299 1484 303
rect 1478 298 1484 299
rect 1518 303 1524 304
rect 1518 299 1519 303
rect 1523 299 1524 303
rect 1518 298 1524 299
rect 1558 303 1564 304
rect 1558 299 1559 303
rect 1563 299 1564 303
rect 1558 298 1564 299
rect 1590 303 1596 304
rect 1590 299 1591 303
rect 1595 299 1596 303
rect 1590 298 1596 299
rect 1622 303 1628 304
rect 1622 299 1623 303
rect 1627 299 1628 303
rect 1622 298 1628 299
rect 1654 303 1660 304
rect 1654 299 1655 303
rect 1659 299 1660 303
rect 1654 298 1660 299
rect 1694 301 1700 302
rect 110 296 116 297
rect 1694 297 1695 301
rect 1699 297 1700 301
rect 1694 296 1700 297
rect 134 286 140 287
rect 110 284 116 285
rect 110 280 111 284
rect 115 280 116 284
rect 134 282 135 286
rect 139 282 140 286
rect 134 281 140 282
rect 166 286 172 287
rect 166 282 167 286
rect 171 282 172 286
rect 166 281 172 282
rect 198 286 204 287
rect 198 282 199 286
rect 203 282 204 286
rect 198 281 204 282
rect 230 286 236 287
rect 230 282 231 286
rect 235 282 236 286
rect 230 281 236 282
rect 262 286 268 287
rect 262 282 263 286
rect 267 282 268 286
rect 262 281 268 282
rect 294 286 300 287
rect 294 282 295 286
rect 299 282 300 286
rect 294 281 300 282
rect 326 286 332 287
rect 326 282 327 286
rect 331 282 332 286
rect 326 281 332 282
rect 358 286 364 287
rect 358 282 359 286
rect 363 282 364 286
rect 358 281 364 282
rect 390 286 396 287
rect 390 282 391 286
rect 395 282 396 286
rect 390 281 396 282
rect 422 286 428 287
rect 422 282 423 286
rect 427 282 428 286
rect 422 281 428 282
rect 454 286 460 287
rect 454 282 455 286
rect 459 282 460 286
rect 454 281 460 282
rect 486 286 492 287
rect 486 282 487 286
rect 491 282 492 286
rect 486 281 492 282
rect 518 286 524 287
rect 518 282 519 286
rect 523 282 524 286
rect 518 281 524 282
rect 550 286 556 287
rect 550 282 551 286
rect 555 282 556 286
rect 550 281 556 282
rect 998 286 1004 287
rect 998 282 999 286
rect 1003 282 1004 286
rect 998 281 1004 282
rect 1030 286 1036 287
rect 1030 282 1031 286
rect 1035 282 1036 286
rect 1030 281 1036 282
rect 1062 286 1068 287
rect 1062 282 1063 286
rect 1067 282 1068 286
rect 1318 286 1324 287
rect 1318 282 1319 286
rect 1323 282 1324 286
rect 1062 281 1068 282
rect 1286 281 1292 282
rect 1318 281 1324 282
rect 1350 286 1356 287
rect 1350 282 1351 286
rect 1355 282 1356 286
rect 1350 281 1356 282
rect 1382 286 1388 287
rect 1382 282 1383 286
rect 1387 282 1388 286
rect 1382 281 1388 282
rect 1414 286 1420 287
rect 1414 282 1415 286
rect 1419 282 1420 286
rect 1414 281 1420 282
rect 1446 286 1452 287
rect 1446 282 1447 286
rect 1451 282 1452 286
rect 1446 281 1452 282
rect 1478 286 1484 287
rect 1478 282 1479 286
rect 1483 282 1484 286
rect 1478 281 1484 282
rect 1518 286 1524 287
rect 1518 282 1519 286
rect 1523 282 1524 286
rect 1518 281 1524 282
rect 1558 286 1564 287
rect 1558 282 1559 286
rect 1563 282 1564 286
rect 1558 281 1564 282
rect 1590 286 1596 287
rect 1590 282 1591 286
rect 1595 282 1596 286
rect 1590 281 1596 282
rect 1622 286 1628 287
rect 1622 282 1623 286
rect 1627 282 1628 286
rect 1622 281 1628 282
rect 1654 286 1660 287
rect 1654 282 1655 286
rect 1659 282 1660 286
rect 1654 281 1660 282
rect 1694 284 1700 285
rect 110 279 116 280
rect 1286 277 1287 281
rect 1291 277 1292 281
rect 1694 280 1695 284
rect 1699 280 1700 284
rect 1694 279 1700 280
rect 1286 276 1292 277
rect 1206 271 1212 272
rect 1206 267 1207 271
rect 1211 267 1212 271
rect 1206 266 1212 267
rect 598 265 604 266
rect 598 261 599 265
rect 603 261 604 265
rect 598 260 604 261
rect 702 265 708 266
rect 702 261 703 265
rect 707 261 708 265
rect 702 260 708 261
rect 806 265 812 266
rect 806 261 807 265
rect 811 261 812 265
rect 806 260 812 261
rect 910 265 916 266
rect 910 261 911 265
rect 915 261 916 265
rect 910 260 916 261
rect 1110 265 1116 266
rect 1110 261 1111 265
rect 1115 261 1116 265
rect 1110 260 1116 261
rect 694 235 700 236
rect 694 231 695 235
rect 699 231 700 235
rect 694 230 700 231
rect 966 235 972 236
rect 966 231 967 235
rect 971 231 972 235
rect 966 230 972 231
rect 838 229 844 230
rect 838 225 839 229
rect 843 225 844 229
rect 838 224 844 225
rect 918 219 924 220
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 918 215 919 219
rect 923 215 924 219
rect 1694 216 1700 217
rect 110 211 116 212
rect 182 214 188 215
rect 182 210 183 214
rect 187 210 188 214
rect 182 209 188 210
rect 214 214 220 215
rect 214 210 215 214
rect 219 210 220 214
rect 214 209 220 210
rect 246 214 252 215
rect 246 210 247 214
rect 251 210 252 214
rect 246 209 252 210
rect 278 214 284 215
rect 278 210 279 214
rect 283 210 284 214
rect 278 209 284 210
rect 310 214 316 215
rect 310 210 311 214
rect 315 210 316 214
rect 310 209 316 210
rect 342 214 348 215
rect 342 210 343 214
rect 347 210 348 214
rect 342 209 348 210
rect 374 214 380 215
rect 374 210 375 214
rect 379 210 380 214
rect 374 209 380 210
rect 406 214 412 215
rect 406 210 407 214
rect 411 210 412 214
rect 406 209 412 210
rect 438 214 444 215
rect 438 210 439 214
rect 443 210 444 214
rect 438 209 444 210
rect 470 214 476 215
rect 470 210 471 214
rect 475 210 476 214
rect 470 209 476 210
rect 502 214 508 215
rect 502 210 503 214
rect 507 210 508 214
rect 502 209 508 210
rect 534 214 540 215
rect 534 210 535 214
rect 539 210 540 214
rect 534 209 540 210
rect 566 214 572 215
rect 566 210 567 214
rect 571 210 572 214
rect 566 209 572 210
rect 598 214 604 215
rect 598 210 599 214
rect 603 210 604 214
rect 598 209 604 210
rect 638 214 644 215
rect 638 210 639 214
rect 643 210 644 214
rect 638 209 644 210
rect 790 214 796 215
rect 918 214 924 215
rect 1062 214 1068 215
rect 790 210 791 214
rect 795 210 796 214
rect 790 209 796 210
rect 1062 210 1063 214
rect 1067 210 1068 214
rect 1062 209 1068 210
rect 1102 214 1108 215
rect 1102 210 1103 214
rect 1107 210 1108 214
rect 1102 209 1108 210
rect 1142 214 1148 215
rect 1142 210 1143 214
rect 1147 210 1148 214
rect 1142 209 1148 210
rect 1182 214 1188 215
rect 1182 210 1183 214
rect 1187 210 1188 214
rect 1182 209 1188 210
rect 1222 214 1228 215
rect 1222 210 1223 214
rect 1227 210 1228 214
rect 1222 209 1228 210
rect 1262 214 1268 215
rect 1262 210 1263 214
rect 1267 210 1268 214
rect 1262 209 1268 210
rect 1302 214 1308 215
rect 1302 210 1303 214
rect 1307 210 1308 214
rect 1302 209 1308 210
rect 1342 214 1348 215
rect 1342 210 1343 214
rect 1347 210 1348 214
rect 1342 209 1348 210
rect 1374 214 1380 215
rect 1374 210 1375 214
rect 1379 210 1380 214
rect 1374 209 1380 210
rect 1406 214 1412 215
rect 1406 210 1407 214
rect 1411 210 1412 214
rect 1406 209 1412 210
rect 1438 214 1444 215
rect 1438 210 1439 214
rect 1443 210 1444 214
rect 1438 209 1444 210
rect 1478 214 1484 215
rect 1478 210 1479 214
rect 1483 210 1484 214
rect 1478 209 1484 210
rect 1518 214 1524 215
rect 1518 210 1519 214
rect 1523 210 1524 214
rect 1518 209 1524 210
rect 1558 214 1564 215
rect 1558 210 1559 214
rect 1563 210 1564 214
rect 1558 209 1564 210
rect 1590 214 1596 215
rect 1590 210 1591 214
rect 1595 210 1596 214
rect 1590 209 1596 210
rect 1622 214 1628 215
rect 1622 210 1623 214
rect 1627 210 1628 214
rect 1622 209 1628 210
rect 1654 214 1660 215
rect 1654 210 1655 214
rect 1659 210 1660 214
rect 1694 212 1695 216
rect 1699 212 1700 216
rect 1694 211 1700 212
rect 1654 209 1660 210
rect 110 199 116 200
rect 110 195 111 199
rect 115 195 116 199
rect 1694 199 1700 200
rect 110 194 116 195
rect 182 197 188 198
rect 182 193 183 197
rect 187 193 188 197
rect 182 192 188 193
rect 214 197 220 198
rect 214 193 215 197
rect 219 193 220 197
rect 214 192 220 193
rect 246 197 252 198
rect 246 193 247 197
rect 251 193 252 197
rect 246 192 252 193
rect 278 197 284 198
rect 278 193 279 197
rect 283 193 284 197
rect 278 192 284 193
rect 310 197 316 198
rect 310 193 311 197
rect 315 193 316 197
rect 310 192 316 193
rect 342 197 348 198
rect 342 193 343 197
rect 347 193 348 197
rect 342 192 348 193
rect 374 197 380 198
rect 374 193 375 197
rect 379 193 380 197
rect 374 192 380 193
rect 406 197 412 198
rect 406 193 407 197
rect 411 193 412 197
rect 406 192 412 193
rect 438 197 444 198
rect 438 193 439 197
rect 443 193 444 197
rect 438 192 444 193
rect 470 197 476 198
rect 470 193 471 197
rect 475 193 476 197
rect 470 192 476 193
rect 502 197 508 198
rect 502 193 503 197
rect 507 193 508 197
rect 502 192 508 193
rect 534 197 540 198
rect 534 193 535 197
rect 539 193 540 197
rect 534 192 540 193
rect 566 197 572 198
rect 566 193 567 197
rect 571 193 572 197
rect 566 192 572 193
rect 598 197 604 198
rect 598 193 599 197
rect 603 193 604 197
rect 598 192 604 193
rect 638 197 644 198
rect 638 193 639 197
rect 643 193 644 197
rect 790 197 796 198
rect 1062 197 1068 198
rect 638 192 644 193
rect 694 194 700 195
rect 694 190 695 194
rect 699 190 700 194
rect 790 193 791 197
rect 795 193 796 197
rect 790 192 796 193
rect 918 196 924 197
rect 918 192 919 196
rect 923 192 924 196
rect 918 191 924 192
rect 966 194 972 195
rect 966 190 967 194
rect 971 190 972 194
rect 1062 193 1063 197
rect 1067 193 1068 197
rect 1062 192 1068 193
rect 1102 197 1108 198
rect 1102 193 1103 197
rect 1107 193 1108 197
rect 1102 192 1108 193
rect 1142 197 1148 198
rect 1142 193 1143 197
rect 1147 193 1148 197
rect 1142 192 1148 193
rect 1182 197 1188 198
rect 1182 193 1183 197
rect 1187 193 1188 197
rect 1182 192 1188 193
rect 1222 197 1228 198
rect 1222 193 1223 197
rect 1227 193 1228 197
rect 1222 192 1228 193
rect 1262 197 1268 198
rect 1262 193 1263 197
rect 1267 193 1268 197
rect 1262 192 1268 193
rect 1302 197 1308 198
rect 1302 193 1303 197
rect 1307 193 1308 197
rect 1302 192 1308 193
rect 1342 197 1348 198
rect 1342 193 1343 197
rect 1347 193 1348 197
rect 1342 192 1348 193
rect 1374 197 1380 198
rect 1374 193 1375 197
rect 1379 193 1380 197
rect 1374 192 1380 193
rect 1406 197 1412 198
rect 1406 193 1407 197
rect 1411 193 1412 197
rect 1406 192 1412 193
rect 1438 197 1444 198
rect 1438 193 1439 197
rect 1443 193 1444 197
rect 1438 192 1444 193
rect 1478 197 1484 198
rect 1478 193 1479 197
rect 1483 193 1484 197
rect 1478 192 1484 193
rect 1518 197 1524 198
rect 1518 193 1519 197
rect 1523 193 1524 197
rect 1518 192 1524 193
rect 1558 197 1564 198
rect 1558 193 1559 197
rect 1563 193 1564 197
rect 1558 192 1564 193
rect 1590 197 1596 198
rect 1590 193 1591 197
rect 1595 193 1596 197
rect 1590 192 1596 193
rect 1622 197 1628 198
rect 1622 193 1623 197
rect 1627 193 1628 197
rect 1622 192 1628 193
rect 1654 197 1660 198
rect 1654 193 1655 197
rect 1659 193 1660 197
rect 1694 195 1695 199
rect 1699 195 1700 199
rect 1694 194 1700 195
rect 1654 192 1660 193
rect 694 189 700 190
rect 830 189 836 190
rect 966 189 972 190
rect 830 185 831 189
rect 835 185 836 189
rect 830 184 836 185
rect 134 167 140 168
rect 110 165 116 166
rect 110 161 111 165
rect 115 161 116 165
rect 134 163 135 167
rect 139 163 140 167
rect 134 162 140 163
rect 166 167 172 168
rect 166 163 167 167
rect 171 163 172 167
rect 166 162 172 163
rect 214 167 220 168
rect 214 163 215 167
rect 219 163 220 167
rect 214 162 220 163
rect 262 167 268 168
rect 262 163 263 167
rect 267 163 268 167
rect 262 162 268 163
rect 310 167 316 168
rect 310 163 311 167
rect 315 163 316 167
rect 310 162 316 163
rect 366 167 372 168
rect 366 163 367 167
rect 371 163 372 167
rect 366 162 372 163
rect 414 167 420 168
rect 414 163 415 167
rect 419 163 420 167
rect 414 162 420 163
rect 470 167 476 168
rect 470 163 471 167
rect 475 163 476 167
rect 470 162 476 163
rect 534 167 540 168
rect 534 163 535 167
rect 539 163 540 167
rect 534 162 540 163
rect 606 167 612 168
rect 606 163 607 167
rect 611 163 612 167
rect 606 162 612 163
rect 686 167 692 168
rect 686 163 687 167
rect 691 163 692 167
rect 686 162 692 163
rect 774 167 780 168
rect 774 163 775 167
rect 779 163 780 167
rect 774 162 780 163
rect 862 167 868 168
rect 862 163 863 167
rect 867 163 868 167
rect 862 162 868 163
rect 958 167 964 168
rect 958 163 959 167
rect 963 163 964 167
rect 958 162 964 163
rect 1054 167 1060 168
rect 1054 163 1055 167
rect 1059 163 1060 167
rect 1054 162 1060 163
rect 1150 167 1156 168
rect 1150 163 1151 167
rect 1155 163 1156 167
rect 1150 162 1156 163
rect 1238 167 1244 168
rect 1238 163 1239 167
rect 1243 163 1244 167
rect 1238 162 1244 163
rect 1326 167 1332 168
rect 1326 163 1327 167
rect 1331 163 1332 167
rect 1326 162 1332 163
rect 1414 167 1420 168
rect 1414 163 1415 167
rect 1419 163 1420 167
rect 1414 162 1420 163
rect 1502 167 1508 168
rect 1502 163 1503 167
rect 1507 163 1508 167
rect 1502 162 1508 163
rect 1590 167 1596 168
rect 1590 163 1591 167
rect 1595 163 1596 167
rect 1590 162 1596 163
rect 1654 167 1660 168
rect 1654 163 1655 167
rect 1659 163 1660 167
rect 1654 162 1660 163
rect 1694 165 1700 166
rect 110 160 116 161
rect 1694 161 1695 165
rect 1699 161 1700 165
rect 1694 160 1700 161
rect 134 150 140 151
rect 110 148 116 149
rect 110 144 111 148
rect 115 144 116 148
rect 134 146 135 150
rect 139 146 140 150
rect 134 145 140 146
rect 166 150 172 151
rect 166 146 167 150
rect 171 146 172 150
rect 166 145 172 146
rect 214 150 220 151
rect 214 146 215 150
rect 219 146 220 150
rect 214 145 220 146
rect 262 150 268 151
rect 262 146 263 150
rect 267 146 268 150
rect 262 145 268 146
rect 310 150 316 151
rect 310 146 311 150
rect 315 146 316 150
rect 310 145 316 146
rect 366 150 372 151
rect 366 146 367 150
rect 371 146 372 150
rect 366 145 372 146
rect 414 150 420 151
rect 414 146 415 150
rect 419 146 420 150
rect 414 145 420 146
rect 470 150 476 151
rect 470 146 471 150
rect 475 146 476 150
rect 470 145 476 146
rect 534 150 540 151
rect 534 146 535 150
rect 539 146 540 150
rect 534 145 540 146
rect 606 150 612 151
rect 606 146 607 150
rect 611 146 612 150
rect 606 145 612 146
rect 686 150 692 151
rect 686 146 687 150
rect 691 146 692 150
rect 686 145 692 146
rect 774 150 780 151
rect 774 146 775 150
rect 779 146 780 150
rect 774 145 780 146
rect 862 150 868 151
rect 862 146 863 150
rect 867 146 868 150
rect 862 145 868 146
rect 958 150 964 151
rect 958 146 959 150
rect 963 146 964 150
rect 958 145 964 146
rect 1054 150 1060 151
rect 1054 146 1055 150
rect 1059 146 1060 150
rect 1054 145 1060 146
rect 1150 150 1156 151
rect 1150 146 1151 150
rect 1155 146 1156 150
rect 1150 145 1156 146
rect 1238 150 1244 151
rect 1238 146 1239 150
rect 1243 146 1244 150
rect 1238 145 1244 146
rect 1326 150 1332 151
rect 1326 146 1327 150
rect 1331 146 1332 150
rect 1326 145 1332 146
rect 1414 150 1420 151
rect 1414 146 1415 150
rect 1419 146 1420 150
rect 1414 145 1420 146
rect 1502 150 1508 151
rect 1502 146 1503 150
rect 1507 146 1508 150
rect 1502 145 1508 146
rect 1590 150 1596 151
rect 1590 146 1591 150
rect 1595 146 1596 150
rect 1590 145 1596 146
rect 1654 150 1660 151
rect 1654 146 1655 150
rect 1659 146 1660 150
rect 1654 145 1660 146
rect 1694 148 1700 149
rect 110 143 116 144
rect 1694 144 1695 148
rect 1699 144 1700 148
rect 1694 143 1700 144
rect 110 108 116 109
rect 110 104 111 108
rect 115 104 116 108
rect 1694 108 1700 109
rect 110 103 116 104
rect 134 106 140 107
rect 134 102 135 106
rect 139 102 140 106
rect 134 101 140 102
rect 166 106 172 107
rect 166 102 167 106
rect 171 102 172 106
rect 166 101 172 102
rect 198 106 204 107
rect 198 102 199 106
rect 203 102 204 106
rect 198 101 204 102
rect 230 106 236 107
rect 230 102 231 106
rect 235 102 236 106
rect 230 101 236 102
rect 262 106 268 107
rect 262 102 263 106
rect 267 102 268 106
rect 262 101 268 102
rect 294 106 300 107
rect 294 102 295 106
rect 299 102 300 106
rect 294 101 300 102
rect 326 106 332 107
rect 326 102 327 106
rect 331 102 332 106
rect 326 101 332 102
rect 358 106 364 107
rect 358 102 359 106
rect 363 102 364 106
rect 358 101 364 102
rect 390 106 396 107
rect 390 102 391 106
rect 395 102 396 106
rect 390 101 396 102
rect 422 106 428 107
rect 422 102 423 106
rect 427 102 428 106
rect 422 101 428 102
rect 454 106 460 107
rect 454 102 455 106
rect 459 102 460 106
rect 454 101 460 102
rect 486 106 492 107
rect 486 102 487 106
rect 491 102 492 106
rect 486 101 492 102
rect 518 106 524 107
rect 518 102 519 106
rect 523 102 524 106
rect 518 101 524 102
rect 550 106 556 107
rect 550 102 551 106
rect 555 102 556 106
rect 550 101 556 102
rect 606 106 612 107
rect 606 102 607 106
rect 611 102 612 106
rect 606 101 612 102
rect 670 106 676 107
rect 670 102 671 106
rect 675 102 676 106
rect 670 101 676 102
rect 742 106 748 107
rect 742 102 743 106
rect 747 102 748 106
rect 742 101 748 102
rect 822 106 828 107
rect 822 102 823 106
rect 827 102 828 106
rect 822 101 828 102
rect 902 106 908 107
rect 902 102 903 106
rect 907 102 908 106
rect 902 101 908 102
rect 982 106 988 107
rect 982 102 983 106
rect 987 102 988 106
rect 982 101 988 102
rect 1054 106 1060 107
rect 1054 102 1055 106
rect 1059 102 1060 106
rect 1054 101 1060 102
rect 1118 106 1124 107
rect 1118 102 1119 106
rect 1123 102 1124 106
rect 1118 101 1124 102
rect 1174 106 1180 107
rect 1174 102 1175 106
rect 1179 102 1180 106
rect 1174 101 1180 102
rect 1222 106 1228 107
rect 1222 102 1223 106
rect 1227 102 1228 106
rect 1222 101 1228 102
rect 1270 106 1276 107
rect 1270 102 1271 106
rect 1275 102 1276 106
rect 1270 101 1276 102
rect 1310 106 1316 107
rect 1310 102 1311 106
rect 1315 102 1316 106
rect 1310 101 1316 102
rect 1342 106 1348 107
rect 1342 102 1343 106
rect 1347 102 1348 106
rect 1342 101 1348 102
rect 1374 106 1380 107
rect 1374 102 1375 106
rect 1379 102 1380 106
rect 1374 101 1380 102
rect 1406 106 1412 107
rect 1406 102 1407 106
rect 1411 102 1412 106
rect 1406 101 1412 102
rect 1438 106 1444 107
rect 1438 102 1439 106
rect 1443 102 1444 106
rect 1438 101 1444 102
rect 1478 106 1484 107
rect 1478 102 1479 106
rect 1483 102 1484 106
rect 1478 101 1484 102
rect 1518 106 1524 107
rect 1518 102 1519 106
rect 1523 102 1524 106
rect 1518 101 1524 102
rect 1558 106 1564 107
rect 1558 102 1559 106
rect 1563 102 1564 106
rect 1558 101 1564 102
rect 1590 106 1596 107
rect 1590 102 1591 106
rect 1595 102 1596 106
rect 1590 101 1596 102
rect 1622 106 1628 107
rect 1622 102 1623 106
rect 1627 102 1628 106
rect 1622 101 1628 102
rect 1654 106 1660 107
rect 1654 102 1655 106
rect 1659 102 1660 106
rect 1694 104 1695 108
rect 1699 104 1700 108
rect 1694 103 1700 104
rect 1654 101 1660 102
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 1694 91 1700 92
rect 110 86 116 87
rect 134 89 140 90
rect 134 85 135 89
rect 139 85 140 89
rect 134 84 140 85
rect 166 89 172 90
rect 166 85 167 89
rect 171 85 172 89
rect 166 84 172 85
rect 198 89 204 90
rect 198 85 199 89
rect 203 85 204 89
rect 198 84 204 85
rect 230 89 236 90
rect 230 85 231 89
rect 235 85 236 89
rect 230 84 236 85
rect 262 89 268 90
rect 262 85 263 89
rect 267 85 268 89
rect 262 84 268 85
rect 294 89 300 90
rect 294 85 295 89
rect 299 85 300 89
rect 294 84 300 85
rect 326 89 332 90
rect 326 85 327 89
rect 331 85 332 89
rect 326 84 332 85
rect 358 89 364 90
rect 358 85 359 89
rect 363 85 364 89
rect 358 84 364 85
rect 390 89 396 90
rect 390 85 391 89
rect 395 85 396 89
rect 390 84 396 85
rect 422 89 428 90
rect 422 85 423 89
rect 427 85 428 89
rect 422 84 428 85
rect 454 89 460 90
rect 454 85 455 89
rect 459 85 460 89
rect 454 84 460 85
rect 486 89 492 90
rect 486 85 487 89
rect 491 85 492 89
rect 486 84 492 85
rect 518 89 524 90
rect 518 85 519 89
rect 523 85 524 89
rect 518 84 524 85
rect 550 89 556 90
rect 550 85 551 89
rect 555 85 556 89
rect 550 84 556 85
rect 606 89 612 90
rect 606 85 607 89
rect 611 85 612 89
rect 606 84 612 85
rect 670 89 676 90
rect 670 85 671 89
rect 675 85 676 89
rect 670 84 676 85
rect 742 89 748 90
rect 742 85 743 89
rect 747 85 748 89
rect 742 84 748 85
rect 822 89 828 90
rect 822 85 823 89
rect 827 85 828 89
rect 822 84 828 85
rect 902 89 908 90
rect 902 85 903 89
rect 907 85 908 89
rect 902 84 908 85
rect 982 89 988 90
rect 982 85 983 89
rect 987 85 988 89
rect 982 84 988 85
rect 1054 89 1060 90
rect 1054 85 1055 89
rect 1059 85 1060 89
rect 1054 84 1060 85
rect 1118 89 1124 90
rect 1118 85 1119 89
rect 1123 85 1124 89
rect 1118 84 1124 85
rect 1174 89 1180 90
rect 1174 85 1175 89
rect 1179 85 1180 89
rect 1174 84 1180 85
rect 1222 89 1228 90
rect 1222 85 1223 89
rect 1227 85 1228 89
rect 1222 84 1228 85
rect 1270 89 1276 90
rect 1270 85 1271 89
rect 1275 85 1276 89
rect 1270 84 1276 85
rect 1310 89 1316 90
rect 1310 85 1311 89
rect 1315 85 1316 89
rect 1310 84 1316 85
rect 1342 89 1348 90
rect 1342 85 1343 89
rect 1347 85 1348 89
rect 1342 84 1348 85
rect 1374 89 1380 90
rect 1374 85 1375 89
rect 1379 85 1380 89
rect 1374 84 1380 85
rect 1406 89 1412 90
rect 1406 85 1407 89
rect 1411 85 1412 89
rect 1406 84 1412 85
rect 1438 89 1444 90
rect 1438 85 1439 89
rect 1443 85 1444 89
rect 1438 84 1444 85
rect 1478 89 1484 90
rect 1478 85 1479 89
rect 1483 85 1484 89
rect 1478 84 1484 85
rect 1518 89 1524 90
rect 1518 85 1519 89
rect 1523 85 1524 89
rect 1518 84 1524 85
rect 1558 89 1564 90
rect 1558 85 1559 89
rect 1563 85 1564 89
rect 1558 84 1564 85
rect 1590 89 1596 90
rect 1590 85 1591 89
rect 1595 85 1596 89
rect 1590 84 1596 85
rect 1622 89 1628 90
rect 1622 85 1623 89
rect 1627 85 1628 89
rect 1622 84 1628 85
rect 1654 89 1660 90
rect 1654 85 1655 89
rect 1659 85 1660 89
rect 1694 87 1695 91
rect 1699 87 1700 91
rect 1694 86 1700 87
rect 1654 84 1660 85
<< m3c >>
rect 111 1749 115 1753
rect 151 1751 155 1755
rect 183 1751 187 1755
rect 215 1751 219 1755
rect 247 1751 251 1755
rect 279 1751 283 1755
rect 311 1751 315 1755
rect 343 1751 347 1755
rect 375 1751 379 1755
rect 407 1751 411 1755
rect 439 1751 443 1755
rect 471 1751 475 1755
rect 503 1751 507 1755
rect 535 1751 539 1755
rect 567 1751 571 1755
rect 599 1751 603 1755
rect 631 1751 635 1755
rect 663 1751 667 1755
rect 695 1751 699 1755
rect 727 1751 731 1755
rect 759 1751 763 1755
rect 791 1751 795 1755
rect 823 1751 827 1755
rect 855 1751 859 1755
rect 887 1751 891 1755
rect 919 1751 923 1755
rect 951 1751 955 1755
rect 983 1751 987 1755
rect 1695 1749 1699 1753
rect 111 1732 115 1736
rect 151 1734 155 1738
rect 183 1734 187 1738
rect 215 1734 219 1738
rect 247 1734 251 1738
rect 279 1734 283 1738
rect 311 1734 315 1738
rect 343 1734 347 1738
rect 375 1734 379 1738
rect 407 1734 411 1738
rect 439 1734 443 1738
rect 471 1734 475 1738
rect 503 1734 507 1738
rect 535 1734 539 1738
rect 567 1734 571 1738
rect 599 1734 603 1738
rect 631 1734 635 1738
rect 663 1734 667 1738
rect 695 1734 699 1738
rect 727 1734 731 1738
rect 759 1734 763 1738
rect 791 1734 795 1738
rect 823 1734 827 1738
rect 855 1734 859 1738
rect 887 1734 891 1738
rect 919 1734 923 1738
rect 951 1734 955 1738
rect 983 1734 987 1738
rect 1695 1732 1699 1736
rect 111 1700 115 1704
rect 191 1698 195 1702
rect 247 1698 251 1702
rect 319 1698 323 1702
rect 415 1698 419 1702
rect 527 1698 531 1702
rect 655 1698 659 1702
rect 791 1698 795 1702
rect 919 1698 923 1702
rect 1047 1698 1051 1702
rect 1159 1698 1163 1702
rect 1255 1698 1259 1702
rect 1335 1698 1339 1702
rect 1407 1698 1411 1702
rect 1463 1698 1467 1702
rect 1519 1698 1523 1702
rect 1567 1698 1571 1702
rect 1623 1698 1627 1702
rect 1655 1698 1659 1702
rect 1695 1700 1699 1704
rect 111 1683 115 1687
rect 191 1681 195 1685
rect 247 1681 251 1685
rect 319 1681 323 1685
rect 415 1681 419 1685
rect 527 1681 531 1685
rect 655 1681 659 1685
rect 791 1681 795 1685
rect 919 1681 923 1685
rect 1047 1681 1051 1685
rect 1159 1681 1163 1685
rect 1255 1681 1259 1685
rect 1335 1681 1339 1685
rect 1407 1681 1411 1685
rect 1463 1681 1467 1685
rect 1519 1681 1523 1685
rect 1567 1681 1571 1685
rect 1623 1681 1627 1685
rect 1655 1681 1659 1685
rect 1695 1683 1699 1687
rect 111 1657 115 1661
rect 135 1659 139 1663
rect 175 1659 179 1663
rect 263 1659 267 1663
rect 391 1659 395 1663
rect 543 1659 547 1663
rect 711 1659 715 1663
rect 879 1659 883 1663
rect 1039 1659 1043 1663
rect 1183 1659 1187 1663
rect 1319 1659 1323 1663
rect 1439 1659 1443 1663
rect 1559 1659 1563 1663
rect 1655 1659 1659 1663
rect 1695 1657 1699 1661
rect 111 1640 115 1644
rect 135 1642 139 1646
rect 175 1642 179 1646
rect 263 1642 267 1646
rect 391 1642 395 1646
rect 543 1642 547 1646
rect 711 1642 715 1646
rect 879 1642 883 1646
rect 1039 1642 1043 1646
rect 1183 1642 1187 1646
rect 1319 1642 1323 1646
rect 1439 1642 1443 1646
rect 1559 1642 1563 1646
rect 1655 1642 1659 1646
rect 1695 1640 1699 1644
rect 111 1604 115 1608
rect 135 1602 139 1606
rect 167 1602 171 1606
rect 199 1602 203 1606
rect 247 1602 251 1606
rect 327 1602 331 1606
rect 439 1602 443 1606
rect 567 1602 571 1606
rect 711 1602 715 1606
rect 855 1602 859 1606
rect 999 1602 1003 1606
rect 1127 1602 1131 1606
rect 1247 1602 1251 1606
rect 1359 1602 1363 1606
rect 1463 1602 1467 1606
rect 1567 1602 1571 1606
rect 1655 1602 1659 1606
rect 1695 1604 1699 1608
rect 111 1587 115 1591
rect 135 1585 139 1589
rect 167 1585 171 1589
rect 199 1585 203 1589
rect 247 1585 251 1589
rect 327 1585 331 1589
rect 439 1585 443 1589
rect 567 1585 571 1589
rect 711 1585 715 1589
rect 855 1585 859 1589
rect 999 1585 1003 1589
rect 1127 1585 1131 1589
rect 1247 1585 1251 1589
rect 1359 1585 1363 1589
rect 1463 1585 1467 1589
rect 1567 1585 1571 1589
rect 1655 1585 1659 1589
rect 1695 1587 1699 1591
rect 111 1569 115 1573
rect 135 1571 139 1575
rect 167 1571 171 1575
rect 231 1571 235 1575
rect 287 1571 291 1575
rect 343 1571 347 1575
rect 399 1571 403 1575
rect 455 1571 459 1575
rect 511 1571 515 1575
rect 575 1571 579 1575
rect 655 1571 659 1575
rect 751 1571 755 1575
rect 855 1571 859 1575
rect 959 1571 963 1575
rect 1063 1571 1067 1575
rect 1159 1571 1163 1575
rect 1247 1571 1251 1575
rect 1327 1571 1331 1575
rect 1399 1571 1403 1575
rect 1471 1571 1475 1575
rect 1535 1571 1539 1575
rect 1607 1571 1611 1575
rect 1655 1571 1659 1575
rect 1695 1569 1699 1573
rect 111 1552 115 1556
rect 135 1554 139 1558
rect 167 1554 171 1558
rect 231 1554 235 1558
rect 287 1554 291 1558
rect 343 1554 347 1558
rect 399 1554 403 1558
rect 455 1554 459 1558
rect 511 1554 515 1558
rect 575 1554 579 1558
rect 655 1554 659 1558
rect 751 1554 755 1558
rect 855 1554 859 1558
rect 959 1554 963 1558
rect 1063 1554 1067 1558
rect 1159 1554 1163 1558
rect 1247 1554 1251 1558
rect 1327 1554 1331 1558
rect 1399 1554 1403 1558
rect 1471 1554 1475 1558
rect 1535 1554 1539 1558
rect 1607 1554 1611 1558
rect 1655 1554 1659 1558
rect 1695 1552 1699 1556
rect 111 1524 115 1528
rect 135 1522 139 1526
rect 175 1522 179 1526
rect 223 1522 227 1526
rect 279 1522 283 1526
rect 335 1522 339 1526
rect 399 1522 403 1526
rect 463 1522 467 1526
rect 535 1522 539 1526
rect 607 1522 611 1526
rect 687 1522 691 1526
rect 775 1522 779 1526
rect 871 1522 875 1526
rect 975 1522 979 1526
rect 1079 1522 1083 1526
rect 1175 1522 1179 1526
rect 1271 1522 1275 1526
rect 1359 1522 1363 1526
rect 1439 1522 1443 1526
rect 1519 1522 1523 1526
rect 1599 1522 1603 1526
rect 1655 1522 1659 1526
rect 1695 1524 1699 1528
rect 111 1507 115 1511
rect 135 1505 139 1509
rect 175 1505 179 1509
rect 223 1505 227 1509
rect 279 1505 283 1509
rect 335 1505 339 1509
rect 399 1505 403 1509
rect 463 1505 467 1509
rect 535 1505 539 1509
rect 607 1505 611 1509
rect 687 1505 691 1509
rect 775 1505 779 1509
rect 871 1505 875 1509
rect 975 1505 979 1509
rect 1079 1505 1083 1509
rect 1175 1505 1179 1509
rect 1271 1505 1275 1509
rect 1359 1505 1363 1509
rect 1439 1505 1443 1509
rect 1519 1505 1523 1509
rect 1599 1505 1603 1509
rect 1655 1505 1659 1509
rect 1695 1507 1699 1511
rect 111 1469 115 1473
rect 175 1471 179 1475
rect 207 1471 211 1475
rect 239 1471 243 1475
rect 271 1471 275 1475
rect 303 1471 307 1475
rect 335 1471 339 1475
rect 367 1471 371 1475
rect 399 1471 403 1475
rect 431 1471 435 1475
rect 463 1471 467 1475
rect 495 1471 499 1475
rect 527 1471 531 1475
rect 559 1471 563 1475
rect 591 1471 595 1475
rect 623 1471 627 1475
rect 663 1471 667 1475
rect 703 1471 707 1475
rect 743 1471 747 1475
rect 775 1471 779 1475
rect 807 1472 811 1476
rect 895 1472 899 1476
rect 935 1472 939 1476
rect 1023 1472 1027 1476
rect 1079 1471 1083 1475
rect 1111 1472 1115 1476
rect 1167 1471 1171 1475
rect 1199 1471 1203 1475
rect 1239 1471 1243 1475
rect 1279 1471 1283 1475
rect 1319 1471 1323 1475
rect 1359 1471 1363 1475
rect 1399 1471 1403 1475
rect 1439 1471 1443 1475
rect 1479 1471 1483 1475
rect 1519 1471 1523 1475
rect 1559 1471 1563 1475
rect 1591 1471 1595 1475
rect 1623 1471 1627 1475
rect 1655 1471 1659 1475
rect 1695 1469 1699 1473
rect 111 1452 115 1456
rect 175 1454 179 1458
rect 207 1454 211 1458
rect 239 1454 243 1458
rect 271 1454 275 1458
rect 303 1454 307 1458
rect 335 1454 339 1458
rect 367 1454 371 1458
rect 399 1454 403 1458
rect 431 1454 435 1458
rect 463 1454 467 1458
rect 495 1454 499 1458
rect 527 1454 531 1458
rect 559 1454 563 1458
rect 591 1454 595 1458
rect 623 1454 627 1458
rect 663 1454 667 1458
rect 703 1454 707 1458
rect 743 1454 747 1458
rect 775 1453 779 1457
rect 807 1453 811 1457
rect 935 1453 939 1457
rect 1039 1451 1043 1455
rect 1079 1454 1083 1458
rect 1127 1451 1131 1455
rect 1167 1454 1171 1458
rect 1199 1454 1203 1458
rect 1239 1454 1243 1458
rect 1279 1453 1283 1457
rect 1319 1454 1323 1458
rect 1359 1454 1363 1458
rect 1399 1454 1403 1458
rect 1439 1454 1443 1458
rect 1479 1454 1483 1458
rect 1519 1454 1523 1458
rect 1559 1454 1563 1458
rect 1591 1454 1595 1458
rect 1623 1454 1627 1458
rect 1655 1454 1659 1458
rect 1695 1452 1699 1456
rect 895 1444 899 1448
rect 767 1411 771 1415
rect 839 1411 843 1415
rect 975 1411 979 1415
rect 895 1406 899 1410
rect 1063 1396 1067 1400
rect 1151 1396 1155 1400
rect 111 1388 115 1392
rect 135 1386 139 1390
rect 167 1386 171 1390
rect 199 1386 203 1390
rect 231 1386 235 1390
rect 263 1386 267 1390
rect 295 1386 299 1390
rect 327 1386 331 1390
rect 359 1386 363 1390
rect 391 1386 395 1390
rect 423 1386 427 1390
rect 455 1386 459 1390
rect 487 1386 491 1390
rect 519 1386 523 1390
rect 551 1386 555 1390
rect 583 1386 587 1390
rect 615 1386 619 1390
rect 647 1386 651 1390
rect 679 1386 683 1390
rect 719 1389 723 1393
rect 807 1391 811 1395
rect 1023 1386 1027 1390
rect 1111 1387 1115 1391
rect 1199 1386 1203 1390
rect 1263 1389 1267 1393
rect 1319 1387 1323 1391
rect 1415 1386 1419 1390
rect 1479 1389 1483 1393
rect 1535 1386 1539 1390
rect 1583 1386 1587 1390
rect 1623 1386 1627 1390
rect 1655 1386 1659 1390
rect 1695 1388 1699 1392
rect 111 1371 115 1375
rect 135 1369 139 1373
rect 167 1369 171 1373
rect 199 1369 203 1373
rect 231 1369 235 1373
rect 263 1369 267 1373
rect 295 1369 299 1373
rect 327 1369 331 1373
rect 359 1369 363 1373
rect 391 1369 395 1373
rect 423 1369 427 1373
rect 455 1369 459 1373
rect 487 1369 491 1373
rect 519 1369 523 1373
rect 551 1369 555 1373
rect 583 1369 587 1373
rect 615 1369 619 1373
rect 647 1369 651 1373
rect 679 1369 683 1373
rect 735 1362 739 1366
rect 767 1364 771 1368
rect 807 1368 811 1372
rect 839 1364 843 1368
rect 887 1368 891 1372
rect 1023 1369 1027 1373
rect 1063 1368 1067 1372
rect 1111 1369 1115 1373
rect 1151 1368 1155 1372
rect 1199 1369 1203 1373
rect 1247 1368 1251 1372
rect 975 1364 979 1368
rect 1319 1368 1323 1372
rect 1415 1369 1419 1373
rect 1463 1368 1467 1372
rect 1535 1369 1539 1373
rect 1583 1369 1587 1373
rect 1623 1369 1627 1373
rect 1655 1369 1659 1373
rect 1695 1371 1699 1375
rect 111 1313 115 1317
rect 135 1315 139 1319
rect 167 1315 171 1319
rect 199 1315 203 1319
rect 231 1315 235 1319
rect 263 1315 267 1319
rect 295 1315 299 1319
rect 327 1315 331 1319
rect 359 1315 363 1319
rect 391 1315 395 1319
rect 423 1315 427 1319
rect 455 1315 459 1319
rect 487 1315 491 1319
rect 519 1315 523 1319
rect 551 1315 555 1319
rect 583 1315 587 1319
rect 615 1315 619 1319
rect 647 1315 651 1319
rect 679 1315 683 1319
rect 711 1315 715 1319
rect 743 1316 747 1320
rect 823 1316 827 1320
rect 903 1316 907 1320
rect 983 1320 987 1324
rect 1023 1316 1027 1320
rect 1063 1316 1067 1320
rect 1159 1316 1163 1320
rect 1215 1316 1219 1320
rect 1303 1316 1307 1320
rect 1391 1315 1395 1319
rect 1423 1315 1427 1319
rect 1455 1316 1459 1320
rect 1495 1315 1499 1319
rect 1527 1315 1531 1319
rect 1559 1315 1563 1319
rect 1591 1315 1595 1319
rect 1623 1315 1627 1319
rect 1655 1315 1659 1319
rect 1695 1313 1699 1317
rect 111 1296 115 1300
rect 135 1298 139 1302
rect 167 1298 171 1302
rect 199 1298 203 1302
rect 231 1298 235 1302
rect 263 1298 267 1302
rect 295 1298 299 1302
rect 327 1298 331 1302
rect 359 1298 363 1302
rect 391 1298 395 1302
rect 423 1298 427 1302
rect 455 1298 459 1302
rect 487 1298 491 1302
rect 519 1298 523 1302
rect 551 1298 555 1302
rect 583 1298 587 1302
rect 615 1298 619 1302
rect 647 1298 651 1302
rect 679 1298 683 1302
rect 711 1298 715 1302
rect 1063 1297 1067 1301
rect 1175 1295 1179 1299
rect 1215 1297 1219 1301
rect 1303 1297 1307 1301
rect 1391 1297 1395 1301
rect 1423 1298 1427 1302
rect 1495 1298 1499 1302
rect 1527 1298 1531 1302
rect 1559 1298 1563 1302
rect 1591 1298 1595 1302
rect 1623 1298 1627 1302
rect 1655 1298 1659 1302
rect 1695 1296 1699 1300
rect 1023 1288 1027 1292
rect 1455 1288 1459 1292
rect 751 1278 755 1282
rect 831 1278 835 1282
rect 911 1278 915 1282
rect 983 1273 987 1277
rect 775 1215 779 1219
rect 1087 1215 1091 1219
rect 1015 1210 1019 1214
rect 111 1192 115 1196
rect 135 1190 139 1194
rect 167 1190 171 1194
rect 199 1190 203 1194
rect 231 1190 235 1194
rect 263 1190 267 1194
rect 295 1190 299 1194
rect 327 1190 331 1194
rect 359 1190 363 1194
rect 391 1190 395 1194
rect 423 1190 427 1194
rect 455 1190 459 1194
rect 487 1190 491 1194
rect 519 1190 523 1194
rect 551 1190 555 1194
rect 583 1190 587 1194
rect 615 1190 619 1194
rect 647 1190 651 1194
rect 679 1190 683 1194
rect 711 1190 715 1194
rect 743 1190 747 1194
rect 811 1191 815 1195
rect 959 1193 963 1197
rect 1127 1190 1131 1194
rect 1159 1190 1163 1194
rect 1215 1193 1219 1197
rect 1255 1190 1259 1194
rect 1295 1193 1299 1197
rect 1343 1190 1347 1194
rect 1375 1190 1379 1194
rect 1407 1190 1411 1194
rect 1439 1190 1443 1194
rect 1479 1190 1483 1194
rect 1519 1190 1523 1194
rect 1559 1190 1563 1194
rect 1591 1190 1595 1194
rect 1623 1190 1627 1194
rect 1655 1190 1659 1194
rect 1695 1192 1699 1196
rect 111 1175 115 1179
rect 135 1173 139 1177
rect 167 1173 171 1177
rect 199 1173 203 1177
rect 231 1173 235 1177
rect 263 1173 267 1177
rect 295 1173 299 1177
rect 327 1173 331 1177
rect 359 1173 363 1177
rect 391 1173 395 1177
rect 423 1173 427 1177
rect 455 1173 459 1177
rect 487 1173 491 1177
rect 519 1173 523 1177
rect 551 1173 555 1177
rect 583 1173 587 1177
rect 615 1173 619 1177
rect 647 1173 651 1177
rect 679 1173 683 1177
rect 711 1173 715 1177
rect 743 1173 747 1177
rect 839 1176 843 1180
rect 775 1168 779 1172
rect 1007 1172 1011 1176
rect 1127 1173 1131 1177
rect 1159 1173 1163 1177
rect 1199 1172 1203 1176
rect 1255 1173 1259 1177
rect 1343 1173 1347 1177
rect 1375 1173 1379 1177
rect 1407 1173 1411 1177
rect 1439 1173 1443 1177
rect 1479 1173 1483 1177
rect 1519 1173 1523 1177
rect 1559 1173 1563 1177
rect 1591 1173 1595 1177
rect 1623 1173 1627 1177
rect 1655 1173 1659 1177
rect 1695 1175 1699 1179
rect 975 1166 979 1170
rect 1087 1168 1091 1172
rect 1311 1166 1315 1170
rect 111 1117 115 1121
rect 135 1119 139 1123
rect 167 1119 171 1123
rect 199 1119 203 1123
rect 231 1119 235 1123
rect 263 1119 267 1123
rect 295 1119 299 1123
rect 327 1119 331 1123
rect 359 1119 363 1123
rect 391 1119 395 1123
rect 423 1119 427 1123
rect 455 1119 459 1123
rect 487 1119 491 1123
rect 519 1119 523 1123
rect 551 1119 555 1123
rect 583 1120 587 1124
rect 687 1116 691 1120
rect 799 1120 803 1124
rect 847 1122 851 1126
rect 935 1119 939 1123
rect 967 1119 971 1123
rect 999 1120 1003 1124
rect 1031 1119 1035 1123
rect 1063 1119 1067 1123
rect 1095 1120 1099 1124
rect 1135 1119 1139 1123
rect 1167 1120 1171 1124
rect 1247 1124 1251 1128
rect 1287 1119 1291 1123
rect 1335 1122 1339 1126
rect 1423 1119 1427 1123
rect 1455 1119 1459 1123
rect 1487 1119 1491 1123
rect 1519 1119 1523 1123
rect 1559 1119 1563 1123
rect 1591 1119 1595 1123
rect 1623 1119 1627 1123
rect 1655 1119 1659 1123
rect 1695 1117 1699 1121
rect 111 1100 115 1104
rect 135 1102 139 1106
rect 167 1102 171 1106
rect 199 1102 203 1106
rect 231 1102 235 1106
rect 263 1102 267 1106
rect 295 1102 299 1106
rect 327 1102 331 1106
rect 359 1102 363 1106
rect 391 1102 395 1106
rect 423 1102 427 1106
rect 455 1102 459 1106
rect 487 1102 491 1106
rect 519 1102 523 1106
rect 551 1102 555 1106
rect 659 1101 663 1105
rect 935 1102 939 1106
rect 967 1102 971 1106
rect 1031 1102 1035 1106
rect 1063 1102 1067 1106
rect 1135 1102 1139 1106
rect 1287 1102 1291 1106
rect 1423 1102 1427 1106
rect 1455 1102 1459 1106
rect 1487 1102 1491 1106
rect 1519 1102 1523 1106
rect 1559 1102 1563 1106
rect 1591 1102 1595 1106
rect 1623 1102 1627 1106
rect 1655 1102 1659 1106
rect 799 1097 803 1101
rect 999 1097 1003 1101
rect 1695 1100 1699 1104
rect 1095 1092 1099 1096
rect 591 1082 595 1086
rect 847 1081 851 1085
rect 1175 1082 1179 1086
rect 1247 1077 1251 1081
rect 1335 1081 1339 1085
rect 503 1015 507 1019
rect 407 1010 411 1014
rect 583 1011 587 1015
rect 711 1011 715 1015
rect 823 1005 827 1009
rect 975 1005 979 1009
rect 1063 1000 1067 1004
rect 1199 1000 1203 1004
rect 1327 1000 1331 1004
rect 1367 1000 1371 1004
rect 111 992 115 996
rect 135 990 139 994
rect 167 990 171 994
rect 199 990 203 994
rect 231 990 235 994
rect 263 990 267 994
rect 327 993 331 997
rect 919 990 923 994
rect 1119 993 1123 997
rect 1167 990 1171 994
rect 1247 993 1251 997
rect 1295 990 1299 994
rect 1407 990 1411 994
rect 1439 990 1443 994
rect 1479 990 1483 994
rect 1519 990 1523 994
rect 1559 990 1563 994
rect 1591 990 1595 994
rect 1623 990 1627 994
rect 1655 990 1659 994
rect 1695 992 1699 996
rect 111 975 115 979
rect 135 973 139 977
rect 167 973 171 977
rect 199 973 203 977
rect 231 973 235 977
rect 263 973 267 977
rect 399 972 403 976
rect 343 966 347 970
rect 503 968 507 972
rect 583 970 587 974
rect 711 970 715 974
rect 919 973 923 977
rect 1063 972 1067 976
rect 1167 973 1171 977
rect 1199 972 1203 976
rect 1295 973 1299 977
rect 1327 972 1331 976
rect 1367 972 1371 976
rect 1407 973 1411 977
rect 1439 973 1443 977
rect 1479 973 1483 977
rect 1519 973 1523 977
rect 1559 973 1563 977
rect 1591 973 1595 977
rect 1623 973 1627 977
rect 1655 973 1659 977
rect 1695 975 1699 979
rect 815 965 819 969
rect 967 965 971 969
rect 1135 966 1139 970
rect 1263 966 1267 970
rect 111 917 115 921
rect 135 919 139 923
rect 167 919 171 923
rect 199 920 203 924
rect 279 924 283 928
rect 319 920 323 924
rect 399 924 403 928
rect 591 922 595 926
rect 463 916 467 920
rect 679 920 683 924
rect 727 922 731 926
rect 815 919 819 923
rect 863 922 867 926
rect 1391 926 1395 930
rect 951 919 955 923
rect 983 920 987 924
rect 1039 919 1043 923
rect 1071 920 1075 924
rect 1111 919 1115 923
rect 1143 920 1147 924
rect 1239 919 1243 923
rect 1271 920 1275 924
rect 1423 919 1427 923
rect 1455 920 1459 924
rect 1519 919 1523 923
rect 1559 919 1563 923
rect 1591 919 1595 923
rect 1623 919 1627 923
rect 1655 919 1659 923
rect 1695 917 1699 921
rect 111 900 115 904
rect 135 902 139 906
rect 167 902 171 906
rect 435 901 439 905
rect 815 902 819 906
rect 951 902 955 906
rect 679 897 683 901
rect 999 899 1003 903
rect 1039 902 1043 906
rect 1111 901 1115 905
rect 1143 901 1147 905
rect 1239 901 1243 905
rect 1271 901 1275 905
rect 1375 899 1379 903
rect 1423 902 1427 906
rect 1471 899 1475 903
rect 1519 902 1523 906
rect 1559 902 1563 906
rect 1591 902 1595 906
rect 1623 902 1627 906
rect 1655 902 1659 906
rect 1695 900 1699 904
rect 1071 892 1075 896
rect 207 882 211 886
rect 327 882 331 886
rect 279 877 283 881
rect 399 877 403 881
rect 591 881 595 885
rect 727 881 731 885
rect 863 881 867 885
rect 231 819 235 823
rect 407 819 411 823
rect 815 819 819 823
rect 663 813 667 817
rect 1423 808 1427 812
rect 1471 808 1475 812
rect 111 800 115 804
rect 951 803 955 807
rect 135 798 139 802
rect 559 798 563 802
rect 1031 801 1035 805
rect 1103 798 1107 802
rect 1167 801 1171 805
rect 1247 801 1251 805
rect 1295 799 1299 803
rect 1327 799 1331 803
rect 1519 798 1523 802
rect 1559 798 1563 802
rect 1591 798 1595 802
rect 1623 798 1627 802
rect 1655 798 1659 802
rect 1695 800 1699 804
rect 111 783 115 787
rect 135 781 139 785
rect 231 778 235 782
rect 407 778 411 782
rect 559 781 563 785
rect 815 778 819 782
rect 951 780 955 784
rect 1015 780 1019 784
rect 1103 781 1107 785
rect 1231 780 1235 784
rect 1295 781 1299 785
rect 1327 780 1331 784
rect 1423 780 1427 784
rect 1471 780 1475 784
rect 1519 781 1523 785
rect 1559 781 1563 785
rect 1591 781 1595 785
rect 1623 781 1627 785
rect 1655 781 1659 785
rect 1695 783 1699 787
rect 655 773 659 777
rect 1183 774 1187 778
rect 111 721 115 725
rect 135 724 139 728
rect 215 728 219 732
rect 287 726 291 730
rect 391 728 395 732
rect 767 731 771 735
rect 999 731 1003 735
rect 615 726 619 730
rect 471 720 475 724
rect 719 724 723 728
rect 863 723 867 727
rect 911 726 915 730
rect 1087 724 1091 728
rect 1167 728 1171 732
rect 1207 724 1211 728
rect 1247 723 1251 727
rect 1279 723 1283 727
rect 1311 723 1315 727
rect 1343 723 1347 727
rect 1375 723 1379 727
rect 1407 723 1411 727
rect 1439 723 1443 727
rect 1479 723 1483 727
rect 1519 723 1523 727
rect 1559 723 1563 727
rect 1591 723 1595 727
rect 1623 723 1627 727
rect 1655 723 1659 727
rect 1695 721 1699 725
rect 111 704 115 708
rect 443 705 447 709
rect 863 706 867 710
rect 1247 706 1251 710
rect 1279 706 1283 710
rect 1311 706 1315 710
rect 1343 706 1347 710
rect 1375 706 1379 710
rect 1407 706 1411 710
rect 1439 706 1443 710
rect 1479 706 1483 710
rect 1519 706 1523 710
rect 1559 706 1563 710
rect 1591 706 1595 710
rect 1623 706 1627 710
rect 1655 706 1659 710
rect 719 701 723 705
rect 1695 704 1699 708
rect 1207 696 1211 700
rect 775 691 779 695
rect 1007 691 1011 695
rect 143 686 147 690
rect 215 681 219 685
rect 287 685 291 689
rect 391 681 395 685
rect 615 685 619 689
rect 911 685 915 689
rect 1095 686 1099 690
rect 1167 681 1171 685
rect 207 623 211 627
rect 287 618 291 622
rect 407 618 411 622
rect 535 619 539 623
rect 767 619 771 623
rect 903 623 907 627
rect 1119 623 1123 627
rect 1335 623 1339 627
rect 999 618 1003 622
rect 1215 618 1219 622
rect 111 600 115 604
rect 135 598 139 602
rect 167 598 171 602
rect 671 598 675 602
rect 1415 598 1419 602
rect 1479 598 1483 602
rect 1543 598 1547 602
rect 1607 598 1611 602
rect 1655 598 1659 602
rect 1695 600 1699 604
rect 111 583 115 587
rect 135 581 139 585
rect 167 581 171 585
rect 207 576 211 580
rect 279 580 283 584
rect 399 580 403 584
rect 535 578 539 582
rect 671 581 675 585
rect 767 578 771 582
rect 903 576 907 580
rect 991 580 995 584
rect 1119 576 1123 580
rect 1207 580 1211 584
rect 1415 581 1419 585
rect 1479 581 1483 585
rect 1543 581 1547 585
rect 1607 581 1611 585
rect 1655 581 1659 585
rect 1695 583 1699 587
rect 1335 576 1339 580
rect 111 529 115 533
rect 135 531 139 535
rect 167 532 171 536
rect 247 536 251 540
rect 303 534 307 538
rect 391 532 395 536
rect 471 536 475 540
rect 535 528 539 532
rect 647 532 651 536
rect 727 536 731 540
rect 775 532 779 536
rect 871 536 875 540
rect 927 532 931 536
rect 1031 536 1035 540
rect 1095 532 1099 536
rect 1199 536 1203 540
rect 1287 528 1291 532
rect 1423 531 1427 535
rect 1479 531 1483 535
rect 1527 531 1531 535
rect 1575 531 1579 535
rect 1623 531 1627 535
rect 1655 531 1659 535
rect 1695 529 1699 533
rect 111 512 115 516
rect 135 514 139 518
rect 507 513 511 517
rect 1259 513 1263 517
rect 1423 514 1427 518
rect 1479 514 1483 518
rect 1527 514 1531 518
rect 1575 514 1579 518
rect 1623 514 1627 518
rect 1655 514 1659 518
rect 1695 512 1699 516
rect 175 494 179 498
rect 247 489 251 493
rect 303 493 307 497
rect 399 494 403 498
rect 655 494 659 498
rect 783 494 787 498
rect 935 494 939 498
rect 1103 494 1107 498
rect 471 489 475 493
rect 727 489 731 493
rect 871 489 875 493
rect 1031 489 1035 493
rect 1199 489 1203 493
rect 375 395 379 399
rect 615 395 619 399
rect 303 390 307 394
rect 543 390 547 394
rect 671 391 675 395
rect 951 390 955 394
rect 1231 391 1235 395
rect 1359 385 1363 389
rect 111 372 115 376
rect 135 370 139 374
rect 167 370 171 374
rect 199 370 203 374
rect 231 370 235 374
rect 263 370 267 374
rect 415 370 419 374
rect 447 370 451 374
rect 487 373 491 377
rect 755 371 759 375
rect 903 370 907 374
rect 1031 373 1035 377
rect 1439 375 1443 379
rect 1075 371 1079 375
rect 1319 370 1323 374
rect 1479 370 1483 374
rect 1519 370 1523 374
rect 1559 370 1563 374
rect 1591 370 1595 374
rect 1623 370 1627 374
rect 1655 370 1659 374
rect 1695 372 1699 376
rect 111 355 115 359
rect 135 353 139 357
rect 167 353 171 357
rect 199 353 203 357
rect 231 353 235 357
rect 263 353 267 357
rect 295 352 299 356
rect 415 353 419 357
rect 447 353 451 357
rect 535 352 539 356
rect 783 356 787 360
rect 375 348 379 352
rect 503 346 507 350
rect 615 348 619 352
rect 671 350 675 354
rect 903 353 907 357
rect 943 352 947 356
rect 1103 356 1107 360
rect 1047 346 1051 350
rect 1231 350 1235 354
rect 1319 353 1323 357
rect 1439 352 1443 356
rect 1479 353 1483 357
rect 1519 353 1523 357
rect 1559 353 1563 357
rect 1591 353 1595 357
rect 1623 353 1627 357
rect 1655 353 1659 357
rect 1695 355 1699 359
rect 1351 345 1355 349
rect 1199 307 1203 311
rect 111 297 115 301
rect 135 299 139 303
rect 167 299 171 303
rect 199 299 203 303
rect 231 299 235 303
rect 263 299 267 303
rect 295 299 299 303
rect 327 299 331 303
rect 359 299 363 303
rect 391 299 395 303
rect 423 299 427 303
rect 455 299 459 303
rect 487 299 491 303
rect 519 299 523 303
rect 551 299 555 303
rect 599 302 603 306
rect 703 302 707 306
rect 807 302 811 306
rect 911 302 915 306
rect 999 299 1003 303
rect 1031 299 1035 303
rect 1063 299 1067 303
rect 1111 302 1115 306
rect 1287 300 1291 304
rect 1319 299 1323 303
rect 1351 299 1355 303
rect 1383 299 1387 303
rect 1415 299 1419 303
rect 1447 299 1451 303
rect 1479 299 1483 303
rect 1519 299 1523 303
rect 1559 299 1563 303
rect 1591 299 1595 303
rect 1623 299 1627 303
rect 1655 299 1659 303
rect 1695 297 1699 301
rect 111 280 115 284
rect 135 282 139 286
rect 167 282 171 286
rect 199 282 203 286
rect 231 282 235 286
rect 263 282 267 286
rect 295 282 299 286
rect 327 282 331 286
rect 359 282 363 286
rect 391 282 395 286
rect 423 282 427 286
rect 455 282 459 286
rect 487 282 491 286
rect 519 282 523 286
rect 551 282 555 286
rect 999 282 1003 286
rect 1031 282 1035 286
rect 1063 282 1067 286
rect 1319 282 1323 286
rect 1351 282 1355 286
rect 1383 282 1387 286
rect 1415 282 1419 286
rect 1447 282 1451 286
rect 1479 282 1483 286
rect 1519 282 1523 286
rect 1559 282 1563 286
rect 1591 282 1595 286
rect 1623 282 1627 286
rect 1655 282 1659 286
rect 1287 277 1291 281
rect 1695 280 1699 284
rect 1207 267 1211 271
rect 599 261 603 265
rect 703 261 707 265
rect 807 261 811 265
rect 911 261 915 265
rect 1111 261 1115 265
rect 695 231 699 235
rect 967 231 971 235
rect 839 225 843 229
rect 111 212 115 216
rect 919 215 923 219
rect 183 210 187 214
rect 215 210 219 214
rect 247 210 251 214
rect 279 210 283 214
rect 311 210 315 214
rect 343 210 347 214
rect 375 210 379 214
rect 407 210 411 214
rect 439 210 443 214
rect 471 210 475 214
rect 503 210 507 214
rect 535 210 539 214
rect 567 210 571 214
rect 599 210 603 214
rect 639 210 643 214
rect 791 210 795 214
rect 1063 210 1067 214
rect 1103 210 1107 214
rect 1143 210 1147 214
rect 1183 210 1187 214
rect 1223 210 1227 214
rect 1263 210 1267 214
rect 1303 210 1307 214
rect 1343 210 1347 214
rect 1375 210 1379 214
rect 1407 210 1411 214
rect 1439 210 1443 214
rect 1479 210 1483 214
rect 1519 210 1523 214
rect 1559 210 1563 214
rect 1591 210 1595 214
rect 1623 210 1627 214
rect 1655 210 1659 214
rect 1695 212 1699 216
rect 111 195 115 199
rect 183 193 187 197
rect 215 193 219 197
rect 247 193 251 197
rect 279 193 283 197
rect 311 193 315 197
rect 343 193 347 197
rect 375 193 379 197
rect 407 193 411 197
rect 439 193 443 197
rect 471 193 475 197
rect 503 193 507 197
rect 535 193 539 197
rect 567 193 571 197
rect 599 193 603 197
rect 639 193 643 197
rect 695 190 699 194
rect 791 193 795 197
rect 919 192 923 196
rect 967 190 971 194
rect 1063 193 1067 197
rect 1103 193 1107 197
rect 1143 193 1147 197
rect 1183 193 1187 197
rect 1223 193 1227 197
rect 1263 193 1267 197
rect 1303 193 1307 197
rect 1343 193 1347 197
rect 1375 193 1379 197
rect 1407 193 1411 197
rect 1439 193 1443 197
rect 1479 193 1483 197
rect 1519 193 1523 197
rect 1559 193 1563 197
rect 1591 193 1595 197
rect 1623 193 1627 197
rect 1655 193 1659 197
rect 1695 195 1699 199
rect 831 185 835 189
rect 111 161 115 165
rect 135 163 139 167
rect 167 163 171 167
rect 215 163 219 167
rect 263 163 267 167
rect 311 163 315 167
rect 367 163 371 167
rect 415 163 419 167
rect 471 163 475 167
rect 535 163 539 167
rect 607 163 611 167
rect 687 163 691 167
rect 775 163 779 167
rect 863 163 867 167
rect 959 163 963 167
rect 1055 163 1059 167
rect 1151 163 1155 167
rect 1239 163 1243 167
rect 1327 163 1331 167
rect 1415 163 1419 167
rect 1503 163 1507 167
rect 1591 163 1595 167
rect 1655 163 1659 167
rect 1695 161 1699 165
rect 111 144 115 148
rect 135 146 139 150
rect 167 146 171 150
rect 215 146 219 150
rect 263 146 267 150
rect 311 146 315 150
rect 367 146 371 150
rect 415 146 419 150
rect 471 146 475 150
rect 535 146 539 150
rect 607 146 611 150
rect 687 146 691 150
rect 775 146 779 150
rect 863 146 867 150
rect 959 146 963 150
rect 1055 146 1059 150
rect 1151 146 1155 150
rect 1239 146 1243 150
rect 1327 146 1331 150
rect 1415 146 1419 150
rect 1503 146 1507 150
rect 1591 146 1595 150
rect 1655 146 1659 150
rect 1695 144 1699 148
rect 111 104 115 108
rect 135 102 139 106
rect 167 102 171 106
rect 199 102 203 106
rect 231 102 235 106
rect 263 102 267 106
rect 295 102 299 106
rect 327 102 331 106
rect 359 102 363 106
rect 391 102 395 106
rect 423 102 427 106
rect 455 102 459 106
rect 487 102 491 106
rect 519 102 523 106
rect 551 102 555 106
rect 607 102 611 106
rect 671 102 675 106
rect 743 102 747 106
rect 823 102 827 106
rect 903 102 907 106
rect 983 102 987 106
rect 1055 102 1059 106
rect 1119 102 1123 106
rect 1175 102 1179 106
rect 1223 102 1227 106
rect 1271 102 1275 106
rect 1311 102 1315 106
rect 1343 102 1347 106
rect 1375 102 1379 106
rect 1407 102 1411 106
rect 1439 102 1443 106
rect 1479 102 1483 106
rect 1519 102 1523 106
rect 1559 102 1563 106
rect 1591 102 1595 106
rect 1623 102 1627 106
rect 1655 102 1659 106
rect 1695 104 1699 108
rect 111 87 115 91
rect 135 85 139 89
rect 167 85 171 89
rect 199 85 203 89
rect 231 85 235 89
rect 263 85 267 89
rect 295 85 299 89
rect 327 85 331 89
rect 359 85 363 89
rect 391 85 395 89
rect 423 85 427 89
rect 455 85 459 89
rect 487 85 491 89
rect 519 85 523 89
rect 551 85 555 89
rect 607 85 611 89
rect 671 85 675 89
rect 743 85 747 89
rect 823 85 827 89
rect 903 85 907 89
rect 983 85 987 89
rect 1055 85 1059 89
rect 1119 85 1123 89
rect 1175 85 1179 89
rect 1223 85 1227 89
rect 1271 85 1275 89
rect 1311 85 1315 89
rect 1343 85 1347 89
rect 1375 85 1379 89
rect 1407 85 1411 89
rect 1439 85 1443 89
rect 1479 85 1483 89
rect 1519 85 1523 89
rect 1559 85 1563 89
rect 1591 85 1595 89
rect 1623 85 1627 89
rect 1655 85 1659 89
rect 1695 87 1699 91
<< m3 >>
rect 111 1762 115 1763
rect 111 1757 115 1758
rect 151 1762 155 1763
rect 112 1754 114 1757
rect 151 1756 155 1758
rect 183 1762 187 1763
rect 183 1756 187 1758
rect 215 1762 219 1763
rect 215 1756 219 1758
rect 247 1762 251 1763
rect 247 1756 251 1758
rect 279 1762 283 1763
rect 279 1756 283 1758
rect 311 1762 315 1763
rect 311 1756 315 1758
rect 343 1762 347 1763
rect 343 1756 347 1758
rect 375 1762 379 1763
rect 375 1756 379 1758
rect 407 1762 411 1763
rect 407 1756 411 1758
rect 439 1762 443 1763
rect 439 1756 443 1758
rect 471 1762 475 1763
rect 471 1756 475 1758
rect 503 1762 507 1763
rect 503 1756 507 1758
rect 535 1762 539 1763
rect 535 1756 539 1758
rect 567 1762 571 1763
rect 567 1756 571 1758
rect 599 1762 603 1763
rect 599 1756 603 1758
rect 631 1762 635 1763
rect 631 1756 635 1758
rect 663 1762 667 1763
rect 663 1756 667 1758
rect 695 1762 699 1763
rect 695 1756 699 1758
rect 727 1762 731 1763
rect 727 1756 731 1758
rect 759 1762 763 1763
rect 759 1756 763 1758
rect 791 1762 795 1763
rect 791 1756 795 1758
rect 823 1762 827 1763
rect 823 1756 827 1758
rect 855 1762 859 1763
rect 855 1756 859 1758
rect 887 1762 891 1763
rect 887 1756 891 1758
rect 919 1762 923 1763
rect 919 1756 923 1758
rect 951 1762 955 1763
rect 951 1756 955 1758
rect 983 1762 987 1763
rect 983 1756 987 1758
rect 1695 1762 1699 1763
rect 1695 1757 1699 1758
rect 150 1755 156 1756
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 150 1751 151 1755
rect 155 1751 156 1755
rect 150 1750 156 1751
rect 182 1755 188 1756
rect 182 1751 183 1755
rect 187 1751 188 1755
rect 182 1750 188 1751
rect 214 1755 220 1756
rect 214 1751 215 1755
rect 219 1751 220 1755
rect 214 1750 220 1751
rect 246 1755 252 1756
rect 246 1751 247 1755
rect 251 1751 252 1755
rect 246 1750 252 1751
rect 278 1755 284 1756
rect 278 1751 279 1755
rect 283 1751 284 1755
rect 278 1750 284 1751
rect 310 1755 316 1756
rect 310 1751 311 1755
rect 315 1751 316 1755
rect 310 1750 316 1751
rect 342 1755 348 1756
rect 342 1751 343 1755
rect 347 1751 348 1755
rect 342 1750 348 1751
rect 374 1755 380 1756
rect 374 1751 375 1755
rect 379 1751 380 1755
rect 374 1750 380 1751
rect 406 1755 412 1756
rect 406 1751 407 1755
rect 411 1751 412 1755
rect 406 1750 412 1751
rect 438 1755 444 1756
rect 438 1751 439 1755
rect 443 1751 444 1755
rect 438 1750 444 1751
rect 470 1755 476 1756
rect 470 1751 471 1755
rect 475 1751 476 1755
rect 470 1750 476 1751
rect 502 1755 508 1756
rect 502 1751 503 1755
rect 507 1751 508 1755
rect 502 1750 508 1751
rect 534 1755 540 1756
rect 534 1751 535 1755
rect 539 1751 540 1755
rect 534 1750 540 1751
rect 566 1755 572 1756
rect 566 1751 567 1755
rect 571 1751 572 1755
rect 566 1750 572 1751
rect 598 1755 604 1756
rect 598 1751 599 1755
rect 603 1751 604 1755
rect 598 1750 604 1751
rect 630 1755 636 1756
rect 630 1751 631 1755
rect 635 1751 636 1755
rect 630 1750 636 1751
rect 662 1755 668 1756
rect 662 1751 663 1755
rect 667 1751 668 1755
rect 662 1750 668 1751
rect 694 1755 700 1756
rect 694 1751 695 1755
rect 699 1751 700 1755
rect 694 1750 700 1751
rect 726 1755 732 1756
rect 726 1751 727 1755
rect 731 1751 732 1755
rect 726 1750 732 1751
rect 758 1755 764 1756
rect 758 1751 759 1755
rect 763 1751 764 1755
rect 758 1750 764 1751
rect 790 1755 796 1756
rect 790 1751 791 1755
rect 795 1751 796 1755
rect 790 1750 796 1751
rect 822 1755 828 1756
rect 822 1751 823 1755
rect 827 1751 828 1755
rect 822 1750 828 1751
rect 854 1755 860 1756
rect 854 1751 855 1755
rect 859 1751 860 1755
rect 854 1750 860 1751
rect 886 1755 892 1756
rect 886 1751 887 1755
rect 891 1751 892 1755
rect 886 1750 892 1751
rect 918 1755 924 1756
rect 918 1751 919 1755
rect 923 1751 924 1755
rect 918 1750 924 1751
rect 950 1755 956 1756
rect 950 1751 951 1755
rect 955 1751 956 1755
rect 950 1750 956 1751
rect 982 1755 988 1756
rect 982 1751 983 1755
rect 987 1751 988 1755
rect 1696 1754 1698 1757
rect 982 1750 988 1751
rect 1694 1753 1700 1754
rect 110 1748 116 1749
rect 1694 1749 1695 1753
rect 1699 1749 1700 1753
rect 1694 1748 1700 1749
rect 150 1738 156 1739
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 150 1734 151 1738
rect 155 1734 156 1738
rect 150 1733 156 1734
rect 182 1738 188 1739
rect 182 1734 183 1738
rect 187 1734 188 1738
rect 182 1733 188 1734
rect 214 1738 220 1739
rect 214 1734 215 1738
rect 219 1734 220 1738
rect 214 1733 220 1734
rect 246 1738 252 1739
rect 246 1734 247 1738
rect 251 1734 252 1738
rect 246 1733 252 1734
rect 278 1738 284 1739
rect 278 1734 279 1738
rect 283 1734 284 1738
rect 278 1733 284 1734
rect 310 1738 316 1739
rect 310 1734 311 1738
rect 315 1734 316 1738
rect 310 1733 316 1734
rect 342 1738 348 1739
rect 342 1734 343 1738
rect 347 1734 348 1738
rect 342 1733 348 1734
rect 374 1738 380 1739
rect 374 1734 375 1738
rect 379 1734 380 1738
rect 374 1733 380 1734
rect 406 1738 412 1739
rect 406 1734 407 1738
rect 411 1734 412 1738
rect 406 1733 412 1734
rect 438 1738 444 1739
rect 438 1734 439 1738
rect 443 1734 444 1738
rect 438 1733 444 1734
rect 470 1738 476 1739
rect 470 1734 471 1738
rect 475 1734 476 1738
rect 470 1733 476 1734
rect 502 1738 508 1739
rect 502 1734 503 1738
rect 507 1734 508 1738
rect 502 1733 508 1734
rect 534 1738 540 1739
rect 534 1734 535 1738
rect 539 1734 540 1738
rect 534 1733 540 1734
rect 566 1738 572 1739
rect 566 1734 567 1738
rect 571 1734 572 1738
rect 566 1733 572 1734
rect 598 1738 604 1739
rect 598 1734 599 1738
rect 603 1734 604 1738
rect 598 1733 604 1734
rect 630 1738 636 1739
rect 630 1734 631 1738
rect 635 1734 636 1738
rect 630 1733 636 1734
rect 662 1738 668 1739
rect 662 1734 663 1738
rect 667 1734 668 1738
rect 662 1733 668 1734
rect 694 1738 700 1739
rect 694 1734 695 1738
rect 699 1734 700 1738
rect 694 1733 700 1734
rect 726 1738 732 1739
rect 726 1734 727 1738
rect 731 1734 732 1738
rect 726 1733 732 1734
rect 758 1738 764 1739
rect 758 1734 759 1738
rect 763 1734 764 1738
rect 758 1733 764 1734
rect 790 1738 796 1739
rect 790 1734 791 1738
rect 795 1734 796 1738
rect 790 1733 796 1734
rect 822 1738 828 1739
rect 822 1734 823 1738
rect 827 1734 828 1738
rect 822 1733 828 1734
rect 854 1738 860 1739
rect 854 1734 855 1738
rect 859 1734 860 1738
rect 854 1733 860 1734
rect 886 1738 892 1739
rect 886 1734 887 1738
rect 891 1734 892 1738
rect 886 1733 892 1734
rect 918 1738 924 1739
rect 918 1734 919 1738
rect 923 1734 924 1738
rect 918 1733 924 1734
rect 950 1738 956 1739
rect 950 1734 951 1738
rect 955 1734 956 1738
rect 950 1733 956 1734
rect 982 1738 988 1739
rect 982 1734 983 1738
rect 987 1734 988 1738
rect 982 1733 988 1734
rect 1694 1736 1700 1737
rect 110 1731 116 1732
rect 112 1719 114 1731
rect 152 1719 154 1733
rect 184 1719 186 1733
rect 216 1719 218 1733
rect 248 1719 250 1733
rect 280 1719 282 1733
rect 312 1719 314 1733
rect 344 1719 346 1733
rect 376 1719 378 1733
rect 408 1719 410 1733
rect 440 1719 442 1733
rect 472 1719 474 1733
rect 504 1719 506 1733
rect 536 1719 538 1733
rect 568 1719 570 1733
rect 600 1719 602 1733
rect 632 1719 634 1733
rect 664 1719 666 1733
rect 696 1719 698 1733
rect 728 1719 730 1733
rect 760 1719 762 1733
rect 792 1719 794 1733
rect 824 1719 826 1733
rect 856 1719 858 1733
rect 888 1719 890 1733
rect 920 1719 922 1733
rect 952 1719 954 1733
rect 984 1719 986 1733
rect 1694 1732 1695 1736
rect 1699 1732 1700 1736
rect 1694 1731 1700 1732
rect 1696 1719 1698 1731
rect 111 1718 115 1719
rect 111 1713 115 1714
rect 151 1718 155 1719
rect 151 1713 155 1714
rect 183 1718 187 1719
rect 183 1713 187 1714
rect 191 1718 195 1719
rect 191 1713 195 1714
rect 215 1718 219 1719
rect 215 1713 219 1714
rect 247 1718 251 1719
rect 247 1713 251 1714
rect 279 1718 283 1719
rect 279 1713 283 1714
rect 311 1718 315 1719
rect 311 1713 315 1714
rect 319 1718 323 1719
rect 319 1713 323 1714
rect 343 1718 347 1719
rect 343 1713 347 1714
rect 375 1718 379 1719
rect 375 1713 379 1714
rect 407 1718 411 1719
rect 407 1713 411 1714
rect 415 1718 419 1719
rect 415 1713 419 1714
rect 439 1718 443 1719
rect 439 1713 443 1714
rect 471 1718 475 1719
rect 471 1713 475 1714
rect 503 1718 507 1719
rect 503 1713 507 1714
rect 527 1718 531 1719
rect 527 1713 531 1714
rect 535 1718 539 1719
rect 535 1713 539 1714
rect 567 1718 571 1719
rect 567 1713 571 1714
rect 599 1718 603 1719
rect 599 1713 603 1714
rect 631 1718 635 1719
rect 631 1713 635 1714
rect 655 1718 659 1719
rect 655 1713 659 1714
rect 663 1718 667 1719
rect 663 1713 667 1714
rect 695 1718 699 1719
rect 695 1713 699 1714
rect 727 1718 731 1719
rect 727 1713 731 1714
rect 759 1718 763 1719
rect 759 1713 763 1714
rect 791 1718 795 1719
rect 791 1713 795 1714
rect 823 1718 827 1719
rect 823 1713 827 1714
rect 855 1718 859 1719
rect 855 1713 859 1714
rect 887 1718 891 1719
rect 887 1713 891 1714
rect 919 1718 923 1719
rect 919 1713 923 1714
rect 951 1718 955 1719
rect 951 1713 955 1714
rect 983 1718 987 1719
rect 983 1713 987 1714
rect 1047 1718 1051 1719
rect 1047 1713 1051 1714
rect 1159 1718 1163 1719
rect 1159 1713 1163 1714
rect 1255 1718 1259 1719
rect 1255 1713 1259 1714
rect 1335 1718 1339 1719
rect 1335 1713 1339 1714
rect 1407 1718 1411 1719
rect 1407 1713 1411 1714
rect 1463 1718 1467 1719
rect 1463 1713 1467 1714
rect 1519 1718 1523 1719
rect 1519 1713 1523 1714
rect 1567 1718 1571 1719
rect 1567 1713 1571 1714
rect 1623 1718 1627 1719
rect 1623 1713 1627 1714
rect 1655 1718 1659 1719
rect 1655 1713 1659 1714
rect 1695 1718 1699 1719
rect 1695 1713 1699 1714
rect 112 1705 114 1713
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 192 1703 194 1713
rect 248 1703 250 1713
rect 320 1703 322 1713
rect 416 1703 418 1713
rect 528 1703 530 1713
rect 656 1703 658 1713
rect 792 1703 794 1713
rect 920 1703 922 1713
rect 1048 1703 1050 1713
rect 1160 1703 1162 1713
rect 1256 1703 1258 1713
rect 1336 1703 1338 1713
rect 1408 1703 1410 1713
rect 1464 1703 1466 1713
rect 1520 1703 1522 1713
rect 1568 1703 1570 1713
rect 1624 1703 1626 1713
rect 1656 1703 1658 1713
rect 1696 1705 1698 1713
rect 1694 1704 1700 1705
rect 110 1699 116 1700
rect 190 1702 196 1703
rect 190 1698 191 1702
rect 195 1698 196 1702
rect 190 1697 196 1698
rect 246 1702 252 1703
rect 246 1698 247 1702
rect 251 1698 252 1702
rect 246 1697 252 1698
rect 318 1702 324 1703
rect 318 1698 319 1702
rect 323 1698 324 1702
rect 318 1697 324 1698
rect 414 1702 420 1703
rect 414 1698 415 1702
rect 419 1698 420 1702
rect 414 1697 420 1698
rect 526 1702 532 1703
rect 526 1698 527 1702
rect 531 1698 532 1702
rect 526 1697 532 1698
rect 654 1702 660 1703
rect 654 1698 655 1702
rect 659 1698 660 1702
rect 654 1697 660 1698
rect 790 1702 796 1703
rect 790 1698 791 1702
rect 795 1698 796 1702
rect 790 1697 796 1698
rect 918 1702 924 1703
rect 918 1698 919 1702
rect 923 1698 924 1702
rect 918 1697 924 1698
rect 1046 1702 1052 1703
rect 1046 1698 1047 1702
rect 1051 1698 1052 1702
rect 1046 1697 1052 1698
rect 1158 1702 1164 1703
rect 1158 1698 1159 1702
rect 1163 1698 1164 1702
rect 1158 1697 1164 1698
rect 1254 1702 1260 1703
rect 1254 1698 1255 1702
rect 1259 1698 1260 1702
rect 1254 1697 1260 1698
rect 1334 1702 1340 1703
rect 1334 1698 1335 1702
rect 1339 1698 1340 1702
rect 1334 1697 1340 1698
rect 1406 1702 1412 1703
rect 1406 1698 1407 1702
rect 1411 1698 1412 1702
rect 1406 1697 1412 1698
rect 1462 1702 1468 1703
rect 1462 1698 1463 1702
rect 1467 1698 1468 1702
rect 1462 1697 1468 1698
rect 1518 1702 1524 1703
rect 1518 1698 1519 1702
rect 1523 1698 1524 1702
rect 1518 1697 1524 1698
rect 1566 1702 1572 1703
rect 1566 1698 1567 1702
rect 1571 1698 1572 1702
rect 1566 1697 1572 1698
rect 1622 1702 1628 1703
rect 1622 1698 1623 1702
rect 1627 1698 1628 1702
rect 1622 1697 1628 1698
rect 1654 1702 1660 1703
rect 1654 1698 1655 1702
rect 1659 1698 1660 1702
rect 1694 1700 1695 1704
rect 1699 1700 1700 1704
rect 1694 1699 1700 1700
rect 1654 1697 1660 1698
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 1694 1687 1700 1688
rect 110 1682 116 1683
rect 190 1685 196 1686
rect 112 1671 114 1682
rect 190 1681 191 1685
rect 195 1681 196 1685
rect 190 1680 196 1681
rect 246 1685 252 1686
rect 246 1681 247 1685
rect 251 1681 252 1685
rect 246 1680 252 1681
rect 318 1685 324 1686
rect 318 1681 319 1685
rect 323 1681 324 1685
rect 318 1680 324 1681
rect 414 1685 420 1686
rect 414 1681 415 1685
rect 419 1681 420 1685
rect 414 1680 420 1681
rect 526 1685 532 1686
rect 526 1681 527 1685
rect 531 1681 532 1685
rect 526 1680 532 1681
rect 654 1685 660 1686
rect 654 1681 655 1685
rect 659 1681 660 1685
rect 654 1680 660 1681
rect 790 1685 796 1686
rect 790 1681 791 1685
rect 795 1681 796 1685
rect 790 1680 796 1681
rect 918 1685 924 1686
rect 918 1681 919 1685
rect 923 1681 924 1685
rect 918 1680 924 1681
rect 1046 1685 1052 1686
rect 1046 1681 1047 1685
rect 1051 1681 1052 1685
rect 1046 1680 1052 1681
rect 1158 1685 1164 1686
rect 1158 1681 1159 1685
rect 1163 1681 1164 1685
rect 1158 1680 1164 1681
rect 1254 1685 1260 1686
rect 1254 1681 1255 1685
rect 1259 1681 1260 1685
rect 1254 1680 1260 1681
rect 1334 1685 1340 1686
rect 1334 1681 1335 1685
rect 1339 1681 1340 1685
rect 1334 1680 1340 1681
rect 1406 1685 1412 1686
rect 1406 1681 1407 1685
rect 1411 1681 1412 1685
rect 1406 1680 1412 1681
rect 1462 1685 1468 1686
rect 1462 1681 1463 1685
rect 1467 1681 1468 1685
rect 1462 1680 1468 1681
rect 1518 1685 1524 1686
rect 1518 1681 1519 1685
rect 1523 1681 1524 1685
rect 1518 1680 1524 1681
rect 1566 1685 1572 1686
rect 1566 1681 1567 1685
rect 1571 1681 1572 1685
rect 1566 1680 1572 1681
rect 1622 1685 1628 1686
rect 1622 1681 1623 1685
rect 1627 1681 1628 1685
rect 1622 1680 1628 1681
rect 1654 1685 1660 1686
rect 1654 1681 1655 1685
rect 1659 1681 1660 1685
rect 1694 1683 1695 1687
rect 1699 1683 1700 1687
rect 1694 1682 1700 1683
rect 1654 1680 1660 1681
rect 192 1671 194 1680
rect 248 1671 250 1680
rect 320 1671 322 1680
rect 416 1671 418 1680
rect 528 1671 530 1680
rect 656 1671 658 1680
rect 792 1671 794 1680
rect 920 1671 922 1680
rect 1048 1671 1050 1680
rect 1160 1671 1162 1680
rect 1256 1671 1258 1680
rect 1336 1671 1338 1680
rect 1408 1671 1410 1680
rect 1464 1671 1466 1680
rect 1520 1671 1522 1680
rect 1568 1671 1570 1680
rect 1624 1671 1626 1680
rect 1656 1671 1658 1680
rect 1696 1671 1698 1682
rect 111 1670 115 1671
rect 111 1665 115 1666
rect 135 1670 139 1671
rect 112 1662 114 1665
rect 135 1664 139 1666
rect 175 1670 179 1671
rect 175 1664 179 1666
rect 191 1670 195 1671
rect 191 1665 195 1666
rect 247 1670 251 1671
rect 247 1665 251 1666
rect 263 1670 267 1671
rect 263 1664 267 1666
rect 319 1670 323 1671
rect 319 1665 323 1666
rect 391 1670 395 1671
rect 391 1664 395 1666
rect 415 1670 419 1671
rect 415 1665 419 1666
rect 527 1670 531 1671
rect 527 1665 531 1666
rect 543 1670 547 1671
rect 543 1664 547 1666
rect 655 1670 659 1671
rect 655 1665 659 1666
rect 711 1670 715 1671
rect 711 1664 715 1666
rect 791 1670 795 1671
rect 791 1665 795 1666
rect 879 1670 883 1671
rect 879 1664 883 1666
rect 919 1670 923 1671
rect 919 1665 923 1666
rect 1039 1670 1043 1671
rect 1039 1664 1043 1666
rect 1047 1670 1051 1671
rect 1047 1665 1051 1666
rect 1159 1670 1163 1671
rect 1159 1665 1163 1666
rect 1183 1670 1187 1671
rect 1183 1664 1187 1666
rect 1255 1670 1259 1671
rect 1255 1665 1259 1666
rect 1319 1670 1323 1671
rect 1319 1664 1323 1666
rect 1335 1670 1339 1671
rect 1335 1665 1339 1666
rect 1407 1670 1411 1671
rect 1407 1665 1411 1666
rect 1439 1670 1443 1671
rect 1439 1664 1443 1666
rect 1463 1670 1467 1671
rect 1463 1665 1467 1666
rect 1519 1670 1523 1671
rect 1519 1665 1523 1666
rect 1559 1670 1563 1671
rect 1559 1664 1563 1666
rect 1567 1670 1571 1671
rect 1567 1665 1571 1666
rect 1623 1670 1627 1671
rect 1623 1665 1627 1666
rect 1655 1670 1659 1671
rect 1655 1664 1659 1666
rect 1695 1670 1699 1671
rect 1695 1665 1699 1666
rect 134 1663 140 1664
rect 110 1661 116 1662
rect 110 1657 111 1661
rect 115 1657 116 1661
rect 134 1659 135 1663
rect 139 1659 140 1663
rect 134 1658 140 1659
rect 174 1663 180 1664
rect 174 1659 175 1663
rect 179 1659 180 1663
rect 174 1658 180 1659
rect 262 1663 268 1664
rect 262 1659 263 1663
rect 267 1659 268 1663
rect 262 1658 268 1659
rect 390 1663 396 1664
rect 390 1659 391 1663
rect 395 1659 396 1663
rect 390 1658 396 1659
rect 542 1663 548 1664
rect 542 1659 543 1663
rect 547 1659 548 1663
rect 542 1658 548 1659
rect 710 1663 716 1664
rect 710 1659 711 1663
rect 715 1659 716 1663
rect 710 1658 716 1659
rect 878 1663 884 1664
rect 878 1659 879 1663
rect 883 1659 884 1663
rect 878 1658 884 1659
rect 1038 1663 1044 1664
rect 1038 1659 1039 1663
rect 1043 1659 1044 1663
rect 1038 1658 1044 1659
rect 1182 1663 1188 1664
rect 1182 1659 1183 1663
rect 1187 1659 1188 1663
rect 1182 1658 1188 1659
rect 1318 1663 1324 1664
rect 1318 1659 1319 1663
rect 1323 1659 1324 1663
rect 1318 1658 1324 1659
rect 1438 1663 1444 1664
rect 1438 1659 1439 1663
rect 1443 1659 1444 1663
rect 1438 1658 1444 1659
rect 1558 1663 1564 1664
rect 1558 1659 1559 1663
rect 1563 1659 1564 1663
rect 1558 1658 1564 1659
rect 1654 1663 1660 1664
rect 1654 1659 1655 1663
rect 1659 1659 1660 1663
rect 1696 1662 1698 1665
rect 1654 1658 1660 1659
rect 1694 1661 1700 1662
rect 110 1656 116 1657
rect 1694 1657 1695 1661
rect 1699 1657 1700 1661
rect 1694 1656 1700 1657
rect 134 1646 140 1647
rect 110 1644 116 1645
rect 110 1640 111 1644
rect 115 1640 116 1644
rect 134 1642 135 1646
rect 139 1642 140 1646
rect 134 1641 140 1642
rect 174 1646 180 1647
rect 174 1642 175 1646
rect 179 1642 180 1646
rect 174 1641 180 1642
rect 262 1646 268 1647
rect 262 1642 263 1646
rect 267 1642 268 1646
rect 262 1641 268 1642
rect 390 1646 396 1647
rect 390 1642 391 1646
rect 395 1642 396 1646
rect 390 1641 396 1642
rect 542 1646 548 1647
rect 542 1642 543 1646
rect 547 1642 548 1646
rect 542 1641 548 1642
rect 710 1646 716 1647
rect 710 1642 711 1646
rect 715 1642 716 1646
rect 710 1641 716 1642
rect 878 1646 884 1647
rect 878 1642 879 1646
rect 883 1642 884 1646
rect 878 1641 884 1642
rect 1038 1646 1044 1647
rect 1038 1642 1039 1646
rect 1043 1642 1044 1646
rect 1038 1641 1044 1642
rect 1182 1646 1188 1647
rect 1182 1642 1183 1646
rect 1187 1642 1188 1646
rect 1182 1641 1188 1642
rect 1318 1646 1324 1647
rect 1318 1642 1319 1646
rect 1323 1642 1324 1646
rect 1318 1641 1324 1642
rect 1438 1646 1444 1647
rect 1438 1642 1439 1646
rect 1443 1642 1444 1646
rect 1438 1641 1444 1642
rect 1558 1646 1564 1647
rect 1558 1642 1559 1646
rect 1563 1642 1564 1646
rect 1558 1641 1564 1642
rect 1654 1646 1660 1647
rect 1654 1642 1655 1646
rect 1659 1642 1660 1646
rect 1654 1641 1660 1642
rect 1694 1644 1700 1645
rect 110 1639 116 1640
rect 112 1623 114 1639
rect 136 1623 138 1641
rect 176 1623 178 1641
rect 264 1623 266 1641
rect 392 1623 394 1641
rect 544 1623 546 1641
rect 712 1623 714 1641
rect 880 1623 882 1641
rect 1040 1623 1042 1641
rect 1184 1623 1186 1641
rect 1320 1623 1322 1641
rect 1440 1623 1442 1641
rect 1560 1623 1562 1641
rect 1656 1623 1658 1641
rect 1694 1640 1695 1644
rect 1699 1640 1700 1644
rect 1694 1639 1700 1640
rect 1696 1623 1698 1639
rect 111 1622 115 1623
rect 111 1617 115 1618
rect 135 1622 139 1623
rect 135 1617 139 1618
rect 167 1622 171 1623
rect 167 1617 171 1618
rect 175 1622 179 1623
rect 175 1617 179 1618
rect 199 1622 203 1623
rect 199 1617 203 1618
rect 247 1622 251 1623
rect 247 1617 251 1618
rect 263 1622 267 1623
rect 263 1617 267 1618
rect 327 1622 331 1623
rect 327 1617 331 1618
rect 391 1622 395 1623
rect 391 1617 395 1618
rect 439 1622 443 1623
rect 439 1617 443 1618
rect 543 1622 547 1623
rect 543 1617 547 1618
rect 567 1622 571 1623
rect 567 1617 571 1618
rect 711 1622 715 1623
rect 711 1617 715 1618
rect 855 1622 859 1623
rect 855 1617 859 1618
rect 879 1622 883 1623
rect 879 1617 883 1618
rect 999 1622 1003 1623
rect 999 1617 1003 1618
rect 1039 1622 1043 1623
rect 1039 1617 1043 1618
rect 1127 1622 1131 1623
rect 1127 1617 1131 1618
rect 1183 1622 1187 1623
rect 1183 1617 1187 1618
rect 1247 1622 1251 1623
rect 1247 1617 1251 1618
rect 1319 1622 1323 1623
rect 1319 1617 1323 1618
rect 1359 1622 1363 1623
rect 1359 1617 1363 1618
rect 1439 1622 1443 1623
rect 1439 1617 1443 1618
rect 1463 1622 1467 1623
rect 1463 1617 1467 1618
rect 1559 1622 1563 1623
rect 1559 1617 1563 1618
rect 1567 1622 1571 1623
rect 1567 1617 1571 1618
rect 1655 1622 1659 1623
rect 1655 1617 1659 1618
rect 1695 1622 1699 1623
rect 1695 1617 1699 1618
rect 112 1609 114 1617
rect 110 1608 116 1609
rect 110 1604 111 1608
rect 115 1604 116 1608
rect 136 1607 138 1617
rect 168 1607 170 1617
rect 200 1607 202 1617
rect 248 1607 250 1617
rect 328 1607 330 1617
rect 440 1607 442 1617
rect 568 1607 570 1617
rect 712 1607 714 1617
rect 856 1607 858 1617
rect 1000 1607 1002 1617
rect 1128 1607 1130 1617
rect 1248 1607 1250 1617
rect 1360 1607 1362 1617
rect 1464 1607 1466 1617
rect 1568 1607 1570 1617
rect 1656 1607 1658 1617
rect 1696 1609 1698 1617
rect 1694 1608 1700 1609
rect 110 1603 116 1604
rect 134 1606 140 1607
rect 134 1602 135 1606
rect 139 1602 140 1606
rect 134 1601 140 1602
rect 166 1606 172 1607
rect 166 1602 167 1606
rect 171 1602 172 1606
rect 166 1601 172 1602
rect 198 1606 204 1607
rect 198 1602 199 1606
rect 203 1602 204 1606
rect 198 1601 204 1602
rect 246 1606 252 1607
rect 246 1602 247 1606
rect 251 1602 252 1606
rect 246 1601 252 1602
rect 326 1606 332 1607
rect 326 1602 327 1606
rect 331 1602 332 1606
rect 326 1601 332 1602
rect 438 1606 444 1607
rect 438 1602 439 1606
rect 443 1602 444 1606
rect 438 1601 444 1602
rect 566 1606 572 1607
rect 566 1602 567 1606
rect 571 1602 572 1606
rect 566 1601 572 1602
rect 710 1606 716 1607
rect 710 1602 711 1606
rect 715 1602 716 1606
rect 710 1601 716 1602
rect 854 1606 860 1607
rect 854 1602 855 1606
rect 859 1602 860 1606
rect 854 1601 860 1602
rect 998 1606 1004 1607
rect 998 1602 999 1606
rect 1003 1602 1004 1606
rect 998 1601 1004 1602
rect 1126 1606 1132 1607
rect 1126 1602 1127 1606
rect 1131 1602 1132 1606
rect 1126 1601 1132 1602
rect 1246 1606 1252 1607
rect 1246 1602 1247 1606
rect 1251 1602 1252 1606
rect 1246 1601 1252 1602
rect 1358 1606 1364 1607
rect 1358 1602 1359 1606
rect 1363 1602 1364 1606
rect 1358 1601 1364 1602
rect 1462 1606 1468 1607
rect 1462 1602 1463 1606
rect 1467 1602 1468 1606
rect 1462 1601 1468 1602
rect 1566 1606 1572 1607
rect 1566 1602 1567 1606
rect 1571 1602 1572 1606
rect 1566 1601 1572 1602
rect 1654 1606 1660 1607
rect 1654 1602 1655 1606
rect 1659 1602 1660 1606
rect 1694 1604 1695 1608
rect 1699 1604 1700 1608
rect 1694 1603 1700 1604
rect 1654 1601 1660 1602
rect 110 1591 116 1592
rect 110 1587 111 1591
rect 115 1587 116 1591
rect 1694 1591 1700 1592
rect 110 1586 116 1587
rect 134 1589 140 1590
rect 112 1583 114 1586
rect 134 1585 135 1589
rect 139 1585 140 1589
rect 134 1584 140 1585
rect 166 1589 172 1590
rect 166 1585 167 1589
rect 171 1585 172 1589
rect 166 1584 172 1585
rect 198 1589 204 1590
rect 198 1585 199 1589
rect 203 1585 204 1589
rect 198 1584 204 1585
rect 246 1589 252 1590
rect 246 1585 247 1589
rect 251 1585 252 1589
rect 246 1584 252 1585
rect 326 1589 332 1590
rect 326 1585 327 1589
rect 331 1585 332 1589
rect 326 1584 332 1585
rect 438 1589 444 1590
rect 438 1585 439 1589
rect 443 1585 444 1589
rect 438 1584 444 1585
rect 566 1589 572 1590
rect 566 1585 567 1589
rect 571 1585 572 1589
rect 566 1584 572 1585
rect 710 1589 716 1590
rect 710 1585 711 1589
rect 715 1585 716 1589
rect 710 1584 716 1585
rect 854 1589 860 1590
rect 854 1585 855 1589
rect 859 1585 860 1589
rect 854 1584 860 1585
rect 998 1589 1004 1590
rect 998 1585 999 1589
rect 1003 1585 1004 1589
rect 998 1584 1004 1585
rect 1126 1589 1132 1590
rect 1126 1585 1127 1589
rect 1131 1585 1132 1589
rect 1126 1584 1132 1585
rect 1246 1589 1252 1590
rect 1246 1585 1247 1589
rect 1251 1585 1252 1589
rect 1246 1584 1252 1585
rect 1358 1589 1364 1590
rect 1358 1585 1359 1589
rect 1363 1585 1364 1589
rect 1358 1584 1364 1585
rect 1462 1589 1468 1590
rect 1462 1585 1463 1589
rect 1467 1585 1468 1589
rect 1462 1584 1468 1585
rect 1566 1589 1572 1590
rect 1566 1585 1567 1589
rect 1571 1585 1572 1589
rect 1566 1584 1572 1585
rect 1654 1589 1660 1590
rect 1654 1585 1655 1589
rect 1659 1585 1660 1589
rect 1694 1587 1695 1591
rect 1699 1587 1700 1591
rect 1694 1586 1700 1587
rect 1654 1584 1660 1585
rect 111 1582 115 1583
rect 111 1577 115 1578
rect 135 1582 139 1584
rect 112 1574 114 1577
rect 135 1576 139 1578
rect 167 1582 171 1584
rect 167 1576 171 1578
rect 199 1582 203 1584
rect 199 1577 203 1578
rect 231 1582 235 1583
rect 231 1576 235 1578
rect 247 1582 251 1584
rect 247 1577 251 1578
rect 287 1582 291 1583
rect 287 1576 291 1578
rect 327 1582 331 1584
rect 327 1577 331 1578
rect 343 1582 347 1583
rect 343 1576 347 1578
rect 399 1582 403 1583
rect 399 1576 403 1578
rect 439 1582 443 1584
rect 439 1577 443 1578
rect 455 1582 459 1583
rect 455 1576 459 1578
rect 511 1582 515 1583
rect 511 1576 515 1578
rect 567 1582 571 1584
rect 567 1577 571 1578
rect 575 1582 579 1583
rect 575 1576 579 1578
rect 655 1582 659 1583
rect 655 1576 659 1578
rect 711 1582 715 1584
rect 711 1577 715 1578
rect 751 1582 755 1583
rect 751 1576 755 1578
rect 855 1582 859 1584
rect 855 1576 859 1578
rect 959 1582 963 1583
rect 959 1576 963 1578
rect 999 1582 1003 1584
rect 999 1577 1003 1578
rect 1063 1582 1067 1583
rect 1063 1576 1067 1578
rect 1127 1582 1131 1584
rect 1127 1577 1131 1578
rect 1159 1582 1163 1583
rect 1159 1576 1163 1578
rect 1247 1582 1251 1584
rect 1247 1576 1251 1578
rect 1327 1582 1331 1583
rect 1327 1576 1331 1578
rect 1359 1582 1363 1584
rect 1359 1577 1363 1578
rect 1399 1582 1403 1583
rect 1399 1576 1403 1578
rect 1463 1582 1467 1584
rect 1463 1577 1467 1578
rect 1471 1582 1475 1583
rect 1471 1576 1475 1578
rect 1535 1582 1539 1583
rect 1535 1576 1539 1578
rect 1567 1582 1571 1584
rect 1567 1577 1571 1578
rect 1607 1582 1611 1583
rect 1607 1576 1611 1578
rect 1655 1582 1659 1584
rect 1696 1583 1698 1586
rect 1655 1576 1659 1578
rect 1695 1582 1699 1583
rect 1695 1577 1699 1578
rect 134 1575 140 1576
rect 110 1573 116 1574
rect 110 1569 111 1573
rect 115 1569 116 1573
rect 134 1571 135 1575
rect 139 1571 140 1575
rect 134 1570 140 1571
rect 166 1575 172 1576
rect 166 1571 167 1575
rect 171 1571 172 1575
rect 166 1570 172 1571
rect 230 1575 236 1576
rect 230 1571 231 1575
rect 235 1571 236 1575
rect 230 1570 236 1571
rect 286 1575 292 1576
rect 286 1571 287 1575
rect 291 1571 292 1575
rect 286 1570 292 1571
rect 342 1575 348 1576
rect 342 1571 343 1575
rect 347 1571 348 1575
rect 342 1570 348 1571
rect 398 1575 404 1576
rect 398 1571 399 1575
rect 403 1571 404 1575
rect 398 1570 404 1571
rect 454 1575 460 1576
rect 454 1571 455 1575
rect 459 1571 460 1575
rect 454 1570 460 1571
rect 510 1575 516 1576
rect 510 1571 511 1575
rect 515 1571 516 1575
rect 510 1570 516 1571
rect 574 1575 580 1576
rect 574 1571 575 1575
rect 579 1571 580 1575
rect 574 1570 580 1571
rect 654 1575 660 1576
rect 654 1571 655 1575
rect 659 1571 660 1575
rect 654 1570 660 1571
rect 750 1575 756 1576
rect 750 1571 751 1575
rect 755 1571 756 1575
rect 750 1570 756 1571
rect 854 1575 860 1576
rect 854 1571 855 1575
rect 859 1571 860 1575
rect 854 1570 860 1571
rect 958 1575 964 1576
rect 958 1571 959 1575
rect 963 1571 964 1575
rect 958 1570 964 1571
rect 1062 1575 1068 1576
rect 1062 1571 1063 1575
rect 1067 1571 1068 1575
rect 1062 1570 1068 1571
rect 1158 1575 1164 1576
rect 1158 1571 1159 1575
rect 1163 1571 1164 1575
rect 1158 1570 1164 1571
rect 1246 1575 1252 1576
rect 1246 1571 1247 1575
rect 1251 1571 1252 1575
rect 1246 1570 1252 1571
rect 1326 1575 1332 1576
rect 1326 1571 1327 1575
rect 1331 1571 1332 1575
rect 1326 1570 1332 1571
rect 1398 1575 1404 1576
rect 1398 1571 1399 1575
rect 1403 1571 1404 1575
rect 1398 1570 1404 1571
rect 1470 1575 1476 1576
rect 1470 1571 1471 1575
rect 1475 1571 1476 1575
rect 1470 1570 1476 1571
rect 1534 1575 1540 1576
rect 1534 1571 1535 1575
rect 1539 1571 1540 1575
rect 1534 1570 1540 1571
rect 1606 1575 1612 1576
rect 1606 1571 1607 1575
rect 1611 1571 1612 1575
rect 1606 1570 1612 1571
rect 1654 1575 1660 1576
rect 1654 1571 1655 1575
rect 1659 1571 1660 1575
rect 1696 1574 1698 1577
rect 1654 1570 1660 1571
rect 1694 1573 1700 1574
rect 110 1568 116 1569
rect 1694 1569 1695 1573
rect 1699 1569 1700 1573
rect 1694 1568 1700 1569
rect 134 1558 140 1559
rect 110 1556 116 1557
rect 110 1552 111 1556
rect 115 1552 116 1556
rect 134 1554 135 1558
rect 139 1554 140 1558
rect 134 1553 140 1554
rect 166 1558 172 1559
rect 166 1554 167 1558
rect 171 1554 172 1558
rect 166 1553 172 1554
rect 230 1558 236 1559
rect 230 1554 231 1558
rect 235 1554 236 1558
rect 230 1553 236 1554
rect 286 1558 292 1559
rect 286 1554 287 1558
rect 291 1554 292 1558
rect 286 1553 292 1554
rect 342 1558 348 1559
rect 342 1554 343 1558
rect 347 1554 348 1558
rect 342 1553 348 1554
rect 398 1558 404 1559
rect 398 1554 399 1558
rect 403 1554 404 1558
rect 398 1553 404 1554
rect 454 1558 460 1559
rect 454 1554 455 1558
rect 459 1554 460 1558
rect 454 1553 460 1554
rect 510 1558 516 1559
rect 510 1554 511 1558
rect 515 1554 516 1558
rect 510 1553 516 1554
rect 574 1558 580 1559
rect 574 1554 575 1558
rect 579 1554 580 1558
rect 574 1553 580 1554
rect 654 1558 660 1559
rect 654 1554 655 1558
rect 659 1554 660 1558
rect 654 1553 660 1554
rect 750 1558 756 1559
rect 750 1554 751 1558
rect 755 1554 756 1558
rect 750 1553 756 1554
rect 854 1558 860 1559
rect 854 1554 855 1558
rect 859 1554 860 1558
rect 854 1553 860 1554
rect 958 1558 964 1559
rect 958 1554 959 1558
rect 963 1554 964 1558
rect 958 1553 964 1554
rect 1062 1558 1068 1559
rect 1062 1554 1063 1558
rect 1067 1554 1068 1558
rect 1062 1553 1068 1554
rect 1158 1558 1164 1559
rect 1158 1554 1159 1558
rect 1163 1554 1164 1558
rect 1158 1553 1164 1554
rect 1246 1558 1252 1559
rect 1246 1554 1247 1558
rect 1251 1554 1252 1558
rect 1246 1553 1252 1554
rect 1326 1558 1332 1559
rect 1326 1554 1327 1558
rect 1331 1554 1332 1558
rect 1326 1553 1332 1554
rect 1398 1558 1404 1559
rect 1398 1554 1399 1558
rect 1403 1554 1404 1558
rect 1398 1553 1404 1554
rect 1470 1558 1476 1559
rect 1470 1554 1471 1558
rect 1475 1554 1476 1558
rect 1470 1553 1476 1554
rect 1534 1558 1540 1559
rect 1534 1554 1535 1558
rect 1539 1554 1540 1558
rect 1534 1553 1540 1554
rect 1606 1558 1612 1559
rect 1606 1554 1607 1558
rect 1611 1554 1612 1558
rect 1606 1553 1612 1554
rect 1654 1558 1660 1559
rect 1654 1554 1655 1558
rect 1659 1554 1660 1558
rect 1654 1553 1660 1554
rect 1694 1556 1700 1557
rect 110 1551 116 1552
rect 112 1543 114 1551
rect 136 1543 138 1553
rect 168 1543 170 1553
rect 232 1543 234 1553
rect 288 1543 290 1553
rect 344 1543 346 1553
rect 400 1543 402 1553
rect 456 1543 458 1553
rect 512 1543 514 1553
rect 576 1543 578 1553
rect 656 1543 658 1553
rect 752 1543 754 1553
rect 856 1543 858 1553
rect 960 1543 962 1553
rect 1064 1543 1066 1553
rect 1160 1543 1162 1553
rect 1248 1543 1250 1553
rect 1328 1543 1330 1553
rect 1400 1543 1402 1553
rect 1472 1543 1474 1553
rect 1536 1543 1538 1553
rect 1608 1543 1610 1553
rect 1656 1543 1658 1553
rect 1694 1552 1695 1556
rect 1699 1552 1700 1556
rect 1694 1551 1700 1552
rect 1696 1543 1698 1551
rect 111 1542 115 1543
rect 111 1537 115 1538
rect 135 1542 139 1543
rect 135 1537 139 1538
rect 167 1542 171 1543
rect 167 1537 171 1538
rect 175 1542 179 1543
rect 175 1537 179 1538
rect 223 1542 227 1543
rect 223 1537 227 1538
rect 231 1542 235 1543
rect 231 1537 235 1538
rect 279 1542 283 1543
rect 279 1537 283 1538
rect 287 1542 291 1543
rect 287 1537 291 1538
rect 335 1542 339 1543
rect 335 1537 339 1538
rect 343 1542 347 1543
rect 343 1537 347 1538
rect 399 1542 403 1543
rect 399 1537 403 1538
rect 455 1542 459 1543
rect 455 1537 459 1538
rect 463 1542 467 1543
rect 463 1537 467 1538
rect 511 1542 515 1543
rect 511 1537 515 1538
rect 535 1542 539 1543
rect 535 1537 539 1538
rect 575 1542 579 1543
rect 575 1537 579 1538
rect 607 1542 611 1543
rect 607 1537 611 1538
rect 655 1542 659 1543
rect 655 1537 659 1538
rect 687 1542 691 1543
rect 687 1537 691 1538
rect 751 1542 755 1543
rect 751 1537 755 1538
rect 775 1542 779 1543
rect 775 1537 779 1538
rect 855 1542 859 1543
rect 855 1537 859 1538
rect 871 1542 875 1543
rect 871 1537 875 1538
rect 959 1542 963 1543
rect 959 1537 963 1538
rect 975 1542 979 1543
rect 975 1537 979 1538
rect 1063 1542 1067 1543
rect 1063 1537 1067 1538
rect 1079 1542 1083 1543
rect 1079 1537 1083 1538
rect 1159 1542 1163 1543
rect 1159 1537 1163 1538
rect 1175 1542 1179 1543
rect 1175 1537 1179 1538
rect 1247 1542 1251 1543
rect 1247 1537 1251 1538
rect 1271 1542 1275 1543
rect 1271 1537 1275 1538
rect 1327 1542 1331 1543
rect 1327 1537 1331 1538
rect 1359 1542 1363 1543
rect 1359 1537 1363 1538
rect 1399 1542 1403 1543
rect 1399 1537 1403 1538
rect 1439 1542 1443 1543
rect 1439 1537 1443 1538
rect 1471 1542 1475 1543
rect 1471 1537 1475 1538
rect 1519 1542 1523 1543
rect 1519 1537 1523 1538
rect 1535 1542 1539 1543
rect 1535 1537 1539 1538
rect 1599 1542 1603 1543
rect 1599 1537 1603 1538
rect 1607 1542 1611 1543
rect 1607 1537 1611 1538
rect 1655 1542 1659 1543
rect 1655 1537 1659 1538
rect 1695 1542 1699 1543
rect 1695 1537 1699 1538
rect 112 1529 114 1537
rect 110 1528 116 1529
rect 110 1524 111 1528
rect 115 1524 116 1528
rect 136 1527 138 1537
rect 176 1527 178 1537
rect 224 1527 226 1537
rect 280 1527 282 1537
rect 336 1527 338 1537
rect 400 1527 402 1537
rect 464 1527 466 1537
rect 536 1527 538 1537
rect 608 1527 610 1537
rect 688 1527 690 1537
rect 776 1527 778 1537
rect 872 1527 874 1537
rect 976 1527 978 1537
rect 1080 1527 1082 1537
rect 1176 1527 1178 1537
rect 1272 1527 1274 1537
rect 1360 1527 1362 1537
rect 1440 1527 1442 1537
rect 1520 1527 1522 1537
rect 1600 1527 1602 1537
rect 1656 1527 1658 1537
rect 1696 1529 1698 1537
rect 1694 1528 1700 1529
rect 110 1523 116 1524
rect 134 1526 140 1527
rect 134 1522 135 1526
rect 139 1522 140 1526
rect 134 1521 140 1522
rect 174 1526 180 1527
rect 174 1522 175 1526
rect 179 1522 180 1526
rect 174 1521 180 1522
rect 222 1526 228 1527
rect 222 1522 223 1526
rect 227 1522 228 1526
rect 222 1521 228 1522
rect 278 1526 284 1527
rect 278 1522 279 1526
rect 283 1522 284 1526
rect 278 1521 284 1522
rect 334 1526 340 1527
rect 334 1522 335 1526
rect 339 1522 340 1526
rect 334 1521 340 1522
rect 398 1526 404 1527
rect 398 1522 399 1526
rect 403 1522 404 1526
rect 398 1521 404 1522
rect 462 1526 468 1527
rect 462 1522 463 1526
rect 467 1522 468 1526
rect 462 1521 468 1522
rect 534 1526 540 1527
rect 534 1522 535 1526
rect 539 1522 540 1526
rect 534 1521 540 1522
rect 606 1526 612 1527
rect 606 1522 607 1526
rect 611 1522 612 1526
rect 606 1521 612 1522
rect 686 1526 692 1527
rect 686 1522 687 1526
rect 691 1522 692 1526
rect 686 1521 692 1522
rect 774 1526 780 1527
rect 774 1522 775 1526
rect 779 1522 780 1526
rect 774 1521 780 1522
rect 870 1526 876 1527
rect 870 1522 871 1526
rect 875 1522 876 1526
rect 870 1521 876 1522
rect 974 1526 980 1527
rect 974 1522 975 1526
rect 979 1522 980 1526
rect 974 1521 980 1522
rect 1078 1526 1084 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1174 1526 1180 1527
rect 1174 1522 1175 1526
rect 1179 1522 1180 1526
rect 1174 1521 1180 1522
rect 1270 1526 1276 1527
rect 1270 1522 1271 1526
rect 1275 1522 1276 1526
rect 1270 1521 1276 1522
rect 1358 1526 1364 1527
rect 1358 1522 1359 1526
rect 1363 1522 1364 1526
rect 1358 1521 1364 1522
rect 1438 1526 1444 1527
rect 1438 1522 1439 1526
rect 1443 1522 1444 1526
rect 1438 1521 1444 1522
rect 1518 1526 1524 1527
rect 1518 1522 1519 1526
rect 1523 1522 1524 1526
rect 1518 1521 1524 1522
rect 1598 1526 1604 1527
rect 1598 1522 1599 1526
rect 1603 1522 1604 1526
rect 1598 1521 1604 1522
rect 1654 1526 1660 1527
rect 1654 1522 1655 1526
rect 1659 1522 1660 1526
rect 1694 1524 1695 1528
rect 1699 1524 1700 1528
rect 1694 1523 1700 1524
rect 1654 1521 1660 1522
rect 110 1511 116 1512
rect 110 1507 111 1511
rect 115 1507 116 1511
rect 1694 1511 1700 1512
rect 110 1506 116 1507
rect 134 1509 140 1510
rect 112 1499 114 1506
rect 134 1505 135 1509
rect 139 1505 140 1509
rect 134 1504 140 1505
rect 174 1509 180 1510
rect 174 1505 175 1509
rect 179 1505 180 1509
rect 174 1504 180 1505
rect 222 1509 228 1510
rect 222 1505 223 1509
rect 227 1505 228 1509
rect 222 1504 228 1505
rect 278 1509 284 1510
rect 278 1505 279 1509
rect 283 1505 284 1509
rect 278 1504 284 1505
rect 334 1509 340 1510
rect 334 1505 335 1509
rect 339 1505 340 1509
rect 334 1504 340 1505
rect 398 1509 404 1510
rect 398 1505 399 1509
rect 403 1505 404 1509
rect 398 1504 404 1505
rect 462 1509 468 1510
rect 462 1505 463 1509
rect 467 1505 468 1509
rect 462 1504 468 1505
rect 534 1509 540 1510
rect 534 1505 535 1509
rect 539 1505 540 1509
rect 534 1504 540 1505
rect 606 1509 612 1510
rect 606 1505 607 1509
rect 611 1505 612 1509
rect 606 1504 612 1505
rect 686 1509 692 1510
rect 686 1505 687 1509
rect 691 1505 692 1509
rect 686 1504 692 1505
rect 774 1509 780 1510
rect 774 1505 775 1509
rect 779 1505 780 1509
rect 774 1504 780 1505
rect 870 1509 876 1510
rect 870 1505 871 1509
rect 875 1505 876 1509
rect 870 1504 876 1505
rect 974 1509 980 1510
rect 974 1505 975 1509
rect 979 1505 980 1509
rect 974 1504 980 1505
rect 1078 1509 1084 1510
rect 1078 1505 1079 1509
rect 1083 1505 1084 1509
rect 1078 1504 1084 1505
rect 1174 1509 1180 1510
rect 1174 1505 1175 1509
rect 1179 1505 1180 1509
rect 1174 1504 1180 1505
rect 1270 1509 1276 1510
rect 1270 1505 1271 1509
rect 1275 1505 1276 1509
rect 1270 1504 1276 1505
rect 1358 1509 1364 1510
rect 1358 1505 1359 1509
rect 1363 1505 1364 1509
rect 1358 1504 1364 1505
rect 1438 1509 1444 1510
rect 1438 1505 1439 1509
rect 1443 1505 1444 1509
rect 1438 1504 1444 1505
rect 1518 1509 1524 1510
rect 1518 1505 1519 1509
rect 1523 1505 1524 1509
rect 1518 1504 1524 1505
rect 1598 1509 1604 1510
rect 1598 1505 1599 1509
rect 1603 1505 1604 1509
rect 1598 1504 1604 1505
rect 1654 1509 1660 1510
rect 1654 1505 1655 1509
rect 1659 1505 1660 1509
rect 1694 1507 1695 1511
rect 1699 1507 1700 1511
rect 1694 1506 1700 1507
rect 1654 1504 1660 1505
rect 136 1499 138 1504
rect 176 1499 178 1504
rect 224 1499 226 1504
rect 280 1499 282 1504
rect 336 1499 338 1504
rect 400 1499 402 1504
rect 464 1499 466 1504
rect 536 1499 538 1504
rect 608 1499 610 1504
rect 688 1499 690 1504
rect 776 1499 778 1504
rect 872 1499 874 1504
rect 976 1499 978 1504
rect 1080 1499 1082 1504
rect 1176 1499 1178 1504
rect 1272 1499 1274 1504
rect 1360 1499 1362 1504
rect 1440 1499 1442 1504
rect 1520 1499 1522 1504
rect 1600 1499 1602 1504
rect 1656 1499 1658 1504
rect 1696 1499 1698 1506
rect 111 1498 115 1499
rect 111 1493 115 1494
rect 135 1498 139 1499
rect 135 1493 139 1494
rect 175 1498 179 1499
rect 175 1493 179 1494
rect 207 1498 211 1499
rect 207 1493 211 1494
rect 223 1498 227 1499
rect 223 1493 227 1494
rect 239 1498 243 1499
rect 239 1493 243 1494
rect 271 1498 275 1499
rect 271 1493 275 1494
rect 279 1498 283 1499
rect 279 1493 283 1494
rect 303 1498 307 1499
rect 303 1493 307 1494
rect 335 1498 339 1499
rect 335 1493 339 1494
rect 367 1498 371 1499
rect 367 1493 371 1494
rect 399 1498 403 1499
rect 399 1493 403 1494
rect 431 1498 435 1499
rect 431 1493 435 1494
rect 463 1498 467 1499
rect 463 1493 467 1494
rect 495 1498 499 1499
rect 495 1493 499 1494
rect 527 1498 531 1499
rect 527 1493 531 1494
rect 535 1498 539 1499
rect 535 1493 539 1494
rect 559 1498 563 1499
rect 559 1493 563 1494
rect 591 1498 595 1499
rect 591 1493 595 1494
rect 607 1498 611 1499
rect 607 1493 611 1494
rect 623 1498 627 1499
rect 623 1493 627 1494
rect 663 1498 667 1499
rect 663 1493 667 1494
rect 687 1498 691 1499
rect 687 1493 691 1494
rect 703 1498 707 1499
rect 703 1493 707 1494
rect 743 1498 747 1499
rect 743 1493 747 1494
rect 775 1498 779 1499
rect 775 1493 779 1494
rect 807 1498 811 1499
rect 807 1493 811 1494
rect 871 1498 875 1499
rect 871 1493 875 1494
rect 895 1498 899 1499
rect 895 1493 899 1494
rect 935 1498 939 1499
rect 935 1493 939 1494
rect 975 1498 979 1499
rect 975 1493 979 1494
rect 1023 1498 1027 1499
rect 1023 1493 1027 1494
rect 1079 1498 1083 1499
rect 1079 1493 1083 1494
rect 1111 1498 1115 1499
rect 1111 1493 1115 1494
rect 1167 1498 1171 1499
rect 1167 1493 1171 1494
rect 1175 1498 1179 1499
rect 1175 1493 1179 1494
rect 1199 1498 1203 1499
rect 1199 1493 1203 1494
rect 1239 1498 1243 1499
rect 1239 1493 1243 1494
rect 1271 1498 1275 1499
rect 1271 1493 1275 1494
rect 1279 1498 1283 1499
rect 1279 1493 1283 1494
rect 1319 1498 1323 1499
rect 1319 1493 1323 1494
rect 1359 1498 1363 1499
rect 1359 1493 1363 1494
rect 1399 1498 1403 1499
rect 1399 1493 1403 1494
rect 1439 1498 1443 1499
rect 1439 1493 1443 1494
rect 1479 1498 1483 1499
rect 1479 1493 1483 1494
rect 1519 1498 1523 1499
rect 1519 1493 1523 1494
rect 1559 1498 1563 1499
rect 1559 1493 1563 1494
rect 1591 1498 1595 1499
rect 1591 1493 1595 1494
rect 1599 1498 1603 1499
rect 1599 1493 1603 1494
rect 1623 1498 1627 1499
rect 1623 1493 1627 1494
rect 1655 1498 1659 1499
rect 1655 1493 1659 1494
rect 1695 1498 1699 1499
rect 1695 1493 1699 1494
rect 112 1474 114 1493
rect 176 1476 178 1493
rect 208 1476 210 1493
rect 240 1476 242 1493
rect 272 1476 274 1493
rect 304 1476 306 1493
rect 336 1476 338 1493
rect 368 1476 370 1493
rect 400 1476 402 1493
rect 432 1476 434 1493
rect 464 1476 466 1493
rect 496 1476 498 1493
rect 528 1476 530 1493
rect 560 1476 562 1493
rect 592 1476 594 1493
rect 624 1476 626 1493
rect 664 1476 666 1493
rect 704 1476 706 1493
rect 744 1476 746 1493
rect 776 1476 778 1493
rect 808 1477 810 1493
rect 896 1477 898 1493
rect 936 1477 938 1493
rect 1024 1477 1026 1493
rect 806 1476 812 1477
rect 174 1475 180 1476
rect 110 1473 116 1474
rect 110 1469 111 1473
rect 115 1469 116 1473
rect 174 1471 175 1475
rect 179 1471 180 1475
rect 174 1470 180 1471
rect 206 1475 212 1476
rect 206 1471 207 1475
rect 211 1471 212 1475
rect 206 1470 212 1471
rect 238 1475 244 1476
rect 238 1471 239 1475
rect 243 1471 244 1475
rect 238 1470 244 1471
rect 270 1475 276 1476
rect 270 1471 271 1475
rect 275 1471 276 1475
rect 270 1470 276 1471
rect 302 1475 308 1476
rect 302 1471 303 1475
rect 307 1471 308 1475
rect 302 1470 308 1471
rect 334 1475 340 1476
rect 334 1471 335 1475
rect 339 1471 340 1475
rect 334 1470 340 1471
rect 366 1475 372 1476
rect 366 1471 367 1475
rect 371 1471 372 1475
rect 366 1470 372 1471
rect 398 1475 404 1476
rect 398 1471 399 1475
rect 403 1471 404 1475
rect 398 1470 404 1471
rect 430 1475 436 1476
rect 430 1471 431 1475
rect 435 1471 436 1475
rect 430 1470 436 1471
rect 462 1475 468 1476
rect 462 1471 463 1475
rect 467 1471 468 1475
rect 462 1470 468 1471
rect 494 1475 500 1476
rect 494 1471 495 1475
rect 499 1471 500 1475
rect 494 1470 500 1471
rect 526 1475 532 1476
rect 526 1471 527 1475
rect 531 1471 532 1475
rect 526 1470 532 1471
rect 558 1475 564 1476
rect 558 1471 559 1475
rect 563 1471 564 1475
rect 558 1470 564 1471
rect 590 1475 596 1476
rect 590 1471 591 1475
rect 595 1471 596 1475
rect 590 1470 596 1471
rect 622 1475 628 1476
rect 622 1471 623 1475
rect 627 1471 628 1475
rect 622 1470 628 1471
rect 662 1475 668 1476
rect 662 1471 663 1475
rect 667 1471 668 1475
rect 662 1470 668 1471
rect 702 1475 708 1476
rect 702 1471 703 1475
rect 707 1471 708 1475
rect 702 1470 708 1471
rect 742 1475 748 1476
rect 742 1471 743 1475
rect 747 1471 748 1475
rect 742 1470 748 1471
rect 774 1475 780 1476
rect 774 1471 775 1475
rect 779 1471 780 1475
rect 806 1472 807 1476
rect 811 1472 812 1476
rect 806 1471 812 1472
rect 894 1476 900 1477
rect 894 1472 895 1476
rect 899 1472 900 1476
rect 894 1471 900 1472
rect 934 1476 940 1477
rect 934 1472 935 1476
rect 939 1472 940 1476
rect 934 1471 940 1472
rect 1022 1476 1028 1477
rect 1080 1476 1082 1493
rect 1112 1477 1114 1493
rect 1110 1476 1116 1477
rect 1168 1476 1170 1493
rect 1200 1476 1202 1493
rect 1240 1476 1242 1493
rect 1280 1476 1282 1493
rect 1320 1476 1322 1493
rect 1360 1476 1362 1493
rect 1400 1476 1402 1493
rect 1440 1476 1442 1493
rect 1480 1476 1482 1493
rect 1520 1476 1522 1493
rect 1560 1476 1562 1493
rect 1592 1476 1594 1493
rect 1624 1476 1626 1493
rect 1656 1476 1658 1493
rect 1022 1472 1023 1476
rect 1027 1472 1028 1476
rect 1022 1471 1028 1472
rect 1078 1475 1084 1476
rect 1078 1471 1079 1475
rect 1083 1471 1084 1475
rect 1110 1472 1111 1476
rect 1115 1472 1116 1476
rect 1110 1471 1116 1472
rect 1166 1475 1172 1476
rect 1166 1471 1167 1475
rect 1171 1471 1172 1475
rect 774 1470 780 1471
rect 1078 1470 1084 1471
rect 1166 1470 1172 1471
rect 1198 1475 1204 1476
rect 1198 1471 1199 1475
rect 1203 1471 1204 1475
rect 1198 1470 1204 1471
rect 1238 1475 1244 1476
rect 1238 1471 1239 1475
rect 1243 1471 1244 1475
rect 1238 1470 1244 1471
rect 1278 1475 1284 1476
rect 1278 1471 1279 1475
rect 1283 1471 1284 1475
rect 1278 1470 1284 1471
rect 1318 1475 1324 1476
rect 1318 1471 1319 1475
rect 1323 1471 1324 1475
rect 1318 1470 1324 1471
rect 1358 1475 1364 1476
rect 1358 1471 1359 1475
rect 1363 1471 1364 1475
rect 1358 1470 1364 1471
rect 1398 1475 1404 1476
rect 1398 1471 1399 1475
rect 1403 1471 1404 1475
rect 1398 1470 1404 1471
rect 1438 1475 1444 1476
rect 1438 1471 1439 1475
rect 1443 1471 1444 1475
rect 1438 1470 1444 1471
rect 1478 1475 1484 1476
rect 1478 1471 1479 1475
rect 1483 1471 1484 1475
rect 1478 1470 1484 1471
rect 1518 1475 1524 1476
rect 1518 1471 1519 1475
rect 1523 1471 1524 1475
rect 1518 1470 1524 1471
rect 1558 1475 1564 1476
rect 1558 1471 1559 1475
rect 1563 1471 1564 1475
rect 1558 1470 1564 1471
rect 1590 1475 1596 1476
rect 1590 1471 1591 1475
rect 1595 1471 1596 1475
rect 1590 1470 1596 1471
rect 1622 1475 1628 1476
rect 1622 1471 1623 1475
rect 1627 1471 1628 1475
rect 1622 1470 1628 1471
rect 1654 1475 1660 1476
rect 1654 1471 1655 1475
rect 1659 1471 1660 1475
rect 1696 1474 1698 1493
rect 1654 1470 1660 1471
rect 1694 1473 1700 1474
rect 110 1468 116 1469
rect 1694 1469 1695 1473
rect 1699 1469 1700 1473
rect 1694 1468 1700 1469
rect 174 1458 180 1459
rect 110 1456 116 1457
rect 110 1452 111 1456
rect 115 1452 116 1456
rect 174 1454 175 1458
rect 179 1454 180 1458
rect 174 1453 180 1454
rect 206 1458 212 1459
rect 206 1454 207 1458
rect 211 1454 212 1458
rect 206 1453 212 1454
rect 238 1458 244 1459
rect 238 1454 239 1458
rect 243 1454 244 1458
rect 238 1453 244 1454
rect 270 1458 276 1459
rect 270 1454 271 1458
rect 275 1454 276 1458
rect 270 1453 276 1454
rect 302 1458 308 1459
rect 302 1454 303 1458
rect 307 1454 308 1458
rect 302 1453 308 1454
rect 334 1458 340 1459
rect 334 1454 335 1458
rect 339 1454 340 1458
rect 334 1453 340 1454
rect 366 1458 372 1459
rect 366 1454 367 1458
rect 371 1454 372 1458
rect 366 1453 372 1454
rect 398 1458 404 1459
rect 398 1454 399 1458
rect 403 1454 404 1458
rect 398 1453 404 1454
rect 430 1458 436 1459
rect 430 1454 431 1458
rect 435 1454 436 1458
rect 430 1453 436 1454
rect 462 1458 468 1459
rect 462 1454 463 1458
rect 467 1454 468 1458
rect 462 1453 468 1454
rect 494 1458 500 1459
rect 494 1454 495 1458
rect 499 1454 500 1458
rect 494 1453 500 1454
rect 526 1458 532 1459
rect 526 1454 527 1458
rect 531 1454 532 1458
rect 526 1453 532 1454
rect 558 1458 564 1459
rect 558 1454 559 1458
rect 563 1454 564 1458
rect 558 1453 564 1454
rect 590 1458 596 1459
rect 590 1454 591 1458
rect 595 1454 596 1458
rect 590 1453 596 1454
rect 622 1458 628 1459
rect 622 1454 623 1458
rect 627 1454 628 1458
rect 622 1453 628 1454
rect 662 1458 668 1459
rect 662 1454 663 1458
rect 667 1454 668 1458
rect 662 1453 668 1454
rect 702 1458 708 1459
rect 702 1454 703 1458
rect 707 1454 708 1458
rect 702 1453 708 1454
rect 742 1458 748 1459
rect 1078 1458 1084 1459
rect 742 1454 743 1458
rect 747 1454 748 1458
rect 742 1453 748 1454
rect 774 1457 780 1458
rect 774 1453 775 1457
rect 779 1453 780 1457
rect 110 1451 116 1452
rect 112 1431 114 1451
rect 176 1431 178 1453
rect 208 1431 210 1453
rect 240 1431 242 1453
rect 272 1431 274 1453
rect 304 1431 306 1453
rect 336 1431 338 1453
rect 368 1431 370 1453
rect 400 1431 402 1453
rect 432 1431 434 1453
rect 464 1431 466 1453
rect 496 1431 498 1453
rect 528 1431 530 1453
rect 560 1431 562 1453
rect 592 1431 594 1453
rect 624 1431 626 1453
rect 664 1431 666 1453
rect 704 1431 706 1453
rect 744 1431 746 1453
rect 774 1452 780 1453
rect 806 1457 812 1458
rect 806 1453 807 1457
rect 811 1453 812 1457
rect 806 1452 812 1453
rect 934 1457 940 1458
rect 934 1453 935 1457
rect 939 1453 940 1457
rect 934 1452 940 1453
rect 1038 1455 1044 1456
rect 776 1431 778 1452
rect 808 1431 810 1452
rect 894 1448 900 1449
rect 894 1444 895 1448
rect 899 1444 900 1448
rect 894 1443 900 1444
rect 896 1431 898 1443
rect 936 1431 938 1452
rect 1038 1451 1039 1455
rect 1043 1451 1044 1455
rect 1078 1454 1079 1458
rect 1083 1454 1084 1458
rect 1166 1458 1172 1459
rect 1078 1453 1084 1454
rect 1126 1455 1132 1456
rect 1038 1450 1044 1451
rect 1040 1431 1042 1450
rect 1080 1431 1082 1453
rect 1126 1451 1127 1455
rect 1131 1451 1132 1455
rect 1166 1454 1167 1458
rect 1171 1454 1172 1458
rect 1166 1453 1172 1454
rect 1198 1458 1204 1459
rect 1198 1454 1199 1458
rect 1203 1454 1204 1458
rect 1198 1453 1204 1454
rect 1238 1458 1244 1459
rect 1318 1458 1324 1459
rect 1238 1454 1239 1458
rect 1243 1454 1244 1458
rect 1238 1453 1244 1454
rect 1278 1457 1284 1458
rect 1278 1453 1279 1457
rect 1283 1453 1284 1457
rect 1318 1454 1319 1458
rect 1323 1454 1324 1458
rect 1318 1453 1324 1454
rect 1358 1458 1364 1459
rect 1358 1454 1359 1458
rect 1363 1454 1364 1458
rect 1358 1453 1364 1454
rect 1398 1458 1404 1459
rect 1398 1454 1399 1458
rect 1403 1454 1404 1458
rect 1398 1453 1404 1454
rect 1438 1458 1444 1459
rect 1438 1454 1439 1458
rect 1443 1454 1444 1458
rect 1438 1453 1444 1454
rect 1478 1458 1484 1459
rect 1478 1454 1479 1458
rect 1483 1454 1484 1458
rect 1478 1453 1484 1454
rect 1518 1458 1524 1459
rect 1518 1454 1519 1458
rect 1523 1454 1524 1458
rect 1518 1453 1524 1454
rect 1558 1458 1564 1459
rect 1558 1454 1559 1458
rect 1563 1454 1564 1458
rect 1558 1453 1564 1454
rect 1590 1458 1596 1459
rect 1590 1454 1591 1458
rect 1595 1454 1596 1458
rect 1590 1453 1596 1454
rect 1622 1458 1628 1459
rect 1622 1454 1623 1458
rect 1627 1454 1628 1458
rect 1622 1453 1628 1454
rect 1654 1458 1660 1459
rect 1654 1454 1655 1458
rect 1659 1454 1660 1458
rect 1654 1453 1660 1454
rect 1694 1456 1700 1457
rect 1126 1450 1132 1451
rect 1128 1431 1130 1450
rect 1168 1431 1170 1453
rect 1200 1431 1202 1453
rect 1240 1431 1242 1453
rect 1278 1452 1284 1453
rect 1280 1431 1282 1452
rect 1320 1431 1322 1453
rect 1360 1431 1362 1453
rect 1400 1431 1402 1453
rect 1440 1431 1442 1453
rect 1480 1431 1482 1453
rect 1520 1431 1522 1453
rect 1560 1431 1562 1453
rect 1592 1431 1594 1453
rect 1624 1431 1626 1453
rect 1656 1431 1658 1453
rect 1694 1452 1695 1456
rect 1699 1452 1700 1456
rect 1694 1451 1700 1452
rect 1696 1431 1698 1451
rect 111 1430 115 1431
rect 111 1425 115 1426
rect 135 1430 139 1431
rect 135 1425 139 1426
rect 167 1430 171 1431
rect 167 1425 171 1426
rect 175 1430 179 1431
rect 175 1425 179 1426
rect 199 1430 203 1431
rect 199 1425 203 1426
rect 207 1430 211 1431
rect 207 1425 211 1426
rect 231 1430 235 1431
rect 231 1425 235 1426
rect 239 1430 243 1431
rect 239 1425 243 1426
rect 263 1430 267 1431
rect 263 1425 267 1426
rect 271 1430 275 1431
rect 271 1425 275 1426
rect 295 1430 299 1431
rect 295 1425 299 1426
rect 303 1430 307 1431
rect 303 1425 307 1426
rect 327 1430 331 1431
rect 327 1425 331 1426
rect 335 1430 339 1431
rect 335 1425 339 1426
rect 359 1430 363 1431
rect 359 1425 363 1426
rect 367 1430 371 1431
rect 367 1425 371 1426
rect 391 1430 395 1431
rect 391 1425 395 1426
rect 399 1430 403 1431
rect 399 1425 403 1426
rect 423 1430 427 1431
rect 423 1425 427 1426
rect 431 1430 435 1431
rect 431 1425 435 1426
rect 455 1430 459 1431
rect 455 1425 459 1426
rect 463 1430 467 1431
rect 463 1425 467 1426
rect 487 1430 491 1431
rect 487 1425 491 1426
rect 495 1430 499 1431
rect 495 1425 499 1426
rect 519 1430 523 1431
rect 519 1425 523 1426
rect 527 1430 531 1431
rect 527 1425 531 1426
rect 551 1430 555 1431
rect 551 1425 555 1426
rect 559 1430 563 1431
rect 559 1425 563 1426
rect 583 1430 587 1431
rect 583 1425 587 1426
rect 591 1430 595 1431
rect 591 1425 595 1426
rect 615 1430 619 1431
rect 615 1425 619 1426
rect 623 1430 627 1431
rect 623 1425 627 1426
rect 647 1430 651 1431
rect 647 1425 651 1426
rect 663 1430 667 1431
rect 663 1425 667 1426
rect 679 1430 683 1431
rect 679 1425 683 1426
rect 703 1430 707 1431
rect 703 1425 707 1426
rect 719 1430 723 1431
rect 719 1425 723 1426
rect 743 1430 747 1431
rect 743 1425 747 1426
rect 767 1430 771 1431
rect 767 1425 771 1426
rect 775 1430 779 1431
rect 775 1425 779 1426
rect 807 1430 811 1431
rect 807 1425 811 1426
rect 839 1430 843 1431
rect 839 1425 843 1426
rect 895 1430 899 1431
rect 895 1425 899 1426
rect 935 1430 939 1431
rect 935 1425 939 1426
rect 975 1430 979 1431
rect 975 1425 979 1426
rect 1023 1430 1027 1431
rect 1023 1425 1027 1426
rect 1039 1430 1043 1431
rect 1039 1425 1043 1426
rect 1063 1430 1067 1431
rect 1063 1425 1067 1426
rect 1079 1430 1083 1431
rect 1079 1425 1083 1426
rect 1111 1430 1115 1431
rect 1111 1425 1115 1426
rect 1127 1430 1131 1431
rect 1127 1425 1131 1426
rect 1151 1430 1155 1431
rect 1151 1425 1155 1426
rect 1167 1430 1171 1431
rect 1167 1425 1171 1426
rect 1199 1430 1203 1431
rect 1199 1425 1203 1426
rect 1239 1430 1243 1431
rect 1239 1425 1243 1426
rect 1263 1430 1267 1431
rect 1263 1425 1267 1426
rect 1279 1430 1283 1431
rect 1279 1425 1283 1426
rect 1319 1430 1323 1431
rect 1319 1425 1323 1426
rect 1359 1430 1363 1431
rect 1359 1425 1363 1426
rect 1399 1430 1403 1431
rect 1399 1425 1403 1426
rect 1415 1430 1419 1431
rect 1415 1425 1419 1426
rect 1439 1430 1443 1431
rect 1439 1425 1443 1426
rect 1479 1430 1483 1431
rect 1479 1425 1483 1426
rect 1519 1430 1523 1431
rect 1519 1425 1523 1426
rect 1535 1430 1539 1431
rect 1535 1425 1539 1426
rect 1559 1430 1563 1431
rect 1559 1425 1563 1426
rect 1583 1430 1587 1431
rect 1583 1425 1587 1426
rect 1591 1430 1595 1431
rect 1591 1425 1595 1426
rect 1623 1430 1627 1431
rect 1623 1425 1627 1426
rect 1655 1430 1659 1431
rect 1655 1425 1659 1426
rect 1695 1430 1699 1431
rect 1695 1425 1699 1426
rect 112 1393 114 1425
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 136 1391 138 1425
rect 168 1391 170 1425
rect 200 1391 202 1425
rect 232 1391 234 1425
rect 264 1391 266 1425
rect 296 1391 298 1425
rect 328 1391 330 1425
rect 360 1391 362 1425
rect 392 1391 394 1425
rect 424 1391 426 1425
rect 456 1391 458 1425
rect 488 1391 490 1425
rect 520 1391 522 1425
rect 552 1391 554 1425
rect 584 1391 586 1425
rect 616 1391 618 1425
rect 648 1391 650 1425
rect 680 1391 682 1425
rect 720 1394 722 1425
rect 768 1416 770 1425
rect 766 1415 772 1416
rect 766 1411 767 1415
rect 771 1411 772 1415
rect 766 1410 772 1411
rect 808 1396 810 1425
rect 840 1416 842 1425
rect 838 1415 844 1416
rect 838 1411 839 1415
rect 843 1411 844 1415
rect 896 1411 898 1425
rect 976 1416 978 1425
rect 974 1415 980 1416
rect 974 1411 975 1415
rect 979 1411 980 1415
rect 838 1410 844 1411
rect 894 1410 900 1411
rect 974 1410 980 1411
rect 894 1406 895 1410
rect 899 1406 900 1410
rect 894 1405 900 1406
rect 806 1395 812 1396
rect 718 1393 724 1394
rect 110 1387 116 1388
rect 134 1390 140 1391
rect 134 1386 135 1390
rect 139 1386 140 1390
rect 134 1385 140 1386
rect 166 1390 172 1391
rect 166 1386 167 1390
rect 171 1386 172 1390
rect 166 1385 172 1386
rect 198 1390 204 1391
rect 198 1386 199 1390
rect 203 1386 204 1390
rect 198 1385 204 1386
rect 230 1390 236 1391
rect 230 1386 231 1390
rect 235 1386 236 1390
rect 230 1385 236 1386
rect 262 1390 268 1391
rect 262 1386 263 1390
rect 267 1386 268 1390
rect 262 1385 268 1386
rect 294 1390 300 1391
rect 294 1386 295 1390
rect 299 1386 300 1390
rect 294 1385 300 1386
rect 326 1390 332 1391
rect 326 1386 327 1390
rect 331 1386 332 1390
rect 326 1385 332 1386
rect 358 1390 364 1391
rect 358 1386 359 1390
rect 363 1386 364 1390
rect 358 1385 364 1386
rect 390 1390 396 1391
rect 390 1386 391 1390
rect 395 1386 396 1390
rect 390 1385 396 1386
rect 422 1390 428 1391
rect 422 1386 423 1390
rect 427 1386 428 1390
rect 422 1385 428 1386
rect 454 1390 460 1391
rect 454 1386 455 1390
rect 459 1386 460 1390
rect 454 1385 460 1386
rect 486 1390 492 1391
rect 486 1386 487 1390
rect 491 1386 492 1390
rect 486 1385 492 1386
rect 518 1390 524 1391
rect 518 1386 519 1390
rect 523 1386 524 1390
rect 518 1385 524 1386
rect 550 1390 556 1391
rect 550 1386 551 1390
rect 555 1386 556 1390
rect 550 1385 556 1386
rect 582 1390 588 1391
rect 582 1386 583 1390
rect 587 1386 588 1390
rect 582 1385 588 1386
rect 614 1390 620 1391
rect 614 1386 615 1390
rect 619 1386 620 1390
rect 614 1385 620 1386
rect 646 1390 652 1391
rect 646 1386 647 1390
rect 651 1386 652 1390
rect 646 1385 652 1386
rect 678 1390 684 1391
rect 678 1386 679 1390
rect 683 1386 684 1390
rect 718 1389 719 1393
rect 723 1389 724 1393
rect 806 1391 807 1395
rect 811 1391 812 1395
rect 1024 1391 1026 1425
rect 1064 1401 1066 1425
rect 1062 1400 1068 1401
rect 1062 1396 1063 1400
rect 1067 1396 1068 1400
rect 1062 1395 1068 1396
rect 1112 1392 1114 1425
rect 1152 1401 1154 1425
rect 1150 1400 1156 1401
rect 1150 1396 1151 1400
rect 1155 1396 1156 1400
rect 1150 1395 1156 1396
rect 1110 1391 1116 1392
rect 1200 1391 1202 1425
rect 1264 1394 1266 1425
rect 1262 1393 1268 1394
rect 806 1390 812 1391
rect 1022 1390 1028 1391
rect 718 1388 724 1389
rect 678 1385 684 1386
rect 1022 1386 1023 1390
rect 1027 1386 1028 1390
rect 1110 1387 1111 1391
rect 1115 1387 1116 1391
rect 1110 1386 1116 1387
rect 1198 1390 1204 1391
rect 1198 1386 1199 1390
rect 1203 1386 1204 1390
rect 1262 1389 1263 1393
rect 1267 1389 1268 1393
rect 1320 1392 1322 1425
rect 1262 1388 1268 1389
rect 1318 1391 1324 1392
rect 1416 1391 1418 1425
rect 1480 1394 1482 1425
rect 1478 1393 1484 1394
rect 1318 1387 1319 1391
rect 1323 1387 1324 1391
rect 1318 1386 1324 1387
rect 1414 1390 1420 1391
rect 1414 1386 1415 1390
rect 1419 1386 1420 1390
rect 1478 1389 1479 1393
rect 1483 1389 1484 1393
rect 1536 1391 1538 1425
rect 1584 1391 1586 1425
rect 1624 1391 1626 1425
rect 1656 1391 1658 1425
rect 1696 1393 1698 1425
rect 1694 1392 1700 1393
rect 1478 1388 1484 1389
rect 1534 1390 1540 1391
rect 1022 1385 1028 1386
rect 1198 1385 1204 1386
rect 1414 1385 1420 1386
rect 1534 1386 1535 1390
rect 1539 1386 1540 1390
rect 1534 1385 1540 1386
rect 1582 1390 1588 1391
rect 1582 1386 1583 1390
rect 1587 1386 1588 1390
rect 1582 1385 1588 1386
rect 1622 1390 1628 1391
rect 1622 1386 1623 1390
rect 1627 1386 1628 1390
rect 1622 1385 1628 1386
rect 1654 1390 1660 1391
rect 1654 1386 1655 1390
rect 1659 1386 1660 1390
rect 1694 1388 1695 1392
rect 1699 1388 1700 1392
rect 1694 1387 1700 1388
rect 1654 1385 1660 1386
rect 110 1375 116 1376
rect 110 1371 111 1375
rect 115 1371 116 1375
rect 1694 1375 1700 1376
rect 110 1370 116 1371
rect 134 1373 140 1374
rect 112 1351 114 1370
rect 134 1369 135 1373
rect 139 1369 140 1373
rect 134 1368 140 1369
rect 166 1373 172 1374
rect 166 1369 167 1373
rect 171 1369 172 1373
rect 166 1368 172 1369
rect 198 1373 204 1374
rect 198 1369 199 1373
rect 203 1369 204 1373
rect 198 1368 204 1369
rect 230 1373 236 1374
rect 230 1369 231 1373
rect 235 1369 236 1373
rect 230 1368 236 1369
rect 262 1373 268 1374
rect 262 1369 263 1373
rect 267 1369 268 1373
rect 262 1368 268 1369
rect 294 1373 300 1374
rect 294 1369 295 1373
rect 299 1369 300 1373
rect 294 1368 300 1369
rect 326 1373 332 1374
rect 326 1369 327 1373
rect 331 1369 332 1373
rect 326 1368 332 1369
rect 358 1373 364 1374
rect 358 1369 359 1373
rect 363 1369 364 1373
rect 358 1368 364 1369
rect 390 1373 396 1374
rect 390 1369 391 1373
rect 395 1369 396 1373
rect 390 1368 396 1369
rect 422 1373 428 1374
rect 422 1369 423 1373
rect 427 1369 428 1373
rect 422 1368 428 1369
rect 454 1373 460 1374
rect 454 1369 455 1373
rect 459 1369 460 1373
rect 454 1368 460 1369
rect 486 1373 492 1374
rect 486 1369 487 1373
rect 491 1369 492 1373
rect 486 1368 492 1369
rect 518 1373 524 1374
rect 518 1369 519 1373
rect 523 1369 524 1373
rect 518 1368 524 1369
rect 550 1373 556 1374
rect 550 1369 551 1373
rect 555 1369 556 1373
rect 550 1368 556 1369
rect 582 1373 588 1374
rect 582 1369 583 1373
rect 587 1369 588 1373
rect 582 1368 588 1369
rect 614 1373 620 1374
rect 614 1369 615 1373
rect 619 1369 620 1373
rect 614 1368 620 1369
rect 646 1373 652 1374
rect 646 1369 647 1373
rect 651 1369 652 1373
rect 646 1368 652 1369
rect 678 1373 684 1374
rect 1022 1373 1028 1374
rect 1110 1373 1116 1374
rect 1198 1373 1204 1374
rect 1414 1373 1420 1374
rect 1534 1373 1540 1374
rect 678 1369 679 1373
rect 683 1369 684 1373
rect 806 1372 812 1373
rect 678 1368 684 1369
rect 766 1368 772 1369
rect 136 1351 138 1368
rect 168 1351 170 1368
rect 200 1351 202 1368
rect 232 1351 234 1368
rect 264 1351 266 1368
rect 296 1351 298 1368
rect 328 1351 330 1368
rect 360 1351 362 1368
rect 392 1351 394 1368
rect 424 1351 426 1368
rect 456 1351 458 1368
rect 488 1351 490 1368
rect 520 1351 522 1368
rect 552 1351 554 1368
rect 584 1351 586 1368
rect 616 1351 618 1368
rect 648 1351 650 1368
rect 680 1351 682 1368
rect 734 1366 740 1367
rect 734 1362 735 1366
rect 739 1362 740 1366
rect 766 1364 767 1368
rect 771 1364 772 1368
rect 806 1368 807 1372
rect 811 1368 812 1372
rect 886 1372 892 1373
rect 806 1367 812 1368
rect 838 1368 844 1369
rect 766 1363 772 1364
rect 734 1361 740 1362
rect 736 1351 738 1361
rect 768 1351 770 1363
rect 808 1351 810 1367
rect 838 1364 839 1368
rect 843 1364 844 1368
rect 886 1368 887 1372
rect 891 1368 892 1372
rect 1022 1369 1023 1373
rect 1027 1369 1028 1373
rect 886 1367 892 1368
rect 974 1368 980 1369
rect 1022 1368 1028 1369
rect 1062 1372 1068 1373
rect 1062 1368 1063 1372
rect 1067 1368 1068 1372
rect 1110 1369 1111 1373
rect 1115 1369 1116 1373
rect 1110 1368 1116 1369
rect 1150 1372 1156 1373
rect 1150 1368 1151 1372
rect 1155 1368 1156 1372
rect 1198 1369 1199 1373
rect 1203 1369 1204 1373
rect 1198 1368 1204 1369
rect 1246 1372 1252 1373
rect 1246 1368 1247 1372
rect 1251 1368 1252 1372
rect 838 1363 844 1364
rect 840 1351 842 1363
rect 888 1351 890 1367
rect 974 1364 975 1368
rect 979 1364 980 1368
rect 974 1363 980 1364
rect 976 1351 978 1363
rect 1024 1351 1026 1368
rect 1062 1367 1068 1368
rect 1064 1351 1066 1367
rect 1112 1351 1114 1368
rect 1150 1367 1156 1368
rect 1152 1351 1154 1367
rect 1200 1351 1202 1368
rect 1246 1367 1252 1368
rect 1318 1372 1324 1373
rect 1318 1368 1319 1372
rect 1323 1368 1324 1372
rect 1414 1369 1415 1373
rect 1419 1369 1420 1373
rect 1414 1368 1420 1369
rect 1462 1372 1468 1373
rect 1462 1368 1463 1372
rect 1467 1368 1468 1372
rect 1534 1369 1535 1373
rect 1539 1369 1540 1373
rect 1534 1368 1540 1369
rect 1582 1373 1588 1374
rect 1582 1369 1583 1373
rect 1587 1369 1588 1373
rect 1582 1368 1588 1369
rect 1622 1373 1628 1374
rect 1622 1369 1623 1373
rect 1627 1369 1628 1373
rect 1622 1368 1628 1369
rect 1654 1373 1660 1374
rect 1654 1369 1655 1373
rect 1659 1369 1660 1373
rect 1694 1371 1695 1375
rect 1699 1371 1700 1375
rect 1694 1370 1700 1371
rect 1654 1368 1660 1369
rect 1318 1367 1324 1368
rect 1248 1351 1250 1367
rect 1320 1351 1322 1367
rect 1416 1351 1418 1368
rect 1462 1367 1468 1368
rect 1464 1351 1466 1367
rect 1536 1351 1538 1368
rect 1584 1351 1586 1368
rect 1624 1351 1626 1368
rect 1656 1351 1658 1368
rect 1696 1351 1698 1370
rect 111 1350 115 1351
rect 111 1345 115 1346
rect 135 1350 139 1351
rect 135 1345 139 1346
rect 167 1350 171 1351
rect 167 1345 171 1346
rect 199 1350 203 1351
rect 199 1345 203 1346
rect 231 1350 235 1351
rect 231 1345 235 1346
rect 263 1350 267 1351
rect 263 1345 267 1346
rect 295 1350 299 1351
rect 295 1345 299 1346
rect 327 1350 331 1351
rect 327 1345 331 1346
rect 359 1350 363 1351
rect 359 1345 363 1346
rect 391 1350 395 1351
rect 391 1345 395 1346
rect 423 1350 427 1351
rect 423 1345 427 1346
rect 455 1350 459 1351
rect 455 1345 459 1346
rect 487 1350 491 1351
rect 487 1345 491 1346
rect 519 1350 523 1351
rect 519 1345 523 1346
rect 551 1350 555 1351
rect 551 1345 555 1346
rect 583 1350 587 1351
rect 583 1345 587 1346
rect 615 1350 619 1351
rect 615 1345 619 1346
rect 647 1350 651 1351
rect 647 1345 651 1346
rect 679 1350 683 1351
rect 679 1345 683 1346
rect 711 1350 715 1351
rect 711 1345 715 1346
rect 735 1350 739 1351
rect 735 1345 739 1346
rect 743 1350 747 1351
rect 743 1345 747 1346
rect 767 1350 771 1351
rect 767 1345 771 1346
rect 807 1350 811 1351
rect 807 1345 811 1346
rect 823 1350 827 1351
rect 823 1345 827 1346
rect 839 1350 843 1351
rect 839 1345 843 1346
rect 887 1350 891 1351
rect 887 1345 891 1346
rect 903 1350 907 1351
rect 903 1345 907 1346
rect 975 1350 979 1351
rect 975 1345 979 1346
rect 983 1350 987 1351
rect 983 1345 987 1346
rect 1023 1350 1027 1351
rect 1023 1345 1027 1346
rect 1063 1350 1067 1351
rect 1063 1345 1067 1346
rect 1111 1350 1115 1351
rect 1111 1345 1115 1346
rect 1151 1350 1155 1351
rect 1151 1345 1155 1346
rect 1159 1350 1163 1351
rect 1159 1345 1163 1346
rect 1199 1350 1203 1351
rect 1199 1345 1203 1346
rect 1215 1350 1219 1351
rect 1215 1345 1219 1346
rect 1247 1350 1251 1351
rect 1247 1345 1251 1346
rect 1303 1350 1307 1351
rect 1303 1345 1307 1346
rect 1319 1350 1323 1351
rect 1319 1345 1323 1346
rect 1391 1350 1395 1351
rect 1391 1345 1395 1346
rect 1415 1350 1419 1351
rect 1415 1345 1419 1346
rect 1423 1350 1427 1351
rect 1423 1345 1427 1346
rect 1455 1350 1459 1351
rect 1455 1345 1459 1346
rect 1463 1350 1467 1351
rect 1463 1345 1467 1346
rect 1495 1350 1499 1351
rect 1495 1345 1499 1346
rect 1527 1350 1531 1351
rect 1527 1345 1531 1346
rect 1535 1350 1539 1351
rect 1535 1345 1539 1346
rect 1559 1350 1563 1351
rect 1559 1345 1563 1346
rect 1583 1350 1587 1351
rect 1583 1345 1587 1346
rect 1591 1350 1595 1351
rect 1591 1345 1595 1346
rect 1623 1350 1627 1351
rect 1623 1345 1627 1346
rect 1655 1350 1659 1351
rect 1655 1345 1659 1346
rect 1695 1350 1699 1351
rect 1695 1345 1699 1346
rect 112 1318 114 1345
rect 136 1320 138 1345
rect 168 1320 170 1345
rect 200 1320 202 1345
rect 232 1320 234 1345
rect 264 1320 266 1345
rect 296 1320 298 1345
rect 328 1320 330 1345
rect 360 1320 362 1345
rect 392 1320 394 1345
rect 424 1320 426 1345
rect 456 1320 458 1345
rect 488 1320 490 1345
rect 520 1320 522 1345
rect 552 1320 554 1345
rect 584 1320 586 1345
rect 616 1320 618 1345
rect 648 1320 650 1345
rect 680 1320 682 1345
rect 712 1320 714 1345
rect 744 1321 746 1345
rect 824 1321 826 1345
rect 904 1321 906 1345
rect 984 1325 986 1345
rect 982 1324 988 1325
rect 742 1320 748 1321
rect 134 1319 140 1320
rect 110 1317 116 1318
rect 110 1313 111 1317
rect 115 1313 116 1317
rect 134 1315 135 1319
rect 139 1315 140 1319
rect 134 1314 140 1315
rect 166 1319 172 1320
rect 166 1315 167 1319
rect 171 1315 172 1319
rect 166 1314 172 1315
rect 198 1319 204 1320
rect 198 1315 199 1319
rect 203 1315 204 1319
rect 198 1314 204 1315
rect 230 1319 236 1320
rect 230 1315 231 1319
rect 235 1315 236 1319
rect 230 1314 236 1315
rect 262 1319 268 1320
rect 262 1315 263 1319
rect 267 1315 268 1319
rect 262 1314 268 1315
rect 294 1319 300 1320
rect 294 1315 295 1319
rect 299 1315 300 1319
rect 294 1314 300 1315
rect 326 1319 332 1320
rect 326 1315 327 1319
rect 331 1315 332 1319
rect 326 1314 332 1315
rect 358 1319 364 1320
rect 358 1315 359 1319
rect 363 1315 364 1319
rect 358 1314 364 1315
rect 390 1319 396 1320
rect 390 1315 391 1319
rect 395 1315 396 1319
rect 390 1314 396 1315
rect 422 1319 428 1320
rect 422 1315 423 1319
rect 427 1315 428 1319
rect 422 1314 428 1315
rect 454 1319 460 1320
rect 454 1315 455 1319
rect 459 1315 460 1319
rect 454 1314 460 1315
rect 486 1319 492 1320
rect 486 1315 487 1319
rect 491 1315 492 1319
rect 486 1314 492 1315
rect 518 1319 524 1320
rect 518 1315 519 1319
rect 523 1315 524 1319
rect 518 1314 524 1315
rect 550 1319 556 1320
rect 550 1315 551 1319
rect 555 1315 556 1319
rect 550 1314 556 1315
rect 582 1319 588 1320
rect 582 1315 583 1319
rect 587 1315 588 1319
rect 582 1314 588 1315
rect 614 1319 620 1320
rect 614 1315 615 1319
rect 619 1315 620 1319
rect 614 1314 620 1315
rect 646 1319 652 1320
rect 646 1315 647 1319
rect 651 1315 652 1319
rect 646 1314 652 1315
rect 678 1319 684 1320
rect 678 1315 679 1319
rect 683 1315 684 1319
rect 678 1314 684 1315
rect 710 1319 716 1320
rect 710 1315 711 1319
rect 715 1315 716 1319
rect 742 1316 743 1320
rect 747 1316 748 1320
rect 742 1315 748 1316
rect 822 1320 828 1321
rect 822 1316 823 1320
rect 827 1316 828 1320
rect 822 1315 828 1316
rect 902 1320 908 1321
rect 902 1316 903 1320
rect 907 1316 908 1320
rect 982 1320 983 1324
rect 987 1320 988 1324
rect 1024 1321 1026 1345
rect 1064 1321 1066 1345
rect 1160 1321 1162 1345
rect 1216 1321 1218 1345
rect 1304 1321 1306 1345
rect 982 1319 988 1320
rect 1022 1320 1028 1321
rect 902 1315 908 1316
rect 1022 1316 1023 1320
rect 1027 1316 1028 1320
rect 1022 1315 1028 1316
rect 1062 1320 1068 1321
rect 1062 1316 1063 1320
rect 1067 1316 1068 1320
rect 1062 1315 1068 1316
rect 1158 1320 1164 1321
rect 1158 1316 1159 1320
rect 1163 1316 1164 1320
rect 1158 1315 1164 1316
rect 1214 1320 1220 1321
rect 1214 1316 1215 1320
rect 1219 1316 1220 1320
rect 1214 1315 1220 1316
rect 1302 1320 1308 1321
rect 1392 1320 1394 1345
rect 1424 1320 1426 1345
rect 1456 1321 1458 1345
rect 1454 1320 1460 1321
rect 1496 1320 1498 1345
rect 1528 1320 1530 1345
rect 1560 1320 1562 1345
rect 1592 1320 1594 1345
rect 1624 1320 1626 1345
rect 1656 1320 1658 1345
rect 1302 1316 1303 1320
rect 1307 1316 1308 1320
rect 1302 1315 1308 1316
rect 1390 1319 1396 1320
rect 1390 1315 1391 1319
rect 1395 1315 1396 1319
rect 710 1314 716 1315
rect 1390 1314 1396 1315
rect 1422 1319 1428 1320
rect 1422 1315 1423 1319
rect 1427 1315 1428 1319
rect 1454 1316 1455 1320
rect 1459 1316 1460 1320
rect 1454 1315 1460 1316
rect 1494 1319 1500 1320
rect 1494 1315 1495 1319
rect 1499 1315 1500 1319
rect 1422 1314 1428 1315
rect 1494 1314 1500 1315
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1558 1319 1564 1320
rect 1558 1315 1559 1319
rect 1563 1315 1564 1319
rect 1558 1314 1564 1315
rect 1590 1319 1596 1320
rect 1590 1315 1591 1319
rect 1595 1315 1596 1319
rect 1590 1314 1596 1315
rect 1622 1319 1628 1320
rect 1622 1315 1623 1319
rect 1627 1315 1628 1319
rect 1622 1314 1628 1315
rect 1654 1319 1660 1320
rect 1654 1315 1655 1319
rect 1659 1315 1660 1319
rect 1696 1318 1698 1345
rect 1654 1314 1660 1315
rect 1694 1317 1700 1318
rect 110 1312 116 1313
rect 1694 1313 1695 1317
rect 1699 1313 1700 1317
rect 1694 1312 1700 1313
rect 134 1302 140 1303
rect 110 1300 116 1301
rect 110 1296 111 1300
rect 115 1296 116 1300
rect 134 1298 135 1302
rect 139 1298 140 1302
rect 134 1297 140 1298
rect 166 1302 172 1303
rect 166 1298 167 1302
rect 171 1298 172 1302
rect 166 1297 172 1298
rect 198 1302 204 1303
rect 198 1298 199 1302
rect 203 1298 204 1302
rect 198 1297 204 1298
rect 230 1302 236 1303
rect 230 1298 231 1302
rect 235 1298 236 1302
rect 230 1297 236 1298
rect 262 1302 268 1303
rect 262 1298 263 1302
rect 267 1298 268 1302
rect 262 1297 268 1298
rect 294 1302 300 1303
rect 294 1298 295 1302
rect 299 1298 300 1302
rect 294 1297 300 1298
rect 326 1302 332 1303
rect 326 1298 327 1302
rect 331 1298 332 1302
rect 326 1297 332 1298
rect 358 1302 364 1303
rect 358 1298 359 1302
rect 363 1298 364 1302
rect 358 1297 364 1298
rect 390 1302 396 1303
rect 390 1298 391 1302
rect 395 1298 396 1302
rect 390 1297 396 1298
rect 422 1302 428 1303
rect 422 1298 423 1302
rect 427 1298 428 1302
rect 422 1297 428 1298
rect 454 1302 460 1303
rect 454 1298 455 1302
rect 459 1298 460 1302
rect 454 1297 460 1298
rect 486 1302 492 1303
rect 486 1298 487 1302
rect 491 1298 492 1302
rect 486 1297 492 1298
rect 518 1302 524 1303
rect 518 1298 519 1302
rect 523 1298 524 1302
rect 518 1297 524 1298
rect 550 1302 556 1303
rect 550 1298 551 1302
rect 555 1298 556 1302
rect 550 1297 556 1298
rect 582 1302 588 1303
rect 582 1298 583 1302
rect 587 1298 588 1302
rect 582 1297 588 1298
rect 614 1302 620 1303
rect 614 1298 615 1302
rect 619 1298 620 1302
rect 614 1297 620 1298
rect 646 1302 652 1303
rect 646 1298 647 1302
rect 651 1298 652 1302
rect 646 1297 652 1298
rect 678 1302 684 1303
rect 678 1298 679 1302
rect 683 1298 684 1302
rect 678 1297 684 1298
rect 710 1302 716 1303
rect 1422 1302 1428 1303
rect 710 1298 711 1302
rect 715 1298 716 1302
rect 710 1297 716 1298
rect 1062 1301 1068 1302
rect 1062 1297 1063 1301
rect 1067 1297 1068 1301
rect 1214 1301 1220 1302
rect 110 1295 116 1296
rect 112 1263 114 1295
rect 136 1263 138 1297
rect 168 1263 170 1297
rect 200 1263 202 1297
rect 232 1263 234 1297
rect 264 1263 266 1297
rect 296 1263 298 1297
rect 328 1263 330 1297
rect 360 1263 362 1297
rect 392 1263 394 1297
rect 424 1263 426 1297
rect 456 1263 458 1297
rect 488 1263 490 1297
rect 520 1263 522 1297
rect 552 1263 554 1297
rect 584 1263 586 1297
rect 616 1263 618 1297
rect 648 1263 650 1297
rect 680 1263 682 1297
rect 712 1263 714 1297
rect 1062 1296 1068 1297
rect 1174 1299 1180 1300
rect 1022 1292 1028 1293
rect 1022 1288 1023 1292
rect 1027 1288 1028 1292
rect 1022 1287 1028 1288
rect 750 1282 756 1283
rect 750 1278 751 1282
rect 755 1278 756 1282
rect 750 1277 756 1278
rect 830 1282 836 1283
rect 830 1278 831 1282
rect 835 1278 836 1282
rect 830 1277 836 1278
rect 910 1282 916 1283
rect 910 1278 911 1282
rect 915 1278 916 1282
rect 910 1277 916 1278
rect 982 1277 988 1278
rect 752 1263 754 1277
rect 832 1263 834 1277
rect 912 1263 914 1277
rect 982 1273 983 1277
rect 987 1273 988 1277
rect 982 1272 988 1273
rect 984 1263 986 1272
rect 1024 1263 1026 1287
rect 1064 1263 1066 1296
rect 1174 1295 1175 1299
rect 1179 1295 1180 1299
rect 1214 1297 1215 1301
rect 1219 1297 1220 1301
rect 1214 1296 1220 1297
rect 1302 1301 1308 1302
rect 1302 1297 1303 1301
rect 1307 1297 1308 1301
rect 1302 1296 1308 1297
rect 1390 1301 1396 1302
rect 1390 1297 1391 1301
rect 1395 1297 1396 1301
rect 1422 1298 1423 1302
rect 1427 1298 1428 1302
rect 1422 1297 1428 1298
rect 1494 1302 1500 1303
rect 1494 1298 1495 1302
rect 1499 1298 1500 1302
rect 1494 1297 1500 1298
rect 1526 1302 1532 1303
rect 1526 1298 1527 1302
rect 1531 1298 1532 1302
rect 1526 1297 1532 1298
rect 1558 1302 1564 1303
rect 1558 1298 1559 1302
rect 1563 1298 1564 1302
rect 1558 1297 1564 1298
rect 1590 1302 1596 1303
rect 1590 1298 1591 1302
rect 1595 1298 1596 1302
rect 1590 1297 1596 1298
rect 1622 1302 1628 1303
rect 1622 1298 1623 1302
rect 1627 1298 1628 1302
rect 1622 1297 1628 1298
rect 1654 1302 1660 1303
rect 1654 1298 1655 1302
rect 1659 1298 1660 1302
rect 1654 1297 1660 1298
rect 1694 1300 1700 1301
rect 1390 1296 1396 1297
rect 1174 1294 1180 1295
rect 1176 1263 1178 1294
rect 1216 1263 1218 1296
rect 1304 1263 1306 1296
rect 1392 1263 1394 1296
rect 1424 1263 1426 1297
rect 1454 1292 1460 1293
rect 1454 1288 1455 1292
rect 1459 1288 1460 1292
rect 1454 1287 1460 1288
rect 1456 1263 1458 1287
rect 1496 1263 1498 1297
rect 1528 1263 1530 1297
rect 1560 1263 1562 1297
rect 1592 1263 1594 1297
rect 1624 1263 1626 1297
rect 1656 1263 1658 1297
rect 1694 1296 1695 1300
rect 1699 1296 1700 1300
rect 1694 1295 1700 1296
rect 1696 1263 1698 1295
rect 111 1262 115 1263
rect 111 1257 115 1258
rect 135 1262 139 1263
rect 135 1257 139 1258
rect 167 1262 171 1263
rect 167 1257 171 1258
rect 199 1262 203 1263
rect 199 1257 203 1258
rect 231 1262 235 1263
rect 231 1257 235 1258
rect 263 1262 267 1263
rect 263 1257 267 1258
rect 295 1262 299 1263
rect 295 1257 299 1258
rect 327 1262 331 1263
rect 327 1257 331 1258
rect 359 1262 363 1263
rect 359 1257 363 1258
rect 391 1262 395 1263
rect 391 1257 395 1258
rect 423 1262 427 1263
rect 423 1257 427 1258
rect 455 1262 459 1263
rect 455 1257 459 1258
rect 487 1262 491 1263
rect 487 1257 491 1258
rect 519 1262 523 1263
rect 519 1257 523 1258
rect 551 1262 555 1263
rect 551 1257 555 1258
rect 583 1262 587 1263
rect 583 1257 587 1258
rect 615 1262 619 1263
rect 615 1257 619 1258
rect 647 1262 651 1263
rect 647 1257 651 1258
rect 679 1262 683 1263
rect 679 1257 683 1258
rect 711 1262 715 1263
rect 711 1257 715 1258
rect 743 1262 747 1263
rect 743 1257 747 1258
rect 751 1262 755 1263
rect 751 1257 755 1258
rect 775 1262 779 1263
rect 775 1257 779 1258
rect 811 1262 815 1263
rect 811 1257 815 1258
rect 831 1262 835 1263
rect 831 1257 835 1258
rect 911 1262 915 1263
rect 911 1257 915 1258
rect 959 1262 963 1263
rect 959 1257 963 1258
rect 983 1262 987 1263
rect 983 1257 987 1258
rect 1015 1262 1019 1263
rect 1015 1257 1019 1258
rect 1023 1262 1027 1263
rect 1023 1257 1027 1258
rect 1063 1262 1067 1263
rect 1063 1257 1067 1258
rect 1087 1262 1091 1263
rect 1087 1257 1091 1258
rect 1127 1262 1131 1263
rect 1127 1257 1131 1258
rect 1159 1262 1163 1263
rect 1159 1257 1163 1258
rect 1175 1262 1179 1263
rect 1175 1257 1179 1258
rect 1215 1262 1219 1263
rect 1215 1257 1219 1258
rect 1255 1262 1259 1263
rect 1255 1257 1259 1258
rect 1295 1262 1299 1263
rect 1295 1257 1299 1258
rect 1303 1262 1307 1263
rect 1303 1257 1307 1258
rect 1343 1262 1347 1263
rect 1343 1257 1347 1258
rect 1375 1262 1379 1263
rect 1375 1257 1379 1258
rect 1391 1262 1395 1263
rect 1391 1257 1395 1258
rect 1407 1262 1411 1263
rect 1407 1257 1411 1258
rect 1423 1262 1427 1263
rect 1423 1257 1427 1258
rect 1439 1262 1443 1263
rect 1439 1257 1443 1258
rect 1455 1262 1459 1263
rect 1455 1257 1459 1258
rect 1479 1262 1483 1263
rect 1479 1257 1483 1258
rect 1495 1262 1499 1263
rect 1495 1257 1499 1258
rect 1519 1262 1523 1263
rect 1519 1257 1523 1258
rect 1527 1262 1531 1263
rect 1527 1257 1531 1258
rect 1559 1262 1563 1263
rect 1559 1257 1563 1258
rect 1591 1262 1595 1263
rect 1591 1257 1595 1258
rect 1623 1262 1627 1263
rect 1623 1257 1627 1258
rect 1655 1262 1659 1263
rect 1655 1257 1659 1258
rect 1695 1262 1699 1263
rect 1695 1257 1699 1258
rect 112 1197 114 1257
rect 110 1196 116 1197
rect 110 1192 111 1196
rect 115 1192 116 1196
rect 136 1195 138 1257
rect 168 1195 170 1257
rect 200 1195 202 1257
rect 232 1195 234 1257
rect 264 1195 266 1257
rect 296 1195 298 1257
rect 328 1195 330 1257
rect 360 1195 362 1257
rect 392 1195 394 1257
rect 424 1195 426 1257
rect 456 1195 458 1257
rect 488 1195 490 1257
rect 520 1195 522 1257
rect 552 1195 554 1257
rect 584 1195 586 1257
rect 616 1195 618 1257
rect 648 1195 650 1257
rect 680 1195 682 1257
rect 712 1195 714 1257
rect 744 1195 746 1257
rect 776 1220 778 1257
rect 774 1219 780 1220
rect 774 1215 775 1219
rect 779 1215 780 1219
rect 774 1214 780 1215
rect 812 1196 814 1257
rect 960 1198 962 1257
rect 1016 1215 1018 1257
rect 1088 1220 1090 1257
rect 1086 1219 1092 1220
rect 1086 1215 1087 1219
rect 1091 1215 1092 1219
rect 1014 1214 1020 1215
rect 1086 1214 1092 1215
rect 1014 1210 1015 1214
rect 1019 1210 1020 1214
rect 1014 1209 1020 1210
rect 958 1197 964 1198
rect 810 1195 816 1196
rect 110 1191 116 1192
rect 134 1194 140 1195
rect 134 1190 135 1194
rect 139 1190 140 1194
rect 134 1189 140 1190
rect 166 1194 172 1195
rect 166 1190 167 1194
rect 171 1190 172 1194
rect 166 1189 172 1190
rect 198 1194 204 1195
rect 198 1190 199 1194
rect 203 1190 204 1194
rect 198 1189 204 1190
rect 230 1194 236 1195
rect 230 1190 231 1194
rect 235 1190 236 1194
rect 230 1189 236 1190
rect 262 1194 268 1195
rect 262 1190 263 1194
rect 267 1190 268 1194
rect 262 1189 268 1190
rect 294 1194 300 1195
rect 294 1190 295 1194
rect 299 1190 300 1194
rect 294 1189 300 1190
rect 326 1194 332 1195
rect 326 1190 327 1194
rect 331 1190 332 1194
rect 326 1189 332 1190
rect 358 1194 364 1195
rect 358 1190 359 1194
rect 363 1190 364 1194
rect 358 1189 364 1190
rect 390 1194 396 1195
rect 390 1190 391 1194
rect 395 1190 396 1194
rect 390 1189 396 1190
rect 422 1194 428 1195
rect 422 1190 423 1194
rect 427 1190 428 1194
rect 422 1189 428 1190
rect 454 1194 460 1195
rect 454 1190 455 1194
rect 459 1190 460 1194
rect 454 1189 460 1190
rect 486 1194 492 1195
rect 486 1190 487 1194
rect 491 1190 492 1194
rect 486 1189 492 1190
rect 518 1194 524 1195
rect 518 1190 519 1194
rect 523 1190 524 1194
rect 518 1189 524 1190
rect 550 1194 556 1195
rect 550 1190 551 1194
rect 555 1190 556 1194
rect 550 1189 556 1190
rect 582 1194 588 1195
rect 582 1190 583 1194
rect 587 1190 588 1194
rect 582 1189 588 1190
rect 614 1194 620 1195
rect 614 1190 615 1194
rect 619 1190 620 1194
rect 614 1189 620 1190
rect 646 1194 652 1195
rect 646 1190 647 1194
rect 651 1190 652 1194
rect 646 1189 652 1190
rect 678 1194 684 1195
rect 678 1190 679 1194
rect 683 1190 684 1194
rect 678 1189 684 1190
rect 710 1194 716 1195
rect 710 1190 711 1194
rect 715 1190 716 1194
rect 710 1189 716 1190
rect 742 1194 748 1195
rect 742 1190 743 1194
rect 747 1190 748 1194
rect 810 1191 811 1195
rect 815 1191 816 1195
rect 958 1193 959 1197
rect 963 1193 964 1197
rect 1128 1195 1130 1257
rect 1160 1195 1162 1257
rect 1216 1198 1218 1257
rect 1214 1197 1220 1198
rect 958 1192 964 1193
rect 1126 1194 1132 1195
rect 810 1190 816 1191
rect 1126 1190 1127 1194
rect 1131 1190 1132 1194
rect 742 1189 748 1190
rect 1126 1189 1132 1190
rect 1158 1194 1164 1195
rect 1158 1190 1159 1194
rect 1163 1190 1164 1194
rect 1214 1193 1215 1197
rect 1219 1193 1220 1197
rect 1256 1195 1258 1257
rect 1296 1198 1298 1257
rect 1294 1197 1300 1198
rect 1214 1192 1220 1193
rect 1254 1194 1260 1195
rect 1158 1189 1164 1190
rect 1254 1190 1255 1194
rect 1259 1190 1260 1194
rect 1294 1193 1295 1197
rect 1299 1193 1300 1197
rect 1344 1195 1346 1257
rect 1376 1195 1378 1257
rect 1408 1195 1410 1257
rect 1440 1195 1442 1257
rect 1480 1195 1482 1257
rect 1520 1195 1522 1257
rect 1560 1195 1562 1257
rect 1592 1195 1594 1257
rect 1624 1195 1626 1257
rect 1656 1195 1658 1257
rect 1696 1197 1698 1257
rect 1694 1196 1700 1197
rect 1294 1192 1300 1193
rect 1342 1194 1348 1195
rect 1254 1189 1260 1190
rect 1342 1190 1343 1194
rect 1347 1190 1348 1194
rect 1342 1189 1348 1190
rect 1374 1194 1380 1195
rect 1374 1190 1375 1194
rect 1379 1190 1380 1194
rect 1374 1189 1380 1190
rect 1406 1194 1412 1195
rect 1406 1190 1407 1194
rect 1411 1190 1412 1194
rect 1406 1189 1412 1190
rect 1438 1194 1444 1195
rect 1438 1190 1439 1194
rect 1443 1190 1444 1194
rect 1438 1189 1444 1190
rect 1478 1194 1484 1195
rect 1478 1190 1479 1194
rect 1483 1190 1484 1194
rect 1478 1189 1484 1190
rect 1518 1194 1524 1195
rect 1518 1190 1519 1194
rect 1523 1190 1524 1194
rect 1518 1189 1524 1190
rect 1558 1194 1564 1195
rect 1558 1190 1559 1194
rect 1563 1190 1564 1194
rect 1558 1189 1564 1190
rect 1590 1194 1596 1195
rect 1590 1190 1591 1194
rect 1595 1190 1596 1194
rect 1590 1189 1596 1190
rect 1622 1194 1628 1195
rect 1622 1190 1623 1194
rect 1627 1190 1628 1194
rect 1622 1189 1628 1190
rect 1654 1194 1660 1195
rect 1654 1190 1655 1194
rect 1659 1190 1660 1194
rect 1694 1192 1695 1196
rect 1699 1192 1700 1196
rect 1694 1191 1700 1192
rect 1654 1189 1660 1190
rect 838 1180 844 1181
rect 110 1179 116 1180
rect 110 1175 111 1179
rect 115 1175 116 1179
rect 110 1174 116 1175
rect 134 1177 140 1178
rect 112 1151 114 1174
rect 134 1173 135 1177
rect 139 1173 140 1177
rect 134 1172 140 1173
rect 166 1177 172 1178
rect 166 1173 167 1177
rect 171 1173 172 1177
rect 166 1172 172 1173
rect 198 1177 204 1178
rect 198 1173 199 1177
rect 203 1173 204 1177
rect 198 1172 204 1173
rect 230 1177 236 1178
rect 230 1173 231 1177
rect 235 1173 236 1177
rect 230 1172 236 1173
rect 262 1177 268 1178
rect 262 1173 263 1177
rect 267 1173 268 1177
rect 262 1172 268 1173
rect 294 1177 300 1178
rect 294 1173 295 1177
rect 299 1173 300 1177
rect 294 1172 300 1173
rect 326 1177 332 1178
rect 326 1173 327 1177
rect 331 1173 332 1177
rect 326 1172 332 1173
rect 358 1177 364 1178
rect 358 1173 359 1177
rect 363 1173 364 1177
rect 358 1172 364 1173
rect 390 1177 396 1178
rect 390 1173 391 1177
rect 395 1173 396 1177
rect 390 1172 396 1173
rect 422 1177 428 1178
rect 422 1173 423 1177
rect 427 1173 428 1177
rect 422 1172 428 1173
rect 454 1177 460 1178
rect 454 1173 455 1177
rect 459 1173 460 1177
rect 454 1172 460 1173
rect 486 1177 492 1178
rect 486 1173 487 1177
rect 491 1173 492 1177
rect 486 1172 492 1173
rect 518 1177 524 1178
rect 518 1173 519 1177
rect 523 1173 524 1177
rect 518 1172 524 1173
rect 550 1177 556 1178
rect 550 1173 551 1177
rect 555 1173 556 1177
rect 550 1172 556 1173
rect 582 1177 588 1178
rect 582 1173 583 1177
rect 587 1173 588 1177
rect 582 1172 588 1173
rect 614 1177 620 1178
rect 614 1173 615 1177
rect 619 1173 620 1177
rect 614 1172 620 1173
rect 646 1177 652 1178
rect 646 1173 647 1177
rect 651 1173 652 1177
rect 646 1172 652 1173
rect 678 1177 684 1178
rect 678 1173 679 1177
rect 683 1173 684 1177
rect 678 1172 684 1173
rect 710 1177 716 1178
rect 710 1173 711 1177
rect 715 1173 716 1177
rect 710 1172 716 1173
rect 742 1177 748 1178
rect 742 1173 743 1177
rect 747 1173 748 1177
rect 838 1176 839 1180
rect 843 1176 844 1180
rect 1694 1179 1700 1180
rect 1126 1177 1132 1178
rect 838 1175 844 1176
rect 1006 1176 1012 1177
rect 742 1172 748 1173
rect 774 1172 780 1173
rect 136 1151 138 1172
rect 168 1151 170 1172
rect 200 1151 202 1172
rect 232 1151 234 1172
rect 264 1151 266 1172
rect 296 1151 298 1172
rect 328 1151 330 1172
rect 360 1151 362 1172
rect 392 1151 394 1172
rect 424 1151 426 1172
rect 456 1151 458 1172
rect 488 1151 490 1172
rect 520 1151 522 1172
rect 552 1151 554 1172
rect 584 1151 586 1172
rect 616 1151 618 1172
rect 648 1151 650 1172
rect 680 1151 682 1172
rect 712 1151 714 1172
rect 744 1151 746 1172
rect 774 1168 775 1172
rect 779 1168 780 1172
rect 774 1167 780 1168
rect 776 1151 778 1167
rect 840 1151 842 1175
rect 1006 1172 1007 1176
rect 1011 1172 1012 1176
rect 1126 1173 1127 1177
rect 1131 1173 1132 1177
rect 1006 1171 1012 1172
rect 1086 1172 1092 1173
rect 1126 1172 1132 1173
rect 1158 1177 1164 1178
rect 1254 1177 1260 1178
rect 1158 1173 1159 1177
rect 1163 1173 1164 1177
rect 1158 1172 1164 1173
rect 1198 1176 1204 1177
rect 1198 1172 1199 1176
rect 1203 1172 1204 1176
rect 1254 1173 1255 1177
rect 1259 1173 1260 1177
rect 1254 1172 1260 1173
rect 1342 1177 1348 1178
rect 1342 1173 1343 1177
rect 1347 1173 1348 1177
rect 1342 1172 1348 1173
rect 1374 1177 1380 1178
rect 1374 1173 1375 1177
rect 1379 1173 1380 1177
rect 1374 1172 1380 1173
rect 1406 1177 1412 1178
rect 1406 1173 1407 1177
rect 1411 1173 1412 1177
rect 1406 1172 1412 1173
rect 1438 1177 1444 1178
rect 1438 1173 1439 1177
rect 1443 1173 1444 1177
rect 1438 1172 1444 1173
rect 1478 1177 1484 1178
rect 1478 1173 1479 1177
rect 1483 1173 1484 1177
rect 1478 1172 1484 1173
rect 1518 1177 1524 1178
rect 1518 1173 1519 1177
rect 1523 1173 1524 1177
rect 1518 1172 1524 1173
rect 1558 1177 1564 1178
rect 1558 1173 1559 1177
rect 1563 1173 1564 1177
rect 1558 1172 1564 1173
rect 1590 1177 1596 1178
rect 1590 1173 1591 1177
rect 1595 1173 1596 1177
rect 1590 1172 1596 1173
rect 1622 1177 1628 1178
rect 1622 1173 1623 1177
rect 1627 1173 1628 1177
rect 1622 1172 1628 1173
rect 1654 1177 1660 1178
rect 1654 1173 1655 1177
rect 1659 1173 1660 1177
rect 1694 1175 1695 1179
rect 1699 1175 1700 1179
rect 1694 1174 1700 1175
rect 1654 1172 1660 1173
rect 974 1170 980 1171
rect 974 1166 975 1170
rect 979 1166 980 1170
rect 974 1165 980 1166
rect 976 1151 978 1165
rect 1008 1151 1010 1171
rect 1086 1168 1087 1172
rect 1091 1168 1092 1172
rect 1086 1167 1092 1168
rect 1088 1151 1090 1167
rect 1128 1151 1130 1172
rect 1160 1151 1162 1172
rect 1198 1171 1204 1172
rect 1200 1151 1202 1171
rect 1256 1151 1258 1172
rect 1310 1170 1316 1171
rect 1310 1166 1311 1170
rect 1315 1166 1316 1170
rect 1310 1165 1316 1166
rect 1312 1151 1314 1165
rect 1344 1151 1346 1172
rect 1376 1151 1378 1172
rect 1408 1151 1410 1172
rect 1440 1151 1442 1172
rect 1480 1151 1482 1172
rect 1520 1151 1522 1172
rect 1560 1151 1562 1172
rect 1592 1151 1594 1172
rect 1624 1151 1626 1172
rect 1656 1151 1658 1172
rect 1696 1151 1698 1174
rect 111 1150 115 1151
rect 111 1145 115 1146
rect 135 1150 139 1151
rect 135 1145 139 1146
rect 167 1150 171 1151
rect 167 1145 171 1146
rect 199 1150 203 1151
rect 199 1145 203 1146
rect 231 1150 235 1151
rect 231 1145 235 1146
rect 263 1150 267 1151
rect 263 1145 267 1146
rect 295 1150 299 1151
rect 295 1145 299 1146
rect 327 1150 331 1151
rect 327 1145 331 1146
rect 359 1150 363 1151
rect 359 1145 363 1146
rect 391 1150 395 1151
rect 391 1145 395 1146
rect 423 1150 427 1151
rect 423 1145 427 1146
rect 455 1150 459 1151
rect 455 1145 459 1146
rect 487 1150 491 1151
rect 487 1145 491 1146
rect 519 1150 523 1151
rect 519 1145 523 1146
rect 551 1150 555 1151
rect 551 1145 555 1146
rect 583 1150 587 1151
rect 583 1145 587 1146
rect 615 1150 619 1151
rect 615 1145 619 1146
rect 647 1150 651 1151
rect 647 1145 651 1146
rect 679 1150 683 1151
rect 679 1145 683 1146
rect 687 1150 691 1151
rect 687 1145 691 1146
rect 711 1150 715 1151
rect 711 1145 715 1146
rect 743 1150 747 1151
rect 743 1145 747 1146
rect 775 1150 779 1151
rect 775 1145 779 1146
rect 799 1150 803 1151
rect 799 1145 803 1146
rect 839 1150 843 1151
rect 839 1145 843 1146
rect 847 1150 851 1151
rect 847 1145 851 1146
rect 935 1150 939 1151
rect 935 1145 939 1146
rect 967 1150 971 1151
rect 967 1145 971 1146
rect 975 1150 979 1151
rect 975 1145 979 1146
rect 999 1150 1003 1151
rect 999 1145 1003 1146
rect 1007 1150 1011 1151
rect 1007 1145 1011 1146
rect 1031 1150 1035 1151
rect 1031 1145 1035 1146
rect 1063 1150 1067 1151
rect 1063 1145 1067 1146
rect 1087 1150 1091 1151
rect 1087 1145 1091 1146
rect 1095 1150 1099 1151
rect 1095 1145 1099 1146
rect 1127 1150 1131 1151
rect 1127 1145 1131 1146
rect 1135 1150 1139 1151
rect 1135 1145 1139 1146
rect 1159 1150 1163 1151
rect 1159 1145 1163 1146
rect 1167 1150 1171 1151
rect 1167 1145 1171 1146
rect 1199 1150 1203 1151
rect 1199 1145 1203 1146
rect 1247 1150 1251 1151
rect 1247 1145 1251 1146
rect 1255 1150 1259 1151
rect 1255 1145 1259 1146
rect 1287 1150 1291 1151
rect 1287 1145 1291 1146
rect 1311 1150 1315 1151
rect 1311 1145 1315 1146
rect 1335 1150 1339 1151
rect 1335 1145 1339 1146
rect 1343 1150 1347 1151
rect 1343 1145 1347 1146
rect 1375 1150 1379 1151
rect 1375 1145 1379 1146
rect 1407 1150 1411 1151
rect 1407 1145 1411 1146
rect 1423 1150 1427 1151
rect 1423 1145 1427 1146
rect 1439 1150 1443 1151
rect 1439 1145 1443 1146
rect 1455 1150 1459 1151
rect 1455 1145 1459 1146
rect 1479 1150 1483 1151
rect 1479 1145 1483 1146
rect 1487 1150 1491 1151
rect 1487 1145 1491 1146
rect 1519 1150 1523 1151
rect 1519 1145 1523 1146
rect 1559 1150 1563 1151
rect 1559 1145 1563 1146
rect 1591 1150 1595 1151
rect 1591 1145 1595 1146
rect 1623 1150 1627 1151
rect 1623 1145 1627 1146
rect 1655 1150 1659 1151
rect 1655 1145 1659 1146
rect 1695 1150 1699 1151
rect 1695 1145 1699 1146
rect 112 1122 114 1145
rect 136 1124 138 1145
rect 168 1124 170 1145
rect 200 1124 202 1145
rect 232 1124 234 1145
rect 264 1124 266 1145
rect 296 1124 298 1145
rect 328 1124 330 1145
rect 360 1124 362 1145
rect 392 1124 394 1145
rect 424 1124 426 1145
rect 456 1124 458 1145
rect 488 1124 490 1145
rect 520 1124 522 1145
rect 552 1124 554 1145
rect 584 1125 586 1145
rect 582 1124 588 1125
rect 134 1123 140 1124
rect 110 1121 116 1122
rect 110 1117 111 1121
rect 115 1117 116 1121
rect 134 1119 135 1123
rect 139 1119 140 1123
rect 134 1118 140 1119
rect 166 1123 172 1124
rect 166 1119 167 1123
rect 171 1119 172 1123
rect 166 1118 172 1119
rect 198 1123 204 1124
rect 198 1119 199 1123
rect 203 1119 204 1123
rect 198 1118 204 1119
rect 230 1123 236 1124
rect 230 1119 231 1123
rect 235 1119 236 1123
rect 230 1118 236 1119
rect 262 1123 268 1124
rect 262 1119 263 1123
rect 267 1119 268 1123
rect 262 1118 268 1119
rect 294 1123 300 1124
rect 294 1119 295 1123
rect 299 1119 300 1123
rect 294 1118 300 1119
rect 326 1123 332 1124
rect 326 1119 327 1123
rect 331 1119 332 1123
rect 326 1118 332 1119
rect 358 1123 364 1124
rect 358 1119 359 1123
rect 363 1119 364 1123
rect 358 1118 364 1119
rect 390 1123 396 1124
rect 390 1119 391 1123
rect 395 1119 396 1123
rect 390 1118 396 1119
rect 422 1123 428 1124
rect 422 1119 423 1123
rect 427 1119 428 1123
rect 422 1118 428 1119
rect 454 1123 460 1124
rect 454 1119 455 1123
rect 459 1119 460 1123
rect 454 1118 460 1119
rect 486 1123 492 1124
rect 486 1119 487 1123
rect 491 1119 492 1123
rect 486 1118 492 1119
rect 518 1123 524 1124
rect 518 1119 519 1123
rect 523 1119 524 1123
rect 518 1118 524 1119
rect 550 1123 556 1124
rect 550 1119 551 1123
rect 555 1119 556 1123
rect 582 1120 583 1124
rect 587 1120 588 1124
rect 688 1121 690 1145
rect 800 1125 802 1145
rect 848 1127 850 1145
rect 846 1126 852 1127
rect 798 1124 804 1125
rect 582 1119 588 1120
rect 686 1120 692 1121
rect 550 1118 556 1119
rect 110 1116 116 1117
rect 686 1116 687 1120
rect 691 1116 692 1120
rect 798 1120 799 1124
rect 803 1120 804 1124
rect 846 1122 847 1126
rect 851 1122 852 1126
rect 936 1124 938 1145
rect 968 1124 970 1145
rect 1000 1125 1002 1145
rect 998 1124 1004 1125
rect 1032 1124 1034 1145
rect 1064 1124 1066 1145
rect 1096 1125 1098 1145
rect 1094 1124 1100 1125
rect 1136 1124 1138 1145
rect 1168 1125 1170 1145
rect 1248 1129 1250 1145
rect 1246 1128 1252 1129
rect 1166 1124 1172 1125
rect 846 1121 852 1122
rect 934 1123 940 1124
rect 798 1119 804 1120
rect 934 1119 935 1123
rect 939 1119 940 1123
rect 934 1118 940 1119
rect 966 1123 972 1124
rect 966 1119 967 1123
rect 971 1119 972 1123
rect 998 1120 999 1124
rect 1003 1120 1004 1124
rect 998 1119 1004 1120
rect 1030 1123 1036 1124
rect 1030 1119 1031 1123
rect 1035 1119 1036 1123
rect 966 1118 972 1119
rect 1030 1118 1036 1119
rect 1062 1123 1068 1124
rect 1062 1119 1063 1123
rect 1067 1119 1068 1123
rect 1094 1120 1095 1124
rect 1099 1120 1100 1124
rect 1094 1119 1100 1120
rect 1134 1123 1140 1124
rect 1134 1119 1135 1123
rect 1139 1119 1140 1123
rect 1166 1120 1167 1124
rect 1171 1120 1172 1124
rect 1246 1124 1247 1128
rect 1251 1124 1252 1128
rect 1288 1124 1290 1145
rect 1336 1127 1338 1145
rect 1334 1126 1340 1127
rect 1246 1123 1252 1124
rect 1286 1123 1292 1124
rect 1166 1119 1172 1120
rect 1286 1119 1287 1123
rect 1291 1119 1292 1123
rect 1334 1122 1335 1126
rect 1339 1122 1340 1126
rect 1424 1124 1426 1145
rect 1456 1124 1458 1145
rect 1488 1124 1490 1145
rect 1520 1124 1522 1145
rect 1560 1124 1562 1145
rect 1592 1124 1594 1145
rect 1624 1124 1626 1145
rect 1656 1124 1658 1145
rect 1334 1121 1340 1122
rect 1422 1123 1428 1124
rect 1062 1118 1068 1119
rect 1134 1118 1140 1119
rect 1286 1118 1292 1119
rect 1422 1119 1423 1123
rect 1427 1119 1428 1123
rect 1422 1118 1428 1119
rect 1454 1123 1460 1124
rect 1454 1119 1455 1123
rect 1459 1119 1460 1123
rect 1454 1118 1460 1119
rect 1486 1123 1492 1124
rect 1486 1119 1487 1123
rect 1491 1119 1492 1123
rect 1486 1118 1492 1119
rect 1518 1123 1524 1124
rect 1518 1119 1519 1123
rect 1523 1119 1524 1123
rect 1518 1118 1524 1119
rect 1558 1123 1564 1124
rect 1558 1119 1559 1123
rect 1563 1119 1564 1123
rect 1558 1118 1564 1119
rect 1590 1123 1596 1124
rect 1590 1119 1591 1123
rect 1595 1119 1596 1123
rect 1590 1118 1596 1119
rect 1622 1123 1628 1124
rect 1622 1119 1623 1123
rect 1627 1119 1628 1123
rect 1622 1118 1628 1119
rect 1654 1123 1660 1124
rect 1654 1119 1655 1123
rect 1659 1119 1660 1123
rect 1696 1122 1698 1145
rect 1654 1118 1660 1119
rect 1694 1121 1700 1122
rect 1694 1117 1695 1121
rect 1699 1117 1700 1121
rect 1694 1116 1700 1117
rect 686 1115 692 1116
rect 134 1106 140 1107
rect 110 1104 116 1105
rect 110 1100 111 1104
rect 115 1100 116 1104
rect 134 1102 135 1106
rect 139 1102 140 1106
rect 134 1101 140 1102
rect 166 1106 172 1107
rect 166 1102 167 1106
rect 171 1102 172 1106
rect 166 1101 172 1102
rect 198 1106 204 1107
rect 198 1102 199 1106
rect 203 1102 204 1106
rect 198 1101 204 1102
rect 230 1106 236 1107
rect 230 1102 231 1106
rect 235 1102 236 1106
rect 230 1101 236 1102
rect 262 1106 268 1107
rect 262 1102 263 1106
rect 267 1102 268 1106
rect 262 1101 268 1102
rect 294 1106 300 1107
rect 294 1102 295 1106
rect 299 1102 300 1106
rect 294 1101 300 1102
rect 326 1106 332 1107
rect 326 1102 327 1106
rect 331 1102 332 1106
rect 326 1101 332 1102
rect 358 1106 364 1107
rect 358 1102 359 1106
rect 363 1102 364 1106
rect 358 1101 364 1102
rect 390 1106 396 1107
rect 390 1102 391 1106
rect 395 1102 396 1106
rect 390 1101 396 1102
rect 422 1106 428 1107
rect 422 1102 423 1106
rect 427 1102 428 1106
rect 422 1101 428 1102
rect 454 1106 460 1107
rect 454 1102 455 1106
rect 459 1102 460 1106
rect 454 1101 460 1102
rect 486 1106 492 1107
rect 486 1102 487 1106
rect 491 1102 492 1106
rect 486 1101 492 1102
rect 518 1106 524 1107
rect 518 1102 519 1106
rect 523 1102 524 1106
rect 518 1101 524 1102
rect 550 1106 556 1107
rect 934 1106 940 1107
rect 550 1102 551 1106
rect 555 1102 556 1106
rect 550 1101 556 1102
rect 658 1105 664 1106
rect 658 1101 659 1105
rect 663 1101 664 1105
rect 934 1102 935 1106
rect 939 1102 940 1106
rect 110 1099 116 1100
rect 112 1035 114 1099
rect 136 1035 138 1101
rect 168 1035 170 1101
rect 200 1035 202 1101
rect 232 1035 234 1101
rect 264 1035 266 1101
rect 296 1035 298 1101
rect 328 1035 330 1101
rect 360 1035 362 1101
rect 392 1035 394 1101
rect 424 1035 426 1101
rect 456 1035 458 1101
rect 488 1035 490 1101
rect 520 1035 522 1101
rect 552 1035 554 1101
rect 658 1100 664 1101
rect 798 1101 804 1102
rect 934 1101 940 1102
rect 966 1106 972 1107
rect 966 1102 967 1106
rect 971 1102 972 1106
rect 1030 1106 1036 1107
rect 1030 1102 1031 1106
rect 1035 1102 1036 1106
rect 966 1101 972 1102
rect 998 1101 1004 1102
rect 1030 1101 1036 1102
rect 1062 1106 1068 1107
rect 1062 1102 1063 1106
rect 1067 1102 1068 1106
rect 1062 1101 1068 1102
rect 1134 1106 1140 1107
rect 1134 1102 1135 1106
rect 1139 1102 1140 1106
rect 1134 1101 1140 1102
rect 1286 1106 1292 1107
rect 1286 1102 1287 1106
rect 1291 1102 1292 1106
rect 1286 1101 1292 1102
rect 1422 1106 1428 1107
rect 1422 1102 1423 1106
rect 1427 1102 1428 1106
rect 1422 1101 1428 1102
rect 1454 1106 1460 1107
rect 1454 1102 1455 1106
rect 1459 1102 1460 1106
rect 1454 1101 1460 1102
rect 1486 1106 1492 1107
rect 1486 1102 1487 1106
rect 1491 1102 1492 1106
rect 1486 1101 1492 1102
rect 1518 1106 1524 1107
rect 1518 1102 1519 1106
rect 1523 1102 1524 1106
rect 1518 1101 1524 1102
rect 1558 1106 1564 1107
rect 1558 1102 1559 1106
rect 1563 1102 1564 1106
rect 1558 1101 1564 1102
rect 1590 1106 1596 1107
rect 1590 1102 1591 1106
rect 1595 1102 1596 1106
rect 1590 1101 1596 1102
rect 1622 1106 1628 1107
rect 1622 1102 1623 1106
rect 1627 1102 1628 1106
rect 1622 1101 1628 1102
rect 1654 1106 1660 1107
rect 1654 1102 1655 1106
rect 1659 1102 1660 1106
rect 1654 1101 1660 1102
rect 1694 1104 1700 1105
rect 590 1086 596 1087
rect 590 1082 591 1086
rect 595 1082 596 1086
rect 590 1081 596 1082
rect 592 1035 594 1081
rect 660 1035 662 1100
rect 798 1097 799 1101
rect 803 1097 804 1101
rect 798 1096 804 1097
rect 800 1035 802 1096
rect 846 1085 852 1086
rect 846 1081 847 1085
rect 851 1081 852 1085
rect 846 1080 852 1081
rect 848 1035 850 1080
rect 936 1035 938 1101
rect 968 1035 970 1101
rect 998 1097 999 1101
rect 1003 1097 1004 1101
rect 998 1096 1004 1097
rect 1000 1035 1002 1096
rect 1032 1035 1034 1101
rect 1064 1035 1066 1101
rect 1094 1096 1100 1097
rect 1094 1092 1095 1096
rect 1099 1092 1100 1096
rect 1094 1091 1100 1092
rect 1096 1035 1098 1091
rect 1136 1035 1138 1101
rect 1174 1086 1180 1087
rect 1174 1082 1175 1086
rect 1179 1082 1180 1086
rect 1174 1081 1180 1082
rect 1246 1081 1252 1082
rect 1176 1035 1178 1081
rect 1246 1077 1247 1081
rect 1251 1077 1252 1081
rect 1246 1076 1252 1077
rect 1248 1035 1250 1076
rect 1288 1035 1290 1101
rect 1334 1085 1340 1086
rect 1334 1081 1335 1085
rect 1339 1081 1340 1085
rect 1334 1080 1340 1081
rect 1336 1035 1338 1080
rect 1424 1035 1426 1101
rect 1456 1035 1458 1101
rect 1488 1035 1490 1101
rect 1520 1035 1522 1101
rect 1560 1035 1562 1101
rect 1592 1035 1594 1101
rect 1624 1035 1626 1101
rect 1656 1035 1658 1101
rect 1694 1100 1695 1104
rect 1699 1100 1700 1104
rect 1694 1099 1700 1100
rect 1696 1035 1698 1099
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 135 1034 139 1035
rect 135 1029 139 1030
rect 167 1034 171 1035
rect 167 1029 171 1030
rect 199 1034 203 1035
rect 199 1029 203 1030
rect 231 1034 235 1035
rect 231 1029 235 1030
rect 263 1034 267 1035
rect 263 1029 267 1030
rect 295 1034 299 1035
rect 295 1029 299 1030
rect 327 1034 331 1035
rect 327 1029 331 1030
rect 359 1034 363 1035
rect 359 1029 363 1030
rect 391 1034 395 1035
rect 391 1029 395 1030
rect 407 1034 411 1035
rect 407 1029 411 1030
rect 423 1034 427 1035
rect 423 1029 427 1030
rect 455 1034 459 1035
rect 455 1029 459 1030
rect 487 1034 491 1035
rect 487 1029 491 1030
rect 503 1034 507 1035
rect 503 1029 507 1030
rect 519 1034 523 1035
rect 519 1029 523 1030
rect 551 1034 555 1035
rect 551 1029 555 1030
rect 583 1034 587 1035
rect 583 1029 587 1030
rect 591 1034 595 1035
rect 591 1029 595 1030
rect 659 1034 663 1035
rect 659 1029 663 1030
rect 711 1034 715 1035
rect 711 1029 715 1030
rect 799 1034 803 1035
rect 799 1029 803 1030
rect 823 1034 827 1035
rect 823 1029 827 1030
rect 847 1034 851 1035
rect 847 1029 851 1030
rect 919 1034 923 1035
rect 919 1029 923 1030
rect 935 1034 939 1035
rect 935 1029 939 1030
rect 967 1034 971 1035
rect 967 1029 971 1030
rect 975 1034 979 1035
rect 975 1029 979 1030
rect 999 1034 1003 1035
rect 999 1029 1003 1030
rect 1031 1034 1035 1035
rect 1031 1029 1035 1030
rect 1063 1034 1067 1035
rect 1063 1029 1067 1030
rect 1095 1034 1099 1035
rect 1095 1029 1099 1030
rect 1119 1034 1123 1035
rect 1119 1029 1123 1030
rect 1135 1034 1139 1035
rect 1135 1029 1139 1030
rect 1167 1034 1171 1035
rect 1167 1029 1171 1030
rect 1175 1034 1179 1035
rect 1175 1029 1179 1030
rect 1199 1034 1203 1035
rect 1199 1029 1203 1030
rect 1247 1034 1251 1035
rect 1247 1029 1251 1030
rect 1287 1034 1291 1035
rect 1287 1029 1291 1030
rect 1295 1034 1299 1035
rect 1295 1029 1299 1030
rect 1327 1034 1331 1035
rect 1327 1029 1331 1030
rect 1335 1034 1339 1035
rect 1335 1029 1339 1030
rect 1367 1034 1371 1035
rect 1367 1029 1371 1030
rect 1407 1034 1411 1035
rect 1407 1029 1411 1030
rect 1423 1034 1427 1035
rect 1423 1029 1427 1030
rect 1439 1034 1443 1035
rect 1439 1029 1443 1030
rect 1455 1034 1459 1035
rect 1455 1029 1459 1030
rect 1479 1034 1483 1035
rect 1479 1029 1483 1030
rect 1487 1034 1491 1035
rect 1487 1029 1491 1030
rect 1519 1034 1523 1035
rect 1519 1029 1523 1030
rect 1559 1034 1563 1035
rect 1559 1029 1563 1030
rect 1591 1034 1595 1035
rect 1591 1029 1595 1030
rect 1623 1034 1627 1035
rect 1623 1029 1627 1030
rect 1655 1034 1659 1035
rect 1655 1029 1659 1030
rect 1695 1034 1699 1035
rect 1695 1029 1699 1030
rect 112 997 114 1029
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 136 995 138 1029
rect 168 995 170 1029
rect 200 995 202 1029
rect 232 995 234 1029
rect 264 995 266 1029
rect 328 998 330 1029
rect 408 1015 410 1029
rect 504 1020 506 1029
rect 502 1019 508 1020
rect 502 1015 503 1019
rect 507 1015 508 1019
rect 584 1016 586 1029
rect 712 1016 714 1029
rect 406 1014 412 1015
rect 502 1014 508 1015
rect 582 1015 588 1016
rect 406 1010 407 1014
rect 411 1010 412 1014
rect 582 1011 583 1015
rect 587 1011 588 1015
rect 582 1010 588 1011
rect 710 1015 716 1016
rect 710 1011 711 1015
rect 715 1011 716 1015
rect 710 1010 716 1011
rect 824 1010 826 1029
rect 406 1009 412 1010
rect 822 1009 828 1010
rect 822 1005 823 1009
rect 827 1005 828 1009
rect 822 1004 828 1005
rect 326 997 332 998
rect 110 991 116 992
rect 134 994 140 995
rect 134 990 135 994
rect 139 990 140 994
rect 134 989 140 990
rect 166 994 172 995
rect 166 990 167 994
rect 171 990 172 994
rect 166 989 172 990
rect 198 994 204 995
rect 198 990 199 994
rect 203 990 204 994
rect 198 989 204 990
rect 230 994 236 995
rect 230 990 231 994
rect 235 990 236 994
rect 230 989 236 990
rect 262 994 268 995
rect 262 990 263 994
rect 267 990 268 994
rect 326 993 327 997
rect 331 993 332 997
rect 920 995 922 1029
rect 976 1010 978 1029
rect 974 1009 980 1010
rect 974 1005 975 1009
rect 979 1005 980 1009
rect 1064 1005 1066 1029
rect 974 1004 980 1005
rect 1062 1004 1068 1005
rect 1062 1000 1063 1004
rect 1067 1000 1068 1004
rect 1062 999 1068 1000
rect 1120 998 1122 1029
rect 1118 997 1124 998
rect 326 992 332 993
rect 918 994 924 995
rect 262 989 268 990
rect 918 990 919 994
rect 923 990 924 994
rect 1118 993 1119 997
rect 1123 993 1124 997
rect 1168 995 1170 1029
rect 1200 1005 1202 1029
rect 1198 1004 1204 1005
rect 1198 1000 1199 1004
rect 1203 1000 1204 1004
rect 1198 999 1204 1000
rect 1248 998 1250 1029
rect 1246 997 1252 998
rect 1118 992 1124 993
rect 1166 994 1172 995
rect 918 989 924 990
rect 1166 990 1167 994
rect 1171 990 1172 994
rect 1246 993 1247 997
rect 1251 993 1252 997
rect 1296 995 1298 1029
rect 1328 1005 1330 1029
rect 1368 1005 1370 1029
rect 1326 1004 1332 1005
rect 1326 1000 1327 1004
rect 1331 1000 1332 1004
rect 1326 999 1332 1000
rect 1366 1004 1372 1005
rect 1366 1000 1367 1004
rect 1371 1000 1372 1004
rect 1366 999 1372 1000
rect 1408 995 1410 1029
rect 1440 995 1442 1029
rect 1480 995 1482 1029
rect 1520 995 1522 1029
rect 1560 995 1562 1029
rect 1592 995 1594 1029
rect 1624 995 1626 1029
rect 1656 995 1658 1029
rect 1696 997 1698 1029
rect 1694 996 1700 997
rect 1246 992 1252 993
rect 1294 994 1300 995
rect 1166 989 1172 990
rect 1294 990 1295 994
rect 1299 990 1300 994
rect 1294 989 1300 990
rect 1406 994 1412 995
rect 1406 990 1407 994
rect 1411 990 1412 994
rect 1406 989 1412 990
rect 1438 994 1444 995
rect 1438 990 1439 994
rect 1443 990 1444 994
rect 1438 989 1444 990
rect 1478 994 1484 995
rect 1478 990 1479 994
rect 1483 990 1484 994
rect 1478 989 1484 990
rect 1518 994 1524 995
rect 1518 990 1519 994
rect 1523 990 1524 994
rect 1518 989 1524 990
rect 1558 994 1564 995
rect 1558 990 1559 994
rect 1563 990 1564 994
rect 1558 989 1564 990
rect 1590 994 1596 995
rect 1590 990 1591 994
rect 1595 990 1596 994
rect 1590 989 1596 990
rect 1622 994 1628 995
rect 1622 990 1623 994
rect 1627 990 1628 994
rect 1622 989 1628 990
rect 1654 994 1660 995
rect 1654 990 1655 994
rect 1659 990 1660 994
rect 1694 992 1695 996
rect 1699 992 1700 996
rect 1694 991 1700 992
rect 1654 989 1660 990
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 1694 979 1700 980
rect 110 974 116 975
rect 134 977 140 978
rect 112 955 114 974
rect 134 973 135 977
rect 139 973 140 977
rect 134 972 140 973
rect 166 977 172 978
rect 166 973 167 977
rect 171 973 172 977
rect 166 972 172 973
rect 198 977 204 978
rect 198 973 199 977
rect 203 973 204 977
rect 198 972 204 973
rect 230 977 236 978
rect 230 973 231 977
rect 235 973 236 977
rect 230 972 236 973
rect 262 977 268 978
rect 918 977 924 978
rect 1166 977 1172 978
rect 1294 977 1300 978
rect 1406 977 1412 978
rect 262 973 263 977
rect 267 973 268 977
rect 262 972 268 973
rect 398 976 404 977
rect 398 972 399 976
rect 403 972 404 976
rect 582 974 588 975
rect 136 955 138 972
rect 168 955 170 972
rect 200 955 202 972
rect 232 955 234 972
rect 264 955 266 972
rect 398 971 404 972
rect 502 972 508 973
rect 342 970 348 971
rect 342 966 343 970
rect 347 966 348 970
rect 342 965 348 966
rect 344 955 346 965
rect 400 955 402 971
rect 502 968 503 972
rect 507 968 508 972
rect 582 970 583 974
rect 587 970 588 974
rect 582 969 588 970
rect 710 974 716 975
rect 710 970 711 974
rect 715 970 716 974
rect 918 973 919 977
rect 923 973 924 977
rect 918 972 924 973
rect 1062 976 1068 977
rect 1062 972 1063 976
rect 1067 972 1068 976
rect 1166 973 1167 977
rect 1171 973 1172 977
rect 1166 972 1172 973
rect 1198 976 1204 977
rect 1198 972 1199 976
rect 1203 972 1204 976
rect 1294 973 1295 977
rect 1299 973 1300 977
rect 1294 972 1300 973
rect 1326 976 1332 977
rect 1326 972 1327 976
rect 1331 972 1332 976
rect 710 969 716 970
rect 814 969 820 970
rect 502 967 508 968
rect 504 955 506 967
rect 584 955 586 969
rect 712 955 714 969
rect 814 965 815 969
rect 819 965 820 969
rect 814 964 820 965
rect 816 955 818 964
rect 920 955 922 972
rect 1062 971 1068 972
rect 966 969 972 970
rect 966 965 967 969
rect 971 965 972 969
rect 966 964 972 965
rect 968 955 970 964
rect 1064 955 1066 971
rect 1134 970 1140 971
rect 1134 966 1135 970
rect 1139 966 1140 970
rect 1134 965 1140 966
rect 1136 955 1138 965
rect 1168 955 1170 972
rect 1198 971 1204 972
rect 1200 955 1202 971
rect 1262 970 1268 971
rect 1262 966 1263 970
rect 1267 966 1268 970
rect 1262 965 1268 966
rect 1264 955 1266 965
rect 1296 955 1298 972
rect 1326 971 1332 972
rect 1366 976 1372 977
rect 1366 972 1367 976
rect 1371 972 1372 976
rect 1406 973 1407 977
rect 1411 973 1412 977
rect 1406 972 1412 973
rect 1438 977 1444 978
rect 1438 973 1439 977
rect 1443 973 1444 977
rect 1438 972 1444 973
rect 1478 977 1484 978
rect 1478 973 1479 977
rect 1483 973 1484 977
rect 1478 972 1484 973
rect 1518 977 1524 978
rect 1518 973 1519 977
rect 1523 973 1524 977
rect 1518 972 1524 973
rect 1558 977 1564 978
rect 1558 973 1559 977
rect 1563 973 1564 977
rect 1558 972 1564 973
rect 1590 977 1596 978
rect 1590 973 1591 977
rect 1595 973 1596 977
rect 1590 972 1596 973
rect 1622 977 1628 978
rect 1622 973 1623 977
rect 1627 973 1628 977
rect 1622 972 1628 973
rect 1654 977 1660 978
rect 1654 973 1655 977
rect 1659 973 1660 977
rect 1694 975 1695 979
rect 1699 975 1700 979
rect 1694 974 1700 975
rect 1654 972 1660 973
rect 1366 971 1372 972
rect 1328 955 1330 971
rect 1368 955 1370 971
rect 1408 955 1410 972
rect 1440 955 1442 972
rect 1480 955 1482 972
rect 1520 955 1522 972
rect 1560 955 1562 972
rect 1592 955 1594 972
rect 1624 955 1626 972
rect 1656 955 1658 972
rect 1696 955 1698 974
rect 111 954 115 955
rect 111 949 115 950
rect 135 954 139 955
rect 135 949 139 950
rect 167 954 171 955
rect 167 949 171 950
rect 199 954 203 955
rect 199 949 203 950
rect 231 954 235 955
rect 231 949 235 950
rect 263 954 267 955
rect 263 949 267 950
rect 279 954 283 955
rect 279 949 283 950
rect 319 954 323 955
rect 319 949 323 950
rect 343 954 347 955
rect 343 949 347 950
rect 399 954 403 955
rect 399 949 403 950
rect 463 954 467 955
rect 463 949 467 950
rect 503 954 507 955
rect 503 949 507 950
rect 583 954 587 955
rect 583 949 587 950
rect 591 954 595 955
rect 591 949 595 950
rect 679 954 683 955
rect 679 949 683 950
rect 711 954 715 955
rect 711 949 715 950
rect 727 954 731 955
rect 727 949 731 950
rect 815 954 819 955
rect 815 949 819 950
rect 863 954 867 955
rect 863 949 867 950
rect 919 954 923 955
rect 919 949 923 950
rect 951 954 955 955
rect 951 949 955 950
rect 967 954 971 955
rect 967 949 971 950
rect 983 954 987 955
rect 983 949 987 950
rect 1039 954 1043 955
rect 1039 949 1043 950
rect 1063 954 1067 955
rect 1063 949 1067 950
rect 1071 954 1075 955
rect 1071 949 1075 950
rect 1111 954 1115 955
rect 1111 949 1115 950
rect 1135 954 1139 955
rect 1135 949 1139 950
rect 1143 954 1147 955
rect 1143 949 1147 950
rect 1167 954 1171 955
rect 1167 949 1171 950
rect 1199 954 1203 955
rect 1199 949 1203 950
rect 1239 954 1243 955
rect 1239 949 1243 950
rect 1263 954 1267 955
rect 1263 949 1267 950
rect 1271 954 1275 955
rect 1271 949 1275 950
rect 1295 954 1299 955
rect 1295 949 1299 950
rect 1327 954 1331 955
rect 1327 949 1331 950
rect 1367 954 1371 955
rect 1367 949 1371 950
rect 1391 954 1395 955
rect 1391 949 1395 950
rect 1407 954 1411 955
rect 1407 949 1411 950
rect 1423 954 1427 955
rect 1423 949 1427 950
rect 1439 954 1443 955
rect 1439 949 1443 950
rect 1455 954 1459 955
rect 1455 949 1459 950
rect 1479 954 1483 955
rect 1479 949 1483 950
rect 1519 954 1523 955
rect 1519 949 1523 950
rect 1559 954 1563 955
rect 1559 949 1563 950
rect 1591 954 1595 955
rect 1591 949 1595 950
rect 1623 954 1627 955
rect 1623 949 1627 950
rect 1655 954 1659 955
rect 1655 949 1659 950
rect 1695 954 1699 955
rect 1695 949 1699 950
rect 112 922 114 949
rect 136 924 138 949
rect 168 924 170 949
rect 200 925 202 949
rect 280 929 282 949
rect 278 928 284 929
rect 198 924 204 925
rect 134 923 140 924
rect 110 921 116 922
rect 110 917 111 921
rect 115 917 116 921
rect 134 919 135 923
rect 139 919 140 923
rect 134 918 140 919
rect 166 923 172 924
rect 166 919 167 923
rect 171 919 172 923
rect 198 920 199 924
rect 203 920 204 924
rect 278 924 279 928
rect 283 924 284 928
rect 320 925 322 949
rect 400 929 402 949
rect 398 928 404 929
rect 278 923 284 924
rect 318 924 324 925
rect 198 919 204 920
rect 318 920 319 924
rect 323 920 324 924
rect 398 924 399 928
rect 403 924 404 928
rect 398 923 404 924
rect 464 921 466 949
rect 592 927 594 949
rect 590 926 596 927
rect 590 922 591 926
rect 595 922 596 926
rect 680 925 682 949
rect 728 927 730 949
rect 726 926 732 927
rect 590 921 596 922
rect 678 924 684 925
rect 318 919 324 920
rect 462 920 468 921
rect 166 918 172 919
rect 110 916 116 917
rect 462 916 463 920
rect 467 916 468 920
rect 678 920 679 924
rect 683 920 684 924
rect 726 922 727 926
rect 731 922 732 926
rect 816 924 818 949
rect 864 927 866 949
rect 862 926 868 927
rect 726 921 732 922
rect 814 923 820 924
rect 678 919 684 920
rect 814 919 815 923
rect 819 919 820 923
rect 862 922 863 926
rect 867 922 868 926
rect 952 924 954 949
rect 984 925 986 949
rect 982 924 988 925
rect 1040 924 1042 949
rect 1072 925 1074 949
rect 1070 924 1076 925
rect 1112 924 1114 949
rect 1144 925 1146 949
rect 1142 924 1148 925
rect 1240 924 1242 949
rect 1272 925 1274 949
rect 1392 931 1394 949
rect 1390 930 1396 931
rect 1390 926 1391 930
rect 1395 926 1396 930
rect 1390 925 1396 926
rect 1270 924 1276 925
rect 1424 924 1426 949
rect 1456 925 1458 949
rect 1454 924 1460 925
rect 1520 924 1522 949
rect 1560 924 1562 949
rect 1592 924 1594 949
rect 1624 924 1626 949
rect 1656 924 1658 949
rect 862 921 868 922
rect 950 923 956 924
rect 814 918 820 919
rect 950 919 951 923
rect 955 919 956 923
rect 982 920 983 924
rect 987 920 988 924
rect 982 919 988 920
rect 1038 923 1044 924
rect 1038 919 1039 923
rect 1043 919 1044 923
rect 1070 920 1071 924
rect 1075 920 1076 924
rect 1070 919 1076 920
rect 1110 923 1116 924
rect 1110 919 1111 923
rect 1115 919 1116 923
rect 1142 920 1143 924
rect 1147 920 1148 924
rect 1142 919 1148 920
rect 1238 923 1244 924
rect 1238 919 1239 923
rect 1243 919 1244 923
rect 1270 920 1271 924
rect 1275 920 1276 924
rect 1270 919 1276 920
rect 1422 923 1428 924
rect 1422 919 1423 923
rect 1427 919 1428 923
rect 1454 920 1455 924
rect 1459 920 1460 924
rect 1454 919 1460 920
rect 1518 923 1524 924
rect 1518 919 1519 923
rect 1523 919 1524 923
rect 950 918 956 919
rect 1038 918 1044 919
rect 1110 918 1116 919
rect 1238 918 1244 919
rect 1422 918 1428 919
rect 1518 918 1524 919
rect 1558 923 1564 924
rect 1558 919 1559 923
rect 1563 919 1564 923
rect 1558 918 1564 919
rect 1590 923 1596 924
rect 1590 919 1591 923
rect 1595 919 1596 923
rect 1590 918 1596 919
rect 1622 923 1628 924
rect 1622 919 1623 923
rect 1627 919 1628 923
rect 1622 918 1628 919
rect 1654 923 1660 924
rect 1654 919 1655 923
rect 1659 919 1660 923
rect 1696 922 1698 949
rect 1654 918 1660 919
rect 1694 921 1700 922
rect 1694 917 1695 921
rect 1699 917 1700 921
rect 1694 916 1700 917
rect 462 915 468 916
rect 134 906 140 907
rect 110 904 116 905
rect 110 900 111 904
rect 115 900 116 904
rect 134 902 135 906
rect 139 902 140 906
rect 134 901 140 902
rect 166 906 172 907
rect 814 906 820 907
rect 166 902 167 906
rect 171 902 172 906
rect 166 901 172 902
rect 434 905 440 906
rect 434 901 435 905
rect 439 901 440 905
rect 814 902 815 906
rect 819 902 820 906
rect 110 899 116 900
rect 112 839 114 899
rect 136 839 138 901
rect 168 839 170 901
rect 434 900 440 901
rect 678 901 684 902
rect 814 901 820 902
rect 950 906 956 907
rect 950 902 951 906
rect 955 902 956 906
rect 1038 906 1044 907
rect 1422 906 1428 907
rect 950 901 956 902
rect 998 903 1004 904
rect 206 886 212 887
rect 206 882 207 886
rect 211 882 212 886
rect 326 886 332 887
rect 326 882 327 886
rect 331 882 332 886
rect 206 881 212 882
rect 278 881 284 882
rect 326 881 332 882
rect 398 881 404 882
rect 208 839 210 881
rect 278 877 279 881
rect 283 877 284 881
rect 278 876 284 877
rect 280 839 282 876
rect 328 839 330 881
rect 398 877 399 881
rect 403 877 404 881
rect 398 876 404 877
rect 400 839 402 876
rect 436 839 438 900
rect 678 897 679 901
rect 683 897 684 901
rect 678 896 684 897
rect 590 885 596 886
rect 590 881 591 885
rect 595 881 596 885
rect 590 880 596 881
rect 592 839 594 880
rect 680 839 682 896
rect 726 885 732 886
rect 726 881 727 885
rect 731 881 732 885
rect 726 880 732 881
rect 728 839 730 880
rect 816 839 818 901
rect 862 885 868 886
rect 862 881 863 885
rect 867 881 868 885
rect 862 880 868 881
rect 864 839 866 880
rect 952 839 954 901
rect 998 899 999 903
rect 1003 899 1004 903
rect 1038 902 1039 906
rect 1043 902 1044 906
rect 1038 901 1044 902
rect 1110 905 1116 906
rect 1110 901 1111 905
rect 1115 901 1116 905
rect 998 898 1004 899
rect 1000 839 1002 898
rect 1040 839 1042 901
rect 1110 900 1116 901
rect 1142 905 1148 906
rect 1142 901 1143 905
rect 1147 901 1148 905
rect 1142 900 1148 901
rect 1238 905 1244 906
rect 1238 901 1239 905
rect 1243 901 1244 905
rect 1238 900 1244 901
rect 1270 905 1276 906
rect 1270 901 1271 905
rect 1275 901 1276 905
rect 1270 900 1276 901
rect 1374 903 1380 904
rect 1070 896 1076 897
rect 1070 892 1071 896
rect 1075 892 1076 896
rect 1070 891 1076 892
rect 1072 839 1074 891
rect 1112 839 1114 900
rect 1144 839 1146 900
rect 1240 839 1242 900
rect 1272 839 1274 900
rect 1374 899 1375 903
rect 1379 899 1380 903
rect 1422 902 1423 906
rect 1427 902 1428 906
rect 1518 906 1524 907
rect 1422 901 1428 902
rect 1470 903 1476 904
rect 1374 898 1380 899
rect 1376 839 1378 898
rect 1424 839 1426 901
rect 1470 899 1471 903
rect 1475 899 1476 903
rect 1518 902 1519 906
rect 1523 902 1524 906
rect 1518 901 1524 902
rect 1558 906 1564 907
rect 1558 902 1559 906
rect 1563 902 1564 906
rect 1558 901 1564 902
rect 1590 906 1596 907
rect 1590 902 1591 906
rect 1595 902 1596 906
rect 1590 901 1596 902
rect 1622 906 1628 907
rect 1622 902 1623 906
rect 1627 902 1628 906
rect 1622 901 1628 902
rect 1654 906 1660 907
rect 1654 902 1655 906
rect 1659 902 1660 906
rect 1654 901 1660 902
rect 1694 904 1700 905
rect 1470 898 1476 899
rect 1472 839 1474 898
rect 1520 839 1522 901
rect 1560 839 1562 901
rect 1592 839 1594 901
rect 1624 839 1626 901
rect 1656 839 1658 901
rect 1694 900 1695 904
rect 1699 900 1700 904
rect 1694 899 1700 900
rect 1696 839 1698 899
rect 111 838 115 839
rect 111 833 115 834
rect 135 838 139 839
rect 135 833 139 834
rect 167 838 171 839
rect 167 833 171 834
rect 207 838 211 839
rect 207 833 211 834
rect 231 838 235 839
rect 231 833 235 834
rect 279 838 283 839
rect 279 833 283 834
rect 327 838 331 839
rect 327 833 331 834
rect 399 838 403 839
rect 399 833 403 834
rect 407 838 411 839
rect 407 833 411 834
rect 435 838 439 839
rect 435 833 439 834
rect 559 838 563 839
rect 559 833 563 834
rect 591 838 595 839
rect 591 833 595 834
rect 663 838 667 839
rect 663 833 667 834
rect 679 838 683 839
rect 679 833 683 834
rect 727 838 731 839
rect 727 833 731 834
rect 815 838 819 839
rect 815 833 819 834
rect 863 838 867 839
rect 863 833 867 834
rect 951 838 955 839
rect 951 833 955 834
rect 999 838 1003 839
rect 999 833 1003 834
rect 1031 838 1035 839
rect 1031 833 1035 834
rect 1039 838 1043 839
rect 1039 833 1043 834
rect 1071 838 1075 839
rect 1071 833 1075 834
rect 1103 838 1107 839
rect 1103 833 1107 834
rect 1111 838 1115 839
rect 1111 833 1115 834
rect 1143 838 1147 839
rect 1143 833 1147 834
rect 1167 838 1171 839
rect 1167 833 1171 834
rect 1239 838 1243 839
rect 1239 833 1243 834
rect 1247 838 1251 839
rect 1247 833 1251 834
rect 1271 838 1275 839
rect 1271 833 1275 834
rect 1295 838 1299 839
rect 1295 833 1299 834
rect 1327 838 1331 839
rect 1327 833 1331 834
rect 1375 838 1379 839
rect 1375 833 1379 834
rect 1423 838 1427 839
rect 1423 833 1427 834
rect 1471 838 1475 839
rect 1471 833 1475 834
rect 1519 838 1523 839
rect 1519 833 1523 834
rect 1559 838 1563 839
rect 1559 833 1563 834
rect 1591 838 1595 839
rect 1591 833 1595 834
rect 1623 838 1627 839
rect 1623 833 1627 834
rect 1655 838 1659 839
rect 1655 833 1659 834
rect 1695 838 1699 839
rect 1695 833 1699 834
rect 112 805 114 833
rect 110 804 116 805
rect 110 800 111 804
rect 115 800 116 804
rect 136 803 138 833
rect 232 824 234 833
rect 408 824 410 833
rect 230 823 236 824
rect 230 819 231 823
rect 235 819 236 823
rect 230 818 236 819
rect 406 823 412 824
rect 406 819 407 823
rect 411 819 412 823
rect 406 818 412 819
rect 560 803 562 833
rect 664 818 666 833
rect 816 824 818 833
rect 814 823 820 824
rect 814 819 815 823
rect 819 819 820 823
rect 814 818 820 819
rect 662 817 668 818
rect 662 813 663 817
rect 667 813 668 817
rect 662 812 668 813
rect 952 808 954 833
rect 950 807 956 808
rect 950 803 951 807
rect 955 803 956 807
rect 1032 806 1034 833
rect 110 799 116 800
rect 134 802 140 803
rect 134 798 135 802
rect 139 798 140 802
rect 134 797 140 798
rect 558 802 564 803
rect 950 802 956 803
rect 1030 805 1036 806
rect 558 798 559 802
rect 563 798 564 802
rect 1030 801 1031 805
rect 1035 801 1036 805
rect 1104 803 1106 833
rect 1168 806 1170 833
rect 1248 806 1250 833
rect 1166 805 1172 806
rect 1030 800 1036 801
rect 1102 802 1108 803
rect 558 797 564 798
rect 1102 798 1103 802
rect 1107 798 1108 802
rect 1166 801 1167 805
rect 1171 801 1172 805
rect 1166 800 1172 801
rect 1246 805 1252 806
rect 1246 801 1247 805
rect 1251 801 1252 805
rect 1296 804 1298 833
rect 1328 804 1330 833
rect 1424 813 1426 833
rect 1472 813 1474 833
rect 1422 812 1428 813
rect 1422 808 1423 812
rect 1427 808 1428 812
rect 1422 807 1428 808
rect 1470 812 1476 813
rect 1470 808 1471 812
rect 1475 808 1476 812
rect 1470 807 1476 808
rect 1246 800 1252 801
rect 1294 803 1300 804
rect 1294 799 1295 803
rect 1299 799 1300 803
rect 1294 798 1300 799
rect 1326 803 1332 804
rect 1520 803 1522 833
rect 1560 803 1562 833
rect 1592 803 1594 833
rect 1624 803 1626 833
rect 1656 803 1658 833
rect 1696 805 1698 833
rect 1694 804 1700 805
rect 1326 799 1327 803
rect 1331 799 1332 803
rect 1326 798 1332 799
rect 1518 802 1524 803
rect 1518 798 1519 802
rect 1523 798 1524 802
rect 1102 797 1108 798
rect 1518 797 1524 798
rect 1558 802 1564 803
rect 1558 798 1559 802
rect 1563 798 1564 802
rect 1558 797 1564 798
rect 1590 802 1596 803
rect 1590 798 1591 802
rect 1595 798 1596 802
rect 1590 797 1596 798
rect 1622 802 1628 803
rect 1622 798 1623 802
rect 1627 798 1628 802
rect 1622 797 1628 798
rect 1654 802 1660 803
rect 1654 798 1655 802
rect 1659 798 1660 802
rect 1694 800 1695 804
rect 1699 800 1700 804
rect 1694 799 1700 800
rect 1654 797 1660 798
rect 110 787 116 788
rect 110 783 111 787
rect 115 783 116 787
rect 1694 787 1700 788
rect 110 782 116 783
rect 134 785 140 786
rect 112 755 114 782
rect 134 781 135 785
rect 139 781 140 785
rect 558 785 564 786
rect 1102 785 1108 786
rect 1294 785 1300 786
rect 1518 785 1524 786
rect 134 780 140 781
rect 230 782 236 783
rect 136 755 138 780
rect 230 778 231 782
rect 235 778 236 782
rect 230 777 236 778
rect 406 782 412 783
rect 406 778 407 782
rect 411 778 412 782
rect 558 781 559 785
rect 563 781 564 785
rect 950 784 956 785
rect 558 780 564 781
rect 814 782 820 783
rect 406 777 412 778
rect 232 755 234 777
rect 408 755 410 777
rect 560 755 562 780
rect 814 778 815 782
rect 819 778 820 782
rect 950 780 951 784
rect 955 780 956 784
rect 950 779 956 780
rect 1014 784 1020 785
rect 1014 780 1015 784
rect 1019 780 1020 784
rect 1102 781 1103 785
rect 1107 781 1108 785
rect 1102 780 1108 781
rect 1230 784 1236 785
rect 1230 780 1231 784
rect 1235 780 1236 784
rect 1294 781 1295 785
rect 1299 781 1300 785
rect 1294 780 1300 781
rect 1326 784 1332 785
rect 1326 780 1327 784
rect 1331 780 1332 784
rect 1014 779 1020 780
rect 654 777 660 778
rect 814 777 820 778
rect 654 773 655 777
rect 659 773 660 777
rect 654 772 660 773
rect 656 755 658 772
rect 816 755 818 777
rect 952 755 954 779
rect 1016 755 1018 779
rect 1104 755 1106 780
rect 1230 779 1236 780
rect 1182 778 1188 779
rect 1182 774 1183 778
rect 1187 774 1188 778
rect 1182 773 1188 774
rect 1184 755 1186 773
rect 1232 755 1234 779
rect 1296 755 1298 780
rect 1326 779 1332 780
rect 1422 784 1428 785
rect 1422 780 1423 784
rect 1427 780 1428 784
rect 1422 779 1428 780
rect 1470 784 1476 785
rect 1470 780 1471 784
rect 1475 780 1476 784
rect 1518 781 1519 785
rect 1523 781 1524 785
rect 1518 780 1524 781
rect 1558 785 1564 786
rect 1558 781 1559 785
rect 1563 781 1564 785
rect 1558 780 1564 781
rect 1590 785 1596 786
rect 1590 781 1591 785
rect 1595 781 1596 785
rect 1590 780 1596 781
rect 1622 785 1628 786
rect 1622 781 1623 785
rect 1627 781 1628 785
rect 1622 780 1628 781
rect 1654 785 1660 786
rect 1654 781 1655 785
rect 1659 781 1660 785
rect 1694 783 1695 787
rect 1699 783 1700 787
rect 1694 782 1700 783
rect 1654 780 1660 781
rect 1470 779 1476 780
rect 1328 755 1330 779
rect 1424 755 1426 779
rect 1472 755 1474 779
rect 1520 755 1522 780
rect 1560 755 1562 780
rect 1592 755 1594 780
rect 1624 755 1626 780
rect 1656 755 1658 780
rect 1696 755 1698 782
rect 111 754 115 755
rect 111 749 115 750
rect 135 754 139 755
rect 135 749 139 750
rect 215 754 219 755
rect 215 749 219 750
rect 231 754 235 755
rect 231 749 235 750
rect 287 754 291 755
rect 287 749 291 750
rect 391 754 395 755
rect 391 749 395 750
rect 407 754 411 755
rect 407 749 411 750
rect 471 754 475 755
rect 471 749 475 750
rect 559 754 563 755
rect 559 749 563 750
rect 615 754 619 755
rect 615 749 619 750
rect 655 754 659 755
rect 655 749 659 750
rect 719 754 723 755
rect 719 749 723 750
rect 767 754 771 755
rect 767 749 771 750
rect 815 754 819 755
rect 815 749 819 750
rect 863 754 867 755
rect 863 749 867 750
rect 911 754 915 755
rect 911 749 915 750
rect 951 754 955 755
rect 951 749 955 750
rect 999 754 1003 755
rect 999 749 1003 750
rect 1015 754 1019 755
rect 1015 749 1019 750
rect 1087 754 1091 755
rect 1087 749 1091 750
rect 1103 754 1107 755
rect 1103 749 1107 750
rect 1167 754 1171 755
rect 1167 749 1171 750
rect 1183 754 1187 755
rect 1183 749 1187 750
rect 1207 754 1211 755
rect 1207 749 1211 750
rect 1231 754 1235 755
rect 1231 749 1235 750
rect 1247 754 1251 755
rect 1247 749 1251 750
rect 1279 754 1283 755
rect 1279 749 1283 750
rect 1295 754 1299 755
rect 1295 749 1299 750
rect 1311 754 1315 755
rect 1311 749 1315 750
rect 1327 754 1331 755
rect 1327 749 1331 750
rect 1343 754 1347 755
rect 1343 749 1347 750
rect 1375 754 1379 755
rect 1375 749 1379 750
rect 1407 754 1411 755
rect 1407 749 1411 750
rect 1423 754 1427 755
rect 1423 749 1427 750
rect 1439 754 1443 755
rect 1439 749 1443 750
rect 1471 754 1475 755
rect 1471 749 1475 750
rect 1479 754 1483 755
rect 1479 749 1483 750
rect 1519 754 1523 755
rect 1519 749 1523 750
rect 1559 754 1563 755
rect 1559 749 1563 750
rect 1591 754 1595 755
rect 1591 749 1595 750
rect 1623 754 1627 755
rect 1623 749 1627 750
rect 1655 754 1659 755
rect 1655 749 1659 750
rect 1695 754 1699 755
rect 1695 749 1699 750
rect 112 726 114 749
rect 136 729 138 749
rect 216 733 218 749
rect 214 732 220 733
rect 134 728 140 729
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 134 724 135 728
rect 139 724 140 728
rect 214 728 215 732
rect 219 728 220 732
rect 288 731 290 749
rect 392 733 394 749
rect 390 732 396 733
rect 214 727 220 728
rect 286 730 292 731
rect 286 726 287 730
rect 291 726 292 730
rect 390 728 391 732
rect 395 728 396 732
rect 390 727 396 728
rect 286 725 292 726
rect 472 725 474 749
rect 616 731 618 749
rect 614 730 620 731
rect 614 726 615 730
rect 619 726 620 730
rect 720 729 722 749
rect 768 736 770 749
rect 766 735 772 736
rect 766 731 767 735
rect 771 731 772 735
rect 766 730 772 731
rect 614 725 620 726
rect 718 728 724 729
rect 864 728 866 749
rect 912 731 914 749
rect 1000 736 1002 749
rect 998 735 1004 736
rect 998 731 999 735
rect 1003 731 1004 735
rect 910 730 916 731
rect 998 730 1004 731
rect 134 723 140 724
rect 470 724 476 725
rect 110 720 116 721
rect 470 720 471 724
rect 475 720 476 724
rect 718 724 719 728
rect 723 724 724 728
rect 718 723 724 724
rect 862 727 868 728
rect 862 723 863 727
rect 867 723 868 727
rect 910 726 911 730
rect 915 726 916 730
rect 1088 729 1090 749
rect 1168 733 1170 749
rect 1166 732 1172 733
rect 910 725 916 726
rect 1086 728 1092 729
rect 1086 724 1087 728
rect 1091 724 1092 728
rect 1166 728 1167 732
rect 1171 728 1172 732
rect 1208 729 1210 749
rect 1166 727 1172 728
rect 1206 728 1212 729
rect 1248 728 1250 749
rect 1280 728 1282 749
rect 1312 728 1314 749
rect 1344 728 1346 749
rect 1376 728 1378 749
rect 1408 728 1410 749
rect 1440 728 1442 749
rect 1480 728 1482 749
rect 1520 728 1522 749
rect 1560 728 1562 749
rect 1592 728 1594 749
rect 1624 728 1626 749
rect 1656 728 1658 749
rect 1086 723 1092 724
rect 1206 724 1207 728
rect 1211 724 1212 728
rect 1206 723 1212 724
rect 1246 727 1252 728
rect 1246 723 1247 727
rect 1251 723 1252 727
rect 862 722 868 723
rect 1246 722 1252 723
rect 1278 727 1284 728
rect 1278 723 1279 727
rect 1283 723 1284 727
rect 1278 722 1284 723
rect 1310 727 1316 728
rect 1310 723 1311 727
rect 1315 723 1316 727
rect 1310 722 1316 723
rect 1342 727 1348 728
rect 1342 723 1343 727
rect 1347 723 1348 727
rect 1342 722 1348 723
rect 1374 727 1380 728
rect 1374 723 1375 727
rect 1379 723 1380 727
rect 1374 722 1380 723
rect 1406 727 1412 728
rect 1406 723 1407 727
rect 1411 723 1412 727
rect 1406 722 1412 723
rect 1438 727 1444 728
rect 1438 723 1439 727
rect 1443 723 1444 727
rect 1438 722 1444 723
rect 1478 727 1484 728
rect 1478 723 1479 727
rect 1483 723 1484 727
rect 1478 722 1484 723
rect 1518 727 1524 728
rect 1518 723 1519 727
rect 1523 723 1524 727
rect 1518 722 1524 723
rect 1558 727 1564 728
rect 1558 723 1559 727
rect 1563 723 1564 727
rect 1558 722 1564 723
rect 1590 727 1596 728
rect 1590 723 1591 727
rect 1595 723 1596 727
rect 1590 722 1596 723
rect 1622 727 1628 728
rect 1622 723 1623 727
rect 1627 723 1628 727
rect 1622 722 1628 723
rect 1654 727 1660 728
rect 1654 723 1655 727
rect 1659 723 1660 727
rect 1696 726 1698 749
rect 1654 722 1660 723
rect 1694 725 1700 726
rect 1694 721 1695 725
rect 1699 721 1700 725
rect 1694 720 1700 721
rect 470 719 476 720
rect 862 710 868 711
rect 442 709 448 710
rect 110 708 116 709
rect 110 704 111 708
rect 115 704 116 708
rect 442 705 443 709
rect 447 705 448 709
rect 862 706 863 710
rect 867 706 868 710
rect 442 704 448 705
rect 718 705 724 706
rect 862 705 868 706
rect 1246 710 1252 711
rect 1246 706 1247 710
rect 1251 706 1252 710
rect 1246 705 1252 706
rect 1278 710 1284 711
rect 1278 706 1279 710
rect 1283 706 1284 710
rect 1278 705 1284 706
rect 1310 710 1316 711
rect 1310 706 1311 710
rect 1315 706 1316 710
rect 1310 705 1316 706
rect 1342 710 1348 711
rect 1342 706 1343 710
rect 1347 706 1348 710
rect 1342 705 1348 706
rect 1374 710 1380 711
rect 1374 706 1375 710
rect 1379 706 1380 710
rect 1374 705 1380 706
rect 1406 710 1412 711
rect 1406 706 1407 710
rect 1411 706 1412 710
rect 1406 705 1412 706
rect 1438 710 1444 711
rect 1438 706 1439 710
rect 1443 706 1444 710
rect 1438 705 1444 706
rect 1478 710 1484 711
rect 1478 706 1479 710
rect 1483 706 1484 710
rect 1478 705 1484 706
rect 1518 710 1524 711
rect 1518 706 1519 710
rect 1523 706 1524 710
rect 1518 705 1524 706
rect 1558 710 1564 711
rect 1558 706 1559 710
rect 1563 706 1564 710
rect 1558 705 1564 706
rect 1590 710 1596 711
rect 1590 706 1591 710
rect 1595 706 1596 710
rect 1590 705 1596 706
rect 1622 710 1628 711
rect 1622 706 1623 710
rect 1627 706 1628 710
rect 1622 705 1628 706
rect 1654 710 1660 711
rect 1654 706 1655 710
rect 1659 706 1660 710
rect 1654 705 1660 706
rect 1694 708 1700 709
rect 110 703 116 704
rect 112 643 114 703
rect 142 690 148 691
rect 142 686 143 690
rect 147 686 148 690
rect 286 689 292 690
rect 142 685 148 686
rect 214 685 220 686
rect 144 643 146 685
rect 214 681 215 685
rect 219 681 220 685
rect 286 685 287 689
rect 291 685 292 689
rect 286 684 292 685
rect 390 685 396 686
rect 214 680 220 681
rect 216 643 218 680
rect 288 643 290 684
rect 390 681 391 685
rect 395 681 396 685
rect 390 680 396 681
rect 392 643 394 680
rect 444 643 446 704
rect 718 701 719 705
rect 723 701 724 705
rect 718 700 724 701
rect 614 689 620 690
rect 614 685 615 689
rect 619 685 620 689
rect 614 684 620 685
rect 616 643 618 684
rect 720 643 722 700
rect 774 695 780 696
rect 774 691 775 695
rect 779 691 780 695
rect 774 690 780 691
rect 776 643 778 690
rect 864 643 866 705
rect 1206 700 1212 701
rect 1206 696 1207 700
rect 1211 696 1212 700
rect 1006 695 1012 696
rect 1206 695 1212 696
rect 1006 691 1007 695
rect 1011 691 1012 695
rect 1006 690 1012 691
rect 1094 690 1100 691
rect 910 689 916 690
rect 910 685 911 689
rect 915 685 916 689
rect 910 684 916 685
rect 912 643 914 684
rect 1008 643 1010 690
rect 1094 686 1095 690
rect 1099 686 1100 690
rect 1094 685 1100 686
rect 1166 685 1172 686
rect 1096 643 1098 685
rect 1166 681 1167 685
rect 1171 681 1172 685
rect 1166 680 1172 681
rect 1168 643 1170 680
rect 1208 643 1210 695
rect 1248 643 1250 705
rect 1280 643 1282 705
rect 1312 643 1314 705
rect 1344 643 1346 705
rect 1376 643 1378 705
rect 1408 643 1410 705
rect 1440 643 1442 705
rect 1480 643 1482 705
rect 1520 643 1522 705
rect 1560 643 1562 705
rect 1592 643 1594 705
rect 1624 643 1626 705
rect 1656 643 1658 705
rect 1694 704 1695 708
rect 1699 704 1700 708
rect 1694 703 1700 704
rect 1696 643 1698 703
rect 111 642 115 643
rect 111 637 115 638
rect 135 642 139 643
rect 135 637 139 638
rect 143 642 147 643
rect 143 637 147 638
rect 167 642 171 643
rect 167 637 171 638
rect 207 642 211 643
rect 207 637 211 638
rect 215 642 219 643
rect 215 637 219 638
rect 287 642 291 643
rect 287 637 291 638
rect 391 642 395 643
rect 391 637 395 638
rect 407 642 411 643
rect 407 637 411 638
rect 443 642 447 643
rect 443 637 447 638
rect 535 642 539 643
rect 535 637 539 638
rect 615 642 619 643
rect 615 637 619 638
rect 671 642 675 643
rect 671 637 675 638
rect 719 642 723 643
rect 719 637 723 638
rect 767 642 771 643
rect 767 637 771 638
rect 775 642 779 643
rect 775 637 779 638
rect 863 642 867 643
rect 863 637 867 638
rect 903 642 907 643
rect 903 637 907 638
rect 911 642 915 643
rect 911 637 915 638
rect 999 642 1003 643
rect 999 637 1003 638
rect 1007 642 1011 643
rect 1007 637 1011 638
rect 1095 642 1099 643
rect 1095 637 1099 638
rect 1119 642 1123 643
rect 1119 637 1123 638
rect 1167 642 1171 643
rect 1167 637 1171 638
rect 1207 642 1211 643
rect 1207 637 1211 638
rect 1215 642 1219 643
rect 1215 637 1219 638
rect 1247 642 1251 643
rect 1247 637 1251 638
rect 1279 642 1283 643
rect 1279 637 1283 638
rect 1311 642 1315 643
rect 1311 637 1315 638
rect 1335 642 1339 643
rect 1335 637 1339 638
rect 1343 642 1347 643
rect 1343 637 1347 638
rect 1375 642 1379 643
rect 1375 637 1379 638
rect 1407 642 1411 643
rect 1407 637 1411 638
rect 1415 642 1419 643
rect 1415 637 1419 638
rect 1439 642 1443 643
rect 1439 637 1443 638
rect 1479 642 1483 643
rect 1479 637 1483 638
rect 1519 642 1523 643
rect 1519 637 1523 638
rect 1543 642 1547 643
rect 1543 637 1547 638
rect 1559 642 1563 643
rect 1559 637 1563 638
rect 1591 642 1595 643
rect 1591 637 1595 638
rect 1607 642 1611 643
rect 1607 637 1611 638
rect 1623 642 1627 643
rect 1623 637 1627 638
rect 1655 642 1659 643
rect 1655 637 1659 638
rect 1695 642 1699 643
rect 1695 637 1699 638
rect 112 605 114 637
rect 110 604 116 605
rect 110 600 111 604
rect 115 600 116 604
rect 136 603 138 637
rect 168 603 170 637
rect 208 628 210 637
rect 206 627 212 628
rect 206 623 207 627
rect 211 623 212 627
rect 288 623 290 637
rect 408 623 410 637
rect 536 624 538 637
rect 534 623 540 624
rect 206 622 212 623
rect 286 622 292 623
rect 286 618 287 622
rect 291 618 292 622
rect 286 617 292 618
rect 406 622 412 623
rect 406 618 407 622
rect 411 618 412 622
rect 534 619 535 623
rect 539 619 540 623
rect 534 618 540 619
rect 406 617 412 618
rect 672 603 674 637
rect 768 624 770 637
rect 904 628 906 637
rect 902 627 908 628
rect 766 623 772 624
rect 766 619 767 623
rect 771 619 772 623
rect 902 623 903 627
rect 907 623 908 627
rect 1000 623 1002 637
rect 1120 628 1122 637
rect 1118 627 1124 628
rect 1118 623 1119 627
rect 1123 623 1124 627
rect 1216 623 1218 637
rect 1336 628 1338 637
rect 1334 627 1340 628
rect 1334 623 1335 627
rect 1339 623 1340 627
rect 902 622 908 623
rect 998 622 1004 623
rect 1118 622 1124 623
rect 1214 622 1220 623
rect 1334 622 1340 623
rect 766 618 772 619
rect 998 618 999 622
rect 1003 618 1004 622
rect 998 617 1004 618
rect 1214 618 1215 622
rect 1219 618 1220 622
rect 1214 617 1220 618
rect 1416 603 1418 637
rect 1480 603 1482 637
rect 1544 603 1546 637
rect 1608 603 1610 637
rect 1656 603 1658 637
rect 1696 605 1698 637
rect 1694 604 1700 605
rect 110 599 116 600
rect 134 602 140 603
rect 134 598 135 602
rect 139 598 140 602
rect 134 597 140 598
rect 166 602 172 603
rect 166 598 167 602
rect 171 598 172 602
rect 166 597 172 598
rect 670 602 676 603
rect 670 598 671 602
rect 675 598 676 602
rect 670 597 676 598
rect 1414 602 1420 603
rect 1414 598 1415 602
rect 1419 598 1420 602
rect 1414 597 1420 598
rect 1478 602 1484 603
rect 1478 598 1479 602
rect 1483 598 1484 602
rect 1478 597 1484 598
rect 1542 602 1548 603
rect 1542 598 1543 602
rect 1547 598 1548 602
rect 1542 597 1548 598
rect 1606 602 1612 603
rect 1606 598 1607 602
rect 1611 598 1612 602
rect 1606 597 1612 598
rect 1654 602 1660 603
rect 1654 598 1655 602
rect 1659 598 1660 602
rect 1694 600 1695 604
rect 1699 600 1700 604
rect 1694 599 1700 600
rect 1654 597 1660 598
rect 110 587 116 588
rect 110 583 111 587
rect 115 583 116 587
rect 1694 587 1700 588
rect 110 582 116 583
rect 134 585 140 586
rect 112 563 114 582
rect 134 581 135 585
rect 139 581 140 585
rect 134 580 140 581
rect 166 585 172 586
rect 670 585 676 586
rect 1414 585 1420 586
rect 166 581 167 585
rect 171 581 172 585
rect 278 584 284 585
rect 166 580 172 581
rect 206 580 212 581
rect 136 563 138 580
rect 168 563 170 580
rect 206 576 207 580
rect 211 576 212 580
rect 278 580 279 584
rect 283 580 284 584
rect 278 579 284 580
rect 398 584 404 585
rect 398 580 399 584
rect 403 580 404 584
rect 398 579 404 580
rect 534 582 540 583
rect 206 575 212 576
rect 208 563 210 575
rect 280 563 282 579
rect 400 563 402 579
rect 534 578 535 582
rect 539 578 540 582
rect 670 581 671 585
rect 675 581 676 585
rect 990 584 996 585
rect 670 580 676 581
rect 766 582 772 583
rect 534 577 540 578
rect 536 563 538 577
rect 672 563 674 580
rect 766 578 767 582
rect 771 578 772 582
rect 766 577 772 578
rect 902 580 908 581
rect 768 563 770 577
rect 902 576 903 580
rect 907 576 908 580
rect 990 580 991 584
rect 995 580 996 584
rect 1206 584 1212 585
rect 990 579 996 580
rect 1118 580 1124 581
rect 902 575 908 576
rect 904 563 906 575
rect 992 563 994 579
rect 1118 576 1119 580
rect 1123 576 1124 580
rect 1206 580 1207 584
rect 1211 580 1212 584
rect 1414 581 1415 585
rect 1419 581 1420 585
rect 1206 579 1212 580
rect 1334 580 1340 581
rect 1414 580 1420 581
rect 1478 585 1484 586
rect 1478 581 1479 585
rect 1483 581 1484 585
rect 1478 580 1484 581
rect 1542 585 1548 586
rect 1542 581 1543 585
rect 1547 581 1548 585
rect 1542 580 1548 581
rect 1606 585 1612 586
rect 1606 581 1607 585
rect 1611 581 1612 585
rect 1606 580 1612 581
rect 1654 585 1660 586
rect 1654 581 1655 585
rect 1659 581 1660 585
rect 1694 583 1695 587
rect 1699 583 1700 587
rect 1694 582 1700 583
rect 1654 580 1660 581
rect 1118 575 1124 576
rect 1120 563 1122 575
rect 1208 563 1210 579
rect 1334 576 1335 580
rect 1339 576 1340 580
rect 1334 575 1340 576
rect 1336 563 1338 575
rect 1416 563 1418 580
rect 1480 563 1482 580
rect 1544 563 1546 580
rect 1608 563 1610 580
rect 1656 563 1658 580
rect 1696 563 1698 582
rect 111 562 115 563
rect 111 557 115 558
rect 135 562 139 563
rect 135 557 139 558
rect 167 562 171 563
rect 167 557 171 558
rect 207 562 211 563
rect 207 557 211 558
rect 247 562 251 563
rect 247 557 251 558
rect 279 562 283 563
rect 279 557 283 558
rect 303 562 307 563
rect 303 557 307 558
rect 391 562 395 563
rect 391 557 395 558
rect 399 562 403 563
rect 399 557 403 558
rect 471 562 475 563
rect 471 557 475 558
rect 535 562 539 563
rect 535 557 539 558
rect 647 562 651 563
rect 647 557 651 558
rect 671 562 675 563
rect 671 557 675 558
rect 727 562 731 563
rect 727 557 731 558
rect 767 562 771 563
rect 767 557 771 558
rect 775 562 779 563
rect 775 557 779 558
rect 871 562 875 563
rect 871 557 875 558
rect 903 562 907 563
rect 903 557 907 558
rect 927 562 931 563
rect 927 557 931 558
rect 991 562 995 563
rect 991 557 995 558
rect 1031 562 1035 563
rect 1031 557 1035 558
rect 1095 562 1099 563
rect 1095 557 1099 558
rect 1119 562 1123 563
rect 1119 557 1123 558
rect 1199 562 1203 563
rect 1199 557 1203 558
rect 1207 562 1211 563
rect 1207 557 1211 558
rect 1287 562 1291 563
rect 1287 557 1291 558
rect 1335 562 1339 563
rect 1335 557 1339 558
rect 1415 562 1419 563
rect 1415 557 1419 558
rect 1423 562 1427 563
rect 1423 557 1427 558
rect 1479 562 1483 563
rect 1479 557 1483 558
rect 1527 562 1531 563
rect 1527 557 1531 558
rect 1543 562 1547 563
rect 1543 557 1547 558
rect 1575 562 1579 563
rect 1575 557 1579 558
rect 1607 562 1611 563
rect 1607 557 1611 558
rect 1623 562 1627 563
rect 1623 557 1627 558
rect 1655 562 1659 563
rect 1655 557 1659 558
rect 1695 562 1699 563
rect 1695 557 1699 558
rect 112 534 114 557
rect 136 536 138 557
rect 168 537 170 557
rect 248 541 250 557
rect 246 540 252 541
rect 166 536 172 537
rect 134 535 140 536
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 134 531 135 535
rect 139 531 140 535
rect 166 532 167 536
rect 171 532 172 536
rect 246 536 247 540
rect 251 536 252 540
rect 304 539 306 557
rect 246 535 252 536
rect 302 538 308 539
rect 302 534 303 538
rect 307 534 308 538
rect 392 537 394 557
rect 472 541 474 557
rect 470 540 476 541
rect 302 533 308 534
rect 390 536 396 537
rect 166 531 172 532
rect 390 532 391 536
rect 395 532 396 536
rect 470 536 471 540
rect 475 536 476 540
rect 470 535 476 536
rect 536 533 538 557
rect 648 537 650 557
rect 728 541 730 557
rect 726 540 732 541
rect 646 536 652 537
rect 390 531 396 532
rect 534 532 540 533
rect 134 530 140 531
rect 110 528 116 529
rect 534 528 535 532
rect 539 528 540 532
rect 646 532 647 536
rect 651 532 652 536
rect 726 536 727 540
rect 731 536 732 540
rect 776 537 778 557
rect 872 541 874 557
rect 870 540 876 541
rect 726 535 732 536
rect 774 536 780 537
rect 646 531 652 532
rect 774 532 775 536
rect 779 532 780 536
rect 870 536 871 540
rect 875 536 876 540
rect 928 537 930 557
rect 1032 541 1034 557
rect 1030 540 1036 541
rect 870 535 876 536
rect 926 536 932 537
rect 774 531 780 532
rect 926 532 927 536
rect 931 532 932 536
rect 1030 536 1031 540
rect 1035 536 1036 540
rect 1096 537 1098 557
rect 1200 541 1202 557
rect 1198 540 1204 541
rect 1030 535 1036 536
rect 1094 536 1100 537
rect 926 531 932 532
rect 1094 532 1095 536
rect 1099 532 1100 536
rect 1198 536 1199 540
rect 1203 536 1204 540
rect 1198 535 1204 536
rect 1288 533 1290 557
rect 1424 536 1426 557
rect 1480 536 1482 557
rect 1528 536 1530 557
rect 1576 536 1578 557
rect 1624 536 1626 557
rect 1656 536 1658 557
rect 1422 535 1428 536
rect 1094 531 1100 532
rect 1286 532 1292 533
rect 534 527 540 528
rect 1286 528 1287 532
rect 1291 528 1292 532
rect 1422 531 1423 535
rect 1427 531 1428 535
rect 1422 530 1428 531
rect 1478 535 1484 536
rect 1478 531 1479 535
rect 1483 531 1484 535
rect 1478 530 1484 531
rect 1526 535 1532 536
rect 1526 531 1527 535
rect 1531 531 1532 535
rect 1526 530 1532 531
rect 1574 535 1580 536
rect 1574 531 1575 535
rect 1579 531 1580 535
rect 1574 530 1580 531
rect 1622 535 1628 536
rect 1622 531 1623 535
rect 1627 531 1628 535
rect 1622 530 1628 531
rect 1654 535 1660 536
rect 1654 531 1655 535
rect 1659 531 1660 535
rect 1696 534 1698 557
rect 1654 530 1660 531
rect 1694 533 1700 534
rect 1694 529 1695 533
rect 1699 529 1700 533
rect 1694 528 1700 529
rect 1286 527 1292 528
rect 134 518 140 519
rect 1422 518 1428 519
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 134 514 135 518
rect 139 514 140 518
rect 134 513 140 514
rect 506 517 512 518
rect 506 513 507 517
rect 511 513 512 517
rect 110 511 116 512
rect 112 443 114 511
rect 136 443 138 513
rect 506 512 512 513
rect 1258 517 1264 518
rect 1258 513 1259 517
rect 1263 513 1264 517
rect 1422 514 1423 518
rect 1427 514 1428 518
rect 1422 513 1428 514
rect 1478 518 1484 519
rect 1478 514 1479 518
rect 1483 514 1484 518
rect 1478 513 1484 514
rect 1526 518 1532 519
rect 1526 514 1527 518
rect 1531 514 1532 518
rect 1526 513 1532 514
rect 1574 518 1580 519
rect 1574 514 1575 518
rect 1579 514 1580 518
rect 1574 513 1580 514
rect 1622 518 1628 519
rect 1622 514 1623 518
rect 1627 514 1628 518
rect 1622 513 1628 514
rect 1654 518 1660 519
rect 1654 514 1655 518
rect 1659 514 1660 518
rect 1654 513 1660 514
rect 1694 516 1700 517
rect 1258 512 1264 513
rect 174 498 180 499
rect 398 498 404 499
rect 174 494 175 498
rect 179 494 180 498
rect 302 497 308 498
rect 174 493 180 494
rect 246 493 252 494
rect 176 443 178 493
rect 246 489 247 493
rect 251 489 252 493
rect 302 493 303 497
rect 307 493 308 497
rect 398 494 399 498
rect 403 494 404 498
rect 398 493 404 494
rect 470 493 476 494
rect 302 492 308 493
rect 246 488 252 489
rect 248 443 250 488
rect 304 443 306 492
rect 400 443 402 493
rect 470 489 471 493
rect 475 489 476 493
rect 470 488 476 489
rect 472 443 474 488
rect 508 443 510 512
rect 654 498 660 499
rect 654 494 655 498
rect 659 494 660 498
rect 782 498 788 499
rect 782 494 783 498
rect 787 494 788 498
rect 934 498 940 499
rect 934 494 935 498
rect 939 494 940 498
rect 1102 498 1108 499
rect 1102 494 1103 498
rect 1107 494 1108 498
rect 654 493 660 494
rect 726 493 732 494
rect 782 493 788 494
rect 870 493 876 494
rect 934 493 940 494
rect 1030 493 1036 494
rect 1102 493 1108 494
rect 1198 493 1204 494
rect 656 443 658 493
rect 726 489 727 493
rect 731 489 732 493
rect 726 488 732 489
rect 728 443 730 488
rect 784 443 786 493
rect 870 489 871 493
rect 875 489 876 493
rect 870 488 876 489
rect 872 443 874 488
rect 936 443 938 493
rect 1030 489 1031 493
rect 1035 489 1036 493
rect 1030 488 1036 489
rect 1032 443 1034 488
rect 1104 443 1106 493
rect 1198 489 1199 493
rect 1203 489 1204 493
rect 1198 488 1204 489
rect 1200 443 1202 488
rect 1260 443 1262 512
rect 1424 443 1426 513
rect 1480 443 1482 513
rect 1528 443 1530 513
rect 1576 443 1578 513
rect 1624 443 1626 513
rect 1656 443 1658 513
rect 1694 512 1695 516
rect 1699 512 1700 516
rect 1694 511 1700 512
rect 1696 443 1698 511
rect 111 442 115 443
rect 111 437 115 438
rect 135 442 139 443
rect 135 437 139 438
rect 167 442 171 443
rect 167 437 171 438
rect 175 442 179 443
rect 175 437 179 438
rect 199 442 203 443
rect 199 437 203 438
rect 231 442 235 443
rect 231 437 235 438
rect 247 442 251 443
rect 247 437 251 438
rect 263 442 267 443
rect 263 437 267 438
rect 303 442 307 443
rect 303 437 307 438
rect 375 442 379 443
rect 375 437 379 438
rect 399 442 403 443
rect 399 437 403 438
rect 415 442 419 443
rect 415 437 419 438
rect 447 442 451 443
rect 447 437 451 438
rect 471 442 475 443
rect 471 437 475 438
rect 487 442 491 443
rect 487 437 491 438
rect 507 442 511 443
rect 507 437 511 438
rect 543 442 547 443
rect 543 437 547 438
rect 615 442 619 443
rect 615 437 619 438
rect 655 442 659 443
rect 655 437 659 438
rect 671 442 675 443
rect 671 437 675 438
rect 727 442 731 443
rect 727 437 731 438
rect 755 442 759 443
rect 755 437 759 438
rect 783 442 787 443
rect 783 437 787 438
rect 871 442 875 443
rect 871 437 875 438
rect 903 442 907 443
rect 903 437 907 438
rect 935 442 939 443
rect 935 437 939 438
rect 951 442 955 443
rect 951 437 955 438
rect 1031 442 1035 443
rect 1031 437 1035 438
rect 1075 442 1079 443
rect 1075 437 1079 438
rect 1103 442 1107 443
rect 1103 437 1107 438
rect 1199 442 1203 443
rect 1199 437 1203 438
rect 1231 442 1235 443
rect 1231 437 1235 438
rect 1259 442 1263 443
rect 1259 437 1263 438
rect 1319 442 1323 443
rect 1319 437 1323 438
rect 1359 442 1363 443
rect 1359 437 1363 438
rect 1423 442 1427 443
rect 1423 437 1427 438
rect 1439 442 1443 443
rect 1439 437 1443 438
rect 1479 442 1483 443
rect 1479 437 1483 438
rect 1519 442 1523 443
rect 1519 437 1523 438
rect 1527 442 1531 443
rect 1527 437 1531 438
rect 1559 442 1563 443
rect 1559 437 1563 438
rect 1575 442 1579 443
rect 1575 437 1579 438
rect 1591 442 1595 443
rect 1591 437 1595 438
rect 1623 442 1627 443
rect 1623 437 1627 438
rect 1655 442 1659 443
rect 1655 437 1659 438
rect 1695 442 1699 443
rect 1695 437 1699 438
rect 112 377 114 437
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 136 375 138 437
rect 168 375 170 437
rect 200 375 202 437
rect 232 375 234 437
rect 264 375 266 437
rect 304 395 306 437
rect 376 400 378 437
rect 374 399 380 400
rect 374 395 375 399
rect 379 395 380 399
rect 302 394 308 395
rect 374 394 380 395
rect 302 390 303 394
rect 307 390 308 394
rect 302 389 308 390
rect 416 375 418 437
rect 448 375 450 437
rect 488 378 490 437
rect 544 395 546 437
rect 616 400 618 437
rect 614 399 620 400
rect 614 395 615 399
rect 619 395 620 399
rect 672 396 674 437
rect 542 394 548 395
rect 614 394 620 395
rect 670 395 676 396
rect 542 390 543 394
rect 547 390 548 394
rect 670 391 671 395
rect 675 391 676 395
rect 670 390 676 391
rect 542 389 548 390
rect 486 377 492 378
rect 110 371 116 372
rect 134 374 140 375
rect 134 370 135 374
rect 139 370 140 374
rect 134 369 140 370
rect 166 374 172 375
rect 166 370 167 374
rect 171 370 172 374
rect 166 369 172 370
rect 198 374 204 375
rect 198 370 199 374
rect 203 370 204 374
rect 198 369 204 370
rect 230 374 236 375
rect 230 370 231 374
rect 235 370 236 374
rect 230 369 236 370
rect 262 374 268 375
rect 262 370 263 374
rect 267 370 268 374
rect 262 369 268 370
rect 414 374 420 375
rect 414 370 415 374
rect 419 370 420 374
rect 414 369 420 370
rect 446 374 452 375
rect 446 370 447 374
rect 451 370 452 374
rect 486 373 487 377
rect 491 373 492 377
rect 756 376 758 437
rect 486 372 492 373
rect 754 375 760 376
rect 904 375 906 437
rect 952 395 954 437
rect 950 394 956 395
rect 950 390 951 394
rect 955 390 956 394
rect 950 389 956 390
rect 1032 378 1034 437
rect 1030 377 1036 378
rect 754 371 755 375
rect 759 371 760 375
rect 754 370 760 371
rect 902 374 908 375
rect 902 370 903 374
rect 907 370 908 374
rect 1030 373 1031 377
rect 1035 373 1036 377
rect 1076 376 1078 437
rect 1232 396 1234 437
rect 1230 395 1236 396
rect 1230 391 1231 395
rect 1235 391 1236 395
rect 1230 390 1236 391
rect 1030 372 1036 373
rect 1074 375 1080 376
rect 1320 375 1322 437
rect 1360 390 1362 437
rect 1358 389 1364 390
rect 1358 385 1359 389
rect 1363 385 1364 389
rect 1358 384 1364 385
rect 1440 380 1442 437
rect 1438 379 1444 380
rect 1438 375 1439 379
rect 1443 375 1444 379
rect 1480 375 1482 437
rect 1520 375 1522 437
rect 1560 375 1562 437
rect 1592 375 1594 437
rect 1624 375 1626 437
rect 1656 375 1658 437
rect 1696 377 1698 437
rect 1694 376 1700 377
rect 1074 371 1075 375
rect 1079 371 1080 375
rect 1074 370 1080 371
rect 1318 374 1324 375
rect 1438 374 1444 375
rect 1478 374 1484 375
rect 1318 370 1319 374
rect 1323 370 1324 374
rect 446 369 452 370
rect 902 369 908 370
rect 1318 369 1324 370
rect 1478 370 1479 374
rect 1483 370 1484 374
rect 1478 369 1484 370
rect 1518 374 1524 375
rect 1518 370 1519 374
rect 1523 370 1524 374
rect 1518 369 1524 370
rect 1558 374 1564 375
rect 1558 370 1559 374
rect 1563 370 1564 374
rect 1558 369 1564 370
rect 1590 374 1596 375
rect 1590 370 1591 374
rect 1595 370 1596 374
rect 1590 369 1596 370
rect 1622 374 1628 375
rect 1622 370 1623 374
rect 1627 370 1628 374
rect 1622 369 1628 370
rect 1654 374 1660 375
rect 1654 370 1655 374
rect 1659 370 1660 374
rect 1694 372 1695 376
rect 1699 372 1700 376
rect 1694 371 1700 372
rect 1654 369 1660 370
rect 782 360 788 361
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 134 357 140 358
rect 112 323 114 354
rect 134 353 135 357
rect 139 353 140 357
rect 134 352 140 353
rect 166 357 172 358
rect 166 353 167 357
rect 171 353 172 357
rect 166 352 172 353
rect 198 357 204 358
rect 198 353 199 357
rect 203 353 204 357
rect 198 352 204 353
rect 230 357 236 358
rect 230 353 231 357
rect 235 353 236 357
rect 230 352 236 353
rect 262 357 268 358
rect 414 357 420 358
rect 262 353 263 357
rect 267 353 268 357
rect 262 352 268 353
rect 294 356 300 357
rect 294 352 295 356
rect 299 352 300 356
rect 414 353 415 357
rect 419 353 420 357
rect 136 323 138 352
rect 168 323 170 352
rect 200 323 202 352
rect 232 323 234 352
rect 264 323 266 352
rect 294 351 300 352
rect 374 352 380 353
rect 414 352 420 353
rect 446 357 452 358
rect 446 353 447 357
rect 451 353 452 357
rect 446 352 452 353
rect 534 356 540 357
rect 534 352 535 356
rect 539 352 540 356
rect 782 356 783 360
rect 787 356 788 360
rect 1102 360 1108 361
rect 782 355 788 356
rect 902 357 908 358
rect 670 354 676 355
rect 296 323 298 351
rect 374 348 375 352
rect 379 348 380 352
rect 374 347 380 348
rect 376 323 378 347
rect 416 323 418 352
rect 448 323 450 352
rect 534 351 540 352
rect 614 352 620 353
rect 502 350 508 351
rect 502 346 503 350
rect 507 346 508 350
rect 502 345 508 346
rect 504 323 506 345
rect 536 323 538 351
rect 614 348 615 352
rect 619 348 620 352
rect 670 350 671 354
rect 675 350 676 354
rect 670 349 676 350
rect 614 347 620 348
rect 616 323 618 347
rect 672 323 674 349
rect 784 323 786 355
rect 902 353 903 357
rect 907 353 908 357
rect 902 352 908 353
rect 942 356 948 357
rect 942 352 943 356
rect 947 352 948 356
rect 1102 356 1103 360
rect 1107 356 1108 360
rect 1694 359 1700 360
rect 1102 355 1108 356
rect 1318 357 1324 358
rect 1478 357 1484 358
rect 904 323 906 352
rect 942 351 948 352
rect 944 323 946 351
rect 1046 350 1052 351
rect 1046 346 1047 350
rect 1051 346 1052 350
rect 1046 345 1052 346
rect 1048 323 1050 345
rect 1104 323 1106 355
rect 1230 354 1236 355
rect 1230 350 1231 354
rect 1235 350 1236 354
rect 1318 353 1319 357
rect 1323 353 1324 357
rect 1318 352 1324 353
rect 1438 356 1444 357
rect 1438 352 1439 356
rect 1443 352 1444 356
rect 1478 353 1479 357
rect 1483 353 1484 357
rect 1478 352 1484 353
rect 1518 357 1524 358
rect 1518 353 1519 357
rect 1523 353 1524 357
rect 1518 352 1524 353
rect 1558 357 1564 358
rect 1558 353 1559 357
rect 1563 353 1564 357
rect 1558 352 1564 353
rect 1590 357 1596 358
rect 1590 353 1591 357
rect 1595 353 1596 357
rect 1590 352 1596 353
rect 1622 357 1628 358
rect 1622 353 1623 357
rect 1627 353 1628 357
rect 1622 352 1628 353
rect 1654 357 1660 358
rect 1654 353 1655 357
rect 1659 353 1660 357
rect 1694 355 1695 359
rect 1699 355 1700 359
rect 1694 354 1700 355
rect 1654 352 1660 353
rect 1230 349 1236 350
rect 1232 323 1234 349
rect 1320 323 1322 352
rect 1438 351 1444 352
rect 1350 349 1356 350
rect 1350 345 1351 349
rect 1355 345 1356 349
rect 1350 344 1356 345
rect 1352 323 1354 344
rect 1440 323 1442 351
rect 1480 323 1482 352
rect 1520 323 1522 352
rect 1560 323 1562 352
rect 1592 323 1594 352
rect 1624 323 1626 352
rect 1656 323 1658 352
rect 1696 323 1698 354
rect 111 322 115 323
rect 111 317 115 318
rect 135 322 139 323
rect 135 317 139 318
rect 167 322 171 323
rect 167 317 171 318
rect 199 322 203 323
rect 199 317 203 318
rect 231 322 235 323
rect 231 317 235 318
rect 263 322 267 323
rect 263 317 267 318
rect 295 322 299 323
rect 295 317 299 318
rect 327 322 331 323
rect 327 317 331 318
rect 359 322 363 323
rect 359 317 363 318
rect 375 322 379 323
rect 375 317 379 318
rect 391 322 395 323
rect 391 317 395 318
rect 415 322 419 323
rect 415 317 419 318
rect 423 322 427 323
rect 423 317 427 318
rect 447 322 451 323
rect 447 317 451 318
rect 455 322 459 323
rect 455 317 459 318
rect 487 322 491 323
rect 487 317 491 318
rect 503 322 507 323
rect 503 317 507 318
rect 519 322 523 323
rect 519 317 523 318
rect 535 322 539 323
rect 535 317 539 318
rect 551 322 555 323
rect 551 317 555 318
rect 599 322 603 323
rect 599 317 603 318
rect 615 322 619 323
rect 615 317 619 318
rect 671 322 675 323
rect 671 317 675 318
rect 703 322 707 323
rect 703 317 707 318
rect 783 322 787 323
rect 783 317 787 318
rect 807 322 811 323
rect 807 317 811 318
rect 903 322 907 323
rect 903 317 907 318
rect 911 322 915 323
rect 911 317 915 318
rect 943 322 947 323
rect 943 317 947 318
rect 999 322 1003 323
rect 999 317 1003 318
rect 1031 322 1035 323
rect 1031 317 1035 318
rect 1047 322 1051 323
rect 1047 317 1051 318
rect 1063 322 1067 323
rect 1063 317 1067 318
rect 1103 322 1107 323
rect 1103 317 1107 318
rect 1111 322 1115 323
rect 1111 317 1115 318
rect 1199 322 1203 323
rect 1199 317 1203 318
rect 1231 322 1235 323
rect 1231 317 1235 318
rect 1287 322 1291 323
rect 1287 317 1291 318
rect 1319 322 1323 323
rect 1319 317 1323 318
rect 1351 322 1355 323
rect 1351 317 1355 318
rect 1383 322 1387 323
rect 1383 317 1387 318
rect 1415 322 1419 323
rect 1415 317 1419 318
rect 1439 322 1443 323
rect 1439 317 1443 318
rect 1447 322 1451 323
rect 1447 317 1451 318
rect 1479 322 1483 323
rect 1479 317 1483 318
rect 1519 322 1523 323
rect 1519 317 1523 318
rect 1559 322 1563 323
rect 1559 317 1563 318
rect 1591 322 1595 323
rect 1591 317 1595 318
rect 1623 322 1627 323
rect 1623 317 1627 318
rect 1655 322 1659 323
rect 1655 317 1659 318
rect 1695 322 1699 323
rect 1695 317 1699 318
rect 112 302 114 317
rect 136 304 138 317
rect 168 304 170 317
rect 200 304 202 317
rect 232 304 234 317
rect 264 304 266 317
rect 296 304 298 317
rect 328 304 330 317
rect 360 304 362 317
rect 392 304 394 317
rect 424 304 426 317
rect 456 304 458 317
rect 488 304 490 317
rect 520 304 522 317
rect 552 304 554 317
rect 600 307 602 317
rect 704 307 706 317
rect 808 307 810 317
rect 912 307 914 317
rect 598 306 604 307
rect 134 303 140 304
rect 110 301 116 302
rect 110 297 111 301
rect 115 297 116 301
rect 134 299 135 303
rect 139 299 140 303
rect 134 298 140 299
rect 166 303 172 304
rect 166 299 167 303
rect 171 299 172 303
rect 166 298 172 299
rect 198 303 204 304
rect 198 299 199 303
rect 203 299 204 303
rect 198 298 204 299
rect 230 303 236 304
rect 230 299 231 303
rect 235 299 236 303
rect 230 298 236 299
rect 262 303 268 304
rect 262 299 263 303
rect 267 299 268 303
rect 262 298 268 299
rect 294 303 300 304
rect 294 299 295 303
rect 299 299 300 303
rect 294 298 300 299
rect 326 303 332 304
rect 326 299 327 303
rect 331 299 332 303
rect 326 298 332 299
rect 358 303 364 304
rect 358 299 359 303
rect 363 299 364 303
rect 358 298 364 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 422 303 428 304
rect 422 299 423 303
rect 427 299 428 303
rect 422 298 428 299
rect 454 303 460 304
rect 454 299 455 303
rect 459 299 460 303
rect 454 298 460 299
rect 486 303 492 304
rect 486 299 487 303
rect 491 299 492 303
rect 486 298 492 299
rect 518 303 524 304
rect 518 299 519 303
rect 523 299 524 303
rect 518 298 524 299
rect 550 303 556 304
rect 550 299 551 303
rect 555 299 556 303
rect 598 302 599 306
rect 603 302 604 306
rect 598 301 604 302
rect 702 306 708 307
rect 702 302 703 306
rect 707 302 708 306
rect 702 301 708 302
rect 806 306 812 307
rect 806 302 807 306
rect 811 302 812 306
rect 806 301 812 302
rect 910 306 916 307
rect 910 302 911 306
rect 915 302 916 306
rect 1000 304 1002 317
rect 1032 304 1034 317
rect 1064 304 1066 317
rect 1112 307 1114 317
rect 1200 312 1202 317
rect 1198 311 1204 312
rect 1198 307 1199 311
rect 1203 307 1204 311
rect 1110 306 1116 307
rect 1198 306 1204 307
rect 910 301 916 302
rect 998 303 1004 304
rect 550 298 556 299
rect 998 299 999 303
rect 1003 299 1004 303
rect 998 298 1004 299
rect 1030 303 1036 304
rect 1030 299 1031 303
rect 1035 299 1036 303
rect 1030 298 1036 299
rect 1062 303 1068 304
rect 1062 299 1063 303
rect 1067 299 1068 303
rect 1110 302 1111 306
rect 1115 302 1116 306
rect 1288 305 1290 317
rect 1110 301 1116 302
rect 1286 304 1292 305
rect 1320 304 1322 317
rect 1352 304 1354 317
rect 1384 304 1386 317
rect 1416 304 1418 317
rect 1448 304 1450 317
rect 1480 304 1482 317
rect 1520 304 1522 317
rect 1560 304 1562 317
rect 1592 304 1594 317
rect 1624 304 1626 317
rect 1656 304 1658 317
rect 1286 300 1287 304
rect 1291 300 1292 304
rect 1286 299 1292 300
rect 1318 303 1324 304
rect 1318 299 1319 303
rect 1323 299 1324 303
rect 1062 298 1068 299
rect 1318 298 1324 299
rect 1350 303 1356 304
rect 1350 299 1351 303
rect 1355 299 1356 303
rect 1350 298 1356 299
rect 1382 303 1388 304
rect 1382 299 1383 303
rect 1387 299 1388 303
rect 1382 298 1388 299
rect 1414 303 1420 304
rect 1414 299 1415 303
rect 1419 299 1420 303
rect 1414 298 1420 299
rect 1446 303 1452 304
rect 1446 299 1447 303
rect 1451 299 1452 303
rect 1446 298 1452 299
rect 1478 303 1484 304
rect 1478 299 1479 303
rect 1483 299 1484 303
rect 1478 298 1484 299
rect 1518 303 1524 304
rect 1518 299 1519 303
rect 1523 299 1524 303
rect 1518 298 1524 299
rect 1558 303 1564 304
rect 1558 299 1559 303
rect 1563 299 1564 303
rect 1558 298 1564 299
rect 1590 303 1596 304
rect 1590 299 1591 303
rect 1595 299 1596 303
rect 1590 298 1596 299
rect 1622 303 1628 304
rect 1622 299 1623 303
rect 1627 299 1628 303
rect 1622 298 1628 299
rect 1654 303 1660 304
rect 1654 299 1655 303
rect 1659 299 1660 303
rect 1696 302 1698 317
rect 1654 298 1660 299
rect 1694 301 1700 302
rect 110 296 116 297
rect 1694 297 1695 301
rect 1699 297 1700 301
rect 1694 296 1700 297
rect 134 286 140 287
rect 110 284 116 285
rect 110 280 111 284
rect 115 280 116 284
rect 134 282 135 286
rect 139 282 140 286
rect 134 281 140 282
rect 166 286 172 287
rect 166 282 167 286
rect 171 282 172 286
rect 166 281 172 282
rect 198 286 204 287
rect 198 282 199 286
rect 203 282 204 286
rect 198 281 204 282
rect 230 286 236 287
rect 230 282 231 286
rect 235 282 236 286
rect 230 281 236 282
rect 262 286 268 287
rect 262 282 263 286
rect 267 282 268 286
rect 262 281 268 282
rect 294 286 300 287
rect 294 282 295 286
rect 299 282 300 286
rect 294 281 300 282
rect 326 286 332 287
rect 326 282 327 286
rect 331 282 332 286
rect 326 281 332 282
rect 358 286 364 287
rect 358 282 359 286
rect 363 282 364 286
rect 358 281 364 282
rect 390 286 396 287
rect 390 282 391 286
rect 395 282 396 286
rect 390 281 396 282
rect 422 286 428 287
rect 422 282 423 286
rect 427 282 428 286
rect 422 281 428 282
rect 454 286 460 287
rect 454 282 455 286
rect 459 282 460 286
rect 454 281 460 282
rect 486 286 492 287
rect 486 282 487 286
rect 491 282 492 286
rect 486 281 492 282
rect 518 286 524 287
rect 518 282 519 286
rect 523 282 524 286
rect 518 281 524 282
rect 550 286 556 287
rect 550 282 551 286
rect 555 282 556 286
rect 550 281 556 282
rect 998 286 1004 287
rect 998 282 999 286
rect 1003 282 1004 286
rect 998 281 1004 282
rect 1030 286 1036 287
rect 1030 282 1031 286
rect 1035 282 1036 286
rect 1030 281 1036 282
rect 1062 286 1068 287
rect 1062 282 1063 286
rect 1067 282 1068 286
rect 1318 286 1324 287
rect 1318 282 1319 286
rect 1323 282 1324 286
rect 1062 281 1068 282
rect 1286 281 1292 282
rect 1318 281 1324 282
rect 1350 286 1356 287
rect 1350 282 1351 286
rect 1355 282 1356 286
rect 1350 281 1356 282
rect 1382 286 1388 287
rect 1382 282 1383 286
rect 1387 282 1388 286
rect 1382 281 1388 282
rect 1414 286 1420 287
rect 1414 282 1415 286
rect 1419 282 1420 286
rect 1414 281 1420 282
rect 1446 286 1452 287
rect 1446 282 1447 286
rect 1451 282 1452 286
rect 1446 281 1452 282
rect 1478 286 1484 287
rect 1478 282 1479 286
rect 1483 282 1484 286
rect 1478 281 1484 282
rect 1518 286 1524 287
rect 1518 282 1519 286
rect 1523 282 1524 286
rect 1518 281 1524 282
rect 1558 286 1564 287
rect 1558 282 1559 286
rect 1563 282 1564 286
rect 1558 281 1564 282
rect 1590 286 1596 287
rect 1590 282 1591 286
rect 1595 282 1596 286
rect 1590 281 1596 282
rect 1622 286 1628 287
rect 1622 282 1623 286
rect 1627 282 1628 286
rect 1622 281 1628 282
rect 1654 286 1660 287
rect 1654 282 1655 286
rect 1659 282 1660 286
rect 1654 281 1660 282
rect 1694 284 1700 285
rect 110 279 116 280
rect 112 251 114 279
rect 136 251 138 281
rect 168 251 170 281
rect 200 251 202 281
rect 232 251 234 281
rect 264 251 266 281
rect 296 251 298 281
rect 328 251 330 281
rect 360 251 362 281
rect 392 251 394 281
rect 424 251 426 281
rect 456 251 458 281
rect 488 251 490 281
rect 520 251 522 281
rect 552 251 554 281
rect 598 265 604 266
rect 598 261 599 265
rect 603 261 604 265
rect 598 260 604 261
rect 702 265 708 266
rect 702 261 703 265
rect 707 261 708 265
rect 702 260 708 261
rect 806 265 812 266
rect 806 261 807 265
rect 811 261 812 265
rect 806 260 812 261
rect 910 265 916 266
rect 910 261 911 265
rect 915 261 916 265
rect 910 260 916 261
rect 600 251 602 260
rect 704 251 706 260
rect 808 251 810 260
rect 912 251 914 260
rect 1000 251 1002 281
rect 1032 251 1034 281
rect 1064 251 1066 281
rect 1286 277 1287 281
rect 1291 277 1292 281
rect 1286 276 1292 277
rect 1206 271 1212 272
rect 1206 267 1207 271
rect 1211 267 1212 271
rect 1206 266 1212 267
rect 1110 265 1116 266
rect 1110 261 1111 265
rect 1115 261 1116 265
rect 1110 260 1116 261
rect 1112 251 1114 260
rect 1208 251 1210 266
rect 1288 251 1290 276
rect 1320 251 1322 281
rect 1352 251 1354 281
rect 1384 251 1386 281
rect 1416 251 1418 281
rect 1448 251 1450 281
rect 1480 251 1482 281
rect 1520 251 1522 281
rect 1560 251 1562 281
rect 1592 251 1594 281
rect 1624 251 1626 281
rect 1656 251 1658 281
rect 1694 280 1695 284
rect 1699 280 1700 284
rect 1694 279 1700 280
rect 1696 251 1698 279
rect 111 250 115 251
rect 111 245 115 246
rect 135 250 139 251
rect 135 245 139 246
rect 167 250 171 251
rect 167 245 171 246
rect 183 250 187 251
rect 183 245 187 246
rect 199 250 203 251
rect 199 245 203 246
rect 215 250 219 251
rect 215 245 219 246
rect 231 250 235 251
rect 231 245 235 246
rect 247 250 251 251
rect 247 245 251 246
rect 263 250 267 251
rect 263 245 267 246
rect 279 250 283 251
rect 279 245 283 246
rect 295 250 299 251
rect 295 245 299 246
rect 311 250 315 251
rect 311 245 315 246
rect 327 250 331 251
rect 327 245 331 246
rect 343 250 347 251
rect 343 245 347 246
rect 359 250 363 251
rect 359 245 363 246
rect 375 250 379 251
rect 375 245 379 246
rect 391 250 395 251
rect 391 245 395 246
rect 407 250 411 251
rect 407 245 411 246
rect 423 250 427 251
rect 423 245 427 246
rect 439 250 443 251
rect 439 245 443 246
rect 455 250 459 251
rect 455 245 459 246
rect 471 250 475 251
rect 471 245 475 246
rect 487 250 491 251
rect 487 245 491 246
rect 503 250 507 251
rect 503 245 507 246
rect 519 250 523 251
rect 519 245 523 246
rect 535 250 539 251
rect 535 245 539 246
rect 551 250 555 251
rect 551 245 555 246
rect 567 250 571 251
rect 567 245 571 246
rect 599 250 603 251
rect 599 245 603 246
rect 639 250 643 251
rect 639 245 643 246
rect 695 250 699 251
rect 695 245 699 246
rect 703 250 707 251
rect 703 245 707 246
rect 791 250 795 251
rect 791 245 795 246
rect 807 250 811 251
rect 807 245 811 246
rect 839 250 843 251
rect 839 245 843 246
rect 911 250 915 251
rect 911 245 915 246
rect 919 250 923 251
rect 919 245 923 246
rect 967 250 971 251
rect 967 245 971 246
rect 999 250 1003 251
rect 999 245 1003 246
rect 1031 250 1035 251
rect 1031 245 1035 246
rect 1063 250 1067 251
rect 1063 245 1067 246
rect 1103 250 1107 251
rect 1103 245 1107 246
rect 1111 250 1115 251
rect 1111 245 1115 246
rect 1143 250 1147 251
rect 1143 245 1147 246
rect 1183 250 1187 251
rect 1183 245 1187 246
rect 1207 250 1211 251
rect 1207 245 1211 246
rect 1223 250 1227 251
rect 1223 245 1227 246
rect 1263 250 1267 251
rect 1263 245 1267 246
rect 1287 250 1291 251
rect 1287 245 1291 246
rect 1303 250 1307 251
rect 1303 245 1307 246
rect 1319 250 1323 251
rect 1319 245 1323 246
rect 1343 250 1347 251
rect 1343 245 1347 246
rect 1351 250 1355 251
rect 1351 245 1355 246
rect 1375 250 1379 251
rect 1375 245 1379 246
rect 1383 250 1387 251
rect 1383 245 1387 246
rect 1407 250 1411 251
rect 1407 245 1411 246
rect 1415 250 1419 251
rect 1415 245 1419 246
rect 1439 250 1443 251
rect 1439 245 1443 246
rect 1447 250 1451 251
rect 1447 245 1451 246
rect 1479 250 1483 251
rect 1479 245 1483 246
rect 1519 250 1523 251
rect 1519 245 1523 246
rect 1559 250 1563 251
rect 1559 245 1563 246
rect 1591 250 1595 251
rect 1591 245 1595 246
rect 1623 250 1627 251
rect 1623 245 1627 246
rect 1655 250 1659 251
rect 1655 245 1659 246
rect 1695 250 1699 251
rect 1695 245 1699 246
rect 112 217 114 245
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 184 215 186 245
rect 216 215 218 245
rect 248 215 250 245
rect 280 215 282 245
rect 312 215 314 245
rect 344 215 346 245
rect 376 215 378 245
rect 408 215 410 245
rect 440 215 442 245
rect 472 215 474 245
rect 504 215 506 245
rect 536 215 538 245
rect 568 215 570 245
rect 600 215 602 245
rect 640 215 642 245
rect 696 236 698 245
rect 694 235 700 236
rect 694 231 695 235
rect 699 231 700 235
rect 694 230 700 231
rect 792 215 794 245
rect 840 230 842 245
rect 838 229 844 230
rect 838 225 839 229
rect 843 225 844 229
rect 838 224 844 225
rect 920 220 922 245
rect 968 236 970 245
rect 966 235 972 236
rect 966 231 967 235
rect 971 231 972 235
rect 966 230 972 231
rect 918 219 924 220
rect 918 215 919 219
rect 923 215 924 219
rect 1064 215 1066 245
rect 1104 215 1106 245
rect 1144 215 1146 245
rect 1184 215 1186 245
rect 1224 215 1226 245
rect 1264 215 1266 245
rect 1304 215 1306 245
rect 1344 215 1346 245
rect 1376 215 1378 245
rect 1408 215 1410 245
rect 1440 215 1442 245
rect 1480 215 1482 245
rect 1520 215 1522 245
rect 1560 215 1562 245
rect 1592 215 1594 245
rect 1624 215 1626 245
rect 1656 215 1658 245
rect 1696 217 1698 245
rect 1694 216 1700 217
rect 110 211 116 212
rect 182 214 188 215
rect 182 210 183 214
rect 187 210 188 214
rect 182 209 188 210
rect 214 214 220 215
rect 214 210 215 214
rect 219 210 220 214
rect 214 209 220 210
rect 246 214 252 215
rect 246 210 247 214
rect 251 210 252 214
rect 246 209 252 210
rect 278 214 284 215
rect 278 210 279 214
rect 283 210 284 214
rect 278 209 284 210
rect 310 214 316 215
rect 310 210 311 214
rect 315 210 316 214
rect 310 209 316 210
rect 342 214 348 215
rect 342 210 343 214
rect 347 210 348 214
rect 342 209 348 210
rect 374 214 380 215
rect 374 210 375 214
rect 379 210 380 214
rect 374 209 380 210
rect 406 214 412 215
rect 406 210 407 214
rect 411 210 412 214
rect 406 209 412 210
rect 438 214 444 215
rect 438 210 439 214
rect 443 210 444 214
rect 438 209 444 210
rect 470 214 476 215
rect 470 210 471 214
rect 475 210 476 214
rect 470 209 476 210
rect 502 214 508 215
rect 502 210 503 214
rect 507 210 508 214
rect 502 209 508 210
rect 534 214 540 215
rect 534 210 535 214
rect 539 210 540 214
rect 534 209 540 210
rect 566 214 572 215
rect 566 210 567 214
rect 571 210 572 214
rect 566 209 572 210
rect 598 214 604 215
rect 598 210 599 214
rect 603 210 604 214
rect 598 209 604 210
rect 638 214 644 215
rect 638 210 639 214
rect 643 210 644 214
rect 638 209 644 210
rect 790 214 796 215
rect 918 214 924 215
rect 1062 214 1068 215
rect 790 210 791 214
rect 795 210 796 214
rect 790 209 796 210
rect 1062 210 1063 214
rect 1067 210 1068 214
rect 1062 209 1068 210
rect 1102 214 1108 215
rect 1102 210 1103 214
rect 1107 210 1108 214
rect 1102 209 1108 210
rect 1142 214 1148 215
rect 1142 210 1143 214
rect 1147 210 1148 214
rect 1142 209 1148 210
rect 1182 214 1188 215
rect 1182 210 1183 214
rect 1187 210 1188 214
rect 1182 209 1188 210
rect 1222 214 1228 215
rect 1222 210 1223 214
rect 1227 210 1228 214
rect 1222 209 1228 210
rect 1262 214 1268 215
rect 1262 210 1263 214
rect 1267 210 1268 214
rect 1262 209 1268 210
rect 1302 214 1308 215
rect 1302 210 1303 214
rect 1307 210 1308 214
rect 1302 209 1308 210
rect 1342 214 1348 215
rect 1342 210 1343 214
rect 1347 210 1348 214
rect 1342 209 1348 210
rect 1374 214 1380 215
rect 1374 210 1375 214
rect 1379 210 1380 214
rect 1374 209 1380 210
rect 1406 214 1412 215
rect 1406 210 1407 214
rect 1411 210 1412 214
rect 1406 209 1412 210
rect 1438 214 1444 215
rect 1438 210 1439 214
rect 1443 210 1444 214
rect 1438 209 1444 210
rect 1478 214 1484 215
rect 1478 210 1479 214
rect 1483 210 1484 214
rect 1478 209 1484 210
rect 1518 214 1524 215
rect 1518 210 1519 214
rect 1523 210 1524 214
rect 1518 209 1524 210
rect 1558 214 1564 215
rect 1558 210 1559 214
rect 1563 210 1564 214
rect 1558 209 1564 210
rect 1590 214 1596 215
rect 1590 210 1591 214
rect 1595 210 1596 214
rect 1590 209 1596 210
rect 1622 214 1628 215
rect 1622 210 1623 214
rect 1627 210 1628 214
rect 1622 209 1628 210
rect 1654 214 1660 215
rect 1654 210 1655 214
rect 1659 210 1660 214
rect 1694 212 1695 216
rect 1699 212 1700 216
rect 1694 211 1700 212
rect 1654 209 1660 210
rect 110 199 116 200
rect 110 195 111 199
rect 115 195 116 199
rect 1694 199 1700 200
rect 110 194 116 195
rect 182 197 188 198
rect 112 175 114 194
rect 182 193 183 197
rect 187 193 188 197
rect 182 192 188 193
rect 214 197 220 198
rect 214 193 215 197
rect 219 193 220 197
rect 214 192 220 193
rect 246 197 252 198
rect 246 193 247 197
rect 251 193 252 197
rect 246 192 252 193
rect 278 197 284 198
rect 278 193 279 197
rect 283 193 284 197
rect 278 192 284 193
rect 310 197 316 198
rect 310 193 311 197
rect 315 193 316 197
rect 310 192 316 193
rect 342 197 348 198
rect 342 193 343 197
rect 347 193 348 197
rect 342 192 348 193
rect 374 197 380 198
rect 374 193 375 197
rect 379 193 380 197
rect 374 192 380 193
rect 406 197 412 198
rect 406 193 407 197
rect 411 193 412 197
rect 406 192 412 193
rect 438 197 444 198
rect 438 193 439 197
rect 443 193 444 197
rect 438 192 444 193
rect 470 197 476 198
rect 470 193 471 197
rect 475 193 476 197
rect 470 192 476 193
rect 502 197 508 198
rect 502 193 503 197
rect 507 193 508 197
rect 502 192 508 193
rect 534 197 540 198
rect 534 193 535 197
rect 539 193 540 197
rect 534 192 540 193
rect 566 197 572 198
rect 566 193 567 197
rect 571 193 572 197
rect 566 192 572 193
rect 598 197 604 198
rect 598 193 599 197
rect 603 193 604 197
rect 598 192 604 193
rect 638 197 644 198
rect 638 193 639 197
rect 643 193 644 197
rect 790 197 796 198
rect 1062 197 1068 198
rect 638 192 644 193
rect 694 194 700 195
rect 184 175 186 192
rect 216 175 218 192
rect 248 175 250 192
rect 280 175 282 192
rect 312 175 314 192
rect 344 175 346 192
rect 376 175 378 192
rect 408 175 410 192
rect 440 175 442 192
rect 472 175 474 192
rect 504 175 506 192
rect 536 175 538 192
rect 568 175 570 192
rect 600 175 602 192
rect 640 175 642 192
rect 694 190 695 194
rect 699 190 700 194
rect 790 193 791 197
rect 795 193 796 197
rect 790 192 796 193
rect 918 196 924 197
rect 918 192 919 196
rect 923 192 924 196
rect 694 189 700 190
rect 696 175 698 189
rect 792 175 794 192
rect 918 191 924 192
rect 966 194 972 195
rect 830 189 836 190
rect 830 185 831 189
rect 835 185 836 189
rect 830 184 836 185
rect 832 175 834 184
rect 920 175 922 191
rect 966 190 967 194
rect 971 190 972 194
rect 1062 193 1063 197
rect 1067 193 1068 197
rect 1062 192 1068 193
rect 1102 197 1108 198
rect 1102 193 1103 197
rect 1107 193 1108 197
rect 1102 192 1108 193
rect 1142 197 1148 198
rect 1142 193 1143 197
rect 1147 193 1148 197
rect 1142 192 1148 193
rect 1182 197 1188 198
rect 1182 193 1183 197
rect 1187 193 1188 197
rect 1182 192 1188 193
rect 1222 197 1228 198
rect 1222 193 1223 197
rect 1227 193 1228 197
rect 1222 192 1228 193
rect 1262 197 1268 198
rect 1262 193 1263 197
rect 1267 193 1268 197
rect 1262 192 1268 193
rect 1302 197 1308 198
rect 1302 193 1303 197
rect 1307 193 1308 197
rect 1302 192 1308 193
rect 1342 197 1348 198
rect 1342 193 1343 197
rect 1347 193 1348 197
rect 1342 192 1348 193
rect 1374 197 1380 198
rect 1374 193 1375 197
rect 1379 193 1380 197
rect 1374 192 1380 193
rect 1406 197 1412 198
rect 1406 193 1407 197
rect 1411 193 1412 197
rect 1406 192 1412 193
rect 1438 197 1444 198
rect 1438 193 1439 197
rect 1443 193 1444 197
rect 1438 192 1444 193
rect 1478 197 1484 198
rect 1478 193 1479 197
rect 1483 193 1484 197
rect 1478 192 1484 193
rect 1518 197 1524 198
rect 1518 193 1519 197
rect 1523 193 1524 197
rect 1518 192 1524 193
rect 1558 197 1564 198
rect 1558 193 1559 197
rect 1563 193 1564 197
rect 1558 192 1564 193
rect 1590 197 1596 198
rect 1590 193 1591 197
rect 1595 193 1596 197
rect 1590 192 1596 193
rect 1622 197 1628 198
rect 1622 193 1623 197
rect 1627 193 1628 197
rect 1622 192 1628 193
rect 1654 197 1660 198
rect 1654 193 1655 197
rect 1659 193 1660 197
rect 1694 195 1695 199
rect 1699 195 1700 199
rect 1694 194 1700 195
rect 1654 192 1660 193
rect 966 189 972 190
rect 968 175 970 189
rect 1064 175 1066 192
rect 1104 175 1106 192
rect 1144 175 1146 192
rect 1184 175 1186 192
rect 1224 175 1226 192
rect 1264 175 1266 192
rect 1304 175 1306 192
rect 1344 175 1346 192
rect 1376 175 1378 192
rect 1408 175 1410 192
rect 1440 175 1442 192
rect 1480 175 1482 192
rect 1520 175 1522 192
rect 1560 175 1562 192
rect 1592 175 1594 192
rect 1624 175 1626 192
rect 1656 175 1658 192
rect 1696 175 1698 194
rect 111 174 115 175
rect 111 169 115 170
rect 135 174 139 175
rect 112 166 114 169
rect 135 168 139 170
rect 167 174 171 175
rect 167 168 171 170
rect 183 174 187 175
rect 183 169 187 170
rect 215 174 219 175
rect 215 168 219 170
rect 247 174 251 175
rect 247 169 251 170
rect 263 174 267 175
rect 263 168 267 170
rect 279 174 283 175
rect 279 169 283 170
rect 311 174 315 175
rect 311 168 315 170
rect 343 174 347 175
rect 343 169 347 170
rect 367 174 371 175
rect 367 168 371 170
rect 375 174 379 175
rect 375 169 379 170
rect 407 174 411 175
rect 407 169 411 170
rect 415 174 419 175
rect 415 168 419 170
rect 439 174 443 175
rect 439 169 443 170
rect 471 174 475 175
rect 471 168 475 170
rect 503 174 507 175
rect 503 169 507 170
rect 535 174 539 175
rect 535 168 539 170
rect 567 174 571 175
rect 567 169 571 170
rect 599 174 603 175
rect 599 169 603 170
rect 607 174 611 175
rect 607 168 611 170
rect 639 174 643 175
rect 639 169 643 170
rect 687 174 691 175
rect 687 168 691 170
rect 695 174 699 175
rect 695 169 699 170
rect 775 174 779 175
rect 775 168 779 170
rect 791 174 795 175
rect 791 169 795 170
rect 831 174 835 175
rect 831 169 835 170
rect 863 174 867 175
rect 863 168 867 170
rect 919 174 923 175
rect 919 169 923 170
rect 959 174 963 175
rect 959 168 963 170
rect 967 174 971 175
rect 967 169 971 170
rect 1055 174 1059 175
rect 1055 168 1059 170
rect 1063 174 1067 175
rect 1063 169 1067 170
rect 1103 174 1107 175
rect 1103 169 1107 170
rect 1143 174 1147 175
rect 1143 169 1147 170
rect 1151 174 1155 175
rect 1151 168 1155 170
rect 1183 174 1187 175
rect 1183 169 1187 170
rect 1223 174 1227 175
rect 1223 169 1227 170
rect 1239 174 1243 175
rect 1239 168 1243 170
rect 1263 174 1267 175
rect 1263 169 1267 170
rect 1303 174 1307 175
rect 1303 169 1307 170
rect 1327 174 1331 175
rect 1327 168 1331 170
rect 1343 174 1347 175
rect 1343 169 1347 170
rect 1375 174 1379 175
rect 1375 169 1379 170
rect 1407 174 1411 175
rect 1407 169 1411 170
rect 1415 174 1419 175
rect 1415 168 1419 170
rect 1439 174 1443 175
rect 1439 169 1443 170
rect 1479 174 1483 175
rect 1479 169 1483 170
rect 1503 174 1507 175
rect 1503 168 1507 170
rect 1519 174 1523 175
rect 1519 169 1523 170
rect 1559 174 1563 175
rect 1559 169 1563 170
rect 1591 174 1595 175
rect 1591 168 1595 170
rect 1623 174 1627 175
rect 1623 169 1627 170
rect 1655 174 1659 175
rect 1655 168 1659 170
rect 1695 174 1699 175
rect 1695 169 1699 170
rect 134 167 140 168
rect 110 165 116 166
rect 110 161 111 165
rect 115 161 116 165
rect 134 163 135 167
rect 139 163 140 167
rect 134 162 140 163
rect 166 167 172 168
rect 166 163 167 167
rect 171 163 172 167
rect 166 162 172 163
rect 214 167 220 168
rect 214 163 215 167
rect 219 163 220 167
rect 214 162 220 163
rect 262 167 268 168
rect 262 163 263 167
rect 267 163 268 167
rect 262 162 268 163
rect 310 167 316 168
rect 310 163 311 167
rect 315 163 316 167
rect 310 162 316 163
rect 366 167 372 168
rect 366 163 367 167
rect 371 163 372 167
rect 366 162 372 163
rect 414 167 420 168
rect 414 163 415 167
rect 419 163 420 167
rect 414 162 420 163
rect 470 167 476 168
rect 470 163 471 167
rect 475 163 476 167
rect 470 162 476 163
rect 534 167 540 168
rect 534 163 535 167
rect 539 163 540 167
rect 534 162 540 163
rect 606 167 612 168
rect 606 163 607 167
rect 611 163 612 167
rect 606 162 612 163
rect 686 167 692 168
rect 686 163 687 167
rect 691 163 692 167
rect 686 162 692 163
rect 774 167 780 168
rect 774 163 775 167
rect 779 163 780 167
rect 774 162 780 163
rect 862 167 868 168
rect 862 163 863 167
rect 867 163 868 167
rect 862 162 868 163
rect 958 167 964 168
rect 958 163 959 167
rect 963 163 964 167
rect 958 162 964 163
rect 1054 167 1060 168
rect 1054 163 1055 167
rect 1059 163 1060 167
rect 1054 162 1060 163
rect 1150 167 1156 168
rect 1150 163 1151 167
rect 1155 163 1156 167
rect 1150 162 1156 163
rect 1238 167 1244 168
rect 1238 163 1239 167
rect 1243 163 1244 167
rect 1238 162 1244 163
rect 1326 167 1332 168
rect 1326 163 1327 167
rect 1331 163 1332 167
rect 1326 162 1332 163
rect 1414 167 1420 168
rect 1414 163 1415 167
rect 1419 163 1420 167
rect 1414 162 1420 163
rect 1502 167 1508 168
rect 1502 163 1503 167
rect 1507 163 1508 167
rect 1502 162 1508 163
rect 1590 167 1596 168
rect 1590 163 1591 167
rect 1595 163 1596 167
rect 1590 162 1596 163
rect 1654 167 1660 168
rect 1654 163 1655 167
rect 1659 163 1660 167
rect 1696 166 1698 169
rect 1654 162 1660 163
rect 1694 165 1700 166
rect 110 160 116 161
rect 1694 161 1695 165
rect 1699 161 1700 165
rect 1694 160 1700 161
rect 134 150 140 151
rect 110 148 116 149
rect 110 144 111 148
rect 115 144 116 148
rect 134 146 135 150
rect 139 146 140 150
rect 134 145 140 146
rect 166 150 172 151
rect 166 146 167 150
rect 171 146 172 150
rect 166 145 172 146
rect 214 150 220 151
rect 214 146 215 150
rect 219 146 220 150
rect 214 145 220 146
rect 262 150 268 151
rect 262 146 263 150
rect 267 146 268 150
rect 262 145 268 146
rect 310 150 316 151
rect 310 146 311 150
rect 315 146 316 150
rect 310 145 316 146
rect 366 150 372 151
rect 366 146 367 150
rect 371 146 372 150
rect 366 145 372 146
rect 414 150 420 151
rect 414 146 415 150
rect 419 146 420 150
rect 414 145 420 146
rect 470 150 476 151
rect 470 146 471 150
rect 475 146 476 150
rect 470 145 476 146
rect 534 150 540 151
rect 534 146 535 150
rect 539 146 540 150
rect 534 145 540 146
rect 606 150 612 151
rect 606 146 607 150
rect 611 146 612 150
rect 606 145 612 146
rect 686 150 692 151
rect 686 146 687 150
rect 691 146 692 150
rect 686 145 692 146
rect 774 150 780 151
rect 774 146 775 150
rect 779 146 780 150
rect 774 145 780 146
rect 862 150 868 151
rect 862 146 863 150
rect 867 146 868 150
rect 862 145 868 146
rect 958 150 964 151
rect 958 146 959 150
rect 963 146 964 150
rect 958 145 964 146
rect 1054 150 1060 151
rect 1054 146 1055 150
rect 1059 146 1060 150
rect 1054 145 1060 146
rect 1150 150 1156 151
rect 1150 146 1151 150
rect 1155 146 1156 150
rect 1150 145 1156 146
rect 1238 150 1244 151
rect 1238 146 1239 150
rect 1243 146 1244 150
rect 1238 145 1244 146
rect 1326 150 1332 151
rect 1326 146 1327 150
rect 1331 146 1332 150
rect 1326 145 1332 146
rect 1414 150 1420 151
rect 1414 146 1415 150
rect 1419 146 1420 150
rect 1414 145 1420 146
rect 1502 150 1508 151
rect 1502 146 1503 150
rect 1507 146 1508 150
rect 1502 145 1508 146
rect 1590 150 1596 151
rect 1590 146 1591 150
rect 1595 146 1596 150
rect 1590 145 1596 146
rect 1654 150 1660 151
rect 1654 146 1655 150
rect 1659 146 1660 150
rect 1654 145 1660 146
rect 1694 148 1700 149
rect 110 143 116 144
rect 112 123 114 143
rect 136 123 138 145
rect 168 123 170 145
rect 216 123 218 145
rect 264 123 266 145
rect 312 123 314 145
rect 368 123 370 145
rect 416 123 418 145
rect 472 123 474 145
rect 536 123 538 145
rect 608 123 610 145
rect 688 123 690 145
rect 776 123 778 145
rect 864 123 866 145
rect 960 123 962 145
rect 1056 123 1058 145
rect 1152 123 1154 145
rect 1240 123 1242 145
rect 1328 123 1330 145
rect 1416 123 1418 145
rect 1504 123 1506 145
rect 1592 123 1594 145
rect 1656 123 1658 145
rect 1694 144 1695 148
rect 1699 144 1700 148
rect 1694 143 1700 144
rect 1696 123 1698 143
rect 111 122 115 123
rect 111 117 115 118
rect 135 122 139 123
rect 135 117 139 118
rect 167 122 171 123
rect 167 117 171 118
rect 199 122 203 123
rect 199 117 203 118
rect 215 122 219 123
rect 215 117 219 118
rect 231 122 235 123
rect 231 117 235 118
rect 263 122 267 123
rect 263 117 267 118
rect 295 122 299 123
rect 295 117 299 118
rect 311 122 315 123
rect 311 117 315 118
rect 327 122 331 123
rect 327 117 331 118
rect 359 122 363 123
rect 359 117 363 118
rect 367 122 371 123
rect 367 117 371 118
rect 391 122 395 123
rect 391 117 395 118
rect 415 122 419 123
rect 415 117 419 118
rect 423 122 427 123
rect 423 117 427 118
rect 455 122 459 123
rect 455 117 459 118
rect 471 122 475 123
rect 471 117 475 118
rect 487 122 491 123
rect 487 117 491 118
rect 519 122 523 123
rect 519 117 523 118
rect 535 122 539 123
rect 535 117 539 118
rect 551 122 555 123
rect 551 117 555 118
rect 607 122 611 123
rect 607 117 611 118
rect 671 122 675 123
rect 671 117 675 118
rect 687 122 691 123
rect 687 117 691 118
rect 743 122 747 123
rect 743 117 747 118
rect 775 122 779 123
rect 775 117 779 118
rect 823 122 827 123
rect 823 117 827 118
rect 863 122 867 123
rect 863 117 867 118
rect 903 122 907 123
rect 903 117 907 118
rect 959 122 963 123
rect 959 117 963 118
rect 983 122 987 123
rect 983 117 987 118
rect 1055 122 1059 123
rect 1055 117 1059 118
rect 1119 122 1123 123
rect 1119 117 1123 118
rect 1151 122 1155 123
rect 1151 117 1155 118
rect 1175 122 1179 123
rect 1175 117 1179 118
rect 1223 122 1227 123
rect 1223 117 1227 118
rect 1239 122 1243 123
rect 1239 117 1243 118
rect 1271 122 1275 123
rect 1271 117 1275 118
rect 1311 122 1315 123
rect 1311 117 1315 118
rect 1327 122 1331 123
rect 1327 117 1331 118
rect 1343 122 1347 123
rect 1343 117 1347 118
rect 1375 122 1379 123
rect 1375 117 1379 118
rect 1407 122 1411 123
rect 1407 117 1411 118
rect 1415 122 1419 123
rect 1415 117 1419 118
rect 1439 122 1443 123
rect 1439 117 1443 118
rect 1479 122 1483 123
rect 1479 117 1483 118
rect 1503 122 1507 123
rect 1503 117 1507 118
rect 1519 122 1523 123
rect 1519 117 1523 118
rect 1559 122 1563 123
rect 1559 117 1563 118
rect 1591 122 1595 123
rect 1591 117 1595 118
rect 1623 122 1627 123
rect 1623 117 1627 118
rect 1655 122 1659 123
rect 1655 117 1659 118
rect 1695 122 1699 123
rect 1695 117 1699 118
rect 112 109 114 117
rect 110 108 116 109
rect 110 104 111 108
rect 115 104 116 108
rect 136 107 138 117
rect 168 107 170 117
rect 200 107 202 117
rect 232 107 234 117
rect 264 107 266 117
rect 296 107 298 117
rect 328 107 330 117
rect 360 107 362 117
rect 392 107 394 117
rect 424 107 426 117
rect 456 107 458 117
rect 488 107 490 117
rect 520 107 522 117
rect 552 107 554 117
rect 608 107 610 117
rect 672 107 674 117
rect 744 107 746 117
rect 824 107 826 117
rect 904 107 906 117
rect 984 107 986 117
rect 1056 107 1058 117
rect 1120 107 1122 117
rect 1176 107 1178 117
rect 1224 107 1226 117
rect 1272 107 1274 117
rect 1312 107 1314 117
rect 1344 107 1346 117
rect 1376 107 1378 117
rect 1408 107 1410 117
rect 1440 107 1442 117
rect 1480 107 1482 117
rect 1520 107 1522 117
rect 1560 107 1562 117
rect 1592 107 1594 117
rect 1624 107 1626 117
rect 1656 107 1658 117
rect 1696 109 1698 117
rect 1694 108 1700 109
rect 110 103 116 104
rect 134 106 140 107
rect 134 102 135 106
rect 139 102 140 106
rect 134 101 140 102
rect 166 106 172 107
rect 166 102 167 106
rect 171 102 172 106
rect 166 101 172 102
rect 198 106 204 107
rect 198 102 199 106
rect 203 102 204 106
rect 198 101 204 102
rect 230 106 236 107
rect 230 102 231 106
rect 235 102 236 106
rect 230 101 236 102
rect 262 106 268 107
rect 262 102 263 106
rect 267 102 268 106
rect 262 101 268 102
rect 294 106 300 107
rect 294 102 295 106
rect 299 102 300 106
rect 294 101 300 102
rect 326 106 332 107
rect 326 102 327 106
rect 331 102 332 106
rect 326 101 332 102
rect 358 106 364 107
rect 358 102 359 106
rect 363 102 364 106
rect 358 101 364 102
rect 390 106 396 107
rect 390 102 391 106
rect 395 102 396 106
rect 390 101 396 102
rect 422 106 428 107
rect 422 102 423 106
rect 427 102 428 106
rect 422 101 428 102
rect 454 106 460 107
rect 454 102 455 106
rect 459 102 460 106
rect 454 101 460 102
rect 486 106 492 107
rect 486 102 487 106
rect 491 102 492 106
rect 486 101 492 102
rect 518 106 524 107
rect 518 102 519 106
rect 523 102 524 106
rect 518 101 524 102
rect 550 106 556 107
rect 550 102 551 106
rect 555 102 556 106
rect 550 101 556 102
rect 606 106 612 107
rect 606 102 607 106
rect 611 102 612 106
rect 606 101 612 102
rect 670 106 676 107
rect 670 102 671 106
rect 675 102 676 106
rect 670 101 676 102
rect 742 106 748 107
rect 742 102 743 106
rect 747 102 748 106
rect 742 101 748 102
rect 822 106 828 107
rect 822 102 823 106
rect 827 102 828 106
rect 822 101 828 102
rect 902 106 908 107
rect 902 102 903 106
rect 907 102 908 106
rect 902 101 908 102
rect 982 106 988 107
rect 982 102 983 106
rect 987 102 988 106
rect 982 101 988 102
rect 1054 106 1060 107
rect 1054 102 1055 106
rect 1059 102 1060 106
rect 1054 101 1060 102
rect 1118 106 1124 107
rect 1118 102 1119 106
rect 1123 102 1124 106
rect 1118 101 1124 102
rect 1174 106 1180 107
rect 1174 102 1175 106
rect 1179 102 1180 106
rect 1174 101 1180 102
rect 1222 106 1228 107
rect 1222 102 1223 106
rect 1227 102 1228 106
rect 1222 101 1228 102
rect 1270 106 1276 107
rect 1270 102 1271 106
rect 1275 102 1276 106
rect 1270 101 1276 102
rect 1310 106 1316 107
rect 1310 102 1311 106
rect 1315 102 1316 106
rect 1310 101 1316 102
rect 1342 106 1348 107
rect 1342 102 1343 106
rect 1347 102 1348 106
rect 1342 101 1348 102
rect 1374 106 1380 107
rect 1374 102 1375 106
rect 1379 102 1380 106
rect 1374 101 1380 102
rect 1406 106 1412 107
rect 1406 102 1407 106
rect 1411 102 1412 106
rect 1406 101 1412 102
rect 1438 106 1444 107
rect 1438 102 1439 106
rect 1443 102 1444 106
rect 1438 101 1444 102
rect 1478 106 1484 107
rect 1478 102 1479 106
rect 1483 102 1484 106
rect 1478 101 1484 102
rect 1518 106 1524 107
rect 1518 102 1519 106
rect 1523 102 1524 106
rect 1518 101 1524 102
rect 1558 106 1564 107
rect 1558 102 1559 106
rect 1563 102 1564 106
rect 1558 101 1564 102
rect 1590 106 1596 107
rect 1590 102 1591 106
rect 1595 102 1596 106
rect 1590 101 1596 102
rect 1622 106 1628 107
rect 1622 102 1623 106
rect 1627 102 1628 106
rect 1622 101 1628 102
rect 1654 106 1660 107
rect 1654 102 1655 106
rect 1659 102 1660 106
rect 1694 104 1695 108
rect 1699 104 1700 108
rect 1694 103 1700 104
rect 1654 101 1660 102
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 1694 91 1700 92
rect 110 86 116 87
rect 134 89 140 90
rect 112 83 114 86
rect 134 85 135 89
rect 139 85 140 89
rect 134 84 140 85
rect 166 89 172 90
rect 166 85 167 89
rect 171 85 172 89
rect 166 84 172 85
rect 198 89 204 90
rect 198 85 199 89
rect 203 85 204 89
rect 198 84 204 85
rect 230 89 236 90
rect 230 85 231 89
rect 235 85 236 89
rect 230 84 236 85
rect 262 89 268 90
rect 262 85 263 89
rect 267 85 268 89
rect 262 84 268 85
rect 294 89 300 90
rect 294 85 295 89
rect 299 85 300 89
rect 294 84 300 85
rect 326 89 332 90
rect 326 85 327 89
rect 331 85 332 89
rect 326 84 332 85
rect 358 89 364 90
rect 358 85 359 89
rect 363 85 364 89
rect 358 84 364 85
rect 390 89 396 90
rect 390 85 391 89
rect 395 85 396 89
rect 390 84 396 85
rect 422 89 428 90
rect 422 85 423 89
rect 427 85 428 89
rect 422 84 428 85
rect 454 89 460 90
rect 454 85 455 89
rect 459 85 460 89
rect 454 84 460 85
rect 486 89 492 90
rect 486 85 487 89
rect 491 85 492 89
rect 486 84 492 85
rect 518 89 524 90
rect 518 85 519 89
rect 523 85 524 89
rect 518 84 524 85
rect 550 89 556 90
rect 550 85 551 89
rect 555 85 556 89
rect 550 84 556 85
rect 606 89 612 90
rect 606 85 607 89
rect 611 85 612 89
rect 606 84 612 85
rect 670 89 676 90
rect 670 85 671 89
rect 675 85 676 89
rect 670 84 676 85
rect 742 89 748 90
rect 742 85 743 89
rect 747 85 748 89
rect 742 84 748 85
rect 822 89 828 90
rect 822 85 823 89
rect 827 85 828 89
rect 822 84 828 85
rect 902 89 908 90
rect 902 85 903 89
rect 907 85 908 89
rect 902 84 908 85
rect 982 89 988 90
rect 982 85 983 89
rect 987 85 988 89
rect 982 84 988 85
rect 1054 89 1060 90
rect 1054 85 1055 89
rect 1059 85 1060 89
rect 1054 84 1060 85
rect 1118 89 1124 90
rect 1118 85 1119 89
rect 1123 85 1124 89
rect 1118 84 1124 85
rect 1174 89 1180 90
rect 1174 85 1175 89
rect 1179 85 1180 89
rect 1174 84 1180 85
rect 1222 89 1228 90
rect 1222 85 1223 89
rect 1227 85 1228 89
rect 1222 84 1228 85
rect 1270 89 1276 90
rect 1270 85 1271 89
rect 1275 85 1276 89
rect 1270 84 1276 85
rect 1310 89 1316 90
rect 1310 85 1311 89
rect 1315 85 1316 89
rect 1310 84 1316 85
rect 1342 89 1348 90
rect 1342 85 1343 89
rect 1347 85 1348 89
rect 1342 84 1348 85
rect 1374 89 1380 90
rect 1374 85 1375 89
rect 1379 85 1380 89
rect 1374 84 1380 85
rect 1406 89 1412 90
rect 1406 85 1407 89
rect 1411 85 1412 89
rect 1406 84 1412 85
rect 1438 89 1444 90
rect 1438 85 1439 89
rect 1443 85 1444 89
rect 1438 84 1444 85
rect 1478 89 1484 90
rect 1478 85 1479 89
rect 1483 85 1484 89
rect 1478 84 1484 85
rect 1518 89 1524 90
rect 1518 85 1519 89
rect 1523 85 1524 89
rect 1518 84 1524 85
rect 1558 89 1564 90
rect 1558 85 1559 89
rect 1563 85 1564 89
rect 1558 84 1564 85
rect 1590 89 1596 90
rect 1590 85 1591 89
rect 1595 85 1596 89
rect 1590 84 1596 85
rect 1622 89 1628 90
rect 1622 85 1623 89
rect 1627 85 1628 89
rect 1622 84 1628 85
rect 1654 89 1660 90
rect 1654 85 1655 89
rect 1659 85 1660 89
rect 1694 87 1695 91
rect 1699 87 1700 91
rect 1694 86 1700 87
rect 1654 84 1660 85
rect 111 82 115 83
rect 111 77 115 78
rect 135 82 139 84
rect 135 77 139 78
rect 167 82 171 84
rect 167 77 171 78
rect 199 82 203 84
rect 199 77 203 78
rect 231 82 235 84
rect 231 77 235 78
rect 263 82 267 84
rect 263 77 267 78
rect 295 82 299 84
rect 295 77 299 78
rect 327 82 331 84
rect 327 77 331 78
rect 359 82 363 84
rect 359 77 363 78
rect 391 82 395 84
rect 391 77 395 78
rect 423 82 427 84
rect 423 77 427 78
rect 455 82 459 84
rect 455 77 459 78
rect 487 82 491 84
rect 487 77 491 78
rect 519 82 523 84
rect 519 77 523 78
rect 551 82 555 84
rect 551 77 555 78
rect 607 82 611 84
rect 607 77 611 78
rect 671 82 675 84
rect 671 77 675 78
rect 743 82 747 84
rect 743 77 747 78
rect 823 82 827 84
rect 823 77 827 78
rect 903 82 907 84
rect 903 77 907 78
rect 983 82 987 84
rect 983 77 987 78
rect 1055 82 1059 84
rect 1055 77 1059 78
rect 1119 82 1123 84
rect 1119 77 1123 78
rect 1175 82 1179 84
rect 1175 77 1179 78
rect 1223 82 1227 84
rect 1223 77 1227 78
rect 1271 82 1275 84
rect 1271 77 1275 78
rect 1311 82 1315 84
rect 1311 77 1315 78
rect 1343 82 1347 84
rect 1343 77 1347 78
rect 1375 82 1379 84
rect 1375 77 1379 78
rect 1407 82 1411 84
rect 1407 77 1411 78
rect 1439 82 1443 84
rect 1439 77 1443 78
rect 1479 82 1483 84
rect 1479 77 1483 78
rect 1519 82 1523 84
rect 1519 77 1523 78
rect 1559 82 1563 84
rect 1559 77 1563 78
rect 1591 82 1595 84
rect 1591 77 1595 78
rect 1623 82 1627 84
rect 1623 77 1627 78
rect 1655 82 1659 84
rect 1696 83 1698 86
rect 1655 77 1659 78
rect 1695 82 1699 83
rect 1695 77 1699 78
<< m4c >>
rect 111 1758 115 1762
rect 151 1758 155 1762
rect 183 1758 187 1762
rect 215 1758 219 1762
rect 247 1758 251 1762
rect 279 1758 283 1762
rect 311 1758 315 1762
rect 343 1758 347 1762
rect 375 1758 379 1762
rect 407 1758 411 1762
rect 439 1758 443 1762
rect 471 1758 475 1762
rect 503 1758 507 1762
rect 535 1758 539 1762
rect 567 1758 571 1762
rect 599 1758 603 1762
rect 631 1758 635 1762
rect 663 1758 667 1762
rect 695 1758 699 1762
rect 727 1758 731 1762
rect 759 1758 763 1762
rect 791 1758 795 1762
rect 823 1758 827 1762
rect 855 1758 859 1762
rect 887 1758 891 1762
rect 919 1758 923 1762
rect 951 1758 955 1762
rect 983 1758 987 1762
rect 1695 1758 1699 1762
rect 111 1714 115 1718
rect 151 1714 155 1718
rect 183 1714 187 1718
rect 191 1714 195 1718
rect 215 1714 219 1718
rect 247 1714 251 1718
rect 279 1714 283 1718
rect 311 1714 315 1718
rect 319 1714 323 1718
rect 343 1714 347 1718
rect 375 1714 379 1718
rect 407 1714 411 1718
rect 415 1714 419 1718
rect 439 1714 443 1718
rect 471 1714 475 1718
rect 503 1714 507 1718
rect 527 1714 531 1718
rect 535 1714 539 1718
rect 567 1714 571 1718
rect 599 1714 603 1718
rect 631 1714 635 1718
rect 655 1714 659 1718
rect 663 1714 667 1718
rect 695 1714 699 1718
rect 727 1714 731 1718
rect 759 1714 763 1718
rect 791 1714 795 1718
rect 823 1714 827 1718
rect 855 1714 859 1718
rect 887 1714 891 1718
rect 919 1714 923 1718
rect 951 1714 955 1718
rect 983 1714 987 1718
rect 1047 1714 1051 1718
rect 1159 1714 1163 1718
rect 1255 1714 1259 1718
rect 1335 1714 1339 1718
rect 1407 1714 1411 1718
rect 1463 1714 1467 1718
rect 1519 1714 1523 1718
rect 1567 1714 1571 1718
rect 1623 1714 1627 1718
rect 1655 1714 1659 1718
rect 1695 1714 1699 1718
rect 111 1666 115 1670
rect 135 1666 139 1670
rect 175 1666 179 1670
rect 191 1666 195 1670
rect 247 1666 251 1670
rect 263 1666 267 1670
rect 319 1666 323 1670
rect 391 1666 395 1670
rect 415 1666 419 1670
rect 527 1666 531 1670
rect 543 1666 547 1670
rect 655 1666 659 1670
rect 711 1666 715 1670
rect 791 1666 795 1670
rect 879 1666 883 1670
rect 919 1666 923 1670
rect 1039 1666 1043 1670
rect 1047 1666 1051 1670
rect 1159 1666 1163 1670
rect 1183 1666 1187 1670
rect 1255 1666 1259 1670
rect 1319 1666 1323 1670
rect 1335 1666 1339 1670
rect 1407 1666 1411 1670
rect 1439 1666 1443 1670
rect 1463 1666 1467 1670
rect 1519 1666 1523 1670
rect 1559 1666 1563 1670
rect 1567 1666 1571 1670
rect 1623 1666 1627 1670
rect 1655 1666 1659 1670
rect 1695 1666 1699 1670
rect 111 1618 115 1622
rect 135 1618 139 1622
rect 167 1618 171 1622
rect 175 1618 179 1622
rect 199 1618 203 1622
rect 247 1618 251 1622
rect 263 1618 267 1622
rect 327 1618 331 1622
rect 391 1618 395 1622
rect 439 1618 443 1622
rect 543 1618 547 1622
rect 567 1618 571 1622
rect 711 1618 715 1622
rect 855 1618 859 1622
rect 879 1618 883 1622
rect 999 1618 1003 1622
rect 1039 1618 1043 1622
rect 1127 1618 1131 1622
rect 1183 1618 1187 1622
rect 1247 1618 1251 1622
rect 1319 1618 1323 1622
rect 1359 1618 1363 1622
rect 1439 1618 1443 1622
rect 1463 1618 1467 1622
rect 1559 1618 1563 1622
rect 1567 1618 1571 1622
rect 1655 1618 1659 1622
rect 1695 1618 1699 1622
rect 111 1578 115 1582
rect 135 1578 139 1582
rect 167 1578 171 1582
rect 199 1578 203 1582
rect 231 1578 235 1582
rect 247 1578 251 1582
rect 287 1578 291 1582
rect 327 1578 331 1582
rect 343 1578 347 1582
rect 399 1578 403 1582
rect 439 1578 443 1582
rect 455 1578 459 1582
rect 511 1578 515 1582
rect 567 1578 571 1582
rect 575 1578 579 1582
rect 655 1578 659 1582
rect 711 1578 715 1582
rect 751 1578 755 1582
rect 855 1578 859 1582
rect 959 1578 963 1582
rect 999 1578 1003 1582
rect 1063 1578 1067 1582
rect 1127 1578 1131 1582
rect 1159 1578 1163 1582
rect 1247 1578 1251 1582
rect 1327 1578 1331 1582
rect 1359 1578 1363 1582
rect 1399 1578 1403 1582
rect 1463 1578 1467 1582
rect 1471 1578 1475 1582
rect 1535 1578 1539 1582
rect 1567 1578 1571 1582
rect 1607 1578 1611 1582
rect 1655 1578 1659 1582
rect 1695 1578 1699 1582
rect 111 1538 115 1542
rect 135 1538 139 1542
rect 167 1538 171 1542
rect 175 1538 179 1542
rect 223 1538 227 1542
rect 231 1538 235 1542
rect 279 1538 283 1542
rect 287 1538 291 1542
rect 335 1538 339 1542
rect 343 1538 347 1542
rect 399 1538 403 1542
rect 455 1538 459 1542
rect 463 1538 467 1542
rect 511 1538 515 1542
rect 535 1538 539 1542
rect 575 1538 579 1542
rect 607 1538 611 1542
rect 655 1538 659 1542
rect 687 1538 691 1542
rect 751 1538 755 1542
rect 775 1538 779 1542
rect 855 1538 859 1542
rect 871 1538 875 1542
rect 959 1538 963 1542
rect 975 1538 979 1542
rect 1063 1538 1067 1542
rect 1079 1538 1083 1542
rect 1159 1538 1163 1542
rect 1175 1538 1179 1542
rect 1247 1538 1251 1542
rect 1271 1538 1275 1542
rect 1327 1538 1331 1542
rect 1359 1538 1363 1542
rect 1399 1538 1403 1542
rect 1439 1538 1443 1542
rect 1471 1538 1475 1542
rect 1519 1538 1523 1542
rect 1535 1538 1539 1542
rect 1599 1538 1603 1542
rect 1607 1538 1611 1542
rect 1655 1538 1659 1542
rect 1695 1538 1699 1542
rect 111 1494 115 1498
rect 135 1494 139 1498
rect 175 1494 179 1498
rect 207 1494 211 1498
rect 223 1494 227 1498
rect 239 1494 243 1498
rect 271 1494 275 1498
rect 279 1494 283 1498
rect 303 1494 307 1498
rect 335 1494 339 1498
rect 367 1494 371 1498
rect 399 1494 403 1498
rect 431 1494 435 1498
rect 463 1494 467 1498
rect 495 1494 499 1498
rect 527 1494 531 1498
rect 535 1494 539 1498
rect 559 1494 563 1498
rect 591 1494 595 1498
rect 607 1494 611 1498
rect 623 1494 627 1498
rect 663 1494 667 1498
rect 687 1494 691 1498
rect 703 1494 707 1498
rect 743 1494 747 1498
rect 775 1494 779 1498
rect 807 1494 811 1498
rect 871 1494 875 1498
rect 895 1494 899 1498
rect 935 1494 939 1498
rect 975 1494 979 1498
rect 1023 1494 1027 1498
rect 1079 1494 1083 1498
rect 1111 1494 1115 1498
rect 1167 1494 1171 1498
rect 1175 1494 1179 1498
rect 1199 1494 1203 1498
rect 1239 1494 1243 1498
rect 1271 1494 1275 1498
rect 1279 1494 1283 1498
rect 1319 1494 1323 1498
rect 1359 1494 1363 1498
rect 1399 1494 1403 1498
rect 1439 1494 1443 1498
rect 1479 1494 1483 1498
rect 1519 1494 1523 1498
rect 1559 1494 1563 1498
rect 1591 1494 1595 1498
rect 1599 1494 1603 1498
rect 1623 1494 1627 1498
rect 1655 1494 1659 1498
rect 1695 1494 1699 1498
rect 111 1426 115 1430
rect 135 1426 139 1430
rect 167 1426 171 1430
rect 175 1426 179 1430
rect 199 1426 203 1430
rect 207 1426 211 1430
rect 231 1426 235 1430
rect 239 1426 243 1430
rect 263 1426 267 1430
rect 271 1426 275 1430
rect 295 1426 299 1430
rect 303 1426 307 1430
rect 327 1426 331 1430
rect 335 1426 339 1430
rect 359 1426 363 1430
rect 367 1426 371 1430
rect 391 1426 395 1430
rect 399 1426 403 1430
rect 423 1426 427 1430
rect 431 1426 435 1430
rect 455 1426 459 1430
rect 463 1426 467 1430
rect 487 1426 491 1430
rect 495 1426 499 1430
rect 519 1426 523 1430
rect 527 1426 531 1430
rect 551 1426 555 1430
rect 559 1426 563 1430
rect 583 1426 587 1430
rect 591 1426 595 1430
rect 615 1426 619 1430
rect 623 1426 627 1430
rect 647 1426 651 1430
rect 663 1426 667 1430
rect 679 1426 683 1430
rect 703 1426 707 1430
rect 719 1426 723 1430
rect 743 1426 747 1430
rect 767 1426 771 1430
rect 775 1426 779 1430
rect 807 1426 811 1430
rect 839 1426 843 1430
rect 895 1426 899 1430
rect 935 1426 939 1430
rect 975 1426 979 1430
rect 1023 1426 1027 1430
rect 1039 1426 1043 1430
rect 1063 1426 1067 1430
rect 1079 1426 1083 1430
rect 1111 1426 1115 1430
rect 1127 1426 1131 1430
rect 1151 1426 1155 1430
rect 1167 1426 1171 1430
rect 1199 1426 1203 1430
rect 1239 1426 1243 1430
rect 1263 1426 1267 1430
rect 1279 1426 1283 1430
rect 1319 1426 1323 1430
rect 1359 1426 1363 1430
rect 1399 1426 1403 1430
rect 1415 1426 1419 1430
rect 1439 1426 1443 1430
rect 1479 1426 1483 1430
rect 1519 1426 1523 1430
rect 1535 1426 1539 1430
rect 1559 1426 1563 1430
rect 1583 1426 1587 1430
rect 1591 1426 1595 1430
rect 1623 1426 1627 1430
rect 1655 1426 1659 1430
rect 1695 1426 1699 1430
rect 111 1346 115 1350
rect 135 1346 139 1350
rect 167 1346 171 1350
rect 199 1346 203 1350
rect 231 1346 235 1350
rect 263 1346 267 1350
rect 295 1346 299 1350
rect 327 1346 331 1350
rect 359 1346 363 1350
rect 391 1346 395 1350
rect 423 1346 427 1350
rect 455 1346 459 1350
rect 487 1346 491 1350
rect 519 1346 523 1350
rect 551 1346 555 1350
rect 583 1346 587 1350
rect 615 1346 619 1350
rect 647 1346 651 1350
rect 679 1346 683 1350
rect 711 1346 715 1350
rect 735 1346 739 1350
rect 743 1346 747 1350
rect 767 1346 771 1350
rect 807 1346 811 1350
rect 823 1346 827 1350
rect 839 1346 843 1350
rect 887 1346 891 1350
rect 903 1346 907 1350
rect 975 1346 979 1350
rect 983 1346 987 1350
rect 1023 1346 1027 1350
rect 1063 1346 1067 1350
rect 1111 1346 1115 1350
rect 1151 1346 1155 1350
rect 1159 1346 1163 1350
rect 1199 1346 1203 1350
rect 1215 1346 1219 1350
rect 1247 1346 1251 1350
rect 1303 1346 1307 1350
rect 1319 1346 1323 1350
rect 1391 1346 1395 1350
rect 1415 1346 1419 1350
rect 1423 1346 1427 1350
rect 1455 1346 1459 1350
rect 1463 1346 1467 1350
rect 1495 1346 1499 1350
rect 1527 1346 1531 1350
rect 1535 1346 1539 1350
rect 1559 1346 1563 1350
rect 1583 1346 1587 1350
rect 1591 1346 1595 1350
rect 1623 1346 1627 1350
rect 1655 1346 1659 1350
rect 1695 1346 1699 1350
rect 111 1258 115 1262
rect 135 1258 139 1262
rect 167 1258 171 1262
rect 199 1258 203 1262
rect 231 1258 235 1262
rect 263 1258 267 1262
rect 295 1258 299 1262
rect 327 1258 331 1262
rect 359 1258 363 1262
rect 391 1258 395 1262
rect 423 1258 427 1262
rect 455 1258 459 1262
rect 487 1258 491 1262
rect 519 1258 523 1262
rect 551 1258 555 1262
rect 583 1258 587 1262
rect 615 1258 619 1262
rect 647 1258 651 1262
rect 679 1258 683 1262
rect 711 1258 715 1262
rect 743 1258 747 1262
rect 751 1258 755 1262
rect 775 1258 779 1262
rect 811 1258 815 1262
rect 831 1258 835 1262
rect 911 1258 915 1262
rect 959 1258 963 1262
rect 983 1258 987 1262
rect 1015 1258 1019 1262
rect 1023 1258 1027 1262
rect 1063 1258 1067 1262
rect 1087 1258 1091 1262
rect 1127 1258 1131 1262
rect 1159 1258 1163 1262
rect 1175 1258 1179 1262
rect 1215 1258 1219 1262
rect 1255 1258 1259 1262
rect 1295 1258 1299 1262
rect 1303 1258 1307 1262
rect 1343 1258 1347 1262
rect 1375 1258 1379 1262
rect 1391 1258 1395 1262
rect 1407 1258 1411 1262
rect 1423 1258 1427 1262
rect 1439 1258 1443 1262
rect 1455 1258 1459 1262
rect 1479 1258 1483 1262
rect 1495 1258 1499 1262
rect 1519 1258 1523 1262
rect 1527 1258 1531 1262
rect 1559 1258 1563 1262
rect 1591 1258 1595 1262
rect 1623 1258 1627 1262
rect 1655 1258 1659 1262
rect 1695 1258 1699 1262
rect 111 1146 115 1150
rect 135 1146 139 1150
rect 167 1146 171 1150
rect 199 1146 203 1150
rect 231 1146 235 1150
rect 263 1146 267 1150
rect 295 1146 299 1150
rect 327 1146 331 1150
rect 359 1146 363 1150
rect 391 1146 395 1150
rect 423 1146 427 1150
rect 455 1146 459 1150
rect 487 1146 491 1150
rect 519 1146 523 1150
rect 551 1146 555 1150
rect 583 1146 587 1150
rect 615 1146 619 1150
rect 647 1146 651 1150
rect 679 1146 683 1150
rect 687 1146 691 1150
rect 711 1146 715 1150
rect 743 1146 747 1150
rect 775 1146 779 1150
rect 799 1146 803 1150
rect 839 1146 843 1150
rect 847 1146 851 1150
rect 935 1146 939 1150
rect 967 1146 971 1150
rect 975 1146 979 1150
rect 999 1146 1003 1150
rect 1007 1146 1011 1150
rect 1031 1146 1035 1150
rect 1063 1146 1067 1150
rect 1087 1146 1091 1150
rect 1095 1146 1099 1150
rect 1127 1146 1131 1150
rect 1135 1146 1139 1150
rect 1159 1146 1163 1150
rect 1167 1146 1171 1150
rect 1199 1146 1203 1150
rect 1247 1146 1251 1150
rect 1255 1146 1259 1150
rect 1287 1146 1291 1150
rect 1311 1146 1315 1150
rect 1335 1146 1339 1150
rect 1343 1146 1347 1150
rect 1375 1146 1379 1150
rect 1407 1146 1411 1150
rect 1423 1146 1427 1150
rect 1439 1146 1443 1150
rect 1455 1146 1459 1150
rect 1479 1146 1483 1150
rect 1487 1146 1491 1150
rect 1519 1146 1523 1150
rect 1559 1146 1563 1150
rect 1591 1146 1595 1150
rect 1623 1146 1627 1150
rect 1655 1146 1659 1150
rect 1695 1146 1699 1150
rect 111 1030 115 1034
rect 135 1030 139 1034
rect 167 1030 171 1034
rect 199 1030 203 1034
rect 231 1030 235 1034
rect 263 1030 267 1034
rect 295 1030 299 1034
rect 327 1030 331 1034
rect 359 1030 363 1034
rect 391 1030 395 1034
rect 407 1030 411 1034
rect 423 1030 427 1034
rect 455 1030 459 1034
rect 487 1030 491 1034
rect 503 1030 507 1034
rect 519 1030 523 1034
rect 551 1030 555 1034
rect 583 1030 587 1034
rect 591 1030 595 1034
rect 659 1030 663 1034
rect 711 1030 715 1034
rect 799 1030 803 1034
rect 823 1030 827 1034
rect 847 1030 851 1034
rect 919 1030 923 1034
rect 935 1030 939 1034
rect 967 1030 971 1034
rect 975 1030 979 1034
rect 999 1030 1003 1034
rect 1031 1030 1035 1034
rect 1063 1030 1067 1034
rect 1095 1030 1099 1034
rect 1119 1030 1123 1034
rect 1135 1030 1139 1034
rect 1167 1030 1171 1034
rect 1175 1030 1179 1034
rect 1199 1030 1203 1034
rect 1247 1030 1251 1034
rect 1287 1030 1291 1034
rect 1295 1030 1299 1034
rect 1327 1030 1331 1034
rect 1335 1030 1339 1034
rect 1367 1030 1371 1034
rect 1407 1030 1411 1034
rect 1423 1030 1427 1034
rect 1439 1030 1443 1034
rect 1455 1030 1459 1034
rect 1479 1030 1483 1034
rect 1487 1030 1491 1034
rect 1519 1030 1523 1034
rect 1559 1030 1563 1034
rect 1591 1030 1595 1034
rect 1623 1030 1627 1034
rect 1655 1030 1659 1034
rect 1695 1030 1699 1034
rect 111 950 115 954
rect 135 950 139 954
rect 167 950 171 954
rect 199 950 203 954
rect 231 950 235 954
rect 263 950 267 954
rect 279 950 283 954
rect 319 950 323 954
rect 343 950 347 954
rect 399 950 403 954
rect 463 950 467 954
rect 503 950 507 954
rect 583 950 587 954
rect 591 950 595 954
rect 679 950 683 954
rect 711 950 715 954
rect 727 950 731 954
rect 815 950 819 954
rect 863 950 867 954
rect 919 950 923 954
rect 951 950 955 954
rect 967 950 971 954
rect 983 950 987 954
rect 1039 950 1043 954
rect 1063 950 1067 954
rect 1071 950 1075 954
rect 1111 950 1115 954
rect 1135 950 1139 954
rect 1143 950 1147 954
rect 1167 950 1171 954
rect 1199 950 1203 954
rect 1239 950 1243 954
rect 1263 950 1267 954
rect 1271 950 1275 954
rect 1295 950 1299 954
rect 1327 950 1331 954
rect 1367 950 1371 954
rect 1391 950 1395 954
rect 1407 950 1411 954
rect 1423 950 1427 954
rect 1439 950 1443 954
rect 1455 950 1459 954
rect 1479 950 1483 954
rect 1519 950 1523 954
rect 1559 950 1563 954
rect 1591 950 1595 954
rect 1623 950 1627 954
rect 1655 950 1659 954
rect 1695 950 1699 954
rect 111 834 115 838
rect 135 834 139 838
rect 167 834 171 838
rect 207 834 211 838
rect 231 834 235 838
rect 279 834 283 838
rect 327 834 331 838
rect 399 834 403 838
rect 407 834 411 838
rect 435 834 439 838
rect 559 834 563 838
rect 591 834 595 838
rect 663 834 667 838
rect 679 834 683 838
rect 727 834 731 838
rect 815 834 819 838
rect 863 834 867 838
rect 951 834 955 838
rect 999 834 1003 838
rect 1031 834 1035 838
rect 1039 834 1043 838
rect 1071 834 1075 838
rect 1103 834 1107 838
rect 1111 834 1115 838
rect 1143 834 1147 838
rect 1167 834 1171 838
rect 1239 834 1243 838
rect 1247 834 1251 838
rect 1271 834 1275 838
rect 1295 834 1299 838
rect 1327 834 1331 838
rect 1375 834 1379 838
rect 1423 834 1427 838
rect 1471 834 1475 838
rect 1519 834 1523 838
rect 1559 834 1563 838
rect 1591 834 1595 838
rect 1623 834 1627 838
rect 1655 834 1659 838
rect 1695 834 1699 838
rect 111 750 115 754
rect 135 750 139 754
rect 215 750 219 754
rect 231 750 235 754
rect 287 750 291 754
rect 391 750 395 754
rect 407 750 411 754
rect 471 750 475 754
rect 559 750 563 754
rect 615 750 619 754
rect 655 750 659 754
rect 719 750 723 754
rect 767 750 771 754
rect 815 750 819 754
rect 863 750 867 754
rect 911 750 915 754
rect 951 750 955 754
rect 999 750 1003 754
rect 1015 750 1019 754
rect 1087 750 1091 754
rect 1103 750 1107 754
rect 1167 750 1171 754
rect 1183 750 1187 754
rect 1207 750 1211 754
rect 1231 750 1235 754
rect 1247 750 1251 754
rect 1279 750 1283 754
rect 1295 750 1299 754
rect 1311 750 1315 754
rect 1327 750 1331 754
rect 1343 750 1347 754
rect 1375 750 1379 754
rect 1407 750 1411 754
rect 1423 750 1427 754
rect 1439 750 1443 754
rect 1471 750 1475 754
rect 1479 750 1483 754
rect 1519 750 1523 754
rect 1559 750 1563 754
rect 1591 750 1595 754
rect 1623 750 1627 754
rect 1655 750 1659 754
rect 1695 750 1699 754
rect 111 638 115 642
rect 135 638 139 642
rect 143 638 147 642
rect 167 638 171 642
rect 207 638 211 642
rect 215 638 219 642
rect 287 638 291 642
rect 391 638 395 642
rect 407 638 411 642
rect 443 638 447 642
rect 535 638 539 642
rect 615 638 619 642
rect 671 638 675 642
rect 719 638 723 642
rect 767 638 771 642
rect 775 638 779 642
rect 863 638 867 642
rect 903 638 907 642
rect 911 638 915 642
rect 999 638 1003 642
rect 1007 638 1011 642
rect 1095 638 1099 642
rect 1119 638 1123 642
rect 1167 638 1171 642
rect 1207 638 1211 642
rect 1215 638 1219 642
rect 1247 638 1251 642
rect 1279 638 1283 642
rect 1311 638 1315 642
rect 1335 638 1339 642
rect 1343 638 1347 642
rect 1375 638 1379 642
rect 1407 638 1411 642
rect 1415 638 1419 642
rect 1439 638 1443 642
rect 1479 638 1483 642
rect 1519 638 1523 642
rect 1543 638 1547 642
rect 1559 638 1563 642
rect 1591 638 1595 642
rect 1607 638 1611 642
rect 1623 638 1627 642
rect 1655 638 1659 642
rect 1695 638 1699 642
rect 111 558 115 562
rect 135 558 139 562
rect 167 558 171 562
rect 207 558 211 562
rect 247 558 251 562
rect 279 558 283 562
rect 303 558 307 562
rect 391 558 395 562
rect 399 558 403 562
rect 471 558 475 562
rect 535 558 539 562
rect 647 558 651 562
rect 671 558 675 562
rect 727 558 731 562
rect 767 558 771 562
rect 775 558 779 562
rect 871 558 875 562
rect 903 558 907 562
rect 927 558 931 562
rect 991 558 995 562
rect 1031 558 1035 562
rect 1095 558 1099 562
rect 1119 558 1123 562
rect 1199 558 1203 562
rect 1207 558 1211 562
rect 1287 558 1291 562
rect 1335 558 1339 562
rect 1415 558 1419 562
rect 1423 558 1427 562
rect 1479 558 1483 562
rect 1527 558 1531 562
rect 1543 558 1547 562
rect 1575 558 1579 562
rect 1607 558 1611 562
rect 1623 558 1627 562
rect 1655 558 1659 562
rect 1695 558 1699 562
rect 111 438 115 442
rect 135 438 139 442
rect 167 438 171 442
rect 175 438 179 442
rect 199 438 203 442
rect 231 438 235 442
rect 247 438 251 442
rect 263 438 267 442
rect 303 438 307 442
rect 375 438 379 442
rect 399 438 403 442
rect 415 438 419 442
rect 447 438 451 442
rect 471 438 475 442
rect 487 438 491 442
rect 507 438 511 442
rect 543 438 547 442
rect 615 438 619 442
rect 655 438 659 442
rect 671 438 675 442
rect 727 438 731 442
rect 755 438 759 442
rect 783 438 787 442
rect 871 438 875 442
rect 903 438 907 442
rect 935 438 939 442
rect 951 438 955 442
rect 1031 438 1035 442
rect 1075 438 1079 442
rect 1103 438 1107 442
rect 1199 438 1203 442
rect 1231 438 1235 442
rect 1259 438 1263 442
rect 1319 438 1323 442
rect 1359 438 1363 442
rect 1423 438 1427 442
rect 1439 438 1443 442
rect 1479 438 1483 442
rect 1519 438 1523 442
rect 1527 438 1531 442
rect 1559 438 1563 442
rect 1575 438 1579 442
rect 1591 438 1595 442
rect 1623 438 1627 442
rect 1655 438 1659 442
rect 1695 438 1699 442
rect 111 318 115 322
rect 135 318 139 322
rect 167 318 171 322
rect 199 318 203 322
rect 231 318 235 322
rect 263 318 267 322
rect 295 318 299 322
rect 327 318 331 322
rect 359 318 363 322
rect 375 318 379 322
rect 391 318 395 322
rect 415 318 419 322
rect 423 318 427 322
rect 447 318 451 322
rect 455 318 459 322
rect 487 318 491 322
rect 503 318 507 322
rect 519 318 523 322
rect 535 318 539 322
rect 551 318 555 322
rect 599 318 603 322
rect 615 318 619 322
rect 671 318 675 322
rect 703 318 707 322
rect 783 318 787 322
rect 807 318 811 322
rect 903 318 907 322
rect 911 318 915 322
rect 943 318 947 322
rect 999 318 1003 322
rect 1031 318 1035 322
rect 1047 318 1051 322
rect 1063 318 1067 322
rect 1103 318 1107 322
rect 1111 318 1115 322
rect 1199 318 1203 322
rect 1231 318 1235 322
rect 1287 318 1291 322
rect 1319 318 1323 322
rect 1351 318 1355 322
rect 1383 318 1387 322
rect 1415 318 1419 322
rect 1439 318 1443 322
rect 1447 318 1451 322
rect 1479 318 1483 322
rect 1519 318 1523 322
rect 1559 318 1563 322
rect 1591 318 1595 322
rect 1623 318 1627 322
rect 1655 318 1659 322
rect 1695 318 1699 322
rect 111 246 115 250
rect 135 246 139 250
rect 167 246 171 250
rect 183 246 187 250
rect 199 246 203 250
rect 215 246 219 250
rect 231 246 235 250
rect 247 246 251 250
rect 263 246 267 250
rect 279 246 283 250
rect 295 246 299 250
rect 311 246 315 250
rect 327 246 331 250
rect 343 246 347 250
rect 359 246 363 250
rect 375 246 379 250
rect 391 246 395 250
rect 407 246 411 250
rect 423 246 427 250
rect 439 246 443 250
rect 455 246 459 250
rect 471 246 475 250
rect 487 246 491 250
rect 503 246 507 250
rect 519 246 523 250
rect 535 246 539 250
rect 551 246 555 250
rect 567 246 571 250
rect 599 246 603 250
rect 639 246 643 250
rect 695 246 699 250
rect 703 246 707 250
rect 791 246 795 250
rect 807 246 811 250
rect 839 246 843 250
rect 911 246 915 250
rect 919 246 923 250
rect 967 246 971 250
rect 999 246 1003 250
rect 1031 246 1035 250
rect 1063 246 1067 250
rect 1103 246 1107 250
rect 1111 246 1115 250
rect 1143 246 1147 250
rect 1183 246 1187 250
rect 1207 246 1211 250
rect 1223 246 1227 250
rect 1263 246 1267 250
rect 1287 246 1291 250
rect 1303 246 1307 250
rect 1319 246 1323 250
rect 1343 246 1347 250
rect 1351 246 1355 250
rect 1375 246 1379 250
rect 1383 246 1387 250
rect 1407 246 1411 250
rect 1415 246 1419 250
rect 1439 246 1443 250
rect 1447 246 1451 250
rect 1479 246 1483 250
rect 1519 246 1523 250
rect 1559 246 1563 250
rect 1591 246 1595 250
rect 1623 246 1627 250
rect 1655 246 1659 250
rect 1695 246 1699 250
rect 111 170 115 174
rect 135 170 139 174
rect 167 170 171 174
rect 183 170 187 174
rect 215 170 219 174
rect 247 170 251 174
rect 263 170 267 174
rect 279 170 283 174
rect 311 170 315 174
rect 343 170 347 174
rect 367 170 371 174
rect 375 170 379 174
rect 407 170 411 174
rect 415 170 419 174
rect 439 170 443 174
rect 471 170 475 174
rect 503 170 507 174
rect 535 170 539 174
rect 567 170 571 174
rect 599 170 603 174
rect 607 170 611 174
rect 639 170 643 174
rect 687 170 691 174
rect 695 170 699 174
rect 775 170 779 174
rect 791 170 795 174
rect 831 170 835 174
rect 863 170 867 174
rect 919 170 923 174
rect 959 170 963 174
rect 967 170 971 174
rect 1055 170 1059 174
rect 1063 170 1067 174
rect 1103 170 1107 174
rect 1143 170 1147 174
rect 1151 170 1155 174
rect 1183 170 1187 174
rect 1223 170 1227 174
rect 1239 170 1243 174
rect 1263 170 1267 174
rect 1303 170 1307 174
rect 1327 170 1331 174
rect 1343 170 1347 174
rect 1375 170 1379 174
rect 1407 170 1411 174
rect 1415 170 1419 174
rect 1439 170 1443 174
rect 1479 170 1483 174
rect 1503 170 1507 174
rect 1519 170 1523 174
rect 1559 170 1563 174
rect 1591 170 1595 174
rect 1623 170 1627 174
rect 1655 170 1659 174
rect 1695 170 1699 174
rect 111 118 115 122
rect 135 118 139 122
rect 167 118 171 122
rect 199 118 203 122
rect 215 118 219 122
rect 231 118 235 122
rect 263 118 267 122
rect 295 118 299 122
rect 311 118 315 122
rect 327 118 331 122
rect 359 118 363 122
rect 367 118 371 122
rect 391 118 395 122
rect 415 118 419 122
rect 423 118 427 122
rect 455 118 459 122
rect 471 118 475 122
rect 487 118 491 122
rect 519 118 523 122
rect 535 118 539 122
rect 551 118 555 122
rect 607 118 611 122
rect 671 118 675 122
rect 687 118 691 122
rect 743 118 747 122
rect 775 118 779 122
rect 823 118 827 122
rect 863 118 867 122
rect 903 118 907 122
rect 959 118 963 122
rect 983 118 987 122
rect 1055 118 1059 122
rect 1119 118 1123 122
rect 1151 118 1155 122
rect 1175 118 1179 122
rect 1223 118 1227 122
rect 1239 118 1243 122
rect 1271 118 1275 122
rect 1311 118 1315 122
rect 1327 118 1331 122
rect 1343 118 1347 122
rect 1375 118 1379 122
rect 1407 118 1411 122
rect 1415 118 1419 122
rect 1439 118 1443 122
rect 1479 118 1483 122
rect 1503 118 1507 122
rect 1519 118 1523 122
rect 1559 118 1563 122
rect 1591 118 1595 122
rect 1623 118 1627 122
rect 1655 118 1659 122
rect 1695 118 1699 122
rect 111 78 115 82
rect 135 78 139 82
rect 167 78 171 82
rect 199 78 203 82
rect 231 78 235 82
rect 263 78 267 82
rect 295 78 299 82
rect 327 78 331 82
rect 359 78 363 82
rect 391 78 395 82
rect 423 78 427 82
rect 455 78 459 82
rect 487 78 491 82
rect 519 78 523 82
rect 551 78 555 82
rect 607 78 611 82
rect 671 78 675 82
rect 743 78 747 82
rect 823 78 827 82
rect 903 78 907 82
rect 983 78 987 82
rect 1055 78 1059 82
rect 1119 78 1123 82
rect 1175 78 1179 82
rect 1223 78 1227 82
rect 1271 78 1275 82
rect 1311 78 1315 82
rect 1343 78 1347 82
rect 1375 78 1379 82
rect 1407 78 1411 82
rect 1439 78 1443 82
rect 1479 78 1483 82
rect 1519 78 1523 82
rect 1559 78 1563 82
rect 1591 78 1595 82
rect 1623 78 1627 82
rect 1655 78 1659 82
rect 1695 78 1699 82
<< m4 >>
rect 84 1757 85 1763
rect 91 1762 1719 1763
rect 91 1758 111 1762
rect 115 1758 151 1762
rect 155 1758 183 1762
rect 187 1758 215 1762
rect 219 1758 247 1762
rect 251 1758 279 1762
rect 283 1758 311 1762
rect 315 1758 343 1762
rect 347 1758 375 1762
rect 379 1758 407 1762
rect 411 1758 439 1762
rect 443 1758 471 1762
rect 475 1758 503 1762
rect 507 1758 535 1762
rect 539 1758 567 1762
rect 571 1758 599 1762
rect 603 1758 631 1762
rect 635 1758 663 1762
rect 667 1758 695 1762
rect 699 1758 727 1762
rect 731 1758 759 1762
rect 763 1758 791 1762
rect 795 1758 823 1762
rect 827 1758 855 1762
rect 859 1758 887 1762
rect 891 1758 919 1762
rect 923 1758 951 1762
rect 955 1758 983 1762
rect 987 1758 1695 1762
rect 1699 1758 1719 1762
rect 91 1757 1719 1758
rect 1725 1757 1726 1763
rect 96 1713 97 1719
rect 103 1718 1731 1719
rect 103 1714 111 1718
rect 115 1714 151 1718
rect 155 1714 183 1718
rect 187 1714 191 1718
rect 195 1714 215 1718
rect 219 1714 247 1718
rect 251 1714 279 1718
rect 283 1714 311 1718
rect 315 1714 319 1718
rect 323 1714 343 1718
rect 347 1714 375 1718
rect 379 1714 407 1718
rect 411 1714 415 1718
rect 419 1714 439 1718
rect 443 1714 471 1718
rect 475 1714 503 1718
rect 507 1714 527 1718
rect 531 1714 535 1718
rect 539 1714 567 1718
rect 571 1714 599 1718
rect 603 1714 631 1718
rect 635 1714 655 1718
rect 659 1714 663 1718
rect 667 1714 695 1718
rect 699 1714 727 1718
rect 731 1714 759 1718
rect 763 1714 791 1718
rect 795 1714 823 1718
rect 827 1714 855 1718
rect 859 1714 887 1718
rect 891 1714 919 1718
rect 923 1714 951 1718
rect 955 1714 983 1718
rect 987 1714 1047 1718
rect 1051 1714 1159 1718
rect 1163 1714 1255 1718
rect 1259 1714 1335 1718
rect 1339 1714 1407 1718
rect 1411 1714 1463 1718
rect 1467 1714 1519 1718
rect 1523 1714 1567 1718
rect 1571 1714 1623 1718
rect 1627 1714 1655 1718
rect 1659 1714 1695 1718
rect 1699 1714 1731 1718
rect 103 1713 1731 1714
rect 1737 1713 1738 1719
rect 84 1665 85 1671
rect 91 1670 1719 1671
rect 91 1666 111 1670
rect 115 1666 135 1670
rect 139 1666 175 1670
rect 179 1666 191 1670
rect 195 1666 247 1670
rect 251 1666 263 1670
rect 267 1666 319 1670
rect 323 1666 391 1670
rect 395 1666 415 1670
rect 419 1666 527 1670
rect 531 1666 543 1670
rect 547 1666 655 1670
rect 659 1666 711 1670
rect 715 1666 791 1670
rect 795 1666 879 1670
rect 883 1666 919 1670
rect 923 1666 1039 1670
rect 1043 1666 1047 1670
rect 1051 1666 1159 1670
rect 1163 1666 1183 1670
rect 1187 1666 1255 1670
rect 1259 1666 1319 1670
rect 1323 1666 1335 1670
rect 1339 1666 1407 1670
rect 1411 1666 1439 1670
rect 1443 1666 1463 1670
rect 1467 1666 1519 1670
rect 1523 1666 1559 1670
rect 1563 1666 1567 1670
rect 1571 1666 1623 1670
rect 1627 1666 1655 1670
rect 1659 1666 1695 1670
rect 1699 1666 1719 1670
rect 91 1665 1719 1666
rect 1725 1665 1726 1671
rect 96 1617 97 1623
rect 103 1622 1731 1623
rect 103 1618 111 1622
rect 115 1618 135 1622
rect 139 1618 167 1622
rect 171 1618 175 1622
rect 179 1618 199 1622
rect 203 1618 247 1622
rect 251 1618 263 1622
rect 267 1618 327 1622
rect 331 1618 391 1622
rect 395 1618 439 1622
rect 443 1618 543 1622
rect 547 1618 567 1622
rect 571 1618 711 1622
rect 715 1618 855 1622
rect 859 1618 879 1622
rect 883 1618 999 1622
rect 1003 1618 1039 1622
rect 1043 1618 1127 1622
rect 1131 1618 1183 1622
rect 1187 1618 1247 1622
rect 1251 1618 1319 1622
rect 1323 1618 1359 1622
rect 1363 1618 1439 1622
rect 1443 1618 1463 1622
rect 1467 1618 1559 1622
rect 1563 1618 1567 1622
rect 1571 1618 1655 1622
rect 1659 1618 1695 1622
rect 1699 1618 1731 1622
rect 103 1617 1731 1618
rect 1737 1617 1738 1623
rect 84 1577 85 1583
rect 91 1582 1719 1583
rect 91 1578 111 1582
rect 115 1578 135 1582
rect 139 1578 167 1582
rect 171 1578 199 1582
rect 203 1578 231 1582
rect 235 1578 247 1582
rect 251 1578 287 1582
rect 291 1578 327 1582
rect 331 1578 343 1582
rect 347 1578 399 1582
rect 403 1578 439 1582
rect 443 1578 455 1582
rect 459 1578 511 1582
rect 515 1578 567 1582
rect 571 1578 575 1582
rect 579 1578 655 1582
rect 659 1578 711 1582
rect 715 1578 751 1582
rect 755 1578 855 1582
rect 859 1578 959 1582
rect 963 1578 999 1582
rect 1003 1578 1063 1582
rect 1067 1578 1127 1582
rect 1131 1578 1159 1582
rect 1163 1578 1247 1582
rect 1251 1578 1327 1582
rect 1331 1578 1359 1582
rect 1363 1578 1399 1582
rect 1403 1578 1463 1582
rect 1467 1578 1471 1582
rect 1475 1578 1535 1582
rect 1539 1578 1567 1582
rect 1571 1578 1607 1582
rect 1611 1578 1655 1582
rect 1659 1578 1695 1582
rect 1699 1578 1719 1582
rect 91 1577 1719 1578
rect 1725 1577 1726 1583
rect 96 1537 97 1543
rect 103 1542 1731 1543
rect 103 1538 111 1542
rect 115 1538 135 1542
rect 139 1538 167 1542
rect 171 1538 175 1542
rect 179 1538 223 1542
rect 227 1538 231 1542
rect 235 1538 279 1542
rect 283 1538 287 1542
rect 291 1538 335 1542
rect 339 1538 343 1542
rect 347 1538 399 1542
rect 403 1538 455 1542
rect 459 1538 463 1542
rect 467 1538 511 1542
rect 515 1538 535 1542
rect 539 1538 575 1542
rect 579 1538 607 1542
rect 611 1538 655 1542
rect 659 1538 687 1542
rect 691 1538 751 1542
rect 755 1538 775 1542
rect 779 1538 855 1542
rect 859 1538 871 1542
rect 875 1538 959 1542
rect 963 1538 975 1542
rect 979 1538 1063 1542
rect 1067 1538 1079 1542
rect 1083 1538 1159 1542
rect 1163 1538 1175 1542
rect 1179 1538 1247 1542
rect 1251 1538 1271 1542
rect 1275 1538 1327 1542
rect 1331 1538 1359 1542
rect 1363 1538 1399 1542
rect 1403 1538 1439 1542
rect 1443 1538 1471 1542
rect 1475 1538 1519 1542
rect 1523 1538 1535 1542
rect 1539 1538 1599 1542
rect 1603 1538 1607 1542
rect 1611 1538 1655 1542
rect 1659 1538 1695 1542
rect 1699 1538 1731 1542
rect 103 1537 1731 1538
rect 1737 1537 1738 1543
rect 84 1493 85 1499
rect 91 1498 1719 1499
rect 91 1494 111 1498
rect 115 1494 135 1498
rect 139 1494 175 1498
rect 179 1494 207 1498
rect 211 1494 223 1498
rect 227 1494 239 1498
rect 243 1494 271 1498
rect 275 1494 279 1498
rect 283 1494 303 1498
rect 307 1494 335 1498
rect 339 1494 367 1498
rect 371 1494 399 1498
rect 403 1494 431 1498
rect 435 1494 463 1498
rect 467 1494 495 1498
rect 499 1494 527 1498
rect 531 1494 535 1498
rect 539 1494 559 1498
rect 563 1494 591 1498
rect 595 1494 607 1498
rect 611 1494 623 1498
rect 627 1494 663 1498
rect 667 1494 687 1498
rect 691 1494 703 1498
rect 707 1494 743 1498
rect 747 1494 775 1498
rect 779 1494 807 1498
rect 811 1494 871 1498
rect 875 1494 895 1498
rect 899 1494 935 1498
rect 939 1494 975 1498
rect 979 1494 1023 1498
rect 1027 1494 1079 1498
rect 1083 1494 1111 1498
rect 1115 1494 1167 1498
rect 1171 1494 1175 1498
rect 1179 1494 1199 1498
rect 1203 1494 1239 1498
rect 1243 1494 1271 1498
rect 1275 1494 1279 1498
rect 1283 1494 1319 1498
rect 1323 1494 1359 1498
rect 1363 1494 1399 1498
rect 1403 1494 1439 1498
rect 1443 1494 1479 1498
rect 1483 1494 1519 1498
rect 1523 1494 1559 1498
rect 1563 1494 1591 1498
rect 1595 1494 1599 1498
rect 1603 1494 1623 1498
rect 1627 1494 1655 1498
rect 1659 1494 1695 1498
rect 1699 1494 1719 1498
rect 91 1493 1719 1494
rect 1725 1493 1726 1499
rect 96 1425 97 1431
rect 103 1430 1731 1431
rect 103 1426 111 1430
rect 115 1426 135 1430
rect 139 1426 167 1430
rect 171 1426 175 1430
rect 179 1426 199 1430
rect 203 1426 207 1430
rect 211 1426 231 1430
rect 235 1426 239 1430
rect 243 1426 263 1430
rect 267 1426 271 1430
rect 275 1426 295 1430
rect 299 1426 303 1430
rect 307 1426 327 1430
rect 331 1426 335 1430
rect 339 1426 359 1430
rect 363 1426 367 1430
rect 371 1426 391 1430
rect 395 1426 399 1430
rect 403 1426 423 1430
rect 427 1426 431 1430
rect 435 1426 455 1430
rect 459 1426 463 1430
rect 467 1426 487 1430
rect 491 1426 495 1430
rect 499 1426 519 1430
rect 523 1426 527 1430
rect 531 1426 551 1430
rect 555 1426 559 1430
rect 563 1426 583 1430
rect 587 1426 591 1430
rect 595 1426 615 1430
rect 619 1426 623 1430
rect 627 1426 647 1430
rect 651 1426 663 1430
rect 667 1426 679 1430
rect 683 1426 703 1430
rect 707 1426 719 1430
rect 723 1426 743 1430
rect 747 1426 767 1430
rect 771 1426 775 1430
rect 779 1426 807 1430
rect 811 1426 839 1430
rect 843 1426 895 1430
rect 899 1426 935 1430
rect 939 1426 975 1430
rect 979 1426 1023 1430
rect 1027 1426 1039 1430
rect 1043 1426 1063 1430
rect 1067 1426 1079 1430
rect 1083 1426 1111 1430
rect 1115 1426 1127 1430
rect 1131 1426 1151 1430
rect 1155 1426 1167 1430
rect 1171 1426 1199 1430
rect 1203 1426 1239 1430
rect 1243 1426 1263 1430
rect 1267 1426 1279 1430
rect 1283 1426 1319 1430
rect 1323 1426 1359 1430
rect 1363 1426 1399 1430
rect 1403 1426 1415 1430
rect 1419 1426 1439 1430
rect 1443 1426 1479 1430
rect 1483 1426 1519 1430
rect 1523 1426 1535 1430
rect 1539 1426 1559 1430
rect 1563 1426 1583 1430
rect 1587 1426 1591 1430
rect 1595 1426 1623 1430
rect 1627 1426 1655 1430
rect 1659 1426 1695 1430
rect 1699 1426 1731 1430
rect 103 1425 1731 1426
rect 1737 1425 1738 1431
rect 84 1345 85 1351
rect 91 1350 1719 1351
rect 91 1346 111 1350
rect 115 1346 135 1350
rect 139 1346 167 1350
rect 171 1346 199 1350
rect 203 1346 231 1350
rect 235 1346 263 1350
rect 267 1346 295 1350
rect 299 1346 327 1350
rect 331 1346 359 1350
rect 363 1346 391 1350
rect 395 1346 423 1350
rect 427 1346 455 1350
rect 459 1346 487 1350
rect 491 1346 519 1350
rect 523 1346 551 1350
rect 555 1346 583 1350
rect 587 1346 615 1350
rect 619 1346 647 1350
rect 651 1346 679 1350
rect 683 1346 711 1350
rect 715 1346 735 1350
rect 739 1346 743 1350
rect 747 1346 767 1350
rect 771 1346 807 1350
rect 811 1346 823 1350
rect 827 1346 839 1350
rect 843 1346 887 1350
rect 891 1346 903 1350
rect 907 1346 975 1350
rect 979 1346 983 1350
rect 987 1346 1023 1350
rect 1027 1346 1063 1350
rect 1067 1346 1111 1350
rect 1115 1346 1151 1350
rect 1155 1346 1159 1350
rect 1163 1346 1199 1350
rect 1203 1346 1215 1350
rect 1219 1346 1247 1350
rect 1251 1346 1303 1350
rect 1307 1346 1319 1350
rect 1323 1346 1391 1350
rect 1395 1346 1415 1350
rect 1419 1346 1423 1350
rect 1427 1346 1455 1350
rect 1459 1346 1463 1350
rect 1467 1346 1495 1350
rect 1499 1346 1527 1350
rect 1531 1346 1535 1350
rect 1539 1346 1559 1350
rect 1563 1346 1583 1350
rect 1587 1346 1591 1350
rect 1595 1346 1623 1350
rect 1627 1346 1655 1350
rect 1659 1346 1695 1350
rect 1699 1346 1719 1350
rect 91 1345 1719 1346
rect 1725 1345 1726 1351
rect 96 1257 97 1263
rect 103 1262 1731 1263
rect 103 1258 111 1262
rect 115 1258 135 1262
rect 139 1258 167 1262
rect 171 1258 199 1262
rect 203 1258 231 1262
rect 235 1258 263 1262
rect 267 1258 295 1262
rect 299 1258 327 1262
rect 331 1258 359 1262
rect 363 1258 391 1262
rect 395 1258 423 1262
rect 427 1258 455 1262
rect 459 1258 487 1262
rect 491 1258 519 1262
rect 523 1258 551 1262
rect 555 1258 583 1262
rect 587 1258 615 1262
rect 619 1258 647 1262
rect 651 1258 679 1262
rect 683 1258 711 1262
rect 715 1258 743 1262
rect 747 1258 751 1262
rect 755 1258 775 1262
rect 779 1258 811 1262
rect 815 1258 831 1262
rect 835 1258 911 1262
rect 915 1258 959 1262
rect 963 1258 983 1262
rect 987 1258 1015 1262
rect 1019 1258 1023 1262
rect 1027 1258 1063 1262
rect 1067 1258 1087 1262
rect 1091 1258 1127 1262
rect 1131 1258 1159 1262
rect 1163 1258 1175 1262
rect 1179 1258 1215 1262
rect 1219 1258 1255 1262
rect 1259 1258 1295 1262
rect 1299 1258 1303 1262
rect 1307 1258 1343 1262
rect 1347 1258 1375 1262
rect 1379 1258 1391 1262
rect 1395 1258 1407 1262
rect 1411 1258 1423 1262
rect 1427 1258 1439 1262
rect 1443 1258 1455 1262
rect 1459 1258 1479 1262
rect 1483 1258 1495 1262
rect 1499 1258 1519 1262
rect 1523 1258 1527 1262
rect 1531 1258 1559 1262
rect 1563 1258 1591 1262
rect 1595 1258 1623 1262
rect 1627 1258 1655 1262
rect 1659 1258 1695 1262
rect 1699 1258 1731 1262
rect 103 1257 1731 1258
rect 1737 1257 1738 1263
rect 84 1145 85 1151
rect 91 1150 1719 1151
rect 91 1146 111 1150
rect 115 1146 135 1150
rect 139 1146 167 1150
rect 171 1146 199 1150
rect 203 1146 231 1150
rect 235 1146 263 1150
rect 267 1146 295 1150
rect 299 1146 327 1150
rect 331 1146 359 1150
rect 363 1146 391 1150
rect 395 1146 423 1150
rect 427 1146 455 1150
rect 459 1146 487 1150
rect 491 1146 519 1150
rect 523 1146 551 1150
rect 555 1146 583 1150
rect 587 1146 615 1150
rect 619 1146 647 1150
rect 651 1146 679 1150
rect 683 1146 687 1150
rect 691 1146 711 1150
rect 715 1146 743 1150
rect 747 1146 775 1150
rect 779 1146 799 1150
rect 803 1146 839 1150
rect 843 1146 847 1150
rect 851 1146 935 1150
rect 939 1146 967 1150
rect 971 1146 975 1150
rect 979 1146 999 1150
rect 1003 1146 1007 1150
rect 1011 1146 1031 1150
rect 1035 1146 1063 1150
rect 1067 1146 1087 1150
rect 1091 1146 1095 1150
rect 1099 1146 1127 1150
rect 1131 1146 1135 1150
rect 1139 1146 1159 1150
rect 1163 1146 1167 1150
rect 1171 1146 1199 1150
rect 1203 1146 1247 1150
rect 1251 1146 1255 1150
rect 1259 1146 1287 1150
rect 1291 1146 1311 1150
rect 1315 1146 1335 1150
rect 1339 1146 1343 1150
rect 1347 1146 1375 1150
rect 1379 1146 1407 1150
rect 1411 1146 1423 1150
rect 1427 1146 1439 1150
rect 1443 1146 1455 1150
rect 1459 1146 1479 1150
rect 1483 1146 1487 1150
rect 1491 1146 1519 1150
rect 1523 1146 1559 1150
rect 1563 1146 1591 1150
rect 1595 1146 1623 1150
rect 1627 1146 1655 1150
rect 1659 1146 1695 1150
rect 1699 1146 1719 1150
rect 91 1145 1719 1146
rect 1725 1145 1726 1151
rect 96 1029 97 1035
rect 103 1034 1731 1035
rect 103 1030 111 1034
rect 115 1030 135 1034
rect 139 1030 167 1034
rect 171 1030 199 1034
rect 203 1030 231 1034
rect 235 1030 263 1034
rect 267 1030 295 1034
rect 299 1030 327 1034
rect 331 1030 359 1034
rect 363 1030 391 1034
rect 395 1030 407 1034
rect 411 1030 423 1034
rect 427 1030 455 1034
rect 459 1030 487 1034
rect 491 1030 503 1034
rect 507 1030 519 1034
rect 523 1030 551 1034
rect 555 1030 583 1034
rect 587 1030 591 1034
rect 595 1030 659 1034
rect 663 1030 711 1034
rect 715 1030 799 1034
rect 803 1030 823 1034
rect 827 1030 847 1034
rect 851 1030 919 1034
rect 923 1030 935 1034
rect 939 1030 967 1034
rect 971 1030 975 1034
rect 979 1030 999 1034
rect 1003 1030 1031 1034
rect 1035 1030 1063 1034
rect 1067 1030 1095 1034
rect 1099 1030 1119 1034
rect 1123 1030 1135 1034
rect 1139 1030 1167 1034
rect 1171 1030 1175 1034
rect 1179 1030 1199 1034
rect 1203 1030 1247 1034
rect 1251 1030 1287 1034
rect 1291 1030 1295 1034
rect 1299 1030 1327 1034
rect 1331 1030 1335 1034
rect 1339 1030 1367 1034
rect 1371 1030 1407 1034
rect 1411 1030 1423 1034
rect 1427 1030 1439 1034
rect 1443 1030 1455 1034
rect 1459 1030 1479 1034
rect 1483 1030 1487 1034
rect 1491 1030 1519 1034
rect 1523 1030 1559 1034
rect 1563 1030 1591 1034
rect 1595 1030 1623 1034
rect 1627 1030 1655 1034
rect 1659 1030 1695 1034
rect 1699 1030 1731 1034
rect 103 1029 1731 1030
rect 1737 1029 1738 1035
rect 84 949 85 955
rect 91 954 1719 955
rect 91 950 111 954
rect 115 950 135 954
rect 139 950 167 954
rect 171 950 199 954
rect 203 950 231 954
rect 235 950 263 954
rect 267 950 279 954
rect 283 950 319 954
rect 323 950 343 954
rect 347 950 399 954
rect 403 950 463 954
rect 467 950 503 954
rect 507 950 583 954
rect 587 950 591 954
rect 595 950 679 954
rect 683 950 711 954
rect 715 950 727 954
rect 731 950 815 954
rect 819 950 863 954
rect 867 950 919 954
rect 923 950 951 954
rect 955 950 967 954
rect 971 950 983 954
rect 987 950 1039 954
rect 1043 950 1063 954
rect 1067 950 1071 954
rect 1075 950 1111 954
rect 1115 950 1135 954
rect 1139 950 1143 954
rect 1147 950 1167 954
rect 1171 950 1199 954
rect 1203 950 1239 954
rect 1243 950 1263 954
rect 1267 950 1271 954
rect 1275 950 1295 954
rect 1299 950 1327 954
rect 1331 950 1367 954
rect 1371 950 1391 954
rect 1395 950 1407 954
rect 1411 950 1423 954
rect 1427 950 1439 954
rect 1443 950 1455 954
rect 1459 950 1479 954
rect 1483 950 1519 954
rect 1523 950 1559 954
rect 1563 950 1591 954
rect 1595 950 1623 954
rect 1627 950 1655 954
rect 1659 950 1695 954
rect 1699 950 1719 954
rect 91 949 1719 950
rect 1725 949 1726 955
rect 96 833 97 839
rect 103 838 1731 839
rect 103 834 111 838
rect 115 834 135 838
rect 139 834 167 838
rect 171 834 207 838
rect 211 834 231 838
rect 235 834 279 838
rect 283 834 327 838
rect 331 834 399 838
rect 403 834 407 838
rect 411 834 435 838
rect 439 834 559 838
rect 563 834 591 838
rect 595 834 663 838
rect 667 834 679 838
rect 683 834 727 838
rect 731 834 815 838
rect 819 834 863 838
rect 867 834 951 838
rect 955 834 999 838
rect 1003 834 1031 838
rect 1035 834 1039 838
rect 1043 834 1071 838
rect 1075 834 1103 838
rect 1107 834 1111 838
rect 1115 834 1143 838
rect 1147 834 1167 838
rect 1171 834 1239 838
rect 1243 834 1247 838
rect 1251 834 1271 838
rect 1275 834 1295 838
rect 1299 834 1327 838
rect 1331 834 1375 838
rect 1379 834 1423 838
rect 1427 834 1471 838
rect 1475 834 1519 838
rect 1523 834 1559 838
rect 1563 834 1591 838
rect 1595 834 1623 838
rect 1627 834 1655 838
rect 1659 834 1695 838
rect 1699 834 1731 838
rect 103 833 1731 834
rect 1737 833 1738 839
rect 84 749 85 755
rect 91 754 1719 755
rect 91 750 111 754
rect 115 750 135 754
rect 139 750 215 754
rect 219 750 231 754
rect 235 750 287 754
rect 291 750 391 754
rect 395 750 407 754
rect 411 750 471 754
rect 475 750 559 754
rect 563 750 615 754
rect 619 750 655 754
rect 659 750 719 754
rect 723 750 767 754
rect 771 750 815 754
rect 819 750 863 754
rect 867 750 911 754
rect 915 750 951 754
rect 955 750 999 754
rect 1003 750 1015 754
rect 1019 750 1087 754
rect 1091 750 1103 754
rect 1107 750 1167 754
rect 1171 750 1183 754
rect 1187 750 1207 754
rect 1211 750 1231 754
rect 1235 750 1247 754
rect 1251 750 1279 754
rect 1283 750 1295 754
rect 1299 750 1311 754
rect 1315 750 1327 754
rect 1331 750 1343 754
rect 1347 750 1375 754
rect 1379 750 1407 754
rect 1411 750 1423 754
rect 1427 750 1439 754
rect 1443 750 1471 754
rect 1475 750 1479 754
rect 1483 750 1519 754
rect 1523 750 1559 754
rect 1563 750 1591 754
rect 1595 750 1623 754
rect 1627 750 1655 754
rect 1659 750 1695 754
rect 1699 750 1719 754
rect 91 749 1719 750
rect 1725 749 1726 755
rect 96 637 97 643
rect 103 642 1731 643
rect 103 638 111 642
rect 115 638 135 642
rect 139 638 143 642
rect 147 638 167 642
rect 171 638 207 642
rect 211 638 215 642
rect 219 638 287 642
rect 291 638 391 642
rect 395 638 407 642
rect 411 638 443 642
rect 447 638 535 642
rect 539 638 615 642
rect 619 638 671 642
rect 675 638 719 642
rect 723 638 767 642
rect 771 638 775 642
rect 779 638 863 642
rect 867 638 903 642
rect 907 638 911 642
rect 915 638 999 642
rect 1003 638 1007 642
rect 1011 638 1095 642
rect 1099 638 1119 642
rect 1123 638 1167 642
rect 1171 638 1207 642
rect 1211 638 1215 642
rect 1219 638 1247 642
rect 1251 638 1279 642
rect 1283 638 1311 642
rect 1315 638 1335 642
rect 1339 638 1343 642
rect 1347 638 1375 642
rect 1379 638 1407 642
rect 1411 638 1415 642
rect 1419 638 1439 642
rect 1443 638 1479 642
rect 1483 638 1519 642
rect 1523 638 1543 642
rect 1547 638 1559 642
rect 1563 638 1591 642
rect 1595 638 1607 642
rect 1611 638 1623 642
rect 1627 638 1655 642
rect 1659 638 1695 642
rect 1699 638 1731 642
rect 103 637 1731 638
rect 1737 637 1738 643
rect 84 557 85 563
rect 91 562 1719 563
rect 91 558 111 562
rect 115 558 135 562
rect 139 558 167 562
rect 171 558 207 562
rect 211 558 247 562
rect 251 558 279 562
rect 283 558 303 562
rect 307 558 391 562
rect 395 558 399 562
rect 403 558 471 562
rect 475 558 535 562
rect 539 558 647 562
rect 651 558 671 562
rect 675 558 727 562
rect 731 558 767 562
rect 771 558 775 562
rect 779 558 871 562
rect 875 558 903 562
rect 907 558 927 562
rect 931 558 991 562
rect 995 558 1031 562
rect 1035 558 1095 562
rect 1099 558 1119 562
rect 1123 558 1199 562
rect 1203 558 1207 562
rect 1211 558 1287 562
rect 1291 558 1335 562
rect 1339 558 1415 562
rect 1419 558 1423 562
rect 1427 558 1479 562
rect 1483 558 1527 562
rect 1531 558 1543 562
rect 1547 558 1575 562
rect 1579 558 1607 562
rect 1611 558 1623 562
rect 1627 558 1655 562
rect 1659 558 1695 562
rect 1699 558 1719 562
rect 91 557 1719 558
rect 1725 557 1726 563
rect 96 437 97 443
rect 103 442 1731 443
rect 103 438 111 442
rect 115 438 135 442
rect 139 438 167 442
rect 171 438 175 442
rect 179 438 199 442
rect 203 438 231 442
rect 235 438 247 442
rect 251 438 263 442
rect 267 438 303 442
rect 307 438 375 442
rect 379 438 399 442
rect 403 438 415 442
rect 419 438 447 442
rect 451 438 471 442
rect 475 438 487 442
rect 491 438 507 442
rect 511 438 543 442
rect 547 438 615 442
rect 619 438 655 442
rect 659 438 671 442
rect 675 438 727 442
rect 731 438 755 442
rect 759 438 783 442
rect 787 438 871 442
rect 875 438 903 442
rect 907 438 935 442
rect 939 438 951 442
rect 955 438 1031 442
rect 1035 438 1075 442
rect 1079 438 1103 442
rect 1107 438 1199 442
rect 1203 438 1231 442
rect 1235 438 1259 442
rect 1263 438 1319 442
rect 1323 438 1359 442
rect 1363 438 1423 442
rect 1427 438 1439 442
rect 1443 438 1479 442
rect 1483 438 1519 442
rect 1523 438 1527 442
rect 1531 438 1559 442
rect 1563 438 1575 442
rect 1579 438 1591 442
rect 1595 438 1623 442
rect 1627 438 1655 442
rect 1659 438 1695 442
rect 1699 438 1731 442
rect 103 437 1731 438
rect 1737 437 1738 443
rect 84 317 85 323
rect 91 322 1719 323
rect 91 318 111 322
rect 115 318 135 322
rect 139 318 167 322
rect 171 318 199 322
rect 203 318 231 322
rect 235 318 263 322
rect 267 318 295 322
rect 299 318 327 322
rect 331 318 359 322
rect 363 318 375 322
rect 379 318 391 322
rect 395 318 415 322
rect 419 318 423 322
rect 427 318 447 322
rect 451 318 455 322
rect 459 318 487 322
rect 491 318 503 322
rect 507 318 519 322
rect 523 318 535 322
rect 539 318 551 322
rect 555 318 599 322
rect 603 318 615 322
rect 619 318 671 322
rect 675 318 703 322
rect 707 318 783 322
rect 787 318 807 322
rect 811 318 903 322
rect 907 318 911 322
rect 915 318 943 322
rect 947 318 999 322
rect 1003 318 1031 322
rect 1035 318 1047 322
rect 1051 318 1063 322
rect 1067 318 1103 322
rect 1107 318 1111 322
rect 1115 318 1199 322
rect 1203 318 1231 322
rect 1235 318 1287 322
rect 1291 318 1319 322
rect 1323 318 1351 322
rect 1355 318 1383 322
rect 1387 318 1415 322
rect 1419 318 1439 322
rect 1443 318 1447 322
rect 1451 318 1479 322
rect 1483 318 1519 322
rect 1523 318 1559 322
rect 1563 318 1591 322
rect 1595 318 1623 322
rect 1627 318 1655 322
rect 1659 318 1695 322
rect 1699 318 1719 322
rect 91 317 1719 318
rect 1725 317 1726 323
rect 96 245 97 251
rect 103 250 1731 251
rect 103 246 111 250
rect 115 246 135 250
rect 139 246 167 250
rect 171 246 183 250
rect 187 246 199 250
rect 203 246 215 250
rect 219 246 231 250
rect 235 246 247 250
rect 251 246 263 250
rect 267 246 279 250
rect 283 246 295 250
rect 299 246 311 250
rect 315 246 327 250
rect 331 246 343 250
rect 347 246 359 250
rect 363 246 375 250
rect 379 246 391 250
rect 395 246 407 250
rect 411 246 423 250
rect 427 246 439 250
rect 443 246 455 250
rect 459 246 471 250
rect 475 246 487 250
rect 491 246 503 250
rect 507 246 519 250
rect 523 246 535 250
rect 539 246 551 250
rect 555 246 567 250
rect 571 246 599 250
rect 603 246 639 250
rect 643 246 695 250
rect 699 246 703 250
rect 707 246 791 250
rect 795 246 807 250
rect 811 246 839 250
rect 843 246 911 250
rect 915 246 919 250
rect 923 246 967 250
rect 971 246 999 250
rect 1003 246 1031 250
rect 1035 246 1063 250
rect 1067 246 1103 250
rect 1107 246 1111 250
rect 1115 246 1143 250
rect 1147 246 1183 250
rect 1187 246 1207 250
rect 1211 246 1223 250
rect 1227 246 1263 250
rect 1267 246 1287 250
rect 1291 246 1303 250
rect 1307 246 1319 250
rect 1323 246 1343 250
rect 1347 246 1351 250
rect 1355 246 1375 250
rect 1379 246 1383 250
rect 1387 246 1407 250
rect 1411 246 1415 250
rect 1419 246 1439 250
rect 1443 246 1447 250
rect 1451 246 1479 250
rect 1483 246 1519 250
rect 1523 246 1559 250
rect 1563 246 1591 250
rect 1595 246 1623 250
rect 1627 246 1655 250
rect 1659 246 1695 250
rect 1699 246 1731 250
rect 103 245 1731 246
rect 1737 245 1738 251
rect 84 169 85 175
rect 91 174 1719 175
rect 91 170 111 174
rect 115 170 135 174
rect 139 170 167 174
rect 171 170 183 174
rect 187 170 215 174
rect 219 170 247 174
rect 251 170 263 174
rect 267 170 279 174
rect 283 170 311 174
rect 315 170 343 174
rect 347 170 367 174
rect 371 170 375 174
rect 379 170 407 174
rect 411 170 415 174
rect 419 170 439 174
rect 443 170 471 174
rect 475 170 503 174
rect 507 170 535 174
rect 539 170 567 174
rect 571 170 599 174
rect 603 170 607 174
rect 611 170 639 174
rect 643 170 687 174
rect 691 170 695 174
rect 699 170 775 174
rect 779 170 791 174
rect 795 170 831 174
rect 835 170 863 174
rect 867 170 919 174
rect 923 170 959 174
rect 963 170 967 174
rect 971 170 1055 174
rect 1059 170 1063 174
rect 1067 170 1103 174
rect 1107 170 1143 174
rect 1147 170 1151 174
rect 1155 170 1183 174
rect 1187 170 1223 174
rect 1227 170 1239 174
rect 1243 170 1263 174
rect 1267 170 1303 174
rect 1307 170 1327 174
rect 1331 170 1343 174
rect 1347 170 1375 174
rect 1379 170 1407 174
rect 1411 170 1415 174
rect 1419 170 1439 174
rect 1443 170 1479 174
rect 1483 170 1503 174
rect 1507 170 1519 174
rect 1523 170 1559 174
rect 1563 170 1591 174
rect 1595 170 1623 174
rect 1627 170 1655 174
rect 1659 170 1695 174
rect 1699 170 1719 174
rect 91 169 1719 170
rect 1725 169 1726 175
rect 96 117 97 123
rect 103 122 1731 123
rect 103 118 111 122
rect 115 118 135 122
rect 139 118 167 122
rect 171 118 199 122
rect 203 118 215 122
rect 219 118 231 122
rect 235 118 263 122
rect 267 118 295 122
rect 299 118 311 122
rect 315 118 327 122
rect 331 118 359 122
rect 363 118 367 122
rect 371 118 391 122
rect 395 118 415 122
rect 419 118 423 122
rect 427 118 455 122
rect 459 118 471 122
rect 475 118 487 122
rect 491 118 519 122
rect 523 118 535 122
rect 539 118 551 122
rect 555 118 607 122
rect 611 118 671 122
rect 675 118 687 122
rect 691 118 743 122
rect 747 118 775 122
rect 779 118 823 122
rect 827 118 863 122
rect 867 118 903 122
rect 907 118 959 122
rect 963 118 983 122
rect 987 118 1055 122
rect 1059 118 1119 122
rect 1123 118 1151 122
rect 1155 118 1175 122
rect 1179 118 1223 122
rect 1227 118 1239 122
rect 1243 118 1271 122
rect 1275 118 1311 122
rect 1315 118 1327 122
rect 1331 118 1343 122
rect 1347 118 1375 122
rect 1379 118 1407 122
rect 1411 118 1415 122
rect 1419 118 1439 122
rect 1443 118 1479 122
rect 1483 118 1503 122
rect 1507 118 1519 122
rect 1523 118 1559 122
rect 1563 118 1591 122
rect 1595 118 1623 122
rect 1627 118 1655 122
rect 1659 118 1695 122
rect 1699 118 1731 122
rect 103 117 1731 118
rect 1737 117 1738 123
rect 84 77 85 83
rect 91 82 1719 83
rect 91 78 111 82
rect 115 78 135 82
rect 139 78 167 82
rect 171 78 199 82
rect 203 78 231 82
rect 235 78 263 82
rect 267 78 295 82
rect 299 78 327 82
rect 331 78 359 82
rect 363 78 391 82
rect 395 78 423 82
rect 427 78 455 82
rect 459 78 487 82
rect 491 78 519 82
rect 523 78 551 82
rect 555 78 607 82
rect 611 78 671 82
rect 675 78 743 82
rect 747 78 823 82
rect 827 78 903 82
rect 907 78 983 82
rect 987 78 1055 82
rect 1059 78 1119 82
rect 1123 78 1175 82
rect 1179 78 1223 82
rect 1227 78 1271 82
rect 1275 78 1311 82
rect 1315 78 1343 82
rect 1347 78 1375 82
rect 1379 78 1407 82
rect 1411 78 1439 82
rect 1443 78 1479 82
rect 1483 78 1519 82
rect 1523 78 1559 82
rect 1563 78 1591 82
rect 1595 78 1623 82
rect 1627 78 1655 82
rect 1659 78 1695 82
rect 1699 78 1719 82
rect 91 77 1719 78
rect 1725 77 1726 83
<< m5c >>
rect 85 1757 91 1763
rect 1719 1757 1725 1763
rect 97 1713 103 1719
rect 1731 1713 1737 1719
rect 85 1665 91 1671
rect 1719 1665 1725 1671
rect 97 1617 103 1623
rect 1731 1617 1737 1623
rect 85 1577 91 1583
rect 1719 1577 1725 1583
rect 97 1537 103 1543
rect 1731 1537 1737 1543
rect 85 1493 91 1499
rect 1719 1493 1725 1499
rect 97 1425 103 1431
rect 1731 1425 1737 1431
rect 85 1345 91 1351
rect 1719 1345 1725 1351
rect 97 1257 103 1263
rect 1731 1257 1737 1263
rect 85 1145 91 1151
rect 1719 1145 1725 1151
rect 97 1029 103 1035
rect 1731 1029 1737 1035
rect 85 949 91 955
rect 1719 949 1725 955
rect 97 833 103 839
rect 1731 833 1737 839
rect 85 749 91 755
rect 1719 749 1725 755
rect 97 637 103 643
rect 1731 637 1737 643
rect 85 557 91 563
rect 1719 557 1725 563
rect 97 437 103 443
rect 1731 437 1737 443
rect 85 317 91 323
rect 1719 317 1725 323
rect 97 245 103 251
rect 1731 245 1737 251
rect 85 169 91 175
rect 1719 169 1725 175
rect 97 117 103 123
rect 1731 117 1737 123
rect 85 77 91 83
rect 1719 77 1725 83
<< m5 >>
rect 84 1763 92 1800
rect 84 1757 85 1763
rect 91 1757 92 1763
rect 84 1671 92 1757
rect 84 1665 85 1671
rect 91 1665 92 1671
rect 84 1583 92 1665
rect 84 1577 85 1583
rect 91 1577 92 1583
rect 84 1499 92 1577
rect 84 1493 85 1499
rect 91 1493 92 1499
rect 84 1351 92 1493
rect 84 1345 85 1351
rect 91 1345 92 1351
rect 84 1151 92 1345
rect 84 1145 85 1151
rect 91 1145 92 1151
rect 84 955 92 1145
rect 84 949 85 955
rect 91 949 92 955
rect 84 755 92 949
rect 84 749 85 755
rect 91 749 92 755
rect 84 563 92 749
rect 84 557 85 563
rect 91 557 92 563
rect 84 323 92 557
rect 84 317 85 323
rect 91 317 92 323
rect 84 175 92 317
rect 84 169 85 175
rect 91 169 92 175
rect 84 83 92 169
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 1719 104 1800
rect 96 1713 97 1719
rect 103 1713 104 1719
rect 96 1623 104 1713
rect 96 1617 97 1623
rect 103 1617 104 1623
rect 96 1543 104 1617
rect 96 1537 97 1543
rect 103 1537 104 1543
rect 96 1431 104 1537
rect 96 1425 97 1431
rect 103 1425 104 1431
rect 96 1263 104 1425
rect 96 1257 97 1263
rect 103 1257 104 1263
rect 96 1035 104 1257
rect 96 1029 97 1035
rect 103 1029 104 1035
rect 96 839 104 1029
rect 96 833 97 839
rect 103 833 104 839
rect 96 643 104 833
rect 96 637 97 643
rect 103 637 104 643
rect 96 443 104 637
rect 96 437 97 443
rect 103 437 104 443
rect 96 251 104 437
rect 96 245 97 251
rect 103 245 104 251
rect 96 123 104 245
rect 96 117 97 123
rect 103 117 104 123
rect 96 72 104 117
rect 1718 1763 1726 1800
rect 1718 1757 1719 1763
rect 1725 1757 1726 1763
rect 1718 1671 1726 1757
rect 1718 1665 1719 1671
rect 1725 1665 1726 1671
rect 1718 1583 1726 1665
rect 1718 1577 1719 1583
rect 1725 1577 1726 1583
rect 1718 1499 1726 1577
rect 1718 1493 1719 1499
rect 1725 1493 1726 1499
rect 1718 1351 1726 1493
rect 1718 1345 1719 1351
rect 1725 1345 1726 1351
rect 1718 1151 1726 1345
rect 1718 1145 1719 1151
rect 1725 1145 1726 1151
rect 1718 955 1726 1145
rect 1718 949 1719 955
rect 1725 949 1726 955
rect 1718 755 1726 949
rect 1718 749 1719 755
rect 1725 749 1726 755
rect 1718 563 1726 749
rect 1718 557 1719 563
rect 1725 557 1726 563
rect 1718 323 1726 557
rect 1718 317 1719 323
rect 1725 317 1726 323
rect 1718 175 1726 317
rect 1718 169 1719 175
rect 1725 169 1726 175
rect 1718 83 1726 169
rect 1718 77 1719 83
rect 1725 77 1726 83
rect 1718 72 1726 77
rect 1730 1719 1738 1800
rect 1730 1713 1731 1719
rect 1737 1713 1738 1719
rect 1730 1623 1738 1713
rect 1730 1617 1731 1623
rect 1737 1617 1738 1623
rect 1730 1543 1738 1617
rect 1730 1537 1731 1543
rect 1737 1537 1738 1543
rect 1730 1431 1738 1537
rect 1730 1425 1731 1431
rect 1737 1425 1738 1431
rect 1730 1263 1738 1425
rect 1730 1257 1731 1263
rect 1737 1257 1738 1263
rect 1730 1035 1738 1257
rect 1730 1029 1731 1035
rect 1737 1029 1738 1035
rect 1730 839 1738 1029
rect 1730 833 1731 839
rect 1737 833 1738 839
rect 1730 643 1738 833
rect 1730 637 1731 643
rect 1737 637 1738 643
rect 1730 443 1738 637
rect 1730 437 1731 443
rect 1737 437 1738 443
rect 1730 251 1738 437
rect 1730 245 1731 251
rect 1737 245 1738 251
rect 1730 123 1738 245
rect 1730 117 1731 123
rect 1737 117 1738 123
rect 1730 72 1738 117
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__43
timestamp 1731220307
transform 1 0 1688 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220307
transform 1 0 104 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220307
transform 1 0 1688 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220307
transform 1 0 104 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220307
transform 1 0 1688 0 -1 1664
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220307
transform 1 0 104 0 -1 1664
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220307
transform 1 0 1688 0 1 1584
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220307
transform 1 0 104 0 1 1584
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220307
transform 1 0 1688 0 -1 1576
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220307
transform 1 0 104 0 -1 1576
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220307
transform 1 0 1688 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220307
transform 1 0 104 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220307
transform 1 0 1688 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220307
transform 1 0 104 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220307
transform 1 0 1688 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220307
transform 1 0 104 0 1 1368
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220307
transform 1 0 1688 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220307
transform 1 0 104 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220307
transform 1 0 1688 0 1 1172
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220307
transform 1 0 104 0 1 1172
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220307
transform 1 0 1688 0 -1 1124
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220307
transform 1 0 104 0 -1 1124
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220307
transform 1 0 1688 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220307
transform 1 0 104 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220307
transform 1 0 1688 0 -1 924
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220307
transform 1 0 104 0 -1 924
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220307
transform 1 0 1688 0 1 780
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220307
transform 1 0 104 0 1 780
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220307
transform 1 0 1688 0 -1 728
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220307
transform 1 0 104 0 -1 728
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220307
transform 1 0 1688 0 1 580
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220307
transform 1 0 104 0 1 580
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220307
transform 1 0 1688 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220307
transform 1 0 104 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220307
transform 1 0 1688 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220307
transform 1 0 104 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220307
transform 1 0 1688 0 -1 304
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220307
transform 1 0 104 0 -1 304
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220307
transform 1 0 1688 0 1 192
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220307
transform 1 0 104 0 1 192
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220307
transform 1 0 1688 0 -1 168
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220307
transform 1 0 104 0 -1 168
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220307
transform 1 0 1688 0 1 84
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220307
transform 1 0 104 0 1 84
box 7 3 12 24
use _0_0std_0_0cells_0_0INVX1  splt_ar0_ai
timestamp 1731220307
transform 1 0 1472 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  splt_ar0_an
timestamp 1731220307
transform 1 0 1464 0 1 776
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_55_6
timestamp 1731220307
transform 1 0 1056 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_54_6
timestamp 1731220307
transform 1 0 1024 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_53_6
timestamp 1731220307
transform 1 0 960 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_52_6
timestamp 1731220307
transform 1 0 928 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_51_6
timestamp 1731220307
transform 1 0 1120 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ad_ainvs_50_6
timestamp 1731220307
transform 1 0 1152 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ac__latch__inv
timestamp 1731220307
transform 1 0 1280 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0OR2X1  splt_ar2_an
timestamp 1731220307
transform 1 0 1448 0 -1 928
box 4 4 48 48
use _0_0std_0_0cells_0_0INVX1  splt_ar1_ai
timestamp 1731220307
transform 1 0 1240 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  splt_ar1_an
timestamp 1731220307
transform 1 0 1200 0 -1 732
box 4 6 36 48
use _0_0cell_0_0ginvx0  splt_ac_acx1
timestamp 1731220307
transform 1 0 1288 0 1 776
box 8 6 28 32
use _0_0cell_0_0gcelem3x0  splt_ac_acx0
timestamp 1731220307
transform 1 0 1320 0 1 752
box 8 5 92 72
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_544_6
timestamp 1731220307
transform 1 0 1024 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_543_6
timestamp 1731220307
transform 1 0 992 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_542_6
timestamp 1731220307
transform 1 0 1056 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_541_6
timestamp 1731220307
transform 1 0 1048 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_540_6
timestamp 1731220307
transform 1 0 976 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_539_6
timestamp 1731220307
transform 1 0 952 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_538_6
timestamp 1731220307
transform 1 0 1144 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_537_6
timestamp 1731220307
transform 1 0 1136 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_536_6
timestamp 1731220307
transform 1 0 1096 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_535_6
timestamp 1731220307
transform 1 0 1176 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_534_6
timestamp 1731220307
transform 1 0 1216 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_533_6
timestamp 1731220307
transform 1 0 1256 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_532_6
timestamp 1731220307
transform 1 0 1320 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_531_6
timestamp 1731220307
transform 1 0 1232 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_530_6
timestamp 1731220307
transform 1 0 1168 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_529_6
timestamp 1731220307
transform 1 0 1112 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_528_6
timestamp 1731220307
transform 1 0 1048 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_527_6
timestamp 1731220307
transform 1 0 1216 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_526_6
timestamp 1731220307
transform 1 0 1264 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_525_6
timestamp 1731220307
transform 1 0 1304 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_524_6
timestamp 1731220307
transform 1 0 1336 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_523_6
timestamp 1731220307
transform 1 0 1368 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_522_6
timestamp 1731220307
transform 1 0 1400 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_521_6
timestamp 1731220307
transform 1 0 1432 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_520_6
timestamp 1731220307
transform 1 0 1472 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_519_6
timestamp 1731220307
transform 1 0 1512 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_518_6
timestamp 1731220307
transform 1 0 1496 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_517_6
timestamp 1731220307
transform 1 0 1408 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_516_6
timestamp 1731220307
transform 1 0 1584 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_515_6
timestamp 1731220307
transform 1 0 1552 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_514_6
timestamp 1731220307
transform 1 0 1512 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_513_6
timestamp 1731220307
transform 1 0 1472 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_512_6
timestamp 1731220307
transform 1 0 1432 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_511_6
timestamp 1731220307
transform 1 0 1400 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_510_6
timestamp 1731220307
transform 1 0 1368 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_59_6
timestamp 1731220307
transform 1 0 1336 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_58_6
timestamp 1731220307
transform 1 0 1296 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_57_6
timestamp 1731220307
transform 1 0 1512 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_56_6
timestamp 1731220307
transform 1 0 1472 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_55_6
timestamp 1731220307
transform 1 0 1440 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_54_6
timestamp 1731220307
transform 1 0 1408 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_53_6
timestamp 1731220307
transform 1 0 1376 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_52_6
timestamp 1731220307
transform 1 0 1344 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_51_6
timestamp 1731220307
transform 1 0 1312 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  splt_ap_ainvs_50_6
timestamp 1731220307
transform 1 0 1312 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  splt_ap_aand
timestamp 1731220307
transform 1 0 1016 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0OR2X1  splt_ar3_an
timestamp 1731220307
transform 1 0 1224 0 1 776
box 4 4 48 48
use _0_0std_0_0cells_0_0AND2X1  splt_ar1__r
timestamp 1731220307
transform 1 0 1232 0 1 956
box 8 4 52 52
use _0_0std_0_0cells_0_0LATCHINV  splt_ac__latch_al
timestamp 1731220307
transform 1 0 1160 0 -1 1144
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  splt_ac__latch_anx
timestamp 1731220307
transform 1 0 1240 0 -1 1132
box 4 6 36 64
use _0_0std_0_0cells_0_0AND2X1  splt_ar2__r
timestamp 1731220307
transform 1 0 1104 0 1 956
box 8 4 52 52
use _0_0std_0_0cells_0_0NOR2X1  splt_anor__ra
timestamp 1731220307
transform 1 0 1416 0 1 776
box 4 6 36 48
use _0_0std_0_0cells_0_0LATCH  splt_alatch_57_6
timestamp 1731220307
transform 1 0 1208 0 1 336
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_56_6
timestamp 1731220307
transform 1 0 1088 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_55_6
timestamp 1731220307
transform 1 0 784 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_54_6
timestamp 1731220307
transform 1 0 744 0 1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_53_6
timestamp 1731220307
transform 1 0 888 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_52_6
timestamp 1731220307
transform 1 0 792 0 1 764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_51_6
timestamp 1731220307
transform 1 0 688 0 1 956
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  splt_alatch_50_6
timestamp 1731220307
transform 1 0 824 0 -1 1140
box 8 5 100 68
use _0_0std_0_0cells_0_0INVX1  snk_ar_ai
timestamp 1731220307
transform 1 0 1288 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  snk_ar_an
timestamp 1731220307
transform 1 0 1320 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_569_6
timestamp 1731220307
transform 1 0 864 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_568_6
timestamp 1731220307
transform 1 0 768 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_567_6
timestamp 1731220307
transform 1 0 648 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_566_6
timestamp 1731220307
transform 1 0 528 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_565_6
timestamp 1731220307
transform 1 0 456 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_564_6
timestamp 1731220307
transform 1 0 360 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_563_6
timestamp 1731220307
transform 1 0 296 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_562_6
timestamp 1731220307
transform 1 0 272 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_561_6
timestamp 1731220307
transform 1 0 216 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_560_6
timestamp 1731220307
transform 1 0 168 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_559_6
timestamp 1731220307
transform 1 0 128 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_558_6
timestamp 1731220307
transform 1 0 280 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_557_6
timestamp 1731220307
transform 1 0 224 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_556_6
timestamp 1731220307
transform 1 0 160 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_555_6
timestamp 1731220307
transform 1 0 128 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_554_6
timestamp 1731220307
transform 1 0 128 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_553_6
timestamp 1731220307
transform 1 0 160 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_552_6
timestamp 1731220307
transform 1 0 192 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_551_6
timestamp 1731220307
transform 1 0 240 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_550_6
timestamp 1731220307
transform 1 0 560 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_549_6
timestamp 1731220307
transform 1 0 432 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_548_6
timestamp 1731220307
transform 1 0 320 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_547_6
timestamp 1731220307
transform 1 0 256 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_546_6
timestamp 1731220307
transform 1 0 168 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_545_6
timestamp 1731220307
transform 1 0 128 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_544_6
timestamp 1731220307
transform 1 0 704 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_543_6
timestamp 1731220307
transform 1 0 536 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_542_6
timestamp 1731220307
transform 1 0 384 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_541_6
timestamp 1731220307
transform 1 0 312 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_540_6
timestamp 1731220307
transform 1 0 240 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_539_6
timestamp 1731220307
transform 1 0 184 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_538_6
timestamp 1731220307
transform 1 0 648 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_537_6
timestamp 1731220307
transform 1 0 520 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_536_6
timestamp 1731220307
transform 1 0 408 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_535_6
timestamp 1731220307
transform 1 0 208 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_534_6
timestamp 1731220307
transform 1 0 176 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_533_6
timestamp 1731220307
transform 1 0 144 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_532_6
timestamp 1731220307
transform 1 0 240 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_531_6
timestamp 1731220307
transform 1 0 272 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_530_6
timestamp 1731220307
transform 1 0 304 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_529_6
timestamp 1731220307
transform 1 0 336 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_528_6
timestamp 1731220307
transform 1 0 368 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_527_6
timestamp 1731220307
transform 1 0 400 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_526_6
timestamp 1731220307
transform 1 0 432 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_525_6
timestamp 1731220307
transform 1 0 464 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_524_6
timestamp 1731220307
transform 1 0 496 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_523_6
timestamp 1731220307
transform 1 0 528 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_522_6
timestamp 1731220307
transform 1 0 560 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_521_6
timestamp 1731220307
transform 1 0 592 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_520_6
timestamp 1731220307
transform 1 0 624 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_519_6
timestamp 1731220307
transform 1 0 656 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_518_6
timestamp 1731220307
transform 1 0 688 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_517_6
timestamp 1731220307
transform 1 0 720 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_516_6
timestamp 1731220307
transform 1 0 752 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_515_6
timestamp 1731220307
transform 1 0 784 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_514_6
timestamp 1731220307
transform 1 0 816 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_513_6
timestamp 1731220307
transform 1 0 848 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_512_6
timestamp 1731220307
transform 1 0 880 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_511_6
timestamp 1731220307
transform 1 0 912 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_510_6
timestamp 1731220307
transform 1 0 944 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_59_6
timestamp 1731220307
transform 1 0 976 0 -1 1760
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_58_6
timestamp 1731220307
transform 1 0 1040 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_57_6
timestamp 1731220307
transform 1 0 912 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_56_6
timestamp 1731220307
transform 1 0 784 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_55_6
timestamp 1731220307
transform 1 0 872 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_54_6
timestamp 1731220307
transform 1 0 1032 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_53_6
timestamp 1731220307
transform 1 0 992 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_52_6
timestamp 1731220307
transform 1 0 1056 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_51_6
timestamp 1731220307
transform 1 0 1072 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad_ainvs_50_6
timestamp 1731220307
transform 1 0 1072 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_57_6
timestamp 1731220307
transform 1 0 896 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_56_6
timestamp 1731220307
transform 1 0 1056 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_55_6
timestamp 1731220307
transform 1 0 784 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_54_6
timestamp 1731220307
transform 1 0 664 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_53_6
timestamp 1731220307
transform 1 0 856 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_52_6
timestamp 1731220307
transform 1 0 552 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_51_6
timestamp 1731220307
transform 1 0 808 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ainv_50_6
timestamp 1731220307
transform 1 0 912 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar2_an
timestamp 1731220307
transform 1 0 1056 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  m_ar1_ai
timestamp 1731220307
transform 1 0 1032 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar1_an
timestamp 1731220307
transform 1 0 1064 0 -1 928
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  m_ar3_ai
timestamp 1731220307
transform 1 0 1432 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar3_an
timestamp 1731220307
transform 1 0 1360 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0AND2X1  m_aand__ct
timestamp 1731220307
transform 1 0 1360 0 -1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0OR2X1  m_aor__ca
timestamp 1731220307
transform 1 0 1008 0 1 776
box 4 4 48 48
use _0_0std_0_0cells_0_0INVX1  m_ar0_ai
timestamp 1731220307
transform 1 0 1160 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar0_an
timestamp 1731220307
transform 1 0 1192 0 1 968
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  m_ar4_ai
timestamp 1731220307
transform 1 0 1128 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  m_ar4_an
timestamp 1731220307
transform 1 0 1088 0 -1 1128
box 4 6 36 48
use _0_0cell_0_0ginvx0  m_ac1_acx1
timestamp 1731220307
transform 1 0 1104 0 -1 928
box 8 6 28 32
use _0_0cell_0_0gcelem3x0  m_ac1_acx0
timestamp 1731220307
transform 1 0 1136 0 -1 952
box 8 5 92 72
use _0_0cell_0_0ginvx0  m_ac0_acx1
timestamp 1731220307
transform 1 0 1232 0 -1 928
box 8 6 28 32
use _0_0cell_0_0gcelem3x0  m_ac0_acx0
timestamp 1731220307
transform 1 0 1264 0 -1 952
box 8 5 92 72
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_544_6
timestamp 1731220307
transform 1 0 544 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_543_6
timestamp 1731220307
transform 1 0 632 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_542_6
timestamp 1731220307
transform 1 0 600 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_541_6
timestamp 1731220307
transform 1 0 680 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_540_6
timestamp 1731220307
transform 1 0 768 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_539_6
timestamp 1731220307
transform 1 0 856 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_538_6
timestamp 1731220307
transform 1 0 896 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_537_6
timestamp 1731220307
transform 1 0 816 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_536_6
timestamp 1731220307
transform 1 0 736 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_535_6
timestamp 1731220307
transform 1 0 664 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_534_6
timestamp 1731220307
transform 1 0 600 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_533_6
timestamp 1731220307
transform 1 0 544 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_532_6
timestamp 1731220307
transform 1 0 512 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_531_6
timestamp 1731220307
transform 1 0 480 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_530_6
timestamp 1731220307
transform 1 0 448 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_529_6
timestamp 1731220307
transform 1 0 416 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_528_6
timestamp 1731220307
transform 1 0 384 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_527_6
timestamp 1731220307
transform 1 0 352 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_526_6
timestamp 1731220307
transform 1 0 320 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_525_6
timestamp 1731220307
transform 1 0 288 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_524_6
timestamp 1731220307
transform 1 0 256 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_523_6
timestamp 1731220307
transform 1 0 224 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_522_6
timestamp 1731220307
transform 1 0 192 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_521_6
timestamp 1731220307
transform 1 0 160 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_520_6
timestamp 1731220307
transform 1 0 128 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_519_6
timestamp 1731220307
transform 1 0 128 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_518_6
timestamp 1731220307
transform 1 0 160 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_517_6
timestamp 1731220307
transform 1 0 208 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_516_6
timestamp 1731220307
transform 1 0 256 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_515_6
timestamp 1731220307
transform 1 0 304 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_514_6
timestamp 1731220307
transform 1 0 360 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_513_6
timestamp 1731220307
transform 1 0 408 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_512_6
timestamp 1731220307
transform 1 0 464 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_511_6
timestamp 1731220307
transform 1 0 528 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_510_6
timestamp 1731220307
transform 1 0 592 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_59_6
timestamp 1731220307
transform 1 0 560 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_58_6
timestamp 1731220307
transform 1 0 528 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_57_6
timestamp 1731220307
transform 1 0 496 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_56_6
timestamp 1731220307
transform 1 0 512 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_55_6
timestamp 1731220307
transform 1 0 480 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_54_6
timestamp 1731220307
transform 1 0 448 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_53_6
timestamp 1731220307
transform 1 0 416 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_52_6
timestamp 1731220307
transform 1 0 384 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_51_6
timestamp 1731220307
transform 1 0 408 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ap_ainvs_50_6
timestamp 1731220307
transform 1 0 440 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  m_ap_aand
timestamp 1731220307
transform 1 0 472 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  m_aand__cf
timestamp 1731220307
transform 1 0 1152 0 1 764
box 8 4 52 52
use _0_0std_0_0cells_0_0INVX1  m_ainv__cd
timestamp 1731220307
transform 1 0 1096 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad__cd_ainvs_51_6
timestamp 1731220307
transform 1 0 1416 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  m_ad__cd_ainvs_50_6
timestamp 1731220307
transform 1 0 1400 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0LATCH  m_alatch_57_6
timestamp 1731220307
transform 1 0 680 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_56_6
timestamp 1731220307
transform 1 0 944 0 1 176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_55_6
timestamp 1731220307
transform 1 0 672 0 1 176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_54_6
timestamp 1731220307
transform 1 0 512 0 1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_53_6
timestamp 1731220307
transform 1 0 592 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_52_6
timestamp 1731220307
transform 1 0 384 0 1 764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_51_6
timestamp 1731220307
transform 1 0 704 0 -1 940
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  m_alatch_50_6
timestamp 1731220307
transform 1 0 840 0 -1 940
box 8 5 100 68
use _0_0std_0_0cells_0_0MUX2X1  m_amux_57_6
timestamp 1731220307
transform 1 0 1344 0 1 336
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_56_6
timestamp 1731220307
transform 1 0 1192 0 -1 320
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_55_6
timestamp 1731220307
transform 1 0 824 0 1 176
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_54_6
timestamp 1731220307
transform 1 0 760 0 -1 744
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_53_6
timestamp 1731220307
transform 1 0 992 0 -1 744
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_52_6
timestamp 1731220307
transform 1 0 648 0 1 764
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_51_6
timestamp 1731220307
transform 1 0 808 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0MUX2X1  m_amux_50_6
timestamp 1731220307
transform 1 0 960 0 1 956
box 8 4 80 64
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_55_6
timestamp 1731220307
transform 1 0 1432 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_54_6
timestamp 1731220307
transform 1 0 1392 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_53_6
timestamp 1731220307
transform 1 0 1312 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_52_6
timestamp 1731220307
transform 1 0 1264 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_51_6
timestamp 1731220307
transform 1 0 1232 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ad_ainvs_50_6
timestamp 1731220307
transform 1 0 1160 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ar0_ai
timestamp 1731220307
transform 1 0 968 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  c_ar0_an
timestamp 1731220307
transform 1 0 888 0 -1 1480
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_544_6
timestamp 1731220307
transform 1 0 256 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_543_6
timestamp 1731220307
transform 1 0 224 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_542_6
timestamp 1731220307
transform 1 0 192 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_541_6
timestamp 1731220307
transform 1 0 224 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_540_6
timestamp 1731220307
transform 1 0 192 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_539_6
timestamp 1731220307
transform 1 0 160 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_538_6
timestamp 1731220307
transform 1 0 128 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_537_6
timestamp 1731220307
transform 1 0 288 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_536_6
timestamp 1731220307
transform 1 0 320 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_535_6
timestamp 1731220307
transform 1 0 352 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_534_6
timestamp 1731220307
transform 1 0 384 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_533_6
timestamp 1731220307
transform 1 0 512 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_532_6
timestamp 1731220307
transform 1 0 480 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_531_6
timestamp 1731220307
transform 1 0 448 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_530_6
timestamp 1731220307
transform 1 0 416 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_529_6
timestamp 1731220307
transform 1 0 480 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_528_6
timestamp 1731220307
transform 1 0 448 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_527_6
timestamp 1731220307
transform 1 0 416 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_526_6
timestamp 1731220307
transform 1 0 384 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_525_6
timestamp 1731220307
transform 1 0 352 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_524_6
timestamp 1731220307
transform 1 0 320 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_523_6
timestamp 1731220307
transform 1 0 288 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_522_6
timestamp 1731220307
transform 1 0 256 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_521_6
timestamp 1731220307
transform 1 0 224 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_520_6
timestamp 1731220307
transform 1 0 192 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_519_6
timestamp 1731220307
transform 1 0 160 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_518_6
timestamp 1731220307
transform 1 0 128 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_517_6
timestamp 1731220307
transform 1 0 128 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_516_6
timestamp 1731220307
transform 1 0 160 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_515_6
timestamp 1731220307
transform 1 0 192 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_514_6
timestamp 1731220307
transform 1 0 224 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_513_6
timestamp 1731220307
transform 1 0 256 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_512_6
timestamp 1731220307
transform 1 0 288 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_511_6
timestamp 1731220307
transform 1 0 320 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_510_6
timestamp 1731220307
transform 1 0 448 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_59_6
timestamp 1731220307
transform 1 0 416 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_58_6
timestamp 1731220307
transform 1 0 384 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_57_6
timestamp 1731220307
transform 1 0 352 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_56_6
timestamp 1731220307
transform 1 0 544 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_55_6
timestamp 1731220307
transform 1 0 512 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_54_6
timestamp 1731220307
transform 1 0 480 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_53_6
timestamp 1731220307
transform 1 0 424 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_52_6
timestamp 1731220307
transform 1 0 392 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_51_6
timestamp 1731220307
transform 1 0 456 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c_ap_ainvs_50_6
timestamp 1731220307
transform 1 0 488 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  c_ap_aand
timestamp 1731220307
transform 1 0 312 0 1 956
box 8 4 52 52
use _0_0cell_0_0ginvx0  c_ac_acx1
timestamp 1731220307
transform 1 0 768 0 -1 1480
box 8 6 28 32
use _0_0cell_0_0gcelem2x0  c_ac_acx0
timestamp 1731220307
transform 1 0 800 0 -1 1496
box 8 4 84 60
use _0_0std_0_0cells_0_0OR2X1  c_ar2_an
timestamp 1731220307
transform 1 0 1016 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  c_ar1_an
timestamp 1731220307
transform 1 0 1104 0 -1 1480
box 4 4 48 48
use _0_0cell_0_0gcelem2x0  c_ac__ra_acx0
timestamp 1731220307
transform 1 0 928 0 -1 1496
box 8 4 84 60
use _0_0std_0_0cells_0_0LATCH  c_alatch_57_6
timestamp 1731220307
transform 1 0 576 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_56_6
timestamp 1731220307
transform 1 0 888 0 -1 320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_55_6
timestamp 1731220307
transform 1 0 648 0 1 336
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_54_6
timestamp 1731220307
transform 1 0 280 0 -1 552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_53_6
timestamp 1731220307
transform 1 0 264 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_52_6
timestamp 1731220307
transform 1 0 208 0 1 764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_51_6
timestamp 1731220307
transform 1 0 568 0 -1 940
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  c_alatch_50_6
timestamp 1731220307
transform 1 0 560 0 1 956
box 8 5 100 68
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_569_6
timestamp 1731220307
transform 1 0 1272 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_568_6
timestamp 1731220307
transform 1 0 1304 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_567_6
timestamp 1731220307
transform 1 0 1336 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_566_6
timestamp 1731220307
transform 1 0 1368 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_565_6
timestamp 1731220307
transform 1 0 1400 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_564_6
timestamp 1731220307
transform 1 0 1432 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_563_6
timestamp 1731220307
transform 1 0 1408 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_562_6
timestamp 1731220307
transform 1 0 1416 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_561_6
timestamp 1731220307
transform 1 0 1472 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_560_6
timestamp 1731220307
transform 1 0 1520 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_559_6
timestamp 1731220307
transform 1 0 1568 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_558_6
timestamp 1731220307
transform 1 0 1552 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_557_6
timestamp 1731220307
transform 1 0 1512 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_556_6
timestamp 1731220307
transform 1 0 1472 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_555_6
timestamp 1731220307
transform 1 0 1552 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_554_6
timestamp 1731220307
transform 1 0 1584 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_553_6
timestamp 1731220307
transform 1 0 1584 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_552_6
timestamp 1731220307
transform 1 0 1584 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_551_6
timestamp 1731220307
transform 1 0 1552 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_550_6
timestamp 1731220307
transform 1 0 1616 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_549_6
timestamp 1731220307
transform 1 0 1648 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_548_6
timestamp 1731220307
transform 1 0 1648 0 -1 172
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_547_6
timestamp 1731220307
transform 1 0 1616 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_546_6
timestamp 1731220307
transform 1 0 1648 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_545_6
timestamp 1731220307
transform 1 0 1648 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_544_6
timestamp 1731220307
transform 1 0 1616 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_543_6
timestamp 1731220307
transform 1 0 1648 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_542_6
timestamp 1731220307
transform 1 0 1616 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_541_6
timestamp 1731220307
transform 1 0 1584 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_540_6
timestamp 1731220307
transform 1 0 1616 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_539_6
timestamp 1731220307
transform 1 0 1648 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_538_6
timestamp 1731220307
transform 1 0 1648 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_537_6
timestamp 1731220307
transform 1 0 1600 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_536_6
timestamp 1731220307
transform 1 0 1536 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_535_6
timestamp 1731220307
transform 1 0 1472 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_534_6
timestamp 1731220307
transform 1 0 1648 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_533_6
timestamp 1731220307
transform 1 0 1616 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_532_6
timestamp 1731220307
transform 1 0 1584 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_531_6
timestamp 1731220307
transform 1 0 1552 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_530_6
timestamp 1731220307
transform 1 0 1512 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_529_6
timestamp 1731220307
transform 1 0 1472 0 -1 732
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_528_6
timestamp 1731220307
transform 1 0 1512 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_527_6
timestamp 1731220307
transform 1 0 1552 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_526_6
timestamp 1731220307
transform 1 0 1584 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_525_6
timestamp 1731220307
transform 1 0 1616 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_524_6
timestamp 1731220307
transform 1 0 1648 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_523_6
timestamp 1731220307
transform 1 0 1648 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_522_6
timestamp 1731220307
transform 1 0 1616 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_521_6
timestamp 1731220307
transform 1 0 1584 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_520_6
timestamp 1731220307
transform 1 0 1552 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_519_6
timestamp 1731220307
transform 1 0 1512 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_518_6
timestamp 1731220307
transform 1 0 1648 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_517_6
timestamp 1731220307
transform 1 0 1616 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_516_6
timestamp 1731220307
transform 1 0 1584 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_515_6
timestamp 1731220307
transform 1 0 1552 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_514_6
timestamp 1731220307
transform 1 0 1512 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_513_6
timestamp 1731220307
transform 1 0 1512 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_512_6
timestamp 1731220307
transform 1 0 1552 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_511_6
timestamp 1731220307
transform 1 0 1552 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_510_6
timestamp 1731220307
transform 1 0 1512 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_59_6
timestamp 1731220307
transform 1 0 1520 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_58_6
timestamp 1731220307
transform 1 0 1528 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_57_6
timestamp 1731220307
transform 1 0 1512 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_56_6
timestamp 1731220307
transform 1 0 1472 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_55_6
timestamp 1731220307
transform 1 0 1512 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_54_6
timestamp 1731220307
transform 1 0 1528 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_53_6
timestamp 1731220307
transform 1 0 1464 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_52_6
timestamp 1731220307
transform 1 0 1392 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_51_6
timestamp 1731220307
transform 1 0 1240 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ad_ainvs_50_6
timestamp 1731220307
transform 1 0 1168 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ar0_ai
timestamp 1731220307
transform 1 0 1016 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  a_ar0_an
timestamp 1731220307
transform 1 0 1056 0 1 1364
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_544_6
timestamp 1731220307
transform 1 0 160 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_543_6
timestamp 1731220307
transform 1 0 160 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_542_6
timestamp 1731220307
transform 1 0 224 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_541_6
timestamp 1731220307
transform 1 0 256 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_540_6
timestamp 1731220307
transform 1 0 288 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_539_6
timestamp 1731220307
transform 1 0 320 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_538_6
timestamp 1731220307
transform 1 0 352 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_537_6
timestamp 1731220307
transform 1 0 336 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_536_6
timestamp 1731220307
transform 1 0 464 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_535_6
timestamp 1731220307
transform 1 0 432 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_534_6
timestamp 1731220307
transform 1 0 400 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_533_6
timestamp 1731220307
transform 1 0 368 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_532_6
timestamp 1731220307
transform 1 0 304 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_531_6
timestamp 1731220307
transform 1 0 272 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_530_6
timestamp 1731220307
transform 1 0 240 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_529_6
timestamp 1731220307
transform 1 0 208 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_528_6
timestamp 1731220307
transform 1 0 176 0 1 188
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_527_6
timestamp 1731220307
transform 1 0 256 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_526_6
timestamp 1731220307
transform 1 0 224 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_525_6
timestamp 1731220307
transform 1 0 192 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_524_6
timestamp 1731220307
transform 1 0 160 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_523_6
timestamp 1731220307
transform 1 0 128 0 -1 308
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_522_6
timestamp 1731220307
transform 1 0 192 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_521_6
timestamp 1731220307
transform 1 0 160 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_520_6
timestamp 1731220307
transform 1 0 128 0 1 348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_519_6
timestamp 1731220307
transform 1 0 128 0 -1 540
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_518_6
timestamp 1731220307
transform 1 0 128 0 1 576
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_517_6
timestamp 1731220307
transform 1 0 128 0 1 776
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_516_6
timestamp 1731220307
transform 1 0 128 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_515_6
timestamp 1731220307
transform 1 0 128 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_514_6
timestamp 1731220307
transform 1 0 160 0 1 968
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_513_6
timestamp 1731220307
transform 1 0 256 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_512_6
timestamp 1731220307
transform 1 0 544 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_511_6
timestamp 1731220307
transform 1 0 544 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_510_6
timestamp 1731220307
transform 1 0 512 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_59_6
timestamp 1731220307
transform 1 0 576 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_58_6
timestamp 1731220307
transform 1 0 608 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_57_6
timestamp 1731220307
transform 1 0 640 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_56_6
timestamp 1731220307
transform 1 0 640 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_55_6
timestamp 1731220307
transform 1 0 608 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_54_6
timestamp 1731220307
transform 1 0 576 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_53_6
timestamp 1731220307
transform 1 0 520 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_52_6
timestamp 1731220307
transform 1 0 552 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_51_6
timestamp 1731220307
transform 1 0 584 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  a_ap_ainvs_50_6
timestamp 1731220307
transform 1 0 736 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  a_ap_aand
timestamp 1731220307
transform 1 0 944 0 1 1156
box 8 4 52 52
use _0_0cell_0_0ginvx0  a_ac_acx1
timestamp 1731220307
transform 1 0 1104 0 1 1364
box 8 6 28 32
use _0_0cell_0_0gcelem3x0  a_ac_acx0
timestamp 1731220307
transform 1 0 1056 0 -1 1348
box 8 5 92 72
use _0_0std_0_0cells_0_0NOR2X1  a_ar2_an
timestamp 1731220307
transform 1 0 1016 0 -1 1324
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  a_ar1_ai
timestamp 1731220307
transform 1 0 1192 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  a_ar1_an
timestamp 1731220307
transform 1 0 1144 0 1 1364
box 4 6 36 48
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_57_6_al
timestamp 1731220307
transform 1 0 1200 0 1 560
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_57_6_anx
timestamp 1731220307
transform 1 0 1328 0 1 572
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_56_6_al
timestamp 1731220307
transform 1 0 1088 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_56_6_anx
timestamp 1731220307
transform 1 0 1192 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_55_6_al
timestamp 1731220307
transform 1 0 640 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_55_6_anx
timestamp 1731220307
transform 1 0 720 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_54_6_al
timestamp 1731220307
transform 1 0 384 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_54_6_anx
timestamp 1731220307
transform 1 0 464 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_53_6_al
timestamp 1731220307
transform 1 0 392 0 1 560
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_53_6_anx
timestamp 1731220307
transform 1 0 384 0 -1 736
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_52_6_al
timestamp 1731220307
transform 1 0 312 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_52_6_anx
timestamp 1731220307
transform 1 0 392 0 -1 932
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_51_6_al
timestamp 1731220307
transform 1 0 1000 0 1 1152
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_51_6_anx
timestamp 1731220307
transform 1 0 1080 0 1 1164
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__b_50_6_al
timestamp 1731220307
transform 1 0 816 0 -1 1340
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__b_50_6_anx
timestamp 1731220307
transform 1 0 832 0 1 1360
box 4 6 36 64
use _0_0std_0_0cells_0_0FAX1  a_aadder_57_6
timestamp 1731220307
transform 1 0 1256 0 -1 560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_56_6
timestamp 1731220307
transform 1 0 1072 0 1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_55_6
timestamp 1731220307
transform 1 0 752 0 1 328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_54_6
timestamp 1731220307
transform 1 0 504 0 -1 560
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_53_6
timestamp 1731220307
transform 1 0 440 0 -1 752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_52_6
timestamp 1731220307
transform 1 0 432 0 -1 948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_51_6
timestamp 1731220307
transform 1 0 656 0 -1 1148
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  a_aadder_50_6
timestamp 1731220307
transform 1 0 808 0 1 1148
box 3 5 132 108
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_57_6_al
timestamp 1731220307
transform 1 0 1080 0 -1 748
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_57_6_anx
timestamp 1731220307
transform 1 0 1160 0 -1 736
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_56_6_al
timestamp 1731220307
transform 1 0 984 0 1 560
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_56_6_anx
timestamp 1731220307
transform 1 0 1112 0 1 572
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_55_6_al
timestamp 1731220307
transform 1 0 768 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_55_6_anx
timestamp 1731220307
transform 1 0 864 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_54_6_al
timestamp 1731220307
transform 1 0 160 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_54_6_anx
timestamp 1731220307
transform 1 0 240 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_53_6_al
timestamp 1731220307
transform 1 0 128 0 -1 748
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_53_6_anx
timestamp 1731220307
transform 1 0 208 0 -1 736
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_52_6_al
timestamp 1731220307
transform 1 0 392 0 1 952
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_52_6_anx
timestamp 1731220307
transform 1 0 496 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_51_6_al
timestamp 1731220307
transform 1 0 896 0 -1 1340
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_51_6_anx
timestamp 1731220307
transform 1 0 976 0 -1 1328
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  a_alatch__a_50_6_al
timestamp 1731220307
transform 1 0 880 0 1 1348
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  a_alatch__a_50_6_anx
timestamp 1731220307
transform 1 0 968 0 1 1360
box 4 6 36 64
use _0_0std_0_0cells_0_0TIELOX1  a_atlo
timestamp 1731220307
transform 1 0 800 0 1 1364
box 8 6 28 37
use _0_0std_0_0cells_0_0OR2X1  i_ar0_an
timestamp 1731220307
transform 1 0 1456 0 1 1364
box 4 4 48 48
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_55_6
timestamp 1731220307
transform 1 0 1352 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_54_6
timestamp 1731220307
transform 1 0 1352 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_53_6
timestamp 1731220307
transform 1 0 1320 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_52_6
timestamp 1731220307
transform 1 0 1240 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_51_6
timestamp 1731220307
transform 1 0 1120 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ad_ainvs_50_6
timestamp 1731220307
transform 1 0 1152 0 -1 1580
box 8 7 28 34
use _0_0cell_0_0ginvx0  i_ac_acx1
timestamp 1731220307
transform 1 0 1272 0 -1 1480
box 8 6 28 32
use _0_0cell_0_0gcelem2x0  i_ac_acx0
timestamp 1731220307
transform 1 0 1312 0 1 1348
box 8 4 84 60
use _0_0std_0_0cells_0_0INVX1  i_ar1_ai
timestamp 1731220307
transform 1 0 1192 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0OR2X1  i_ar1_an
timestamp 1731220307
transform 1 0 1240 0 1 1364
box 4 4 48 48
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_544_6
timestamp 1731220307
transform 1 0 656 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_543_6
timestamp 1731220307
transform 1 0 696 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_542_6
timestamp 1731220307
transform 1 0 680 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_541_6
timestamp 1731220307
transform 1 0 600 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_540_6
timestamp 1731220307
transform 1 0 616 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_539_6
timestamp 1731220307
transform 1 0 672 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_538_6
timestamp 1731220307
transform 1 0 672 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_537_6
timestamp 1731220307
transform 1 0 704 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_536_6
timestamp 1731220307
transform 1 0 736 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_535_6
timestamp 1731220307
transform 1 0 704 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_534_6
timestamp 1731220307
transform 1 0 672 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_533_6
timestamp 1731220307
transform 1 0 640 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_532_6
timestamp 1731220307
transform 1 0 608 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_531_6
timestamp 1731220307
transform 1 0 576 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_530_6
timestamp 1731220307
transform 1 0 544 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_529_6
timestamp 1731220307
transform 1 0 512 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_528_6
timestamp 1731220307
transform 1 0 480 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_527_6
timestamp 1731220307
transform 1 0 448 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_526_6
timestamp 1731220307
transform 1 0 416 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_525_6
timestamp 1731220307
transform 1 0 384 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_524_6
timestamp 1731220307
transform 1 0 352 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_523_6
timestamp 1731220307
transform 1 0 320 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_522_6
timestamp 1731220307
transform 1 0 288 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_521_6
timestamp 1731220307
transform 1 0 256 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_520_6
timestamp 1731220307
transform 1 0 224 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_519_6
timestamp 1731220307
transform 1 0 192 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_518_6
timestamp 1731220307
transform 1 0 160 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_517_6
timestamp 1731220307
transform 1 0 128 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_516_6
timestamp 1731220307
transform 1 0 168 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_515_6
timestamp 1731220307
transform 1 0 200 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_514_6
timestamp 1731220307
transform 1 0 232 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_513_6
timestamp 1731220307
transform 1 0 264 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_512_6
timestamp 1731220307
transform 1 0 328 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_511_6
timestamp 1731220307
transform 1 0 328 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_510_6
timestamp 1731220307
transform 1 0 392 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_59_6
timestamp 1731220307
transform 1 0 336 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_58_6
timestamp 1731220307
transform 1 0 392 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_57_6
timestamp 1731220307
transform 1 0 448 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_56_6
timestamp 1731220307
transform 1 0 504 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_55_6
timestamp 1731220307
transform 1 0 568 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_54_6
timestamp 1731220307
transform 1 0 704 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_53_6
timestamp 1731220307
transform 1 0 848 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_52_6
timestamp 1731220307
transform 1 0 952 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_51_6
timestamp 1731220307
transform 1 0 848 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  i_ap_ainvs_50_6
timestamp 1731220307
transform 1 0 744 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  i_ap_aand
timestamp 1731220307
transform 1 0 704 0 1 1352
box 8 4 52 52
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_57_6_al
timestamp 1731220307
transform 1 0 920 0 -1 556
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_57_6_anx
timestamp 1731220307
transform 1 0 896 0 1 572
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_56_6_al
timestamp 1731220307
transform 1 0 936 0 1 332
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_56_6_anx
timestamp 1731220307
transform 1 0 1024 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_55_6_al
timestamp 1731220307
transform 1 0 528 0 1 332
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_55_6_anx
timestamp 1731220307
transform 1 0 608 0 1 344
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_54_6_al
timestamp 1731220307
transform 1 0 288 0 1 332
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_54_6_anx
timestamp 1731220307
transform 1 0 368 0 1 344
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_53_6_al
timestamp 1731220307
transform 1 0 272 0 1 560
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_53_6_anx
timestamp 1731220307
transform 1 0 200 0 1 572
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_52_6_al
timestamp 1731220307
transform 1 0 192 0 -1 944
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_52_6_anx
timestamp 1731220307
transform 1 0 272 0 -1 932
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_51_6_al
timestamp 1731220307
transform 1 0 576 0 -1 1144
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_51_6_anx
timestamp 1731220307
transform 1 0 768 0 1 1164
box 4 6 36 64
use _0_0std_0_0cells_0_0LATCHINV  i_alatch_50_6_al
timestamp 1731220307
transform 1 0 736 0 -1 1340
box 8 4 70 72
use _0_0std_0_0cells_0_0NOR2X2  i_alatch_50_6_anx
timestamp 1731220307
transform 1 0 760 0 1 1360
box 4 6 36 64
use _0_0std_0_0cells_0_0INVX1  src_ar_ai
timestamp 1731220307
transform 1 0 944 0 -1 928
box 8 7 28 34
use _0_0std_0_0cells_0_0OR2X1  src_ar_an
timestamp 1731220307
transform 1 0 976 0 -1 928
box 4 4 48 48
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_57_6
timestamp 1731220307
transform 1 0 1432 0 1 348
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_56_6
timestamp 1731220307
transform 1 0 1280 0 -1 308
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_55_6
timestamp 1731220307
transform 1 0 912 0 1 188
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_54_6
timestamp 1731220307
transform 1 0 712 0 -1 732
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_53_6
timestamp 1731220307
transform 1 0 944 0 1 776
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_52_6
timestamp 1731220307
transform 1 0 672 0 -1 928
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_51_6
timestamp 1731220307
transform 1 0 792 0 -1 1128
box 8 6 28 37
use _0_0std_0_0cells_0_0TIELOX1  src_atlo_50_6
timestamp 1731220307
transform 1 0 992 0 -1 1128
box 8 6 28 37
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_55_6
timestamp 1731220307
transform 1 0 1448 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_54_6
timestamp 1731220307
transform 1 0 1416 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_53_6
timestamp 1731220307
transform 1 0 1368 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_52_6
timestamp 1731220307
transform 1 0 1336 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_51_6
timestamp 1731220307
transform 1 0 1400 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ad_ainvs_50_6
timestamp 1731220307
transform 1 0 1416 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ar0_ai
timestamp 1731220307
transform 1 0 1488 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0NOR2X1  c__copy_ar0_an
timestamp 1731220307
transform 1 0 1448 0 -1 1324
box 4 6 36 48
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_544_6
timestamp 1731220307
transform 1 0 1248 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_543_6
timestamp 1731220307
transform 1 0 1432 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_542_6
timestamp 1731220307
transform 1 0 1472 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_541_6
timestamp 1731220307
transform 1 0 1480 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_540_6
timestamp 1731220307
transform 1 0 1584 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_539_6
timestamp 1731220307
transform 1 0 1648 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_538_6
timestamp 1731220307
transform 1 0 1616 0 -1 1128
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_537_6
timestamp 1731220307
transform 1 0 1584 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_536_6
timestamp 1731220307
transform 1 0 1616 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_535_6
timestamp 1731220307
transform 1 0 1648 0 1 1168
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_534_6
timestamp 1731220307
transform 1 0 1648 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_533_6
timestamp 1731220307
transform 1 0 1616 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_532_6
timestamp 1731220307
transform 1 0 1584 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_531_6
timestamp 1731220307
transform 1 0 1552 0 -1 1324
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_530_6
timestamp 1731220307
transform 1 0 1648 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_529_6
timestamp 1731220307
transform 1 0 1616 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_528_6
timestamp 1731220307
transform 1 0 1576 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_527_6
timestamp 1731220307
transform 1 0 1552 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_526_6
timestamp 1731220307
transform 1 0 1584 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_525_6
timestamp 1731220307
transform 1 0 1648 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_524_6
timestamp 1731220307
transform 1 0 1616 0 -1 1480
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_523_6
timestamp 1731220307
transform 1 0 1592 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_522_6
timestamp 1731220307
transform 1 0 1648 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_521_6
timestamp 1731220307
transform 1 0 1648 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_520_6
timestamp 1731220307
transform 1 0 1600 0 -1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_519_6
timestamp 1731220307
transform 1 0 1560 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_518_6
timestamp 1731220307
transform 1 0 1648 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_517_6
timestamp 1731220307
transform 1 0 1648 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_516_6
timestamp 1731220307
transform 1 0 1552 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_515_6
timestamp 1731220307
transform 1 0 1432 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_514_6
timestamp 1731220307
transform 1 0 1648 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_513_6
timestamp 1731220307
transform 1 0 1616 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_512_6
timestamp 1731220307
transform 1 0 1560 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_511_6
timestamp 1731220307
transform 1 0 1512 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_510_6
timestamp 1731220307
transform 1 0 1456 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_59_6
timestamp 1731220307
transform 1 0 1400 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_58_6
timestamp 1731220307
transform 1 0 1328 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_57_6
timestamp 1731220307
transform 1 0 1248 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_56_6
timestamp 1731220307
transform 1 0 1152 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_55_6
timestamp 1731220307
transform 1 0 1176 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_54_6
timestamp 1731220307
transform 1 0 1312 0 -1 1668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_53_6
timestamp 1731220307
transform 1 0 1352 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_52_6
timestamp 1731220307
transform 1 0 1456 0 1 1580
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_51_6
timestamp 1731220307
transform 1 0 1432 0 1 1500
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  c__copy_ap_ainvs_50_6
timestamp 1731220307
transform 1 0 1408 0 1 1364
box 8 7 28 34
use _0_0std_0_0cells_0_0AND2X1  c__copy_ap_aand
timestamp 1731220307
transform 1 0 1280 0 1 1156
box 8 4 52 52
use _0_0cell_0_0ginvx0  c__copy_ac_acx1
timestamp 1731220307
transform 1 0 1384 0 -1 1324
box 8 6 28 32
use _0_0cell_0_0gcelem2x0  c__copy_ac_acx0
timestamp 1731220307
transform 1 0 1296 0 -1 1340
box 8 4 84 60
use _0_0std_0_0cells_0_0OR2X1  c__copy_ar2_an
timestamp 1731220307
transform 1 0 1152 0 -1 1324
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  c__copy_ar1_an
timestamp 1731220307
transform 1 0 1192 0 1 1168
box 4 4 48 48
use _0_0cell_0_0gcelem2x0  c__copy_ac__ra_acx0
timestamp 1731220307
transform 1 0 1208 0 -1 1340
box 8 4 84 60
use _0_0std_0_0cells_0_0LATCH  c__copy_alatch_50_6
timestamp 1731220307
transform 1 0 1312 0 -1 1140
box 8 5 100 68
<< labels >>
rlabel m1 s 638 1796 642 1800 6 L.d[0]
port 0 nsew signal input
rlabel m1 s 80 1666 84 1670 6 L.d[1]
port 1 nsew signal input
rlabel m1 s 80 1398 84 1402 6 L.d[2]
port 2 nsew signal input
rlabel m1 s 80 866 84 870 6 L.d[3]
port 3 nsew signal input
rlabel m1 s 80 470 84 474 6 L.d[4]
port 4 nsew signal input
rlabel m1 s 80 602 84 606 6 L.d[5]
port 5 nsew signal input
rlabel m1 s 1748 262 1752 266 6 L.d[6]
port 6 nsew signal input
rlabel m1 s 1748 454 1752 458 6 L.d[7]
port 7 nsew signal input
rlabel m1 s 1748 1222 1752 1226 6 L.r
port 8 nsew signal input
rlabel m1 s 1190 1796 1194 1800 6 L.a
port 9 nsew signal tristate
rlabel m1 s 1748 646 1752 650 6 C.d[0]
port 10 nsew signal input
rlabel m1 s 1748 838 1752 842 6 C.r
port 11 nsew signal input
rlabel m1 s 1748 1030 1752 1034 6 C.a
port 12 nsew signal tristate
rlabel m1 s 80 1534 84 1538 6 R.d[0]
port 13 nsew signal tristate
rlabel m1 s 80 1266 84 1270 6 R.d[1]
port 14 nsew signal tristate
rlabel m1 s 80 1002 84 1006 6 R.d[2]
port 15 nsew signal tristate
rlabel m1 s 80 734 84 738 6 R.d[3]
port 16 nsew signal tristate
rlabel m1 s 80 334 84 338 6 R.d[4]
port 17 nsew signal tristate
rlabel m1 s 80 202 84 206 6 R.d[5]
port 18 nsew signal tristate
rlabel m1 s 1190 72 1194 76 6 R.d[6]
port 19 nsew signal tristate
rlabel m1 s 638 72 642 76 6 R.d[7]
port 20 nsew signal tristate
rlabel m1 s 1748 1414 1752 1418 6 R.r
port 21 nsew signal tristate
rlabel m1 s 1748 1606 1752 1610 6 R.a
port 22 nsew signal input
rlabel m1 s 80 1134 84 1138 6 Reset
port 23 nsew signal input
<< end >>
