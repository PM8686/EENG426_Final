magic
tech sky130l
timestamp 1728952526
<< ndiffusion >>
rect -5 28 8 29
rect -5 25 -1 28
rect 2 25 8 28
rect -5 23 8 25
rect 11 27 17 29
rect 11 24 12 27
rect 15 24 17 27
rect 11 23 17 24
rect 20 28 45 29
rect 20 25 25 28
rect 28 25 45 28
rect 20 23 45 25
rect 49 27 58 29
rect 49 24 52 27
rect 55 24 58 27
rect 49 23 58 24
<< ndc >>
rect -1 25 2 28
rect 12 24 15 27
rect 25 25 28 28
rect 52 24 55 27
<< ntransistor >>
rect 8 23 11 29
rect 17 23 20 29
rect 45 23 49 29
<< pdiffusion >>
rect -5 14 8 16
rect -5 11 2 14
rect 5 11 8 14
rect -5 10 8 11
rect 11 10 17 16
rect 20 14 45 16
rect 20 11 33 14
rect 36 11 45 14
rect 20 10 45 11
rect 49 14 58 16
rect 49 11 52 14
rect 55 11 58 14
rect 49 10 58 11
<< pdc >>
rect 2 11 5 14
rect 33 11 36 14
rect 52 11 55 14
<< ptransistor >>
rect 8 10 11 16
rect 17 10 20 16
rect 45 10 49 16
<< polysilicon >>
rect 7 36 12 37
rect 7 33 8 36
rect 11 33 12 36
rect 7 32 12 33
rect 16 36 21 37
rect 16 33 17 36
rect 20 33 21 36
rect 16 32 21 33
rect 8 29 11 32
rect 17 29 20 32
rect 45 29 49 36
rect 8 16 11 23
rect 17 16 20 23
rect 45 16 49 23
rect 8 8 11 10
rect 17 7 20 10
rect 45 8 49 10
rect 44 6 49 8
rect 44 3 45 6
rect 48 3 49 6
rect 44 2 49 3
<< pc >>
rect 8 33 11 36
rect 17 33 20 36
rect 45 3 48 6
<< m1 >>
rect -2 41 -1 44
rect 2 41 3 44
rect -2 28 3 41
rect 24 41 25 44
rect 28 41 29 44
rect 7 36 12 37
rect 7 33 8 36
rect 11 33 12 36
rect 7 32 12 33
rect 16 36 21 37
rect 16 33 17 36
rect 20 33 21 36
rect 16 32 21 33
rect 24 28 29 41
rect -2 25 -1 28
rect 2 25 3 28
rect -2 23 3 25
rect 11 27 16 28
rect 11 24 12 27
rect 15 24 16 27
rect 24 25 25 28
rect 28 25 29 28
rect 24 24 29 25
rect 11 23 16 24
rect 1 14 6 15
rect 1 11 2 14
rect 5 11 6 14
rect 1 7 5 11
rect 13 8 16 23
rect 32 14 36 36
rect 52 27 56 28
rect 55 24 56 27
rect 52 14 56 24
rect 32 11 33 14
rect 36 11 37 14
rect 55 11 56 14
rect 1 4 2 7
rect 12 7 16 8
rect 15 4 16 7
rect 44 6 49 8
rect 44 3 45 6
rect 48 3 49 6
rect 52 5 56 11
rect 44 2 49 3
<< m2c >>
rect -1 41 2 44
rect 25 41 28 44
rect 2 4 5 7
rect 12 4 15 7
rect 45 3 48 6
<< m2 >>
rect -2 44 29 45
rect -2 41 -1 44
rect 2 41 25 44
rect 28 41 29 44
rect -2 40 29 41
rect 1 7 49 8
rect 1 4 2 7
rect 5 4 12 7
rect 15 6 49 7
rect 15 4 45 6
rect 1 3 45 4
rect 48 3 49 6
rect 44 2 49 3
<< labels >>
rlabel m1 s 8 32 12 36 6 A
port 1 nsew signal input
rlabel m1 s 16 32 20 36 6 B
port 2 nsew signal input
rlabel m1 32 32 36 36 1 Vdd
rlabel m1 24 32 28 36 1 GND
rlabel m1 52 5 56 9 8 Y
<< properties >>
string LEFsite CoreSite
string LEFclass CORE
string FIXED_BBOX 0 0 40 40
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
