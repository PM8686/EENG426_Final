magic
tech sky130l
timestamp 1729031399
<< ndiffusion >>
rect 8 10 13 16
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 15 20 16
rect 15 12 16 15
rect 19 12 20 15
rect 15 6 20 12
rect 22 10 27 16
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
<< ndc >>
rect 9 7 12 10
rect 16 12 19 15
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
<< pdiffusion >>
rect 8 52 13 53
rect 8 49 9 52
rect 12 49 13 52
rect 8 23 13 49
rect 15 23 20 53
rect 22 27 27 53
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
<< pdc >>
rect 9 49 12 52
rect 23 24 26 27
<< ptransistor >>
rect 13 23 15 53
rect 20 23 22 53
<< polysilicon >>
rect 13 64 20 65
rect 13 61 16 64
rect 19 61 20 64
rect 13 60 20 61
rect 24 61 29 62
rect 13 53 15 60
rect 24 58 25 61
rect 28 58 29 61
rect 24 56 29 58
rect 20 54 29 56
rect 20 53 22 54
rect 13 16 15 23
rect 20 16 22 23
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 16 61 19 64
rect 25 58 28 61
<< m1 >>
rect 16 64 20 65
rect 19 61 20 64
rect 8 59 12 60
rect 11 56 12 59
rect 16 56 20 61
rect 24 61 28 62
rect 24 58 25 61
rect 24 56 28 58
rect 8 52 12 56
rect 8 49 9 52
rect 8 48 12 49
rect 16 24 23 27
rect 26 24 27 27
rect 16 15 20 24
rect 19 12 20 15
rect 8 10 12 11
rect 8 7 9 10
rect 8 4 12 7
rect 16 4 20 12
rect 23 10 26 11
rect 23 6 26 7
<< m2c >>
rect 8 56 11 59
rect 9 7 12 10
rect 23 7 26 10
<< m2 >>
rect 7 59 12 60
rect 7 56 8 59
rect 11 56 12 59
rect 7 55 12 56
rect 8 10 27 11
rect 8 7 9 10
rect 12 7 23 10
rect 26 7 27 10
rect 8 6 27 7
<< labels >>
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 24 23 24 3 Y
rlabel polysilicon 21 17 21 17 3 B
rlabel polysilicon 21 22 21 22 3 B
rlabel ndiffusion 16 7 16 7 3 Y
rlabel polysilicon 14 17 14 17 3 A
rlabel polysilicon 14 22 14 22 3 A
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m1 9 5 9 5 3 GND
rlabel m2 9 7 9 7 3 GND
rlabel m1 17 5 17 5 3 Y
rlabel m1 17 57 17 57 3 A
rlabel m1 25 57 25 57 3 B
rlabel m2c 9 57 9 57 3 Vdd
<< end >>
