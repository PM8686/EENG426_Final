magic
tech sky130l
timestamp 1729225234
<< ndiffusion >>
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 6 13 8
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
rect 22 11 27 12
rect 22 8 23 11
rect 26 8 27 11
rect 22 6 27 8
rect 29 11 44 12
rect 29 8 40 11
rect 43 8 44 11
rect 29 6 44 8
<< ndc >>
rect 9 8 12 11
rect 16 7 19 10
rect 23 8 26 11
rect 40 8 43 11
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
rect 27 6 29 12
<< pdiffusion >>
rect 8 27 13 34
rect 8 24 9 27
rect 12 24 13 27
rect 8 19 13 24
rect 15 19 20 34
rect 22 27 26 34
rect 22 25 27 27
rect 22 22 23 25
rect 26 22 27 25
rect 22 19 27 22
rect 29 25 34 27
rect 29 23 44 25
rect 29 20 40 23
rect 43 20 44 23
rect 29 19 44 20
<< pdc >>
rect 9 24 12 27
rect 23 22 26 25
rect 40 20 43 23
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
rect 27 19 29 27
<< polysilicon >>
rect 10 41 15 42
rect 10 38 11 41
rect 14 38 15 41
rect 10 37 15 38
rect 18 41 23 42
rect 18 38 19 41
rect 22 38 23 41
rect 18 37 23 38
rect 13 34 15 37
rect 20 34 22 37
rect 27 27 29 29
rect 13 12 15 19
rect 20 12 22 19
rect 27 12 29 19
rect 13 4 15 6
rect 20 4 22 6
rect 27 -4 29 6
rect 25 -5 30 -4
rect 25 -8 26 -5
rect 29 -8 30 -5
rect 25 -9 30 -8
<< pc >>
rect 11 38 14 41
rect 19 38 22 41
rect 26 -8 29 -5
<< m1 >>
rect 10 41 15 42
rect 10 38 11 41
rect 14 38 15 41
rect 10 37 15 38
rect 18 41 22 42
rect 18 38 19 41
rect 18 37 22 38
rect 25 36 29 40
rect 32 36 36 40
rect 25 32 28 36
rect 23 29 28 32
rect 9 27 12 28
rect 9 19 12 24
rect 23 25 26 29
rect 23 21 26 22
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 7 13 8
rect 16 10 19 16
rect 22 11 27 12
rect 22 8 23 11
rect 26 8 27 11
rect 22 7 27 8
rect 33 11 36 36
rect 33 7 36 8
rect 40 23 43 24
rect 40 11 43 20
rect 8 3 12 4
rect 11 0 12 3
rect 16 -5 19 7
rect 40 3 43 8
rect 25 -5 30 -4
rect 25 -8 26 -5
rect 29 -8 30 -5
rect 25 -9 30 -8
<< m2c >>
rect 9 16 12 19
rect 16 16 19 19
rect 9 8 12 11
rect 23 8 26 11
rect 33 8 36 11
rect 8 0 11 3
rect 40 0 43 3
rect 16 -8 19 -5
rect 26 -8 29 -5
<< m2 >>
rect 8 19 20 20
rect 8 16 9 19
rect 12 16 16 19
rect 19 16 20 19
rect 8 15 20 16
rect 8 11 13 12
rect 8 8 9 11
rect 12 10 13 11
rect 22 11 27 12
rect 22 10 23 11
rect 12 8 23 10
rect 26 10 27 11
rect 32 11 37 12
rect 32 10 33 11
rect 26 8 33 10
rect 36 8 37 11
rect 8 7 37 8
rect 7 3 12 4
rect 39 3 44 4
rect 7 0 8 3
rect 11 0 40 3
rect 43 0 44 3
rect 7 -1 12 0
rect 39 -1 44 0
rect 15 -5 30 -4
rect 15 -8 16 -5
rect 19 -8 26 -5
rect 29 -8 30 -5
rect 15 -9 30 -8
<< labels >>
rlabel pdiffusion 30 20 30 20 3 Y
rlabel ndiffusion 30 7 30 7 3 Y
rlabel polysilicon 28 13 28 13 3 _Y
rlabel polysilicon 28 18 28 18 3 _Y
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 20 23 20 3 Vdd
rlabel polysilicon 21 13 21 13 3 A
rlabel polysilicon 21 18 21 18 3 A
rlabel ndiffusion 16 7 16 7 3 _Y
rlabel polysilicon 14 13 14 13 3 B
rlabel polysilicon 14 18 14 18 3 B
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 _Y
rlabel m1 33 37 33 37 3 GND
port 1 e
rlabel m1 26 37 27 38 5 Vdd
rlabel m2c 9 1 10 2 2 Y
rlabel m1 34 37 35 38 5 GND
rlabel pc 12 39 13 40 4 B
rlabel pc 20 39 21 40 5 A
<< end >>
