magic
tech sky130l
timestamp 1731220379
<< m2 >>
rect 158 2650 164 2651
rect 158 2646 159 2650
rect 163 2646 164 2650
rect 158 2645 164 2646
rect 214 2650 220 2651
rect 214 2646 215 2650
rect 219 2646 220 2650
rect 214 2645 220 2646
rect 270 2650 276 2651
rect 270 2646 271 2650
rect 275 2646 276 2650
rect 270 2645 276 2646
rect 326 2650 332 2651
rect 326 2646 327 2650
rect 331 2646 332 2650
rect 326 2645 332 2646
rect 110 2641 116 2642
rect 110 2637 111 2641
rect 115 2637 116 2641
rect 110 2636 116 2637
rect 1326 2641 1332 2642
rect 1326 2637 1327 2641
rect 1331 2637 1332 2641
rect 1326 2636 1332 2637
rect 110 2624 116 2625
rect 1326 2624 1332 2625
rect 110 2620 111 2624
rect 115 2620 116 2624
rect 110 2619 116 2620
rect 142 2623 148 2624
rect 142 2619 143 2623
rect 147 2619 148 2623
rect 142 2618 148 2619
rect 198 2623 204 2624
rect 198 2619 199 2623
rect 203 2619 204 2623
rect 198 2618 204 2619
rect 254 2623 260 2624
rect 254 2619 255 2623
rect 259 2619 260 2623
rect 254 2618 260 2619
rect 310 2623 316 2624
rect 310 2619 311 2623
rect 315 2619 316 2623
rect 1326 2620 1327 2624
rect 1331 2620 1332 2624
rect 1326 2619 1332 2620
rect 310 2618 316 2619
rect 1414 2598 1420 2599
rect 1414 2594 1415 2598
rect 1419 2594 1420 2598
rect 1414 2593 1420 2594
rect 1470 2598 1476 2599
rect 1470 2594 1471 2598
rect 1475 2594 1476 2598
rect 1470 2593 1476 2594
rect 1526 2598 1532 2599
rect 1526 2594 1527 2598
rect 1531 2594 1532 2598
rect 1526 2593 1532 2594
rect 1582 2598 1588 2599
rect 1582 2594 1583 2598
rect 1587 2594 1588 2598
rect 1582 2593 1588 2594
rect 1638 2598 1644 2599
rect 1638 2594 1639 2598
rect 1643 2594 1644 2598
rect 1638 2593 1644 2594
rect 1694 2598 1700 2599
rect 1694 2594 1695 2598
rect 1699 2594 1700 2598
rect 1694 2593 1700 2594
rect 142 2589 148 2590
rect 110 2588 116 2589
rect 110 2584 111 2588
rect 115 2584 116 2588
rect 142 2585 143 2589
rect 147 2585 148 2589
rect 142 2584 148 2585
rect 198 2589 204 2590
rect 198 2585 199 2589
rect 203 2585 204 2589
rect 198 2584 204 2585
rect 262 2589 268 2590
rect 262 2585 263 2589
rect 267 2585 268 2589
rect 262 2584 268 2585
rect 342 2589 348 2590
rect 342 2585 343 2589
rect 347 2585 348 2589
rect 342 2584 348 2585
rect 430 2589 436 2590
rect 430 2585 431 2589
rect 435 2585 436 2589
rect 430 2584 436 2585
rect 518 2589 524 2590
rect 518 2585 519 2589
rect 523 2585 524 2589
rect 518 2584 524 2585
rect 606 2589 612 2590
rect 606 2585 607 2589
rect 611 2585 612 2589
rect 606 2584 612 2585
rect 686 2589 692 2590
rect 686 2585 687 2589
rect 691 2585 692 2589
rect 686 2584 692 2585
rect 766 2589 772 2590
rect 766 2585 767 2589
rect 771 2585 772 2589
rect 766 2584 772 2585
rect 838 2589 844 2590
rect 838 2585 839 2589
rect 843 2585 844 2589
rect 838 2584 844 2585
rect 902 2589 908 2590
rect 902 2585 903 2589
rect 907 2585 908 2589
rect 902 2584 908 2585
rect 966 2589 972 2590
rect 966 2585 967 2589
rect 971 2585 972 2589
rect 966 2584 972 2585
rect 1030 2589 1036 2590
rect 1030 2585 1031 2589
rect 1035 2585 1036 2589
rect 1030 2584 1036 2585
rect 1094 2589 1100 2590
rect 1094 2585 1095 2589
rect 1099 2585 1100 2589
rect 1094 2584 1100 2585
rect 1158 2589 1164 2590
rect 1158 2585 1159 2589
rect 1163 2585 1164 2589
rect 1158 2584 1164 2585
rect 1214 2589 1220 2590
rect 1214 2585 1215 2589
rect 1219 2585 1220 2589
rect 1214 2584 1220 2585
rect 1270 2589 1276 2590
rect 1366 2589 1372 2590
rect 1270 2585 1271 2589
rect 1275 2585 1276 2589
rect 1270 2584 1276 2585
rect 1326 2588 1332 2589
rect 1326 2584 1327 2588
rect 1331 2584 1332 2588
rect 1366 2585 1367 2589
rect 1371 2585 1372 2589
rect 1366 2584 1372 2585
rect 2582 2589 2588 2590
rect 2582 2585 2583 2589
rect 2587 2585 2588 2589
rect 2582 2584 2588 2585
rect 110 2583 116 2584
rect 1326 2583 1332 2584
rect 1366 2572 1372 2573
rect 2582 2572 2588 2573
rect 110 2571 116 2572
rect 110 2567 111 2571
rect 115 2567 116 2571
rect 110 2566 116 2567
rect 1326 2571 1332 2572
rect 1326 2567 1327 2571
rect 1331 2567 1332 2571
rect 1366 2568 1367 2572
rect 1371 2568 1372 2572
rect 1366 2567 1372 2568
rect 1398 2571 1404 2572
rect 1398 2567 1399 2571
rect 1403 2567 1404 2571
rect 1326 2566 1332 2567
rect 1398 2566 1404 2567
rect 1454 2571 1460 2572
rect 1454 2567 1455 2571
rect 1459 2567 1460 2571
rect 1454 2566 1460 2567
rect 1510 2571 1516 2572
rect 1510 2567 1511 2571
rect 1515 2567 1516 2571
rect 1510 2566 1516 2567
rect 1566 2571 1572 2572
rect 1566 2567 1567 2571
rect 1571 2567 1572 2571
rect 1566 2566 1572 2567
rect 1622 2571 1628 2572
rect 1622 2567 1623 2571
rect 1627 2567 1628 2571
rect 1622 2566 1628 2567
rect 1678 2571 1684 2572
rect 1678 2567 1679 2571
rect 1683 2567 1684 2571
rect 2582 2568 2583 2572
rect 2587 2568 2588 2572
rect 2582 2567 2588 2568
rect 1678 2566 1684 2567
rect 158 2562 164 2563
rect 158 2558 159 2562
rect 163 2558 164 2562
rect 158 2557 164 2558
rect 214 2562 220 2563
rect 214 2558 215 2562
rect 219 2558 220 2562
rect 214 2557 220 2558
rect 278 2562 284 2563
rect 278 2558 279 2562
rect 283 2558 284 2562
rect 278 2557 284 2558
rect 358 2562 364 2563
rect 358 2558 359 2562
rect 363 2558 364 2562
rect 358 2557 364 2558
rect 446 2562 452 2563
rect 446 2558 447 2562
rect 451 2558 452 2562
rect 446 2557 452 2558
rect 534 2562 540 2563
rect 534 2558 535 2562
rect 539 2558 540 2562
rect 534 2557 540 2558
rect 622 2562 628 2563
rect 622 2558 623 2562
rect 627 2558 628 2562
rect 622 2557 628 2558
rect 702 2562 708 2563
rect 702 2558 703 2562
rect 707 2558 708 2562
rect 702 2557 708 2558
rect 782 2562 788 2563
rect 782 2558 783 2562
rect 787 2558 788 2562
rect 782 2557 788 2558
rect 854 2562 860 2563
rect 854 2558 855 2562
rect 859 2558 860 2562
rect 854 2557 860 2558
rect 918 2562 924 2563
rect 918 2558 919 2562
rect 923 2558 924 2562
rect 918 2557 924 2558
rect 982 2562 988 2563
rect 982 2558 983 2562
rect 987 2558 988 2562
rect 982 2557 988 2558
rect 1046 2562 1052 2563
rect 1046 2558 1047 2562
rect 1051 2558 1052 2562
rect 1046 2557 1052 2558
rect 1110 2562 1116 2563
rect 1110 2558 1111 2562
rect 1115 2558 1116 2562
rect 1110 2557 1116 2558
rect 1174 2562 1180 2563
rect 1174 2558 1175 2562
rect 1179 2558 1180 2562
rect 1174 2557 1180 2558
rect 1230 2562 1236 2563
rect 1230 2558 1231 2562
rect 1235 2558 1236 2562
rect 1230 2557 1236 2558
rect 1286 2562 1292 2563
rect 1286 2558 1287 2562
rect 1291 2558 1292 2562
rect 1286 2557 1292 2558
rect 1398 2537 1404 2538
rect 1366 2536 1372 2537
rect 1366 2532 1367 2536
rect 1371 2532 1372 2536
rect 1398 2533 1399 2537
rect 1403 2533 1404 2537
rect 1398 2532 1404 2533
rect 1454 2537 1460 2538
rect 1454 2533 1455 2537
rect 1459 2533 1460 2537
rect 1454 2532 1460 2533
rect 1510 2537 1516 2538
rect 1510 2533 1511 2537
rect 1515 2533 1516 2537
rect 1510 2532 1516 2533
rect 1566 2537 1572 2538
rect 1566 2533 1567 2537
rect 1571 2533 1572 2537
rect 1566 2532 1572 2533
rect 1622 2537 1628 2538
rect 1622 2533 1623 2537
rect 1627 2533 1628 2537
rect 1622 2532 1628 2533
rect 1678 2537 1684 2538
rect 1678 2533 1679 2537
rect 1683 2533 1684 2537
rect 1678 2532 1684 2533
rect 1734 2537 1740 2538
rect 1734 2533 1735 2537
rect 1739 2533 1740 2537
rect 1734 2532 1740 2533
rect 2582 2536 2588 2537
rect 2582 2532 2583 2536
rect 2587 2532 2588 2536
rect 1366 2531 1372 2532
rect 2582 2531 2588 2532
rect 158 2526 164 2527
rect 158 2522 159 2526
rect 163 2522 164 2526
rect 158 2521 164 2522
rect 214 2526 220 2527
rect 214 2522 215 2526
rect 219 2522 220 2526
rect 214 2521 220 2522
rect 318 2526 324 2527
rect 318 2522 319 2526
rect 323 2522 324 2526
rect 318 2521 324 2522
rect 430 2526 436 2527
rect 430 2522 431 2526
rect 435 2522 436 2526
rect 430 2521 436 2522
rect 550 2526 556 2527
rect 550 2522 551 2526
rect 555 2522 556 2526
rect 550 2521 556 2522
rect 670 2526 676 2527
rect 670 2522 671 2526
rect 675 2522 676 2526
rect 670 2521 676 2522
rect 790 2526 796 2527
rect 790 2522 791 2526
rect 795 2522 796 2526
rect 790 2521 796 2522
rect 902 2526 908 2527
rect 902 2522 903 2526
rect 907 2522 908 2526
rect 902 2521 908 2522
rect 1006 2526 1012 2527
rect 1006 2522 1007 2526
rect 1011 2522 1012 2526
rect 1006 2521 1012 2522
rect 1102 2526 1108 2527
rect 1102 2522 1103 2526
rect 1107 2522 1108 2526
rect 1102 2521 1108 2522
rect 1206 2526 1212 2527
rect 1206 2522 1207 2526
rect 1211 2522 1212 2526
rect 1206 2521 1212 2522
rect 1286 2526 1292 2527
rect 1286 2522 1287 2526
rect 1291 2522 1292 2526
rect 1286 2521 1292 2522
rect 1366 2519 1372 2520
rect 110 2517 116 2518
rect 110 2513 111 2517
rect 115 2513 116 2517
rect 110 2512 116 2513
rect 1326 2517 1332 2518
rect 1326 2513 1327 2517
rect 1331 2513 1332 2517
rect 1366 2515 1367 2519
rect 1371 2515 1372 2519
rect 1366 2514 1372 2515
rect 2582 2519 2588 2520
rect 2582 2515 2583 2519
rect 2587 2515 2588 2519
rect 2582 2514 2588 2515
rect 1326 2512 1332 2513
rect 1414 2510 1420 2511
rect 1414 2506 1415 2510
rect 1419 2506 1420 2510
rect 1414 2505 1420 2506
rect 1470 2510 1476 2511
rect 1470 2506 1471 2510
rect 1475 2506 1476 2510
rect 1470 2505 1476 2506
rect 1526 2510 1532 2511
rect 1526 2506 1527 2510
rect 1531 2506 1532 2510
rect 1526 2505 1532 2506
rect 1582 2510 1588 2511
rect 1582 2506 1583 2510
rect 1587 2506 1588 2510
rect 1582 2505 1588 2506
rect 1638 2510 1644 2511
rect 1638 2506 1639 2510
rect 1643 2506 1644 2510
rect 1638 2505 1644 2506
rect 1694 2510 1700 2511
rect 1694 2506 1695 2510
rect 1699 2506 1700 2510
rect 1694 2505 1700 2506
rect 1750 2510 1756 2511
rect 1750 2506 1751 2510
rect 1755 2506 1756 2510
rect 1750 2505 1756 2506
rect 110 2500 116 2501
rect 1326 2500 1332 2501
rect 110 2496 111 2500
rect 115 2496 116 2500
rect 110 2495 116 2496
rect 142 2499 148 2500
rect 142 2495 143 2499
rect 147 2495 148 2499
rect 142 2494 148 2495
rect 198 2499 204 2500
rect 198 2495 199 2499
rect 203 2495 204 2499
rect 198 2494 204 2495
rect 302 2499 308 2500
rect 302 2495 303 2499
rect 307 2495 308 2499
rect 302 2494 308 2495
rect 414 2499 420 2500
rect 414 2495 415 2499
rect 419 2495 420 2499
rect 414 2494 420 2495
rect 534 2499 540 2500
rect 534 2495 535 2499
rect 539 2495 540 2499
rect 534 2494 540 2495
rect 654 2499 660 2500
rect 654 2495 655 2499
rect 659 2495 660 2499
rect 654 2494 660 2495
rect 774 2499 780 2500
rect 774 2495 775 2499
rect 779 2495 780 2499
rect 774 2494 780 2495
rect 886 2499 892 2500
rect 886 2495 887 2499
rect 891 2495 892 2499
rect 886 2494 892 2495
rect 990 2499 996 2500
rect 990 2495 991 2499
rect 995 2495 996 2499
rect 990 2494 996 2495
rect 1086 2499 1092 2500
rect 1086 2495 1087 2499
rect 1091 2495 1092 2499
rect 1086 2494 1092 2495
rect 1190 2499 1196 2500
rect 1190 2495 1191 2499
rect 1195 2495 1196 2499
rect 1190 2494 1196 2495
rect 1270 2499 1276 2500
rect 1270 2495 1271 2499
rect 1275 2495 1276 2499
rect 1326 2496 1327 2500
rect 1331 2496 1332 2500
rect 1326 2495 1332 2496
rect 1270 2494 1276 2495
rect 1470 2482 1476 2483
rect 1470 2478 1471 2482
rect 1475 2478 1476 2482
rect 1470 2477 1476 2478
rect 1526 2482 1532 2483
rect 1526 2478 1527 2482
rect 1531 2478 1532 2482
rect 1526 2477 1532 2478
rect 1582 2482 1588 2483
rect 1582 2478 1583 2482
rect 1587 2478 1588 2482
rect 1582 2477 1588 2478
rect 1638 2482 1644 2483
rect 1638 2478 1639 2482
rect 1643 2478 1644 2482
rect 1638 2477 1644 2478
rect 1694 2482 1700 2483
rect 1694 2478 1695 2482
rect 1699 2478 1700 2482
rect 1694 2477 1700 2478
rect 1750 2482 1756 2483
rect 1750 2478 1751 2482
rect 1755 2478 1756 2482
rect 1750 2477 1756 2478
rect 1366 2473 1372 2474
rect 1366 2469 1367 2473
rect 1371 2469 1372 2473
rect 1366 2468 1372 2469
rect 2582 2473 2588 2474
rect 2582 2469 2583 2473
rect 2587 2469 2588 2473
rect 2582 2468 2588 2469
rect 142 2457 148 2458
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 142 2453 143 2457
rect 147 2453 148 2457
rect 142 2452 148 2453
rect 198 2457 204 2458
rect 198 2453 199 2457
rect 203 2453 204 2457
rect 198 2452 204 2453
rect 294 2457 300 2458
rect 294 2453 295 2457
rect 299 2453 300 2457
rect 294 2452 300 2453
rect 406 2457 412 2458
rect 406 2453 407 2457
rect 411 2453 412 2457
rect 406 2452 412 2453
rect 518 2457 524 2458
rect 518 2453 519 2457
rect 523 2453 524 2457
rect 518 2452 524 2453
rect 638 2457 644 2458
rect 638 2453 639 2457
rect 643 2453 644 2457
rect 638 2452 644 2453
rect 750 2457 756 2458
rect 750 2453 751 2457
rect 755 2453 756 2457
rect 750 2452 756 2453
rect 854 2457 860 2458
rect 854 2453 855 2457
rect 859 2453 860 2457
rect 854 2452 860 2453
rect 950 2457 956 2458
rect 950 2453 951 2457
rect 955 2453 956 2457
rect 950 2452 956 2453
rect 1046 2457 1052 2458
rect 1046 2453 1047 2457
rect 1051 2453 1052 2457
rect 1046 2452 1052 2453
rect 1142 2457 1148 2458
rect 1142 2453 1143 2457
rect 1147 2453 1148 2457
rect 1142 2452 1148 2453
rect 1238 2457 1244 2458
rect 1238 2453 1239 2457
rect 1243 2453 1244 2457
rect 1238 2452 1244 2453
rect 1326 2456 1332 2457
rect 1326 2452 1327 2456
rect 1331 2452 1332 2456
rect 110 2451 116 2452
rect 1326 2451 1332 2452
rect 1366 2456 1372 2457
rect 2582 2456 2588 2457
rect 1366 2452 1367 2456
rect 1371 2452 1372 2456
rect 1366 2451 1372 2452
rect 1454 2455 1460 2456
rect 1454 2451 1455 2455
rect 1459 2451 1460 2455
rect 1454 2450 1460 2451
rect 1510 2455 1516 2456
rect 1510 2451 1511 2455
rect 1515 2451 1516 2455
rect 1510 2450 1516 2451
rect 1566 2455 1572 2456
rect 1566 2451 1567 2455
rect 1571 2451 1572 2455
rect 1566 2450 1572 2451
rect 1622 2455 1628 2456
rect 1622 2451 1623 2455
rect 1627 2451 1628 2455
rect 1622 2450 1628 2451
rect 1678 2455 1684 2456
rect 1678 2451 1679 2455
rect 1683 2451 1684 2455
rect 1678 2450 1684 2451
rect 1734 2455 1740 2456
rect 1734 2451 1735 2455
rect 1739 2451 1740 2455
rect 2582 2452 2583 2456
rect 2587 2452 2588 2456
rect 2582 2451 2588 2452
rect 1734 2450 1740 2451
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 1326 2439 1332 2440
rect 1326 2435 1327 2439
rect 1331 2435 1332 2439
rect 1326 2434 1332 2435
rect 158 2430 164 2431
rect 158 2426 159 2430
rect 163 2426 164 2430
rect 158 2425 164 2426
rect 214 2430 220 2431
rect 214 2426 215 2430
rect 219 2426 220 2430
rect 214 2425 220 2426
rect 310 2430 316 2431
rect 310 2426 311 2430
rect 315 2426 316 2430
rect 310 2425 316 2426
rect 422 2430 428 2431
rect 422 2426 423 2430
rect 427 2426 428 2430
rect 422 2425 428 2426
rect 534 2430 540 2431
rect 534 2426 535 2430
rect 539 2426 540 2430
rect 534 2425 540 2426
rect 654 2430 660 2431
rect 654 2426 655 2430
rect 659 2426 660 2430
rect 654 2425 660 2426
rect 766 2430 772 2431
rect 766 2426 767 2430
rect 771 2426 772 2430
rect 766 2425 772 2426
rect 870 2430 876 2431
rect 870 2426 871 2430
rect 875 2426 876 2430
rect 870 2425 876 2426
rect 966 2430 972 2431
rect 966 2426 967 2430
rect 971 2426 972 2430
rect 966 2425 972 2426
rect 1062 2430 1068 2431
rect 1062 2426 1063 2430
rect 1067 2426 1068 2430
rect 1062 2425 1068 2426
rect 1158 2430 1164 2431
rect 1158 2426 1159 2430
rect 1163 2426 1164 2430
rect 1158 2425 1164 2426
rect 1254 2430 1260 2431
rect 1254 2426 1255 2430
rect 1259 2426 1260 2430
rect 1254 2425 1260 2426
rect 1478 2413 1484 2414
rect 1366 2412 1372 2413
rect 1366 2408 1367 2412
rect 1371 2408 1372 2412
rect 1478 2409 1479 2413
rect 1483 2409 1484 2413
rect 1478 2408 1484 2409
rect 1534 2413 1540 2414
rect 1534 2409 1535 2413
rect 1539 2409 1540 2413
rect 1534 2408 1540 2409
rect 1590 2413 1596 2414
rect 1590 2409 1591 2413
rect 1595 2409 1596 2413
rect 1590 2408 1596 2409
rect 1646 2413 1652 2414
rect 1646 2409 1647 2413
rect 1651 2409 1652 2413
rect 1646 2408 1652 2409
rect 1702 2413 1708 2414
rect 1702 2409 1703 2413
rect 1707 2409 1708 2413
rect 1702 2408 1708 2409
rect 1758 2413 1764 2414
rect 1758 2409 1759 2413
rect 1763 2409 1764 2413
rect 1758 2408 1764 2409
rect 2582 2412 2588 2413
rect 2582 2408 2583 2412
rect 2587 2408 2588 2412
rect 1366 2407 1372 2408
rect 2582 2407 2588 2408
rect 222 2398 228 2399
rect 222 2394 223 2398
rect 227 2394 228 2398
rect 222 2393 228 2394
rect 286 2398 292 2399
rect 286 2394 287 2398
rect 291 2394 292 2398
rect 286 2393 292 2394
rect 366 2398 372 2399
rect 366 2394 367 2398
rect 371 2394 372 2398
rect 366 2393 372 2394
rect 454 2398 460 2399
rect 454 2394 455 2398
rect 459 2394 460 2398
rect 454 2393 460 2394
rect 542 2398 548 2399
rect 542 2394 543 2398
rect 547 2394 548 2398
rect 542 2393 548 2394
rect 638 2398 644 2399
rect 638 2394 639 2398
rect 643 2394 644 2398
rect 638 2393 644 2394
rect 726 2398 732 2399
rect 726 2394 727 2398
rect 731 2394 732 2398
rect 726 2393 732 2394
rect 814 2398 820 2399
rect 814 2394 815 2398
rect 819 2394 820 2398
rect 814 2393 820 2394
rect 894 2398 900 2399
rect 894 2394 895 2398
rect 899 2394 900 2398
rect 894 2393 900 2394
rect 974 2398 980 2399
rect 974 2394 975 2398
rect 979 2394 980 2398
rect 974 2393 980 2394
rect 1054 2398 1060 2399
rect 1054 2394 1055 2398
rect 1059 2394 1060 2398
rect 1054 2393 1060 2394
rect 1142 2398 1148 2399
rect 1142 2394 1143 2398
rect 1147 2394 1148 2398
rect 1142 2393 1148 2394
rect 1366 2395 1372 2396
rect 1366 2391 1367 2395
rect 1371 2391 1372 2395
rect 1366 2390 1372 2391
rect 2582 2395 2588 2396
rect 2582 2391 2583 2395
rect 2587 2391 2588 2395
rect 2582 2390 2588 2391
rect 110 2389 116 2390
rect 110 2385 111 2389
rect 115 2385 116 2389
rect 110 2384 116 2385
rect 1326 2389 1332 2390
rect 1326 2385 1327 2389
rect 1331 2385 1332 2389
rect 1326 2384 1332 2385
rect 1494 2386 1500 2387
rect 1494 2382 1495 2386
rect 1499 2382 1500 2386
rect 1494 2381 1500 2382
rect 1550 2386 1556 2387
rect 1550 2382 1551 2386
rect 1555 2382 1556 2386
rect 1550 2381 1556 2382
rect 1606 2386 1612 2387
rect 1606 2382 1607 2386
rect 1611 2382 1612 2386
rect 1606 2381 1612 2382
rect 1662 2386 1668 2387
rect 1662 2382 1663 2386
rect 1667 2382 1668 2386
rect 1662 2381 1668 2382
rect 1718 2386 1724 2387
rect 1718 2382 1719 2386
rect 1723 2382 1724 2386
rect 1718 2381 1724 2382
rect 1774 2386 1780 2387
rect 1774 2382 1775 2386
rect 1779 2382 1780 2386
rect 1774 2381 1780 2382
rect 110 2372 116 2373
rect 1326 2372 1332 2373
rect 110 2368 111 2372
rect 115 2368 116 2372
rect 110 2367 116 2368
rect 206 2371 212 2372
rect 206 2367 207 2371
rect 211 2367 212 2371
rect 206 2366 212 2367
rect 270 2371 276 2372
rect 270 2367 271 2371
rect 275 2367 276 2371
rect 270 2366 276 2367
rect 350 2371 356 2372
rect 350 2367 351 2371
rect 355 2367 356 2371
rect 350 2366 356 2367
rect 438 2371 444 2372
rect 438 2367 439 2371
rect 443 2367 444 2371
rect 438 2366 444 2367
rect 526 2371 532 2372
rect 526 2367 527 2371
rect 531 2367 532 2371
rect 526 2366 532 2367
rect 622 2371 628 2372
rect 622 2367 623 2371
rect 627 2367 628 2371
rect 622 2366 628 2367
rect 710 2371 716 2372
rect 710 2367 711 2371
rect 715 2367 716 2371
rect 710 2366 716 2367
rect 798 2371 804 2372
rect 798 2367 799 2371
rect 803 2367 804 2371
rect 798 2366 804 2367
rect 878 2371 884 2372
rect 878 2367 879 2371
rect 883 2367 884 2371
rect 878 2366 884 2367
rect 958 2371 964 2372
rect 958 2367 959 2371
rect 963 2367 964 2371
rect 958 2366 964 2367
rect 1038 2371 1044 2372
rect 1038 2367 1039 2371
rect 1043 2367 1044 2371
rect 1038 2366 1044 2367
rect 1126 2371 1132 2372
rect 1126 2367 1127 2371
rect 1131 2367 1132 2371
rect 1326 2368 1327 2372
rect 1331 2368 1332 2372
rect 1326 2367 1332 2368
rect 1126 2366 1132 2367
rect 1470 2358 1476 2359
rect 1470 2354 1471 2358
rect 1475 2354 1476 2358
rect 1470 2353 1476 2354
rect 1526 2358 1532 2359
rect 1526 2354 1527 2358
rect 1531 2354 1532 2358
rect 1526 2353 1532 2354
rect 1582 2358 1588 2359
rect 1582 2354 1583 2358
rect 1587 2354 1588 2358
rect 1582 2353 1588 2354
rect 1638 2358 1644 2359
rect 1638 2354 1639 2358
rect 1643 2354 1644 2358
rect 1638 2353 1644 2354
rect 1694 2358 1700 2359
rect 1694 2354 1695 2358
rect 1699 2354 1700 2358
rect 1694 2353 1700 2354
rect 1366 2349 1372 2350
rect 1366 2345 1367 2349
rect 1371 2345 1372 2349
rect 1366 2344 1372 2345
rect 2582 2349 2588 2350
rect 2582 2345 2583 2349
rect 2587 2345 2588 2349
rect 2582 2344 2588 2345
rect 1366 2332 1372 2333
rect 2582 2332 2588 2333
rect 326 2329 332 2330
rect 110 2328 116 2329
rect 110 2324 111 2328
rect 115 2324 116 2328
rect 326 2325 327 2329
rect 331 2325 332 2329
rect 326 2324 332 2325
rect 382 2329 388 2330
rect 382 2325 383 2329
rect 387 2325 388 2329
rect 382 2324 388 2325
rect 438 2329 444 2330
rect 438 2325 439 2329
rect 443 2325 444 2329
rect 438 2324 444 2325
rect 502 2329 508 2330
rect 502 2325 503 2329
rect 507 2325 508 2329
rect 502 2324 508 2325
rect 566 2329 572 2330
rect 566 2325 567 2329
rect 571 2325 572 2329
rect 566 2324 572 2325
rect 630 2329 636 2330
rect 630 2325 631 2329
rect 635 2325 636 2329
rect 630 2324 636 2325
rect 694 2329 700 2330
rect 694 2325 695 2329
rect 699 2325 700 2329
rect 694 2324 700 2325
rect 758 2329 764 2330
rect 758 2325 759 2329
rect 763 2325 764 2329
rect 758 2324 764 2325
rect 822 2329 828 2330
rect 822 2325 823 2329
rect 827 2325 828 2329
rect 822 2324 828 2325
rect 886 2329 892 2330
rect 886 2325 887 2329
rect 891 2325 892 2329
rect 886 2324 892 2325
rect 950 2329 956 2330
rect 950 2325 951 2329
rect 955 2325 956 2329
rect 950 2324 956 2325
rect 1014 2329 1020 2330
rect 1014 2325 1015 2329
rect 1019 2325 1020 2329
rect 1014 2324 1020 2325
rect 1326 2328 1332 2329
rect 1326 2324 1327 2328
rect 1331 2324 1332 2328
rect 1366 2328 1367 2332
rect 1371 2328 1372 2332
rect 1366 2327 1372 2328
rect 1454 2331 1460 2332
rect 1454 2327 1455 2331
rect 1459 2327 1460 2331
rect 1454 2326 1460 2327
rect 1510 2331 1516 2332
rect 1510 2327 1511 2331
rect 1515 2327 1516 2331
rect 1510 2326 1516 2327
rect 1566 2331 1572 2332
rect 1566 2327 1567 2331
rect 1571 2327 1572 2331
rect 1566 2326 1572 2327
rect 1622 2331 1628 2332
rect 1622 2327 1623 2331
rect 1627 2327 1628 2331
rect 1622 2326 1628 2327
rect 1678 2331 1684 2332
rect 1678 2327 1679 2331
rect 1683 2327 1684 2331
rect 2582 2328 2583 2332
rect 2587 2328 2588 2332
rect 2582 2327 2588 2328
rect 1678 2326 1684 2327
rect 110 2323 116 2324
rect 1326 2323 1332 2324
rect 110 2311 116 2312
rect 110 2307 111 2311
rect 115 2307 116 2311
rect 110 2306 116 2307
rect 1326 2311 1332 2312
rect 1326 2307 1327 2311
rect 1331 2307 1332 2311
rect 1326 2306 1332 2307
rect 342 2302 348 2303
rect 342 2298 343 2302
rect 347 2298 348 2302
rect 342 2297 348 2298
rect 398 2302 404 2303
rect 398 2298 399 2302
rect 403 2298 404 2302
rect 398 2297 404 2298
rect 454 2302 460 2303
rect 454 2298 455 2302
rect 459 2298 460 2302
rect 454 2297 460 2298
rect 518 2302 524 2303
rect 518 2298 519 2302
rect 523 2298 524 2302
rect 518 2297 524 2298
rect 582 2302 588 2303
rect 582 2298 583 2302
rect 587 2298 588 2302
rect 582 2297 588 2298
rect 646 2302 652 2303
rect 646 2298 647 2302
rect 651 2298 652 2302
rect 646 2297 652 2298
rect 710 2302 716 2303
rect 710 2298 711 2302
rect 715 2298 716 2302
rect 710 2297 716 2298
rect 774 2302 780 2303
rect 774 2298 775 2302
rect 779 2298 780 2302
rect 774 2297 780 2298
rect 838 2302 844 2303
rect 838 2298 839 2302
rect 843 2298 844 2302
rect 838 2297 844 2298
rect 902 2302 908 2303
rect 902 2298 903 2302
rect 907 2298 908 2302
rect 902 2297 908 2298
rect 966 2302 972 2303
rect 966 2298 967 2302
rect 971 2298 972 2302
rect 966 2297 972 2298
rect 1030 2302 1036 2303
rect 1030 2298 1031 2302
rect 1035 2298 1036 2302
rect 1030 2297 1036 2298
rect 1398 2297 1404 2298
rect 1366 2296 1372 2297
rect 1366 2292 1367 2296
rect 1371 2292 1372 2296
rect 1398 2293 1399 2297
rect 1403 2293 1404 2297
rect 1398 2292 1404 2293
rect 1454 2297 1460 2298
rect 1454 2293 1455 2297
rect 1459 2293 1460 2297
rect 1454 2292 1460 2293
rect 1510 2297 1516 2298
rect 1510 2293 1511 2297
rect 1515 2293 1516 2297
rect 1510 2292 1516 2293
rect 1566 2297 1572 2298
rect 1566 2293 1567 2297
rect 1571 2293 1572 2297
rect 1566 2292 1572 2293
rect 1622 2297 1628 2298
rect 1622 2293 1623 2297
rect 1627 2293 1628 2297
rect 1622 2292 1628 2293
rect 1678 2297 1684 2298
rect 1678 2293 1679 2297
rect 1683 2293 1684 2297
rect 1678 2292 1684 2293
rect 1734 2297 1740 2298
rect 1734 2293 1735 2297
rect 1739 2293 1740 2297
rect 1734 2292 1740 2293
rect 1790 2297 1796 2298
rect 1790 2293 1791 2297
rect 1795 2293 1796 2297
rect 1790 2292 1796 2293
rect 1846 2297 1852 2298
rect 1846 2293 1847 2297
rect 1851 2293 1852 2297
rect 1846 2292 1852 2293
rect 1902 2297 1908 2298
rect 1902 2293 1903 2297
rect 1907 2293 1908 2297
rect 1902 2292 1908 2293
rect 1958 2297 1964 2298
rect 1958 2293 1959 2297
rect 1963 2293 1964 2297
rect 1958 2292 1964 2293
rect 2014 2297 2020 2298
rect 2014 2293 2015 2297
rect 2019 2293 2020 2297
rect 2014 2292 2020 2293
rect 2070 2297 2076 2298
rect 2070 2293 2071 2297
rect 2075 2293 2076 2297
rect 2070 2292 2076 2293
rect 2126 2297 2132 2298
rect 2126 2293 2127 2297
rect 2131 2293 2132 2297
rect 2126 2292 2132 2293
rect 2182 2297 2188 2298
rect 2182 2293 2183 2297
rect 2187 2293 2188 2297
rect 2182 2292 2188 2293
rect 2246 2297 2252 2298
rect 2246 2293 2247 2297
rect 2251 2293 2252 2297
rect 2246 2292 2252 2293
rect 2310 2297 2316 2298
rect 2310 2293 2311 2297
rect 2315 2293 2316 2297
rect 2310 2292 2316 2293
rect 2374 2297 2380 2298
rect 2374 2293 2375 2297
rect 2379 2293 2380 2297
rect 2374 2292 2380 2293
rect 2438 2297 2444 2298
rect 2438 2293 2439 2297
rect 2443 2293 2444 2297
rect 2438 2292 2444 2293
rect 2582 2296 2588 2297
rect 2582 2292 2583 2296
rect 2587 2292 2588 2296
rect 1366 2291 1372 2292
rect 2582 2291 2588 2292
rect 1366 2279 1372 2280
rect 1366 2275 1367 2279
rect 1371 2275 1372 2279
rect 1366 2274 1372 2275
rect 2582 2279 2588 2280
rect 2582 2275 2583 2279
rect 2587 2275 2588 2279
rect 2582 2274 2588 2275
rect 406 2270 412 2271
rect 406 2266 407 2270
rect 411 2266 412 2270
rect 406 2265 412 2266
rect 462 2270 468 2271
rect 462 2266 463 2270
rect 467 2266 468 2270
rect 462 2265 468 2266
rect 518 2270 524 2271
rect 518 2266 519 2270
rect 523 2266 524 2270
rect 518 2265 524 2266
rect 574 2270 580 2271
rect 574 2266 575 2270
rect 579 2266 580 2270
rect 574 2265 580 2266
rect 630 2270 636 2271
rect 630 2266 631 2270
rect 635 2266 636 2270
rect 630 2265 636 2266
rect 686 2270 692 2271
rect 686 2266 687 2270
rect 691 2266 692 2270
rect 686 2265 692 2266
rect 742 2270 748 2271
rect 742 2266 743 2270
rect 747 2266 748 2270
rect 742 2265 748 2266
rect 798 2270 804 2271
rect 798 2266 799 2270
rect 803 2266 804 2270
rect 798 2265 804 2266
rect 854 2270 860 2271
rect 854 2266 855 2270
rect 859 2266 860 2270
rect 854 2265 860 2266
rect 910 2270 916 2271
rect 910 2266 911 2270
rect 915 2266 916 2270
rect 910 2265 916 2266
rect 966 2270 972 2271
rect 966 2266 967 2270
rect 971 2266 972 2270
rect 966 2265 972 2266
rect 1414 2270 1420 2271
rect 1414 2266 1415 2270
rect 1419 2266 1420 2270
rect 1414 2265 1420 2266
rect 1470 2270 1476 2271
rect 1470 2266 1471 2270
rect 1475 2266 1476 2270
rect 1470 2265 1476 2266
rect 1526 2270 1532 2271
rect 1526 2266 1527 2270
rect 1531 2266 1532 2270
rect 1526 2265 1532 2266
rect 1582 2270 1588 2271
rect 1582 2266 1583 2270
rect 1587 2266 1588 2270
rect 1582 2265 1588 2266
rect 1638 2270 1644 2271
rect 1638 2266 1639 2270
rect 1643 2266 1644 2270
rect 1638 2265 1644 2266
rect 1694 2270 1700 2271
rect 1694 2266 1695 2270
rect 1699 2266 1700 2270
rect 1694 2265 1700 2266
rect 1750 2270 1756 2271
rect 1750 2266 1751 2270
rect 1755 2266 1756 2270
rect 1750 2265 1756 2266
rect 1806 2270 1812 2271
rect 1806 2266 1807 2270
rect 1811 2266 1812 2270
rect 1806 2265 1812 2266
rect 1862 2270 1868 2271
rect 1862 2266 1863 2270
rect 1867 2266 1868 2270
rect 1862 2265 1868 2266
rect 1918 2270 1924 2271
rect 1918 2266 1919 2270
rect 1923 2266 1924 2270
rect 1918 2265 1924 2266
rect 1974 2270 1980 2271
rect 1974 2266 1975 2270
rect 1979 2266 1980 2270
rect 1974 2265 1980 2266
rect 2030 2270 2036 2271
rect 2030 2266 2031 2270
rect 2035 2266 2036 2270
rect 2030 2265 2036 2266
rect 2086 2270 2092 2271
rect 2086 2266 2087 2270
rect 2091 2266 2092 2270
rect 2086 2265 2092 2266
rect 2142 2270 2148 2271
rect 2142 2266 2143 2270
rect 2147 2266 2148 2270
rect 2142 2265 2148 2266
rect 2198 2270 2204 2271
rect 2198 2266 2199 2270
rect 2203 2266 2204 2270
rect 2198 2265 2204 2266
rect 2262 2270 2268 2271
rect 2262 2266 2263 2270
rect 2267 2266 2268 2270
rect 2262 2265 2268 2266
rect 2326 2270 2332 2271
rect 2326 2266 2327 2270
rect 2331 2266 2332 2270
rect 2326 2265 2332 2266
rect 2390 2270 2396 2271
rect 2390 2266 2391 2270
rect 2395 2266 2396 2270
rect 2390 2265 2396 2266
rect 2454 2270 2460 2271
rect 2454 2266 2455 2270
rect 2459 2266 2460 2270
rect 2454 2265 2460 2266
rect 110 2261 116 2262
rect 110 2257 111 2261
rect 115 2257 116 2261
rect 110 2256 116 2257
rect 1326 2261 1332 2262
rect 1326 2257 1327 2261
rect 1331 2257 1332 2261
rect 1326 2256 1332 2257
rect 1414 2246 1420 2247
rect 110 2244 116 2245
rect 1326 2244 1332 2245
rect 110 2240 111 2244
rect 115 2240 116 2244
rect 110 2239 116 2240
rect 390 2243 396 2244
rect 390 2239 391 2243
rect 395 2239 396 2243
rect 390 2238 396 2239
rect 446 2243 452 2244
rect 446 2239 447 2243
rect 451 2239 452 2243
rect 446 2238 452 2239
rect 502 2243 508 2244
rect 502 2239 503 2243
rect 507 2239 508 2243
rect 502 2238 508 2239
rect 558 2243 564 2244
rect 558 2239 559 2243
rect 563 2239 564 2243
rect 558 2238 564 2239
rect 614 2243 620 2244
rect 614 2239 615 2243
rect 619 2239 620 2243
rect 614 2238 620 2239
rect 670 2243 676 2244
rect 670 2239 671 2243
rect 675 2239 676 2243
rect 670 2238 676 2239
rect 726 2243 732 2244
rect 726 2239 727 2243
rect 731 2239 732 2243
rect 726 2238 732 2239
rect 782 2243 788 2244
rect 782 2239 783 2243
rect 787 2239 788 2243
rect 782 2238 788 2239
rect 838 2243 844 2244
rect 838 2239 839 2243
rect 843 2239 844 2243
rect 838 2238 844 2239
rect 894 2243 900 2244
rect 894 2239 895 2243
rect 899 2239 900 2243
rect 894 2238 900 2239
rect 950 2243 956 2244
rect 950 2239 951 2243
rect 955 2239 956 2243
rect 1326 2240 1327 2244
rect 1331 2240 1332 2244
rect 1414 2242 1415 2246
rect 1419 2242 1420 2246
rect 1414 2241 1420 2242
rect 1510 2246 1516 2247
rect 1510 2242 1511 2246
rect 1515 2242 1516 2246
rect 1510 2241 1516 2242
rect 1622 2246 1628 2247
rect 1622 2242 1623 2246
rect 1627 2242 1628 2246
rect 1622 2241 1628 2242
rect 1726 2246 1732 2247
rect 1726 2242 1727 2246
rect 1731 2242 1732 2246
rect 1726 2241 1732 2242
rect 1822 2246 1828 2247
rect 1822 2242 1823 2246
rect 1827 2242 1828 2246
rect 1822 2241 1828 2242
rect 1902 2246 1908 2247
rect 1902 2242 1903 2246
rect 1907 2242 1908 2246
rect 1902 2241 1908 2242
rect 1982 2246 1988 2247
rect 1982 2242 1983 2246
rect 1987 2242 1988 2246
rect 1982 2241 1988 2242
rect 2054 2246 2060 2247
rect 2054 2242 2055 2246
rect 2059 2242 2060 2246
rect 2054 2241 2060 2242
rect 2118 2246 2124 2247
rect 2118 2242 2119 2246
rect 2123 2242 2124 2246
rect 2118 2241 2124 2242
rect 2190 2246 2196 2247
rect 2190 2242 2191 2246
rect 2195 2242 2196 2246
rect 2190 2241 2196 2242
rect 2262 2246 2268 2247
rect 2262 2242 2263 2246
rect 2267 2242 2268 2246
rect 2262 2241 2268 2242
rect 2334 2246 2340 2247
rect 2334 2242 2335 2246
rect 2339 2242 2340 2246
rect 2334 2241 2340 2242
rect 1326 2239 1332 2240
rect 950 2238 956 2239
rect 1366 2237 1372 2238
rect 1366 2233 1367 2237
rect 1371 2233 1372 2237
rect 1366 2232 1372 2233
rect 2582 2237 2588 2238
rect 2582 2233 2583 2237
rect 2587 2233 2588 2237
rect 2582 2232 2588 2233
rect 1366 2220 1372 2221
rect 2582 2220 2588 2221
rect 1366 2216 1367 2220
rect 1371 2216 1372 2220
rect 1366 2215 1372 2216
rect 1398 2219 1404 2220
rect 1398 2215 1399 2219
rect 1403 2215 1404 2219
rect 1398 2214 1404 2215
rect 1494 2219 1500 2220
rect 1494 2215 1495 2219
rect 1499 2215 1500 2219
rect 1494 2214 1500 2215
rect 1606 2219 1612 2220
rect 1606 2215 1607 2219
rect 1611 2215 1612 2219
rect 1606 2214 1612 2215
rect 1710 2219 1716 2220
rect 1710 2215 1711 2219
rect 1715 2215 1716 2219
rect 1710 2214 1716 2215
rect 1806 2219 1812 2220
rect 1806 2215 1807 2219
rect 1811 2215 1812 2219
rect 1806 2214 1812 2215
rect 1886 2219 1892 2220
rect 1886 2215 1887 2219
rect 1891 2215 1892 2219
rect 1886 2214 1892 2215
rect 1966 2219 1972 2220
rect 1966 2215 1967 2219
rect 1971 2215 1972 2219
rect 1966 2214 1972 2215
rect 2038 2219 2044 2220
rect 2038 2215 2039 2219
rect 2043 2215 2044 2219
rect 2038 2214 2044 2215
rect 2102 2219 2108 2220
rect 2102 2215 2103 2219
rect 2107 2215 2108 2219
rect 2102 2214 2108 2215
rect 2174 2219 2180 2220
rect 2174 2215 2175 2219
rect 2179 2215 2180 2219
rect 2174 2214 2180 2215
rect 2246 2219 2252 2220
rect 2246 2215 2247 2219
rect 2251 2215 2252 2219
rect 2246 2214 2252 2215
rect 2318 2219 2324 2220
rect 2318 2215 2319 2219
rect 2323 2215 2324 2219
rect 2582 2216 2583 2220
rect 2587 2216 2588 2220
rect 2582 2215 2588 2216
rect 2318 2214 2324 2215
rect 422 2205 428 2206
rect 110 2204 116 2205
rect 110 2200 111 2204
rect 115 2200 116 2204
rect 422 2201 423 2205
rect 427 2201 428 2205
rect 422 2200 428 2201
rect 478 2205 484 2206
rect 478 2201 479 2205
rect 483 2201 484 2205
rect 478 2200 484 2201
rect 534 2205 540 2206
rect 534 2201 535 2205
rect 539 2201 540 2205
rect 534 2200 540 2201
rect 590 2205 596 2206
rect 590 2201 591 2205
rect 595 2201 596 2205
rect 590 2200 596 2201
rect 646 2205 652 2206
rect 646 2201 647 2205
rect 651 2201 652 2205
rect 646 2200 652 2201
rect 710 2205 716 2206
rect 710 2201 711 2205
rect 715 2201 716 2205
rect 710 2200 716 2201
rect 782 2205 788 2206
rect 782 2201 783 2205
rect 787 2201 788 2205
rect 782 2200 788 2201
rect 854 2205 860 2206
rect 854 2201 855 2205
rect 859 2201 860 2205
rect 854 2200 860 2201
rect 926 2205 932 2206
rect 926 2201 927 2205
rect 931 2201 932 2205
rect 926 2200 932 2201
rect 998 2205 1004 2206
rect 998 2201 999 2205
rect 1003 2201 1004 2205
rect 998 2200 1004 2201
rect 1070 2205 1076 2206
rect 1070 2201 1071 2205
rect 1075 2201 1076 2205
rect 1070 2200 1076 2201
rect 1142 2205 1148 2206
rect 1142 2201 1143 2205
rect 1147 2201 1148 2205
rect 1142 2200 1148 2201
rect 1214 2205 1220 2206
rect 1214 2201 1215 2205
rect 1219 2201 1220 2205
rect 1214 2200 1220 2201
rect 1270 2205 1276 2206
rect 1270 2201 1271 2205
rect 1275 2201 1276 2205
rect 1270 2200 1276 2201
rect 1326 2204 1332 2205
rect 1326 2200 1327 2204
rect 1331 2200 1332 2204
rect 110 2199 116 2200
rect 1326 2199 1332 2200
rect 110 2187 116 2188
rect 110 2183 111 2187
rect 115 2183 116 2187
rect 110 2182 116 2183
rect 1326 2187 1332 2188
rect 1326 2183 1327 2187
rect 1331 2183 1332 2187
rect 1326 2182 1332 2183
rect 1750 2181 1756 2182
rect 1366 2180 1372 2181
rect 438 2178 444 2179
rect 438 2174 439 2178
rect 443 2174 444 2178
rect 438 2173 444 2174
rect 494 2178 500 2179
rect 494 2174 495 2178
rect 499 2174 500 2178
rect 494 2173 500 2174
rect 550 2178 556 2179
rect 550 2174 551 2178
rect 555 2174 556 2178
rect 550 2173 556 2174
rect 606 2178 612 2179
rect 606 2174 607 2178
rect 611 2174 612 2178
rect 606 2173 612 2174
rect 662 2178 668 2179
rect 662 2174 663 2178
rect 667 2174 668 2178
rect 662 2173 668 2174
rect 726 2178 732 2179
rect 726 2174 727 2178
rect 731 2174 732 2178
rect 726 2173 732 2174
rect 798 2178 804 2179
rect 798 2174 799 2178
rect 803 2174 804 2178
rect 798 2173 804 2174
rect 870 2178 876 2179
rect 870 2174 871 2178
rect 875 2174 876 2178
rect 870 2173 876 2174
rect 942 2178 948 2179
rect 942 2174 943 2178
rect 947 2174 948 2178
rect 942 2173 948 2174
rect 1014 2178 1020 2179
rect 1014 2174 1015 2178
rect 1019 2174 1020 2178
rect 1014 2173 1020 2174
rect 1086 2178 1092 2179
rect 1086 2174 1087 2178
rect 1091 2174 1092 2178
rect 1086 2173 1092 2174
rect 1158 2178 1164 2179
rect 1158 2174 1159 2178
rect 1163 2174 1164 2178
rect 1158 2173 1164 2174
rect 1230 2178 1236 2179
rect 1230 2174 1231 2178
rect 1235 2174 1236 2178
rect 1230 2173 1236 2174
rect 1286 2178 1292 2179
rect 1286 2174 1287 2178
rect 1291 2174 1292 2178
rect 1366 2176 1367 2180
rect 1371 2176 1372 2180
rect 1750 2177 1751 2181
rect 1755 2177 1756 2181
rect 1750 2176 1756 2177
rect 1838 2181 1844 2182
rect 1838 2177 1839 2181
rect 1843 2177 1844 2181
rect 1838 2176 1844 2177
rect 1926 2181 1932 2182
rect 1926 2177 1927 2181
rect 1931 2177 1932 2181
rect 1926 2176 1932 2177
rect 2006 2181 2012 2182
rect 2006 2177 2007 2181
rect 2011 2177 2012 2181
rect 2006 2176 2012 2177
rect 2086 2181 2092 2182
rect 2086 2177 2087 2181
rect 2091 2177 2092 2181
rect 2086 2176 2092 2177
rect 2166 2181 2172 2182
rect 2166 2177 2167 2181
rect 2171 2177 2172 2181
rect 2166 2176 2172 2177
rect 2246 2181 2252 2182
rect 2246 2177 2247 2181
rect 2251 2177 2252 2181
rect 2246 2176 2252 2177
rect 2334 2181 2340 2182
rect 2334 2177 2335 2181
rect 2339 2177 2340 2181
rect 2334 2176 2340 2177
rect 2422 2181 2428 2182
rect 2422 2177 2423 2181
rect 2427 2177 2428 2181
rect 2422 2176 2428 2177
rect 2582 2180 2588 2181
rect 2582 2176 2583 2180
rect 2587 2176 2588 2180
rect 1366 2175 1372 2176
rect 2582 2175 2588 2176
rect 1286 2173 1292 2174
rect 1366 2163 1372 2164
rect 1366 2159 1367 2163
rect 1371 2159 1372 2163
rect 1366 2158 1372 2159
rect 2582 2163 2588 2164
rect 2582 2159 2583 2163
rect 2587 2159 2588 2163
rect 2582 2158 2588 2159
rect 1766 2154 1772 2155
rect 1766 2150 1767 2154
rect 1771 2150 1772 2154
rect 1766 2149 1772 2150
rect 1854 2154 1860 2155
rect 1854 2150 1855 2154
rect 1859 2150 1860 2154
rect 1854 2149 1860 2150
rect 1942 2154 1948 2155
rect 1942 2150 1943 2154
rect 1947 2150 1948 2154
rect 1942 2149 1948 2150
rect 2022 2154 2028 2155
rect 2022 2150 2023 2154
rect 2027 2150 2028 2154
rect 2022 2149 2028 2150
rect 2102 2154 2108 2155
rect 2102 2150 2103 2154
rect 2107 2150 2108 2154
rect 2102 2149 2108 2150
rect 2182 2154 2188 2155
rect 2182 2150 2183 2154
rect 2187 2150 2188 2154
rect 2182 2149 2188 2150
rect 2262 2154 2268 2155
rect 2262 2150 2263 2154
rect 2267 2150 2268 2154
rect 2262 2149 2268 2150
rect 2350 2154 2356 2155
rect 2350 2150 2351 2154
rect 2355 2150 2356 2154
rect 2350 2149 2356 2150
rect 2438 2154 2444 2155
rect 2438 2150 2439 2154
rect 2443 2150 2444 2154
rect 2438 2149 2444 2150
rect 198 2146 204 2147
rect 198 2142 199 2146
rect 203 2142 204 2146
rect 198 2141 204 2142
rect 270 2146 276 2147
rect 270 2142 271 2146
rect 275 2142 276 2146
rect 270 2141 276 2142
rect 350 2146 356 2147
rect 350 2142 351 2146
rect 355 2142 356 2146
rect 350 2141 356 2142
rect 446 2146 452 2147
rect 446 2142 447 2146
rect 451 2142 452 2146
rect 446 2141 452 2142
rect 550 2146 556 2147
rect 550 2142 551 2146
rect 555 2142 556 2146
rect 550 2141 556 2142
rect 662 2146 668 2147
rect 662 2142 663 2146
rect 667 2142 668 2146
rect 662 2141 668 2142
rect 774 2146 780 2147
rect 774 2142 775 2146
rect 779 2142 780 2146
rect 774 2141 780 2142
rect 878 2146 884 2147
rect 878 2142 879 2146
rect 883 2142 884 2146
rect 878 2141 884 2142
rect 982 2146 988 2147
rect 982 2142 983 2146
rect 987 2142 988 2146
rect 982 2141 988 2142
rect 1078 2146 1084 2147
rect 1078 2142 1079 2146
rect 1083 2142 1084 2146
rect 1078 2141 1084 2142
rect 1182 2146 1188 2147
rect 1182 2142 1183 2146
rect 1187 2142 1188 2146
rect 1182 2141 1188 2142
rect 1286 2146 1292 2147
rect 1286 2142 1287 2146
rect 1291 2142 1292 2146
rect 1286 2141 1292 2142
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 110 2132 116 2133
rect 1326 2137 1332 2138
rect 1326 2133 1327 2137
rect 1331 2133 1332 2137
rect 1326 2132 1332 2133
rect 1606 2130 1612 2131
rect 1606 2126 1607 2130
rect 1611 2126 1612 2130
rect 1606 2125 1612 2126
rect 1678 2130 1684 2131
rect 1678 2126 1679 2130
rect 1683 2126 1684 2130
rect 1678 2125 1684 2126
rect 1766 2130 1772 2131
rect 1766 2126 1767 2130
rect 1771 2126 1772 2130
rect 1766 2125 1772 2126
rect 1862 2130 1868 2131
rect 1862 2126 1863 2130
rect 1867 2126 1868 2130
rect 1862 2125 1868 2126
rect 1958 2130 1964 2131
rect 1958 2126 1959 2130
rect 1963 2126 1964 2130
rect 1958 2125 1964 2126
rect 2062 2130 2068 2131
rect 2062 2126 2063 2130
rect 2067 2126 2068 2130
rect 2062 2125 2068 2126
rect 2158 2130 2164 2131
rect 2158 2126 2159 2130
rect 2163 2126 2164 2130
rect 2158 2125 2164 2126
rect 2254 2130 2260 2131
rect 2254 2126 2255 2130
rect 2259 2126 2260 2130
rect 2254 2125 2260 2126
rect 2350 2130 2356 2131
rect 2350 2126 2351 2130
rect 2355 2126 2356 2130
rect 2350 2125 2356 2126
rect 2446 2130 2452 2131
rect 2446 2126 2447 2130
rect 2451 2126 2452 2130
rect 2446 2125 2452 2126
rect 2542 2130 2548 2131
rect 2542 2126 2543 2130
rect 2547 2126 2548 2130
rect 2542 2125 2548 2126
rect 1366 2121 1372 2122
rect 110 2120 116 2121
rect 1326 2120 1332 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 110 2115 116 2116
rect 182 2119 188 2120
rect 182 2115 183 2119
rect 187 2115 188 2119
rect 182 2114 188 2115
rect 254 2119 260 2120
rect 254 2115 255 2119
rect 259 2115 260 2119
rect 254 2114 260 2115
rect 334 2119 340 2120
rect 334 2115 335 2119
rect 339 2115 340 2119
rect 334 2114 340 2115
rect 430 2119 436 2120
rect 430 2115 431 2119
rect 435 2115 436 2119
rect 430 2114 436 2115
rect 534 2119 540 2120
rect 534 2115 535 2119
rect 539 2115 540 2119
rect 534 2114 540 2115
rect 646 2119 652 2120
rect 646 2115 647 2119
rect 651 2115 652 2119
rect 646 2114 652 2115
rect 758 2119 764 2120
rect 758 2115 759 2119
rect 763 2115 764 2119
rect 758 2114 764 2115
rect 862 2119 868 2120
rect 862 2115 863 2119
rect 867 2115 868 2119
rect 862 2114 868 2115
rect 966 2119 972 2120
rect 966 2115 967 2119
rect 971 2115 972 2119
rect 966 2114 972 2115
rect 1062 2119 1068 2120
rect 1062 2115 1063 2119
rect 1067 2115 1068 2119
rect 1062 2114 1068 2115
rect 1166 2119 1172 2120
rect 1166 2115 1167 2119
rect 1171 2115 1172 2119
rect 1166 2114 1172 2115
rect 1270 2119 1276 2120
rect 1270 2115 1271 2119
rect 1275 2115 1276 2119
rect 1326 2116 1327 2120
rect 1331 2116 1332 2120
rect 1366 2117 1367 2121
rect 1371 2117 1372 2121
rect 1366 2116 1372 2117
rect 2582 2121 2588 2122
rect 2582 2117 2583 2121
rect 2587 2117 2588 2121
rect 2582 2116 2588 2117
rect 1326 2115 1332 2116
rect 1270 2114 1276 2115
rect 1366 2104 1372 2105
rect 2582 2104 2588 2105
rect 1366 2100 1367 2104
rect 1371 2100 1372 2104
rect 1366 2099 1372 2100
rect 1590 2103 1596 2104
rect 1590 2099 1591 2103
rect 1595 2099 1596 2103
rect 1590 2098 1596 2099
rect 1662 2103 1668 2104
rect 1662 2099 1663 2103
rect 1667 2099 1668 2103
rect 1662 2098 1668 2099
rect 1750 2103 1756 2104
rect 1750 2099 1751 2103
rect 1755 2099 1756 2103
rect 1750 2098 1756 2099
rect 1846 2103 1852 2104
rect 1846 2099 1847 2103
rect 1851 2099 1852 2103
rect 1846 2098 1852 2099
rect 1942 2103 1948 2104
rect 1942 2099 1943 2103
rect 1947 2099 1948 2103
rect 1942 2098 1948 2099
rect 2046 2103 2052 2104
rect 2046 2099 2047 2103
rect 2051 2099 2052 2103
rect 2046 2098 2052 2099
rect 2142 2103 2148 2104
rect 2142 2099 2143 2103
rect 2147 2099 2148 2103
rect 2142 2098 2148 2099
rect 2238 2103 2244 2104
rect 2238 2099 2239 2103
rect 2243 2099 2244 2103
rect 2238 2098 2244 2099
rect 2334 2103 2340 2104
rect 2334 2099 2335 2103
rect 2339 2099 2340 2103
rect 2334 2098 2340 2099
rect 2430 2103 2436 2104
rect 2430 2099 2431 2103
rect 2435 2099 2436 2103
rect 2430 2098 2436 2099
rect 2526 2103 2532 2104
rect 2526 2099 2527 2103
rect 2531 2099 2532 2103
rect 2582 2100 2583 2104
rect 2587 2100 2588 2104
rect 2582 2099 2588 2100
rect 2526 2098 2532 2099
rect 142 2073 148 2074
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 142 2069 143 2073
rect 147 2069 148 2073
rect 142 2068 148 2069
rect 198 2073 204 2074
rect 198 2069 199 2073
rect 203 2069 204 2073
rect 198 2068 204 2069
rect 270 2073 276 2074
rect 270 2069 271 2073
rect 275 2069 276 2073
rect 270 2068 276 2069
rect 366 2073 372 2074
rect 366 2069 367 2073
rect 371 2069 372 2073
rect 366 2068 372 2069
rect 462 2073 468 2074
rect 462 2069 463 2073
rect 467 2069 468 2073
rect 462 2068 468 2069
rect 566 2073 572 2074
rect 566 2069 567 2073
rect 571 2069 572 2073
rect 566 2068 572 2069
rect 662 2073 668 2074
rect 662 2069 663 2073
rect 667 2069 668 2073
rect 662 2068 668 2069
rect 758 2073 764 2074
rect 758 2069 759 2073
rect 763 2069 764 2073
rect 758 2068 764 2069
rect 846 2073 852 2074
rect 846 2069 847 2073
rect 851 2069 852 2073
rect 846 2068 852 2069
rect 926 2073 932 2074
rect 926 2069 927 2073
rect 931 2069 932 2073
rect 926 2068 932 2069
rect 1006 2073 1012 2074
rect 1006 2069 1007 2073
rect 1011 2069 1012 2073
rect 1006 2068 1012 2069
rect 1094 2073 1100 2074
rect 1094 2069 1095 2073
rect 1099 2069 1100 2073
rect 1094 2068 1100 2069
rect 1182 2073 1188 2074
rect 1182 2069 1183 2073
rect 1187 2069 1188 2073
rect 1182 2068 1188 2069
rect 1326 2072 1332 2073
rect 1326 2068 1327 2072
rect 1331 2068 1332 2072
rect 1486 2069 1492 2070
rect 110 2067 116 2068
rect 1326 2067 1332 2068
rect 1366 2068 1372 2069
rect 1366 2064 1367 2068
rect 1371 2064 1372 2068
rect 1486 2065 1487 2069
rect 1491 2065 1492 2069
rect 1486 2064 1492 2065
rect 1582 2069 1588 2070
rect 1582 2065 1583 2069
rect 1587 2065 1588 2069
rect 1582 2064 1588 2065
rect 1678 2069 1684 2070
rect 1678 2065 1679 2069
rect 1683 2065 1684 2069
rect 1678 2064 1684 2065
rect 1782 2069 1788 2070
rect 1782 2065 1783 2069
rect 1787 2065 1788 2069
rect 1782 2064 1788 2065
rect 1886 2069 1892 2070
rect 1886 2065 1887 2069
rect 1891 2065 1892 2069
rect 1886 2064 1892 2065
rect 1982 2069 1988 2070
rect 1982 2065 1983 2069
rect 1987 2065 1988 2069
rect 1982 2064 1988 2065
rect 2078 2069 2084 2070
rect 2078 2065 2079 2069
rect 2083 2065 2084 2069
rect 2078 2064 2084 2065
rect 2166 2069 2172 2070
rect 2166 2065 2167 2069
rect 2171 2065 2172 2069
rect 2166 2064 2172 2065
rect 2254 2069 2260 2070
rect 2254 2065 2255 2069
rect 2259 2065 2260 2069
rect 2254 2064 2260 2065
rect 2342 2069 2348 2070
rect 2342 2065 2343 2069
rect 2347 2065 2348 2069
rect 2342 2064 2348 2065
rect 2438 2069 2444 2070
rect 2438 2065 2439 2069
rect 2443 2065 2444 2069
rect 2438 2064 2444 2065
rect 2526 2069 2532 2070
rect 2526 2065 2527 2069
rect 2531 2065 2532 2069
rect 2526 2064 2532 2065
rect 2582 2068 2588 2069
rect 2582 2064 2583 2068
rect 2587 2064 2588 2068
rect 1366 2063 1372 2064
rect 2582 2063 2588 2064
rect 110 2055 116 2056
rect 110 2051 111 2055
rect 115 2051 116 2055
rect 110 2050 116 2051
rect 1326 2055 1332 2056
rect 1326 2051 1327 2055
rect 1331 2051 1332 2055
rect 1326 2050 1332 2051
rect 1366 2051 1372 2052
rect 1366 2047 1367 2051
rect 1371 2047 1372 2051
rect 158 2046 164 2047
rect 158 2042 159 2046
rect 163 2042 164 2046
rect 158 2041 164 2042
rect 214 2046 220 2047
rect 214 2042 215 2046
rect 219 2042 220 2046
rect 214 2041 220 2042
rect 286 2046 292 2047
rect 286 2042 287 2046
rect 291 2042 292 2046
rect 286 2041 292 2042
rect 382 2046 388 2047
rect 382 2042 383 2046
rect 387 2042 388 2046
rect 382 2041 388 2042
rect 478 2046 484 2047
rect 478 2042 479 2046
rect 483 2042 484 2046
rect 478 2041 484 2042
rect 582 2046 588 2047
rect 582 2042 583 2046
rect 587 2042 588 2046
rect 582 2041 588 2042
rect 678 2046 684 2047
rect 678 2042 679 2046
rect 683 2042 684 2046
rect 678 2041 684 2042
rect 774 2046 780 2047
rect 774 2042 775 2046
rect 779 2042 780 2046
rect 774 2041 780 2042
rect 862 2046 868 2047
rect 862 2042 863 2046
rect 867 2042 868 2046
rect 862 2041 868 2042
rect 942 2046 948 2047
rect 942 2042 943 2046
rect 947 2042 948 2046
rect 942 2041 948 2042
rect 1022 2046 1028 2047
rect 1022 2042 1023 2046
rect 1027 2042 1028 2046
rect 1022 2041 1028 2042
rect 1110 2046 1116 2047
rect 1110 2042 1111 2046
rect 1115 2042 1116 2046
rect 1110 2041 1116 2042
rect 1198 2046 1204 2047
rect 1366 2046 1372 2047
rect 2582 2051 2588 2052
rect 2582 2047 2583 2051
rect 2587 2047 2588 2051
rect 2582 2046 2588 2047
rect 1198 2042 1199 2046
rect 1203 2042 1204 2046
rect 1198 2041 1204 2042
rect 1502 2042 1508 2043
rect 1502 2038 1503 2042
rect 1507 2038 1508 2042
rect 1502 2037 1508 2038
rect 1598 2042 1604 2043
rect 1598 2038 1599 2042
rect 1603 2038 1604 2042
rect 1598 2037 1604 2038
rect 1694 2042 1700 2043
rect 1694 2038 1695 2042
rect 1699 2038 1700 2042
rect 1694 2037 1700 2038
rect 1798 2042 1804 2043
rect 1798 2038 1799 2042
rect 1803 2038 1804 2042
rect 1798 2037 1804 2038
rect 1902 2042 1908 2043
rect 1902 2038 1903 2042
rect 1907 2038 1908 2042
rect 1902 2037 1908 2038
rect 1998 2042 2004 2043
rect 1998 2038 1999 2042
rect 2003 2038 2004 2042
rect 1998 2037 2004 2038
rect 2094 2042 2100 2043
rect 2094 2038 2095 2042
rect 2099 2038 2100 2042
rect 2094 2037 2100 2038
rect 2182 2042 2188 2043
rect 2182 2038 2183 2042
rect 2187 2038 2188 2042
rect 2182 2037 2188 2038
rect 2270 2042 2276 2043
rect 2270 2038 2271 2042
rect 2275 2038 2276 2042
rect 2270 2037 2276 2038
rect 2358 2042 2364 2043
rect 2358 2038 2359 2042
rect 2363 2038 2364 2042
rect 2358 2037 2364 2038
rect 2454 2042 2460 2043
rect 2454 2038 2455 2042
rect 2459 2038 2460 2042
rect 2454 2037 2460 2038
rect 2542 2042 2548 2043
rect 2542 2038 2543 2042
rect 2547 2038 2548 2042
rect 2542 2037 2548 2038
rect 1414 2018 1420 2019
rect 174 2014 180 2015
rect 174 2010 175 2014
rect 179 2010 180 2014
rect 174 2009 180 2010
rect 238 2014 244 2015
rect 238 2010 239 2014
rect 243 2010 244 2014
rect 238 2009 244 2010
rect 310 2014 316 2015
rect 310 2010 311 2014
rect 315 2010 316 2014
rect 310 2009 316 2010
rect 390 2014 396 2015
rect 390 2010 391 2014
rect 395 2010 396 2014
rect 390 2009 396 2010
rect 470 2014 476 2015
rect 470 2010 471 2014
rect 475 2010 476 2014
rect 470 2009 476 2010
rect 558 2014 564 2015
rect 558 2010 559 2014
rect 563 2010 564 2014
rect 558 2009 564 2010
rect 646 2014 652 2015
rect 646 2010 647 2014
rect 651 2010 652 2014
rect 646 2009 652 2010
rect 734 2014 740 2015
rect 734 2010 735 2014
rect 739 2010 740 2014
rect 734 2009 740 2010
rect 822 2014 828 2015
rect 822 2010 823 2014
rect 827 2010 828 2014
rect 822 2009 828 2010
rect 910 2014 916 2015
rect 910 2010 911 2014
rect 915 2010 916 2014
rect 910 2009 916 2010
rect 1006 2014 1012 2015
rect 1006 2010 1007 2014
rect 1011 2010 1012 2014
rect 1006 2009 1012 2010
rect 1102 2014 1108 2015
rect 1102 2010 1103 2014
rect 1107 2010 1108 2014
rect 1414 2014 1415 2018
rect 1419 2014 1420 2018
rect 1414 2013 1420 2014
rect 1470 2018 1476 2019
rect 1470 2014 1471 2018
rect 1475 2014 1476 2018
rect 1470 2013 1476 2014
rect 1534 2018 1540 2019
rect 1534 2014 1535 2018
rect 1539 2014 1540 2018
rect 1534 2013 1540 2014
rect 1614 2018 1620 2019
rect 1614 2014 1615 2018
rect 1619 2014 1620 2018
rect 1614 2013 1620 2014
rect 1702 2018 1708 2019
rect 1702 2014 1703 2018
rect 1707 2014 1708 2018
rect 1702 2013 1708 2014
rect 1790 2018 1796 2019
rect 1790 2014 1791 2018
rect 1795 2014 1796 2018
rect 1790 2013 1796 2014
rect 1886 2018 1892 2019
rect 1886 2014 1887 2018
rect 1891 2014 1892 2018
rect 1886 2013 1892 2014
rect 1982 2018 1988 2019
rect 1982 2014 1983 2018
rect 1987 2014 1988 2018
rect 1982 2013 1988 2014
rect 2078 2018 2084 2019
rect 2078 2014 2079 2018
rect 2083 2014 2084 2018
rect 2078 2013 2084 2014
rect 2174 2018 2180 2019
rect 2174 2014 2175 2018
rect 2179 2014 2180 2018
rect 2174 2013 2180 2014
rect 2270 2018 2276 2019
rect 2270 2014 2271 2018
rect 2275 2014 2276 2018
rect 2270 2013 2276 2014
rect 2366 2018 2372 2019
rect 2366 2014 2367 2018
rect 2371 2014 2372 2018
rect 2366 2013 2372 2014
rect 2462 2018 2468 2019
rect 2462 2014 2463 2018
rect 2467 2014 2468 2018
rect 2462 2013 2468 2014
rect 2542 2018 2548 2019
rect 2542 2014 2543 2018
rect 2547 2014 2548 2018
rect 2542 2013 2548 2014
rect 1102 2009 1108 2010
rect 1366 2009 1372 2010
rect 110 2005 116 2006
rect 110 2001 111 2005
rect 115 2001 116 2005
rect 110 2000 116 2001
rect 1326 2005 1332 2006
rect 1326 2001 1327 2005
rect 1331 2001 1332 2005
rect 1366 2005 1367 2009
rect 1371 2005 1372 2009
rect 1366 2004 1372 2005
rect 2582 2009 2588 2010
rect 2582 2005 2583 2009
rect 2587 2005 2588 2009
rect 2582 2004 2588 2005
rect 1326 2000 1332 2001
rect 1366 1992 1372 1993
rect 2582 1992 2588 1993
rect 110 1988 116 1989
rect 1326 1988 1332 1989
rect 110 1984 111 1988
rect 115 1984 116 1988
rect 110 1983 116 1984
rect 158 1987 164 1988
rect 158 1983 159 1987
rect 163 1983 164 1987
rect 158 1982 164 1983
rect 222 1987 228 1988
rect 222 1983 223 1987
rect 227 1983 228 1987
rect 222 1982 228 1983
rect 294 1987 300 1988
rect 294 1983 295 1987
rect 299 1983 300 1987
rect 294 1982 300 1983
rect 374 1987 380 1988
rect 374 1983 375 1987
rect 379 1983 380 1987
rect 374 1982 380 1983
rect 454 1987 460 1988
rect 454 1983 455 1987
rect 459 1983 460 1987
rect 454 1982 460 1983
rect 542 1987 548 1988
rect 542 1983 543 1987
rect 547 1983 548 1987
rect 542 1982 548 1983
rect 630 1987 636 1988
rect 630 1983 631 1987
rect 635 1983 636 1987
rect 630 1982 636 1983
rect 718 1987 724 1988
rect 718 1983 719 1987
rect 723 1983 724 1987
rect 718 1982 724 1983
rect 806 1987 812 1988
rect 806 1983 807 1987
rect 811 1983 812 1987
rect 806 1982 812 1983
rect 894 1987 900 1988
rect 894 1983 895 1987
rect 899 1983 900 1987
rect 894 1982 900 1983
rect 990 1987 996 1988
rect 990 1983 991 1987
rect 995 1983 996 1987
rect 990 1982 996 1983
rect 1086 1987 1092 1988
rect 1086 1983 1087 1987
rect 1091 1983 1092 1987
rect 1326 1984 1327 1988
rect 1331 1984 1332 1988
rect 1366 1988 1367 1992
rect 1371 1988 1372 1992
rect 1366 1987 1372 1988
rect 1398 1991 1404 1992
rect 1398 1987 1399 1991
rect 1403 1987 1404 1991
rect 1398 1986 1404 1987
rect 1454 1991 1460 1992
rect 1454 1987 1455 1991
rect 1459 1987 1460 1991
rect 1454 1986 1460 1987
rect 1518 1991 1524 1992
rect 1518 1987 1519 1991
rect 1523 1987 1524 1991
rect 1518 1986 1524 1987
rect 1598 1991 1604 1992
rect 1598 1987 1599 1991
rect 1603 1987 1604 1991
rect 1598 1986 1604 1987
rect 1686 1991 1692 1992
rect 1686 1987 1687 1991
rect 1691 1987 1692 1991
rect 1686 1986 1692 1987
rect 1774 1991 1780 1992
rect 1774 1987 1775 1991
rect 1779 1987 1780 1991
rect 1774 1986 1780 1987
rect 1870 1991 1876 1992
rect 1870 1987 1871 1991
rect 1875 1987 1876 1991
rect 1870 1986 1876 1987
rect 1966 1991 1972 1992
rect 1966 1987 1967 1991
rect 1971 1987 1972 1991
rect 1966 1986 1972 1987
rect 2062 1991 2068 1992
rect 2062 1987 2063 1991
rect 2067 1987 2068 1991
rect 2062 1986 2068 1987
rect 2158 1991 2164 1992
rect 2158 1987 2159 1991
rect 2163 1987 2164 1991
rect 2158 1986 2164 1987
rect 2254 1991 2260 1992
rect 2254 1987 2255 1991
rect 2259 1987 2260 1991
rect 2254 1986 2260 1987
rect 2350 1991 2356 1992
rect 2350 1987 2351 1991
rect 2355 1987 2356 1991
rect 2350 1986 2356 1987
rect 2446 1991 2452 1992
rect 2446 1987 2447 1991
rect 2451 1987 2452 1991
rect 2446 1986 2452 1987
rect 2526 1991 2532 1992
rect 2526 1987 2527 1991
rect 2531 1987 2532 1991
rect 2582 1988 2583 1992
rect 2587 1988 2588 1992
rect 2582 1987 2588 1988
rect 2526 1986 2532 1987
rect 1326 1983 1332 1984
rect 1086 1982 1092 1983
rect 382 1953 388 1954
rect 110 1952 116 1953
rect 110 1948 111 1952
rect 115 1948 116 1952
rect 382 1949 383 1953
rect 387 1949 388 1953
rect 382 1948 388 1949
rect 438 1953 444 1954
rect 438 1949 439 1953
rect 443 1949 444 1953
rect 438 1948 444 1949
rect 494 1953 500 1954
rect 494 1949 495 1953
rect 499 1949 500 1953
rect 494 1948 500 1949
rect 550 1953 556 1954
rect 550 1949 551 1953
rect 555 1949 556 1953
rect 550 1948 556 1949
rect 606 1953 612 1954
rect 606 1949 607 1953
rect 611 1949 612 1953
rect 606 1948 612 1949
rect 670 1953 676 1954
rect 670 1949 671 1953
rect 675 1949 676 1953
rect 670 1948 676 1949
rect 734 1953 740 1954
rect 734 1949 735 1953
rect 739 1949 740 1953
rect 734 1948 740 1949
rect 806 1953 812 1954
rect 806 1949 807 1953
rect 811 1949 812 1953
rect 806 1948 812 1949
rect 878 1953 884 1954
rect 878 1949 879 1953
rect 883 1949 884 1953
rect 878 1948 884 1949
rect 950 1953 956 1954
rect 950 1949 951 1953
rect 955 1949 956 1953
rect 950 1948 956 1949
rect 1022 1953 1028 1954
rect 1398 1953 1404 1954
rect 1022 1949 1023 1953
rect 1027 1949 1028 1953
rect 1022 1948 1028 1949
rect 1326 1952 1332 1953
rect 1326 1948 1327 1952
rect 1331 1948 1332 1952
rect 110 1947 116 1948
rect 1326 1947 1332 1948
rect 1366 1952 1372 1953
rect 1366 1948 1367 1952
rect 1371 1948 1372 1952
rect 1398 1949 1399 1953
rect 1403 1949 1404 1953
rect 1398 1948 1404 1949
rect 1454 1953 1460 1954
rect 1454 1949 1455 1953
rect 1459 1949 1460 1953
rect 1454 1948 1460 1949
rect 1518 1953 1524 1954
rect 1518 1949 1519 1953
rect 1523 1949 1524 1953
rect 1518 1948 1524 1949
rect 1598 1953 1604 1954
rect 1598 1949 1599 1953
rect 1603 1949 1604 1953
rect 1598 1948 1604 1949
rect 1678 1953 1684 1954
rect 1678 1949 1679 1953
rect 1683 1949 1684 1953
rect 1678 1948 1684 1949
rect 1758 1953 1764 1954
rect 1758 1949 1759 1953
rect 1763 1949 1764 1953
rect 1758 1948 1764 1949
rect 1854 1953 1860 1954
rect 1854 1949 1855 1953
rect 1859 1949 1860 1953
rect 1854 1948 1860 1949
rect 1966 1953 1972 1954
rect 1966 1949 1967 1953
rect 1971 1949 1972 1953
rect 1966 1948 1972 1949
rect 2094 1953 2100 1954
rect 2094 1949 2095 1953
rect 2099 1949 2100 1953
rect 2094 1948 2100 1949
rect 2238 1953 2244 1954
rect 2238 1949 2239 1953
rect 2243 1949 2244 1953
rect 2238 1948 2244 1949
rect 2390 1953 2396 1954
rect 2390 1949 2391 1953
rect 2395 1949 2396 1953
rect 2390 1948 2396 1949
rect 2526 1953 2532 1954
rect 2526 1949 2527 1953
rect 2531 1949 2532 1953
rect 2526 1948 2532 1949
rect 2582 1952 2588 1953
rect 2582 1948 2583 1952
rect 2587 1948 2588 1952
rect 1366 1947 1372 1948
rect 2582 1947 2588 1948
rect 110 1935 116 1936
rect 110 1931 111 1935
rect 115 1931 116 1935
rect 110 1930 116 1931
rect 1326 1935 1332 1936
rect 1326 1931 1327 1935
rect 1331 1931 1332 1935
rect 1326 1930 1332 1931
rect 1366 1935 1372 1936
rect 1366 1931 1367 1935
rect 1371 1931 1372 1935
rect 1366 1930 1372 1931
rect 2582 1935 2588 1936
rect 2582 1931 2583 1935
rect 2587 1931 2588 1935
rect 2582 1930 2588 1931
rect 398 1926 404 1927
rect 398 1922 399 1926
rect 403 1922 404 1926
rect 398 1921 404 1922
rect 454 1926 460 1927
rect 454 1922 455 1926
rect 459 1922 460 1926
rect 454 1921 460 1922
rect 510 1926 516 1927
rect 510 1922 511 1926
rect 515 1922 516 1926
rect 510 1921 516 1922
rect 566 1926 572 1927
rect 566 1922 567 1926
rect 571 1922 572 1926
rect 566 1921 572 1922
rect 622 1926 628 1927
rect 622 1922 623 1926
rect 627 1922 628 1926
rect 622 1921 628 1922
rect 686 1926 692 1927
rect 686 1922 687 1926
rect 691 1922 692 1926
rect 686 1921 692 1922
rect 750 1926 756 1927
rect 750 1922 751 1926
rect 755 1922 756 1926
rect 750 1921 756 1922
rect 822 1926 828 1927
rect 822 1922 823 1926
rect 827 1922 828 1926
rect 822 1921 828 1922
rect 894 1926 900 1927
rect 894 1922 895 1926
rect 899 1922 900 1926
rect 894 1921 900 1922
rect 966 1926 972 1927
rect 966 1922 967 1926
rect 971 1922 972 1926
rect 966 1921 972 1922
rect 1038 1926 1044 1927
rect 1038 1922 1039 1926
rect 1043 1922 1044 1926
rect 1038 1921 1044 1922
rect 1414 1926 1420 1927
rect 1414 1922 1415 1926
rect 1419 1922 1420 1926
rect 1414 1921 1420 1922
rect 1470 1926 1476 1927
rect 1470 1922 1471 1926
rect 1475 1922 1476 1926
rect 1470 1921 1476 1922
rect 1534 1926 1540 1927
rect 1534 1922 1535 1926
rect 1539 1922 1540 1926
rect 1534 1921 1540 1922
rect 1614 1926 1620 1927
rect 1614 1922 1615 1926
rect 1619 1922 1620 1926
rect 1614 1921 1620 1922
rect 1694 1926 1700 1927
rect 1694 1922 1695 1926
rect 1699 1922 1700 1926
rect 1694 1921 1700 1922
rect 1774 1926 1780 1927
rect 1774 1922 1775 1926
rect 1779 1922 1780 1926
rect 1774 1921 1780 1922
rect 1870 1926 1876 1927
rect 1870 1922 1871 1926
rect 1875 1922 1876 1926
rect 1870 1921 1876 1922
rect 1982 1926 1988 1927
rect 1982 1922 1983 1926
rect 1987 1922 1988 1926
rect 1982 1921 1988 1922
rect 2110 1926 2116 1927
rect 2110 1922 2111 1926
rect 2115 1922 2116 1926
rect 2110 1921 2116 1922
rect 2254 1926 2260 1927
rect 2254 1922 2255 1926
rect 2259 1922 2260 1926
rect 2254 1921 2260 1922
rect 2406 1926 2412 1927
rect 2406 1922 2407 1926
rect 2411 1922 2412 1926
rect 2406 1921 2412 1922
rect 2542 1926 2548 1927
rect 2542 1922 2543 1926
rect 2547 1922 2548 1926
rect 2542 1921 2548 1922
rect 518 1902 524 1903
rect 518 1898 519 1902
rect 523 1898 524 1902
rect 518 1897 524 1898
rect 574 1902 580 1903
rect 574 1898 575 1902
rect 579 1898 580 1902
rect 574 1897 580 1898
rect 630 1902 636 1903
rect 630 1898 631 1902
rect 635 1898 636 1902
rect 630 1897 636 1898
rect 686 1902 692 1903
rect 686 1898 687 1902
rect 691 1898 692 1902
rect 686 1897 692 1898
rect 742 1902 748 1903
rect 742 1898 743 1902
rect 747 1898 748 1902
rect 742 1897 748 1898
rect 806 1902 812 1903
rect 806 1898 807 1902
rect 811 1898 812 1902
rect 806 1897 812 1898
rect 870 1902 876 1903
rect 870 1898 871 1902
rect 875 1898 876 1902
rect 870 1897 876 1898
rect 934 1902 940 1903
rect 934 1898 935 1902
rect 939 1898 940 1902
rect 934 1897 940 1898
rect 998 1902 1004 1903
rect 998 1898 999 1902
rect 1003 1898 1004 1902
rect 998 1897 1004 1898
rect 1574 1902 1580 1903
rect 1574 1898 1575 1902
rect 1579 1898 1580 1902
rect 1574 1897 1580 1898
rect 1630 1902 1636 1903
rect 1630 1898 1631 1902
rect 1635 1898 1636 1902
rect 1630 1897 1636 1898
rect 1686 1902 1692 1903
rect 1686 1898 1687 1902
rect 1691 1898 1692 1902
rect 1686 1897 1692 1898
rect 1742 1902 1748 1903
rect 1742 1898 1743 1902
rect 1747 1898 1748 1902
rect 1742 1897 1748 1898
rect 1798 1902 1804 1903
rect 1798 1898 1799 1902
rect 1803 1898 1804 1902
rect 1798 1897 1804 1898
rect 1854 1902 1860 1903
rect 1854 1898 1855 1902
rect 1859 1898 1860 1902
rect 1854 1897 1860 1898
rect 1926 1902 1932 1903
rect 1926 1898 1927 1902
rect 1931 1898 1932 1902
rect 1926 1897 1932 1898
rect 2014 1902 2020 1903
rect 2014 1898 2015 1902
rect 2019 1898 2020 1902
rect 2014 1897 2020 1898
rect 2126 1902 2132 1903
rect 2126 1898 2127 1902
rect 2131 1898 2132 1902
rect 2126 1897 2132 1898
rect 2246 1902 2252 1903
rect 2246 1898 2247 1902
rect 2251 1898 2252 1902
rect 2246 1897 2252 1898
rect 2382 1902 2388 1903
rect 2382 1898 2383 1902
rect 2387 1898 2388 1902
rect 2382 1897 2388 1898
rect 2518 1902 2524 1903
rect 2518 1898 2519 1902
rect 2523 1898 2524 1902
rect 2518 1897 2524 1898
rect 110 1893 116 1894
rect 110 1889 111 1893
rect 115 1889 116 1893
rect 110 1888 116 1889
rect 1326 1893 1332 1894
rect 1326 1889 1327 1893
rect 1331 1889 1332 1893
rect 1326 1888 1332 1889
rect 1366 1893 1372 1894
rect 1366 1889 1367 1893
rect 1371 1889 1372 1893
rect 1366 1888 1372 1889
rect 2582 1893 2588 1894
rect 2582 1889 2583 1893
rect 2587 1889 2588 1893
rect 2582 1888 2588 1889
rect 110 1876 116 1877
rect 1326 1876 1332 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 502 1875 508 1876
rect 502 1871 503 1875
rect 507 1871 508 1875
rect 502 1870 508 1871
rect 558 1875 564 1876
rect 558 1871 559 1875
rect 563 1871 564 1875
rect 558 1870 564 1871
rect 614 1875 620 1876
rect 614 1871 615 1875
rect 619 1871 620 1875
rect 614 1870 620 1871
rect 670 1875 676 1876
rect 670 1871 671 1875
rect 675 1871 676 1875
rect 670 1870 676 1871
rect 726 1875 732 1876
rect 726 1871 727 1875
rect 731 1871 732 1875
rect 726 1870 732 1871
rect 790 1875 796 1876
rect 790 1871 791 1875
rect 795 1871 796 1875
rect 790 1870 796 1871
rect 854 1875 860 1876
rect 854 1871 855 1875
rect 859 1871 860 1875
rect 854 1870 860 1871
rect 918 1875 924 1876
rect 918 1871 919 1875
rect 923 1871 924 1875
rect 918 1870 924 1871
rect 982 1875 988 1876
rect 982 1871 983 1875
rect 987 1871 988 1875
rect 1326 1872 1327 1876
rect 1331 1872 1332 1876
rect 1326 1871 1332 1872
rect 1366 1876 1372 1877
rect 2582 1876 2588 1877
rect 1366 1872 1367 1876
rect 1371 1872 1372 1876
rect 1366 1871 1372 1872
rect 1558 1875 1564 1876
rect 1558 1871 1559 1875
rect 1563 1871 1564 1875
rect 982 1870 988 1871
rect 1558 1870 1564 1871
rect 1614 1875 1620 1876
rect 1614 1871 1615 1875
rect 1619 1871 1620 1875
rect 1614 1870 1620 1871
rect 1670 1875 1676 1876
rect 1670 1871 1671 1875
rect 1675 1871 1676 1875
rect 1670 1870 1676 1871
rect 1726 1875 1732 1876
rect 1726 1871 1727 1875
rect 1731 1871 1732 1875
rect 1726 1870 1732 1871
rect 1782 1875 1788 1876
rect 1782 1871 1783 1875
rect 1787 1871 1788 1875
rect 1782 1870 1788 1871
rect 1838 1875 1844 1876
rect 1838 1871 1839 1875
rect 1843 1871 1844 1875
rect 1838 1870 1844 1871
rect 1910 1875 1916 1876
rect 1910 1871 1911 1875
rect 1915 1871 1916 1875
rect 1910 1870 1916 1871
rect 1998 1875 2004 1876
rect 1998 1871 1999 1875
rect 2003 1871 2004 1875
rect 1998 1870 2004 1871
rect 2110 1875 2116 1876
rect 2110 1871 2111 1875
rect 2115 1871 2116 1875
rect 2110 1870 2116 1871
rect 2230 1875 2236 1876
rect 2230 1871 2231 1875
rect 2235 1871 2236 1875
rect 2230 1870 2236 1871
rect 2366 1875 2372 1876
rect 2366 1871 2367 1875
rect 2371 1871 2372 1875
rect 2366 1870 2372 1871
rect 2502 1875 2508 1876
rect 2502 1871 2503 1875
rect 2507 1871 2508 1875
rect 2582 1872 2583 1876
rect 2587 1872 2588 1876
rect 2582 1871 2588 1872
rect 2502 1870 2508 1871
rect 142 1837 148 1838
rect 110 1836 116 1837
rect 110 1832 111 1836
rect 115 1832 116 1836
rect 142 1833 143 1837
rect 147 1833 148 1837
rect 142 1832 148 1833
rect 198 1837 204 1838
rect 198 1833 199 1837
rect 203 1833 204 1837
rect 198 1832 204 1833
rect 254 1837 260 1838
rect 254 1833 255 1837
rect 259 1833 260 1837
rect 254 1832 260 1833
rect 310 1837 316 1838
rect 310 1833 311 1837
rect 315 1833 316 1837
rect 310 1832 316 1833
rect 374 1837 380 1838
rect 374 1833 375 1837
rect 379 1833 380 1837
rect 374 1832 380 1833
rect 454 1837 460 1838
rect 454 1833 455 1837
rect 459 1833 460 1837
rect 454 1832 460 1833
rect 542 1837 548 1838
rect 542 1833 543 1837
rect 547 1833 548 1837
rect 542 1832 548 1833
rect 630 1837 636 1838
rect 630 1833 631 1837
rect 635 1833 636 1837
rect 630 1832 636 1833
rect 718 1837 724 1838
rect 718 1833 719 1837
rect 723 1833 724 1837
rect 718 1832 724 1833
rect 798 1837 804 1838
rect 798 1833 799 1837
rect 803 1833 804 1837
rect 798 1832 804 1833
rect 886 1837 892 1838
rect 886 1833 887 1837
rect 891 1833 892 1837
rect 886 1832 892 1833
rect 974 1837 980 1838
rect 974 1833 975 1837
rect 979 1833 980 1837
rect 974 1832 980 1833
rect 1062 1837 1068 1838
rect 1062 1833 1063 1837
rect 1067 1833 1068 1837
rect 1062 1832 1068 1833
rect 1326 1836 1332 1837
rect 1326 1832 1327 1836
rect 1331 1832 1332 1836
rect 1622 1833 1628 1834
rect 110 1831 116 1832
rect 1326 1831 1332 1832
rect 1366 1832 1372 1833
rect 1366 1828 1367 1832
rect 1371 1828 1372 1832
rect 1622 1829 1623 1833
rect 1627 1829 1628 1833
rect 1622 1828 1628 1829
rect 1678 1833 1684 1834
rect 1678 1829 1679 1833
rect 1683 1829 1684 1833
rect 1678 1828 1684 1829
rect 1734 1833 1740 1834
rect 1734 1829 1735 1833
rect 1739 1829 1740 1833
rect 1734 1828 1740 1829
rect 1790 1833 1796 1834
rect 1790 1829 1791 1833
rect 1795 1829 1796 1833
rect 1790 1828 1796 1829
rect 1846 1833 1852 1834
rect 1846 1829 1847 1833
rect 1851 1829 1852 1833
rect 1846 1828 1852 1829
rect 1902 1833 1908 1834
rect 1902 1829 1903 1833
rect 1907 1829 1908 1833
rect 1902 1828 1908 1829
rect 1966 1833 1972 1834
rect 1966 1829 1967 1833
rect 1971 1829 1972 1833
rect 1966 1828 1972 1829
rect 2038 1833 2044 1834
rect 2038 1829 2039 1833
rect 2043 1829 2044 1833
rect 2038 1828 2044 1829
rect 2126 1833 2132 1834
rect 2126 1829 2127 1833
rect 2131 1829 2132 1833
rect 2126 1828 2132 1829
rect 2222 1833 2228 1834
rect 2222 1829 2223 1833
rect 2227 1829 2228 1833
rect 2222 1828 2228 1829
rect 2326 1833 2332 1834
rect 2326 1829 2327 1833
rect 2331 1829 2332 1833
rect 2326 1828 2332 1829
rect 2438 1833 2444 1834
rect 2438 1829 2439 1833
rect 2443 1829 2444 1833
rect 2438 1828 2444 1829
rect 2526 1833 2532 1834
rect 2526 1829 2527 1833
rect 2531 1829 2532 1833
rect 2526 1828 2532 1829
rect 2582 1832 2588 1833
rect 2582 1828 2583 1832
rect 2587 1828 2588 1832
rect 1366 1827 1372 1828
rect 2582 1827 2588 1828
rect 110 1819 116 1820
rect 110 1815 111 1819
rect 115 1815 116 1819
rect 110 1814 116 1815
rect 1326 1819 1332 1820
rect 1326 1815 1327 1819
rect 1331 1815 1332 1819
rect 1326 1814 1332 1815
rect 1366 1815 1372 1816
rect 1366 1811 1367 1815
rect 1371 1811 1372 1815
rect 158 1810 164 1811
rect 158 1806 159 1810
rect 163 1806 164 1810
rect 158 1805 164 1806
rect 214 1810 220 1811
rect 214 1806 215 1810
rect 219 1806 220 1810
rect 214 1805 220 1806
rect 270 1810 276 1811
rect 270 1806 271 1810
rect 275 1806 276 1810
rect 270 1805 276 1806
rect 326 1810 332 1811
rect 326 1806 327 1810
rect 331 1806 332 1810
rect 326 1805 332 1806
rect 390 1810 396 1811
rect 390 1806 391 1810
rect 395 1806 396 1810
rect 390 1805 396 1806
rect 470 1810 476 1811
rect 470 1806 471 1810
rect 475 1806 476 1810
rect 470 1805 476 1806
rect 558 1810 564 1811
rect 558 1806 559 1810
rect 563 1806 564 1810
rect 558 1805 564 1806
rect 646 1810 652 1811
rect 646 1806 647 1810
rect 651 1806 652 1810
rect 646 1805 652 1806
rect 734 1810 740 1811
rect 734 1806 735 1810
rect 739 1806 740 1810
rect 734 1805 740 1806
rect 814 1810 820 1811
rect 814 1806 815 1810
rect 819 1806 820 1810
rect 814 1805 820 1806
rect 902 1810 908 1811
rect 902 1806 903 1810
rect 907 1806 908 1810
rect 902 1805 908 1806
rect 990 1810 996 1811
rect 990 1806 991 1810
rect 995 1806 996 1810
rect 990 1805 996 1806
rect 1078 1810 1084 1811
rect 1366 1810 1372 1811
rect 2582 1815 2588 1816
rect 2582 1811 2583 1815
rect 2587 1811 2588 1815
rect 2582 1810 2588 1811
rect 1078 1806 1079 1810
rect 1083 1806 1084 1810
rect 1078 1805 1084 1806
rect 1638 1806 1644 1807
rect 1638 1802 1639 1806
rect 1643 1802 1644 1806
rect 1638 1801 1644 1802
rect 1694 1806 1700 1807
rect 1694 1802 1695 1806
rect 1699 1802 1700 1806
rect 1694 1801 1700 1802
rect 1750 1806 1756 1807
rect 1750 1802 1751 1806
rect 1755 1802 1756 1806
rect 1750 1801 1756 1802
rect 1806 1806 1812 1807
rect 1806 1802 1807 1806
rect 1811 1802 1812 1806
rect 1806 1801 1812 1802
rect 1862 1806 1868 1807
rect 1862 1802 1863 1806
rect 1867 1802 1868 1806
rect 1862 1801 1868 1802
rect 1918 1806 1924 1807
rect 1918 1802 1919 1806
rect 1923 1802 1924 1806
rect 1918 1801 1924 1802
rect 1982 1806 1988 1807
rect 1982 1802 1983 1806
rect 1987 1802 1988 1806
rect 1982 1801 1988 1802
rect 2054 1806 2060 1807
rect 2054 1802 2055 1806
rect 2059 1802 2060 1806
rect 2054 1801 2060 1802
rect 2142 1806 2148 1807
rect 2142 1802 2143 1806
rect 2147 1802 2148 1806
rect 2142 1801 2148 1802
rect 2238 1806 2244 1807
rect 2238 1802 2239 1806
rect 2243 1802 2244 1806
rect 2238 1801 2244 1802
rect 2342 1806 2348 1807
rect 2342 1802 2343 1806
rect 2347 1802 2348 1806
rect 2342 1801 2348 1802
rect 2454 1806 2460 1807
rect 2454 1802 2455 1806
rect 2459 1802 2460 1806
rect 2454 1801 2460 1802
rect 2542 1806 2548 1807
rect 2542 1802 2543 1806
rect 2547 1802 2548 1806
rect 2542 1801 2548 1802
rect 158 1778 164 1779
rect 158 1774 159 1778
rect 163 1774 164 1778
rect 158 1773 164 1774
rect 254 1778 260 1779
rect 254 1774 255 1778
rect 259 1774 260 1778
rect 254 1773 260 1774
rect 374 1778 380 1779
rect 374 1774 375 1778
rect 379 1774 380 1778
rect 374 1773 380 1774
rect 502 1778 508 1779
rect 502 1774 503 1778
rect 507 1774 508 1778
rect 502 1773 508 1774
rect 622 1778 628 1779
rect 622 1774 623 1778
rect 627 1774 628 1778
rect 622 1773 628 1774
rect 742 1778 748 1779
rect 742 1774 743 1778
rect 747 1774 748 1778
rect 742 1773 748 1774
rect 854 1778 860 1779
rect 854 1774 855 1778
rect 859 1774 860 1778
rect 854 1773 860 1774
rect 958 1778 964 1779
rect 958 1774 959 1778
rect 963 1774 964 1778
rect 958 1773 964 1774
rect 1054 1778 1060 1779
rect 1054 1774 1055 1778
rect 1059 1774 1060 1778
rect 1054 1773 1060 1774
rect 1150 1778 1156 1779
rect 1150 1774 1151 1778
rect 1155 1774 1156 1778
rect 1150 1773 1156 1774
rect 1246 1778 1252 1779
rect 1246 1774 1247 1778
rect 1251 1774 1252 1778
rect 1246 1773 1252 1774
rect 1470 1774 1476 1775
rect 1470 1770 1471 1774
rect 1475 1770 1476 1774
rect 110 1769 116 1770
rect 110 1765 111 1769
rect 115 1765 116 1769
rect 110 1764 116 1765
rect 1326 1769 1332 1770
rect 1470 1769 1476 1770
rect 1534 1774 1540 1775
rect 1534 1770 1535 1774
rect 1539 1770 1540 1774
rect 1534 1769 1540 1770
rect 1614 1774 1620 1775
rect 1614 1770 1615 1774
rect 1619 1770 1620 1774
rect 1614 1769 1620 1770
rect 1694 1774 1700 1775
rect 1694 1770 1695 1774
rect 1699 1770 1700 1774
rect 1694 1769 1700 1770
rect 1782 1774 1788 1775
rect 1782 1770 1783 1774
rect 1787 1770 1788 1774
rect 1782 1769 1788 1770
rect 1878 1774 1884 1775
rect 1878 1770 1879 1774
rect 1883 1770 1884 1774
rect 1878 1769 1884 1770
rect 1974 1774 1980 1775
rect 1974 1770 1975 1774
rect 1979 1770 1980 1774
rect 1974 1769 1980 1770
rect 2070 1774 2076 1775
rect 2070 1770 2071 1774
rect 2075 1770 2076 1774
rect 2070 1769 2076 1770
rect 2166 1774 2172 1775
rect 2166 1770 2167 1774
rect 2171 1770 2172 1774
rect 2166 1769 2172 1770
rect 2262 1774 2268 1775
rect 2262 1770 2263 1774
rect 2267 1770 2268 1774
rect 2262 1769 2268 1770
rect 2358 1774 2364 1775
rect 2358 1770 2359 1774
rect 2363 1770 2364 1774
rect 2358 1769 2364 1770
rect 2462 1774 2468 1775
rect 2462 1770 2463 1774
rect 2467 1770 2468 1774
rect 2462 1769 2468 1770
rect 2542 1774 2548 1775
rect 2542 1770 2543 1774
rect 2547 1770 2548 1774
rect 2542 1769 2548 1770
rect 1326 1765 1327 1769
rect 1331 1765 1332 1769
rect 1326 1764 1332 1765
rect 1366 1765 1372 1766
rect 1366 1761 1367 1765
rect 1371 1761 1372 1765
rect 1366 1760 1372 1761
rect 2582 1765 2588 1766
rect 2582 1761 2583 1765
rect 2587 1761 2588 1765
rect 2582 1760 2588 1761
rect 110 1752 116 1753
rect 1326 1752 1332 1753
rect 110 1748 111 1752
rect 115 1748 116 1752
rect 110 1747 116 1748
rect 142 1751 148 1752
rect 142 1747 143 1751
rect 147 1747 148 1751
rect 142 1746 148 1747
rect 238 1751 244 1752
rect 238 1747 239 1751
rect 243 1747 244 1751
rect 238 1746 244 1747
rect 358 1751 364 1752
rect 358 1747 359 1751
rect 363 1747 364 1751
rect 358 1746 364 1747
rect 486 1751 492 1752
rect 486 1747 487 1751
rect 491 1747 492 1751
rect 486 1746 492 1747
rect 606 1751 612 1752
rect 606 1747 607 1751
rect 611 1747 612 1751
rect 606 1746 612 1747
rect 726 1751 732 1752
rect 726 1747 727 1751
rect 731 1747 732 1751
rect 726 1746 732 1747
rect 838 1751 844 1752
rect 838 1747 839 1751
rect 843 1747 844 1751
rect 838 1746 844 1747
rect 942 1751 948 1752
rect 942 1747 943 1751
rect 947 1747 948 1751
rect 942 1746 948 1747
rect 1038 1751 1044 1752
rect 1038 1747 1039 1751
rect 1043 1747 1044 1751
rect 1038 1746 1044 1747
rect 1134 1751 1140 1752
rect 1134 1747 1135 1751
rect 1139 1747 1140 1751
rect 1134 1746 1140 1747
rect 1230 1751 1236 1752
rect 1230 1747 1231 1751
rect 1235 1747 1236 1751
rect 1326 1748 1327 1752
rect 1331 1748 1332 1752
rect 1326 1747 1332 1748
rect 1366 1748 1372 1749
rect 2582 1748 2588 1749
rect 1230 1746 1236 1747
rect 1366 1744 1367 1748
rect 1371 1744 1372 1748
rect 1366 1743 1372 1744
rect 1454 1747 1460 1748
rect 1454 1743 1455 1747
rect 1459 1743 1460 1747
rect 1454 1742 1460 1743
rect 1518 1747 1524 1748
rect 1518 1743 1519 1747
rect 1523 1743 1524 1747
rect 1518 1742 1524 1743
rect 1598 1747 1604 1748
rect 1598 1743 1599 1747
rect 1603 1743 1604 1747
rect 1598 1742 1604 1743
rect 1678 1747 1684 1748
rect 1678 1743 1679 1747
rect 1683 1743 1684 1747
rect 1678 1742 1684 1743
rect 1766 1747 1772 1748
rect 1766 1743 1767 1747
rect 1771 1743 1772 1747
rect 1766 1742 1772 1743
rect 1862 1747 1868 1748
rect 1862 1743 1863 1747
rect 1867 1743 1868 1747
rect 1862 1742 1868 1743
rect 1958 1747 1964 1748
rect 1958 1743 1959 1747
rect 1963 1743 1964 1747
rect 1958 1742 1964 1743
rect 2054 1747 2060 1748
rect 2054 1743 2055 1747
rect 2059 1743 2060 1747
rect 2054 1742 2060 1743
rect 2150 1747 2156 1748
rect 2150 1743 2151 1747
rect 2155 1743 2156 1747
rect 2150 1742 2156 1743
rect 2246 1747 2252 1748
rect 2246 1743 2247 1747
rect 2251 1743 2252 1747
rect 2246 1742 2252 1743
rect 2342 1747 2348 1748
rect 2342 1743 2343 1747
rect 2347 1743 2348 1747
rect 2342 1742 2348 1743
rect 2446 1747 2452 1748
rect 2446 1743 2447 1747
rect 2451 1743 2452 1747
rect 2446 1742 2452 1743
rect 2526 1747 2532 1748
rect 2526 1743 2527 1747
rect 2531 1743 2532 1747
rect 2582 1744 2583 1748
rect 2587 1744 2588 1748
rect 2582 1743 2588 1744
rect 2526 1742 2532 1743
rect 142 1717 148 1718
rect 110 1716 116 1717
rect 110 1712 111 1716
rect 115 1712 116 1716
rect 142 1713 143 1717
rect 147 1713 148 1717
rect 142 1712 148 1713
rect 262 1717 268 1718
rect 262 1713 263 1717
rect 267 1713 268 1717
rect 262 1712 268 1713
rect 414 1717 420 1718
rect 414 1713 415 1717
rect 419 1713 420 1717
rect 414 1712 420 1713
rect 566 1717 572 1718
rect 566 1713 567 1717
rect 571 1713 572 1717
rect 566 1712 572 1713
rect 710 1717 716 1718
rect 710 1713 711 1717
rect 715 1713 716 1717
rect 710 1712 716 1713
rect 854 1717 860 1718
rect 854 1713 855 1717
rect 859 1713 860 1717
rect 854 1712 860 1713
rect 998 1717 1004 1718
rect 998 1713 999 1717
rect 1003 1713 1004 1717
rect 998 1712 1004 1713
rect 1142 1717 1148 1718
rect 1142 1713 1143 1717
rect 1147 1713 1148 1717
rect 1142 1712 1148 1713
rect 1270 1717 1276 1718
rect 1270 1713 1271 1717
rect 1275 1713 1276 1717
rect 1270 1712 1276 1713
rect 1326 1716 1332 1717
rect 1326 1712 1327 1716
rect 1331 1712 1332 1716
rect 110 1711 116 1712
rect 1326 1711 1332 1712
rect 1398 1709 1404 1710
rect 1366 1708 1372 1709
rect 1366 1704 1367 1708
rect 1371 1704 1372 1708
rect 1398 1705 1399 1709
rect 1403 1705 1404 1709
rect 1398 1704 1404 1705
rect 1478 1709 1484 1710
rect 1478 1705 1479 1709
rect 1483 1705 1484 1709
rect 1478 1704 1484 1705
rect 1598 1709 1604 1710
rect 1598 1705 1599 1709
rect 1603 1705 1604 1709
rect 1598 1704 1604 1705
rect 1718 1709 1724 1710
rect 1718 1705 1719 1709
rect 1723 1705 1724 1709
rect 1718 1704 1724 1705
rect 1838 1709 1844 1710
rect 1838 1705 1839 1709
rect 1843 1705 1844 1709
rect 1838 1704 1844 1705
rect 1950 1709 1956 1710
rect 1950 1705 1951 1709
rect 1955 1705 1956 1709
rect 1950 1704 1956 1705
rect 2054 1709 2060 1710
rect 2054 1705 2055 1709
rect 2059 1705 2060 1709
rect 2054 1704 2060 1705
rect 2158 1709 2164 1710
rect 2158 1705 2159 1709
rect 2163 1705 2164 1709
rect 2158 1704 2164 1705
rect 2254 1709 2260 1710
rect 2254 1705 2255 1709
rect 2259 1705 2260 1709
rect 2254 1704 2260 1705
rect 2350 1709 2356 1710
rect 2350 1705 2351 1709
rect 2355 1705 2356 1709
rect 2350 1704 2356 1705
rect 2446 1709 2452 1710
rect 2446 1705 2447 1709
rect 2451 1705 2452 1709
rect 2446 1704 2452 1705
rect 2526 1709 2532 1710
rect 2526 1705 2527 1709
rect 2531 1705 2532 1709
rect 2526 1704 2532 1705
rect 2582 1708 2588 1709
rect 2582 1704 2583 1708
rect 2587 1704 2588 1708
rect 1366 1703 1372 1704
rect 2582 1703 2588 1704
rect 110 1699 116 1700
rect 110 1695 111 1699
rect 115 1695 116 1699
rect 110 1694 116 1695
rect 1326 1699 1332 1700
rect 1326 1695 1327 1699
rect 1331 1695 1332 1699
rect 1326 1694 1332 1695
rect 1366 1691 1372 1692
rect 158 1690 164 1691
rect 158 1686 159 1690
rect 163 1686 164 1690
rect 158 1685 164 1686
rect 278 1690 284 1691
rect 278 1686 279 1690
rect 283 1686 284 1690
rect 278 1685 284 1686
rect 430 1690 436 1691
rect 430 1686 431 1690
rect 435 1686 436 1690
rect 430 1685 436 1686
rect 582 1690 588 1691
rect 582 1686 583 1690
rect 587 1686 588 1690
rect 582 1685 588 1686
rect 726 1690 732 1691
rect 726 1686 727 1690
rect 731 1686 732 1690
rect 726 1685 732 1686
rect 870 1690 876 1691
rect 870 1686 871 1690
rect 875 1686 876 1690
rect 870 1685 876 1686
rect 1014 1690 1020 1691
rect 1014 1686 1015 1690
rect 1019 1686 1020 1690
rect 1014 1685 1020 1686
rect 1158 1690 1164 1691
rect 1158 1686 1159 1690
rect 1163 1686 1164 1690
rect 1158 1685 1164 1686
rect 1286 1690 1292 1691
rect 1286 1686 1287 1690
rect 1291 1686 1292 1690
rect 1366 1687 1367 1691
rect 1371 1687 1372 1691
rect 1366 1686 1372 1687
rect 2582 1691 2588 1692
rect 2582 1687 2583 1691
rect 2587 1687 2588 1691
rect 2582 1686 2588 1687
rect 1286 1685 1292 1686
rect 1414 1682 1420 1683
rect 1414 1678 1415 1682
rect 1419 1678 1420 1682
rect 1414 1677 1420 1678
rect 1494 1682 1500 1683
rect 1494 1678 1495 1682
rect 1499 1678 1500 1682
rect 1494 1677 1500 1678
rect 1614 1682 1620 1683
rect 1614 1678 1615 1682
rect 1619 1678 1620 1682
rect 1614 1677 1620 1678
rect 1734 1682 1740 1683
rect 1734 1678 1735 1682
rect 1739 1678 1740 1682
rect 1734 1677 1740 1678
rect 1854 1682 1860 1683
rect 1854 1678 1855 1682
rect 1859 1678 1860 1682
rect 1854 1677 1860 1678
rect 1966 1682 1972 1683
rect 1966 1678 1967 1682
rect 1971 1678 1972 1682
rect 1966 1677 1972 1678
rect 2070 1682 2076 1683
rect 2070 1678 2071 1682
rect 2075 1678 2076 1682
rect 2070 1677 2076 1678
rect 2174 1682 2180 1683
rect 2174 1678 2175 1682
rect 2179 1678 2180 1682
rect 2174 1677 2180 1678
rect 2270 1682 2276 1683
rect 2270 1678 2271 1682
rect 2275 1678 2276 1682
rect 2270 1677 2276 1678
rect 2366 1682 2372 1683
rect 2366 1678 2367 1682
rect 2371 1678 2372 1682
rect 2366 1677 2372 1678
rect 2462 1682 2468 1683
rect 2462 1678 2463 1682
rect 2467 1678 2468 1682
rect 2462 1677 2468 1678
rect 2542 1682 2548 1683
rect 2542 1678 2543 1682
rect 2547 1678 2548 1682
rect 2542 1677 2548 1678
rect 158 1662 164 1663
rect 158 1658 159 1662
rect 163 1658 164 1662
rect 158 1657 164 1658
rect 222 1662 228 1663
rect 222 1658 223 1662
rect 227 1658 228 1662
rect 222 1657 228 1658
rect 302 1662 308 1663
rect 302 1658 303 1662
rect 307 1658 308 1662
rect 302 1657 308 1658
rect 382 1662 388 1663
rect 382 1658 383 1662
rect 387 1658 388 1662
rect 382 1657 388 1658
rect 462 1662 468 1663
rect 462 1658 463 1662
rect 467 1658 468 1662
rect 462 1657 468 1658
rect 534 1662 540 1663
rect 534 1658 535 1662
rect 539 1658 540 1662
rect 534 1657 540 1658
rect 606 1662 612 1663
rect 606 1658 607 1662
rect 611 1658 612 1662
rect 606 1657 612 1658
rect 678 1662 684 1663
rect 678 1658 679 1662
rect 683 1658 684 1662
rect 678 1657 684 1658
rect 766 1662 772 1663
rect 766 1658 767 1662
rect 771 1658 772 1662
rect 766 1657 772 1658
rect 862 1662 868 1663
rect 862 1658 863 1662
rect 867 1658 868 1662
rect 862 1657 868 1658
rect 966 1662 972 1663
rect 966 1658 967 1662
rect 971 1658 972 1662
rect 966 1657 972 1658
rect 1078 1662 1084 1663
rect 1078 1658 1079 1662
rect 1083 1658 1084 1662
rect 1078 1657 1084 1658
rect 1190 1662 1196 1663
rect 1190 1658 1191 1662
rect 1195 1658 1196 1662
rect 1190 1657 1196 1658
rect 1286 1662 1292 1663
rect 1286 1658 1287 1662
rect 1291 1658 1292 1662
rect 1286 1657 1292 1658
rect 1414 1658 1420 1659
rect 1414 1654 1415 1658
rect 1419 1654 1420 1658
rect 110 1653 116 1654
rect 110 1649 111 1653
rect 115 1649 116 1653
rect 110 1648 116 1649
rect 1326 1653 1332 1654
rect 1414 1653 1420 1654
rect 1502 1658 1508 1659
rect 1502 1654 1503 1658
rect 1507 1654 1508 1658
rect 1502 1653 1508 1654
rect 1622 1658 1628 1659
rect 1622 1654 1623 1658
rect 1627 1654 1628 1658
rect 1622 1653 1628 1654
rect 1750 1658 1756 1659
rect 1750 1654 1751 1658
rect 1755 1654 1756 1658
rect 1750 1653 1756 1654
rect 1878 1658 1884 1659
rect 1878 1654 1879 1658
rect 1883 1654 1884 1658
rect 1878 1653 1884 1654
rect 1998 1658 2004 1659
rect 1998 1654 1999 1658
rect 2003 1654 2004 1658
rect 1998 1653 2004 1654
rect 2118 1658 2124 1659
rect 2118 1654 2119 1658
rect 2123 1654 2124 1658
rect 2118 1653 2124 1654
rect 2230 1658 2236 1659
rect 2230 1654 2231 1658
rect 2235 1654 2236 1658
rect 2230 1653 2236 1654
rect 2342 1658 2348 1659
rect 2342 1654 2343 1658
rect 2347 1654 2348 1658
rect 2342 1653 2348 1654
rect 2454 1658 2460 1659
rect 2454 1654 2455 1658
rect 2459 1654 2460 1658
rect 2454 1653 2460 1654
rect 2542 1658 2548 1659
rect 2542 1654 2543 1658
rect 2547 1654 2548 1658
rect 2542 1653 2548 1654
rect 1326 1649 1327 1653
rect 1331 1649 1332 1653
rect 1326 1648 1332 1649
rect 1366 1649 1372 1650
rect 1366 1645 1367 1649
rect 1371 1645 1372 1649
rect 1366 1644 1372 1645
rect 2582 1649 2588 1650
rect 2582 1645 2583 1649
rect 2587 1645 2588 1649
rect 2582 1644 2588 1645
rect 110 1636 116 1637
rect 1326 1636 1332 1637
rect 110 1632 111 1636
rect 115 1632 116 1636
rect 110 1631 116 1632
rect 142 1635 148 1636
rect 142 1631 143 1635
rect 147 1631 148 1635
rect 142 1630 148 1631
rect 206 1635 212 1636
rect 206 1631 207 1635
rect 211 1631 212 1635
rect 206 1630 212 1631
rect 286 1635 292 1636
rect 286 1631 287 1635
rect 291 1631 292 1635
rect 286 1630 292 1631
rect 366 1635 372 1636
rect 366 1631 367 1635
rect 371 1631 372 1635
rect 366 1630 372 1631
rect 446 1635 452 1636
rect 446 1631 447 1635
rect 451 1631 452 1635
rect 446 1630 452 1631
rect 518 1635 524 1636
rect 518 1631 519 1635
rect 523 1631 524 1635
rect 518 1630 524 1631
rect 590 1635 596 1636
rect 590 1631 591 1635
rect 595 1631 596 1635
rect 590 1630 596 1631
rect 662 1635 668 1636
rect 662 1631 663 1635
rect 667 1631 668 1635
rect 662 1630 668 1631
rect 750 1635 756 1636
rect 750 1631 751 1635
rect 755 1631 756 1635
rect 750 1630 756 1631
rect 846 1635 852 1636
rect 846 1631 847 1635
rect 851 1631 852 1635
rect 846 1630 852 1631
rect 950 1635 956 1636
rect 950 1631 951 1635
rect 955 1631 956 1635
rect 950 1630 956 1631
rect 1062 1635 1068 1636
rect 1062 1631 1063 1635
rect 1067 1631 1068 1635
rect 1062 1630 1068 1631
rect 1174 1635 1180 1636
rect 1174 1631 1175 1635
rect 1179 1631 1180 1635
rect 1174 1630 1180 1631
rect 1270 1635 1276 1636
rect 1270 1631 1271 1635
rect 1275 1631 1276 1635
rect 1326 1632 1327 1636
rect 1331 1632 1332 1636
rect 1326 1631 1332 1632
rect 1366 1632 1372 1633
rect 2582 1632 2588 1633
rect 1270 1630 1276 1631
rect 1366 1628 1367 1632
rect 1371 1628 1372 1632
rect 1366 1627 1372 1628
rect 1398 1631 1404 1632
rect 1398 1627 1399 1631
rect 1403 1627 1404 1631
rect 1398 1626 1404 1627
rect 1486 1631 1492 1632
rect 1486 1627 1487 1631
rect 1491 1627 1492 1631
rect 1486 1626 1492 1627
rect 1606 1631 1612 1632
rect 1606 1627 1607 1631
rect 1611 1627 1612 1631
rect 1606 1626 1612 1627
rect 1734 1631 1740 1632
rect 1734 1627 1735 1631
rect 1739 1627 1740 1631
rect 1734 1626 1740 1627
rect 1862 1631 1868 1632
rect 1862 1627 1863 1631
rect 1867 1627 1868 1631
rect 1862 1626 1868 1627
rect 1982 1631 1988 1632
rect 1982 1627 1983 1631
rect 1987 1627 1988 1631
rect 1982 1626 1988 1627
rect 2102 1631 2108 1632
rect 2102 1627 2103 1631
rect 2107 1627 2108 1631
rect 2102 1626 2108 1627
rect 2214 1631 2220 1632
rect 2214 1627 2215 1631
rect 2219 1627 2220 1631
rect 2214 1626 2220 1627
rect 2326 1631 2332 1632
rect 2326 1627 2327 1631
rect 2331 1627 2332 1631
rect 2326 1626 2332 1627
rect 2438 1631 2444 1632
rect 2438 1627 2439 1631
rect 2443 1627 2444 1631
rect 2438 1626 2444 1627
rect 2526 1631 2532 1632
rect 2526 1627 2527 1631
rect 2531 1627 2532 1631
rect 2582 1628 2583 1632
rect 2587 1628 2588 1632
rect 2582 1627 2588 1628
rect 2526 1626 2532 1627
rect 142 1601 148 1602
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 142 1597 143 1601
rect 147 1597 148 1601
rect 142 1596 148 1597
rect 246 1601 252 1602
rect 246 1597 247 1601
rect 251 1597 252 1601
rect 246 1596 252 1597
rect 366 1601 372 1602
rect 366 1597 367 1601
rect 371 1597 372 1601
rect 366 1596 372 1597
rect 478 1601 484 1602
rect 478 1597 479 1601
rect 483 1597 484 1601
rect 478 1596 484 1597
rect 574 1601 580 1602
rect 574 1597 575 1601
rect 579 1597 580 1601
rect 574 1596 580 1597
rect 670 1601 676 1602
rect 670 1597 671 1601
rect 675 1597 676 1601
rect 670 1596 676 1597
rect 766 1601 772 1602
rect 766 1597 767 1601
rect 771 1597 772 1601
rect 766 1596 772 1597
rect 862 1601 868 1602
rect 862 1597 863 1601
rect 867 1597 868 1601
rect 862 1596 868 1597
rect 958 1601 964 1602
rect 958 1597 959 1601
rect 963 1597 964 1601
rect 958 1596 964 1597
rect 1062 1601 1068 1602
rect 1062 1597 1063 1601
rect 1067 1597 1068 1601
rect 1062 1596 1068 1597
rect 1174 1601 1180 1602
rect 1174 1597 1175 1601
rect 1179 1597 1180 1601
rect 1174 1596 1180 1597
rect 1270 1601 1276 1602
rect 1270 1597 1271 1601
rect 1275 1597 1276 1601
rect 1270 1596 1276 1597
rect 1326 1600 1332 1601
rect 1326 1596 1327 1600
rect 1331 1596 1332 1600
rect 110 1595 116 1596
rect 1326 1595 1332 1596
rect 1398 1585 1404 1586
rect 1366 1584 1372 1585
rect 110 1583 116 1584
rect 110 1579 111 1583
rect 115 1579 116 1583
rect 110 1578 116 1579
rect 1326 1583 1332 1584
rect 1326 1579 1327 1583
rect 1331 1579 1332 1583
rect 1366 1580 1367 1584
rect 1371 1580 1372 1584
rect 1398 1581 1399 1585
rect 1403 1581 1404 1585
rect 1398 1580 1404 1581
rect 1494 1585 1500 1586
rect 1494 1581 1495 1585
rect 1499 1581 1500 1585
rect 1494 1580 1500 1581
rect 1614 1585 1620 1586
rect 1614 1581 1615 1585
rect 1619 1581 1620 1585
rect 1614 1580 1620 1581
rect 1742 1585 1748 1586
rect 1742 1581 1743 1585
rect 1747 1581 1748 1585
rect 1742 1580 1748 1581
rect 1862 1585 1868 1586
rect 1862 1581 1863 1585
rect 1867 1581 1868 1585
rect 1862 1580 1868 1581
rect 1982 1585 1988 1586
rect 1982 1581 1983 1585
rect 1987 1581 1988 1585
rect 1982 1580 1988 1581
rect 2094 1585 2100 1586
rect 2094 1581 2095 1585
rect 2099 1581 2100 1585
rect 2094 1580 2100 1581
rect 2198 1585 2204 1586
rect 2198 1581 2199 1585
rect 2203 1581 2204 1585
rect 2198 1580 2204 1581
rect 2294 1585 2300 1586
rect 2294 1581 2295 1585
rect 2299 1581 2300 1585
rect 2294 1580 2300 1581
rect 2390 1585 2396 1586
rect 2390 1581 2391 1585
rect 2395 1581 2396 1585
rect 2390 1580 2396 1581
rect 2494 1585 2500 1586
rect 2494 1581 2495 1585
rect 2499 1581 2500 1585
rect 2494 1580 2500 1581
rect 2582 1584 2588 1585
rect 2582 1580 2583 1584
rect 2587 1580 2588 1584
rect 1366 1579 1372 1580
rect 2582 1579 2588 1580
rect 1326 1578 1332 1579
rect 158 1574 164 1575
rect 158 1570 159 1574
rect 163 1570 164 1574
rect 158 1569 164 1570
rect 262 1574 268 1575
rect 262 1570 263 1574
rect 267 1570 268 1574
rect 262 1569 268 1570
rect 382 1574 388 1575
rect 382 1570 383 1574
rect 387 1570 388 1574
rect 382 1569 388 1570
rect 494 1574 500 1575
rect 494 1570 495 1574
rect 499 1570 500 1574
rect 494 1569 500 1570
rect 590 1574 596 1575
rect 590 1570 591 1574
rect 595 1570 596 1574
rect 590 1569 596 1570
rect 686 1574 692 1575
rect 686 1570 687 1574
rect 691 1570 692 1574
rect 686 1569 692 1570
rect 782 1574 788 1575
rect 782 1570 783 1574
rect 787 1570 788 1574
rect 782 1569 788 1570
rect 878 1574 884 1575
rect 878 1570 879 1574
rect 883 1570 884 1574
rect 878 1569 884 1570
rect 974 1574 980 1575
rect 974 1570 975 1574
rect 979 1570 980 1574
rect 974 1569 980 1570
rect 1078 1574 1084 1575
rect 1078 1570 1079 1574
rect 1083 1570 1084 1574
rect 1078 1569 1084 1570
rect 1190 1574 1196 1575
rect 1190 1570 1191 1574
rect 1195 1570 1196 1574
rect 1190 1569 1196 1570
rect 1286 1574 1292 1575
rect 1286 1570 1287 1574
rect 1291 1570 1292 1574
rect 1286 1569 1292 1570
rect 1366 1567 1372 1568
rect 1366 1563 1367 1567
rect 1371 1563 1372 1567
rect 1366 1562 1372 1563
rect 2582 1567 2588 1568
rect 2582 1563 2583 1567
rect 2587 1563 2588 1567
rect 2582 1562 2588 1563
rect 1414 1558 1420 1559
rect 1414 1554 1415 1558
rect 1419 1554 1420 1558
rect 1414 1553 1420 1554
rect 1510 1558 1516 1559
rect 1510 1554 1511 1558
rect 1515 1554 1516 1558
rect 1510 1553 1516 1554
rect 1630 1558 1636 1559
rect 1630 1554 1631 1558
rect 1635 1554 1636 1558
rect 1630 1553 1636 1554
rect 1758 1558 1764 1559
rect 1758 1554 1759 1558
rect 1763 1554 1764 1558
rect 1758 1553 1764 1554
rect 1878 1558 1884 1559
rect 1878 1554 1879 1558
rect 1883 1554 1884 1558
rect 1878 1553 1884 1554
rect 1998 1558 2004 1559
rect 1998 1554 1999 1558
rect 2003 1554 2004 1558
rect 1998 1553 2004 1554
rect 2110 1558 2116 1559
rect 2110 1554 2111 1558
rect 2115 1554 2116 1558
rect 2110 1553 2116 1554
rect 2214 1558 2220 1559
rect 2214 1554 2215 1558
rect 2219 1554 2220 1558
rect 2214 1553 2220 1554
rect 2310 1558 2316 1559
rect 2310 1554 2311 1558
rect 2315 1554 2316 1558
rect 2310 1553 2316 1554
rect 2406 1558 2412 1559
rect 2406 1554 2407 1558
rect 2411 1554 2412 1558
rect 2406 1553 2412 1554
rect 2510 1558 2516 1559
rect 2510 1554 2511 1558
rect 2515 1554 2516 1558
rect 2510 1553 2516 1554
rect 158 1546 164 1547
rect 158 1542 159 1546
rect 163 1542 164 1546
rect 158 1541 164 1542
rect 230 1546 236 1547
rect 230 1542 231 1546
rect 235 1542 236 1546
rect 230 1541 236 1542
rect 334 1546 340 1547
rect 334 1542 335 1546
rect 339 1542 340 1546
rect 334 1541 340 1542
rect 454 1546 460 1547
rect 454 1542 455 1546
rect 459 1542 460 1546
rect 454 1541 460 1542
rect 582 1546 588 1547
rect 582 1542 583 1546
rect 587 1542 588 1546
rect 582 1541 588 1542
rect 718 1546 724 1547
rect 718 1542 719 1546
rect 723 1542 724 1546
rect 718 1541 724 1542
rect 862 1546 868 1547
rect 862 1542 863 1546
rect 867 1542 868 1546
rect 862 1541 868 1542
rect 1006 1546 1012 1547
rect 1006 1542 1007 1546
rect 1011 1542 1012 1546
rect 1006 1541 1012 1542
rect 1150 1546 1156 1547
rect 1150 1542 1151 1546
rect 1155 1542 1156 1546
rect 1150 1541 1156 1542
rect 1286 1546 1292 1547
rect 1286 1542 1287 1546
rect 1291 1542 1292 1546
rect 1286 1541 1292 1542
rect 110 1537 116 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 110 1532 116 1533
rect 1326 1537 1332 1538
rect 1326 1533 1327 1537
rect 1331 1533 1332 1537
rect 1326 1532 1332 1533
rect 1414 1530 1420 1531
rect 1414 1526 1415 1530
rect 1419 1526 1420 1530
rect 1414 1525 1420 1526
rect 1526 1530 1532 1531
rect 1526 1526 1527 1530
rect 1531 1526 1532 1530
rect 1526 1525 1532 1526
rect 1646 1530 1652 1531
rect 1646 1526 1647 1530
rect 1651 1526 1652 1530
rect 1646 1525 1652 1526
rect 1766 1530 1772 1531
rect 1766 1526 1767 1530
rect 1771 1526 1772 1530
rect 1766 1525 1772 1526
rect 1878 1530 1884 1531
rect 1878 1526 1879 1530
rect 1883 1526 1884 1530
rect 1878 1525 1884 1526
rect 1982 1530 1988 1531
rect 1982 1526 1983 1530
rect 1987 1526 1988 1530
rect 1982 1525 1988 1526
rect 2078 1530 2084 1531
rect 2078 1526 2079 1530
rect 2083 1526 2084 1530
rect 2078 1525 2084 1526
rect 2166 1530 2172 1531
rect 2166 1526 2167 1530
rect 2171 1526 2172 1530
rect 2166 1525 2172 1526
rect 2254 1530 2260 1531
rect 2254 1526 2255 1530
rect 2259 1526 2260 1530
rect 2254 1525 2260 1526
rect 2334 1530 2340 1531
rect 2334 1526 2335 1530
rect 2339 1526 2340 1530
rect 2334 1525 2340 1526
rect 2406 1530 2412 1531
rect 2406 1526 2407 1530
rect 2411 1526 2412 1530
rect 2406 1525 2412 1526
rect 2486 1530 2492 1531
rect 2486 1526 2487 1530
rect 2491 1526 2492 1530
rect 2486 1525 2492 1526
rect 2542 1530 2548 1531
rect 2542 1526 2543 1530
rect 2547 1526 2548 1530
rect 2542 1525 2548 1526
rect 1366 1521 1372 1522
rect 110 1520 116 1521
rect 1326 1520 1332 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 110 1515 116 1516
rect 142 1519 148 1520
rect 142 1515 143 1519
rect 147 1515 148 1519
rect 142 1514 148 1515
rect 214 1519 220 1520
rect 214 1515 215 1519
rect 219 1515 220 1519
rect 214 1514 220 1515
rect 318 1519 324 1520
rect 318 1515 319 1519
rect 323 1515 324 1519
rect 318 1514 324 1515
rect 438 1519 444 1520
rect 438 1515 439 1519
rect 443 1515 444 1519
rect 438 1514 444 1515
rect 566 1519 572 1520
rect 566 1515 567 1519
rect 571 1515 572 1519
rect 566 1514 572 1515
rect 702 1519 708 1520
rect 702 1515 703 1519
rect 707 1515 708 1519
rect 702 1514 708 1515
rect 846 1519 852 1520
rect 846 1515 847 1519
rect 851 1515 852 1519
rect 846 1514 852 1515
rect 990 1519 996 1520
rect 990 1515 991 1519
rect 995 1515 996 1519
rect 990 1514 996 1515
rect 1134 1519 1140 1520
rect 1134 1515 1135 1519
rect 1139 1515 1140 1519
rect 1134 1514 1140 1515
rect 1270 1519 1276 1520
rect 1270 1515 1271 1519
rect 1275 1515 1276 1519
rect 1326 1516 1327 1520
rect 1331 1516 1332 1520
rect 1366 1517 1367 1521
rect 1371 1517 1372 1521
rect 1366 1516 1372 1517
rect 2582 1521 2588 1522
rect 2582 1517 2583 1521
rect 2587 1517 2588 1521
rect 2582 1516 2588 1517
rect 1326 1515 1332 1516
rect 1270 1514 1276 1515
rect 1366 1504 1372 1505
rect 2582 1504 2588 1505
rect 1366 1500 1367 1504
rect 1371 1500 1372 1504
rect 1366 1499 1372 1500
rect 1398 1503 1404 1504
rect 1398 1499 1399 1503
rect 1403 1499 1404 1503
rect 1398 1498 1404 1499
rect 1510 1503 1516 1504
rect 1510 1499 1511 1503
rect 1515 1499 1516 1503
rect 1510 1498 1516 1499
rect 1630 1503 1636 1504
rect 1630 1499 1631 1503
rect 1635 1499 1636 1503
rect 1630 1498 1636 1499
rect 1750 1503 1756 1504
rect 1750 1499 1751 1503
rect 1755 1499 1756 1503
rect 1750 1498 1756 1499
rect 1862 1503 1868 1504
rect 1862 1499 1863 1503
rect 1867 1499 1868 1503
rect 1862 1498 1868 1499
rect 1966 1503 1972 1504
rect 1966 1499 1967 1503
rect 1971 1499 1972 1503
rect 1966 1498 1972 1499
rect 2062 1503 2068 1504
rect 2062 1499 2063 1503
rect 2067 1499 2068 1503
rect 2062 1498 2068 1499
rect 2150 1503 2156 1504
rect 2150 1499 2151 1503
rect 2155 1499 2156 1503
rect 2150 1498 2156 1499
rect 2238 1503 2244 1504
rect 2238 1499 2239 1503
rect 2243 1499 2244 1503
rect 2238 1498 2244 1499
rect 2318 1503 2324 1504
rect 2318 1499 2319 1503
rect 2323 1499 2324 1503
rect 2318 1498 2324 1499
rect 2390 1503 2396 1504
rect 2390 1499 2391 1503
rect 2395 1499 2396 1503
rect 2390 1498 2396 1499
rect 2470 1503 2476 1504
rect 2470 1499 2471 1503
rect 2475 1499 2476 1503
rect 2470 1498 2476 1499
rect 2526 1503 2532 1504
rect 2526 1499 2527 1503
rect 2531 1499 2532 1503
rect 2582 1500 2583 1504
rect 2587 1500 2588 1504
rect 2582 1499 2588 1500
rect 2526 1498 2532 1499
rect 142 1485 148 1486
rect 110 1484 116 1485
rect 110 1480 111 1484
rect 115 1480 116 1484
rect 142 1481 143 1485
rect 147 1481 148 1485
rect 142 1480 148 1481
rect 198 1485 204 1486
rect 198 1481 199 1485
rect 203 1481 204 1485
rect 198 1480 204 1481
rect 270 1485 276 1486
rect 270 1481 271 1485
rect 275 1481 276 1485
rect 270 1480 276 1481
rect 366 1485 372 1486
rect 366 1481 367 1485
rect 371 1481 372 1485
rect 366 1480 372 1481
rect 478 1485 484 1486
rect 478 1481 479 1485
rect 483 1481 484 1485
rect 478 1480 484 1481
rect 590 1485 596 1486
rect 590 1481 591 1485
rect 595 1481 596 1485
rect 590 1480 596 1481
rect 702 1485 708 1486
rect 702 1481 703 1485
rect 707 1481 708 1485
rect 702 1480 708 1481
rect 806 1485 812 1486
rect 806 1481 807 1485
rect 811 1481 812 1485
rect 806 1480 812 1481
rect 910 1485 916 1486
rect 910 1481 911 1485
rect 915 1481 916 1485
rect 910 1480 916 1481
rect 1006 1485 1012 1486
rect 1006 1481 1007 1485
rect 1011 1481 1012 1485
rect 1006 1480 1012 1481
rect 1102 1485 1108 1486
rect 1102 1481 1103 1485
rect 1107 1481 1108 1485
rect 1102 1480 1108 1481
rect 1198 1485 1204 1486
rect 1198 1481 1199 1485
rect 1203 1481 1204 1485
rect 1198 1480 1204 1481
rect 1270 1485 1276 1486
rect 1270 1481 1271 1485
rect 1275 1481 1276 1485
rect 1270 1480 1276 1481
rect 1326 1484 1332 1485
rect 1326 1480 1327 1484
rect 1331 1480 1332 1484
rect 110 1479 116 1480
rect 1326 1479 1332 1480
rect 110 1467 116 1468
rect 110 1463 111 1467
rect 115 1463 116 1467
rect 110 1462 116 1463
rect 1326 1467 1332 1468
rect 1326 1463 1327 1467
rect 1331 1463 1332 1467
rect 1326 1462 1332 1463
rect 1398 1461 1404 1462
rect 1366 1460 1372 1461
rect 158 1458 164 1459
rect 158 1454 159 1458
rect 163 1454 164 1458
rect 158 1453 164 1454
rect 214 1458 220 1459
rect 214 1454 215 1458
rect 219 1454 220 1458
rect 214 1453 220 1454
rect 286 1458 292 1459
rect 286 1454 287 1458
rect 291 1454 292 1458
rect 286 1453 292 1454
rect 382 1458 388 1459
rect 382 1454 383 1458
rect 387 1454 388 1458
rect 382 1453 388 1454
rect 494 1458 500 1459
rect 494 1454 495 1458
rect 499 1454 500 1458
rect 494 1453 500 1454
rect 606 1458 612 1459
rect 606 1454 607 1458
rect 611 1454 612 1458
rect 606 1453 612 1454
rect 718 1458 724 1459
rect 718 1454 719 1458
rect 723 1454 724 1458
rect 718 1453 724 1454
rect 822 1458 828 1459
rect 822 1454 823 1458
rect 827 1454 828 1458
rect 822 1453 828 1454
rect 926 1458 932 1459
rect 926 1454 927 1458
rect 931 1454 932 1458
rect 926 1453 932 1454
rect 1022 1458 1028 1459
rect 1022 1454 1023 1458
rect 1027 1454 1028 1458
rect 1022 1453 1028 1454
rect 1118 1458 1124 1459
rect 1118 1454 1119 1458
rect 1123 1454 1124 1458
rect 1118 1453 1124 1454
rect 1214 1458 1220 1459
rect 1214 1454 1215 1458
rect 1219 1454 1220 1458
rect 1214 1453 1220 1454
rect 1286 1458 1292 1459
rect 1286 1454 1287 1458
rect 1291 1454 1292 1458
rect 1366 1456 1367 1460
rect 1371 1456 1372 1460
rect 1398 1457 1399 1461
rect 1403 1457 1404 1461
rect 1398 1456 1404 1457
rect 1502 1461 1508 1462
rect 1502 1457 1503 1461
rect 1507 1457 1508 1461
rect 1502 1456 1508 1457
rect 1630 1461 1636 1462
rect 1630 1457 1631 1461
rect 1635 1457 1636 1461
rect 1630 1456 1636 1457
rect 1750 1461 1756 1462
rect 1750 1457 1751 1461
rect 1755 1457 1756 1461
rect 1750 1456 1756 1457
rect 1870 1461 1876 1462
rect 1870 1457 1871 1461
rect 1875 1457 1876 1461
rect 1870 1456 1876 1457
rect 1982 1461 1988 1462
rect 1982 1457 1983 1461
rect 1987 1457 1988 1461
rect 1982 1456 1988 1457
rect 2086 1461 2092 1462
rect 2086 1457 2087 1461
rect 2091 1457 2092 1461
rect 2086 1456 2092 1457
rect 2182 1461 2188 1462
rect 2182 1457 2183 1461
rect 2187 1457 2188 1461
rect 2182 1456 2188 1457
rect 2270 1461 2276 1462
rect 2270 1457 2271 1461
rect 2275 1457 2276 1461
rect 2270 1456 2276 1457
rect 2358 1461 2364 1462
rect 2358 1457 2359 1461
rect 2363 1457 2364 1461
rect 2358 1456 2364 1457
rect 2454 1461 2460 1462
rect 2454 1457 2455 1461
rect 2459 1457 2460 1461
rect 2454 1456 2460 1457
rect 2526 1461 2532 1462
rect 2526 1457 2527 1461
rect 2531 1457 2532 1461
rect 2526 1456 2532 1457
rect 2582 1460 2588 1461
rect 2582 1456 2583 1460
rect 2587 1456 2588 1460
rect 1366 1455 1372 1456
rect 2582 1455 2588 1456
rect 1286 1453 1292 1454
rect 1366 1443 1372 1444
rect 1366 1439 1367 1443
rect 1371 1439 1372 1443
rect 1366 1438 1372 1439
rect 2582 1443 2588 1444
rect 2582 1439 2583 1443
rect 2587 1439 2588 1443
rect 2582 1438 2588 1439
rect 1414 1434 1420 1435
rect 254 1430 260 1431
rect 254 1426 255 1430
rect 259 1426 260 1430
rect 254 1425 260 1426
rect 310 1430 316 1431
rect 310 1426 311 1430
rect 315 1426 316 1430
rect 310 1425 316 1426
rect 374 1430 380 1431
rect 374 1426 375 1430
rect 379 1426 380 1430
rect 374 1425 380 1426
rect 446 1430 452 1431
rect 446 1426 447 1430
rect 451 1426 452 1430
rect 446 1425 452 1426
rect 526 1430 532 1431
rect 526 1426 527 1430
rect 531 1426 532 1430
rect 526 1425 532 1426
rect 606 1430 612 1431
rect 606 1426 607 1430
rect 611 1426 612 1430
rect 606 1425 612 1426
rect 694 1430 700 1431
rect 694 1426 695 1430
rect 699 1426 700 1430
rect 694 1425 700 1426
rect 782 1430 788 1431
rect 782 1426 783 1430
rect 787 1426 788 1430
rect 782 1425 788 1426
rect 870 1430 876 1431
rect 870 1426 871 1430
rect 875 1426 876 1430
rect 870 1425 876 1426
rect 958 1430 964 1431
rect 958 1426 959 1430
rect 963 1426 964 1430
rect 958 1425 964 1426
rect 1054 1430 1060 1431
rect 1054 1426 1055 1430
rect 1059 1426 1060 1430
rect 1054 1425 1060 1426
rect 1150 1430 1156 1431
rect 1150 1426 1151 1430
rect 1155 1426 1156 1430
rect 1414 1430 1415 1434
rect 1419 1430 1420 1434
rect 1414 1429 1420 1430
rect 1518 1434 1524 1435
rect 1518 1430 1519 1434
rect 1523 1430 1524 1434
rect 1518 1429 1524 1430
rect 1646 1434 1652 1435
rect 1646 1430 1647 1434
rect 1651 1430 1652 1434
rect 1646 1429 1652 1430
rect 1766 1434 1772 1435
rect 1766 1430 1767 1434
rect 1771 1430 1772 1434
rect 1766 1429 1772 1430
rect 1886 1434 1892 1435
rect 1886 1430 1887 1434
rect 1891 1430 1892 1434
rect 1886 1429 1892 1430
rect 1998 1434 2004 1435
rect 1998 1430 1999 1434
rect 2003 1430 2004 1434
rect 1998 1429 2004 1430
rect 2102 1434 2108 1435
rect 2102 1430 2103 1434
rect 2107 1430 2108 1434
rect 2102 1429 2108 1430
rect 2198 1434 2204 1435
rect 2198 1430 2199 1434
rect 2203 1430 2204 1434
rect 2198 1429 2204 1430
rect 2286 1434 2292 1435
rect 2286 1430 2287 1434
rect 2291 1430 2292 1434
rect 2286 1429 2292 1430
rect 2374 1434 2380 1435
rect 2374 1430 2375 1434
rect 2379 1430 2380 1434
rect 2374 1429 2380 1430
rect 2470 1434 2476 1435
rect 2470 1430 2471 1434
rect 2475 1430 2476 1434
rect 2470 1429 2476 1430
rect 2542 1434 2548 1435
rect 2542 1430 2543 1434
rect 2547 1430 2548 1434
rect 2542 1429 2548 1430
rect 1150 1425 1156 1426
rect 110 1421 116 1422
rect 110 1417 111 1421
rect 115 1417 116 1421
rect 110 1416 116 1417
rect 1326 1421 1332 1422
rect 1326 1417 1327 1421
rect 1331 1417 1332 1421
rect 1326 1416 1332 1417
rect 1414 1406 1420 1407
rect 110 1404 116 1405
rect 1326 1404 1332 1405
rect 110 1400 111 1404
rect 115 1400 116 1404
rect 110 1399 116 1400
rect 238 1403 244 1404
rect 238 1399 239 1403
rect 243 1399 244 1403
rect 238 1398 244 1399
rect 294 1403 300 1404
rect 294 1399 295 1403
rect 299 1399 300 1403
rect 294 1398 300 1399
rect 358 1403 364 1404
rect 358 1399 359 1403
rect 363 1399 364 1403
rect 358 1398 364 1399
rect 430 1403 436 1404
rect 430 1399 431 1403
rect 435 1399 436 1403
rect 430 1398 436 1399
rect 510 1403 516 1404
rect 510 1399 511 1403
rect 515 1399 516 1403
rect 510 1398 516 1399
rect 590 1403 596 1404
rect 590 1399 591 1403
rect 595 1399 596 1403
rect 590 1398 596 1399
rect 678 1403 684 1404
rect 678 1399 679 1403
rect 683 1399 684 1403
rect 678 1398 684 1399
rect 766 1403 772 1404
rect 766 1399 767 1403
rect 771 1399 772 1403
rect 766 1398 772 1399
rect 854 1403 860 1404
rect 854 1399 855 1403
rect 859 1399 860 1403
rect 854 1398 860 1399
rect 942 1403 948 1404
rect 942 1399 943 1403
rect 947 1399 948 1403
rect 942 1398 948 1399
rect 1038 1403 1044 1404
rect 1038 1399 1039 1403
rect 1043 1399 1044 1403
rect 1038 1398 1044 1399
rect 1134 1403 1140 1404
rect 1134 1399 1135 1403
rect 1139 1399 1140 1403
rect 1326 1400 1327 1404
rect 1331 1400 1332 1404
rect 1414 1402 1415 1406
rect 1419 1402 1420 1406
rect 1414 1401 1420 1402
rect 1470 1406 1476 1407
rect 1470 1402 1471 1406
rect 1475 1402 1476 1406
rect 1470 1401 1476 1402
rect 1550 1406 1556 1407
rect 1550 1402 1551 1406
rect 1555 1402 1556 1406
rect 1550 1401 1556 1402
rect 1630 1406 1636 1407
rect 1630 1402 1631 1406
rect 1635 1402 1636 1406
rect 1630 1401 1636 1402
rect 1710 1406 1716 1407
rect 1710 1402 1711 1406
rect 1715 1402 1716 1406
rect 1710 1401 1716 1402
rect 1790 1406 1796 1407
rect 1790 1402 1791 1406
rect 1795 1402 1796 1406
rect 1790 1401 1796 1402
rect 1870 1406 1876 1407
rect 1870 1402 1871 1406
rect 1875 1402 1876 1406
rect 1870 1401 1876 1402
rect 1958 1406 1964 1407
rect 1958 1402 1959 1406
rect 1963 1402 1964 1406
rect 1958 1401 1964 1402
rect 2054 1406 2060 1407
rect 2054 1402 2055 1406
rect 2059 1402 2060 1406
rect 2054 1401 2060 1402
rect 2166 1406 2172 1407
rect 2166 1402 2167 1406
rect 2171 1402 2172 1406
rect 2166 1401 2172 1402
rect 2294 1406 2300 1407
rect 2294 1402 2295 1406
rect 2299 1402 2300 1406
rect 2294 1401 2300 1402
rect 2430 1406 2436 1407
rect 2430 1402 2431 1406
rect 2435 1402 2436 1406
rect 2430 1401 2436 1402
rect 2542 1406 2548 1407
rect 2542 1402 2543 1406
rect 2547 1402 2548 1406
rect 2542 1401 2548 1402
rect 1326 1399 1332 1400
rect 1134 1398 1140 1399
rect 1366 1397 1372 1398
rect 1366 1393 1367 1397
rect 1371 1393 1372 1397
rect 1366 1392 1372 1393
rect 2582 1397 2588 1398
rect 2582 1393 2583 1397
rect 2587 1393 2588 1397
rect 2582 1392 2588 1393
rect 1366 1380 1372 1381
rect 2582 1380 2588 1381
rect 1366 1376 1367 1380
rect 1371 1376 1372 1380
rect 1366 1375 1372 1376
rect 1398 1379 1404 1380
rect 1398 1375 1399 1379
rect 1403 1375 1404 1379
rect 1398 1374 1404 1375
rect 1454 1379 1460 1380
rect 1454 1375 1455 1379
rect 1459 1375 1460 1379
rect 1454 1374 1460 1375
rect 1534 1379 1540 1380
rect 1534 1375 1535 1379
rect 1539 1375 1540 1379
rect 1534 1374 1540 1375
rect 1614 1379 1620 1380
rect 1614 1375 1615 1379
rect 1619 1375 1620 1379
rect 1614 1374 1620 1375
rect 1694 1379 1700 1380
rect 1694 1375 1695 1379
rect 1699 1375 1700 1379
rect 1694 1374 1700 1375
rect 1774 1379 1780 1380
rect 1774 1375 1775 1379
rect 1779 1375 1780 1379
rect 1774 1374 1780 1375
rect 1854 1379 1860 1380
rect 1854 1375 1855 1379
rect 1859 1375 1860 1379
rect 1854 1374 1860 1375
rect 1942 1379 1948 1380
rect 1942 1375 1943 1379
rect 1947 1375 1948 1379
rect 1942 1374 1948 1375
rect 2038 1379 2044 1380
rect 2038 1375 2039 1379
rect 2043 1375 2044 1379
rect 2038 1374 2044 1375
rect 2150 1379 2156 1380
rect 2150 1375 2151 1379
rect 2155 1375 2156 1379
rect 2150 1374 2156 1375
rect 2278 1379 2284 1380
rect 2278 1375 2279 1379
rect 2283 1375 2284 1379
rect 2278 1374 2284 1375
rect 2414 1379 2420 1380
rect 2414 1375 2415 1379
rect 2419 1375 2420 1379
rect 2414 1374 2420 1375
rect 2526 1379 2532 1380
rect 2526 1375 2527 1379
rect 2531 1375 2532 1379
rect 2582 1376 2583 1380
rect 2587 1376 2588 1380
rect 2582 1375 2588 1376
rect 2526 1374 2532 1375
rect 358 1361 364 1362
rect 110 1360 116 1361
rect 110 1356 111 1360
rect 115 1356 116 1360
rect 358 1357 359 1361
rect 363 1357 364 1361
rect 358 1356 364 1357
rect 414 1361 420 1362
rect 414 1357 415 1361
rect 419 1357 420 1361
rect 414 1356 420 1357
rect 470 1361 476 1362
rect 470 1357 471 1361
rect 475 1357 476 1361
rect 470 1356 476 1357
rect 526 1361 532 1362
rect 526 1357 527 1361
rect 531 1357 532 1361
rect 526 1356 532 1357
rect 590 1361 596 1362
rect 590 1357 591 1361
rect 595 1357 596 1361
rect 590 1356 596 1357
rect 670 1361 676 1362
rect 670 1357 671 1361
rect 675 1357 676 1361
rect 670 1356 676 1357
rect 750 1361 756 1362
rect 750 1357 751 1361
rect 755 1357 756 1361
rect 750 1356 756 1357
rect 838 1361 844 1362
rect 838 1357 839 1361
rect 843 1357 844 1361
rect 838 1356 844 1357
rect 934 1361 940 1362
rect 934 1357 935 1361
rect 939 1357 940 1361
rect 934 1356 940 1357
rect 1030 1361 1036 1362
rect 1030 1357 1031 1361
rect 1035 1357 1036 1361
rect 1030 1356 1036 1357
rect 1126 1361 1132 1362
rect 1126 1357 1127 1361
rect 1131 1357 1132 1361
rect 1126 1356 1132 1357
rect 1230 1361 1236 1362
rect 1230 1357 1231 1361
rect 1235 1357 1236 1361
rect 1230 1356 1236 1357
rect 1326 1360 1332 1361
rect 1326 1356 1327 1360
rect 1331 1356 1332 1360
rect 110 1355 116 1356
rect 1326 1355 1332 1356
rect 1422 1345 1428 1346
rect 1366 1344 1372 1345
rect 110 1343 116 1344
rect 110 1339 111 1343
rect 115 1339 116 1343
rect 110 1338 116 1339
rect 1326 1343 1332 1344
rect 1326 1339 1327 1343
rect 1331 1339 1332 1343
rect 1366 1340 1367 1344
rect 1371 1340 1372 1344
rect 1422 1341 1423 1345
rect 1427 1341 1428 1345
rect 1422 1340 1428 1341
rect 1494 1345 1500 1346
rect 1494 1341 1495 1345
rect 1499 1341 1500 1345
rect 1494 1340 1500 1341
rect 1574 1345 1580 1346
rect 1574 1341 1575 1345
rect 1579 1341 1580 1345
rect 1574 1340 1580 1341
rect 1654 1345 1660 1346
rect 1654 1341 1655 1345
rect 1659 1341 1660 1345
rect 1654 1340 1660 1341
rect 1758 1345 1764 1346
rect 1758 1341 1759 1345
rect 1763 1341 1764 1345
rect 1758 1340 1764 1341
rect 1878 1345 1884 1346
rect 1878 1341 1879 1345
rect 1883 1341 1884 1345
rect 1878 1340 1884 1341
rect 2022 1345 2028 1346
rect 2022 1341 2023 1345
rect 2027 1341 2028 1345
rect 2022 1340 2028 1341
rect 2182 1345 2188 1346
rect 2182 1341 2183 1345
rect 2187 1341 2188 1345
rect 2182 1340 2188 1341
rect 2358 1345 2364 1346
rect 2358 1341 2359 1345
rect 2363 1341 2364 1345
rect 2358 1340 2364 1341
rect 2526 1345 2532 1346
rect 2526 1341 2527 1345
rect 2531 1341 2532 1345
rect 2526 1340 2532 1341
rect 2582 1344 2588 1345
rect 2582 1340 2583 1344
rect 2587 1340 2588 1344
rect 1366 1339 1372 1340
rect 2582 1339 2588 1340
rect 1326 1338 1332 1339
rect 374 1334 380 1335
rect 374 1330 375 1334
rect 379 1330 380 1334
rect 374 1329 380 1330
rect 430 1334 436 1335
rect 430 1330 431 1334
rect 435 1330 436 1334
rect 430 1329 436 1330
rect 486 1334 492 1335
rect 486 1330 487 1334
rect 491 1330 492 1334
rect 486 1329 492 1330
rect 542 1334 548 1335
rect 542 1330 543 1334
rect 547 1330 548 1334
rect 542 1329 548 1330
rect 606 1334 612 1335
rect 606 1330 607 1334
rect 611 1330 612 1334
rect 606 1329 612 1330
rect 686 1334 692 1335
rect 686 1330 687 1334
rect 691 1330 692 1334
rect 686 1329 692 1330
rect 766 1334 772 1335
rect 766 1330 767 1334
rect 771 1330 772 1334
rect 766 1329 772 1330
rect 854 1334 860 1335
rect 854 1330 855 1334
rect 859 1330 860 1334
rect 854 1329 860 1330
rect 950 1334 956 1335
rect 950 1330 951 1334
rect 955 1330 956 1334
rect 950 1329 956 1330
rect 1046 1334 1052 1335
rect 1046 1330 1047 1334
rect 1051 1330 1052 1334
rect 1046 1329 1052 1330
rect 1142 1334 1148 1335
rect 1142 1330 1143 1334
rect 1147 1330 1148 1334
rect 1142 1329 1148 1330
rect 1246 1334 1252 1335
rect 1246 1330 1247 1334
rect 1251 1330 1252 1334
rect 1246 1329 1252 1330
rect 1366 1327 1372 1328
rect 1366 1323 1367 1327
rect 1371 1323 1372 1327
rect 1366 1322 1372 1323
rect 2582 1327 2588 1328
rect 2582 1323 2583 1327
rect 2587 1323 2588 1327
rect 2582 1322 2588 1323
rect 1438 1318 1444 1319
rect 1438 1314 1439 1318
rect 1443 1314 1444 1318
rect 1438 1313 1444 1314
rect 1510 1318 1516 1319
rect 1510 1314 1511 1318
rect 1515 1314 1516 1318
rect 1510 1313 1516 1314
rect 1590 1318 1596 1319
rect 1590 1314 1591 1318
rect 1595 1314 1596 1318
rect 1590 1313 1596 1314
rect 1670 1318 1676 1319
rect 1670 1314 1671 1318
rect 1675 1314 1676 1318
rect 1670 1313 1676 1314
rect 1774 1318 1780 1319
rect 1774 1314 1775 1318
rect 1779 1314 1780 1318
rect 1774 1313 1780 1314
rect 1894 1318 1900 1319
rect 1894 1314 1895 1318
rect 1899 1314 1900 1318
rect 1894 1313 1900 1314
rect 2038 1318 2044 1319
rect 2038 1314 2039 1318
rect 2043 1314 2044 1318
rect 2038 1313 2044 1314
rect 2198 1318 2204 1319
rect 2198 1314 2199 1318
rect 2203 1314 2204 1318
rect 2198 1313 2204 1314
rect 2374 1318 2380 1319
rect 2374 1314 2375 1318
rect 2379 1314 2380 1318
rect 2374 1313 2380 1314
rect 2542 1318 2548 1319
rect 2542 1314 2543 1318
rect 2547 1314 2548 1318
rect 2542 1313 2548 1314
rect 470 1302 476 1303
rect 470 1298 471 1302
rect 475 1298 476 1302
rect 470 1297 476 1298
rect 526 1302 532 1303
rect 526 1298 527 1302
rect 531 1298 532 1302
rect 526 1297 532 1298
rect 582 1302 588 1303
rect 582 1298 583 1302
rect 587 1298 588 1302
rect 582 1297 588 1298
rect 646 1302 652 1303
rect 646 1298 647 1302
rect 651 1298 652 1302
rect 646 1297 652 1298
rect 726 1302 732 1303
rect 726 1298 727 1302
rect 731 1298 732 1302
rect 726 1297 732 1298
rect 806 1302 812 1303
rect 806 1298 807 1302
rect 811 1298 812 1302
rect 806 1297 812 1298
rect 894 1302 900 1303
rect 894 1298 895 1302
rect 899 1298 900 1302
rect 894 1297 900 1298
rect 990 1302 996 1303
rect 990 1298 991 1302
rect 995 1298 996 1302
rect 990 1297 996 1298
rect 1094 1302 1100 1303
rect 1094 1298 1095 1302
rect 1099 1298 1100 1302
rect 1094 1297 1100 1298
rect 1198 1302 1204 1303
rect 1198 1298 1199 1302
rect 1203 1298 1204 1302
rect 1198 1297 1204 1298
rect 1286 1302 1292 1303
rect 1286 1298 1287 1302
rect 1291 1298 1292 1302
rect 1286 1297 1292 1298
rect 1430 1294 1436 1295
rect 110 1293 116 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 1326 1293 1332 1294
rect 1326 1289 1327 1293
rect 1331 1289 1332 1293
rect 1430 1290 1431 1294
rect 1435 1290 1436 1294
rect 1430 1289 1436 1290
rect 1494 1294 1500 1295
rect 1494 1290 1495 1294
rect 1499 1290 1500 1294
rect 1494 1289 1500 1290
rect 1558 1294 1564 1295
rect 1558 1290 1559 1294
rect 1563 1290 1564 1294
rect 1558 1289 1564 1290
rect 1630 1294 1636 1295
rect 1630 1290 1631 1294
rect 1635 1290 1636 1294
rect 1630 1289 1636 1290
rect 1702 1294 1708 1295
rect 1702 1290 1703 1294
rect 1707 1290 1708 1294
rect 1702 1289 1708 1290
rect 1774 1294 1780 1295
rect 1774 1290 1775 1294
rect 1779 1290 1780 1294
rect 1774 1289 1780 1290
rect 1854 1294 1860 1295
rect 1854 1290 1855 1294
rect 1859 1290 1860 1294
rect 1854 1289 1860 1290
rect 1942 1294 1948 1295
rect 1942 1290 1943 1294
rect 1947 1290 1948 1294
rect 1942 1289 1948 1290
rect 2046 1294 2052 1295
rect 2046 1290 2047 1294
rect 2051 1290 2052 1294
rect 2046 1289 2052 1290
rect 2158 1294 2164 1295
rect 2158 1290 2159 1294
rect 2163 1290 2164 1294
rect 2158 1289 2164 1290
rect 2286 1294 2292 1295
rect 2286 1290 2287 1294
rect 2291 1290 2292 1294
rect 2286 1289 2292 1290
rect 2422 1294 2428 1295
rect 2422 1290 2423 1294
rect 2427 1290 2428 1294
rect 2422 1289 2428 1290
rect 2542 1294 2548 1295
rect 2542 1290 2543 1294
rect 2547 1290 2548 1294
rect 2542 1289 2548 1290
rect 1326 1288 1332 1289
rect 1366 1285 1372 1286
rect 1366 1281 1367 1285
rect 1371 1281 1372 1285
rect 1366 1280 1372 1281
rect 2582 1285 2588 1286
rect 2582 1281 2583 1285
rect 2587 1281 2588 1285
rect 2582 1280 2588 1281
rect 110 1276 116 1277
rect 1326 1276 1332 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 110 1271 116 1272
rect 454 1275 460 1276
rect 454 1271 455 1275
rect 459 1271 460 1275
rect 454 1270 460 1271
rect 510 1275 516 1276
rect 510 1271 511 1275
rect 515 1271 516 1275
rect 510 1270 516 1271
rect 566 1275 572 1276
rect 566 1271 567 1275
rect 571 1271 572 1275
rect 566 1270 572 1271
rect 630 1275 636 1276
rect 630 1271 631 1275
rect 635 1271 636 1275
rect 630 1270 636 1271
rect 710 1275 716 1276
rect 710 1271 711 1275
rect 715 1271 716 1275
rect 710 1270 716 1271
rect 790 1275 796 1276
rect 790 1271 791 1275
rect 795 1271 796 1275
rect 790 1270 796 1271
rect 878 1275 884 1276
rect 878 1271 879 1275
rect 883 1271 884 1275
rect 878 1270 884 1271
rect 974 1275 980 1276
rect 974 1271 975 1275
rect 979 1271 980 1275
rect 974 1270 980 1271
rect 1078 1275 1084 1276
rect 1078 1271 1079 1275
rect 1083 1271 1084 1275
rect 1078 1270 1084 1271
rect 1182 1275 1188 1276
rect 1182 1271 1183 1275
rect 1187 1271 1188 1275
rect 1182 1270 1188 1271
rect 1270 1275 1276 1276
rect 1270 1271 1271 1275
rect 1275 1271 1276 1275
rect 1326 1272 1327 1276
rect 1331 1272 1332 1276
rect 1326 1271 1332 1272
rect 1270 1270 1276 1271
rect 1366 1268 1372 1269
rect 2582 1268 2588 1269
rect 1366 1264 1367 1268
rect 1371 1264 1372 1268
rect 1366 1263 1372 1264
rect 1414 1267 1420 1268
rect 1414 1263 1415 1267
rect 1419 1263 1420 1267
rect 1414 1262 1420 1263
rect 1478 1267 1484 1268
rect 1478 1263 1479 1267
rect 1483 1263 1484 1267
rect 1478 1262 1484 1263
rect 1542 1267 1548 1268
rect 1542 1263 1543 1267
rect 1547 1263 1548 1267
rect 1542 1262 1548 1263
rect 1614 1267 1620 1268
rect 1614 1263 1615 1267
rect 1619 1263 1620 1267
rect 1614 1262 1620 1263
rect 1686 1267 1692 1268
rect 1686 1263 1687 1267
rect 1691 1263 1692 1267
rect 1686 1262 1692 1263
rect 1758 1267 1764 1268
rect 1758 1263 1759 1267
rect 1763 1263 1764 1267
rect 1758 1262 1764 1263
rect 1838 1267 1844 1268
rect 1838 1263 1839 1267
rect 1843 1263 1844 1267
rect 1838 1262 1844 1263
rect 1926 1267 1932 1268
rect 1926 1263 1927 1267
rect 1931 1263 1932 1267
rect 1926 1262 1932 1263
rect 2030 1267 2036 1268
rect 2030 1263 2031 1267
rect 2035 1263 2036 1267
rect 2030 1262 2036 1263
rect 2142 1267 2148 1268
rect 2142 1263 2143 1267
rect 2147 1263 2148 1267
rect 2142 1262 2148 1263
rect 2270 1267 2276 1268
rect 2270 1263 2271 1267
rect 2275 1263 2276 1267
rect 2270 1262 2276 1263
rect 2406 1267 2412 1268
rect 2406 1263 2407 1267
rect 2411 1263 2412 1267
rect 2406 1262 2412 1263
rect 2526 1267 2532 1268
rect 2526 1263 2527 1267
rect 2531 1263 2532 1267
rect 2582 1264 2583 1268
rect 2587 1264 2588 1268
rect 2582 1263 2588 1264
rect 2526 1262 2532 1263
rect 382 1237 388 1238
rect 110 1236 116 1237
rect 110 1232 111 1236
rect 115 1232 116 1236
rect 382 1233 383 1237
rect 387 1233 388 1237
rect 382 1232 388 1233
rect 438 1237 444 1238
rect 438 1233 439 1237
rect 443 1233 444 1237
rect 438 1232 444 1233
rect 502 1237 508 1238
rect 502 1233 503 1237
rect 507 1233 508 1237
rect 502 1232 508 1233
rect 574 1237 580 1238
rect 574 1233 575 1237
rect 579 1233 580 1237
rect 574 1232 580 1233
rect 646 1237 652 1238
rect 646 1233 647 1237
rect 651 1233 652 1237
rect 646 1232 652 1233
rect 726 1237 732 1238
rect 726 1233 727 1237
rect 731 1233 732 1237
rect 726 1232 732 1233
rect 814 1237 820 1238
rect 814 1233 815 1237
rect 819 1233 820 1237
rect 814 1232 820 1233
rect 902 1237 908 1238
rect 902 1233 903 1237
rect 907 1233 908 1237
rect 902 1232 908 1233
rect 990 1237 996 1238
rect 990 1233 991 1237
rect 995 1233 996 1237
rect 990 1232 996 1233
rect 1078 1237 1084 1238
rect 1078 1233 1079 1237
rect 1083 1233 1084 1237
rect 1078 1232 1084 1233
rect 1174 1237 1180 1238
rect 1174 1233 1175 1237
rect 1179 1233 1180 1237
rect 1174 1232 1180 1233
rect 1270 1237 1276 1238
rect 1270 1233 1271 1237
rect 1275 1233 1276 1237
rect 1270 1232 1276 1233
rect 1326 1236 1332 1237
rect 1326 1232 1327 1236
rect 1331 1232 1332 1236
rect 110 1231 116 1232
rect 1326 1231 1332 1232
rect 1398 1229 1404 1230
rect 1366 1228 1372 1229
rect 1366 1224 1367 1228
rect 1371 1224 1372 1228
rect 1398 1225 1399 1229
rect 1403 1225 1404 1229
rect 1398 1224 1404 1225
rect 1454 1229 1460 1230
rect 1454 1225 1455 1229
rect 1459 1225 1460 1229
rect 1454 1224 1460 1225
rect 1534 1229 1540 1230
rect 1534 1225 1535 1229
rect 1539 1225 1540 1229
rect 1534 1224 1540 1225
rect 1614 1229 1620 1230
rect 1614 1225 1615 1229
rect 1619 1225 1620 1229
rect 1614 1224 1620 1225
rect 1694 1229 1700 1230
rect 1694 1225 1695 1229
rect 1699 1225 1700 1229
rect 1694 1224 1700 1225
rect 1774 1229 1780 1230
rect 1774 1225 1775 1229
rect 1779 1225 1780 1229
rect 1774 1224 1780 1225
rect 1854 1229 1860 1230
rect 1854 1225 1855 1229
rect 1859 1225 1860 1229
rect 1854 1224 1860 1225
rect 1942 1229 1948 1230
rect 1942 1225 1943 1229
rect 1947 1225 1948 1229
rect 1942 1224 1948 1225
rect 2038 1229 2044 1230
rect 2038 1225 2039 1229
rect 2043 1225 2044 1229
rect 2038 1224 2044 1225
rect 2150 1229 2156 1230
rect 2150 1225 2151 1229
rect 2155 1225 2156 1229
rect 2150 1224 2156 1225
rect 2278 1229 2284 1230
rect 2278 1225 2279 1229
rect 2283 1225 2284 1229
rect 2278 1224 2284 1225
rect 2414 1229 2420 1230
rect 2414 1225 2415 1229
rect 2419 1225 2420 1229
rect 2414 1224 2420 1225
rect 2526 1229 2532 1230
rect 2526 1225 2527 1229
rect 2531 1225 2532 1229
rect 2526 1224 2532 1225
rect 2582 1228 2588 1229
rect 2582 1224 2583 1228
rect 2587 1224 2588 1228
rect 1366 1223 1372 1224
rect 2582 1223 2588 1224
rect 110 1219 116 1220
rect 110 1215 111 1219
rect 115 1215 116 1219
rect 110 1214 116 1215
rect 1326 1219 1332 1220
rect 1326 1215 1327 1219
rect 1331 1215 1332 1219
rect 1326 1214 1332 1215
rect 1366 1211 1372 1212
rect 398 1210 404 1211
rect 398 1206 399 1210
rect 403 1206 404 1210
rect 398 1205 404 1206
rect 454 1210 460 1211
rect 454 1206 455 1210
rect 459 1206 460 1210
rect 454 1205 460 1206
rect 518 1210 524 1211
rect 518 1206 519 1210
rect 523 1206 524 1210
rect 518 1205 524 1206
rect 590 1210 596 1211
rect 590 1206 591 1210
rect 595 1206 596 1210
rect 590 1205 596 1206
rect 662 1210 668 1211
rect 662 1206 663 1210
rect 667 1206 668 1210
rect 662 1205 668 1206
rect 742 1210 748 1211
rect 742 1206 743 1210
rect 747 1206 748 1210
rect 742 1205 748 1206
rect 830 1210 836 1211
rect 830 1206 831 1210
rect 835 1206 836 1210
rect 830 1205 836 1206
rect 918 1210 924 1211
rect 918 1206 919 1210
rect 923 1206 924 1210
rect 918 1205 924 1206
rect 1006 1210 1012 1211
rect 1006 1206 1007 1210
rect 1011 1206 1012 1210
rect 1006 1205 1012 1206
rect 1094 1210 1100 1211
rect 1094 1206 1095 1210
rect 1099 1206 1100 1210
rect 1094 1205 1100 1206
rect 1190 1210 1196 1211
rect 1190 1206 1191 1210
rect 1195 1206 1196 1210
rect 1190 1205 1196 1206
rect 1286 1210 1292 1211
rect 1286 1206 1287 1210
rect 1291 1206 1292 1210
rect 1366 1207 1367 1211
rect 1371 1207 1372 1211
rect 1366 1206 1372 1207
rect 2582 1211 2588 1212
rect 2582 1207 2583 1211
rect 2587 1207 2588 1211
rect 2582 1206 2588 1207
rect 1286 1205 1292 1206
rect 1414 1202 1420 1203
rect 1414 1198 1415 1202
rect 1419 1198 1420 1202
rect 1414 1197 1420 1198
rect 1470 1202 1476 1203
rect 1470 1198 1471 1202
rect 1475 1198 1476 1202
rect 1470 1197 1476 1198
rect 1550 1202 1556 1203
rect 1550 1198 1551 1202
rect 1555 1198 1556 1202
rect 1550 1197 1556 1198
rect 1630 1202 1636 1203
rect 1630 1198 1631 1202
rect 1635 1198 1636 1202
rect 1630 1197 1636 1198
rect 1710 1202 1716 1203
rect 1710 1198 1711 1202
rect 1715 1198 1716 1202
rect 1710 1197 1716 1198
rect 1790 1202 1796 1203
rect 1790 1198 1791 1202
rect 1795 1198 1796 1202
rect 1790 1197 1796 1198
rect 1870 1202 1876 1203
rect 1870 1198 1871 1202
rect 1875 1198 1876 1202
rect 1870 1197 1876 1198
rect 1958 1202 1964 1203
rect 1958 1198 1959 1202
rect 1963 1198 1964 1202
rect 1958 1197 1964 1198
rect 2054 1202 2060 1203
rect 2054 1198 2055 1202
rect 2059 1198 2060 1202
rect 2054 1197 2060 1198
rect 2166 1202 2172 1203
rect 2166 1198 2167 1202
rect 2171 1198 2172 1202
rect 2166 1197 2172 1198
rect 2294 1202 2300 1203
rect 2294 1198 2295 1202
rect 2299 1198 2300 1202
rect 2294 1197 2300 1198
rect 2430 1202 2436 1203
rect 2430 1198 2431 1202
rect 2435 1198 2436 1202
rect 2430 1197 2436 1198
rect 2542 1202 2548 1203
rect 2542 1198 2543 1202
rect 2547 1198 2548 1202
rect 2542 1197 2548 1198
rect 278 1182 284 1183
rect 278 1178 279 1182
rect 283 1178 284 1182
rect 278 1177 284 1178
rect 342 1182 348 1183
rect 342 1178 343 1182
rect 347 1178 348 1182
rect 342 1177 348 1178
rect 414 1182 420 1183
rect 414 1178 415 1182
rect 419 1178 420 1182
rect 414 1177 420 1178
rect 494 1182 500 1183
rect 494 1178 495 1182
rect 499 1178 500 1182
rect 494 1177 500 1178
rect 582 1182 588 1183
rect 582 1178 583 1182
rect 587 1178 588 1182
rect 582 1177 588 1178
rect 670 1182 676 1183
rect 670 1178 671 1182
rect 675 1178 676 1182
rect 670 1177 676 1178
rect 758 1182 764 1183
rect 758 1178 759 1182
rect 763 1178 764 1182
rect 758 1177 764 1178
rect 846 1182 852 1183
rect 846 1178 847 1182
rect 851 1178 852 1182
rect 846 1177 852 1178
rect 934 1182 940 1183
rect 934 1178 935 1182
rect 939 1178 940 1182
rect 934 1177 940 1178
rect 1014 1182 1020 1183
rect 1014 1178 1015 1182
rect 1019 1178 1020 1182
rect 1014 1177 1020 1178
rect 1086 1182 1092 1183
rect 1086 1178 1087 1182
rect 1091 1178 1092 1182
rect 1086 1177 1092 1178
rect 1158 1182 1164 1183
rect 1158 1178 1159 1182
rect 1163 1178 1164 1182
rect 1158 1177 1164 1178
rect 1230 1182 1236 1183
rect 1230 1178 1231 1182
rect 1235 1178 1236 1182
rect 1230 1177 1236 1178
rect 1286 1182 1292 1183
rect 1286 1178 1287 1182
rect 1291 1178 1292 1182
rect 1286 1177 1292 1178
rect 110 1173 116 1174
rect 110 1169 111 1173
rect 115 1169 116 1173
rect 110 1168 116 1169
rect 1326 1173 1332 1174
rect 1326 1169 1327 1173
rect 1331 1169 1332 1173
rect 1326 1168 1332 1169
rect 1694 1170 1700 1171
rect 1694 1166 1695 1170
rect 1699 1166 1700 1170
rect 1694 1165 1700 1166
rect 1766 1170 1772 1171
rect 1766 1166 1767 1170
rect 1771 1166 1772 1170
rect 1766 1165 1772 1166
rect 1846 1170 1852 1171
rect 1846 1166 1847 1170
rect 1851 1166 1852 1170
rect 1846 1165 1852 1166
rect 1918 1170 1924 1171
rect 1918 1166 1919 1170
rect 1923 1166 1924 1170
rect 1918 1165 1924 1166
rect 1990 1170 1996 1171
rect 1990 1166 1991 1170
rect 1995 1166 1996 1170
rect 1990 1165 1996 1166
rect 2062 1170 2068 1171
rect 2062 1166 2063 1170
rect 2067 1166 2068 1170
rect 2062 1165 2068 1166
rect 2134 1170 2140 1171
rect 2134 1166 2135 1170
rect 2139 1166 2140 1170
rect 2134 1165 2140 1166
rect 2206 1170 2212 1171
rect 2206 1166 2207 1170
rect 2211 1166 2212 1170
rect 2206 1165 2212 1166
rect 2286 1170 2292 1171
rect 2286 1166 2287 1170
rect 2291 1166 2292 1170
rect 2286 1165 2292 1166
rect 2366 1170 2372 1171
rect 2366 1166 2367 1170
rect 2371 1166 2372 1170
rect 2366 1165 2372 1166
rect 1366 1161 1372 1162
rect 1366 1157 1367 1161
rect 1371 1157 1372 1161
rect 110 1156 116 1157
rect 1326 1156 1332 1157
rect 1366 1156 1372 1157
rect 2582 1161 2588 1162
rect 2582 1157 2583 1161
rect 2587 1157 2588 1161
rect 2582 1156 2588 1157
rect 110 1152 111 1156
rect 115 1152 116 1156
rect 110 1151 116 1152
rect 262 1155 268 1156
rect 262 1151 263 1155
rect 267 1151 268 1155
rect 262 1150 268 1151
rect 326 1155 332 1156
rect 326 1151 327 1155
rect 331 1151 332 1155
rect 326 1150 332 1151
rect 398 1155 404 1156
rect 398 1151 399 1155
rect 403 1151 404 1155
rect 398 1150 404 1151
rect 478 1155 484 1156
rect 478 1151 479 1155
rect 483 1151 484 1155
rect 478 1150 484 1151
rect 566 1155 572 1156
rect 566 1151 567 1155
rect 571 1151 572 1155
rect 566 1150 572 1151
rect 654 1155 660 1156
rect 654 1151 655 1155
rect 659 1151 660 1155
rect 654 1150 660 1151
rect 742 1155 748 1156
rect 742 1151 743 1155
rect 747 1151 748 1155
rect 742 1150 748 1151
rect 830 1155 836 1156
rect 830 1151 831 1155
rect 835 1151 836 1155
rect 830 1150 836 1151
rect 918 1155 924 1156
rect 918 1151 919 1155
rect 923 1151 924 1155
rect 918 1150 924 1151
rect 998 1155 1004 1156
rect 998 1151 999 1155
rect 1003 1151 1004 1155
rect 998 1150 1004 1151
rect 1070 1155 1076 1156
rect 1070 1151 1071 1155
rect 1075 1151 1076 1155
rect 1070 1150 1076 1151
rect 1142 1155 1148 1156
rect 1142 1151 1143 1155
rect 1147 1151 1148 1155
rect 1142 1150 1148 1151
rect 1214 1155 1220 1156
rect 1214 1151 1215 1155
rect 1219 1151 1220 1155
rect 1214 1150 1220 1151
rect 1270 1155 1276 1156
rect 1270 1151 1271 1155
rect 1275 1151 1276 1155
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1326 1151 1332 1152
rect 1270 1150 1276 1151
rect 1366 1144 1372 1145
rect 2582 1144 2588 1145
rect 1366 1140 1367 1144
rect 1371 1140 1372 1144
rect 1366 1139 1372 1140
rect 1678 1143 1684 1144
rect 1678 1139 1679 1143
rect 1683 1139 1684 1143
rect 1678 1138 1684 1139
rect 1750 1143 1756 1144
rect 1750 1139 1751 1143
rect 1755 1139 1756 1143
rect 1750 1138 1756 1139
rect 1830 1143 1836 1144
rect 1830 1139 1831 1143
rect 1835 1139 1836 1143
rect 1830 1138 1836 1139
rect 1902 1143 1908 1144
rect 1902 1139 1903 1143
rect 1907 1139 1908 1143
rect 1902 1138 1908 1139
rect 1974 1143 1980 1144
rect 1974 1139 1975 1143
rect 1979 1139 1980 1143
rect 1974 1138 1980 1139
rect 2046 1143 2052 1144
rect 2046 1139 2047 1143
rect 2051 1139 2052 1143
rect 2046 1138 2052 1139
rect 2118 1143 2124 1144
rect 2118 1139 2119 1143
rect 2123 1139 2124 1143
rect 2118 1138 2124 1139
rect 2190 1143 2196 1144
rect 2190 1139 2191 1143
rect 2195 1139 2196 1143
rect 2190 1138 2196 1139
rect 2270 1143 2276 1144
rect 2270 1139 2271 1143
rect 2275 1139 2276 1143
rect 2270 1138 2276 1139
rect 2350 1143 2356 1144
rect 2350 1139 2351 1143
rect 2355 1139 2356 1143
rect 2582 1140 2583 1144
rect 2587 1140 2588 1144
rect 2582 1139 2588 1140
rect 2350 1138 2356 1139
rect 142 1113 148 1114
rect 110 1112 116 1113
rect 110 1108 111 1112
rect 115 1108 116 1112
rect 142 1109 143 1113
rect 147 1109 148 1113
rect 142 1108 148 1109
rect 206 1113 212 1114
rect 206 1109 207 1113
rect 211 1109 212 1113
rect 206 1108 212 1109
rect 270 1113 276 1114
rect 270 1109 271 1113
rect 275 1109 276 1113
rect 270 1108 276 1109
rect 342 1113 348 1114
rect 342 1109 343 1113
rect 347 1109 348 1113
rect 342 1108 348 1109
rect 422 1113 428 1114
rect 422 1109 423 1113
rect 427 1109 428 1113
rect 422 1108 428 1109
rect 502 1113 508 1114
rect 502 1109 503 1113
rect 507 1109 508 1113
rect 502 1108 508 1109
rect 582 1113 588 1114
rect 582 1109 583 1113
rect 587 1109 588 1113
rect 582 1108 588 1109
rect 662 1113 668 1114
rect 662 1109 663 1113
rect 667 1109 668 1113
rect 662 1108 668 1109
rect 742 1113 748 1114
rect 742 1109 743 1113
rect 747 1109 748 1113
rect 742 1108 748 1109
rect 830 1113 836 1114
rect 830 1109 831 1113
rect 835 1109 836 1113
rect 830 1108 836 1109
rect 918 1113 924 1114
rect 918 1109 919 1113
rect 923 1109 924 1113
rect 918 1108 924 1109
rect 1006 1113 1012 1114
rect 1006 1109 1007 1113
rect 1011 1109 1012 1113
rect 1006 1108 1012 1109
rect 1326 1112 1332 1113
rect 1326 1108 1327 1112
rect 1331 1108 1332 1112
rect 1398 1109 1404 1110
rect 110 1107 116 1108
rect 1326 1107 1332 1108
rect 1366 1108 1372 1109
rect 1366 1104 1367 1108
rect 1371 1104 1372 1108
rect 1398 1105 1399 1109
rect 1403 1105 1404 1109
rect 1398 1104 1404 1105
rect 1478 1109 1484 1110
rect 1478 1105 1479 1109
rect 1483 1105 1484 1109
rect 1478 1104 1484 1105
rect 1582 1109 1588 1110
rect 1582 1105 1583 1109
rect 1587 1105 1588 1109
rect 1582 1104 1588 1105
rect 1686 1109 1692 1110
rect 1686 1105 1687 1109
rect 1691 1105 1692 1109
rect 1686 1104 1692 1105
rect 1782 1109 1788 1110
rect 1782 1105 1783 1109
rect 1787 1105 1788 1109
rect 1782 1104 1788 1105
rect 1878 1109 1884 1110
rect 1878 1105 1879 1109
rect 1883 1105 1884 1109
rect 1878 1104 1884 1105
rect 1974 1109 1980 1110
rect 1974 1105 1975 1109
rect 1979 1105 1980 1109
rect 1974 1104 1980 1105
rect 2062 1109 2068 1110
rect 2062 1105 2063 1109
rect 2067 1105 2068 1109
rect 2062 1104 2068 1105
rect 2150 1109 2156 1110
rect 2150 1105 2151 1109
rect 2155 1105 2156 1109
rect 2150 1104 2156 1105
rect 2238 1109 2244 1110
rect 2238 1105 2239 1109
rect 2243 1105 2244 1109
rect 2238 1104 2244 1105
rect 2326 1109 2332 1110
rect 2326 1105 2327 1109
rect 2331 1105 2332 1109
rect 2326 1104 2332 1105
rect 2414 1109 2420 1110
rect 2414 1105 2415 1109
rect 2419 1105 2420 1109
rect 2414 1104 2420 1105
rect 2582 1108 2588 1109
rect 2582 1104 2583 1108
rect 2587 1104 2588 1108
rect 1366 1103 1372 1104
rect 2582 1103 2588 1104
rect 110 1095 116 1096
rect 110 1091 111 1095
rect 115 1091 116 1095
rect 110 1090 116 1091
rect 1326 1095 1332 1096
rect 1326 1091 1327 1095
rect 1331 1091 1332 1095
rect 1326 1090 1332 1091
rect 1366 1091 1372 1092
rect 1366 1087 1367 1091
rect 1371 1087 1372 1091
rect 158 1086 164 1087
rect 158 1082 159 1086
rect 163 1082 164 1086
rect 158 1081 164 1082
rect 222 1086 228 1087
rect 222 1082 223 1086
rect 227 1082 228 1086
rect 222 1081 228 1082
rect 286 1086 292 1087
rect 286 1082 287 1086
rect 291 1082 292 1086
rect 286 1081 292 1082
rect 358 1086 364 1087
rect 358 1082 359 1086
rect 363 1082 364 1086
rect 358 1081 364 1082
rect 438 1086 444 1087
rect 438 1082 439 1086
rect 443 1082 444 1086
rect 438 1081 444 1082
rect 518 1086 524 1087
rect 518 1082 519 1086
rect 523 1082 524 1086
rect 518 1081 524 1082
rect 598 1086 604 1087
rect 598 1082 599 1086
rect 603 1082 604 1086
rect 598 1081 604 1082
rect 678 1086 684 1087
rect 678 1082 679 1086
rect 683 1082 684 1086
rect 678 1081 684 1082
rect 758 1086 764 1087
rect 758 1082 759 1086
rect 763 1082 764 1086
rect 758 1081 764 1082
rect 846 1086 852 1087
rect 846 1082 847 1086
rect 851 1082 852 1086
rect 846 1081 852 1082
rect 934 1086 940 1087
rect 934 1082 935 1086
rect 939 1082 940 1086
rect 934 1081 940 1082
rect 1022 1086 1028 1087
rect 1366 1086 1372 1087
rect 2582 1091 2588 1092
rect 2582 1087 2583 1091
rect 2587 1087 2588 1091
rect 2582 1086 2588 1087
rect 1022 1082 1023 1086
rect 1027 1082 1028 1086
rect 1022 1081 1028 1082
rect 1414 1082 1420 1083
rect 1414 1078 1415 1082
rect 1419 1078 1420 1082
rect 1414 1077 1420 1078
rect 1494 1082 1500 1083
rect 1494 1078 1495 1082
rect 1499 1078 1500 1082
rect 1494 1077 1500 1078
rect 1598 1082 1604 1083
rect 1598 1078 1599 1082
rect 1603 1078 1604 1082
rect 1598 1077 1604 1078
rect 1702 1082 1708 1083
rect 1702 1078 1703 1082
rect 1707 1078 1708 1082
rect 1702 1077 1708 1078
rect 1798 1082 1804 1083
rect 1798 1078 1799 1082
rect 1803 1078 1804 1082
rect 1798 1077 1804 1078
rect 1894 1082 1900 1083
rect 1894 1078 1895 1082
rect 1899 1078 1900 1082
rect 1894 1077 1900 1078
rect 1990 1082 1996 1083
rect 1990 1078 1991 1082
rect 1995 1078 1996 1082
rect 1990 1077 1996 1078
rect 2078 1082 2084 1083
rect 2078 1078 2079 1082
rect 2083 1078 2084 1082
rect 2078 1077 2084 1078
rect 2166 1082 2172 1083
rect 2166 1078 2167 1082
rect 2171 1078 2172 1082
rect 2166 1077 2172 1078
rect 2254 1082 2260 1083
rect 2254 1078 2255 1082
rect 2259 1078 2260 1082
rect 2254 1077 2260 1078
rect 2342 1082 2348 1083
rect 2342 1078 2343 1082
rect 2347 1078 2348 1082
rect 2342 1077 2348 1078
rect 2430 1082 2436 1083
rect 2430 1078 2431 1082
rect 2435 1078 2436 1082
rect 2430 1077 2436 1078
rect 158 1058 164 1059
rect 158 1054 159 1058
rect 163 1054 164 1058
rect 158 1053 164 1054
rect 214 1058 220 1059
rect 214 1054 215 1058
rect 219 1054 220 1058
rect 214 1053 220 1054
rect 286 1058 292 1059
rect 286 1054 287 1058
rect 291 1054 292 1058
rect 286 1053 292 1054
rect 382 1058 388 1059
rect 382 1054 383 1058
rect 387 1054 388 1058
rect 382 1053 388 1054
rect 478 1058 484 1059
rect 478 1054 479 1058
rect 483 1054 484 1058
rect 478 1053 484 1054
rect 582 1058 588 1059
rect 582 1054 583 1058
rect 587 1054 588 1058
rect 582 1053 588 1054
rect 686 1058 692 1059
rect 686 1054 687 1058
rect 691 1054 692 1058
rect 686 1053 692 1054
rect 782 1058 788 1059
rect 782 1054 783 1058
rect 787 1054 788 1058
rect 782 1053 788 1054
rect 878 1058 884 1059
rect 878 1054 879 1058
rect 883 1054 884 1058
rect 878 1053 884 1054
rect 966 1058 972 1059
rect 966 1054 967 1058
rect 971 1054 972 1058
rect 966 1053 972 1054
rect 1062 1058 1068 1059
rect 1062 1054 1063 1058
rect 1067 1054 1068 1058
rect 1062 1053 1068 1054
rect 1158 1058 1164 1059
rect 1158 1054 1159 1058
rect 1163 1054 1164 1058
rect 1158 1053 1164 1054
rect 1414 1058 1420 1059
rect 1414 1054 1415 1058
rect 1419 1054 1420 1058
rect 1414 1053 1420 1054
rect 1510 1058 1516 1059
rect 1510 1054 1511 1058
rect 1515 1054 1516 1058
rect 1510 1053 1516 1054
rect 1630 1058 1636 1059
rect 1630 1054 1631 1058
rect 1635 1054 1636 1058
rect 1630 1053 1636 1054
rect 1750 1058 1756 1059
rect 1750 1054 1751 1058
rect 1755 1054 1756 1058
rect 1750 1053 1756 1054
rect 1870 1058 1876 1059
rect 1870 1054 1871 1058
rect 1875 1054 1876 1058
rect 1870 1053 1876 1054
rect 1990 1058 1996 1059
rect 1990 1054 1991 1058
rect 1995 1054 1996 1058
rect 1990 1053 1996 1054
rect 2102 1058 2108 1059
rect 2102 1054 2103 1058
rect 2107 1054 2108 1058
rect 2102 1053 2108 1054
rect 2198 1058 2204 1059
rect 2198 1054 2199 1058
rect 2203 1054 2204 1058
rect 2198 1053 2204 1054
rect 2294 1058 2300 1059
rect 2294 1054 2295 1058
rect 2299 1054 2300 1058
rect 2294 1053 2300 1054
rect 2382 1058 2388 1059
rect 2382 1054 2383 1058
rect 2387 1054 2388 1058
rect 2382 1053 2388 1054
rect 2470 1058 2476 1059
rect 2470 1054 2471 1058
rect 2475 1054 2476 1058
rect 2470 1053 2476 1054
rect 2542 1058 2548 1059
rect 2542 1054 2543 1058
rect 2547 1054 2548 1058
rect 2542 1053 2548 1054
rect 110 1049 116 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 1326 1049 1332 1050
rect 1326 1045 1327 1049
rect 1331 1045 1332 1049
rect 1326 1044 1332 1045
rect 1366 1049 1372 1050
rect 1366 1045 1367 1049
rect 1371 1045 1372 1049
rect 1366 1044 1372 1045
rect 2582 1049 2588 1050
rect 2582 1045 2583 1049
rect 2587 1045 2588 1049
rect 2582 1044 2588 1045
rect 110 1032 116 1033
rect 1326 1032 1332 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 110 1027 116 1028
rect 142 1031 148 1032
rect 142 1027 143 1031
rect 147 1027 148 1031
rect 142 1026 148 1027
rect 198 1031 204 1032
rect 198 1027 199 1031
rect 203 1027 204 1031
rect 198 1026 204 1027
rect 270 1031 276 1032
rect 270 1027 271 1031
rect 275 1027 276 1031
rect 270 1026 276 1027
rect 366 1031 372 1032
rect 366 1027 367 1031
rect 371 1027 372 1031
rect 366 1026 372 1027
rect 462 1031 468 1032
rect 462 1027 463 1031
rect 467 1027 468 1031
rect 462 1026 468 1027
rect 566 1031 572 1032
rect 566 1027 567 1031
rect 571 1027 572 1031
rect 566 1026 572 1027
rect 670 1031 676 1032
rect 670 1027 671 1031
rect 675 1027 676 1031
rect 670 1026 676 1027
rect 766 1031 772 1032
rect 766 1027 767 1031
rect 771 1027 772 1031
rect 766 1026 772 1027
rect 862 1031 868 1032
rect 862 1027 863 1031
rect 867 1027 868 1031
rect 862 1026 868 1027
rect 950 1031 956 1032
rect 950 1027 951 1031
rect 955 1027 956 1031
rect 950 1026 956 1027
rect 1046 1031 1052 1032
rect 1046 1027 1047 1031
rect 1051 1027 1052 1031
rect 1046 1026 1052 1027
rect 1142 1031 1148 1032
rect 1142 1027 1143 1031
rect 1147 1027 1148 1031
rect 1326 1028 1327 1032
rect 1331 1028 1332 1032
rect 1326 1027 1332 1028
rect 1366 1032 1372 1033
rect 2582 1032 2588 1033
rect 1366 1028 1367 1032
rect 1371 1028 1372 1032
rect 1366 1027 1372 1028
rect 1398 1031 1404 1032
rect 1398 1027 1399 1031
rect 1403 1027 1404 1031
rect 1142 1026 1148 1027
rect 1398 1026 1404 1027
rect 1494 1031 1500 1032
rect 1494 1027 1495 1031
rect 1499 1027 1500 1031
rect 1494 1026 1500 1027
rect 1614 1031 1620 1032
rect 1614 1027 1615 1031
rect 1619 1027 1620 1031
rect 1614 1026 1620 1027
rect 1734 1031 1740 1032
rect 1734 1027 1735 1031
rect 1739 1027 1740 1031
rect 1734 1026 1740 1027
rect 1854 1031 1860 1032
rect 1854 1027 1855 1031
rect 1859 1027 1860 1031
rect 1854 1026 1860 1027
rect 1974 1031 1980 1032
rect 1974 1027 1975 1031
rect 1979 1027 1980 1031
rect 1974 1026 1980 1027
rect 2086 1031 2092 1032
rect 2086 1027 2087 1031
rect 2091 1027 2092 1031
rect 2086 1026 2092 1027
rect 2182 1031 2188 1032
rect 2182 1027 2183 1031
rect 2187 1027 2188 1031
rect 2182 1026 2188 1027
rect 2278 1031 2284 1032
rect 2278 1027 2279 1031
rect 2283 1027 2284 1031
rect 2278 1026 2284 1027
rect 2366 1031 2372 1032
rect 2366 1027 2367 1031
rect 2371 1027 2372 1031
rect 2366 1026 2372 1027
rect 2454 1031 2460 1032
rect 2454 1027 2455 1031
rect 2459 1027 2460 1031
rect 2454 1026 2460 1027
rect 2526 1031 2532 1032
rect 2526 1027 2527 1031
rect 2531 1027 2532 1031
rect 2582 1028 2583 1032
rect 2587 1028 2588 1032
rect 2582 1027 2588 1028
rect 2526 1026 2532 1027
rect 142 993 148 994
rect 110 992 116 993
rect 110 988 111 992
rect 115 988 116 992
rect 142 989 143 993
rect 147 989 148 993
rect 142 988 148 989
rect 198 993 204 994
rect 198 989 199 993
rect 203 989 204 993
rect 198 988 204 989
rect 278 993 284 994
rect 278 989 279 993
rect 283 989 284 993
rect 278 988 284 989
rect 382 993 388 994
rect 382 989 383 993
rect 387 989 388 993
rect 382 988 388 989
rect 494 993 500 994
rect 494 989 495 993
rect 499 989 500 993
rect 494 988 500 989
rect 614 993 620 994
rect 614 989 615 993
rect 619 989 620 993
rect 614 988 620 989
rect 726 993 732 994
rect 726 989 727 993
rect 731 989 732 993
rect 726 988 732 989
rect 838 993 844 994
rect 838 989 839 993
rect 843 989 844 993
rect 838 988 844 989
rect 950 993 956 994
rect 950 989 951 993
rect 955 989 956 993
rect 950 988 956 989
rect 1054 993 1060 994
rect 1054 989 1055 993
rect 1059 989 1060 993
rect 1054 988 1060 989
rect 1158 993 1164 994
rect 1158 989 1159 993
rect 1163 989 1164 993
rect 1158 988 1164 989
rect 1270 993 1276 994
rect 1486 993 1492 994
rect 1270 989 1271 993
rect 1275 989 1276 993
rect 1270 988 1276 989
rect 1326 992 1332 993
rect 1326 988 1327 992
rect 1331 988 1332 992
rect 110 987 116 988
rect 1326 987 1332 988
rect 1366 992 1372 993
rect 1366 988 1367 992
rect 1371 988 1372 992
rect 1486 989 1487 993
rect 1491 989 1492 993
rect 1486 988 1492 989
rect 1582 993 1588 994
rect 1582 989 1583 993
rect 1587 989 1588 993
rect 1582 988 1588 989
rect 1694 993 1700 994
rect 1694 989 1695 993
rect 1699 989 1700 993
rect 1694 988 1700 989
rect 1806 993 1812 994
rect 1806 989 1807 993
rect 1811 989 1812 993
rect 1806 988 1812 989
rect 1918 993 1924 994
rect 1918 989 1919 993
rect 1923 989 1924 993
rect 1918 988 1924 989
rect 2022 993 2028 994
rect 2022 989 2023 993
rect 2027 989 2028 993
rect 2022 988 2028 989
rect 2118 993 2124 994
rect 2118 989 2119 993
rect 2123 989 2124 993
rect 2118 988 2124 989
rect 2214 993 2220 994
rect 2214 989 2215 993
rect 2219 989 2220 993
rect 2214 988 2220 989
rect 2302 993 2308 994
rect 2302 989 2303 993
rect 2307 989 2308 993
rect 2302 988 2308 989
rect 2382 993 2388 994
rect 2382 989 2383 993
rect 2387 989 2388 993
rect 2382 988 2388 989
rect 2462 993 2468 994
rect 2462 989 2463 993
rect 2467 989 2468 993
rect 2462 988 2468 989
rect 2526 993 2532 994
rect 2526 989 2527 993
rect 2531 989 2532 993
rect 2526 988 2532 989
rect 2582 992 2588 993
rect 2582 988 2583 992
rect 2587 988 2588 992
rect 1366 987 1372 988
rect 2582 987 2588 988
rect 110 975 116 976
rect 110 971 111 975
rect 115 971 116 975
rect 110 970 116 971
rect 1326 975 1332 976
rect 1326 971 1327 975
rect 1331 971 1332 975
rect 1326 970 1332 971
rect 1366 975 1372 976
rect 1366 971 1367 975
rect 1371 971 1372 975
rect 1366 970 1372 971
rect 2582 975 2588 976
rect 2582 971 2583 975
rect 2587 971 2588 975
rect 2582 970 2588 971
rect 158 966 164 967
rect 158 962 159 966
rect 163 962 164 966
rect 158 961 164 962
rect 214 966 220 967
rect 214 962 215 966
rect 219 962 220 966
rect 214 961 220 962
rect 294 966 300 967
rect 294 962 295 966
rect 299 962 300 966
rect 294 961 300 962
rect 398 966 404 967
rect 398 962 399 966
rect 403 962 404 966
rect 398 961 404 962
rect 510 966 516 967
rect 510 962 511 966
rect 515 962 516 966
rect 510 961 516 962
rect 630 966 636 967
rect 630 962 631 966
rect 635 962 636 966
rect 630 961 636 962
rect 742 966 748 967
rect 742 962 743 966
rect 747 962 748 966
rect 742 961 748 962
rect 854 966 860 967
rect 854 962 855 966
rect 859 962 860 966
rect 854 961 860 962
rect 966 966 972 967
rect 966 962 967 966
rect 971 962 972 966
rect 966 961 972 962
rect 1070 966 1076 967
rect 1070 962 1071 966
rect 1075 962 1076 966
rect 1070 961 1076 962
rect 1174 966 1180 967
rect 1174 962 1175 966
rect 1179 962 1180 966
rect 1174 961 1180 962
rect 1286 966 1292 967
rect 1286 962 1287 966
rect 1291 962 1292 966
rect 1286 961 1292 962
rect 1502 966 1508 967
rect 1502 962 1503 966
rect 1507 962 1508 966
rect 1502 961 1508 962
rect 1598 966 1604 967
rect 1598 962 1599 966
rect 1603 962 1604 966
rect 1598 961 1604 962
rect 1710 966 1716 967
rect 1710 962 1711 966
rect 1715 962 1716 966
rect 1710 961 1716 962
rect 1822 966 1828 967
rect 1822 962 1823 966
rect 1827 962 1828 966
rect 1822 961 1828 962
rect 1934 966 1940 967
rect 1934 962 1935 966
rect 1939 962 1940 966
rect 1934 961 1940 962
rect 2038 966 2044 967
rect 2038 962 2039 966
rect 2043 962 2044 966
rect 2038 961 2044 962
rect 2134 966 2140 967
rect 2134 962 2135 966
rect 2139 962 2140 966
rect 2134 961 2140 962
rect 2230 966 2236 967
rect 2230 962 2231 966
rect 2235 962 2236 966
rect 2230 961 2236 962
rect 2318 966 2324 967
rect 2318 962 2319 966
rect 2323 962 2324 966
rect 2318 961 2324 962
rect 2398 966 2404 967
rect 2398 962 2399 966
rect 2403 962 2404 966
rect 2398 961 2404 962
rect 2478 966 2484 967
rect 2478 962 2479 966
rect 2483 962 2484 966
rect 2478 961 2484 962
rect 2542 966 2548 967
rect 2542 962 2543 966
rect 2547 962 2548 966
rect 2542 961 2548 962
rect 158 934 164 935
rect 158 930 159 934
rect 163 930 164 934
rect 158 929 164 930
rect 214 934 220 935
rect 214 930 215 934
rect 219 930 220 934
rect 214 929 220 930
rect 286 934 292 935
rect 286 930 287 934
rect 291 930 292 934
rect 286 929 292 930
rect 374 934 380 935
rect 374 930 375 934
rect 379 930 380 934
rect 374 929 380 930
rect 470 934 476 935
rect 470 930 471 934
rect 475 930 476 934
rect 470 929 476 930
rect 566 934 572 935
rect 566 930 567 934
rect 571 930 572 934
rect 566 929 572 930
rect 670 934 676 935
rect 670 930 671 934
rect 675 930 676 934
rect 670 929 676 930
rect 766 934 772 935
rect 766 930 767 934
rect 771 930 772 934
rect 766 929 772 930
rect 862 934 868 935
rect 862 930 863 934
rect 867 930 868 934
rect 862 929 868 930
rect 958 934 964 935
rect 958 930 959 934
rect 963 930 964 934
rect 958 929 964 930
rect 1046 934 1052 935
rect 1046 930 1047 934
rect 1051 930 1052 934
rect 1046 929 1052 930
rect 1134 934 1140 935
rect 1134 930 1135 934
rect 1139 930 1140 934
rect 1134 929 1140 930
rect 1222 934 1228 935
rect 1222 930 1223 934
rect 1227 930 1228 934
rect 1222 929 1228 930
rect 1286 934 1292 935
rect 1286 930 1287 934
rect 1291 930 1292 934
rect 1286 929 1292 930
rect 1414 934 1420 935
rect 1414 930 1415 934
rect 1419 930 1420 934
rect 1414 929 1420 930
rect 1534 934 1540 935
rect 1534 930 1535 934
rect 1539 930 1540 934
rect 1534 929 1540 930
rect 1670 934 1676 935
rect 1670 930 1671 934
rect 1675 930 1676 934
rect 1670 929 1676 930
rect 1806 934 1812 935
rect 1806 930 1807 934
rect 1811 930 1812 934
rect 1806 929 1812 930
rect 1934 934 1940 935
rect 1934 930 1935 934
rect 1939 930 1940 934
rect 1934 929 1940 930
rect 2054 934 2060 935
rect 2054 930 2055 934
rect 2059 930 2060 934
rect 2054 929 2060 930
rect 2166 934 2172 935
rect 2166 930 2167 934
rect 2171 930 2172 934
rect 2166 929 2172 930
rect 2270 934 2276 935
rect 2270 930 2271 934
rect 2275 930 2276 934
rect 2270 929 2276 930
rect 2366 934 2372 935
rect 2366 930 2367 934
rect 2371 930 2372 934
rect 2366 929 2372 930
rect 2462 934 2468 935
rect 2462 930 2463 934
rect 2467 930 2468 934
rect 2462 929 2468 930
rect 2542 934 2548 935
rect 2542 930 2543 934
rect 2547 930 2548 934
rect 2542 929 2548 930
rect 110 925 116 926
rect 110 921 111 925
rect 115 921 116 925
rect 110 920 116 921
rect 1326 925 1332 926
rect 1326 921 1327 925
rect 1331 921 1332 925
rect 1326 920 1332 921
rect 1366 925 1372 926
rect 1366 921 1367 925
rect 1371 921 1372 925
rect 1366 920 1372 921
rect 2582 925 2588 926
rect 2582 921 2583 925
rect 2587 921 2588 925
rect 2582 920 2588 921
rect 110 908 116 909
rect 1326 908 1332 909
rect 110 904 111 908
rect 115 904 116 908
rect 110 903 116 904
rect 142 907 148 908
rect 142 903 143 907
rect 147 903 148 907
rect 142 902 148 903
rect 198 907 204 908
rect 198 903 199 907
rect 203 903 204 907
rect 198 902 204 903
rect 270 907 276 908
rect 270 903 271 907
rect 275 903 276 907
rect 270 902 276 903
rect 358 907 364 908
rect 358 903 359 907
rect 363 903 364 907
rect 358 902 364 903
rect 454 907 460 908
rect 454 903 455 907
rect 459 903 460 907
rect 454 902 460 903
rect 550 907 556 908
rect 550 903 551 907
rect 555 903 556 907
rect 550 902 556 903
rect 654 907 660 908
rect 654 903 655 907
rect 659 903 660 907
rect 654 902 660 903
rect 750 907 756 908
rect 750 903 751 907
rect 755 903 756 907
rect 750 902 756 903
rect 846 907 852 908
rect 846 903 847 907
rect 851 903 852 907
rect 846 902 852 903
rect 942 907 948 908
rect 942 903 943 907
rect 947 903 948 907
rect 942 902 948 903
rect 1030 907 1036 908
rect 1030 903 1031 907
rect 1035 903 1036 907
rect 1030 902 1036 903
rect 1118 907 1124 908
rect 1118 903 1119 907
rect 1123 903 1124 907
rect 1118 902 1124 903
rect 1206 907 1212 908
rect 1206 903 1207 907
rect 1211 903 1212 907
rect 1206 902 1212 903
rect 1270 907 1276 908
rect 1270 903 1271 907
rect 1275 903 1276 907
rect 1326 904 1327 908
rect 1331 904 1332 908
rect 1326 903 1332 904
rect 1366 908 1372 909
rect 2582 908 2588 909
rect 1366 904 1367 908
rect 1371 904 1372 908
rect 1366 903 1372 904
rect 1398 907 1404 908
rect 1398 903 1399 907
rect 1403 903 1404 907
rect 1270 902 1276 903
rect 1398 902 1404 903
rect 1518 907 1524 908
rect 1518 903 1519 907
rect 1523 903 1524 907
rect 1518 902 1524 903
rect 1654 907 1660 908
rect 1654 903 1655 907
rect 1659 903 1660 907
rect 1654 902 1660 903
rect 1790 907 1796 908
rect 1790 903 1791 907
rect 1795 903 1796 907
rect 1790 902 1796 903
rect 1918 907 1924 908
rect 1918 903 1919 907
rect 1923 903 1924 907
rect 1918 902 1924 903
rect 2038 907 2044 908
rect 2038 903 2039 907
rect 2043 903 2044 907
rect 2038 902 2044 903
rect 2150 907 2156 908
rect 2150 903 2151 907
rect 2155 903 2156 907
rect 2150 902 2156 903
rect 2254 907 2260 908
rect 2254 903 2255 907
rect 2259 903 2260 907
rect 2254 902 2260 903
rect 2350 907 2356 908
rect 2350 903 2351 907
rect 2355 903 2356 907
rect 2350 902 2356 903
rect 2446 907 2452 908
rect 2446 903 2447 907
rect 2451 903 2452 907
rect 2446 902 2452 903
rect 2526 907 2532 908
rect 2526 903 2527 907
rect 2531 903 2532 907
rect 2582 904 2583 908
rect 2587 904 2588 908
rect 2582 903 2588 904
rect 2526 902 2532 903
rect 182 869 188 870
rect 110 868 116 869
rect 110 864 111 868
rect 115 864 116 868
rect 182 865 183 869
rect 187 865 188 869
rect 182 864 188 865
rect 238 869 244 870
rect 238 865 239 869
rect 243 865 244 869
rect 238 864 244 865
rect 302 869 308 870
rect 302 865 303 869
rect 307 865 308 869
rect 302 864 308 865
rect 374 869 380 870
rect 374 865 375 869
rect 379 865 380 869
rect 374 864 380 865
rect 454 869 460 870
rect 454 865 455 869
rect 459 865 460 869
rect 454 864 460 865
rect 542 869 548 870
rect 542 865 543 869
rect 547 865 548 869
rect 542 864 548 865
rect 638 869 644 870
rect 638 865 639 869
rect 643 865 644 869
rect 638 864 644 865
rect 742 869 748 870
rect 742 865 743 869
rect 747 865 748 869
rect 742 864 748 865
rect 854 869 860 870
rect 854 865 855 869
rect 859 865 860 869
rect 854 864 860 865
rect 966 869 972 870
rect 966 865 967 869
rect 971 865 972 869
rect 966 864 972 865
rect 1086 869 1092 870
rect 1086 865 1087 869
rect 1091 865 1092 869
rect 1086 864 1092 865
rect 1214 869 1220 870
rect 1398 869 1404 870
rect 1214 865 1215 869
rect 1219 865 1220 869
rect 1214 864 1220 865
rect 1326 868 1332 869
rect 1326 864 1327 868
rect 1331 864 1332 868
rect 110 863 116 864
rect 1326 863 1332 864
rect 1366 868 1372 869
rect 1366 864 1367 868
rect 1371 864 1372 868
rect 1398 865 1399 869
rect 1403 865 1404 869
rect 1398 864 1404 865
rect 1454 869 1460 870
rect 1454 865 1455 869
rect 1459 865 1460 869
rect 1454 864 1460 865
rect 1518 869 1524 870
rect 1518 865 1519 869
rect 1523 865 1524 869
rect 1518 864 1524 865
rect 1606 869 1612 870
rect 1606 865 1607 869
rect 1611 865 1612 869
rect 1606 864 1612 865
rect 1694 869 1700 870
rect 1694 865 1695 869
rect 1699 865 1700 869
rect 1694 864 1700 865
rect 1790 869 1796 870
rect 1790 865 1791 869
rect 1795 865 1796 869
rect 1790 864 1796 865
rect 1894 869 1900 870
rect 1894 865 1895 869
rect 1899 865 1900 869
rect 1894 864 1900 865
rect 1998 869 2004 870
rect 1998 865 1999 869
rect 2003 865 2004 869
rect 1998 864 2004 865
rect 2102 869 2108 870
rect 2102 865 2103 869
rect 2107 865 2108 869
rect 2102 864 2108 865
rect 2206 869 2212 870
rect 2206 865 2207 869
rect 2211 865 2212 869
rect 2206 864 2212 865
rect 2310 869 2316 870
rect 2310 865 2311 869
rect 2315 865 2316 869
rect 2310 864 2316 865
rect 2422 869 2428 870
rect 2422 865 2423 869
rect 2427 865 2428 869
rect 2422 864 2428 865
rect 2526 869 2532 870
rect 2526 865 2527 869
rect 2531 865 2532 869
rect 2526 864 2532 865
rect 2582 868 2588 869
rect 2582 864 2583 868
rect 2587 864 2588 868
rect 1366 863 1372 864
rect 2582 863 2588 864
rect 110 851 116 852
rect 110 847 111 851
rect 115 847 116 851
rect 110 846 116 847
rect 1326 851 1332 852
rect 1326 847 1327 851
rect 1331 847 1332 851
rect 1326 846 1332 847
rect 1366 851 1372 852
rect 1366 847 1367 851
rect 1371 847 1372 851
rect 1366 846 1372 847
rect 2582 851 2588 852
rect 2582 847 2583 851
rect 2587 847 2588 851
rect 2582 846 2588 847
rect 198 842 204 843
rect 198 838 199 842
rect 203 838 204 842
rect 198 837 204 838
rect 254 842 260 843
rect 254 838 255 842
rect 259 838 260 842
rect 254 837 260 838
rect 318 842 324 843
rect 318 838 319 842
rect 323 838 324 842
rect 318 837 324 838
rect 390 842 396 843
rect 390 838 391 842
rect 395 838 396 842
rect 390 837 396 838
rect 470 842 476 843
rect 470 838 471 842
rect 475 838 476 842
rect 470 837 476 838
rect 558 842 564 843
rect 558 838 559 842
rect 563 838 564 842
rect 558 837 564 838
rect 654 842 660 843
rect 654 838 655 842
rect 659 838 660 842
rect 654 837 660 838
rect 758 842 764 843
rect 758 838 759 842
rect 763 838 764 842
rect 758 837 764 838
rect 870 842 876 843
rect 870 838 871 842
rect 875 838 876 842
rect 870 837 876 838
rect 982 842 988 843
rect 982 838 983 842
rect 987 838 988 842
rect 982 837 988 838
rect 1102 842 1108 843
rect 1102 838 1103 842
rect 1107 838 1108 842
rect 1102 837 1108 838
rect 1230 842 1236 843
rect 1230 838 1231 842
rect 1235 838 1236 842
rect 1230 837 1236 838
rect 1414 842 1420 843
rect 1414 838 1415 842
rect 1419 838 1420 842
rect 1414 837 1420 838
rect 1470 842 1476 843
rect 1470 838 1471 842
rect 1475 838 1476 842
rect 1470 837 1476 838
rect 1534 842 1540 843
rect 1534 838 1535 842
rect 1539 838 1540 842
rect 1534 837 1540 838
rect 1622 842 1628 843
rect 1622 838 1623 842
rect 1627 838 1628 842
rect 1622 837 1628 838
rect 1710 842 1716 843
rect 1710 838 1711 842
rect 1715 838 1716 842
rect 1710 837 1716 838
rect 1806 842 1812 843
rect 1806 838 1807 842
rect 1811 838 1812 842
rect 1806 837 1812 838
rect 1910 842 1916 843
rect 1910 838 1911 842
rect 1915 838 1916 842
rect 1910 837 1916 838
rect 2014 842 2020 843
rect 2014 838 2015 842
rect 2019 838 2020 842
rect 2014 837 2020 838
rect 2118 842 2124 843
rect 2118 838 2119 842
rect 2123 838 2124 842
rect 2118 837 2124 838
rect 2222 842 2228 843
rect 2222 838 2223 842
rect 2227 838 2228 842
rect 2222 837 2228 838
rect 2326 842 2332 843
rect 2326 838 2327 842
rect 2331 838 2332 842
rect 2326 837 2332 838
rect 2438 842 2444 843
rect 2438 838 2439 842
rect 2443 838 2444 842
rect 2438 837 2444 838
rect 2542 842 2548 843
rect 2542 838 2543 842
rect 2547 838 2548 842
rect 2542 837 2548 838
rect 1526 814 1532 815
rect 382 810 388 811
rect 382 806 383 810
rect 387 806 388 810
rect 382 805 388 806
rect 438 810 444 811
rect 438 806 439 810
rect 443 806 444 810
rect 438 805 444 806
rect 494 810 500 811
rect 494 806 495 810
rect 499 806 500 810
rect 494 805 500 806
rect 558 810 564 811
rect 558 806 559 810
rect 563 806 564 810
rect 558 805 564 806
rect 630 810 636 811
rect 630 806 631 810
rect 635 806 636 810
rect 630 805 636 806
rect 702 810 708 811
rect 702 806 703 810
rect 707 806 708 810
rect 702 805 708 806
rect 782 810 788 811
rect 782 806 783 810
rect 787 806 788 810
rect 782 805 788 806
rect 870 810 876 811
rect 870 806 871 810
rect 875 806 876 810
rect 870 805 876 806
rect 958 810 964 811
rect 958 806 959 810
rect 963 806 964 810
rect 958 805 964 806
rect 1046 810 1052 811
rect 1046 806 1047 810
rect 1051 806 1052 810
rect 1046 805 1052 806
rect 1134 810 1140 811
rect 1134 806 1135 810
rect 1139 806 1140 810
rect 1134 805 1140 806
rect 1222 810 1228 811
rect 1222 806 1223 810
rect 1227 806 1228 810
rect 1526 810 1527 814
rect 1531 810 1532 814
rect 1526 809 1532 810
rect 1582 814 1588 815
rect 1582 810 1583 814
rect 1587 810 1588 814
rect 1582 809 1588 810
rect 1638 814 1644 815
rect 1638 810 1639 814
rect 1643 810 1644 814
rect 1638 809 1644 810
rect 1694 814 1700 815
rect 1694 810 1695 814
rect 1699 810 1700 814
rect 1694 809 1700 810
rect 1750 814 1756 815
rect 1750 810 1751 814
rect 1755 810 1756 814
rect 1750 809 1756 810
rect 1806 814 1812 815
rect 1806 810 1807 814
rect 1811 810 1812 814
rect 1806 809 1812 810
rect 1878 814 1884 815
rect 1878 810 1879 814
rect 1883 810 1884 814
rect 1878 809 1884 810
rect 1958 814 1964 815
rect 1958 810 1959 814
rect 1963 810 1964 814
rect 1958 809 1964 810
rect 2054 814 2060 815
rect 2054 810 2055 814
rect 2059 810 2060 814
rect 2054 809 2060 810
rect 2166 814 2172 815
rect 2166 810 2167 814
rect 2171 810 2172 814
rect 2166 809 2172 810
rect 2294 814 2300 815
rect 2294 810 2295 814
rect 2299 810 2300 814
rect 2294 809 2300 810
rect 2430 814 2436 815
rect 2430 810 2431 814
rect 2435 810 2436 814
rect 2430 809 2436 810
rect 2542 814 2548 815
rect 2542 810 2543 814
rect 2547 810 2548 814
rect 2542 809 2548 810
rect 1222 805 1228 806
rect 1366 805 1372 806
rect 110 801 116 802
rect 110 797 111 801
rect 115 797 116 801
rect 110 796 116 797
rect 1326 801 1332 802
rect 1326 797 1327 801
rect 1331 797 1332 801
rect 1366 801 1367 805
rect 1371 801 1372 805
rect 1366 800 1372 801
rect 2582 805 2588 806
rect 2582 801 2583 805
rect 2587 801 2588 805
rect 2582 800 2588 801
rect 1326 796 1332 797
rect 1366 788 1372 789
rect 2582 788 2588 789
rect 110 784 116 785
rect 1326 784 1332 785
rect 110 780 111 784
rect 115 780 116 784
rect 110 779 116 780
rect 366 783 372 784
rect 366 779 367 783
rect 371 779 372 783
rect 366 778 372 779
rect 422 783 428 784
rect 422 779 423 783
rect 427 779 428 783
rect 422 778 428 779
rect 478 783 484 784
rect 478 779 479 783
rect 483 779 484 783
rect 478 778 484 779
rect 542 783 548 784
rect 542 779 543 783
rect 547 779 548 783
rect 542 778 548 779
rect 614 783 620 784
rect 614 779 615 783
rect 619 779 620 783
rect 614 778 620 779
rect 686 783 692 784
rect 686 779 687 783
rect 691 779 692 783
rect 686 778 692 779
rect 766 783 772 784
rect 766 779 767 783
rect 771 779 772 783
rect 766 778 772 779
rect 854 783 860 784
rect 854 779 855 783
rect 859 779 860 783
rect 854 778 860 779
rect 942 783 948 784
rect 942 779 943 783
rect 947 779 948 783
rect 942 778 948 779
rect 1030 783 1036 784
rect 1030 779 1031 783
rect 1035 779 1036 783
rect 1030 778 1036 779
rect 1118 783 1124 784
rect 1118 779 1119 783
rect 1123 779 1124 783
rect 1118 778 1124 779
rect 1206 783 1212 784
rect 1206 779 1207 783
rect 1211 779 1212 783
rect 1326 780 1327 784
rect 1331 780 1332 784
rect 1366 784 1367 788
rect 1371 784 1372 788
rect 1366 783 1372 784
rect 1510 787 1516 788
rect 1510 783 1511 787
rect 1515 783 1516 787
rect 1510 782 1516 783
rect 1566 787 1572 788
rect 1566 783 1567 787
rect 1571 783 1572 787
rect 1566 782 1572 783
rect 1622 787 1628 788
rect 1622 783 1623 787
rect 1627 783 1628 787
rect 1622 782 1628 783
rect 1678 787 1684 788
rect 1678 783 1679 787
rect 1683 783 1684 787
rect 1678 782 1684 783
rect 1734 787 1740 788
rect 1734 783 1735 787
rect 1739 783 1740 787
rect 1734 782 1740 783
rect 1790 787 1796 788
rect 1790 783 1791 787
rect 1795 783 1796 787
rect 1790 782 1796 783
rect 1862 787 1868 788
rect 1862 783 1863 787
rect 1867 783 1868 787
rect 1862 782 1868 783
rect 1942 787 1948 788
rect 1942 783 1943 787
rect 1947 783 1948 787
rect 1942 782 1948 783
rect 2038 787 2044 788
rect 2038 783 2039 787
rect 2043 783 2044 787
rect 2038 782 2044 783
rect 2150 787 2156 788
rect 2150 783 2151 787
rect 2155 783 2156 787
rect 2150 782 2156 783
rect 2278 787 2284 788
rect 2278 783 2279 787
rect 2283 783 2284 787
rect 2278 782 2284 783
rect 2414 787 2420 788
rect 2414 783 2415 787
rect 2419 783 2420 787
rect 2414 782 2420 783
rect 2526 787 2532 788
rect 2526 783 2527 787
rect 2531 783 2532 787
rect 2582 784 2583 788
rect 2587 784 2588 788
rect 2582 783 2588 784
rect 2526 782 2532 783
rect 1326 779 1332 780
rect 1206 778 1212 779
rect 382 749 388 750
rect 110 748 116 749
rect 110 744 111 748
rect 115 744 116 748
rect 382 745 383 749
rect 387 745 388 749
rect 382 744 388 745
rect 438 749 444 750
rect 438 745 439 749
rect 443 745 444 749
rect 438 744 444 745
rect 494 749 500 750
rect 494 745 495 749
rect 499 745 500 749
rect 494 744 500 745
rect 558 749 564 750
rect 558 745 559 749
rect 563 745 564 749
rect 558 744 564 745
rect 630 749 636 750
rect 630 745 631 749
rect 635 745 636 749
rect 630 744 636 745
rect 710 749 716 750
rect 710 745 711 749
rect 715 745 716 749
rect 710 744 716 745
rect 790 749 796 750
rect 790 745 791 749
rect 795 745 796 749
rect 790 744 796 745
rect 870 749 876 750
rect 870 745 871 749
rect 875 745 876 749
rect 870 744 876 745
rect 950 749 956 750
rect 950 745 951 749
rect 955 745 956 749
rect 950 744 956 745
rect 1038 749 1044 750
rect 1038 745 1039 749
rect 1043 745 1044 749
rect 1038 744 1044 745
rect 1126 749 1132 750
rect 1126 745 1127 749
rect 1131 745 1132 749
rect 1126 744 1132 745
rect 1326 748 1332 749
rect 1326 744 1327 748
rect 1331 744 1332 748
rect 1646 745 1652 746
rect 110 743 116 744
rect 1326 743 1332 744
rect 1366 744 1372 745
rect 1366 740 1367 744
rect 1371 740 1372 744
rect 1646 741 1647 745
rect 1651 741 1652 745
rect 1646 740 1652 741
rect 1702 745 1708 746
rect 1702 741 1703 745
rect 1707 741 1708 745
rect 1702 740 1708 741
rect 1758 745 1764 746
rect 1758 741 1759 745
rect 1763 741 1764 745
rect 1758 740 1764 741
rect 1814 745 1820 746
rect 1814 741 1815 745
rect 1819 741 1820 745
rect 1814 740 1820 741
rect 1870 745 1876 746
rect 1870 741 1871 745
rect 1875 741 1876 745
rect 1870 740 1876 741
rect 1926 745 1932 746
rect 1926 741 1927 745
rect 1931 741 1932 745
rect 1926 740 1932 741
rect 1990 745 1996 746
rect 1990 741 1991 745
rect 1995 741 1996 745
rect 1990 740 1996 741
rect 2062 745 2068 746
rect 2062 741 2063 745
rect 2067 741 2068 745
rect 2062 740 2068 741
rect 2142 745 2148 746
rect 2142 741 2143 745
rect 2147 741 2148 745
rect 2142 740 2148 741
rect 2230 745 2236 746
rect 2230 741 2231 745
rect 2235 741 2236 745
rect 2230 740 2236 741
rect 2334 745 2340 746
rect 2334 741 2335 745
rect 2339 741 2340 745
rect 2334 740 2340 741
rect 2438 745 2444 746
rect 2438 741 2439 745
rect 2443 741 2444 745
rect 2438 740 2444 741
rect 2526 745 2532 746
rect 2526 741 2527 745
rect 2531 741 2532 745
rect 2526 740 2532 741
rect 2582 744 2588 745
rect 2582 740 2583 744
rect 2587 740 2588 744
rect 1366 739 1372 740
rect 2582 739 2588 740
rect 110 731 116 732
rect 110 727 111 731
rect 115 727 116 731
rect 110 726 116 727
rect 1326 731 1332 732
rect 1326 727 1327 731
rect 1331 727 1332 731
rect 1326 726 1332 727
rect 1366 727 1372 728
rect 1366 723 1367 727
rect 1371 723 1372 727
rect 398 722 404 723
rect 398 718 399 722
rect 403 718 404 722
rect 398 717 404 718
rect 454 722 460 723
rect 454 718 455 722
rect 459 718 460 722
rect 454 717 460 718
rect 510 722 516 723
rect 510 718 511 722
rect 515 718 516 722
rect 510 717 516 718
rect 574 722 580 723
rect 574 718 575 722
rect 579 718 580 722
rect 574 717 580 718
rect 646 722 652 723
rect 646 718 647 722
rect 651 718 652 722
rect 646 717 652 718
rect 726 722 732 723
rect 726 718 727 722
rect 731 718 732 722
rect 726 717 732 718
rect 806 722 812 723
rect 806 718 807 722
rect 811 718 812 722
rect 806 717 812 718
rect 886 722 892 723
rect 886 718 887 722
rect 891 718 892 722
rect 886 717 892 718
rect 966 722 972 723
rect 966 718 967 722
rect 971 718 972 722
rect 966 717 972 718
rect 1054 722 1060 723
rect 1054 718 1055 722
rect 1059 718 1060 722
rect 1054 717 1060 718
rect 1142 722 1148 723
rect 1366 722 1372 723
rect 2582 727 2588 728
rect 2582 723 2583 727
rect 2587 723 2588 727
rect 2582 722 2588 723
rect 1142 718 1143 722
rect 1147 718 1148 722
rect 1142 717 1148 718
rect 1662 718 1668 719
rect 1662 714 1663 718
rect 1667 714 1668 718
rect 1662 713 1668 714
rect 1718 718 1724 719
rect 1718 714 1719 718
rect 1723 714 1724 718
rect 1718 713 1724 714
rect 1774 718 1780 719
rect 1774 714 1775 718
rect 1779 714 1780 718
rect 1774 713 1780 714
rect 1830 718 1836 719
rect 1830 714 1831 718
rect 1835 714 1836 718
rect 1830 713 1836 714
rect 1886 718 1892 719
rect 1886 714 1887 718
rect 1891 714 1892 718
rect 1886 713 1892 714
rect 1942 718 1948 719
rect 1942 714 1943 718
rect 1947 714 1948 718
rect 1942 713 1948 714
rect 2006 718 2012 719
rect 2006 714 2007 718
rect 2011 714 2012 718
rect 2006 713 2012 714
rect 2078 718 2084 719
rect 2078 714 2079 718
rect 2083 714 2084 718
rect 2078 713 2084 714
rect 2158 718 2164 719
rect 2158 714 2159 718
rect 2163 714 2164 718
rect 2158 713 2164 714
rect 2246 718 2252 719
rect 2246 714 2247 718
rect 2251 714 2252 718
rect 2246 713 2252 714
rect 2350 718 2356 719
rect 2350 714 2351 718
rect 2355 714 2356 718
rect 2350 713 2356 714
rect 2454 718 2460 719
rect 2454 714 2455 718
rect 2459 714 2460 718
rect 2454 713 2460 714
rect 2542 718 2548 719
rect 2542 714 2543 718
rect 2547 714 2548 718
rect 2542 713 2548 714
rect 342 698 348 699
rect 342 694 343 698
rect 347 694 348 698
rect 342 693 348 694
rect 414 698 420 699
rect 414 694 415 698
rect 419 694 420 698
rect 414 693 420 694
rect 486 698 492 699
rect 486 694 487 698
rect 491 694 492 698
rect 486 693 492 694
rect 558 698 564 699
rect 558 694 559 698
rect 563 694 564 698
rect 558 693 564 694
rect 630 698 636 699
rect 630 694 631 698
rect 635 694 636 698
rect 630 693 636 694
rect 694 698 700 699
rect 694 694 695 698
rect 699 694 700 698
rect 694 693 700 694
rect 758 698 764 699
rect 758 694 759 698
rect 763 694 764 698
rect 758 693 764 694
rect 822 698 828 699
rect 822 694 823 698
rect 827 694 828 698
rect 822 693 828 694
rect 886 698 892 699
rect 886 694 887 698
rect 891 694 892 698
rect 886 693 892 694
rect 950 698 956 699
rect 950 694 951 698
rect 955 694 956 698
rect 950 693 956 694
rect 1022 698 1028 699
rect 1022 694 1023 698
rect 1027 694 1028 698
rect 1022 693 1028 694
rect 1734 690 1740 691
rect 110 689 116 690
rect 110 685 111 689
rect 115 685 116 689
rect 110 684 116 685
rect 1326 689 1332 690
rect 1326 685 1327 689
rect 1331 685 1332 689
rect 1734 686 1735 690
rect 1739 686 1740 690
rect 1734 685 1740 686
rect 1790 690 1796 691
rect 1790 686 1791 690
rect 1795 686 1796 690
rect 1790 685 1796 686
rect 1854 690 1860 691
rect 1854 686 1855 690
rect 1859 686 1860 690
rect 1854 685 1860 686
rect 1918 690 1924 691
rect 1918 686 1919 690
rect 1923 686 1924 690
rect 1918 685 1924 686
rect 1990 690 1996 691
rect 1990 686 1991 690
rect 1995 686 1996 690
rect 1990 685 1996 686
rect 2062 690 2068 691
rect 2062 686 2063 690
rect 2067 686 2068 690
rect 2062 685 2068 686
rect 2126 690 2132 691
rect 2126 686 2127 690
rect 2131 686 2132 690
rect 2126 685 2132 686
rect 2198 690 2204 691
rect 2198 686 2199 690
rect 2203 686 2204 690
rect 2198 685 2204 686
rect 2270 690 2276 691
rect 2270 686 2271 690
rect 2275 686 2276 690
rect 2270 685 2276 686
rect 2342 690 2348 691
rect 2342 686 2343 690
rect 2347 686 2348 690
rect 2342 685 2348 686
rect 2414 690 2420 691
rect 2414 686 2415 690
rect 2419 686 2420 690
rect 2414 685 2420 686
rect 2486 690 2492 691
rect 2486 686 2487 690
rect 2491 686 2492 690
rect 2486 685 2492 686
rect 2542 690 2548 691
rect 2542 686 2543 690
rect 2547 686 2548 690
rect 2542 685 2548 686
rect 1326 684 1332 685
rect 1366 681 1372 682
rect 1366 677 1367 681
rect 1371 677 1372 681
rect 1366 676 1372 677
rect 2582 681 2588 682
rect 2582 677 2583 681
rect 2587 677 2588 681
rect 2582 676 2588 677
rect 110 672 116 673
rect 1326 672 1332 673
rect 110 668 111 672
rect 115 668 116 672
rect 110 667 116 668
rect 326 671 332 672
rect 326 667 327 671
rect 331 667 332 671
rect 326 666 332 667
rect 398 671 404 672
rect 398 667 399 671
rect 403 667 404 671
rect 398 666 404 667
rect 470 671 476 672
rect 470 667 471 671
rect 475 667 476 671
rect 470 666 476 667
rect 542 671 548 672
rect 542 667 543 671
rect 547 667 548 671
rect 542 666 548 667
rect 614 671 620 672
rect 614 667 615 671
rect 619 667 620 671
rect 614 666 620 667
rect 678 671 684 672
rect 678 667 679 671
rect 683 667 684 671
rect 678 666 684 667
rect 742 671 748 672
rect 742 667 743 671
rect 747 667 748 671
rect 742 666 748 667
rect 806 671 812 672
rect 806 667 807 671
rect 811 667 812 671
rect 806 666 812 667
rect 870 671 876 672
rect 870 667 871 671
rect 875 667 876 671
rect 870 666 876 667
rect 934 671 940 672
rect 934 667 935 671
rect 939 667 940 671
rect 934 666 940 667
rect 1006 671 1012 672
rect 1006 667 1007 671
rect 1011 667 1012 671
rect 1326 668 1327 672
rect 1331 668 1332 672
rect 1326 667 1332 668
rect 1006 666 1012 667
rect 1366 664 1372 665
rect 2582 664 2588 665
rect 1366 660 1367 664
rect 1371 660 1372 664
rect 1366 659 1372 660
rect 1718 663 1724 664
rect 1718 659 1719 663
rect 1723 659 1724 663
rect 1718 658 1724 659
rect 1774 663 1780 664
rect 1774 659 1775 663
rect 1779 659 1780 663
rect 1774 658 1780 659
rect 1838 663 1844 664
rect 1838 659 1839 663
rect 1843 659 1844 663
rect 1838 658 1844 659
rect 1902 663 1908 664
rect 1902 659 1903 663
rect 1907 659 1908 663
rect 1902 658 1908 659
rect 1974 663 1980 664
rect 1974 659 1975 663
rect 1979 659 1980 663
rect 1974 658 1980 659
rect 2046 663 2052 664
rect 2046 659 2047 663
rect 2051 659 2052 663
rect 2046 658 2052 659
rect 2110 663 2116 664
rect 2110 659 2111 663
rect 2115 659 2116 663
rect 2110 658 2116 659
rect 2182 663 2188 664
rect 2182 659 2183 663
rect 2187 659 2188 663
rect 2182 658 2188 659
rect 2254 663 2260 664
rect 2254 659 2255 663
rect 2259 659 2260 663
rect 2254 658 2260 659
rect 2326 663 2332 664
rect 2326 659 2327 663
rect 2331 659 2332 663
rect 2326 658 2332 659
rect 2398 663 2404 664
rect 2398 659 2399 663
rect 2403 659 2404 663
rect 2398 658 2404 659
rect 2470 663 2476 664
rect 2470 659 2471 663
rect 2475 659 2476 663
rect 2470 658 2476 659
rect 2526 663 2532 664
rect 2526 659 2527 663
rect 2531 659 2532 663
rect 2582 660 2583 664
rect 2587 660 2588 664
rect 2582 659 2588 660
rect 2526 658 2532 659
rect 230 633 236 634
rect 110 632 116 633
rect 110 628 111 632
rect 115 628 116 632
rect 230 629 231 633
rect 235 629 236 633
rect 230 628 236 629
rect 294 633 300 634
rect 294 629 295 633
rect 299 629 300 633
rect 294 628 300 629
rect 358 633 364 634
rect 358 629 359 633
rect 363 629 364 633
rect 358 628 364 629
rect 422 633 428 634
rect 422 629 423 633
rect 427 629 428 633
rect 422 628 428 629
rect 478 633 484 634
rect 478 629 479 633
rect 483 629 484 633
rect 478 628 484 629
rect 534 633 540 634
rect 534 629 535 633
rect 539 629 540 633
rect 534 628 540 629
rect 598 633 604 634
rect 598 629 599 633
rect 603 629 604 633
rect 598 628 604 629
rect 662 633 668 634
rect 662 629 663 633
rect 667 629 668 633
rect 662 628 668 629
rect 726 633 732 634
rect 726 629 727 633
rect 731 629 732 633
rect 726 628 732 629
rect 790 633 796 634
rect 790 629 791 633
rect 795 629 796 633
rect 790 628 796 629
rect 854 633 860 634
rect 854 629 855 633
rect 859 629 860 633
rect 854 628 860 629
rect 918 633 924 634
rect 918 629 919 633
rect 923 629 924 633
rect 918 628 924 629
rect 1326 632 1332 633
rect 1326 628 1327 632
rect 1331 628 1332 632
rect 110 627 116 628
rect 1326 627 1332 628
rect 1614 625 1620 626
rect 1366 624 1372 625
rect 1366 620 1367 624
rect 1371 620 1372 624
rect 1614 621 1615 625
rect 1619 621 1620 625
rect 1614 620 1620 621
rect 1678 625 1684 626
rect 1678 621 1679 625
rect 1683 621 1684 625
rect 1678 620 1684 621
rect 1758 625 1764 626
rect 1758 621 1759 625
rect 1763 621 1764 625
rect 1758 620 1764 621
rect 1838 625 1844 626
rect 1838 621 1839 625
rect 1843 621 1844 625
rect 1838 620 1844 621
rect 1926 625 1932 626
rect 1926 621 1927 625
rect 1931 621 1932 625
rect 1926 620 1932 621
rect 2014 625 2020 626
rect 2014 621 2015 625
rect 2019 621 2020 625
rect 2014 620 2020 621
rect 2094 625 2100 626
rect 2094 621 2095 625
rect 2099 621 2100 625
rect 2094 620 2100 621
rect 2174 625 2180 626
rect 2174 621 2175 625
rect 2179 621 2180 625
rect 2174 620 2180 621
rect 2254 625 2260 626
rect 2254 621 2255 625
rect 2259 621 2260 625
rect 2254 620 2260 621
rect 2326 625 2332 626
rect 2326 621 2327 625
rect 2331 621 2332 625
rect 2326 620 2332 621
rect 2398 625 2404 626
rect 2398 621 2399 625
rect 2403 621 2404 625
rect 2398 620 2404 621
rect 2470 625 2476 626
rect 2470 621 2471 625
rect 2475 621 2476 625
rect 2470 620 2476 621
rect 2526 625 2532 626
rect 2526 621 2527 625
rect 2531 621 2532 625
rect 2526 620 2532 621
rect 2582 624 2588 625
rect 2582 620 2583 624
rect 2587 620 2588 624
rect 1366 619 1372 620
rect 2582 619 2588 620
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 110 610 116 611
rect 1326 615 1332 616
rect 1326 611 1327 615
rect 1331 611 1332 615
rect 1326 610 1332 611
rect 1366 607 1372 608
rect 246 606 252 607
rect 246 602 247 606
rect 251 602 252 606
rect 246 601 252 602
rect 310 606 316 607
rect 310 602 311 606
rect 315 602 316 606
rect 310 601 316 602
rect 374 606 380 607
rect 374 602 375 606
rect 379 602 380 606
rect 374 601 380 602
rect 438 606 444 607
rect 438 602 439 606
rect 443 602 444 606
rect 438 601 444 602
rect 494 606 500 607
rect 494 602 495 606
rect 499 602 500 606
rect 494 601 500 602
rect 550 606 556 607
rect 550 602 551 606
rect 555 602 556 606
rect 550 601 556 602
rect 614 606 620 607
rect 614 602 615 606
rect 619 602 620 606
rect 614 601 620 602
rect 678 606 684 607
rect 678 602 679 606
rect 683 602 684 606
rect 678 601 684 602
rect 742 606 748 607
rect 742 602 743 606
rect 747 602 748 606
rect 742 601 748 602
rect 806 606 812 607
rect 806 602 807 606
rect 811 602 812 606
rect 806 601 812 602
rect 870 606 876 607
rect 870 602 871 606
rect 875 602 876 606
rect 870 601 876 602
rect 934 606 940 607
rect 934 602 935 606
rect 939 602 940 606
rect 1366 603 1367 607
rect 1371 603 1372 607
rect 1366 602 1372 603
rect 2582 607 2588 608
rect 2582 603 2583 607
rect 2587 603 2588 607
rect 2582 602 2588 603
rect 934 601 940 602
rect 1630 598 1636 599
rect 1630 594 1631 598
rect 1635 594 1636 598
rect 1630 593 1636 594
rect 1694 598 1700 599
rect 1694 594 1695 598
rect 1699 594 1700 598
rect 1694 593 1700 594
rect 1774 598 1780 599
rect 1774 594 1775 598
rect 1779 594 1780 598
rect 1774 593 1780 594
rect 1854 598 1860 599
rect 1854 594 1855 598
rect 1859 594 1860 598
rect 1854 593 1860 594
rect 1942 598 1948 599
rect 1942 594 1943 598
rect 1947 594 1948 598
rect 1942 593 1948 594
rect 2030 598 2036 599
rect 2030 594 2031 598
rect 2035 594 2036 598
rect 2030 593 2036 594
rect 2110 598 2116 599
rect 2110 594 2111 598
rect 2115 594 2116 598
rect 2110 593 2116 594
rect 2190 598 2196 599
rect 2190 594 2191 598
rect 2195 594 2196 598
rect 2190 593 2196 594
rect 2270 598 2276 599
rect 2270 594 2271 598
rect 2275 594 2276 598
rect 2270 593 2276 594
rect 2342 598 2348 599
rect 2342 594 2343 598
rect 2347 594 2348 598
rect 2342 593 2348 594
rect 2414 598 2420 599
rect 2414 594 2415 598
rect 2419 594 2420 598
rect 2414 593 2420 594
rect 2486 598 2492 599
rect 2486 594 2487 598
rect 2491 594 2492 598
rect 2486 593 2492 594
rect 2542 598 2548 599
rect 2542 594 2543 598
rect 2547 594 2548 598
rect 2542 593 2548 594
rect 190 574 196 575
rect 190 570 191 574
rect 195 570 196 574
rect 190 569 196 570
rect 278 574 284 575
rect 278 570 279 574
rect 283 570 284 574
rect 278 569 284 570
rect 366 574 372 575
rect 366 570 367 574
rect 371 570 372 574
rect 366 569 372 570
rect 462 574 468 575
rect 462 570 463 574
rect 467 570 468 574
rect 462 569 468 570
rect 558 574 564 575
rect 558 570 559 574
rect 563 570 564 574
rect 558 569 564 570
rect 646 574 652 575
rect 646 570 647 574
rect 651 570 652 574
rect 646 569 652 570
rect 734 574 740 575
rect 734 570 735 574
rect 739 570 740 574
rect 734 569 740 570
rect 814 574 820 575
rect 814 570 815 574
rect 819 570 820 574
rect 814 569 820 570
rect 886 574 892 575
rect 886 570 887 574
rect 891 570 892 574
rect 886 569 892 570
rect 966 574 972 575
rect 966 570 967 574
rect 971 570 972 574
rect 966 569 972 570
rect 1046 574 1052 575
rect 1046 570 1047 574
rect 1051 570 1052 574
rect 1046 569 1052 570
rect 1126 574 1132 575
rect 1126 570 1127 574
rect 1131 570 1132 574
rect 1126 569 1132 570
rect 1510 566 1516 567
rect 110 565 116 566
rect 110 561 111 565
rect 115 561 116 565
rect 110 560 116 561
rect 1326 565 1332 566
rect 1326 561 1327 565
rect 1331 561 1332 565
rect 1510 562 1511 566
rect 1515 562 1516 566
rect 1510 561 1516 562
rect 1574 566 1580 567
rect 1574 562 1575 566
rect 1579 562 1580 566
rect 1574 561 1580 562
rect 1654 566 1660 567
rect 1654 562 1655 566
rect 1659 562 1660 566
rect 1654 561 1660 562
rect 1734 566 1740 567
rect 1734 562 1735 566
rect 1739 562 1740 566
rect 1734 561 1740 562
rect 1822 566 1828 567
rect 1822 562 1823 566
rect 1827 562 1828 566
rect 1822 561 1828 562
rect 1910 566 1916 567
rect 1910 562 1911 566
rect 1915 562 1916 566
rect 1910 561 1916 562
rect 1998 566 2004 567
rect 1998 562 1999 566
rect 2003 562 2004 566
rect 1998 561 2004 562
rect 2086 566 2092 567
rect 2086 562 2087 566
rect 2091 562 2092 566
rect 2086 561 2092 562
rect 2174 566 2180 567
rect 2174 562 2175 566
rect 2179 562 2180 566
rect 2174 561 2180 562
rect 2270 566 2276 567
rect 2270 562 2271 566
rect 2275 562 2276 566
rect 2270 561 2276 562
rect 2366 566 2372 567
rect 2366 562 2367 566
rect 2371 562 2372 566
rect 2366 561 2372 562
rect 2462 566 2468 567
rect 2462 562 2463 566
rect 2467 562 2468 566
rect 2462 561 2468 562
rect 2542 566 2548 567
rect 2542 562 2543 566
rect 2547 562 2548 566
rect 2542 561 2548 562
rect 1326 560 1332 561
rect 1366 557 1372 558
rect 1366 553 1367 557
rect 1371 553 1372 557
rect 1366 552 1372 553
rect 2582 557 2588 558
rect 2582 553 2583 557
rect 2587 553 2588 557
rect 2582 552 2588 553
rect 110 548 116 549
rect 1326 548 1332 549
rect 110 544 111 548
rect 115 544 116 548
rect 110 543 116 544
rect 174 547 180 548
rect 174 543 175 547
rect 179 543 180 547
rect 174 542 180 543
rect 262 547 268 548
rect 262 543 263 547
rect 267 543 268 547
rect 262 542 268 543
rect 350 547 356 548
rect 350 543 351 547
rect 355 543 356 547
rect 350 542 356 543
rect 446 547 452 548
rect 446 543 447 547
rect 451 543 452 547
rect 446 542 452 543
rect 542 547 548 548
rect 542 543 543 547
rect 547 543 548 547
rect 542 542 548 543
rect 630 547 636 548
rect 630 543 631 547
rect 635 543 636 547
rect 630 542 636 543
rect 718 547 724 548
rect 718 543 719 547
rect 723 543 724 547
rect 718 542 724 543
rect 798 547 804 548
rect 798 543 799 547
rect 803 543 804 547
rect 798 542 804 543
rect 870 547 876 548
rect 870 543 871 547
rect 875 543 876 547
rect 870 542 876 543
rect 950 547 956 548
rect 950 543 951 547
rect 955 543 956 547
rect 950 542 956 543
rect 1030 547 1036 548
rect 1030 543 1031 547
rect 1035 543 1036 547
rect 1030 542 1036 543
rect 1110 547 1116 548
rect 1110 543 1111 547
rect 1115 543 1116 547
rect 1326 544 1327 548
rect 1331 544 1332 548
rect 1326 543 1332 544
rect 1110 542 1116 543
rect 1366 540 1372 541
rect 2582 540 2588 541
rect 1366 536 1367 540
rect 1371 536 1372 540
rect 1366 535 1372 536
rect 1494 539 1500 540
rect 1494 535 1495 539
rect 1499 535 1500 539
rect 1494 534 1500 535
rect 1558 539 1564 540
rect 1558 535 1559 539
rect 1563 535 1564 539
rect 1558 534 1564 535
rect 1638 539 1644 540
rect 1638 535 1639 539
rect 1643 535 1644 539
rect 1638 534 1644 535
rect 1718 539 1724 540
rect 1718 535 1719 539
rect 1723 535 1724 539
rect 1718 534 1724 535
rect 1806 539 1812 540
rect 1806 535 1807 539
rect 1811 535 1812 539
rect 1806 534 1812 535
rect 1894 539 1900 540
rect 1894 535 1895 539
rect 1899 535 1900 539
rect 1894 534 1900 535
rect 1982 539 1988 540
rect 1982 535 1983 539
rect 1987 535 1988 539
rect 1982 534 1988 535
rect 2070 539 2076 540
rect 2070 535 2071 539
rect 2075 535 2076 539
rect 2070 534 2076 535
rect 2158 539 2164 540
rect 2158 535 2159 539
rect 2163 535 2164 539
rect 2158 534 2164 535
rect 2254 539 2260 540
rect 2254 535 2255 539
rect 2259 535 2260 539
rect 2254 534 2260 535
rect 2350 539 2356 540
rect 2350 535 2351 539
rect 2355 535 2356 539
rect 2350 534 2356 535
rect 2446 539 2452 540
rect 2446 535 2447 539
rect 2451 535 2452 539
rect 2446 534 2452 535
rect 2526 539 2532 540
rect 2526 535 2527 539
rect 2531 535 2532 539
rect 2582 536 2583 540
rect 2587 536 2588 540
rect 2582 535 2588 536
rect 2526 534 2532 535
rect 142 509 148 510
rect 110 508 116 509
rect 110 504 111 508
rect 115 504 116 508
rect 142 505 143 509
rect 147 505 148 509
rect 142 504 148 505
rect 206 509 212 510
rect 206 505 207 509
rect 211 505 212 509
rect 206 504 212 505
rect 310 509 316 510
rect 310 505 311 509
rect 315 505 316 509
rect 310 504 316 505
rect 430 509 436 510
rect 430 505 431 509
rect 435 505 436 509
rect 430 504 436 505
rect 550 509 556 510
rect 550 505 551 509
rect 555 505 556 509
rect 550 504 556 505
rect 670 509 676 510
rect 670 505 671 509
rect 675 505 676 509
rect 670 504 676 505
rect 790 509 796 510
rect 790 505 791 509
rect 795 505 796 509
rect 790 504 796 505
rect 902 509 908 510
rect 902 505 903 509
rect 907 505 908 509
rect 902 504 908 505
rect 1006 509 1012 510
rect 1006 505 1007 509
rect 1011 505 1012 509
rect 1006 504 1012 505
rect 1102 509 1108 510
rect 1102 505 1103 509
rect 1107 505 1108 509
rect 1102 504 1108 505
rect 1198 509 1204 510
rect 1198 505 1199 509
rect 1203 505 1204 509
rect 1198 504 1204 505
rect 1270 509 1276 510
rect 1270 505 1271 509
rect 1275 505 1276 509
rect 1270 504 1276 505
rect 1326 508 1332 509
rect 1326 504 1327 508
rect 1331 504 1332 508
rect 110 503 116 504
rect 1326 503 1332 504
rect 1398 501 1404 502
rect 1366 500 1372 501
rect 1366 496 1367 500
rect 1371 496 1372 500
rect 1398 497 1399 501
rect 1403 497 1404 501
rect 1398 496 1404 497
rect 1454 501 1460 502
rect 1454 497 1455 501
rect 1459 497 1460 501
rect 1454 496 1460 497
rect 1518 501 1524 502
rect 1518 497 1519 501
rect 1523 497 1524 501
rect 1518 496 1524 497
rect 1606 501 1612 502
rect 1606 497 1607 501
rect 1611 497 1612 501
rect 1606 496 1612 497
rect 1694 501 1700 502
rect 1694 497 1695 501
rect 1699 497 1700 501
rect 1694 496 1700 497
rect 1790 501 1796 502
rect 1790 497 1791 501
rect 1795 497 1796 501
rect 1790 496 1796 497
rect 1886 501 1892 502
rect 1886 497 1887 501
rect 1891 497 1892 501
rect 1886 496 1892 497
rect 1982 501 1988 502
rect 1982 497 1983 501
rect 1987 497 1988 501
rect 1982 496 1988 497
rect 2086 501 2092 502
rect 2086 497 2087 501
rect 2091 497 2092 501
rect 2086 496 2092 497
rect 2198 501 2204 502
rect 2198 497 2199 501
rect 2203 497 2204 501
rect 2198 496 2204 497
rect 2310 501 2316 502
rect 2310 497 2311 501
rect 2315 497 2316 501
rect 2310 496 2316 497
rect 2430 501 2436 502
rect 2430 497 2431 501
rect 2435 497 2436 501
rect 2430 496 2436 497
rect 2526 501 2532 502
rect 2526 497 2527 501
rect 2531 497 2532 501
rect 2526 496 2532 497
rect 2582 500 2588 501
rect 2582 496 2583 500
rect 2587 496 2588 500
rect 1366 495 1372 496
rect 2582 495 2588 496
rect 110 491 116 492
rect 110 487 111 491
rect 115 487 116 491
rect 110 486 116 487
rect 1326 491 1332 492
rect 1326 487 1327 491
rect 1331 487 1332 491
rect 1326 486 1332 487
rect 1366 483 1372 484
rect 158 482 164 483
rect 158 478 159 482
rect 163 478 164 482
rect 158 477 164 478
rect 222 482 228 483
rect 222 478 223 482
rect 227 478 228 482
rect 222 477 228 478
rect 326 482 332 483
rect 326 478 327 482
rect 331 478 332 482
rect 326 477 332 478
rect 446 482 452 483
rect 446 478 447 482
rect 451 478 452 482
rect 446 477 452 478
rect 566 482 572 483
rect 566 478 567 482
rect 571 478 572 482
rect 566 477 572 478
rect 686 482 692 483
rect 686 478 687 482
rect 691 478 692 482
rect 686 477 692 478
rect 806 482 812 483
rect 806 478 807 482
rect 811 478 812 482
rect 806 477 812 478
rect 918 482 924 483
rect 918 478 919 482
rect 923 478 924 482
rect 918 477 924 478
rect 1022 482 1028 483
rect 1022 478 1023 482
rect 1027 478 1028 482
rect 1022 477 1028 478
rect 1118 482 1124 483
rect 1118 478 1119 482
rect 1123 478 1124 482
rect 1118 477 1124 478
rect 1214 482 1220 483
rect 1214 478 1215 482
rect 1219 478 1220 482
rect 1214 477 1220 478
rect 1286 482 1292 483
rect 1286 478 1287 482
rect 1291 478 1292 482
rect 1366 479 1367 483
rect 1371 479 1372 483
rect 1366 478 1372 479
rect 2582 483 2588 484
rect 2582 479 2583 483
rect 2587 479 2588 483
rect 2582 478 2588 479
rect 1286 477 1292 478
rect 1414 474 1420 475
rect 1414 470 1415 474
rect 1419 470 1420 474
rect 1414 469 1420 470
rect 1470 474 1476 475
rect 1470 470 1471 474
rect 1475 470 1476 474
rect 1470 469 1476 470
rect 1534 474 1540 475
rect 1534 470 1535 474
rect 1539 470 1540 474
rect 1534 469 1540 470
rect 1622 474 1628 475
rect 1622 470 1623 474
rect 1627 470 1628 474
rect 1622 469 1628 470
rect 1710 474 1716 475
rect 1710 470 1711 474
rect 1715 470 1716 474
rect 1710 469 1716 470
rect 1806 474 1812 475
rect 1806 470 1807 474
rect 1811 470 1812 474
rect 1806 469 1812 470
rect 1902 474 1908 475
rect 1902 470 1903 474
rect 1907 470 1908 474
rect 1902 469 1908 470
rect 1998 474 2004 475
rect 1998 470 1999 474
rect 2003 470 2004 474
rect 1998 469 2004 470
rect 2102 474 2108 475
rect 2102 470 2103 474
rect 2107 470 2108 474
rect 2102 469 2108 470
rect 2214 474 2220 475
rect 2214 470 2215 474
rect 2219 470 2220 474
rect 2214 469 2220 470
rect 2326 474 2332 475
rect 2326 470 2327 474
rect 2331 470 2332 474
rect 2326 469 2332 470
rect 2446 474 2452 475
rect 2446 470 2447 474
rect 2451 470 2452 474
rect 2446 469 2452 470
rect 2542 474 2548 475
rect 2542 470 2543 474
rect 2547 470 2548 474
rect 2542 469 2548 470
rect 158 454 164 455
rect 158 450 159 454
rect 163 450 164 454
rect 158 449 164 450
rect 222 454 228 455
rect 222 450 223 454
rect 227 450 228 454
rect 222 449 228 450
rect 318 454 324 455
rect 318 450 319 454
rect 323 450 324 454
rect 318 449 324 450
rect 422 454 428 455
rect 422 450 423 454
rect 427 450 428 454
rect 422 449 428 450
rect 534 454 540 455
rect 534 450 535 454
rect 539 450 540 454
rect 534 449 540 450
rect 638 454 644 455
rect 638 450 639 454
rect 643 450 644 454
rect 638 449 644 450
rect 742 454 748 455
rect 742 450 743 454
rect 747 450 748 454
rect 742 449 748 450
rect 838 454 844 455
rect 838 450 839 454
rect 843 450 844 454
rect 838 449 844 450
rect 926 454 932 455
rect 926 450 927 454
rect 931 450 932 454
rect 926 449 932 450
rect 1006 454 1012 455
rect 1006 450 1007 454
rect 1011 450 1012 454
rect 1006 449 1012 450
rect 1078 454 1084 455
rect 1078 450 1079 454
rect 1083 450 1084 454
rect 1078 449 1084 450
rect 1150 454 1156 455
rect 1150 450 1151 454
rect 1155 450 1156 454
rect 1150 449 1156 450
rect 1230 454 1236 455
rect 1230 450 1231 454
rect 1235 450 1236 454
rect 1230 449 1236 450
rect 1286 454 1292 455
rect 1286 450 1287 454
rect 1291 450 1292 454
rect 1286 449 1292 450
rect 110 445 116 446
rect 110 441 111 445
rect 115 441 116 445
rect 110 440 116 441
rect 1326 445 1332 446
rect 1326 441 1327 445
rect 1331 441 1332 445
rect 1326 440 1332 441
rect 1414 442 1420 443
rect 1414 438 1415 442
rect 1419 438 1420 442
rect 1414 437 1420 438
rect 1486 442 1492 443
rect 1486 438 1487 442
rect 1491 438 1492 442
rect 1486 437 1492 438
rect 1574 442 1580 443
rect 1574 438 1575 442
rect 1579 438 1580 442
rect 1574 437 1580 438
rect 1662 442 1668 443
rect 1662 438 1663 442
rect 1667 438 1668 442
rect 1662 437 1668 438
rect 1758 442 1764 443
rect 1758 438 1759 442
rect 1763 438 1764 442
rect 1758 437 1764 438
rect 1862 442 1868 443
rect 1862 438 1863 442
rect 1867 438 1868 442
rect 1862 437 1868 438
rect 1974 442 1980 443
rect 1974 438 1975 442
rect 1979 438 1980 442
rect 1974 437 1980 438
rect 2110 442 2116 443
rect 2110 438 2111 442
rect 2115 438 2116 442
rect 2110 437 2116 438
rect 2254 442 2260 443
rect 2254 438 2255 442
rect 2259 438 2260 442
rect 2254 437 2260 438
rect 2406 442 2412 443
rect 2406 438 2407 442
rect 2411 438 2412 442
rect 2406 437 2412 438
rect 2542 442 2548 443
rect 2542 438 2543 442
rect 2547 438 2548 442
rect 2542 437 2548 438
rect 1366 433 1372 434
rect 1366 429 1367 433
rect 1371 429 1372 433
rect 110 428 116 429
rect 1326 428 1332 429
rect 1366 428 1372 429
rect 2582 433 2588 434
rect 2582 429 2583 433
rect 2587 429 2588 433
rect 2582 428 2588 429
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 142 427 148 428
rect 142 423 143 427
rect 147 423 148 427
rect 142 422 148 423
rect 206 427 212 428
rect 206 423 207 427
rect 211 423 212 427
rect 206 422 212 423
rect 302 427 308 428
rect 302 423 303 427
rect 307 423 308 427
rect 302 422 308 423
rect 406 427 412 428
rect 406 423 407 427
rect 411 423 412 427
rect 406 422 412 423
rect 518 427 524 428
rect 518 423 519 427
rect 523 423 524 427
rect 518 422 524 423
rect 622 427 628 428
rect 622 423 623 427
rect 627 423 628 427
rect 622 422 628 423
rect 726 427 732 428
rect 726 423 727 427
rect 731 423 732 427
rect 726 422 732 423
rect 822 427 828 428
rect 822 423 823 427
rect 827 423 828 427
rect 822 422 828 423
rect 910 427 916 428
rect 910 423 911 427
rect 915 423 916 427
rect 910 422 916 423
rect 990 427 996 428
rect 990 423 991 427
rect 995 423 996 427
rect 990 422 996 423
rect 1062 427 1068 428
rect 1062 423 1063 427
rect 1067 423 1068 427
rect 1062 422 1068 423
rect 1134 427 1140 428
rect 1134 423 1135 427
rect 1139 423 1140 427
rect 1134 422 1140 423
rect 1214 427 1220 428
rect 1214 423 1215 427
rect 1219 423 1220 427
rect 1214 422 1220 423
rect 1270 427 1276 428
rect 1270 423 1271 427
rect 1275 423 1276 427
rect 1326 424 1327 428
rect 1331 424 1332 428
rect 1326 423 1332 424
rect 1270 422 1276 423
rect 1366 416 1372 417
rect 2582 416 2588 417
rect 1366 412 1367 416
rect 1371 412 1372 416
rect 1366 411 1372 412
rect 1398 415 1404 416
rect 1398 411 1399 415
rect 1403 411 1404 415
rect 1398 410 1404 411
rect 1470 415 1476 416
rect 1470 411 1471 415
rect 1475 411 1476 415
rect 1470 410 1476 411
rect 1558 415 1564 416
rect 1558 411 1559 415
rect 1563 411 1564 415
rect 1558 410 1564 411
rect 1646 415 1652 416
rect 1646 411 1647 415
rect 1651 411 1652 415
rect 1646 410 1652 411
rect 1742 415 1748 416
rect 1742 411 1743 415
rect 1747 411 1748 415
rect 1742 410 1748 411
rect 1846 415 1852 416
rect 1846 411 1847 415
rect 1851 411 1852 415
rect 1846 410 1852 411
rect 1958 415 1964 416
rect 1958 411 1959 415
rect 1963 411 1964 415
rect 1958 410 1964 411
rect 2094 415 2100 416
rect 2094 411 2095 415
rect 2099 411 2100 415
rect 2094 410 2100 411
rect 2238 415 2244 416
rect 2238 411 2239 415
rect 2243 411 2244 415
rect 2238 410 2244 411
rect 2390 415 2396 416
rect 2390 411 2391 415
rect 2395 411 2396 415
rect 2390 410 2396 411
rect 2526 415 2532 416
rect 2526 411 2527 415
rect 2531 411 2532 415
rect 2582 412 2583 416
rect 2587 412 2588 416
rect 2582 411 2588 412
rect 2526 410 2532 411
rect 142 385 148 386
rect 110 384 116 385
rect 110 380 111 384
rect 115 380 116 384
rect 142 381 143 385
rect 147 381 148 385
rect 142 380 148 381
rect 206 385 212 386
rect 206 381 207 385
rect 211 381 212 385
rect 206 380 212 381
rect 302 385 308 386
rect 302 381 303 385
rect 307 381 308 385
rect 302 380 308 381
rect 398 385 404 386
rect 398 381 399 385
rect 403 381 404 385
rect 398 380 404 381
rect 494 385 500 386
rect 494 381 495 385
rect 499 381 500 385
rect 494 380 500 381
rect 582 385 588 386
rect 582 381 583 385
rect 587 381 588 385
rect 582 380 588 381
rect 670 385 676 386
rect 670 381 671 385
rect 675 381 676 385
rect 670 380 676 381
rect 750 385 756 386
rect 750 381 751 385
rect 755 381 756 385
rect 750 380 756 381
rect 822 385 828 386
rect 822 381 823 385
rect 827 381 828 385
rect 822 380 828 381
rect 894 385 900 386
rect 894 381 895 385
rect 899 381 900 385
rect 894 380 900 381
rect 966 385 972 386
rect 966 381 967 385
rect 971 381 972 385
rect 966 380 972 381
rect 1046 385 1052 386
rect 1046 381 1047 385
rect 1051 381 1052 385
rect 1046 380 1052 381
rect 1326 384 1332 385
rect 1326 380 1327 384
rect 1331 380 1332 384
rect 110 379 116 380
rect 1326 379 1332 380
rect 1398 377 1404 378
rect 1366 376 1372 377
rect 1366 372 1367 376
rect 1371 372 1372 376
rect 1398 373 1399 377
rect 1403 373 1404 377
rect 1398 372 1404 373
rect 1454 377 1460 378
rect 1454 373 1455 377
rect 1459 373 1460 377
rect 1454 372 1460 373
rect 1510 377 1516 378
rect 1510 373 1511 377
rect 1515 373 1516 377
rect 1510 372 1516 373
rect 1566 377 1572 378
rect 1566 373 1567 377
rect 1571 373 1572 377
rect 1566 372 1572 373
rect 1630 377 1636 378
rect 1630 373 1631 377
rect 1635 373 1636 377
rect 1630 372 1636 373
rect 1694 377 1700 378
rect 1694 373 1695 377
rect 1699 373 1700 377
rect 1694 372 1700 373
rect 1758 377 1764 378
rect 1758 373 1759 377
rect 1763 373 1764 377
rect 1758 372 1764 373
rect 1838 377 1844 378
rect 1838 373 1839 377
rect 1843 373 1844 377
rect 1838 372 1844 373
rect 1942 377 1948 378
rect 1942 373 1943 377
rect 1947 373 1948 377
rect 1942 372 1948 373
rect 2070 377 2076 378
rect 2070 373 2071 377
rect 2075 373 2076 377
rect 2070 372 2076 373
rect 2214 377 2220 378
rect 2214 373 2215 377
rect 2219 373 2220 377
rect 2214 372 2220 373
rect 2366 377 2372 378
rect 2366 373 2367 377
rect 2371 373 2372 377
rect 2366 372 2372 373
rect 2526 377 2532 378
rect 2526 373 2527 377
rect 2531 373 2532 377
rect 2526 372 2532 373
rect 2582 376 2588 377
rect 2582 372 2583 376
rect 2587 372 2588 376
rect 1366 371 1372 372
rect 2582 371 2588 372
rect 110 367 116 368
rect 110 363 111 367
rect 115 363 116 367
rect 110 362 116 363
rect 1326 367 1332 368
rect 1326 363 1327 367
rect 1331 363 1332 367
rect 1326 362 1332 363
rect 1366 359 1372 360
rect 158 358 164 359
rect 158 354 159 358
rect 163 354 164 358
rect 158 353 164 354
rect 222 358 228 359
rect 222 354 223 358
rect 227 354 228 358
rect 222 353 228 354
rect 318 358 324 359
rect 318 354 319 358
rect 323 354 324 358
rect 318 353 324 354
rect 414 358 420 359
rect 414 354 415 358
rect 419 354 420 358
rect 414 353 420 354
rect 510 358 516 359
rect 510 354 511 358
rect 515 354 516 358
rect 510 353 516 354
rect 598 358 604 359
rect 598 354 599 358
rect 603 354 604 358
rect 598 353 604 354
rect 686 358 692 359
rect 686 354 687 358
rect 691 354 692 358
rect 686 353 692 354
rect 766 358 772 359
rect 766 354 767 358
rect 771 354 772 358
rect 766 353 772 354
rect 838 358 844 359
rect 838 354 839 358
rect 843 354 844 358
rect 838 353 844 354
rect 910 358 916 359
rect 910 354 911 358
rect 915 354 916 358
rect 910 353 916 354
rect 982 358 988 359
rect 982 354 983 358
rect 987 354 988 358
rect 982 353 988 354
rect 1062 358 1068 359
rect 1062 354 1063 358
rect 1067 354 1068 358
rect 1366 355 1367 359
rect 1371 355 1372 359
rect 1366 354 1372 355
rect 2582 359 2588 360
rect 2582 355 2583 359
rect 2587 355 2588 359
rect 2582 354 2588 355
rect 1062 353 1068 354
rect 1414 350 1420 351
rect 1414 346 1415 350
rect 1419 346 1420 350
rect 1414 345 1420 346
rect 1470 350 1476 351
rect 1470 346 1471 350
rect 1475 346 1476 350
rect 1470 345 1476 346
rect 1526 350 1532 351
rect 1526 346 1527 350
rect 1531 346 1532 350
rect 1526 345 1532 346
rect 1582 350 1588 351
rect 1582 346 1583 350
rect 1587 346 1588 350
rect 1582 345 1588 346
rect 1646 350 1652 351
rect 1646 346 1647 350
rect 1651 346 1652 350
rect 1646 345 1652 346
rect 1710 350 1716 351
rect 1710 346 1711 350
rect 1715 346 1716 350
rect 1710 345 1716 346
rect 1774 350 1780 351
rect 1774 346 1775 350
rect 1779 346 1780 350
rect 1774 345 1780 346
rect 1854 350 1860 351
rect 1854 346 1855 350
rect 1859 346 1860 350
rect 1854 345 1860 346
rect 1958 350 1964 351
rect 1958 346 1959 350
rect 1963 346 1964 350
rect 1958 345 1964 346
rect 2086 350 2092 351
rect 2086 346 2087 350
rect 2091 346 2092 350
rect 2086 345 2092 346
rect 2230 350 2236 351
rect 2230 346 2231 350
rect 2235 346 2236 350
rect 2230 345 2236 346
rect 2382 350 2388 351
rect 2382 346 2383 350
rect 2387 346 2388 350
rect 2382 345 2388 346
rect 2542 350 2548 351
rect 2542 346 2543 350
rect 2547 346 2548 350
rect 2542 345 2548 346
rect 158 330 164 331
rect 158 326 159 330
rect 163 326 164 330
rect 158 325 164 326
rect 222 330 228 331
rect 222 326 223 330
rect 227 326 228 330
rect 222 325 228 326
rect 310 330 316 331
rect 310 326 311 330
rect 315 326 316 330
rect 310 325 316 326
rect 390 330 396 331
rect 390 326 391 330
rect 395 326 396 330
rect 390 325 396 326
rect 470 330 476 331
rect 470 326 471 330
rect 475 326 476 330
rect 470 325 476 326
rect 542 330 548 331
rect 542 326 543 330
rect 547 326 548 330
rect 542 325 548 326
rect 606 330 612 331
rect 606 326 607 330
rect 611 326 612 330
rect 606 325 612 326
rect 670 330 676 331
rect 670 326 671 330
rect 675 326 676 330
rect 670 325 676 326
rect 734 330 740 331
rect 734 326 735 330
rect 739 326 740 330
rect 734 325 740 326
rect 798 330 804 331
rect 798 326 799 330
rect 803 326 804 330
rect 798 325 804 326
rect 862 330 868 331
rect 862 326 863 330
rect 867 326 868 330
rect 862 325 868 326
rect 934 330 940 331
rect 934 326 935 330
rect 939 326 940 330
rect 934 325 940 326
rect 1606 322 1612 323
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 110 316 116 317
rect 1326 321 1332 322
rect 1326 317 1327 321
rect 1331 317 1332 321
rect 1606 318 1607 322
rect 1611 318 1612 322
rect 1606 317 1612 318
rect 1662 322 1668 323
rect 1662 318 1663 322
rect 1667 318 1668 322
rect 1662 317 1668 318
rect 1718 322 1724 323
rect 1718 318 1719 322
rect 1723 318 1724 322
rect 1718 317 1724 318
rect 1774 322 1780 323
rect 1774 318 1775 322
rect 1779 318 1780 322
rect 1774 317 1780 318
rect 1830 322 1836 323
rect 1830 318 1831 322
rect 1835 318 1836 322
rect 1830 317 1836 318
rect 1886 322 1892 323
rect 1886 318 1887 322
rect 1891 318 1892 322
rect 1886 317 1892 318
rect 1950 322 1956 323
rect 1950 318 1951 322
rect 1955 318 1956 322
rect 1950 317 1956 318
rect 2030 322 2036 323
rect 2030 318 2031 322
rect 2035 318 2036 322
rect 2030 317 2036 318
rect 2118 322 2124 323
rect 2118 318 2119 322
rect 2123 318 2124 322
rect 2118 317 2124 318
rect 2222 322 2228 323
rect 2222 318 2223 322
rect 2227 318 2228 322
rect 2222 317 2228 318
rect 2334 322 2340 323
rect 2334 318 2335 322
rect 2339 318 2340 322
rect 2334 317 2340 318
rect 2446 322 2452 323
rect 2446 318 2447 322
rect 2451 318 2452 322
rect 2446 317 2452 318
rect 2542 322 2548 323
rect 2542 318 2543 322
rect 2547 318 2548 322
rect 2542 317 2548 318
rect 1326 316 1332 317
rect 1366 313 1372 314
rect 1366 309 1367 313
rect 1371 309 1372 313
rect 1366 308 1372 309
rect 2582 313 2588 314
rect 2582 309 2583 313
rect 2587 309 2588 313
rect 2582 308 2588 309
rect 110 304 116 305
rect 1326 304 1332 305
rect 110 300 111 304
rect 115 300 116 304
rect 110 299 116 300
rect 142 303 148 304
rect 142 299 143 303
rect 147 299 148 303
rect 142 298 148 299
rect 206 303 212 304
rect 206 299 207 303
rect 211 299 212 303
rect 206 298 212 299
rect 294 303 300 304
rect 294 299 295 303
rect 299 299 300 303
rect 294 298 300 299
rect 374 303 380 304
rect 374 299 375 303
rect 379 299 380 303
rect 374 298 380 299
rect 454 303 460 304
rect 454 299 455 303
rect 459 299 460 303
rect 454 298 460 299
rect 526 303 532 304
rect 526 299 527 303
rect 531 299 532 303
rect 526 298 532 299
rect 590 303 596 304
rect 590 299 591 303
rect 595 299 596 303
rect 590 298 596 299
rect 654 303 660 304
rect 654 299 655 303
rect 659 299 660 303
rect 654 298 660 299
rect 718 303 724 304
rect 718 299 719 303
rect 723 299 724 303
rect 718 298 724 299
rect 782 303 788 304
rect 782 299 783 303
rect 787 299 788 303
rect 782 298 788 299
rect 846 303 852 304
rect 846 299 847 303
rect 851 299 852 303
rect 846 298 852 299
rect 918 303 924 304
rect 918 299 919 303
rect 923 299 924 303
rect 1326 300 1327 304
rect 1331 300 1332 304
rect 1326 299 1332 300
rect 918 298 924 299
rect 1366 296 1372 297
rect 2582 296 2588 297
rect 1366 292 1367 296
rect 1371 292 1372 296
rect 1366 291 1372 292
rect 1590 295 1596 296
rect 1590 291 1591 295
rect 1595 291 1596 295
rect 1590 290 1596 291
rect 1646 295 1652 296
rect 1646 291 1647 295
rect 1651 291 1652 295
rect 1646 290 1652 291
rect 1702 295 1708 296
rect 1702 291 1703 295
rect 1707 291 1708 295
rect 1702 290 1708 291
rect 1758 295 1764 296
rect 1758 291 1759 295
rect 1763 291 1764 295
rect 1758 290 1764 291
rect 1814 295 1820 296
rect 1814 291 1815 295
rect 1819 291 1820 295
rect 1814 290 1820 291
rect 1870 295 1876 296
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 1870 290 1876 291
rect 1934 295 1940 296
rect 1934 291 1935 295
rect 1939 291 1940 295
rect 1934 290 1940 291
rect 2014 295 2020 296
rect 2014 291 2015 295
rect 2019 291 2020 295
rect 2014 290 2020 291
rect 2102 295 2108 296
rect 2102 291 2103 295
rect 2107 291 2108 295
rect 2102 290 2108 291
rect 2206 295 2212 296
rect 2206 291 2207 295
rect 2211 291 2212 295
rect 2206 290 2212 291
rect 2318 295 2324 296
rect 2318 291 2319 295
rect 2323 291 2324 295
rect 2318 290 2324 291
rect 2430 295 2436 296
rect 2430 291 2431 295
rect 2435 291 2436 295
rect 2430 290 2436 291
rect 2526 295 2532 296
rect 2526 291 2527 295
rect 2531 291 2532 295
rect 2582 292 2583 296
rect 2587 292 2588 296
rect 2582 291 2588 292
rect 2526 290 2532 291
rect 142 261 148 262
rect 110 260 116 261
rect 110 256 111 260
rect 115 256 116 260
rect 142 257 143 261
rect 147 257 148 261
rect 142 256 148 257
rect 230 261 236 262
rect 230 257 231 261
rect 235 257 236 261
rect 230 256 236 257
rect 334 261 340 262
rect 334 257 335 261
rect 339 257 340 261
rect 334 256 340 257
rect 430 261 436 262
rect 430 257 431 261
rect 435 257 436 261
rect 430 256 436 257
rect 518 261 524 262
rect 518 257 519 261
rect 523 257 524 261
rect 518 256 524 257
rect 598 261 604 262
rect 598 257 599 261
rect 603 257 604 261
rect 598 256 604 257
rect 678 261 684 262
rect 678 257 679 261
rect 683 257 684 261
rect 678 256 684 257
rect 750 261 756 262
rect 750 257 751 261
rect 755 257 756 261
rect 750 256 756 257
rect 814 261 820 262
rect 814 257 815 261
rect 819 257 820 261
rect 814 256 820 257
rect 886 261 892 262
rect 886 257 887 261
rect 891 257 892 261
rect 886 256 892 257
rect 958 261 964 262
rect 958 257 959 261
rect 963 257 964 261
rect 958 256 964 257
rect 1030 261 1036 262
rect 1030 257 1031 261
rect 1035 257 1036 261
rect 1030 256 1036 257
rect 1326 260 1332 261
rect 1326 256 1327 260
rect 1331 256 1332 260
rect 1726 257 1732 258
rect 110 255 116 256
rect 1326 255 1332 256
rect 1366 256 1372 257
rect 1366 252 1367 256
rect 1371 252 1372 256
rect 1726 253 1727 257
rect 1731 253 1732 257
rect 1726 252 1732 253
rect 1782 257 1788 258
rect 1782 253 1783 257
rect 1787 253 1788 257
rect 1782 252 1788 253
rect 1838 257 1844 258
rect 1838 253 1839 257
rect 1843 253 1844 257
rect 1838 252 1844 253
rect 1894 257 1900 258
rect 1894 253 1895 257
rect 1899 253 1900 257
rect 1894 252 1900 253
rect 1950 257 1956 258
rect 1950 253 1951 257
rect 1955 253 1956 257
rect 1950 252 1956 253
rect 2006 257 2012 258
rect 2006 253 2007 257
rect 2011 253 2012 257
rect 2006 252 2012 253
rect 2070 257 2076 258
rect 2070 253 2071 257
rect 2075 253 2076 257
rect 2070 252 2076 253
rect 2142 257 2148 258
rect 2142 253 2143 257
rect 2147 253 2148 257
rect 2142 252 2148 253
rect 2230 257 2236 258
rect 2230 253 2231 257
rect 2235 253 2236 257
rect 2230 252 2236 253
rect 2334 257 2340 258
rect 2334 253 2335 257
rect 2339 253 2340 257
rect 2334 252 2340 253
rect 2438 257 2444 258
rect 2438 253 2439 257
rect 2443 253 2444 257
rect 2438 252 2444 253
rect 2526 257 2532 258
rect 2526 253 2527 257
rect 2531 253 2532 257
rect 2526 252 2532 253
rect 2582 256 2588 257
rect 2582 252 2583 256
rect 2587 252 2588 256
rect 1366 251 1372 252
rect 2582 251 2588 252
rect 110 243 116 244
rect 110 239 111 243
rect 115 239 116 243
rect 110 238 116 239
rect 1326 243 1332 244
rect 1326 239 1327 243
rect 1331 239 1332 243
rect 1326 238 1332 239
rect 1366 239 1372 240
rect 1366 235 1367 239
rect 1371 235 1372 239
rect 158 234 164 235
rect 158 230 159 234
rect 163 230 164 234
rect 158 229 164 230
rect 246 234 252 235
rect 246 230 247 234
rect 251 230 252 234
rect 246 229 252 230
rect 350 234 356 235
rect 350 230 351 234
rect 355 230 356 234
rect 350 229 356 230
rect 446 234 452 235
rect 446 230 447 234
rect 451 230 452 234
rect 446 229 452 230
rect 534 234 540 235
rect 534 230 535 234
rect 539 230 540 234
rect 534 229 540 230
rect 614 234 620 235
rect 614 230 615 234
rect 619 230 620 234
rect 614 229 620 230
rect 694 234 700 235
rect 694 230 695 234
rect 699 230 700 234
rect 694 229 700 230
rect 766 234 772 235
rect 766 230 767 234
rect 771 230 772 234
rect 766 229 772 230
rect 830 234 836 235
rect 830 230 831 234
rect 835 230 836 234
rect 830 229 836 230
rect 902 234 908 235
rect 902 230 903 234
rect 907 230 908 234
rect 902 229 908 230
rect 974 234 980 235
rect 974 230 975 234
rect 979 230 980 234
rect 974 229 980 230
rect 1046 234 1052 235
rect 1366 234 1372 235
rect 2582 239 2588 240
rect 2582 235 2583 239
rect 2587 235 2588 239
rect 2582 234 2588 235
rect 1046 230 1047 234
rect 1051 230 1052 234
rect 1046 229 1052 230
rect 1742 230 1748 231
rect 1742 226 1743 230
rect 1747 226 1748 230
rect 1742 225 1748 226
rect 1798 230 1804 231
rect 1798 226 1799 230
rect 1803 226 1804 230
rect 1798 225 1804 226
rect 1854 230 1860 231
rect 1854 226 1855 230
rect 1859 226 1860 230
rect 1854 225 1860 226
rect 1910 230 1916 231
rect 1910 226 1911 230
rect 1915 226 1916 230
rect 1910 225 1916 226
rect 1966 230 1972 231
rect 1966 226 1967 230
rect 1971 226 1972 230
rect 1966 225 1972 226
rect 2022 230 2028 231
rect 2022 226 2023 230
rect 2027 226 2028 230
rect 2022 225 2028 226
rect 2086 230 2092 231
rect 2086 226 2087 230
rect 2091 226 2092 230
rect 2086 225 2092 226
rect 2158 230 2164 231
rect 2158 226 2159 230
rect 2163 226 2164 230
rect 2158 225 2164 226
rect 2246 230 2252 231
rect 2246 226 2247 230
rect 2251 226 2252 230
rect 2246 225 2252 226
rect 2350 230 2356 231
rect 2350 226 2351 230
rect 2355 226 2356 230
rect 2350 225 2356 226
rect 2454 230 2460 231
rect 2454 226 2455 230
rect 2459 226 2460 230
rect 2454 225 2460 226
rect 2542 230 2548 231
rect 2542 226 2543 230
rect 2547 226 2548 230
rect 2542 225 2548 226
rect 166 206 172 207
rect 166 202 167 206
rect 171 202 172 206
rect 166 201 172 202
rect 254 206 260 207
rect 254 202 255 206
rect 259 202 260 206
rect 254 201 260 202
rect 350 206 356 207
rect 350 202 351 206
rect 355 202 356 206
rect 350 201 356 202
rect 446 206 452 207
rect 446 202 447 206
rect 451 202 452 206
rect 446 201 452 202
rect 550 206 556 207
rect 550 202 551 206
rect 555 202 556 206
rect 550 201 556 202
rect 654 206 660 207
rect 654 202 655 206
rect 659 202 660 206
rect 654 201 660 202
rect 750 206 756 207
rect 750 202 751 206
rect 755 202 756 206
rect 750 201 756 202
rect 846 206 852 207
rect 846 202 847 206
rect 851 202 852 206
rect 846 201 852 202
rect 934 206 940 207
rect 934 202 935 206
rect 939 202 940 206
rect 934 201 940 202
rect 1022 206 1028 207
rect 1022 202 1023 206
rect 1027 202 1028 206
rect 1022 201 1028 202
rect 1110 206 1116 207
rect 1110 202 1111 206
rect 1115 202 1116 206
rect 1110 201 1116 202
rect 1198 206 1204 207
rect 1198 202 1199 206
rect 1203 202 1204 206
rect 1198 201 1204 202
rect 1462 206 1468 207
rect 1462 202 1463 206
rect 1467 202 1468 206
rect 1462 201 1468 202
rect 1534 206 1540 207
rect 1534 202 1535 206
rect 1539 202 1540 206
rect 1534 201 1540 202
rect 1622 206 1628 207
rect 1622 202 1623 206
rect 1627 202 1628 206
rect 1622 201 1628 202
rect 1718 206 1724 207
rect 1718 202 1719 206
rect 1723 202 1724 206
rect 1718 201 1724 202
rect 1822 206 1828 207
rect 1822 202 1823 206
rect 1827 202 1828 206
rect 1822 201 1828 202
rect 1926 206 1932 207
rect 1926 202 1927 206
rect 1931 202 1932 206
rect 1926 201 1932 202
rect 2030 206 2036 207
rect 2030 202 2031 206
rect 2035 202 2036 206
rect 2030 201 2036 202
rect 2134 206 2140 207
rect 2134 202 2135 206
rect 2139 202 2140 206
rect 2134 201 2140 202
rect 2238 206 2244 207
rect 2238 202 2239 206
rect 2243 202 2244 206
rect 2238 201 2244 202
rect 2342 206 2348 207
rect 2342 202 2343 206
rect 2347 202 2348 206
rect 2342 201 2348 202
rect 2454 206 2460 207
rect 2454 202 2455 206
rect 2459 202 2460 206
rect 2454 201 2460 202
rect 2542 206 2548 207
rect 2542 202 2543 206
rect 2547 202 2548 206
rect 2542 201 2548 202
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 110 192 116 193
rect 1326 197 1332 198
rect 1326 193 1327 197
rect 1331 193 1332 197
rect 1326 192 1332 193
rect 1366 197 1372 198
rect 1366 193 1367 197
rect 1371 193 1372 197
rect 1366 192 1372 193
rect 2582 197 2588 198
rect 2582 193 2583 197
rect 2587 193 2588 197
rect 2582 192 2588 193
rect 110 180 116 181
rect 1326 180 1332 181
rect 110 176 111 180
rect 115 176 116 180
rect 110 175 116 176
rect 150 179 156 180
rect 150 175 151 179
rect 155 175 156 179
rect 150 174 156 175
rect 238 179 244 180
rect 238 175 239 179
rect 243 175 244 179
rect 238 174 244 175
rect 334 179 340 180
rect 334 175 335 179
rect 339 175 340 179
rect 334 174 340 175
rect 430 179 436 180
rect 430 175 431 179
rect 435 175 436 179
rect 430 174 436 175
rect 534 179 540 180
rect 534 175 535 179
rect 539 175 540 179
rect 534 174 540 175
rect 638 179 644 180
rect 638 175 639 179
rect 643 175 644 179
rect 638 174 644 175
rect 734 179 740 180
rect 734 175 735 179
rect 739 175 740 179
rect 734 174 740 175
rect 830 179 836 180
rect 830 175 831 179
rect 835 175 836 179
rect 830 174 836 175
rect 918 179 924 180
rect 918 175 919 179
rect 923 175 924 179
rect 918 174 924 175
rect 1006 179 1012 180
rect 1006 175 1007 179
rect 1011 175 1012 179
rect 1006 174 1012 175
rect 1094 179 1100 180
rect 1094 175 1095 179
rect 1099 175 1100 179
rect 1094 174 1100 175
rect 1182 179 1188 180
rect 1182 175 1183 179
rect 1187 175 1188 179
rect 1326 176 1327 180
rect 1331 176 1332 180
rect 1326 175 1332 176
rect 1366 180 1372 181
rect 2582 180 2588 181
rect 1366 176 1367 180
rect 1371 176 1372 180
rect 1366 175 1372 176
rect 1446 179 1452 180
rect 1446 175 1447 179
rect 1451 175 1452 179
rect 1182 174 1188 175
rect 1446 174 1452 175
rect 1518 179 1524 180
rect 1518 175 1519 179
rect 1523 175 1524 179
rect 1518 174 1524 175
rect 1606 179 1612 180
rect 1606 175 1607 179
rect 1611 175 1612 179
rect 1606 174 1612 175
rect 1702 179 1708 180
rect 1702 175 1703 179
rect 1707 175 1708 179
rect 1702 174 1708 175
rect 1806 179 1812 180
rect 1806 175 1807 179
rect 1811 175 1812 179
rect 1806 174 1812 175
rect 1910 179 1916 180
rect 1910 175 1911 179
rect 1915 175 1916 179
rect 1910 174 1916 175
rect 2014 179 2020 180
rect 2014 175 2015 179
rect 2019 175 2020 179
rect 2014 174 2020 175
rect 2118 179 2124 180
rect 2118 175 2119 179
rect 2123 175 2124 179
rect 2118 174 2124 175
rect 2222 179 2228 180
rect 2222 175 2223 179
rect 2227 175 2228 179
rect 2222 174 2228 175
rect 2326 179 2332 180
rect 2326 175 2327 179
rect 2331 175 2332 179
rect 2326 174 2332 175
rect 2438 179 2444 180
rect 2438 175 2439 179
rect 2443 175 2444 179
rect 2438 174 2444 175
rect 2526 179 2532 180
rect 2526 175 2527 179
rect 2531 175 2532 179
rect 2582 176 2583 180
rect 2587 176 2588 180
rect 2582 175 2588 176
rect 2526 174 2532 175
rect 1398 129 1404 130
rect 1366 128 1372 129
rect 1366 124 1367 128
rect 1371 124 1372 128
rect 1398 125 1399 129
rect 1403 125 1404 129
rect 1398 124 1404 125
rect 1454 129 1460 130
rect 1454 125 1455 129
rect 1459 125 1460 129
rect 1454 124 1460 125
rect 1510 129 1516 130
rect 1510 125 1511 129
rect 1515 125 1516 129
rect 1510 124 1516 125
rect 1566 129 1572 130
rect 1566 125 1567 129
rect 1571 125 1572 129
rect 1566 124 1572 125
rect 1638 129 1644 130
rect 1638 125 1639 129
rect 1643 125 1644 129
rect 1638 124 1644 125
rect 1718 129 1724 130
rect 1718 125 1719 129
rect 1723 125 1724 129
rect 1718 124 1724 125
rect 1798 129 1804 130
rect 1798 125 1799 129
rect 1803 125 1804 129
rect 1798 124 1804 125
rect 1878 129 1884 130
rect 1878 125 1879 129
rect 1883 125 1884 129
rect 1878 124 1884 125
rect 1958 129 1964 130
rect 1958 125 1959 129
rect 1963 125 1964 129
rect 1958 124 1964 125
rect 2030 129 2036 130
rect 2030 125 2031 129
rect 2035 125 2036 129
rect 2030 124 2036 125
rect 2102 129 2108 130
rect 2102 125 2103 129
rect 2107 125 2108 129
rect 2102 124 2108 125
rect 2166 129 2172 130
rect 2166 125 2167 129
rect 2171 125 2172 129
rect 2166 124 2172 125
rect 2230 129 2236 130
rect 2230 125 2231 129
rect 2235 125 2236 129
rect 2230 124 2236 125
rect 2294 129 2300 130
rect 2294 125 2295 129
rect 2299 125 2300 129
rect 2294 124 2300 125
rect 2358 129 2364 130
rect 2358 125 2359 129
rect 2363 125 2364 129
rect 2358 124 2364 125
rect 2414 129 2420 130
rect 2414 125 2415 129
rect 2419 125 2420 129
rect 2414 124 2420 125
rect 2470 129 2476 130
rect 2470 125 2471 129
rect 2475 125 2476 129
rect 2470 124 2476 125
rect 2526 129 2532 130
rect 2526 125 2527 129
rect 2531 125 2532 129
rect 2526 124 2532 125
rect 2582 128 2588 129
rect 2582 124 2583 128
rect 2587 124 2588 128
rect 1366 123 1372 124
rect 2582 123 2588 124
rect 142 121 148 122
rect 110 120 116 121
rect 110 116 111 120
rect 115 116 116 120
rect 142 117 143 121
rect 147 117 148 121
rect 142 116 148 117
rect 198 121 204 122
rect 198 117 199 121
rect 203 117 204 121
rect 198 116 204 117
rect 254 121 260 122
rect 254 117 255 121
rect 259 117 260 121
rect 254 116 260 117
rect 310 121 316 122
rect 310 117 311 121
rect 315 117 316 121
rect 310 116 316 117
rect 366 121 372 122
rect 366 117 367 121
rect 371 117 372 121
rect 366 116 372 117
rect 422 121 428 122
rect 422 117 423 121
rect 427 117 428 121
rect 422 116 428 117
rect 478 121 484 122
rect 478 117 479 121
rect 483 117 484 121
rect 478 116 484 117
rect 534 121 540 122
rect 534 117 535 121
rect 539 117 540 121
rect 534 116 540 117
rect 606 121 612 122
rect 606 117 607 121
rect 611 117 612 121
rect 606 116 612 117
rect 670 121 676 122
rect 670 117 671 121
rect 675 117 676 121
rect 670 116 676 117
rect 734 121 740 122
rect 734 117 735 121
rect 739 117 740 121
rect 734 116 740 117
rect 798 121 804 122
rect 798 117 799 121
rect 803 117 804 121
rect 798 116 804 117
rect 854 121 860 122
rect 854 117 855 121
rect 859 117 860 121
rect 854 116 860 117
rect 910 121 916 122
rect 910 117 911 121
rect 915 117 916 121
rect 910 116 916 117
rect 974 121 980 122
rect 974 117 975 121
rect 979 117 980 121
rect 974 116 980 117
rect 1038 121 1044 122
rect 1038 117 1039 121
rect 1043 117 1044 121
rect 1038 116 1044 117
rect 1102 121 1108 122
rect 1102 117 1103 121
rect 1107 117 1108 121
rect 1102 116 1108 117
rect 1158 121 1164 122
rect 1158 117 1159 121
rect 1163 117 1164 121
rect 1158 116 1164 117
rect 1214 121 1220 122
rect 1214 117 1215 121
rect 1219 117 1220 121
rect 1214 116 1220 117
rect 1270 121 1276 122
rect 1270 117 1271 121
rect 1275 117 1276 121
rect 1270 116 1276 117
rect 1326 120 1332 121
rect 1326 116 1327 120
rect 1331 116 1332 120
rect 110 115 116 116
rect 1326 115 1332 116
rect 1366 111 1372 112
rect 1366 107 1367 111
rect 1371 107 1372 111
rect 1366 106 1372 107
rect 2582 111 2588 112
rect 2582 107 2583 111
rect 2587 107 2588 111
rect 2582 106 2588 107
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 110 98 116 99
rect 1326 103 1332 104
rect 1326 99 1327 103
rect 1331 99 1332 103
rect 1326 98 1332 99
rect 1414 102 1420 103
rect 1414 98 1415 102
rect 1419 98 1420 102
rect 1414 97 1420 98
rect 1470 102 1476 103
rect 1470 98 1471 102
rect 1475 98 1476 102
rect 1470 97 1476 98
rect 1526 102 1532 103
rect 1526 98 1527 102
rect 1531 98 1532 102
rect 1526 97 1532 98
rect 1582 102 1588 103
rect 1582 98 1583 102
rect 1587 98 1588 102
rect 1582 97 1588 98
rect 1654 102 1660 103
rect 1654 98 1655 102
rect 1659 98 1660 102
rect 1654 97 1660 98
rect 1734 102 1740 103
rect 1734 98 1735 102
rect 1739 98 1740 102
rect 1734 97 1740 98
rect 1814 102 1820 103
rect 1814 98 1815 102
rect 1819 98 1820 102
rect 1814 97 1820 98
rect 1894 102 1900 103
rect 1894 98 1895 102
rect 1899 98 1900 102
rect 1894 97 1900 98
rect 1974 102 1980 103
rect 1974 98 1975 102
rect 1979 98 1980 102
rect 1974 97 1980 98
rect 2046 102 2052 103
rect 2046 98 2047 102
rect 2051 98 2052 102
rect 2046 97 2052 98
rect 2118 102 2124 103
rect 2118 98 2119 102
rect 2123 98 2124 102
rect 2118 97 2124 98
rect 2182 102 2188 103
rect 2182 98 2183 102
rect 2187 98 2188 102
rect 2182 97 2188 98
rect 2246 102 2252 103
rect 2246 98 2247 102
rect 2251 98 2252 102
rect 2246 97 2252 98
rect 2310 102 2316 103
rect 2310 98 2311 102
rect 2315 98 2316 102
rect 2310 97 2316 98
rect 2374 102 2380 103
rect 2374 98 2375 102
rect 2379 98 2380 102
rect 2374 97 2380 98
rect 2430 102 2436 103
rect 2430 98 2431 102
rect 2435 98 2436 102
rect 2430 97 2436 98
rect 2486 102 2492 103
rect 2486 98 2487 102
rect 2491 98 2492 102
rect 2486 97 2492 98
rect 2542 102 2548 103
rect 2542 98 2543 102
rect 2547 98 2548 102
rect 2542 97 2548 98
rect 158 94 164 95
rect 158 90 159 94
rect 163 90 164 94
rect 158 89 164 90
rect 214 94 220 95
rect 214 90 215 94
rect 219 90 220 94
rect 214 89 220 90
rect 270 94 276 95
rect 270 90 271 94
rect 275 90 276 94
rect 270 89 276 90
rect 326 94 332 95
rect 326 90 327 94
rect 331 90 332 94
rect 326 89 332 90
rect 382 94 388 95
rect 382 90 383 94
rect 387 90 388 94
rect 382 89 388 90
rect 438 94 444 95
rect 438 90 439 94
rect 443 90 444 94
rect 438 89 444 90
rect 494 94 500 95
rect 494 90 495 94
rect 499 90 500 94
rect 494 89 500 90
rect 550 94 556 95
rect 550 90 551 94
rect 555 90 556 94
rect 550 89 556 90
rect 622 94 628 95
rect 622 90 623 94
rect 627 90 628 94
rect 622 89 628 90
rect 686 94 692 95
rect 686 90 687 94
rect 691 90 692 94
rect 686 89 692 90
rect 750 94 756 95
rect 750 90 751 94
rect 755 90 756 94
rect 750 89 756 90
rect 814 94 820 95
rect 814 90 815 94
rect 819 90 820 94
rect 814 89 820 90
rect 870 94 876 95
rect 870 90 871 94
rect 875 90 876 94
rect 870 89 876 90
rect 926 94 932 95
rect 926 90 927 94
rect 931 90 932 94
rect 926 89 932 90
rect 990 94 996 95
rect 990 90 991 94
rect 995 90 996 94
rect 990 89 996 90
rect 1054 94 1060 95
rect 1054 90 1055 94
rect 1059 90 1060 94
rect 1054 89 1060 90
rect 1118 94 1124 95
rect 1118 90 1119 94
rect 1123 90 1124 94
rect 1118 89 1124 90
rect 1174 94 1180 95
rect 1174 90 1175 94
rect 1179 90 1180 94
rect 1174 89 1180 90
rect 1230 94 1236 95
rect 1230 90 1231 94
rect 1235 90 1236 94
rect 1230 89 1236 90
rect 1286 94 1292 95
rect 1286 90 1287 94
rect 1291 90 1292 94
rect 1286 89 1292 90
<< m3c >>
rect 159 2646 163 2650
rect 215 2646 219 2650
rect 271 2646 275 2650
rect 327 2646 331 2650
rect 111 2637 115 2641
rect 1327 2637 1331 2641
rect 111 2620 115 2624
rect 143 2619 147 2623
rect 199 2619 203 2623
rect 255 2619 259 2623
rect 311 2619 315 2623
rect 1327 2620 1331 2624
rect 1415 2594 1419 2598
rect 1471 2594 1475 2598
rect 1527 2594 1531 2598
rect 1583 2594 1587 2598
rect 1639 2594 1643 2598
rect 1695 2594 1699 2598
rect 111 2584 115 2588
rect 143 2585 147 2589
rect 199 2585 203 2589
rect 263 2585 267 2589
rect 343 2585 347 2589
rect 431 2585 435 2589
rect 519 2585 523 2589
rect 607 2585 611 2589
rect 687 2585 691 2589
rect 767 2585 771 2589
rect 839 2585 843 2589
rect 903 2585 907 2589
rect 967 2585 971 2589
rect 1031 2585 1035 2589
rect 1095 2585 1099 2589
rect 1159 2585 1163 2589
rect 1215 2585 1219 2589
rect 1271 2585 1275 2589
rect 1327 2584 1331 2588
rect 1367 2585 1371 2589
rect 2583 2585 2587 2589
rect 111 2567 115 2571
rect 1327 2567 1331 2571
rect 1367 2568 1371 2572
rect 1399 2567 1403 2571
rect 1455 2567 1459 2571
rect 1511 2567 1515 2571
rect 1567 2567 1571 2571
rect 1623 2567 1627 2571
rect 1679 2567 1683 2571
rect 2583 2568 2587 2572
rect 159 2558 163 2562
rect 215 2558 219 2562
rect 279 2558 283 2562
rect 359 2558 363 2562
rect 447 2558 451 2562
rect 535 2558 539 2562
rect 623 2558 627 2562
rect 703 2558 707 2562
rect 783 2558 787 2562
rect 855 2558 859 2562
rect 919 2558 923 2562
rect 983 2558 987 2562
rect 1047 2558 1051 2562
rect 1111 2558 1115 2562
rect 1175 2558 1179 2562
rect 1231 2558 1235 2562
rect 1287 2558 1291 2562
rect 1367 2532 1371 2536
rect 1399 2533 1403 2537
rect 1455 2533 1459 2537
rect 1511 2533 1515 2537
rect 1567 2533 1571 2537
rect 1623 2533 1627 2537
rect 1679 2533 1683 2537
rect 1735 2533 1739 2537
rect 2583 2532 2587 2536
rect 159 2522 163 2526
rect 215 2522 219 2526
rect 319 2522 323 2526
rect 431 2522 435 2526
rect 551 2522 555 2526
rect 671 2522 675 2526
rect 791 2522 795 2526
rect 903 2522 907 2526
rect 1007 2522 1011 2526
rect 1103 2522 1107 2526
rect 1207 2522 1211 2526
rect 1287 2522 1291 2526
rect 111 2513 115 2517
rect 1327 2513 1331 2517
rect 1367 2515 1371 2519
rect 2583 2515 2587 2519
rect 1415 2506 1419 2510
rect 1471 2506 1475 2510
rect 1527 2506 1531 2510
rect 1583 2506 1587 2510
rect 1639 2506 1643 2510
rect 1695 2506 1699 2510
rect 1751 2506 1755 2510
rect 111 2496 115 2500
rect 143 2495 147 2499
rect 199 2495 203 2499
rect 303 2495 307 2499
rect 415 2495 419 2499
rect 535 2495 539 2499
rect 655 2495 659 2499
rect 775 2495 779 2499
rect 887 2495 891 2499
rect 991 2495 995 2499
rect 1087 2495 1091 2499
rect 1191 2495 1195 2499
rect 1271 2495 1275 2499
rect 1327 2496 1331 2500
rect 1471 2478 1475 2482
rect 1527 2478 1531 2482
rect 1583 2478 1587 2482
rect 1639 2478 1643 2482
rect 1695 2478 1699 2482
rect 1751 2478 1755 2482
rect 1367 2469 1371 2473
rect 2583 2469 2587 2473
rect 111 2452 115 2456
rect 143 2453 147 2457
rect 199 2453 203 2457
rect 295 2453 299 2457
rect 407 2453 411 2457
rect 519 2453 523 2457
rect 639 2453 643 2457
rect 751 2453 755 2457
rect 855 2453 859 2457
rect 951 2453 955 2457
rect 1047 2453 1051 2457
rect 1143 2453 1147 2457
rect 1239 2453 1243 2457
rect 1327 2452 1331 2456
rect 1367 2452 1371 2456
rect 1455 2451 1459 2455
rect 1511 2451 1515 2455
rect 1567 2451 1571 2455
rect 1623 2451 1627 2455
rect 1679 2451 1683 2455
rect 1735 2451 1739 2455
rect 2583 2452 2587 2456
rect 111 2435 115 2439
rect 1327 2435 1331 2439
rect 159 2426 163 2430
rect 215 2426 219 2430
rect 311 2426 315 2430
rect 423 2426 427 2430
rect 535 2426 539 2430
rect 655 2426 659 2430
rect 767 2426 771 2430
rect 871 2426 875 2430
rect 967 2426 971 2430
rect 1063 2426 1067 2430
rect 1159 2426 1163 2430
rect 1255 2426 1259 2430
rect 1367 2408 1371 2412
rect 1479 2409 1483 2413
rect 1535 2409 1539 2413
rect 1591 2409 1595 2413
rect 1647 2409 1651 2413
rect 1703 2409 1707 2413
rect 1759 2409 1763 2413
rect 2583 2408 2587 2412
rect 223 2394 227 2398
rect 287 2394 291 2398
rect 367 2394 371 2398
rect 455 2394 459 2398
rect 543 2394 547 2398
rect 639 2394 643 2398
rect 727 2394 731 2398
rect 815 2394 819 2398
rect 895 2394 899 2398
rect 975 2394 979 2398
rect 1055 2394 1059 2398
rect 1143 2394 1147 2398
rect 1367 2391 1371 2395
rect 2583 2391 2587 2395
rect 111 2385 115 2389
rect 1327 2385 1331 2389
rect 1495 2382 1499 2386
rect 1551 2382 1555 2386
rect 1607 2382 1611 2386
rect 1663 2382 1667 2386
rect 1719 2382 1723 2386
rect 1775 2382 1779 2386
rect 111 2368 115 2372
rect 207 2367 211 2371
rect 271 2367 275 2371
rect 351 2367 355 2371
rect 439 2367 443 2371
rect 527 2367 531 2371
rect 623 2367 627 2371
rect 711 2367 715 2371
rect 799 2367 803 2371
rect 879 2367 883 2371
rect 959 2367 963 2371
rect 1039 2367 1043 2371
rect 1127 2367 1131 2371
rect 1327 2368 1331 2372
rect 1471 2354 1475 2358
rect 1527 2354 1531 2358
rect 1583 2354 1587 2358
rect 1639 2354 1643 2358
rect 1695 2354 1699 2358
rect 1367 2345 1371 2349
rect 2583 2345 2587 2349
rect 111 2324 115 2328
rect 327 2325 331 2329
rect 383 2325 387 2329
rect 439 2325 443 2329
rect 503 2325 507 2329
rect 567 2325 571 2329
rect 631 2325 635 2329
rect 695 2325 699 2329
rect 759 2325 763 2329
rect 823 2325 827 2329
rect 887 2325 891 2329
rect 951 2325 955 2329
rect 1015 2325 1019 2329
rect 1327 2324 1331 2328
rect 1367 2328 1371 2332
rect 1455 2327 1459 2331
rect 1511 2327 1515 2331
rect 1567 2327 1571 2331
rect 1623 2327 1627 2331
rect 1679 2327 1683 2331
rect 2583 2328 2587 2332
rect 111 2307 115 2311
rect 1327 2307 1331 2311
rect 343 2298 347 2302
rect 399 2298 403 2302
rect 455 2298 459 2302
rect 519 2298 523 2302
rect 583 2298 587 2302
rect 647 2298 651 2302
rect 711 2298 715 2302
rect 775 2298 779 2302
rect 839 2298 843 2302
rect 903 2298 907 2302
rect 967 2298 971 2302
rect 1031 2298 1035 2302
rect 1367 2292 1371 2296
rect 1399 2293 1403 2297
rect 1455 2293 1459 2297
rect 1511 2293 1515 2297
rect 1567 2293 1571 2297
rect 1623 2293 1627 2297
rect 1679 2293 1683 2297
rect 1735 2293 1739 2297
rect 1791 2293 1795 2297
rect 1847 2293 1851 2297
rect 1903 2293 1907 2297
rect 1959 2293 1963 2297
rect 2015 2293 2019 2297
rect 2071 2293 2075 2297
rect 2127 2293 2131 2297
rect 2183 2293 2187 2297
rect 2247 2293 2251 2297
rect 2311 2293 2315 2297
rect 2375 2293 2379 2297
rect 2439 2293 2443 2297
rect 2583 2292 2587 2296
rect 1367 2275 1371 2279
rect 2583 2275 2587 2279
rect 407 2266 411 2270
rect 463 2266 467 2270
rect 519 2266 523 2270
rect 575 2266 579 2270
rect 631 2266 635 2270
rect 687 2266 691 2270
rect 743 2266 747 2270
rect 799 2266 803 2270
rect 855 2266 859 2270
rect 911 2266 915 2270
rect 967 2266 971 2270
rect 1415 2266 1419 2270
rect 1471 2266 1475 2270
rect 1527 2266 1531 2270
rect 1583 2266 1587 2270
rect 1639 2266 1643 2270
rect 1695 2266 1699 2270
rect 1751 2266 1755 2270
rect 1807 2266 1811 2270
rect 1863 2266 1867 2270
rect 1919 2266 1923 2270
rect 1975 2266 1979 2270
rect 2031 2266 2035 2270
rect 2087 2266 2091 2270
rect 2143 2266 2147 2270
rect 2199 2266 2203 2270
rect 2263 2266 2267 2270
rect 2327 2266 2331 2270
rect 2391 2266 2395 2270
rect 2455 2266 2459 2270
rect 111 2257 115 2261
rect 1327 2257 1331 2261
rect 111 2240 115 2244
rect 391 2239 395 2243
rect 447 2239 451 2243
rect 503 2239 507 2243
rect 559 2239 563 2243
rect 615 2239 619 2243
rect 671 2239 675 2243
rect 727 2239 731 2243
rect 783 2239 787 2243
rect 839 2239 843 2243
rect 895 2239 899 2243
rect 951 2239 955 2243
rect 1327 2240 1331 2244
rect 1415 2242 1419 2246
rect 1511 2242 1515 2246
rect 1623 2242 1627 2246
rect 1727 2242 1731 2246
rect 1823 2242 1827 2246
rect 1903 2242 1907 2246
rect 1983 2242 1987 2246
rect 2055 2242 2059 2246
rect 2119 2242 2123 2246
rect 2191 2242 2195 2246
rect 2263 2242 2267 2246
rect 2335 2242 2339 2246
rect 1367 2233 1371 2237
rect 2583 2233 2587 2237
rect 1367 2216 1371 2220
rect 1399 2215 1403 2219
rect 1495 2215 1499 2219
rect 1607 2215 1611 2219
rect 1711 2215 1715 2219
rect 1807 2215 1811 2219
rect 1887 2215 1891 2219
rect 1967 2215 1971 2219
rect 2039 2215 2043 2219
rect 2103 2215 2107 2219
rect 2175 2215 2179 2219
rect 2247 2215 2251 2219
rect 2319 2215 2323 2219
rect 2583 2216 2587 2220
rect 111 2200 115 2204
rect 423 2201 427 2205
rect 479 2201 483 2205
rect 535 2201 539 2205
rect 591 2201 595 2205
rect 647 2201 651 2205
rect 711 2201 715 2205
rect 783 2201 787 2205
rect 855 2201 859 2205
rect 927 2201 931 2205
rect 999 2201 1003 2205
rect 1071 2201 1075 2205
rect 1143 2201 1147 2205
rect 1215 2201 1219 2205
rect 1271 2201 1275 2205
rect 1327 2200 1331 2204
rect 111 2183 115 2187
rect 1327 2183 1331 2187
rect 439 2174 443 2178
rect 495 2174 499 2178
rect 551 2174 555 2178
rect 607 2174 611 2178
rect 663 2174 667 2178
rect 727 2174 731 2178
rect 799 2174 803 2178
rect 871 2174 875 2178
rect 943 2174 947 2178
rect 1015 2174 1019 2178
rect 1087 2174 1091 2178
rect 1159 2174 1163 2178
rect 1231 2174 1235 2178
rect 1287 2174 1291 2178
rect 1367 2176 1371 2180
rect 1751 2177 1755 2181
rect 1839 2177 1843 2181
rect 1927 2177 1931 2181
rect 2007 2177 2011 2181
rect 2087 2177 2091 2181
rect 2167 2177 2171 2181
rect 2247 2177 2251 2181
rect 2335 2177 2339 2181
rect 2423 2177 2427 2181
rect 2583 2176 2587 2180
rect 1367 2159 1371 2163
rect 2583 2159 2587 2163
rect 1767 2150 1771 2154
rect 1855 2150 1859 2154
rect 1943 2150 1947 2154
rect 2023 2150 2027 2154
rect 2103 2150 2107 2154
rect 2183 2150 2187 2154
rect 2263 2150 2267 2154
rect 2351 2150 2355 2154
rect 2439 2150 2443 2154
rect 199 2142 203 2146
rect 271 2142 275 2146
rect 351 2142 355 2146
rect 447 2142 451 2146
rect 551 2142 555 2146
rect 663 2142 667 2146
rect 775 2142 779 2146
rect 879 2142 883 2146
rect 983 2142 987 2146
rect 1079 2142 1083 2146
rect 1183 2142 1187 2146
rect 1287 2142 1291 2146
rect 111 2133 115 2137
rect 1327 2133 1331 2137
rect 1607 2126 1611 2130
rect 1679 2126 1683 2130
rect 1767 2126 1771 2130
rect 1863 2126 1867 2130
rect 1959 2126 1963 2130
rect 2063 2126 2067 2130
rect 2159 2126 2163 2130
rect 2255 2126 2259 2130
rect 2351 2126 2355 2130
rect 2447 2126 2451 2130
rect 2543 2126 2547 2130
rect 111 2116 115 2120
rect 183 2115 187 2119
rect 255 2115 259 2119
rect 335 2115 339 2119
rect 431 2115 435 2119
rect 535 2115 539 2119
rect 647 2115 651 2119
rect 759 2115 763 2119
rect 863 2115 867 2119
rect 967 2115 971 2119
rect 1063 2115 1067 2119
rect 1167 2115 1171 2119
rect 1271 2115 1275 2119
rect 1327 2116 1331 2120
rect 1367 2117 1371 2121
rect 2583 2117 2587 2121
rect 1367 2100 1371 2104
rect 1591 2099 1595 2103
rect 1663 2099 1667 2103
rect 1751 2099 1755 2103
rect 1847 2099 1851 2103
rect 1943 2099 1947 2103
rect 2047 2099 2051 2103
rect 2143 2099 2147 2103
rect 2239 2099 2243 2103
rect 2335 2099 2339 2103
rect 2431 2099 2435 2103
rect 2527 2099 2531 2103
rect 2583 2100 2587 2104
rect 111 2068 115 2072
rect 143 2069 147 2073
rect 199 2069 203 2073
rect 271 2069 275 2073
rect 367 2069 371 2073
rect 463 2069 467 2073
rect 567 2069 571 2073
rect 663 2069 667 2073
rect 759 2069 763 2073
rect 847 2069 851 2073
rect 927 2069 931 2073
rect 1007 2069 1011 2073
rect 1095 2069 1099 2073
rect 1183 2069 1187 2073
rect 1327 2068 1331 2072
rect 1367 2064 1371 2068
rect 1487 2065 1491 2069
rect 1583 2065 1587 2069
rect 1679 2065 1683 2069
rect 1783 2065 1787 2069
rect 1887 2065 1891 2069
rect 1983 2065 1987 2069
rect 2079 2065 2083 2069
rect 2167 2065 2171 2069
rect 2255 2065 2259 2069
rect 2343 2065 2347 2069
rect 2439 2065 2443 2069
rect 2527 2065 2531 2069
rect 2583 2064 2587 2068
rect 111 2051 115 2055
rect 1327 2051 1331 2055
rect 1367 2047 1371 2051
rect 159 2042 163 2046
rect 215 2042 219 2046
rect 287 2042 291 2046
rect 383 2042 387 2046
rect 479 2042 483 2046
rect 583 2042 587 2046
rect 679 2042 683 2046
rect 775 2042 779 2046
rect 863 2042 867 2046
rect 943 2042 947 2046
rect 1023 2042 1027 2046
rect 1111 2042 1115 2046
rect 2583 2047 2587 2051
rect 1199 2042 1203 2046
rect 1503 2038 1507 2042
rect 1599 2038 1603 2042
rect 1695 2038 1699 2042
rect 1799 2038 1803 2042
rect 1903 2038 1907 2042
rect 1999 2038 2003 2042
rect 2095 2038 2099 2042
rect 2183 2038 2187 2042
rect 2271 2038 2275 2042
rect 2359 2038 2363 2042
rect 2455 2038 2459 2042
rect 2543 2038 2547 2042
rect 175 2010 179 2014
rect 239 2010 243 2014
rect 311 2010 315 2014
rect 391 2010 395 2014
rect 471 2010 475 2014
rect 559 2010 563 2014
rect 647 2010 651 2014
rect 735 2010 739 2014
rect 823 2010 827 2014
rect 911 2010 915 2014
rect 1007 2010 1011 2014
rect 1103 2010 1107 2014
rect 1415 2014 1419 2018
rect 1471 2014 1475 2018
rect 1535 2014 1539 2018
rect 1615 2014 1619 2018
rect 1703 2014 1707 2018
rect 1791 2014 1795 2018
rect 1887 2014 1891 2018
rect 1983 2014 1987 2018
rect 2079 2014 2083 2018
rect 2175 2014 2179 2018
rect 2271 2014 2275 2018
rect 2367 2014 2371 2018
rect 2463 2014 2467 2018
rect 2543 2014 2547 2018
rect 111 2001 115 2005
rect 1327 2001 1331 2005
rect 1367 2005 1371 2009
rect 2583 2005 2587 2009
rect 111 1984 115 1988
rect 159 1983 163 1987
rect 223 1983 227 1987
rect 295 1983 299 1987
rect 375 1983 379 1987
rect 455 1983 459 1987
rect 543 1983 547 1987
rect 631 1983 635 1987
rect 719 1983 723 1987
rect 807 1983 811 1987
rect 895 1983 899 1987
rect 991 1983 995 1987
rect 1087 1983 1091 1987
rect 1327 1984 1331 1988
rect 1367 1988 1371 1992
rect 1399 1987 1403 1991
rect 1455 1987 1459 1991
rect 1519 1987 1523 1991
rect 1599 1987 1603 1991
rect 1687 1987 1691 1991
rect 1775 1987 1779 1991
rect 1871 1987 1875 1991
rect 1967 1987 1971 1991
rect 2063 1987 2067 1991
rect 2159 1987 2163 1991
rect 2255 1987 2259 1991
rect 2351 1987 2355 1991
rect 2447 1987 2451 1991
rect 2527 1987 2531 1991
rect 2583 1988 2587 1992
rect 111 1948 115 1952
rect 383 1949 387 1953
rect 439 1949 443 1953
rect 495 1949 499 1953
rect 551 1949 555 1953
rect 607 1949 611 1953
rect 671 1949 675 1953
rect 735 1949 739 1953
rect 807 1949 811 1953
rect 879 1949 883 1953
rect 951 1949 955 1953
rect 1023 1949 1027 1953
rect 1327 1948 1331 1952
rect 1367 1948 1371 1952
rect 1399 1949 1403 1953
rect 1455 1949 1459 1953
rect 1519 1949 1523 1953
rect 1599 1949 1603 1953
rect 1679 1949 1683 1953
rect 1759 1949 1763 1953
rect 1855 1949 1859 1953
rect 1967 1949 1971 1953
rect 2095 1949 2099 1953
rect 2239 1949 2243 1953
rect 2391 1949 2395 1953
rect 2527 1949 2531 1953
rect 2583 1948 2587 1952
rect 111 1931 115 1935
rect 1327 1931 1331 1935
rect 1367 1931 1371 1935
rect 2583 1931 2587 1935
rect 399 1922 403 1926
rect 455 1922 459 1926
rect 511 1922 515 1926
rect 567 1922 571 1926
rect 623 1922 627 1926
rect 687 1922 691 1926
rect 751 1922 755 1926
rect 823 1922 827 1926
rect 895 1922 899 1926
rect 967 1922 971 1926
rect 1039 1922 1043 1926
rect 1415 1922 1419 1926
rect 1471 1922 1475 1926
rect 1535 1922 1539 1926
rect 1615 1922 1619 1926
rect 1695 1922 1699 1926
rect 1775 1922 1779 1926
rect 1871 1922 1875 1926
rect 1983 1922 1987 1926
rect 2111 1922 2115 1926
rect 2255 1922 2259 1926
rect 2407 1922 2411 1926
rect 2543 1922 2547 1926
rect 519 1898 523 1902
rect 575 1898 579 1902
rect 631 1898 635 1902
rect 687 1898 691 1902
rect 743 1898 747 1902
rect 807 1898 811 1902
rect 871 1898 875 1902
rect 935 1898 939 1902
rect 999 1898 1003 1902
rect 1575 1898 1579 1902
rect 1631 1898 1635 1902
rect 1687 1898 1691 1902
rect 1743 1898 1747 1902
rect 1799 1898 1803 1902
rect 1855 1898 1859 1902
rect 1927 1898 1931 1902
rect 2015 1898 2019 1902
rect 2127 1898 2131 1902
rect 2247 1898 2251 1902
rect 2383 1898 2387 1902
rect 2519 1898 2523 1902
rect 111 1889 115 1893
rect 1327 1889 1331 1893
rect 1367 1889 1371 1893
rect 2583 1889 2587 1893
rect 111 1872 115 1876
rect 503 1871 507 1875
rect 559 1871 563 1875
rect 615 1871 619 1875
rect 671 1871 675 1875
rect 727 1871 731 1875
rect 791 1871 795 1875
rect 855 1871 859 1875
rect 919 1871 923 1875
rect 983 1871 987 1875
rect 1327 1872 1331 1876
rect 1367 1872 1371 1876
rect 1559 1871 1563 1875
rect 1615 1871 1619 1875
rect 1671 1871 1675 1875
rect 1727 1871 1731 1875
rect 1783 1871 1787 1875
rect 1839 1871 1843 1875
rect 1911 1871 1915 1875
rect 1999 1871 2003 1875
rect 2111 1871 2115 1875
rect 2231 1871 2235 1875
rect 2367 1871 2371 1875
rect 2503 1871 2507 1875
rect 2583 1872 2587 1876
rect 111 1832 115 1836
rect 143 1833 147 1837
rect 199 1833 203 1837
rect 255 1833 259 1837
rect 311 1833 315 1837
rect 375 1833 379 1837
rect 455 1833 459 1837
rect 543 1833 547 1837
rect 631 1833 635 1837
rect 719 1833 723 1837
rect 799 1833 803 1837
rect 887 1833 891 1837
rect 975 1833 979 1837
rect 1063 1833 1067 1837
rect 1327 1832 1331 1836
rect 1367 1828 1371 1832
rect 1623 1829 1627 1833
rect 1679 1829 1683 1833
rect 1735 1829 1739 1833
rect 1791 1829 1795 1833
rect 1847 1829 1851 1833
rect 1903 1829 1907 1833
rect 1967 1829 1971 1833
rect 2039 1829 2043 1833
rect 2127 1829 2131 1833
rect 2223 1829 2227 1833
rect 2327 1829 2331 1833
rect 2439 1829 2443 1833
rect 2527 1829 2531 1833
rect 2583 1828 2587 1832
rect 111 1815 115 1819
rect 1327 1815 1331 1819
rect 1367 1811 1371 1815
rect 159 1806 163 1810
rect 215 1806 219 1810
rect 271 1806 275 1810
rect 327 1806 331 1810
rect 391 1806 395 1810
rect 471 1806 475 1810
rect 559 1806 563 1810
rect 647 1806 651 1810
rect 735 1806 739 1810
rect 815 1806 819 1810
rect 903 1806 907 1810
rect 991 1806 995 1810
rect 2583 1811 2587 1815
rect 1079 1806 1083 1810
rect 1639 1802 1643 1806
rect 1695 1802 1699 1806
rect 1751 1802 1755 1806
rect 1807 1802 1811 1806
rect 1863 1802 1867 1806
rect 1919 1802 1923 1806
rect 1983 1802 1987 1806
rect 2055 1802 2059 1806
rect 2143 1802 2147 1806
rect 2239 1802 2243 1806
rect 2343 1802 2347 1806
rect 2455 1802 2459 1806
rect 2543 1802 2547 1806
rect 159 1774 163 1778
rect 255 1774 259 1778
rect 375 1774 379 1778
rect 503 1774 507 1778
rect 623 1774 627 1778
rect 743 1774 747 1778
rect 855 1774 859 1778
rect 959 1774 963 1778
rect 1055 1774 1059 1778
rect 1151 1774 1155 1778
rect 1247 1774 1251 1778
rect 1471 1770 1475 1774
rect 111 1765 115 1769
rect 1535 1770 1539 1774
rect 1615 1770 1619 1774
rect 1695 1770 1699 1774
rect 1783 1770 1787 1774
rect 1879 1770 1883 1774
rect 1975 1770 1979 1774
rect 2071 1770 2075 1774
rect 2167 1770 2171 1774
rect 2263 1770 2267 1774
rect 2359 1770 2363 1774
rect 2463 1770 2467 1774
rect 2543 1770 2547 1774
rect 1327 1765 1331 1769
rect 1367 1761 1371 1765
rect 2583 1761 2587 1765
rect 111 1748 115 1752
rect 143 1747 147 1751
rect 239 1747 243 1751
rect 359 1747 363 1751
rect 487 1747 491 1751
rect 607 1747 611 1751
rect 727 1747 731 1751
rect 839 1747 843 1751
rect 943 1747 947 1751
rect 1039 1747 1043 1751
rect 1135 1747 1139 1751
rect 1231 1747 1235 1751
rect 1327 1748 1331 1752
rect 1367 1744 1371 1748
rect 1455 1743 1459 1747
rect 1519 1743 1523 1747
rect 1599 1743 1603 1747
rect 1679 1743 1683 1747
rect 1767 1743 1771 1747
rect 1863 1743 1867 1747
rect 1959 1743 1963 1747
rect 2055 1743 2059 1747
rect 2151 1743 2155 1747
rect 2247 1743 2251 1747
rect 2343 1743 2347 1747
rect 2447 1743 2451 1747
rect 2527 1743 2531 1747
rect 2583 1744 2587 1748
rect 111 1712 115 1716
rect 143 1713 147 1717
rect 263 1713 267 1717
rect 415 1713 419 1717
rect 567 1713 571 1717
rect 711 1713 715 1717
rect 855 1713 859 1717
rect 999 1713 1003 1717
rect 1143 1713 1147 1717
rect 1271 1713 1275 1717
rect 1327 1712 1331 1716
rect 1367 1704 1371 1708
rect 1399 1705 1403 1709
rect 1479 1705 1483 1709
rect 1599 1705 1603 1709
rect 1719 1705 1723 1709
rect 1839 1705 1843 1709
rect 1951 1705 1955 1709
rect 2055 1705 2059 1709
rect 2159 1705 2163 1709
rect 2255 1705 2259 1709
rect 2351 1705 2355 1709
rect 2447 1705 2451 1709
rect 2527 1705 2531 1709
rect 2583 1704 2587 1708
rect 111 1695 115 1699
rect 1327 1695 1331 1699
rect 159 1686 163 1690
rect 279 1686 283 1690
rect 431 1686 435 1690
rect 583 1686 587 1690
rect 727 1686 731 1690
rect 871 1686 875 1690
rect 1015 1686 1019 1690
rect 1159 1686 1163 1690
rect 1287 1686 1291 1690
rect 1367 1687 1371 1691
rect 2583 1687 2587 1691
rect 1415 1678 1419 1682
rect 1495 1678 1499 1682
rect 1615 1678 1619 1682
rect 1735 1678 1739 1682
rect 1855 1678 1859 1682
rect 1967 1678 1971 1682
rect 2071 1678 2075 1682
rect 2175 1678 2179 1682
rect 2271 1678 2275 1682
rect 2367 1678 2371 1682
rect 2463 1678 2467 1682
rect 2543 1678 2547 1682
rect 159 1658 163 1662
rect 223 1658 227 1662
rect 303 1658 307 1662
rect 383 1658 387 1662
rect 463 1658 467 1662
rect 535 1658 539 1662
rect 607 1658 611 1662
rect 679 1658 683 1662
rect 767 1658 771 1662
rect 863 1658 867 1662
rect 967 1658 971 1662
rect 1079 1658 1083 1662
rect 1191 1658 1195 1662
rect 1287 1658 1291 1662
rect 1415 1654 1419 1658
rect 111 1649 115 1653
rect 1503 1654 1507 1658
rect 1623 1654 1627 1658
rect 1751 1654 1755 1658
rect 1879 1654 1883 1658
rect 1999 1654 2003 1658
rect 2119 1654 2123 1658
rect 2231 1654 2235 1658
rect 2343 1654 2347 1658
rect 2455 1654 2459 1658
rect 2543 1654 2547 1658
rect 1327 1649 1331 1653
rect 1367 1645 1371 1649
rect 2583 1645 2587 1649
rect 111 1632 115 1636
rect 143 1631 147 1635
rect 207 1631 211 1635
rect 287 1631 291 1635
rect 367 1631 371 1635
rect 447 1631 451 1635
rect 519 1631 523 1635
rect 591 1631 595 1635
rect 663 1631 667 1635
rect 751 1631 755 1635
rect 847 1631 851 1635
rect 951 1631 955 1635
rect 1063 1631 1067 1635
rect 1175 1631 1179 1635
rect 1271 1631 1275 1635
rect 1327 1632 1331 1636
rect 1367 1628 1371 1632
rect 1399 1627 1403 1631
rect 1487 1627 1491 1631
rect 1607 1627 1611 1631
rect 1735 1627 1739 1631
rect 1863 1627 1867 1631
rect 1983 1627 1987 1631
rect 2103 1627 2107 1631
rect 2215 1627 2219 1631
rect 2327 1627 2331 1631
rect 2439 1627 2443 1631
rect 2527 1627 2531 1631
rect 2583 1628 2587 1632
rect 111 1596 115 1600
rect 143 1597 147 1601
rect 247 1597 251 1601
rect 367 1597 371 1601
rect 479 1597 483 1601
rect 575 1597 579 1601
rect 671 1597 675 1601
rect 767 1597 771 1601
rect 863 1597 867 1601
rect 959 1597 963 1601
rect 1063 1597 1067 1601
rect 1175 1597 1179 1601
rect 1271 1597 1275 1601
rect 1327 1596 1331 1600
rect 111 1579 115 1583
rect 1327 1579 1331 1583
rect 1367 1580 1371 1584
rect 1399 1581 1403 1585
rect 1495 1581 1499 1585
rect 1615 1581 1619 1585
rect 1743 1581 1747 1585
rect 1863 1581 1867 1585
rect 1983 1581 1987 1585
rect 2095 1581 2099 1585
rect 2199 1581 2203 1585
rect 2295 1581 2299 1585
rect 2391 1581 2395 1585
rect 2495 1581 2499 1585
rect 2583 1580 2587 1584
rect 159 1570 163 1574
rect 263 1570 267 1574
rect 383 1570 387 1574
rect 495 1570 499 1574
rect 591 1570 595 1574
rect 687 1570 691 1574
rect 783 1570 787 1574
rect 879 1570 883 1574
rect 975 1570 979 1574
rect 1079 1570 1083 1574
rect 1191 1570 1195 1574
rect 1287 1570 1291 1574
rect 1367 1563 1371 1567
rect 2583 1563 2587 1567
rect 1415 1554 1419 1558
rect 1511 1554 1515 1558
rect 1631 1554 1635 1558
rect 1759 1554 1763 1558
rect 1879 1554 1883 1558
rect 1999 1554 2003 1558
rect 2111 1554 2115 1558
rect 2215 1554 2219 1558
rect 2311 1554 2315 1558
rect 2407 1554 2411 1558
rect 2511 1554 2515 1558
rect 159 1542 163 1546
rect 231 1542 235 1546
rect 335 1542 339 1546
rect 455 1542 459 1546
rect 583 1542 587 1546
rect 719 1542 723 1546
rect 863 1542 867 1546
rect 1007 1542 1011 1546
rect 1151 1542 1155 1546
rect 1287 1542 1291 1546
rect 111 1533 115 1537
rect 1327 1533 1331 1537
rect 1415 1526 1419 1530
rect 1527 1526 1531 1530
rect 1647 1526 1651 1530
rect 1767 1526 1771 1530
rect 1879 1526 1883 1530
rect 1983 1526 1987 1530
rect 2079 1526 2083 1530
rect 2167 1526 2171 1530
rect 2255 1526 2259 1530
rect 2335 1526 2339 1530
rect 2407 1526 2411 1530
rect 2487 1526 2491 1530
rect 2543 1526 2547 1530
rect 111 1516 115 1520
rect 143 1515 147 1519
rect 215 1515 219 1519
rect 319 1515 323 1519
rect 439 1515 443 1519
rect 567 1515 571 1519
rect 703 1515 707 1519
rect 847 1515 851 1519
rect 991 1515 995 1519
rect 1135 1515 1139 1519
rect 1271 1515 1275 1519
rect 1327 1516 1331 1520
rect 1367 1517 1371 1521
rect 2583 1517 2587 1521
rect 1367 1500 1371 1504
rect 1399 1499 1403 1503
rect 1511 1499 1515 1503
rect 1631 1499 1635 1503
rect 1751 1499 1755 1503
rect 1863 1499 1867 1503
rect 1967 1499 1971 1503
rect 2063 1499 2067 1503
rect 2151 1499 2155 1503
rect 2239 1499 2243 1503
rect 2319 1499 2323 1503
rect 2391 1499 2395 1503
rect 2471 1499 2475 1503
rect 2527 1499 2531 1503
rect 2583 1500 2587 1504
rect 111 1480 115 1484
rect 143 1481 147 1485
rect 199 1481 203 1485
rect 271 1481 275 1485
rect 367 1481 371 1485
rect 479 1481 483 1485
rect 591 1481 595 1485
rect 703 1481 707 1485
rect 807 1481 811 1485
rect 911 1481 915 1485
rect 1007 1481 1011 1485
rect 1103 1481 1107 1485
rect 1199 1481 1203 1485
rect 1271 1481 1275 1485
rect 1327 1480 1331 1484
rect 111 1463 115 1467
rect 1327 1463 1331 1467
rect 159 1454 163 1458
rect 215 1454 219 1458
rect 287 1454 291 1458
rect 383 1454 387 1458
rect 495 1454 499 1458
rect 607 1454 611 1458
rect 719 1454 723 1458
rect 823 1454 827 1458
rect 927 1454 931 1458
rect 1023 1454 1027 1458
rect 1119 1454 1123 1458
rect 1215 1454 1219 1458
rect 1287 1454 1291 1458
rect 1367 1456 1371 1460
rect 1399 1457 1403 1461
rect 1503 1457 1507 1461
rect 1631 1457 1635 1461
rect 1751 1457 1755 1461
rect 1871 1457 1875 1461
rect 1983 1457 1987 1461
rect 2087 1457 2091 1461
rect 2183 1457 2187 1461
rect 2271 1457 2275 1461
rect 2359 1457 2363 1461
rect 2455 1457 2459 1461
rect 2527 1457 2531 1461
rect 2583 1456 2587 1460
rect 1367 1439 1371 1443
rect 2583 1439 2587 1443
rect 255 1426 259 1430
rect 311 1426 315 1430
rect 375 1426 379 1430
rect 447 1426 451 1430
rect 527 1426 531 1430
rect 607 1426 611 1430
rect 695 1426 699 1430
rect 783 1426 787 1430
rect 871 1426 875 1430
rect 959 1426 963 1430
rect 1055 1426 1059 1430
rect 1151 1426 1155 1430
rect 1415 1430 1419 1434
rect 1519 1430 1523 1434
rect 1647 1430 1651 1434
rect 1767 1430 1771 1434
rect 1887 1430 1891 1434
rect 1999 1430 2003 1434
rect 2103 1430 2107 1434
rect 2199 1430 2203 1434
rect 2287 1430 2291 1434
rect 2375 1430 2379 1434
rect 2471 1430 2475 1434
rect 2543 1430 2547 1434
rect 111 1417 115 1421
rect 1327 1417 1331 1421
rect 111 1400 115 1404
rect 239 1399 243 1403
rect 295 1399 299 1403
rect 359 1399 363 1403
rect 431 1399 435 1403
rect 511 1399 515 1403
rect 591 1399 595 1403
rect 679 1399 683 1403
rect 767 1399 771 1403
rect 855 1399 859 1403
rect 943 1399 947 1403
rect 1039 1399 1043 1403
rect 1135 1399 1139 1403
rect 1327 1400 1331 1404
rect 1415 1402 1419 1406
rect 1471 1402 1475 1406
rect 1551 1402 1555 1406
rect 1631 1402 1635 1406
rect 1711 1402 1715 1406
rect 1791 1402 1795 1406
rect 1871 1402 1875 1406
rect 1959 1402 1963 1406
rect 2055 1402 2059 1406
rect 2167 1402 2171 1406
rect 2295 1402 2299 1406
rect 2431 1402 2435 1406
rect 2543 1402 2547 1406
rect 1367 1393 1371 1397
rect 2583 1393 2587 1397
rect 1367 1376 1371 1380
rect 1399 1375 1403 1379
rect 1455 1375 1459 1379
rect 1535 1375 1539 1379
rect 1615 1375 1619 1379
rect 1695 1375 1699 1379
rect 1775 1375 1779 1379
rect 1855 1375 1859 1379
rect 1943 1375 1947 1379
rect 2039 1375 2043 1379
rect 2151 1375 2155 1379
rect 2279 1375 2283 1379
rect 2415 1375 2419 1379
rect 2527 1375 2531 1379
rect 2583 1376 2587 1380
rect 111 1356 115 1360
rect 359 1357 363 1361
rect 415 1357 419 1361
rect 471 1357 475 1361
rect 527 1357 531 1361
rect 591 1357 595 1361
rect 671 1357 675 1361
rect 751 1357 755 1361
rect 839 1357 843 1361
rect 935 1357 939 1361
rect 1031 1357 1035 1361
rect 1127 1357 1131 1361
rect 1231 1357 1235 1361
rect 1327 1356 1331 1360
rect 111 1339 115 1343
rect 1327 1339 1331 1343
rect 1367 1340 1371 1344
rect 1423 1341 1427 1345
rect 1495 1341 1499 1345
rect 1575 1341 1579 1345
rect 1655 1341 1659 1345
rect 1759 1341 1763 1345
rect 1879 1341 1883 1345
rect 2023 1341 2027 1345
rect 2183 1341 2187 1345
rect 2359 1341 2363 1345
rect 2527 1341 2531 1345
rect 2583 1340 2587 1344
rect 375 1330 379 1334
rect 431 1330 435 1334
rect 487 1330 491 1334
rect 543 1330 547 1334
rect 607 1330 611 1334
rect 687 1330 691 1334
rect 767 1330 771 1334
rect 855 1330 859 1334
rect 951 1330 955 1334
rect 1047 1330 1051 1334
rect 1143 1330 1147 1334
rect 1247 1330 1251 1334
rect 1367 1323 1371 1327
rect 2583 1323 2587 1327
rect 1439 1314 1443 1318
rect 1511 1314 1515 1318
rect 1591 1314 1595 1318
rect 1671 1314 1675 1318
rect 1775 1314 1779 1318
rect 1895 1314 1899 1318
rect 2039 1314 2043 1318
rect 2199 1314 2203 1318
rect 2375 1314 2379 1318
rect 2543 1314 2547 1318
rect 471 1298 475 1302
rect 527 1298 531 1302
rect 583 1298 587 1302
rect 647 1298 651 1302
rect 727 1298 731 1302
rect 807 1298 811 1302
rect 895 1298 899 1302
rect 991 1298 995 1302
rect 1095 1298 1099 1302
rect 1199 1298 1203 1302
rect 1287 1298 1291 1302
rect 111 1289 115 1293
rect 1327 1289 1331 1293
rect 1431 1290 1435 1294
rect 1495 1290 1499 1294
rect 1559 1290 1563 1294
rect 1631 1290 1635 1294
rect 1703 1290 1707 1294
rect 1775 1290 1779 1294
rect 1855 1290 1859 1294
rect 1943 1290 1947 1294
rect 2047 1290 2051 1294
rect 2159 1290 2163 1294
rect 2287 1290 2291 1294
rect 2423 1290 2427 1294
rect 2543 1290 2547 1294
rect 1367 1281 1371 1285
rect 2583 1281 2587 1285
rect 111 1272 115 1276
rect 455 1271 459 1275
rect 511 1271 515 1275
rect 567 1271 571 1275
rect 631 1271 635 1275
rect 711 1271 715 1275
rect 791 1271 795 1275
rect 879 1271 883 1275
rect 975 1271 979 1275
rect 1079 1271 1083 1275
rect 1183 1271 1187 1275
rect 1271 1271 1275 1275
rect 1327 1272 1331 1276
rect 1367 1264 1371 1268
rect 1415 1263 1419 1267
rect 1479 1263 1483 1267
rect 1543 1263 1547 1267
rect 1615 1263 1619 1267
rect 1687 1263 1691 1267
rect 1759 1263 1763 1267
rect 1839 1263 1843 1267
rect 1927 1263 1931 1267
rect 2031 1263 2035 1267
rect 2143 1263 2147 1267
rect 2271 1263 2275 1267
rect 2407 1263 2411 1267
rect 2527 1263 2531 1267
rect 2583 1264 2587 1268
rect 111 1232 115 1236
rect 383 1233 387 1237
rect 439 1233 443 1237
rect 503 1233 507 1237
rect 575 1233 579 1237
rect 647 1233 651 1237
rect 727 1233 731 1237
rect 815 1233 819 1237
rect 903 1233 907 1237
rect 991 1233 995 1237
rect 1079 1233 1083 1237
rect 1175 1233 1179 1237
rect 1271 1233 1275 1237
rect 1327 1232 1331 1236
rect 1367 1224 1371 1228
rect 1399 1225 1403 1229
rect 1455 1225 1459 1229
rect 1535 1225 1539 1229
rect 1615 1225 1619 1229
rect 1695 1225 1699 1229
rect 1775 1225 1779 1229
rect 1855 1225 1859 1229
rect 1943 1225 1947 1229
rect 2039 1225 2043 1229
rect 2151 1225 2155 1229
rect 2279 1225 2283 1229
rect 2415 1225 2419 1229
rect 2527 1225 2531 1229
rect 2583 1224 2587 1228
rect 111 1215 115 1219
rect 1327 1215 1331 1219
rect 399 1206 403 1210
rect 455 1206 459 1210
rect 519 1206 523 1210
rect 591 1206 595 1210
rect 663 1206 667 1210
rect 743 1206 747 1210
rect 831 1206 835 1210
rect 919 1206 923 1210
rect 1007 1206 1011 1210
rect 1095 1206 1099 1210
rect 1191 1206 1195 1210
rect 1287 1206 1291 1210
rect 1367 1207 1371 1211
rect 2583 1207 2587 1211
rect 1415 1198 1419 1202
rect 1471 1198 1475 1202
rect 1551 1198 1555 1202
rect 1631 1198 1635 1202
rect 1711 1198 1715 1202
rect 1791 1198 1795 1202
rect 1871 1198 1875 1202
rect 1959 1198 1963 1202
rect 2055 1198 2059 1202
rect 2167 1198 2171 1202
rect 2295 1198 2299 1202
rect 2431 1198 2435 1202
rect 2543 1198 2547 1202
rect 279 1178 283 1182
rect 343 1178 347 1182
rect 415 1178 419 1182
rect 495 1178 499 1182
rect 583 1178 587 1182
rect 671 1178 675 1182
rect 759 1178 763 1182
rect 847 1178 851 1182
rect 935 1178 939 1182
rect 1015 1178 1019 1182
rect 1087 1178 1091 1182
rect 1159 1178 1163 1182
rect 1231 1178 1235 1182
rect 1287 1178 1291 1182
rect 111 1169 115 1173
rect 1327 1169 1331 1173
rect 1695 1166 1699 1170
rect 1767 1166 1771 1170
rect 1847 1166 1851 1170
rect 1919 1166 1923 1170
rect 1991 1166 1995 1170
rect 2063 1166 2067 1170
rect 2135 1166 2139 1170
rect 2207 1166 2211 1170
rect 2287 1166 2291 1170
rect 2367 1166 2371 1170
rect 1367 1157 1371 1161
rect 2583 1157 2587 1161
rect 111 1152 115 1156
rect 263 1151 267 1155
rect 327 1151 331 1155
rect 399 1151 403 1155
rect 479 1151 483 1155
rect 567 1151 571 1155
rect 655 1151 659 1155
rect 743 1151 747 1155
rect 831 1151 835 1155
rect 919 1151 923 1155
rect 999 1151 1003 1155
rect 1071 1151 1075 1155
rect 1143 1151 1147 1155
rect 1215 1151 1219 1155
rect 1271 1151 1275 1155
rect 1327 1152 1331 1156
rect 1367 1140 1371 1144
rect 1679 1139 1683 1143
rect 1751 1139 1755 1143
rect 1831 1139 1835 1143
rect 1903 1139 1907 1143
rect 1975 1139 1979 1143
rect 2047 1139 2051 1143
rect 2119 1139 2123 1143
rect 2191 1139 2195 1143
rect 2271 1139 2275 1143
rect 2351 1139 2355 1143
rect 2583 1140 2587 1144
rect 111 1108 115 1112
rect 143 1109 147 1113
rect 207 1109 211 1113
rect 271 1109 275 1113
rect 343 1109 347 1113
rect 423 1109 427 1113
rect 503 1109 507 1113
rect 583 1109 587 1113
rect 663 1109 667 1113
rect 743 1109 747 1113
rect 831 1109 835 1113
rect 919 1109 923 1113
rect 1007 1109 1011 1113
rect 1327 1108 1331 1112
rect 1367 1104 1371 1108
rect 1399 1105 1403 1109
rect 1479 1105 1483 1109
rect 1583 1105 1587 1109
rect 1687 1105 1691 1109
rect 1783 1105 1787 1109
rect 1879 1105 1883 1109
rect 1975 1105 1979 1109
rect 2063 1105 2067 1109
rect 2151 1105 2155 1109
rect 2239 1105 2243 1109
rect 2327 1105 2331 1109
rect 2415 1105 2419 1109
rect 2583 1104 2587 1108
rect 111 1091 115 1095
rect 1327 1091 1331 1095
rect 1367 1087 1371 1091
rect 159 1082 163 1086
rect 223 1082 227 1086
rect 287 1082 291 1086
rect 359 1082 363 1086
rect 439 1082 443 1086
rect 519 1082 523 1086
rect 599 1082 603 1086
rect 679 1082 683 1086
rect 759 1082 763 1086
rect 847 1082 851 1086
rect 935 1082 939 1086
rect 2583 1087 2587 1091
rect 1023 1082 1027 1086
rect 1415 1078 1419 1082
rect 1495 1078 1499 1082
rect 1599 1078 1603 1082
rect 1703 1078 1707 1082
rect 1799 1078 1803 1082
rect 1895 1078 1899 1082
rect 1991 1078 1995 1082
rect 2079 1078 2083 1082
rect 2167 1078 2171 1082
rect 2255 1078 2259 1082
rect 2343 1078 2347 1082
rect 2431 1078 2435 1082
rect 159 1054 163 1058
rect 215 1054 219 1058
rect 287 1054 291 1058
rect 383 1054 387 1058
rect 479 1054 483 1058
rect 583 1054 587 1058
rect 687 1054 691 1058
rect 783 1054 787 1058
rect 879 1054 883 1058
rect 967 1054 971 1058
rect 1063 1054 1067 1058
rect 1159 1054 1163 1058
rect 1415 1054 1419 1058
rect 1511 1054 1515 1058
rect 1631 1054 1635 1058
rect 1751 1054 1755 1058
rect 1871 1054 1875 1058
rect 1991 1054 1995 1058
rect 2103 1054 2107 1058
rect 2199 1054 2203 1058
rect 2295 1054 2299 1058
rect 2383 1054 2387 1058
rect 2471 1054 2475 1058
rect 2543 1054 2547 1058
rect 111 1045 115 1049
rect 1327 1045 1331 1049
rect 1367 1045 1371 1049
rect 2583 1045 2587 1049
rect 111 1028 115 1032
rect 143 1027 147 1031
rect 199 1027 203 1031
rect 271 1027 275 1031
rect 367 1027 371 1031
rect 463 1027 467 1031
rect 567 1027 571 1031
rect 671 1027 675 1031
rect 767 1027 771 1031
rect 863 1027 867 1031
rect 951 1027 955 1031
rect 1047 1027 1051 1031
rect 1143 1027 1147 1031
rect 1327 1028 1331 1032
rect 1367 1028 1371 1032
rect 1399 1027 1403 1031
rect 1495 1027 1499 1031
rect 1615 1027 1619 1031
rect 1735 1027 1739 1031
rect 1855 1027 1859 1031
rect 1975 1027 1979 1031
rect 2087 1027 2091 1031
rect 2183 1027 2187 1031
rect 2279 1027 2283 1031
rect 2367 1027 2371 1031
rect 2455 1027 2459 1031
rect 2527 1027 2531 1031
rect 2583 1028 2587 1032
rect 111 988 115 992
rect 143 989 147 993
rect 199 989 203 993
rect 279 989 283 993
rect 383 989 387 993
rect 495 989 499 993
rect 615 989 619 993
rect 727 989 731 993
rect 839 989 843 993
rect 951 989 955 993
rect 1055 989 1059 993
rect 1159 989 1163 993
rect 1271 989 1275 993
rect 1327 988 1331 992
rect 1367 988 1371 992
rect 1487 989 1491 993
rect 1583 989 1587 993
rect 1695 989 1699 993
rect 1807 989 1811 993
rect 1919 989 1923 993
rect 2023 989 2027 993
rect 2119 989 2123 993
rect 2215 989 2219 993
rect 2303 989 2307 993
rect 2383 989 2387 993
rect 2463 989 2467 993
rect 2527 989 2531 993
rect 2583 988 2587 992
rect 111 971 115 975
rect 1327 971 1331 975
rect 1367 971 1371 975
rect 2583 971 2587 975
rect 159 962 163 966
rect 215 962 219 966
rect 295 962 299 966
rect 399 962 403 966
rect 511 962 515 966
rect 631 962 635 966
rect 743 962 747 966
rect 855 962 859 966
rect 967 962 971 966
rect 1071 962 1075 966
rect 1175 962 1179 966
rect 1287 962 1291 966
rect 1503 962 1507 966
rect 1599 962 1603 966
rect 1711 962 1715 966
rect 1823 962 1827 966
rect 1935 962 1939 966
rect 2039 962 2043 966
rect 2135 962 2139 966
rect 2231 962 2235 966
rect 2319 962 2323 966
rect 2399 962 2403 966
rect 2479 962 2483 966
rect 2543 962 2547 966
rect 159 930 163 934
rect 215 930 219 934
rect 287 930 291 934
rect 375 930 379 934
rect 471 930 475 934
rect 567 930 571 934
rect 671 930 675 934
rect 767 930 771 934
rect 863 930 867 934
rect 959 930 963 934
rect 1047 930 1051 934
rect 1135 930 1139 934
rect 1223 930 1227 934
rect 1287 930 1291 934
rect 1415 930 1419 934
rect 1535 930 1539 934
rect 1671 930 1675 934
rect 1807 930 1811 934
rect 1935 930 1939 934
rect 2055 930 2059 934
rect 2167 930 2171 934
rect 2271 930 2275 934
rect 2367 930 2371 934
rect 2463 930 2467 934
rect 2543 930 2547 934
rect 111 921 115 925
rect 1327 921 1331 925
rect 1367 921 1371 925
rect 2583 921 2587 925
rect 111 904 115 908
rect 143 903 147 907
rect 199 903 203 907
rect 271 903 275 907
rect 359 903 363 907
rect 455 903 459 907
rect 551 903 555 907
rect 655 903 659 907
rect 751 903 755 907
rect 847 903 851 907
rect 943 903 947 907
rect 1031 903 1035 907
rect 1119 903 1123 907
rect 1207 903 1211 907
rect 1271 903 1275 907
rect 1327 904 1331 908
rect 1367 904 1371 908
rect 1399 903 1403 907
rect 1519 903 1523 907
rect 1655 903 1659 907
rect 1791 903 1795 907
rect 1919 903 1923 907
rect 2039 903 2043 907
rect 2151 903 2155 907
rect 2255 903 2259 907
rect 2351 903 2355 907
rect 2447 903 2451 907
rect 2527 903 2531 907
rect 2583 904 2587 908
rect 111 864 115 868
rect 183 865 187 869
rect 239 865 243 869
rect 303 865 307 869
rect 375 865 379 869
rect 455 865 459 869
rect 543 865 547 869
rect 639 865 643 869
rect 743 865 747 869
rect 855 865 859 869
rect 967 865 971 869
rect 1087 865 1091 869
rect 1215 865 1219 869
rect 1327 864 1331 868
rect 1367 864 1371 868
rect 1399 865 1403 869
rect 1455 865 1459 869
rect 1519 865 1523 869
rect 1607 865 1611 869
rect 1695 865 1699 869
rect 1791 865 1795 869
rect 1895 865 1899 869
rect 1999 865 2003 869
rect 2103 865 2107 869
rect 2207 865 2211 869
rect 2311 865 2315 869
rect 2423 865 2427 869
rect 2527 865 2531 869
rect 2583 864 2587 868
rect 111 847 115 851
rect 1327 847 1331 851
rect 1367 847 1371 851
rect 2583 847 2587 851
rect 199 838 203 842
rect 255 838 259 842
rect 319 838 323 842
rect 391 838 395 842
rect 471 838 475 842
rect 559 838 563 842
rect 655 838 659 842
rect 759 838 763 842
rect 871 838 875 842
rect 983 838 987 842
rect 1103 838 1107 842
rect 1231 838 1235 842
rect 1415 838 1419 842
rect 1471 838 1475 842
rect 1535 838 1539 842
rect 1623 838 1627 842
rect 1711 838 1715 842
rect 1807 838 1811 842
rect 1911 838 1915 842
rect 2015 838 2019 842
rect 2119 838 2123 842
rect 2223 838 2227 842
rect 2327 838 2331 842
rect 2439 838 2443 842
rect 2543 838 2547 842
rect 383 806 387 810
rect 439 806 443 810
rect 495 806 499 810
rect 559 806 563 810
rect 631 806 635 810
rect 703 806 707 810
rect 783 806 787 810
rect 871 806 875 810
rect 959 806 963 810
rect 1047 806 1051 810
rect 1135 806 1139 810
rect 1223 806 1227 810
rect 1527 810 1531 814
rect 1583 810 1587 814
rect 1639 810 1643 814
rect 1695 810 1699 814
rect 1751 810 1755 814
rect 1807 810 1811 814
rect 1879 810 1883 814
rect 1959 810 1963 814
rect 2055 810 2059 814
rect 2167 810 2171 814
rect 2295 810 2299 814
rect 2431 810 2435 814
rect 2543 810 2547 814
rect 111 797 115 801
rect 1327 797 1331 801
rect 1367 801 1371 805
rect 2583 801 2587 805
rect 111 780 115 784
rect 367 779 371 783
rect 423 779 427 783
rect 479 779 483 783
rect 543 779 547 783
rect 615 779 619 783
rect 687 779 691 783
rect 767 779 771 783
rect 855 779 859 783
rect 943 779 947 783
rect 1031 779 1035 783
rect 1119 779 1123 783
rect 1207 779 1211 783
rect 1327 780 1331 784
rect 1367 784 1371 788
rect 1511 783 1515 787
rect 1567 783 1571 787
rect 1623 783 1627 787
rect 1679 783 1683 787
rect 1735 783 1739 787
rect 1791 783 1795 787
rect 1863 783 1867 787
rect 1943 783 1947 787
rect 2039 783 2043 787
rect 2151 783 2155 787
rect 2279 783 2283 787
rect 2415 783 2419 787
rect 2527 783 2531 787
rect 2583 784 2587 788
rect 111 744 115 748
rect 383 745 387 749
rect 439 745 443 749
rect 495 745 499 749
rect 559 745 563 749
rect 631 745 635 749
rect 711 745 715 749
rect 791 745 795 749
rect 871 745 875 749
rect 951 745 955 749
rect 1039 745 1043 749
rect 1127 745 1131 749
rect 1327 744 1331 748
rect 1367 740 1371 744
rect 1647 741 1651 745
rect 1703 741 1707 745
rect 1759 741 1763 745
rect 1815 741 1819 745
rect 1871 741 1875 745
rect 1927 741 1931 745
rect 1991 741 1995 745
rect 2063 741 2067 745
rect 2143 741 2147 745
rect 2231 741 2235 745
rect 2335 741 2339 745
rect 2439 741 2443 745
rect 2527 741 2531 745
rect 2583 740 2587 744
rect 111 727 115 731
rect 1327 727 1331 731
rect 1367 723 1371 727
rect 399 718 403 722
rect 455 718 459 722
rect 511 718 515 722
rect 575 718 579 722
rect 647 718 651 722
rect 727 718 731 722
rect 807 718 811 722
rect 887 718 891 722
rect 967 718 971 722
rect 1055 718 1059 722
rect 2583 723 2587 727
rect 1143 718 1147 722
rect 1663 714 1667 718
rect 1719 714 1723 718
rect 1775 714 1779 718
rect 1831 714 1835 718
rect 1887 714 1891 718
rect 1943 714 1947 718
rect 2007 714 2011 718
rect 2079 714 2083 718
rect 2159 714 2163 718
rect 2247 714 2251 718
rect 2351 714 2355 718
rect 2455 714 2459 718
rect 2543 714 2547 718
rect 343 694 347 698
rect 415 694 419 698
rect 487 694 491 698
rect 559 694 563 698
rect 631 694 635 698
rect 695 694 699 698
rect 759 694 763 698
rect 823 694 827 698
rect 887 694 891 698
rect 951 694 955 698
rect 1023 694 1027 698
rect 111 685 115 689
rect 1327 685 1331 689
rect 1735 686 1739 690
rect 1791 686 1795 690
rect 1855 686 1859 690
rect 1919 686 1923 690
rect 1991 686 1995 690
rect 2063 686 2067 690
rect 2127 686 2131 690
rect 2199 686 2203 690
rect 2271 686 2275 690
rect 2343 686 2347 690
rect 2415 686 2419 690
rect 2487 686 2491 690
rect 2543 686 2547 690
rect 1367 677 1371 681
rect 2583 677 2587 681
rect 111 668 115 672
rect 327 667 331 671
rect 399 667 403 671
rect 471 667 475 671
rect 543 667 547 671
rect 615 667 619 671
rect 679 667 683 671
rect 743 667 747 671
rect 807 667 811 671
rect 871 667 875 671
rect 935 667 939 671
rect 1007 667 1011 671
rect 1327 668 1331 672
rect 1367 660 1371 664
rect 1719 659 1723 663
rect 1775 659 1779 663
rect 1839 659 1843 663
rect 1903 659 1907 663
rect 1975 659 1979 663
rect 2047 659 2051 663
rect 2111 659 2115 663
rect 2183 659 2187 663
rect 2255 659 2259 663
rect 2327 659 2331 663
rect 2399 659 2403 663
rect 2471 659 2475 663
rect 2527 659 2531 663
rect 2583 660 2587 664
rect 111 628 115 632
rect 231 629 235 633
rect 295 629 299 633
rect 359 629 363 633
rect 423 629 427 633
rect 479 629 483 633
rect 535 629 539 633
rect 599 629 603 633
rect 663 629 667 633
rect 727 629 731 633
rect 791 629 795 633
rect 855 629 859 633
rect 919 629 923 633
rect 1327 628 1331 632
rect 1367 620 1371 624
rect 1615 621 1619 625
rect 1679 621 1683 625
rect 1759 621 1763 625
rect 1839 621 1843 625
rect 1927 621 1931 625
rect 2015 621 2019 625
rect 2095 621 2099 625
rect 2175 621 2179 625
rect 2255 621 2259 625
rect 2327 621 2331 625
rect 2399 621 2403 625
rect 2471 621 2475 625
rect 2527 621 2531 625
rect 2583 620 2587 624
rect 111 611 115 615
rect 1327 611 1331 615
rect 247 602 251 606
rect 311 602 315 606
rect 375 602 379 606
rect 439 602 443 606
rect 495 602 499 606
rect 551 602 555 606
rect 615 602 619 606
rect 679 602 683 606
rect 743 602 747 606
rect 807 602 811 606
rect 871 602 875 606
rect 935 602 939 606
rect 1367 603 1371 607
rect 2583 603 2587 607
rect 1631 594 1635 598
rect 1695 594 1699 598
rect 1775 594 1779 598
rect 1855 594 1859 598
rect 1943 594 1947 598
rect 2031 594 2035 598
rect 2111 594 2115 598
rect 2191 594 2195 598
rect 2271 594 2275 598
rect 2343 594 2347 598
rect 2415 594 2419 598
rect 2487 594 2491 598
rect 2543 594 2547 598
rect 191 570 195 574
rect 279 570 283 574
rect 367 570 371 574
rect 463 570 467 574
rect 559 570 563 574
rect 647 570 651 574
rect 735 570 739 574
rect 815 570 819 574
rect 887 570 891 574
rect 967 570 971 574
rect 1047 570 1051 574
rect 1127 570 1131 574
rect 111 561 115 565
rect 1327 561 1331 565
rect 1511 562 1515 566
rect 1575 562 1579 566
rect 1655 562 1659 566
rect 1735 562 1739 566
rect 1823 562 1827 566
rect 1911 562 1915 566
rect 1999 562 2003 566
rect 2087 562 2091 566
rect 2175 562 2179 566
rect 2271 562 2275 566
rect 2367 562 2371 566
rect 2463 562 2467 566
rect 2543 562 2547 566
rect 1367 553 1371 557
rect 2583 553 2587 557
rect 111 544 115 548
rect 175 543 179 547
rect 263 543 267 547
rect 351 543 355 547
rect 447 543 451 547
rect 543 543 547 547
rect 631 543 635 547
rect 719 543 723 547
rect 799 543 803 547
rect 871 543 875 547
rect 951 543 955 547
rect 1031 543 1035 547
rect 1111 543 1115 547
rect 1327 544 1331 548
rect 1367 536 1371 540
rect 1495 535 1499 539
rect 1559 535 1563 539
rect 1639 535 1643 539
rect 1719 535 1723 539
rect 1807 535 1811 539
rect 1895 535 1899 539
rect 1983 535 1987 539
rect 2071 535 2075 539
rect 2159 535 2163 539
rect 2255 535 2259 539
rect 2351 535 2355 539
rect 2447 535 2451 539
rect 2527 535 2531 539
rect 2583 536 2587 540
rect 111 504 115 508
rect 143 505 147 509
rect 207 505 211 509
rect 311 505 315 509
rect 431 505 435 509
rect 551 505 555 509
rect 671 505 675 509
rect 791 505 795 509
rect 903 505 907 509
rect 1007 505 1011 509
rect 1103 505 1107 509
rect 1199 505 1203 509
rect 1271 505 1275 509
rect 1327 504 1331 508
rect 1367 496 1371 500
rect 1399 497 1403 501
rect 1455 497 1459 501
rect 1519 497 1523 501
rect 1607 497 1611 501
rect 1695 497 1699 501
rect 1791 497 1795 501
rect 1887 497 1891 501
rect 1983 497 1987 501
rect 2087 497 2091 501
rect 2199 497 2203 501
rect 2311 497 2315 501
rect 2431 497 2435 501
rect 2527 497 2531 501
rect 2583 496 2587 500
rect 111 487 115 491
rect 1327 487 1331 491
rect 159 478 163 482
rect 223 478 227 482
rect 327 478 331 482
rect 447 478 451 482
rect 567 478 571 482
rect 687 478 691 482
rect 807 478 811 482
rect 919 478 923 482
rect 1023 478 1027 482
rect 1119 478 1123 482
rect 1215 478 1219 482
rect 1287 478 1291 482
rect 1367 479 1371 483
rect 2583 479 2587 483
rect 1415 470 1419 474
rect 1471 470 1475 474
rect 1535 470 1539 474
rect 1623 470 1627 474
rect 1711 470 1715 474
rect 1807 470 1811 474
rect 1903 470 1907 474
rect 1999 470 2003 474
rect 2103 470 2107 474
rect 2215 470 2219 474
rect 2327 470 2331 474
rect 2447 470 2451 474
rect 2543 470 2547 474
rect 159 450 163 454
rect 223 450 227 454
rect 319 450 323 454
rect 423 450 427 454
rect 535 450 539 454
rect 639 450 643 454
rect 743 450 747 454
rect 839 450 843 454
rect 927 450 931 454
rect 1007 450 1011 454
rect 1079 450 1083 454
rect 1151 450 1155 454
rect 1231 450 1235 454
rect 1287 450 1291 454
rect 111 441 115 445
rect 1327 441 1331 445
rect 1415 438 1419 442
rect 1487 438 1491 442
rect 1575 438 1579 442
rect 1663 438 1667 442
rect 1759 438 1763 442
rect 1863 438 1867 442
rect 1975 438 1979 442
rect 2111 438 2115 442
rect 2255 438 2259 442
rect 2407 438 2411 442
rect 2543 438 2547 442
rect 1367 429 1371 433
rect 2583 429 2587 433
rect 111 424 115 428
rect 143 423 147 427
rect 207 423 211 427
rect 303 423 307 427
rect 407 423 411 427
rect 519 423 523 427
rect 623 423 627 427
rect 727 423 731 427
rect 823 423 827 427
rect 911 423 915 427
rect 991 423 995 427
rect 1063 423 1067 427
rect 1135 423 1139 427
rect 1215 423 1219 427
rect 1271 423 1275 427
rect 1327 424 1331 428
rect 1367 412 1371 416
rect 1399 411 1403 415
rect 1471 411 1475 415
rect 1559 411 1563 415
rect 1647 411 1651 415
rect 1743 411 1747 415
rect 1847 411 1851 415
rect 1959 411 1963 415
rect 2095 411 2099 415
rect 2239 411 2243 415
rect 2391 411 2395 415
rect 2527 411 2531 415
rect 2583 412 2587 416
rect 111 380 115 384
rect 143 381 147 385
rect 207 381 211 385
rect 303 381 307 385
rect 399 381 403 385
rect 495 381 499 385
rect 583 381 587 385
rect 671 381 675 385
rect 751 381 755 385
rect 823 381 827 385
rect 895 381 899 385
rect 967 381 971 385
rect 1047 381 1051 385
rect 1327 380 1331 384
rect 1367 372 1371 376
rect 1399 373 1403 377
rect 1455 373 1459 377
rect 1511 373 1515 377
rect 1567 373 1571 377
rect 1631 373 1635 377
rect 1695 373 1699 377
rect 1759 373 1763 377
rect 1839 373 1843 377
rect 1943 373 1947 377
rect 2071 373 2075 377
rect 2215 373 2219 377
rect 2367 373 2371 377
rect 2527 373 2531 377
rect 2583 372 2587 376
rect 111 363 115 367
rect 1327 363 1331 367
rect 159 354 163 358
rect 223 354 227 358
rect 319 354 323 358
rect 415 354 419 358
rect 511 354 515 358
rect 599 354 603 358
rect 687 354 691 358
rect 767 354 771 358
rect 839 354 843 358
rect 911 354 915 358
rect 983 354 987 358
rect 1063 354 1067 358
rect 1367 355 1371 359
rect 2583 355 2587 359
rect 1415 346 1419 350
rect 1471 346 1475 350
rect 1527 346 1531 350
rect 1583 346 1587 350
rect 1647 346 1651 350
rect 1711 346 1715 350
rect 1775 346 1779 350
rect 1855 346 1859 350
rect 1959 346 1963 350
rect 2087 346 2091 350
rect 2231 346 2235 350
rect 2383 346 2387 350
rect 2543 346 2547 350
rect 159 326 163 330
rect 223 326 227 330
rect 311 326 315 330
rect 391 326 395 330
rect 471 326 475 330
rect 543 326 547 330
rect 607 326 611 330
rect 671 326 675 330
rect 735 326 739 330
rect 799 326 803 330
rect 863 326 867 330
rect 935 326 939 330
rect 111 317 115 321
rect 1327 317 1331 321
rect 1607 318 1611 322
rect 1663 318 1667 322
rect 1719 318 1723 322
rect 1775 318 1779 322
rect 1831 318 1835 322
rect 1887 318 1891 322
rect 1951 318 1955 322
rect 2031 318 2035 322
rect 2119 318 2123 322
rect 2223 318 2227 322
rect 2335 318 2339 322
rect 2447 318 2451 322
rect 2543 318 2547 322
rect 1367 309 1371 313
rect 2583 309 2587 313
rect 111 300 115 304
rect 143 299 147 303
rect 207 299 211 303
rect 295 299 299 303
rect 375 299 379 303
rect 455 299 459 303
rect 527 299 531 303
rect 591 299 595 303
rect 655 299 659 303
rect 719 299 723 303
rect 783 299 787 303
rect 847 299 851 303
rect 919 299 923 303
rect 1327 300 1331 304
rect 1367 292 1371 296
rect 1591 291 1595 295
rect 1647 291 1651 295
rect 1703 291 1707 295
rect 1759 291 1763 295
rect 1815 291 1819 295
rect 1871 291 1875 295
rect 1935 291 1939 295
rect 2015 291 2019 295
rect 2103 291 2107 295
rect 2207 291 2211 295
rect 2319 291 2323 295
rect 2431 291 2435 295
rect 2527 291 2531 295
rect 2583 292 2587 296
rect 111 256 115 260
rect 143 257 147 261
rect 231 257 235 261
rect 335 257 339 261
rect 431 257 435 261
rect 519 257 523 261
rect 599 257 603 261
rect 679 257 683 261
rect 751 257 755 261
rect 815 257 819 261
rect 887 257 891 261
rect 959 257 963 261
rect 1031 257 1035 261
rect 1327 256 1331 260
rect 1367 252 1371 256
rect 1727 253 1731 257
rect 1783 253 1787 257
rect 1839 253 1843 257
rect 1895 253 1899 257
rect 1951 253 1955 257
rect 2007 253 2011 257
rect 2071 253 2075 257
rect 2143 253 2147 257
rect 2231 253 2235 257
rect 2335 253 2339 257
rect 2439 253 2443 257
rect 2527 253 2531 257
rect 2583 252 2587 256
rect 111 239 115 243
rect 1327 239 1331 243
rect 1367 235 1371 239
rect 159 230 163 234
rect 247 230 251 234
rect 351 230 355 234
rect 447 230 451 234
rect 535 230 539 234
rect 615 230 619 234
rect 695 230 699 234
rect 767 230 771 234
rect 831 230 835 234
rect 903 230 907 234
rect 975 230 979 234
rect 2583 235 2587 239
rect 1047 230 1051 234
rect 1743 226 1747 230
rect 1799 226 1803 230
rect 1855 226 1859 230
rect 1911 226 1915 230
rect 1967 226 1971 230
rect 2023 226 2027 230
rect 2087 226 2091 230
rect 2159 226 2163 230
rect 2247 226 2251 230
rect 2351 226 2355 230
rect 2455 226 2459 230
rect 2543 226 2547 230
rect 167 202 171 206
rect 255 202 259 206
rect 351 202 355 206
rect 447 202 451 206
rect 551 202 555 206
rect 655 202 659 206
rect 751 202 755 206
rect 847 202 851 206
rect 935 202 939 206
rect 1023 202 1027 206
rect 1111 202 1115 206
rect 1199 202 1203 206
rect 1463 202 1467 206
rect 1535 202 1539 206
rect 1623 202 1627 206
rect 1719 202 1723 206
rect 1823 202 1827 206
rect 1927 202 1931 206
rect 2031 202 2035 206
rect 2135 202 2139 206
rect 2239 202 2243 206
rect 2343 202 2347 206
rect 2455 202 2459 206
rect 2543 202 2547 206
rect 111 193 115 197
rect 1327 193 1331 197
rect 1367 193 1371 197
rect 2583 193 2587 197
rect 111 176 115 180
rect 151 175 155 179
rect 239 175 243 179
rect 335 175 339 179
rect 431 175 435 179
rect 535 175 539 179
rect 639 175 643 179
rect 735 175 739 179
rect 831 175 835 179
rect 919 175 923 179
rect 1007 175 1011 179
rect 1095 175 1099 179
rect 1183 175 1187 179
rect 1327 176 1331 180
rect 1367 176 1371 180
rect 1447 175 1451 179
rect 1519 175 1523 179
rect 1607 175 1611 179
rect 1703 175 1707 179
rect 1807 175 1811 179
rect 1911 175 1915 179
rect 2015 175 2019 179
rect 2119 175 2123 179
rect 2223 175 2227 179
rect 2327 175 2331 179
rect 2439 175 2443 179
rect 2527 175 2531 179
rect 2583 176 2587 180
rect 1367 124 1371 128
rect 1399 125 1403 129
rect 1455 125 1459 129
rect 1511 125 1515 129
rect 1567 125 1571 129
rect 1639 125 1643 129
rect 1719 125 1723 129
rect 1799 125 1803 129
rect 1879 125 1883 129
rect 1959 125 1963 129
rect 2031 125 2035 129
rect 2103 125 2107 129
rect 2167 125 2171 129
rect 2231 125 2235 129
rect 2295 125 2299 129
rect 2359 125 2363 129
rect 2415 125 2419 129
rect 2471 125 2475 129
rect 2527 125 2531 129
rect 2583 124 2587 128
rect 111 116 115 120
rect 143 117 147 121
rect 199 117 203 121
rect 255 117 259 121
rect 311 117 315 121
rect 367 117 371 121
rect 423 117 427 121
rect 479 117 483 121
rect 535 117 539 121
rect 607 117 611 121
rect 671 117 675 121
rect 735 117 739 121
rect 799 117 803 121
rect 855 117 859 121
rect 911 117 915 121
rect 975 117 979 121
rect 1039 117 1043 121
rect 1103 117 1107 121
rect 1159 117 1163 121
rect 1215 117 1219 121
rect 1271 117 1275 121
rect 1327 116 1331 120
rect 1367 107 1371 111
rect 2583 107 2587 111
rect 111 99 115 103
rect 1327 99 1331 103
rect 1415 98 1419 102
rect 1471 98 1475 102
rect 1527 98 1531 102
rect 1583 98 1587 102
rect 1655 98 1659 102
rect 1735 98 1739 102
rect 1815 98 1819 102
rect 1895 98 1899 102
rect 1975 98 1979 102
rect 2047 98 2051 102
rect 2119 98 2123 102
rect 2183 98 2187 102
rect 2247 98 2251 102
rect 2311 98 2315 102
rect 2375 98 2379 102
rect 2431 98 2435 102
rect 2487 98 2491 102
rect 2543 98 2547 102
rect 159 90 163 94
rect 215 90 219 94
rect 271 90 275 94
rect 327 90 331 94
rect 383 90 387 94
rect 439 90 443 94
rect 495 90 499 94
rect 551 90 555 94
rect 623 90 627 94
rect 687 90 691 94
rect 751 90 755 94
rect 815 90 819 94
rect 871 90 875 94
rect 927 90 931 94
rect 991 90 995 94
rect 1055 90 1059 94
rect 1119 90 1123 94
rect 1175 90 1179 94
rect 1231 90 1235 94
rect 1287 90 1291 94
<< m3 >>
rect 111 2662 115 2663
rect 111 2657 115 2658
rect 159 2662 163 2663
rect 159 2657 163 2658
rect 215 2662 219 2663
rect 215 2657 219 2658
rect 271 2662 275 2663
rect 271 2657 275 2658
rect 327 2662 331 2663
rect 327 2657 331 2658
rect 1327 2662 1331 2663
rect 1327 2657 1331 2658
rect 112 2642 114 2657
rect 160 2651 162 2657
rect 216 2651 218 2657
rect 272 2651 274 2657
rect 328 2651 330 2657
rect 158 2650 164 2651
rect 158 2646 159 2650
rect 163 2646 164 2650
rect 158 2645 164 2646
rect 214 2650 220 2651
rect 214 2646 215 2650
rect 219 2646 220 2650
rect 214 2645 220 2646
rect 270 2650 276 2651
rect 270 2646 271 2650
rect 275 2646 276 2650
rect 270 2645 276 2646
rect 326 2650 332 2651
rect 326 2646 327 2650
rect 331 2646 332 2650
rect 326 2645 332 2646
rect 1328 2642 1330 2657
rect 110 2641 116 2642
rect 110 2637 111 2641
rect 115 2637 116 2641
rect 110 2636 116 2637
rect 1326 2641 1332 2642
rect 1326 2637 1327 2641
rect 1331 2637 1332 2641
rect 1326 2636 1332 2637
rect 110 2624 116 2625
rect 1326 2624 1332 2625
rect 110 2620 111 2624
rect 115 2620 116 2624
rect 110 2619 116 2620
rect 142 2623 148 2624
rect 142 2619 143 2623
rect 147 2619 148 2623
rect 112 2607 114 2619
rect 142 2618 148 2619
rect 198 2623 204 2624
rect 198 2619 199 2623
rect 203 2619 204 2623
rect 198 2618 204 2619
rect 254 2623 260 2624
rect 254 2619 255 2623
rect 259 2619 260 2623
rect 254 2618 260 2619
rect 310 2623 316 2624
rect 310 2619 311 2623
rect 315 2619 316 2623
rect 1326 2620 1327 2624
rect 1331 2620 1332 2624
rect 1326 2619 1332 2620
rect 310 2618 316 2619
rect 144 2607 146 2618
rect 200 2607 202 2618
rect 256 2607 258 2618
rect 312 2607 314 2618
rect 1328 2607 1330 2619
rect 1367 2610 1371 2611
rect 111 2606 115 2607
rect 111 2601 115 2602
rect 143 2606 147 2607
rect 143 2601 147 2602
rect 199 2606 203 2607
rect 199 2601 203 2602
rect 255 2606 259 2607
rect 255 2601 259 2602
rect 263 2606 267 2607
rect 263 2601 267 2602
rect 311 2606 315 2607
rect 311 2601 315 2602
rect 343 2606 347 2607
rect 343 2601 347 2602
rect 431 2606 435 2607
rect 431 2601 435 2602
rect 519 2606 523 2607
rect 519 2601 523 2602
rect 607 2606 611 2607
rect 607 2601 611 2602
rect 687 2606 691 2607
rect 687 2601 691 2602
rect 767 2606 771 2607
rect 767 2601 771 2602
rect 839 2606 843 2607
rect 839 2601 843 2602
rect 903 2606 907 2607
rect 903 2601 907 2602
rect 967 2606 971 2607
rect 967 2601 971 2602
rect 1031 2606 1035 2607
rect 1031 2601 1035 2602
rect 1095 2606 1099 2607
rect 1095 2601 1099 2602
rect 1159 2606 1163 2607
rect 1159 2601 1163 2602
rect 1215 2606 1219 2607
rect 1215 2601 1219 2602
rect 1271 2606 1275 2607
rect 1271 2601 1275 2602
rect 1327 2606 1331 2607
rect 1367 2605 1371 2606
rect 1415 2610 1419 2611
rect 1415 2605 1419 2606
rect 1471 2610 1475 2611
rect 1471 2605 1475 2606
rect 1527 2610 1531 2611
rect 1527 2605 1531 2606
rect 1583 2610 1587 2611
rect 1583 2605 1587 2606
rect 1639 2610 1643 2611
rect 1639 2605 1643 2606
rect 1695 2610 1699 2611
rect 1695 2605 1699 2606
rect 2583 2610 2587 2611
rect 2583 2605 2587 2606
rect 1327 2601 1331 2602
rect 112 2589 114 2601
rect 144 2590 146 2601
rect 200 2590 202 2601
rect 264 2590 266 2601
rect 344 2590 346 2601
rect 432 2590 434 2601
rect 520 2590 522 2601
rect 608 2590 610 2601
rect 688 2590 690 2601
rect 768 2590 770 2601
rect 840 2590 842 2601
rect 904 2590 906 2601
rect 968 2590 970 2601
rect 1032 2590 1034 2601
rect 1096 2590 1098 2601
rect 1160 2590 1162 2601
rect 1216 2590 1218 2601
rect 1272 2590 1274 2601
rect 142 2589 148 2590
rect 110 2588 116 2589
rect 110 2584 111 2588
rect 115 2584 116 2588
rect 142 2585 143 2589
rect 147 2585 148 2589
rect 142 2584 148 2585
rect 198 2589 204 2590
rect 198 2585 199 2589
rect 203 2585 204 2589
rect 198 2584 204 2585
rect 262 2589 268 2590
rect 262 2585 263 2589
rect 267 2585 268 2589
rect 262 2584 268 2585
rect 342 2589 348 2590
rect 342 2585 343 2589
rect 347 2585 348 2589
rect 342 2584 348 2585
rect 430 2589 436 2590
rect 430 2585 431 2589
rect 435 2585 436 2589
rect 430 2584 436 2585
rect 518 2589 524 2590
rect 518 2585 519 2589
rect 523 2585 524 2589
rect 518 2584 524 2585
rect 606 2589 612 2590
rect 606 2585 607 2589
rect 611 2585 612 2589
rect 606 2584 612 2585
rect 686 2589 692 2590
rect 686 2585 687 2589
rect 691 2585 692 2589
rect 686 2584 692 2585
rect 766 2589 772 2590
rect 766 2585 767 2589
rect 771 2585 772 2589
rect 766 2584 772 2585
rect 838 2589 844 2590
rect 838 2585 839 2589
rect 843 2585 844 2589
rect 838 2584 844 2585
rect 902 2589 908 2590
rect 902 2585 903 2589
rect 907 2585 908 2589
rect 902 2584 908 2585
rect 966 2589 972 2590
rect 966 2585 967 2589
rect 971 2585 972 2589
rect 966 2584 972 2585
rect 1030 2589 1036 2590
rect 1030 2585 1031 2589
rect 1035 2585 1036 2589
rect 1030 2584 1036 2585
rect 1094 2589 1100 2590
rect 1094 2585 1095 2589
rect 1099 2585 1100 2589
rect 1094 2584 1100 2585
rect 1158 2589 1164 2590
rect 1158 2585 1159 2589
rect 1163 2585 1164 2589
rect 1158 2584 1164 2585
rect 1214 2589 1220 2590
rect 1214 2585 1215 2589
rect 1219 2585 1220 2589
rect 1214 2584 1220 2585
rect 1270 2589 1276 2590
rect 1328 2589 1330 2601
rect 1368 2590 1370 2605
rect 1416 2599 1418 2605
rect 1472 2599 1474 2605
rect 1528 2599 1530 2605
rect 1584 2599 1586 2605
rect 1640 2599 1642 2605
rect 1696 2599 1698 2605
rect 1414 2598 1420 2599
rect 1414 2594 1415 2598
rect 1419 2594 1420 2598
rect 1414 2593 1420 2594
rect 1470 2598 1476 2599
rect 1470 2594 1471 2598
rect 1475 2594 1476 2598
rect 1470 2593 1476 2594
rect 1526 2598 1532 2599
rect 1526 2594 1527 2598
rect 1531 2594 1532 2598
rect 1526 2593 1532 2594
rect 1582 2598 1588 2599
rect 1582 2594 1583 2598
rect 1587 2594 1588 2598
rect 1582 2593 1588 2594
rect 1638 2598 1644 2599
rect 1638 2594 1639 2598
rect 1643 2594 1644 2598
rect 1638 2593 1644 2594
rect 1694 2598 1700 2599
rect 1694 2594 1695 2598
rect 1699 2594 1700 2598
rect 1694 2593 1700 2594
rect 2584 2590 2586 2605
rect 1366 2589 1372 2590
rect 1270 2585 1271 2589
rect 1275 2585 1276 2589
rect 1270 2584 1276 2585
rect 1326 2588 1332 2589
rect 1326 2584 1327 2588
rect 1331 2584 1332 2588
rect 1366 2585 1367 2589
rect 1371 2585 1372 2589
rect 1366 2584 1372 2585
rect 2582 2589 2588 2590
rect 2582 2585 2583 2589
rect 2587 2585 2588 2589
rect 2582 2584 2588 2585
rect 110 2583 116 2584
rect 1326 2583 1332 2584
rect 1366 2572 1372 2573
rect 2582 2572 2588 2573
rect 110 2571 116 2572
rect 110 2567 111 2571
rect 115 2567 116 2571
rect 110 2566 116 2567
rect 1326 2571 1332 2572
rect 1326 2567 1327 2571
rect 1331 2567 1332 2571
rect 1366 2568 1367 2572
rect 1371 2568 1372 2572
rect 1366 2567 1372 2568
rect 1398 2571 1404 2572
rect 1398 2567 1399 2571
rect 1403 2567 1404 2571
rect 1326 2566 1332 2567
rect 112 2539 114 2566
rect 158 2562 164 2563
rect 158 2558 159 2562
rect 163 2558 164 2562
rect 158 2557 164 2558
rect 214 2562 220 2563
rect 214 2558 215 2562
rect 219 2558 220 2562
rect 214 2557 220 2558
rect 278 2562 284 2563
rect 278 2558 279 2562
rect 283 2558 284 2562
rect 278 2557 284 2558
rect 358 2562 364 2563
rect 358 2558 359 2562
rect 363 2558 364 2562
rect 358 2557 364 2558
rect 446 2562 452 2563
rect 446 2558 447 2562
rect 451 2558 452 2562
rect 446 2557 452 2558
rect 534 2562 540 2563
rect 534 2558 535 2562
rect 539 2558 540 2562
rect 534 2557 540 2558
rect 622 2562 628 2563
rect 622 2558 623 2562
rect 627 2558 628 2562
rect 622 2557 628 2558
rect 702 2562 708 2563
rect 702 2558 703 2562
rect 707 2558 708 2562
rect 702 2557 708 2558
rect 782 2562 788 2563
rect 782 2558 783 2562
rect 787 2558 788 2562
rect 782 2557 788 2558
rect 854 2562 860 2563
rect 854 2558 855 2562
rect 859 2558 860 2562
rect 854 2557 860 2558
rect 918 2562 924 2563
rect 918 2558 919 2562
rect 923 2558 924 2562
rect 918 2557 924 2558
rect 982 2562 988 2563
rect 982 2558 983 2562
rect 987 2558 988 2562
rect 982 2557 988 2558
rect 1046 2562 1052 2563
rect 1046 2558 1047 2562
rect 1051 2558 1052 2562
rect 1046 2557 1052 2558
rect 1110 2562 1116 2563
rect 1110 2558 1111 2562
rect 1115 2558 1116 2562
rect 1110 2557 1116 2558
rect 1174 2562 1180 2563
rect 1174 2558 1175 2562
rect 1179 2558 1180 2562
rect 1174 2557 1180 2558
rect 1230 2562 1236 2563
rect 1230 2558 1231 2562
rect 1235 2558 1236 2562
rect 1230 2557 1236 2558
rect 1286 2562 1292 2563
rect 1286 2558 1287 2562
rect 1291 2558 1292 2562
rect 1286 2557 1292 2558
rect 160 2539 162 2557
rect 216 2539 218 2557
rect 280 2539 282 2557
rect 360 2539 362 2557
rect 448 2539 450 2557
rect 536 2539 538 2557
rect 624 2539 626 2557
rect 704 2539 706 2557
rect 784 2539 786 2557
rect 856 2539 858 2557
rect 920 2539 922 2557
rect 984 2539 986 2557
rect 1048 2539 1050 2557
rect 1112 2539 1114 2557
rect 1176 2539 1178 2557
rect 1232 2539 1234 2557
rect 1288 2539 1290 2557
rect 1328 2539 1330 2566
rect 1368 2555 1370 2567
rect 1398 2566 1404 2567
rect 1454 2571 1460 2572
rect 1454 2567 1455 2571
rect 1459 2567 1460 2571
rect 1454 2566 1460 2567
rect 1510 2571 1516 2572
rect 1510 2567 1511 2571
rect 1515 2567 1516 2571
rect 1510 2566 1516 2567
rect 1566 2571 1572 2572
rect 1566 2567 1567 2571
rect 1571 2567 1572 2571
rect 1566 2566 1572 2567
rect 1622 2571 1628 2572
rect 1622 2567 1623 2571
rect 1627 2567 1628 2571
rect 1622 2566 1628 2567
rect 1678 2571 1684 2572
rect 1678 2567 1679 2571
rect 1683 2567 1684 2571
rect 2582 2568 2583 2572
rect 2587 2568 2588 2572
rect 2582 2567 2588 2568
rect 1678 2566 1684 2567
rect 1400 2555 1402 2566
rect 1456 2555 1458 2566
rect 1512 2555 1514 2566
rect 1568 2555 1570 2566
rect 1624 2555 1626 2566
rect 1680 2555 1682 2566
rect 2584 2555 2586 2567
rect 1367 2554 1371 2555
rect 1367 2549 1371 2550
rect 1399 2554 1403 2555
rect 1399 2549 1403 2550
rect 1455 2554 1459 2555
rect 1455 2549 1459 2550
rect 1511 2554 1515 2555
rect 1511 2549 1515 2550
rect 1567 2554 1571 2555
rect 1567 2549 1571 2550
rect 1623 2554 1627 2555
rect 1623 2549 1627 2550
rect 1679 2554 1683 2555
rect 1679 2549 1683 2550
rect 1735 2554 1739 2555
rect 1735 2549 1739 2550
rect 2583 2554 2587 2555
rect 2583 2549 2587 2550
rect 111 2538 115 2539
rect 111 2533 115 2534
rect 159 2538 163 2539
rect 159 2533 163 2534
rect 215 2538 219 2539
rect 215 2533 219 2534
rect 279 2538 283 2539
rect 279 2533 283 2534
rect 319 2538 323 2539
rect 319 2533 323 2534
rect 359 2538 363 2539
rect 359 2533 363 2534
rect 431 2538 435 2539
rect 431 2533 435 2534
rect 447 2538 451 2539
rect 447 2533 451 2534
rect 535 2538 539 2539
rect 535 2533 539 2534
rect 551 2538 555 2539
rect 551 2533 555 2534
rect 623 2538 627 2539
rect 623 2533 627 2534
rect 671 2538 675 2539
rect 671 2533 675 2534
rect 703 2538 707 2539
rect 703 2533 707 2534
rect 783 2538 787 2539
rect 783 2533 787 2534
rect 791 2538 795 2539
rect 791 2533 795 2534
rect 855 2538 859 2539
rect 855 2533 859 2534
rect 903 2538 907 2539
rect 903 2533 907 2534
rect 919 2538 923 2539
rect 919 2533 923 2534
rect 983 2538 987 2539
rect 983 2533 987 2534
rect 1007 2538 1011 2539
rect 1007 2533 1011 2534
rect 1047 2538 1051 2539
rect 1047 2533 1051 2534
rect 1103 2538 1107 2539
rect 1103 2533 1107 2534
rect 1111 2538 1115 2539
rect 1111 2533 1115 2534
rect 1175 2538 1179 2539
rect 1175 2533 1179 2534
rect 1207 2538 1211 2539
rect 1207 2533 1211 2534
rect 1231 2538 1235 2539
rect 1231 2533 1235 2534
rect 1287 2538 1291 2539
rect 1287 2533 1291 2534
rect 1327 2538 1331 2539
rect 1368 2537 1370 2549
rect 1400 2538 1402 2549
rect 1456 2538 1458 2549
rect 1512 2538 1514 2549
rect 1568 2538 1570 2549
rect 1624 2538 1626 2549
rect 1680 2538 1682 2549
rect 1736 2538 1738 2549
rect 1398 2537 1404 2538
rect 1327 2533 1331 2534
rect 1366 2536 1372 2537
rect 112 2518 114 2533
rect 160 2527 162 2533
rect 216 2527 218 2533
rect 320 2527 322 2533
rect 432 2527 434 2533
rect 552 2527 554 2533
rect 672 2527 674 2533
rect 792 2527 794 2533
rect 904 2527 906 2533
rect 1008 2527 1010 2533
rect 1104 2527 1106 2533
rect 1208 2527 1210 2533
rect 1288 2527 1290 2533
rect 158 2526 164 2527
rect 158 2522 159 2526
rect 163 2522 164 2526
rect 158 2521 164 2522
rect 214 2526 220 2527
rect 214 2522 215 2526
rect 219 2522 220 2526
rect 214 2521 220 2522
rect 318 2526 324 2527
rect 318 2522 319 2526
rect 323 2522 324 2526
rect 318 2521 324 2522
rect 430 2526 436 2527
rect 430 2522 431 2526
rect 435 2522 436 2526
rect 430 2521 436 2522
rect 550 2526 556 2527
rect 550 2522 551 2526
rect 555 2522 556 2526
rect 550 2521 556 2522
rect 670 2526 676 2527
rect 670 2522 671 2526
rect 675 2522 676 2526
rect 670 2521 676 2522
rect 790 2526 796 2527
rect 790 2522 791 2526
rect 795 2522 796 2526
rect 790 2521 796 2522
rect 902 2526 908 2527
rect 902 2522 903 2526
rect 907 2522 908 2526
rect 902 2521 908 2522
rect 1006 2526 1012 2527
rect 1006 2522 1007 2526
rect 1011 2522 1012 2526
rect 1006 2521 1012 2522
rect 1102 2526 1108 2527
rect 1102 2522 1103 2526
rect 1107 2522 1108 2526
rect 1102 2521 1108 2522
rect 1206 2526 1212 2527
rect 1206 2522 1207 2526
rect 1211 2522 1212 2526
rect 1206 2521 1212 2522
rect 1286 2526 1292 2527
rect 1286 2522 1287 2526
rect 1291 2522 1292 2526
rect 1286 2521 1292 2522
rect 1328 2518 1330 2533
rect 1366 2532 1367 2536
rect 1371 2532 1372 2536
rect 1398 2533 1399 2537
rect 1403 2533 1404 2537
rect 1398 2532 1404 2533
rect 1454 2537 1460 2538
rect 1454 2533 1455 2537
rect 1459 2533 1460 2537
rect 1454 2532 1460 2533
rect 1510 2537 1516 2538
rect 1510 2533 1511 2537
rect 1515 2533 1516 2537
rect 1510 2532 1516 2533
rect 1566 2537 1572 2538
rect 1566 2533 1567 2537
rect 1571 2533 1572 2537
rect 1566 2532 1572 2533
rect 1622 2537 1628 2538
rect 1622 2533 1623 2537
rect 1627 2533 1628 2537
rect 1622 2532 1628 2533
rect 1678 2537 1684 2538
rect 1678 2533 1679 2537
rect 1683 2533 1684 2537
rect 1678 2532 1684 2533
rect 1734 2537 1740 2538
rect 2584 2537 2586 2549
rect 1734 2533 1735 2537
rect 1739 2533 1740 2537
rect 1734 2532 1740 2533
rect 2582 2536 2588 2537
rect 2582 2532 2583 2536
rect 2587 2532 2588 2536
rect 1366 2531 1372 2532
rect 2582 2531 2588 2532
rect 1366 2519 1372 2520
rect 110 2517 116 2518
rect 110 2513 111 2517
rect 115 2513 116 2517
rect 110 2512 116 2513
rect 1326 2517 1332 2518
rect 1326 2513 1327 2517
rect 1331 2513 1332 2517
rect 1366 2515 1367 2519
rect 1371 2515 1372 2519
rect 1366 2514 1372 2515
rect 2582 2519 2588 2520
rect 2582 2515 2583 2519
rect 2587 2515 2588 2519
rect 2582 2514 2588 2515
rect 1326 2512 1332 2513
rect 110 2500 116 2501
rect 1326 2500 1332 2501
rect 110 2496 111 2500
rect 115 2496 116 2500
rect 110 2495 116 2496
rect 142 2499 148 2500
rect 142 2495 143 2499
rect 147 2495 148 2499
rect 112 2475 114 2495
rect 142 2494 148 2495
rect 198 2499 204 2500
rect 198 2495 199 2499
rect 203 2495 204 2499
rect 198 2494 204 2495
rect 302 2499 308 2500
rect 302 2495 303 2499
rect 307 2495 308 2499
rect 302 2494 308 2495
rect 414 2499 420 2500
rect 414 2495 415 2499
rect 419 2495 420 2499
rect 414 2494 420 2495
rect 534 2499 540 2500
rect 534 2495 535 2499
rect 539 2495 540 2499
rect 534 2494 540 2495
rect 654 2499 660 2500
rect 654 2495 655 2499
rect 659 2495 660 2499
rect 654 2494 660 2495
rect 774 2499 780 2500
rect 774 2495 775 2499
rect 779 2495 780 2499
rect 774 2494 780 2495
rect 886 2499 892 2500
rect 886 2495 887 2499
rect 891 2495 892 2499
rect 886 2494 892 2495
rect 990 2499 996 2500
rect 990 2495 991 2499
rect 995 2495 996 2499
rect 990 2494 996 2495
rect 1086 2499 1092 2500
rect 1086 2495 1087 2499
rect 1091 2495 1092 2499
rect 1086 2494 1092 2495
rect 1190 2499 1196 2500
rect 1190 2495 1191 2499
rect 1195 2495 1196 2499
rect 1190 2494 1196 2495
rect 1270 2499 1276 2500
rect 1270 2495 1271 2499
rect 1275 2495 1276 2499
rect 1326 2496 1327 2500
rect 1331 2496 1332 2500
rect 1326 2495 1332 2496
rect 1368 2495 1370 2514
rect 1414 2510 1420 2511
rect 1414 2506 1415 2510
rect 1419 2506 1420 2510
rect 1414 2505 1420 2506
rect 1470 2510 1476 2511
rect 1470 2506 1471 2510
rect 1475 2506 1476 2510
rect 1470 2505 1476 2506
rect 1526 2510 1532 2511
rect 1526 2506 1527 2510
rect 1531 2506 1532 2510
rect 1526 2505 1532 2506
rect 1582 2510 1588 2511
rect 1582 2506 1583 2510
rect 1587 2506 1588 2510
rect 1582 2505 1588 2506
rect 1638 2510 1644 2511
rect 1638 2506 1639 2510
rect 1643 2506 1644 2510
rect 1638 2505 1644 2506
rect 1694 2510 1700 2511
rect 1694 2506 1695 2510
rect 1699 2506 1700 2510
rect 1694 2505 1700 2506
rect 1750 2510 1756 2511
rect 1750 2506 1751 2510
rect 1755 2506 1756 2510
rect 1750 2505 1756 2506
rect 1416 2495 1418 2505
rect 1472 2495 1474 2505
rect 1528 2495 1530 2505
rect 1584 2495 1586 2505
rect 1640 2495 1642 2505
rect 1696 2495 1698 2505
rect 1752 2495 1754 2505
rect 2584 2495 2586 2514
rect 1270 2494 1276 2495
rect 144 2475 146 2494
rect 200 2475 202 2494
rect 304 2475 306 2494
rect 416 2475 418 2494
rect 536 2475 538 2494
rect 656 2475 658 2494
rect 776 2475 778 2494
rect 888 2475 890 2494
rect 992 2475 994 2494
rect 1088 2475 1090 2494
rect 1192 2475 1194 2494
rect 1272 2475 1274 2494
rect 1328 2475 1330 2495
rect 1367 2494 1371 2495
rect 1367 2489 1371 2490
rect 1415 2494 1419 2495
rect 1415 2489 1419 2490
rect 1471 2494 1475 2495
rect 1471 2489 1475 2490
rect 1527 2494 1531 2495
rect 1527 2489 1531 2490
rect 1583 2494 1587 2495
rect 1583 2489 1587 2490
rect 1639 2494 1643 2495
rect 1639 2489 1643 2490
rect 1695 2494 1699 2495
rect 1695 2489 1699 2490
rect 1751 2494 1755 2495
rect 1751 2489 1755 2490
rect 2583 2494 2587 2495
rect 2583 2489 2587 2490
rect 111 2474 115 2475
rect 111 2469 115 2470
rect 143 2474 147 2475
rect 143 2469 147 2470
rect 199 2474 203 2475
rect 199 2469 203 2470
rect 295 2474 299 2475
rect 295 2469 299 2470
rect 303 2474 307 2475
rect 303 2469 307 2470
rect 407 2474 411 2475
rect 407 2469 411 2470
rect 415 2474 419 2475
rect 415 2469 419 2470
rect 519 2474 523 2475
rect 519 2469 523 2470
rect 535 2474 539 2475
rect 535 2469 539 2470
rect 639 2474 643 2475
rect 639 2469 643 2470
rect 655 2474 659 2475
rect 655 2469 659 2470
rect 751 2474 755 2475
rect 751 2469 755 2470
rect 775 2474 779 2475
rect 775 2469 779 2470
rect 855 2474 859 2475
rect 855 2469 859 2470
rect 887 2474 891 2475
rect 887 2469 891 2470
rect 951 2474 955 2475
rect 951 2469 955 2470
rect 991 2474 995 2475
rect 991 2469 995 2470
rect 1047 2474 1051 2475
rect 1047 2469 1051 2470
rect 1087 2474 1091 2475
rect 1087 2469 1091 2470
rect 1143 2474 1147 2475
rect 1143 2469 1147 2470
rect 1191 2474 1195 2475
rect 1191 2469 1195 2470
rect 1239 2474 1243 2475
rect 1239 2469 1243 2470
rect 1271 2474 1275 2475
rect 1271 2469 1275 2470
rect 1327 2474 1331 2475
rect 1368 2474 1370 2489
rect 1472 2483 1474 2489
rect 1528 2483 1530 2489
rect 1584 2483 1586 2489
rect 1640 2483 1642 2489
rect 1696 2483 1698 2489
rect 1752 2483 1754 2489
rect 1470 2482 1476 2483
rect 1470 2478 1471 2482
rect 1475 2478 1476 2482
rect 1470 2477 1476 2478
rect 1526 2482 1532 2483
rect 1526 2478 1527 2482
rect 1531 2478 1532 2482
rect 1526 2477 1532 2478
rect 1582 2482 1588 2483
rect 1582 2478 1583 2482
rect 1587 2478 1588 2482
rect 1582 2477 1588 2478
rect 1638 2482 1644 2483
rect 1638 2478 1639 2482
rect 1643 2478 1644 2482
rect 1638 2477 1644 2478
rect 1694 2482 1700 2483
rect 1694 2478 1695 2482
rect 1699 2478 1700 2482
rect 1694 2477 1700 2478
rect 1750 2482 1756 2483
rect 1750 2478 1751 2482
rect 1755 2478 1756 2482
rect 1750 2477 1756 2478
rect 2584 2474 2586 2489
rect 1327 2469 1331 2470
rect 1366 2473 1372 2474
rect 1366 2469 1367 2473
rect 1371 2469 1372 2473
rect 112 2457 114 2469
rect 144 2458 146 2469
rect 200 2458 202 2469
rect 296 2458 298 2469
rect 408 2458 410 2469
rect 520 2458 522 2469
rect 640 2458 642 2469
rect 752 2458 754 2469
rect 856 2458 858 2469
rect 952 2458 954 2469
rect 1048 2458 1050 2469
rect 1144 2458 1146 2469
rect 1240 2458 1242 2469
rect 142 2457 148 2458
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 142 2453 143 2457
rect 147 2453 148 2457
rect 142 2452 148 2453
rect 198 2457 204 2458
rect 198 2453 199 2457
rect 203 2453 204 2457
rect 198 2452 204 2453
rect 294 2457 300 2458
rect 294 2453 295 2457
rect 299 2453 300 2457
rect 294 2452 300 2453
rect 406 2457 412 2458
rect 406 2453 407 2457
rect 411 2453 412 2457
rect 406 2452 412 2453
rect 518 2457 524 2458
rect 518 2453 519 2457
rect 523 2453 524 2457
rect 518 2452 524 2453
rect 638 2457 644 2458
rect 638 2453 639 2457
rect 643 2453 644 2457
rect 638 2452 644 2453
rect 750 2457 756 2458
rect 750 2453 751 2457
rect 755 2453 756 2457
rect 750 2452 756 2453
rect 854 2457 860 2458
rect 854 2453 855 2457
rect 859 2453 860 2457
rect 854 2452 860 2453
rect 950 2457 956 2458
rect 950 2453 951 2457
rect 955 2453 956 2457
rect 950 2452 956 2453
rect 1046 2457 1052 2458
rect 1046 2453 1047 2457
rect 1051 2453 1052 2457
rect 1046 2452 1052 2453
rect 1142 2457 1148 2458
rect 1142 2453 1143 2457
rect 1147 2453 1148 2457
rect 1142 2452 1148 2453
rect 1238 2457 1244 2458
rect 1328 2457 1330 2469
rect 1366 2468 1372 2469
rect 2582 2473 2588 2474
rect 2582 2469 2583 2473
rect 2587 2469 2588 2473
rect 2582 2468 2588 2469
rect 1238 2453 1239 2457
rect 1243 2453 1244 2457
rect 1238 2452 1244 2453
rect 1326 2456 1332 2457
rect 1326 2452 1327 2456
rect 1331 2452 1332 2456
rect 110 2451 116 2452
rect 1326 2451 1332 2452
rect 1366 2456 1372 2457
rect 2582 2456 2588 2457
rect 1366 2452 1367 2456
rect 1371 2452 1372 2456
rect 1366 2451 1372 2452
rect 1454 2455 1460 2456
rect 1454 2451 1455 2455
rect 1459 2451 1460 2455
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 1326 2439 1332 2440
rect 1326 2435 1327 2439
rect 1331 2435 1332 2439
rect 1326 2434 1332 2435
rect 112 2411 114 2434
rect 158 2430 164 2431
rect 158 2426 159 2430
rect 163 2426 164 2430
rect 158 2425 164 2426
rect 214 2430 220 2431
rect 214 2426 215 2430
rect 219 2426 220 2430
rect 214 2425 220 2426
rect 310 2430 316 2431
rect 310 2426 311 2430
rect 315 2426 316 2430
rect 310 2425 316 2426
rect 422 2430 428 2431
rect 422 2426 423 2430
rect 427 2426 428 2430
rect 422 2425 428 2426
rect 534 2430 540 2431
rect 534 2426 535 2430
rect 539 2426 540 2430
rect 534 2425 540 2426
rect 654 2430 660 2431
rect 654 2426 655 2430
rect 659 2426 660 2430
rect 654 2425 660 2426
rect 766 2430 772 2431
rect 766 2426 767 2430
rect 771 2426 772 2430
rect 766 2425 772 2426
rect 870 2430 876 2431
rect 870 2426 871 2430
rect 875 2426 876 2430
rect 870 2425 876 2426
rect 966 2430 972 2431
rect 966 2426 967 2430
rect 971 2426 972 2430
rect 966 2425 972 2426
rect 1062 2430 1068 2431
rect 1062 2426 1063 2430
rect 1067 2426 1068 2430
rect 1062 2425 1068 2426
rect 1158 2430 1164 2431
rect 1158 2426 1159 2430
rect 1163 2426 1164 2430
rect 1158 2425 1164 2426
rect 1254 2430 1260 2431
rect 1254 2426 1255 2430
rect 1259 2426 1260 2430
rect 1254 2425 1260 2426
rect 160 2411 162 2425
rect 216 2411 218 2425
rect 312 2411 314 2425
rect 424 2411 426 2425
rect 536 2411 538 2425
rect 656 2411 658 2425
rect 768 2411 770 2425
rect 872 2411 874 2425
rect 968 2411 970 2425
rect 1064 2411 1066 2425
rect 1160 2411 1162 2425
rect 1256 2411 1258 2425
rect 1328 2411 1330 2434
rect 1368 2431 1370 2451
rect 1454 2450 1460 2451
rect 1510 2455 1516 2456
rect 1510 2451 1511 2455
rect 1515 2451 1516 2455
rect 1510 2450 1516 2451
rect 1566 2455 1572 2456
rect 1566 2451 1567 2455
rect 1571 2451 1572 2455
rect 1566 2450 1572 2451
rect 1622 2455 1628 2456
rect 1622 2451 1623 2455
rect 1627 2451 1628 2455
rect 1622 2450 1628 2451
rect 1678 2455 1684 2456
rect 1678 2451 1679 2455
rect 1683 2451 1684 2455
rect 1678 2450 1684 2451
rect 1734 2455 1740 2456
rect 1734 2451 1735 2455
rect 1739 2451 1740 2455
rect 2582 2452 2583 2456
rect 2587 2452 2588 2456
rect 2582 2451 2588 2452
rect 1734 2450 1740 2451
rect 1456 2431 1458 2450
rect 1512 2431 1514 2450
rect 1568 2431 1570 2450
rect 1624 2431 1626 2450
rect 1680 2431 1682 2450
rect 1736 2431 1738 2450
rect 2584 2431 2586 2451
rect 1367 2430 1371 2431
rect 1367 2425 1371 2426
rect 1455 2430 1459 2431
rect 1455 2425 1459 2426
rect 1479 2430 1483 2431
rect 1479 2425 1483 2426
rect 1511 2430 1515 2431
rect 1511 2425 1515 2426
rect 1535 2430 1539 2431
rect 1535 2425 1539 2426
rect 1567 2430 1571 2431
rect 1567 2425 1571 2426
rect 1591 2430 1595 2431
rect 1591 2425 1595 2426
rect 1623 2430 1627 2431
rect 1623 2425 1627 2426
rect 1647 2430 1651 2431
rect 1647 2425 1651 2426
rect 1679 2430 1683 2431
rect 1679 2425 1683 2426
rect 1703 2430 1707 2431
rect 1703 2425 1707 2426
rect 1735 2430 1739 2431
rect 1735 2425 1739 2426
rect 1759 2430 1763 2431
rect 1759 2425 1763 2426
rect 2583 2430 2587 2431
rect 2583 2425 2587 2426
rect 1368 2413 1370 2425
rect 1480 2414 1482 2425
rect 1536 2414 1538 2425
rect 1592 2414 1594 2425
rect 1648 2414 1650 2425
rect 1704 2414 1706 2425
rect 1760 2414 1762 2425
rect 1478 2413 1484 2414
rect 1366 2412 1372 2413
rect 111 2410 115 2411
rect 111 2405 115 2406
rect 159 2410 163 2411
rect 159 2405 163 2406
rect 215 2410 219 2411
rect 215 2405 219 2406
rect 223 2410 227 2411
rect 223 2405 227 2406
rect 287 2410 291 2411
rect 287 2405 291 2406
rect 311 2410 315 2411
rect 311 2405 315 2406
rect 367 2410 371 2411
rect 367 2405 371 2406
rect 423 2410 427 2411
rect 423 2405 427 2406
rect 455 2410 459 2411
rect 455 2405 459 2406
rect 535 2410 539 2411
rect 535 2405 539 2406
rect 543 2410 547 2411
rect 543 2405 547 2406
rect 639 2410 643 2411
rect 639 2405 643 2406
rect 655 2410 659 2411
rect 655 2405 659 2406
rect 727 2410 731 2411
rect 727 2405 731 2406
rect 767 2410 771 2411
rect 767 2405 771 2406
rect 815 2410 819 2411
rect 815 2405 819 2406
rect 871 2410 875 2411
rect 871 2405 875 2406
rect 895 2410 899 2411
rect 895 2405 899 2406
rect 967 2410 971 2411
rect 967 2405 971 2406
rect 975 2410 979 2411
rect 975 2405 979 2406
rect 1055 2410 1059 2411
rect 1055 2405 1059 2406
rect 1063 2410 1067 2411
rect 1063 2405 1067 2406
rect 1143 2410 1147 2411
rect 1143 2405 1147 2406
rect 1159 2410 1163 2411
rect 1159 2405 1163 2406
rect 1255 2410 1259 2411
rect 1255 2405 1259 2406
rect 1327 2410 1331 2411
rect 1366 2408 1367 2412
rect 1371 2408 1372 2412
rect 1478 2409 1479 2413
rect 1483 2409 1484 2413
rect 1478 2408 1484 2409
rect 1534 2413 1540 2414
rect 1534 2409 1535 2413
rect 1539 2409 1540 2413
rect 1534 2408 1540 2409
rect 1590 2413 1596 2414
rect 1590 2409 1591 2413
rect 1595 2409 1596 2413
rect 1590 2408 1596 2409
rect 1646 2413 1652 2414
rect 1646 2409 1647 2413
rect 1651 2409 1652 2413
rect 1646 2408 1652 2409
rect 1702 2413 1708 2414
rect 1702 2409 1703 2413
rect 1707 2409 1708 2413
rect 1702 2408 1708 2409
rect 1758 2413 1764 2414
rect 2584 2413 2586 2425
rect 1758 2409 1759 2413
rect 1763 2409 1764 2413
rect 1758 2408 1764 2409
rect 2582 2412 2588 2413
rect 2582 2408 2583 2412
rect 2587 2408 2588 2412
rect 1366 2407 1372 2408
rect 2582 2407 2588 2408
rect 1327 2405 1331 2406
rect 112 2390 114 2405
rect 224 2399 226 2405
rect 288 2399 290 2405
rect 368 2399 370 2405
rect 456 2399 458 2405
rect 544 2399 546 2405
rect 640 2399 642 2405
rect 728 2399 730 2405
rect 816 2399 818 2405
rect 896 2399 898 2405
rect 976 2399 978 2405
rect 1056 2399 1058 2405
rect 1144 2399 1146 2405
rect 222 2398 228 2399
rect 222 2394 223 2398
rect 227 2394 228 2398
rect 222 2393 228 2394
rect 286 2398 292 2399
rect 286 2394 287 2398
rect 291 2394 292 2398
rect 286 2393 292 2394
rect 366 2398 372 2399
rect 366 2394 367 2398
rect 371 2394 372 2398
rect 366 2393 372 2394
rect 454 2398 460 2399
rect 454 2394 455 2398
rect 459 2394 460 2398
rect 454 2393 460 2394
rect 542 2398 548 2399
rect 542 2394 543 2398
rect 547 2394 548 2398
rect 542 2393 548 2394
rect 638 2398 644 2399
rect 638 2394 639 2398
rect 643 2394 644 2398
rect 638 2393 644 2394
rect 726 2398 732 2399
rect 726 2394 727 2398
rect 731 2394 732 2398
rect 726 2393 732 2394
rect 814 2398 820 2399
rect 814 2394 815 2398
rect 819 2394 820 2398
rect 814 2393 820 2394
rect 894 2398 900 2399
rect 894 2394 895 2398
rect 899 2394 900 2398
rect 894 2393 900 2394
rect 974 2398 980 2399
rect 974 2394 975 2398
rect 979 2394 980 2398
rect 974 2393 980 2394
rect 1054 2398 1060 2399
rect 1054 2394 1055 2398
rect 1059 2394 1060 2398
rect 1054 2393 1060 2394
rect 1142 2398 1148 2399
rect 1142 2394 1143 2398
rect 1147 2394 1148 2398
rect 1142 2393 1148 2394
rect 1328 2390 1330 2405
rect 1366 2395 1372 2396
rect 1366 2391 1367 2395
rect 1371 2391 1372 2395
rect 1366 2390 1372 2391
rect 2582 2395 2588 2396
rect 2582 2391 2583 2395
rect 2587 2391 2588 2395
rect 2582 2390 2588 2391
rect 110 2389 116 2390
rect 110 2385 111 2389
rect 115 2385 116 2389
rect 110 2384 116 2385
rect 1326 2389 1332 2390
rect 1326 2385 1327 2389
rect 1331 2385 1332 2389
rect 1326 2384 1332 2385
rect 110 2372 116 2373
rect 1326 2372 1332 2373
rect 110 2368 111 2372
rect 115 2368 116 2372
rect 110 2367 116 2368
rect 206 2371 212 2372
rect 206 2367 207 2371
rect 211 2367 212 2371
rect 112 2347 114 2367
rect 206 2366 212 2367
rect 270 2371 276 2372
rect 270 2367 271 2371
rect 275 2367 276 2371
rect 270 2366 276 2367
rect 350 2371 356 2372
rect 350 2367 351 2371
rect 355 2367 356 2371
rect 350 2366 356 2367
rect 438 2371 444 2372
rect 438 2367 439 2371
rect 443 2367 444 2371
rect 438 2366 444 2367
rect 526 2371 532 2372
rect 526 2367 527 2371
rect 531 2367 532 2371
rect 526 2366 532 2367
rect 622 2371 628 2372
rect 622 2367 623 2371
rect 627 2367 628 2371
rect 622 2366 628 2367
rect 710 2371 716 2372
rect 710 2367 711 2371
rect 715 2367 716 2371
rect 710 2366 716 2367
rect 798 2371 804 2372
rect 798 2367 799 2371
rect 803 2367 804 2371
rect 798 2366 804 2367
rect 878 2371 884 2372
rect 878 2367 879 2371
rect 883 2367 884 2371
rect 878 2366 884 2367
rect 958 2371 964 2372
rect 958 2367 959 2371
rect 963 2367 964 2371
rect 958 2366 964 2367
rect 1038 2371 1044 2372
rect 1038 2367 1039 2371
rect 1043 2367 1044 2371
rect 1038 2366 1044 2367
rect 1126 2371 1132 2372
rect 1126 2367 1127 2371
rect 1131 2367 1132 2371
rect 1326 2368 1327 2372
rect 1331 2368 1332 2372
rect 1368 2371 1370 2390
rect 1494 2386 1500 2387
rect 1494 2382 1495 2386
rect 1499 2382 1500 2386
rect 1494 2381 1500 2382
rect 1550 2386 1556 2387
rect 1550 2382 1551 2386
rect 1555 2382 1556 2386
rect 1550 2381 1556 2382
rect 1606 2386 1612 2387
rect 1606 2382 1607 2386
rect 1611 2382 1612 2386
rect 1606 2381 1612 2382
rect 1662 2386 1668 2387
rect 1662 2382 1663 2386
rect 1667 2382 1668 2386
rect 1662 2381 1668 2382
rect 1718 2386 1724 2387
rect 1718 2382 1719 2386
rect 1723 2382 1724 2386
rect 1718 2381 1724 2382
rect 1774 2386 1780 2387
rect 1774 2382 1775 2386
rect 1779 2382 1780 2386
rect 1774 2381 1780 2382
rect 1496 2371 1498 2381
rect 1552 2371 1554 2381
rect 1608 2371 1610 2381
rect 1664 2371 1666 2381
rect 1720 2371 1722 2381
rect 1776 2371 1778 2381
rect 2584 2371 2586 2390
rect 1326 2367 1332 2368
rect 1367 2370 1371 2371
rect 1126 2366 1132 2367
rect 208 2347 210 2366
rect 272 2347 274 2366
rect 352 2347 354 2366
rect 440 2347 442 2366
rect 528 2347 530 2366
rect 624 2347 626 2366
rect 712 2347 714 2366
rect 800 2347 802 2366
rect 880 2347 882 2366
rect 960 2347 962 2366
rect 1040 2347 1042 2366
rect 1128 2347 1130 2366
rect 1328 2347 1330 2367
rect 1367 2365 1371 2366
rect 1471 2370 1475 2371
rect 1471 2365 1475 2366
rect 1495 2370 1499 2371
rect 1495 2365 1499 2366
rect 1527 2370 1531 2371
rect 1527 2365 1531 2366
rect 1551 2370 1555 2371
rect 1551 2365 1555 2366
rect 1583 2370 1587 2371
rect 1583 2365 1587 2366
rect 1607 2370 1611 2371
rect 1607 2365 1611 2366
rect 1639 2370 1643 2371
rect 1639 2365 1643 2366
rect 1663 2370 1667 2371
rect 1663 2365 1667 2366
rect 1695 2370 1699 2371
rect 1695 2365 1699 2366
rect 1719 2370 1723 2371
rect 1719 2365 1723 2366
rect 1775 2370 1779 2371
rect 1775 2365 1779 2366
rect 2583 2370 2587 2371
rect 2583 2365 2587 2366
rect 1368 2350 1370 2365
rect 1472 2359 1474 2365
rect 1528 2359 1530 2365
rect 1584 2359 1586 2365
rect 1640 2359 1642 2365
rect 1696 2359 1698 2365
rect 1470 2358 1476 2359
rect 1470 2354 1471 2358
rect 1475 2354 1476 2358
rect 1470 2353 1476 2354
rect 1526 2358 1532 2359
rect 1526 2354 1527 2358
rect 1531 2354 1532 2358
rect 1526 2353 1532 2354
rect 1582 2358 1588 2359
rect 1582 2354 1583 2358
rect 1587 2354 1588 2358
rect 1582 2353 1588 2354
rect 1638 2358 1644 2359
rect 1638 2354 1639 2358
rect 1643 2354 1644 2358
rect 1638 2353 1644 2354
rect 1694 2358 1700 2359
rect 1694 2354 1695 2358
rect 1699 2354 1700 2358
rect 1694 2353 1700 2354
rect 2584 2350 2586 2365
rect 1366 2349 1372 2350
rect 111 2346 115 2347
rect 111 2341 115 2342
rect 207 2346 211 2347
rect 207 2341 211 2342
rect 271 2346 275 2347
rect 271 2341 275 2342
rect 327 2346 331 2347
rect 327 2341 331 2342
rect 351 2346 355 2347
rect 351 2341 355 2342
rect 383 2346 387 2347
rect 383 2341 387 2342
rect 439 2346 443 2347
rect 439 2341 443 2342
rect 503 2346 507 2347
rect 503 2341 507 2342
rect 527 2346 531 2347
rect 527 2341 531 2342
rect 567 2346 571 2347
rect 567 2341 571 2342
rect 623 2346 627 2347
rect 623 2341 627 2342
rect 631 2346 635 2347
rect 631 2341 635 2342
rect 695 2346 699 2347
rect 695 2341 699 2342
rect 711 2346 715 2347
rect 711 2341 715 2342
rect 759 2346 763 2347
rect 759 2341 763 2342
rect 799 2346 803 2347
rect 799 2341 803 2342
rect 823 2346 827 2347
rect 823 2341 827 2342
rect 879 2346 883 2347
rect 879 2341 883 2342
rect 887 2346 891 2347
rect 887 2341 891 2342
rect 951 2346 955 2347
rect 951 2341 955 2342
rect 959 2346 963 2347
rect 959 2341 963 2342
rect 1015 2346 1019 2347
rect 1015 2341 1019 2342
rect 1039 2346 1043 2347
rect 1039 2341 1043 2342
rect 1127 2346 1131 2347
rect 1127 2341 1131 2342
rect 1327 2346 1331 2347
rect 1366 2345 1367 2349
rect 1371 2345 1372 2349
rect 1366 2344 1372 2345
rect 2582 2349 2588 2350
rect 2582 2345 2583 2349
rect 2587 2345 2588 2349
rect 2582 2344 2588 2345
rect 1327 2341 1331 2342
rect 112 2329 114 2341
rect 328 2330 330 2341
rect 384 2330 386 2341
rect 440 2330 442 2341
rect 504 2330 506 2341
rect 568 2330 570 2341
rect 632 2330 634 2341
rect 696 2330 698 2341
rect 760 2330 762 2341
rect 824 2330 826 2341
rect 888 2330 890 2341
rect 952 2330 954 2341
rect 1016 2330 1018 2341
rect 326 2329 332 2330
rect 110 2328 116 2329
rect 110 2324 111 2328
rect 115 2324 116 2328
rect 326 2325 327 2329
rect 331 2325 332 2329
rect 326 2324 332 2325
rect 382 2329 388 2330
rect 382 2325 383 2329
rect 387 2325 388 2329
rect 382 2324 388 2325
rect 438 2329 444 2330
rect 438 2325 439 2329
rect 443 2325 444 2329
rect 438 2324 444 2325
rect 502 2329 508 2330
rect 502 2325 503 2329
rect 507 2325 508 2329
rect 502 2324 508 2325
rect 566 2329 572 2330
rect 566 2325 567 2329
rect 571 2325 572 2329
rect 566 2324 572 2325
rect 630 2329 636 2330
rect 630 2325 631 2329
rect 635 2325 636 2329
rect 630 2324 636 2325
rect 694 2329 700 2330
rect 694 2325 695 2329
rect 699 2325 700 2329
rect 694 2324 700 2325
rect 758 2329 764 2330
rect 758 2325 759 2329
rect 763 2325 764 2329
rect 758 2324 764 2325
rect 822 2329 828 2330
rect 822 2325 823 2329
rect 827 2325 828 2329
rect 822 2324 828 2325
rect 886 2329 892 2330
rect 886 2325 887 2329
rect 891 2325 892 2329
rect 886 2324 892 2325
rect 950 2329 956 2330
rect 950 2325 951 2329
rect 955 2325 956 2329
rect 950 2324 956 2325
rect 1014 2329 1020 2330
rect 1328 2329 1330 2341
rect 1366 2332 1372 2333
rect 2582 2332 2588 2333
rect 1014 2325 1015 2329
rect 1019 2325 1020 2329
rect 1014 2324 1020 2325
rect 1326 2328 1332 2329
rect 1326 2324 1327 2328
rect 1331 2324 1332 2328
rect 1366 2328 1367 2332
rect 1371 2328 1372 2332
rect 1366 2327 1372 2328
rect 1454 2331 1460 2332
rect 1454 2327 1455 2331
rect 1459 2327 1460 2331
rect 110 2323 116 2324
rect 1326 2323 1332 2324
rect 1368 2315 1370 2327
rect 1454 2326 1460 2327
rect 1510 2331 1516 2332
rect 1510 2327 1511 2331
rect 1515 2327 1516 2331
rect 1510 2326 1516 2327
rect 1566 2331 1572 2332
rect 1566 2327 1567 2331
rect 1571 2327 1572 2331
rect 1566 2326 1572 2327
rect 1622 2331 1628 2332
rect 1622 2327 1623 2331
rect 1627 2327 1628 2331
rect 1622 2326 1628 2327
rect 1678 2331 1684 2332
rect 1678 2327 1679 2331
rect 1683 2327 1684 2331
rect 2582 2328 2583 2332
rect 2587 2328 2588 2332
rect 2582 2327 2588 2328
rect 1678 2326 1684 2327
rect 1456 2315 1458 2326
rect 1512 2315 1514 2326
rect 1568 2315 1570 2326
rect 1624 2315 1626 2326
rect 1680 2315 1682 2326
rect 2584 2315 2586 2327
rect 1367 2314 1371 2315
rect 110 2311 116 2312
rect 110 2307 111 2311
rect 115 2307 116 2311
rect 110 2306 116 2307
rect 1326 2311 1332 2312
rect 1326 2307 1327 2311
rect 1331 2307 1332 2311
rect 1367 2309 1371 2310
rect 1399 2314 1403 2315
rect 1399 2309 1403 2310
rect 1455 2314 1459 2315
rect 1455 2309 1459 2310
rect 1511 2314 1515 2315
rect 1511 2309 1515 2310
rect 1567 2314 1571 2315
rect 1567 2309 1571 2310
rect 1623 2314 1627 2315
rect 1623 2309 1627 2310
rect 1679 2314 1683 2315
rect 1679 2309 1683 2310
rect 1735 2314 1739 2315
rect 1735 2309 1739 2310
rect 1791 2314 1795 2315
rect 1791 2309 1795 2310
rect 1847 2314 1851 2315
rect 1847 2309 1851 2310
rect 1903 2314 1907 2315
rect 1903 2309 1907 2310
rect 1959 2314 1963 2315
rect 1959 2309 1963 2310
rect 2015 2314 2019 2315
rect 2015 2309 2019 2310
rect 2071 2314 2075 2315
rect 2071 2309 2075 2310
rect 2127 2314 2131 2315
rect 2127 2309 2131 2310
rect 2183 2314 2187 2315
rect 2183 2309 2187 2310
rect 2247 2314 2251 2315
rect 2247 2309 2251 2310
rect 2311 2314 2315 2315
rect 2311 2309 2315 2310
rect 2375 2314 2379 2315
rect 2375 2309 2379 2310
rect 2439 2314 2443 2315
rect 2439 2309 2443 2310
rect 2583 2314 2587 2315
rect 2583 2309 2587 2310
rect 1326 2306 1332 2307
rect 112 2283 114 2306
rect 342 2302 348 2303
rect 342 2298 343 2302
rect 347 2298 348 2302
rect 342 2297 348 2298
rect 398 2302 404 2303
rect 398 2298 399 2302
rect 403 2298 404 2302
rect 398 2297 404 2298
rect 454 2302 460 2303
rect 454 2298 455 2302
rect 459 2298 460 2302
rect 454 2297 460 2298
rect 518 2302 524 2303
rect 518 2298 519 2302
rect 523 2298 524 2302
rect 518 2297 524 2298
rect 582 2302 588 2303
rect 582 2298 583 2302
rect 587 2298 588 2302
rect 582 2297 588 2298
rect 646 2302 652 2303
rect 646 2298 647 2302
rect 651 2298 652 2302
rect 646 2297 652 2298
rect 710 2302 716 2303
rect 710 2298 711 2302
rect 715 2298 716 2302
rect 710 2297 716 2298
rect 774 2302 780 2303
rect 774 2298 775 2302
rect 779 2298 780 2302
rect 774 2297 780 2298
rect 838 2302 844 2303
rect 838 2298 839 2302
rect 843 2298 844 2302
rect 838 2297 844 2298
rect 902 2302 908 2303
rect 902 2298 903 2302
rect 907 2298 908 2302
rect 902 2297 908 2298
rect 966 2302 972 2303
rect 966 2298 967 2302
rect 971 2298 972 2302
rect 966 2297 972 2298
rect 1030 2302 1036 2303
rect 1030 2298 1031 2302
rect 1035 2298 1036 2302
rect 1030 2297 1036 2298
rect 344 2283 346 2297
rect 400 2283 402 2297
rect 456 2283 458 2297
rect 520 2283 522 2297
rect 584 2283 586 2297
rect 648 2283 650 2297
rect 712 2283 714 2297
rect 776 2283 778 2297
rect 840 2283 842 2297
rect 904 2283 906 2297
rect 968 2283 970 2297
rect 1032 2283 1034 2297
rect 1328 2283 1330 2306
rect 1368 2297 1370 2309
rect 1400 2298 1402 2309
rect 1456 2298 1458 2309
rect 1512 2298 1514 2309
rect 1568 2298 1570 2309
rect 1624 2298 1626 2309
rect 1680 2298 1682 2309
rect 1736 2298 1738 2309
rect 1792 2298 1794 2309
rect 1848 2298 1850 2309
rect 1904 2298 1906 2309
rect 1960 2298 1962 2309
rect 2016 2298 2018 2309
rect 2072 2298 2074 2309
rect 2128 2298 2130 2309
rect 2184 2298 2186 2309
rect 2248 2298 2250 2309
rect 2312 2298 2314 2309
rect 2376 2298 2378 2309
rect 2440 2298 2442 2309
rect 1398 2297 1404 2298
rect 1366 2296 1372 2297
rect 1366 2292 1367 2296
rect 1371 2292 1372 2296
rect 1398 2293 1399 2297
rect 1403 2293 1404 2297
rect 1398 2292 1404 2293
rect 1454 2297 1460 2298
rect 1454 2293 1455 2297
rect 1459 2293 1460 2297
rect 1454 2292 1460 2293
rect 1510 2297 1516 2298
rect 1510 2293 1511 2297
rect 1515 2293 1516 2297
rect 1510 2292 1516 2293
rect 1566 2297 1572 2298
rect 1566 2293 1567 2297
rect 1571 2293 1572 2297
rect 1566 2292 1572 2293
rect 1622 2297 1628 2298
rect 1622 2293 1623 2297
rect 1627 2293 1628 2297
rect 1622 2292 1628 2293
rect 1678 2297 1684 2298
rect 1678 2293 1679 2297
rect 1683 2293 1684 2297
rect 1678 2292 1684 2293
rect 1734 2297 1740 2298
rect 1734 2293 1735 2297
rect 1739 2293 1740 2297
rect 1734 2292 1740 2293
rect 1790 2297 1796 2298
rect 1790 2293 1791 2297
rect 1795 2293 1796 2297
rect 1790 2292 1796 2293
rect 1846 2297 1852 2298
rect 1846 2293 1847 2297
rect 1851 2293 1852 2297
rect 1846 2292 1852 2293
rect 1902 2297 1908 2298
rect 1902 2293 1903 2297
rect 1907 2293 1908 2297
rect 1902 2292 1908 2293
rect 1958 2297 1964 2298
rect 1958 2293 1959 2297
rect 1963 2293 1964 2297
rect 1958 2292 1964 2293
rect 2014 2297 2020 2298
rect 2014 2293 2015 2297
rect 2019 2293 2020 2297
rect 2014 2292 2020 2293
rect 2070 2297 2076 2298
rect 2070 2293 2071 2297
rect 2075 2293 2076 2297
rect 2070 2292 2076 2293
rect 2126 2297 2132 2298
rect 2126 2293 2127 2297
rect 2131 2293 2132 2297
rect 2126 2292 2132 2293
rect 2182 2297 2188 2298
rect 2182 2293 2183 2297
rect 2187 2293 2188 2297
rect 2182 2292 2188 2293
rect 2246 2297 2252 2298
rect 2246 2293 2247 2297
rect 2251 2293 2252 2297
rect 2246 2292 2252 2293
rect 2310 2297 2316 2298
rect 2310 2293 2311 2297
rect 2315 2293 2316 2297
rect 2310 2292 2316 2293
rect 2374 2297 2380 2298
rect 2374 2293 2375 2297
rect 2379 2293 2380 2297
rect 2374 2292 2380 2293
rect 2438 2297 2444 2298
rect 2584 2297 2586 2309
rect 2438 2293 2439 2297
rect 2443 2293 2444 2297
rect 2438 2292 2444 2293
rect 2582 2296 2588 2297
rect 2582 2292 2583 2296
rect 2587 2292 2588 2296
rect 1366 2291 1372 2292
rect 2582 2291 2588 2292
rect 111 2282 115 2283
rect 111 2277 115 2278
rect 343 2282 347 2283
rect 343 2277 347 2278
rect 399 2282 403 2283
rect 399 2277 403 2278
rect 407 2282 411 2283
rect 407 2277 411 2278
rect 455 2282 459 2283
rect 455 2277 459 2278
rect 463 2282 467 2283
rect 463 2277 467 2278
rect 519 2282 523 2283
rect 519 2277 523 2278
rect 575 2282 579 2283
rect 575 2277 579 2278
rect 583 2282 587 2283
rect 583 2277 587 2278
rect 631 2282 635 2283
rect 631 2277 635 2278
rect 647 2282 651 2283
rect 647 2277 651 2278
rect 687 2282 691 2283
rect 687 2277 691 2278
rect 711 2282 715 2283
rect 711 2277 715 2278
rect 743 2282 747 2283
rect 743 2277 747 2278
rect 775 2282 779 2283
rect 775 2277 779 2278
rect 799 2282 803 2283
rect 799 2277 803 2278
rect 839 2282 843 2283
rect 839 2277 843 2278
rect 855 2282 859 2283
rect 855 2277 859 2278
rect 903 2282 907 2283
rect 903 2277 907 2278
rect 911 2282 915 2283
rect 911 2277 915 2278
rect 967 2282 971 2283
rect 967 2277 971 2278
rect 1031 2282 1035 2283
rect 1031 2277 1035 2278
rect 1327 2282 1331 2283
rect 1327 2277 1331 2278
rect 1366 2279 1372 2280
rect 112 2262 114 2277
rect 408 2271 410 2277
rect 464 2271 466 2277
rect 520 2271 522 2277
rect 576 2271 578 2277
rect 632 2271 634 2277
rect 688 2271 690 2277
rect 744 2271 746 2277
rect 800 2271 802 2277
rect 856 2271 858 2277
rect 912 2271 914 2277
rect 968 2271 970 2277
rect 406 2270 412 2271
rect 406 2266 407 2270
rect 411 2266 412 2270
rect 406 2265 412 2266
rect 462 2270 468 2271
rect 462 2266 463 2270
rect 467 2266 468 2270
rect 462 2265 468 2266
rect 518 2270 524 2271
rect 518 2266 519 2270
rect 523 2266 524 2270
rect 518 2265 524 2266
rect 574 2270 580 2271
rect 574 2266 575 2270
rect 579 2266 580 2270
rect 574 2265 580 2266
rect 630 2270 636 2271
rect 630 2266 631 2270
rect 635 2266 636 2270
rect 630 2265 636 2266
rect 686 2270 692 2271
rect 686 2266 687 2270
rect 691 2266 692 2270
rect 686 2265 692 2266
rect 742 2270 748 2271
rect 742 2266 743 2270
rect 747 2266 748 2270
rect 742 2265 748 2266
rect 798 2270 804 2271
rect 798 2266 799 2270
rect 803 2266 804 2270
rect 798 2265 804 2266
rect 854 2270 860 2271
rect 854 2266 855 2270
rect 859 2266 860 2270
rect 854 2265 860 2266
rect 910 2270 916 2271
rect 910 2266 911 2270
rect 915 2266 916 2270
rect 910 2265 916 2266
rect 966 2270 972 2271
rect 966 2266 967 2270
rect 971 2266 972 2270
rect 966 2265 972 2266
rect 1328 2262 1330 2277
rect 1366 2275 1367 2279
rect 1371 2275 1372 2279
rect 1366 2274 1372 2275
rect 2582 2279 2588 2280
rect 2582 2275 2583 2279
rect 2587 2275 2588 2279
rect 2582 2274 2588 2275
rect 110 2261 116 2262
rect 110 2257 111 2261
rect 115 2257 116 2261
rect 110 2256 116 2257
rect 1326 2261 1332 2262
rect 1326 2257 1327 2261
rect 1331 2257 1332 2261
rect 1368 2259 1370 2274
rect 1414 2270 1420 2271
rect 1414 2266 1415 2270
rect 1419 2266 1420 2270
rect 1414 2265 1420 2266
rect 1470 2270 1476 2271
rect 1470 2266 1471 2270
rect 1475 2266 1476 2270
rect 1470 2265 1476 2266
rect 1526 2270 1532 2271
rect 1526 2266 1527 2270
rect 1531 2266 1532 2270
rect 1526 2265 1532 2266
rect 1582 2270 1588 2271
rect 1582 2266 1583 2270
rect 1587 2266 1588 2270
rect 1582 2265 1588 2266
rect 1638 2270 1644 2271
rect 1638 2266 1639 2270
rect 1643 2266 1644 2270
rect 1638 2265 1644 2266
rect 1694 2270 1700 2271
rect 1694 2266 1695 2270
rect 1699 2266 1700 2270
rect 1694 2265 1700 2266
rect 1750 2270 1756 2271
rect 1750 2266 1751 2270
rect 1755 2266 1756 2270
rect 1750 2265 1756 2266
rect 1806 2270 1812 2271
rect 1806 2266 1807 2270
rect 1811 2266 1812 2270
rect 1806 2265 1812 2266
rect 1862 2270 1868 2271
rect 1862 2266 1863 2270
rect 1867 2266 1868 2270
rect 1862 2265 1868 2266
rect 1918 2270 1924 2271
rect 1918 2266 1919 2270
rect 1923 2266 1924 2270
rect 1918 2265 1924 2266
rect 1974 2270 1980 2271
rect 1974 2266 1975 2270
rect 1979 2266 1980 2270
rect 1974 2265 1980 2266
rect 2030 2270 2036 2271
rect 2030 2266 2031 2270
rect 2035 2266 2036 2270
rect 2030 2265 2036 2266
rect 2086 2270 2092 2271
rect 2086 2266 2087 2270
rect 2091 2266 2092 2270
rect 2086 2265 2092 2266
rect 2142 2270 2148 2271
rect 2142 2266 2143 2270
rect 2147 2266 2148 2270
rect 2142 2265 2148 2266
rect 2198 2270 2204 2271
rect 2198 2266 2199 2270
rect 2203 2266 2204 2270
rect 2198 2265 2204 2266
rect 2262 2270 2268 2271
rect 2262 2266 2263 2270
rect 2267 2266 2268 2270
rect 2262 2265 2268 2266
rect 2326 2270 2332 2271
rect 2326 2266 2327 2270
rect 2331 2266 2332 2270
rect 2326 2265 2332 2266
rect 2390 2270 2396 2271
rect 2390 2266 2391 2270
rect 2395 2266 2396 2270
rect 2390 2265 2396 2266
rect 2454 2270 2460 2271
rect 2454 2266 2455 2270
rect 2459 2266 2460 2270
rect 2454 2265 2460 2266
rect 1416 2259 1418 2265
rect 1472 2259 1474 2265
rect 1528 2259 1530 2265
rect 1584 2259 1586 2265
rect 1640 2259 1642 2265
rect 1696 2259 1698 2265
rect 1752 2259 1754 2265
rect 1808 2259 1810 2265
rect 1864 2259 1866 2265
rect 1920 2259 1922 2265
rect 1976 2259 1978 2265
rect 2032 2259 2034 2265
rect 2088 2259 2090 2265
rect 2144 2259 2146 2265
rect 2200 2259 2202 2265
rect 2264 2259 2266 2265
rect 2328 2259 2330 2265
rect 2392 2259 2394 2265
rect 2456 2259 2458 2265
rect 2584 2259 2586 2274
rect 1326 2256 1332 2257
rect 1367 2258 1371 2259
rect 1367 2253 1371 2254
rect 1415 2258 1419 2259
rect 1415 2253 1419 2254
rect 1471 2258 1475 2259
rect 1471 2253 1475 2254
rect 1511 2258 1515 2259
rect 1511 2253 1515 2254
rect 1527 2258 1531 2259
rect 1527 2253 1531 2254
rect 1583 2258 1587 2259
rect 1583 2253 1587 2254
rect 1623 2258 1627 2259
rect 1623 2253 1627 2254
rect 1639 2258 1643 2259
rect 1639 2253 1643 2254
rect 1695 2258 1699 2259
rect 1695 2253 1699 2254
rect 1727 2258 1731 2259
rect 1727 2253 1731 2254
rect 1751 2258 1755 2259
rect 1751 2253 1755 2254
rect 1807 2258 1811 2259
rect 1807 2253 1811 2254
rect 1823 2258 1827 2259
rect 1823 2253 1827 2254
rect 1863 2258 1867 2259
rect 1863 2253 1867 2254
rect 1903 2258 1907 2259
rect 1903 2253 1907 2254
rect 1919 2258 1923 2259
rect 1919 2253 1923 2254
rect 1975 2258 1979 2259
rect 1975 2253 1979 2254
rect 1983 2258 1987 2259
rect 1983 2253 1987 2254
rect 2031 2258 2035 2259
rect 2031 2253 2035 2254
rect 2055 2258 2059 2259
rect 2055 2253 2059 2254
rect 2087 2258 2091 2259
rect 2087 2253 2091 2254
rect 2119 2258 2123 2259
rect 2119 2253 2123 2254
rect 2143 2258 2147 2259
rect 2143 2253 2147 2254
rect 2191 2258 2195 2259
rect 2191 2253 2195 2254
rect 2199 2258 2203 2259
rect 2199 2253 2203 2254
rect 2263 2258 2267 2259
rect 2263 2253 2267 2254
rect 2327 2258 2331 2259
rect 2327 2253 2331 2254
rect 2335 2258 2339 2259
rect 2335 2253 2339 2254
rect 2391 2258 2395 2259
rect 2391 2253 2395 2254
rect 2455 2258 2459 2259
rect 2455 2253 2459 2254
rect 2583 2258 2587 2259
rect 2583 2253 2587 2254
rect 110 2244 116 2245
rect 1326 2244 1332 2245
rect 110 2240 111 2244
rect 115 2240 116 2244
rect 110 2239 116 2240
rect 390 2243 396 2244
rect 390 2239 391 2243
rect 395 2239 396 2243
rect 112 2223 114 2239
rect 390 2238 396 2239
rect 446 2243 452 2244
rect 446 2239 447 2243
rect 451 2239 452 2243
rect 446 2238 452 2239
rect 502 2243 508 2244
rect 502 2239 503 2243
rect 507 2239 508 2243
rect 502 2238 508 2239
rect 558 2243 564 2244
rect 558 2239 559 2243
rect 563 2239 564 2243
rect 558 2238 564 2239
rect 614 2243 620 2244
rect 614 2239 615 2243
rect 619 2239 620 2243
rect 614 2238 620 2239
rect 670 2243 676 2244
rect 670 2239 671 2243
rect 675 2239 676 2243
rect 670 2238 676 2239
rect 726 2243 732 2244
rect 726 2239 727 2243
rect 731 2239 732 2243
rect 726 2238 732 2239
rect 782 2243 788 2244
rect 782 2239 783 2243
rect 787 2239 788 2243
rect 782 2238 788 2239
rect 838 2243 844 2244
rect 838 2239 839 2243
rect 843 2239 844 2243
rect 838 2238 844 2239
rect 894 2243 900 2244
rect 894 2239 895 2243
rect 899 2239 900 2243
rect 894 2238 900 2239
rect 950 2243 956 2244
rect 950 2239 951 2243
rect 955 2239 956 2243
rect 1326 2240 1327 2244
rect 1331 2240 1332 2244
rect 1326 2239 1332 2240
rect 950 2238 956 2239
rect 392 2223 394 2238
rect 448 2223 450 2238
rect 504 2223 506 2238
rect 560 2223 562 2238
rect 616 2223 618 2238
rect 672 2223 674 2238
rect 728 2223 730 2238
rect 784 2223 786 2238
rect 840 2223 842 2238
rect 896 2223 898 2238
rect 952 2223 954 2238
rect 1328 2223 1330 2239
rect 1368 2238 1370 2253
rect 1416 2247 1418 2253
rect 1512 2247 1514 2253
rect 1624 2247 1626 2253
rect 1728 2247 1730 2253
rect 1824 2247 1826 2253
rect 1904 2247 1906 2253
rect 1984 2247 1986 2253
rect 2056 2247 2058 2253
rect 2120 2247 2122 2253
rect 2192 2247 2194 2253
rect 2264 2247 2266 2253
rect 2336 2247 2338 2253
rect 1414 2246 1420 2247
rect 1414 2242 1415 2246
rect 1419 2242 1420 2246
rect 1414 2241 1420 2242
rect 1510 2246 1516 2247
rect 1510 2242 1511 2246
rect 1515 2242 1516 2246
rect 1510 2241 1516 2242
rect 1622 2246 1628 2247
rect 1622 2242 1623 2246
rect 1627 2242 1628 2246
rect 1622 2241 1628 2242
rect 1726 2246 1732 2247
rect 1726 2242 1727 2246
rect 1731 2242 1732 2246
rect 1726 2241 1732 2242
rect 1822 2246 1828 2247
rect 1822 2242 1823 2246
rect 1827 2242 1828 2246
rect 1822 2241 1828 2242
rect 1902 2246 1908 2247
rect 1902 2242 1903 2246
rect 1907 2242 1908 2246
rect 1902 2241 1908 2242
rect 1982 2246 1988 2247
rect 1982 2242 1983 2246
rect 1987 2242 1988 2246
rect 1982 2241 1988 2242
rect 2054 2246 2060 2247
rect 2054 2242 2055 2246
rect 2059 2242 2060 2246
rect 2054 2241 2060 2242
rect 2118 2246 2124 2247
rect 2118 2242 2119 2246
rect 2123 2242 2124 2246
rect 2118 2241 2124 2242
rect 2190 2246 2196 2247
rect 2190 2242 2191 2246
rect 2195 2242 2196 2246
rect 2190 2241 2196 2242
rect 2262 2246 2268 2247
rect 2262 2242 2263 2246
rect 2267 2242 2268 2246
rect 2262 2241 2268 2242
rect 2334 2246 2340 2247
rect 2334 2242 2335 2246
rect 2339 2242 2340 2246
rect 2334 2241 2340 2242
rect 2584 2238 2586 2253
rect 1366 2237 1372 2238
rect 1366 2233 1367 2237
rect 1371 2233 1372 2237
rect 1366 2232 1372 2233
rect 2582 2237 2588 2238
rect 2582 2233 2583 2237
rect 2587 2233 2588 2237
rect 2582 2232 2588 2233
rect 111 2222 115 2223
rect 111 2217 115 2218
rect 391 2222 395 2223
rect 391 2217 395 2218
rect 423 2222 427 2223
rect 423 2217 427 2218
rect 447 2222 451 2223
rect 447 2217 451 2218
rect 479 2222 483 2223
rect 479 2217 483 2218
rect 503 2222 507 2223
rect 503 2217 507 2218
rect 535 2222 539 2223
rect 535 2217 539 2218
rect 559 2222 563 2223
rect 559 2217 563 2218
rect 591 2222 595 2223
rect 591 2217 595 2218
rect 615 2222 619 2223
rect 615 2217 619 2218
rect 647 2222 651 2223
rect 647 2217 651 2218
rect 671 2222 675 2223
rect 671 2217 675 2218
rect 711 2222 715 2223
rect 711 2217 715 2218
rect 727 2222 731 2223
rect 727 2217 731 2218
rect 783 2222 787 2223
rect 783 2217 787 2218
rect 839 2222 843 2223
rect 839 2217 843 2218
rect 855 2222 859 2223
rect 855 2217 859 2218
rect 895 2222 899 2223
rect 895 2217 899 2218
rect 927 2222 931 2223
rect 927 2217 931 2218
rect 951 2222 955 2223
rect 951 2217 955 2218
rect 999 2222 1003 2223
rect 999 2217 1003 2218
rect 1071 2222 1075 2223
rect 1071 2217 1075 2218
rect 1143 2222 1147 2223
rect 1143 2217 1147 2218
rect 1215 2222 1219 2223
rect 1215 2217 1219 2218
rect 1271 2222 1275 2223
rect 1271 2217 1275 2218
rect 1327 2222 1331 2223
rect 1327 2217 1331 2218
rect 1366 2220 1372 2221
rect 2582 2220 2588 2221
rect 112 2205 114 2217
rect 424 2206 426 2217
rect 480 2206 482 2217
rect 536 2206 538 2217
rect 592 2206 594 2217
rect 648 2206 650 2217
rect 712 2206 714 2217
rect 784 2206 786 2217
rect 856 2206 858 2217
rect 928 2206 930 2217
rect 1000 2206 1002 2217
rect 1072 2206 1074 2217
rect 1144 2206 1146 2217
rect 1216 2206 1218 2217
rect 1272 2206 1274 2217
rect 422 2205 428 2206
rect 110 2204 116 2205
rect 110 2200 111 2204
rect 115 2200 116 2204
rect 422 2201 423 2205
rect 427 2201 428 2205
rect 422 2200 428 2201
rect 478 2205 484 2206
rect 478 2201 479 2205
rect 483 2201 484 2205
rect 478 2200 484 2201
rect 534 2205 540 2206
rect 534 2201 535 2205
rect 539 2201 540 2205
rect 534 2200 540 2201
rect 590 2205 596 2206
rect 590 2201 591 2205
rect 595 2201 596 2205
rect 590 2200 596 2201
rect 646 2205 652 2206
rect 646 2201 647 2205
rect 651 2201 652 2205
rect 646 2200 652 2201
rect 710 2205 716 2206
rect 710 2201 711 2205
rect 715 2201 716 2205
rect 710 2200 716 2201
rect 782 2205 788 2206
rect 782 2201 783 2205
rect 787 2201 788 2205
rect 782 2200 788 2201
rect 854 2205 860 2206
rect 854 2201 855 2205
rect 859 2201 860 2205
rect 854 2200 860 2201
rect 926 2205 932 2206
rect 926 2201 927 2205
rect 931 2201 932 2205
rect 926 2200 932 2201
rect 998 2205 1004 2206
rect 998 2201 999 2205
rect 1003 2201 1004 2205
rect 998 2200 1004 2201
rect 1070 2205 1076 2206
rect 1070 2201 1071 2205
rect 1075 2201 1076 2205
rect 1070 2200 1076 2201
rect 1142 2205 1148 2206
rect 1142 2201 1143 2205
rect 1147 2201 1148 2205
rect 1142 2200 1148 2201
rect 1214 2205 1220 2206
rect 1214 2201 1215 2205
rect 1219 2201 1220 2205
rect 1214 2200 1220 2201
rect 1270 2205 1276 2206
rect 1328 2205 1330 2217
rect 1366 2216 1367 2220
rect 1371 2216 1372 2220
rect 1366 2215 1372 2216
rect 1398 2219 1404 2220
rect 1398 2215 1399 2219
rect 1403 2215 1404 2219
rect 1270 2201 1271 2205
rect 1275 2201 1276 2205
rect 1270 2200 1276 2201
rect 1326 2204 1332 2205
rect 1326 2200 1327 2204
rect 1331 2200 1332 2204
rect 110 2199 116 2200
rect 1326 2199 1332 2200
rect 1368 2199 1370 2215
rect 1398 2214 1404 2215
rect 1494 2219 1500 2220
rect 1494 2215 1495 2219
rect 1499 2215 1500 2219
rect 1494 2214 1500 2215
rect 1606 2219 1612 2220
rect 1606 2215 1607 2219
rect 1611 2215 1612 2219
rect 1606 2214 1612 2215
rect 1710 2219 1716 2220
rect 1710 2215 1711 2219
rect 1715 2215 1716 2219
rect 1710 2214 1716 2215
rect 1806 2219 1812 2220
rect 1806 2215 1807 2219
rect 1811 2215 1812 2219
rect 1806 2214 1812 2215
rect 1886 2219 1892 2220
rect 1886 2215 1887 2219
rect 1891 2215 1892 2219
rect 1886 2214 1892 2215
rect 1966 2219 1972 2220
rect 1966 2215 1967 2219
rect 1971 2215 1972 2219
rect 1966 2214 1972 2215
rect 2038 2219 2044 2220
rect 2038 2215 2039 2219
rect 2043 2215 2044 2219
rect 2038 2214 2044 2215
rect 2102 2219 2108 2220
rect 2102 2215 2103 2219
rect 2107 2215 2108 2219
rect 2102 2214 2108 2215
rect 2174 2219 2180 2220
rect 2174 2215 2175 2219
rect 2179 2215 2180 2219
rect 2174 2214 2180 2215
rect 2246 2219 2252 2220
rect 2246 2215 2247 2219
rect 2251 2215 2252 2219
rect 2246 2214 2252 2215
rect 2318 2219 2324 2220
rect 2318 2215 2319 2219
rect 2323 2215 2324 2219
rect 2582 2216 2583 2220
rect 2587 2216 2588 2220
rect 2582 2215 2588 2216
rect 2318 2214 2324 2215
rect 1400 2199 1402 2214
rect 1496 2199 1498 2214
rect 1608 2199 1610 2214
rect 1712 2199 1714 2214
rect 1808 2199 1810 2214
rect 1888 2199 1890 2214
rect 1968 2199 1970 2214
rect 2040 2199 2042 2214
rect 2104 2199 2106 2214
rect 2176 2199 2178 2214
rect 2248 2199 2250 2214
rect 2320 2199 2322 2214
rect 2584 2199 2586 2215
rect 1367 2198 1371 2199
rect 1367 2193 1371 2194
rect 1399 2198 1403 2199
rect 1399 2193 1403 2194
rect 1495 2198 1499 2199
rect 1495 2193 1499 2194
rect 1607 2198 1611 2199
rect 1607 2193 1611 2194
rect 1711 2198 1715 2199
rect 1711 2193 1715 2194
rect 1751 2198 1755 2199
rect 1751 2193 1755 2194
rect 1807 2198 1811 2199
rect 1807 2193 1811 2194
rect 1839 2198 1843 2199
rect 1839 2193 1843 2194
rect 1887 2198 1891 2199
rect 1887 2193 1891 2194
rect 1927 2198 1931 2199
rect 1927 2193 1931 2194
rect 1967 2198 1971 2199
rect 1967 2193 1971 2194
rect 2007 2198 2011 2199
rect 2007 2193 2011 2194
rect 2039 2198 2043 2199
rect 2039 2193 2043 2194
rect 2087 2198 2091 2199
rect 2087 2193 2091 2194
rect 2103 2198 2107 2199
rect 2103 2193 2107 2194
rect 2167 2198 2171 2199
rect 2167 2193 2171 2194
rect 2175 2198 2179 2199
rect 2175 2193 2179 2194
rect 2247 2198 2251 2199
rect 2247 2193 2251 2194
rect 2319 2198 2323 2199
rect 2319 2193 2323 2194
rect 2335 2198 2339 2199
rect 2335 2193 2339 2194
rect 2423 2198 2427 2199
rect 2423 2193 2427 2194
rect 2583 2198 2587 2199
rect 2583 2193 2587 2194
rect 110 2187 116 2188
rect 110 2183 111 2187
rect 115 2183 116 2187
rect 110 2182 116 2183
rect 1326 2187 1332 2188
rect 1326 2183 1327 2187
rect 1331 2183 1332 2187
rect 1326 2182 1332 2183
rect 112 2159 114 2182
rect 438 2178 444 2179
rect 438 2174 439 2178
rect 443 2174 444 2178
rect 438 2173 444 2174
rect 494 2178 500 2179
rect 494 2174 495 2178
rect 499 2174 500 2178
rect 494 2173 500 2174
rect 550 2178 556 2179
rect 550 2174 551 2178
rect 555 2174 556 2178
rect 550 2173 556 2174
rect 606 2178 612 2179
rect 606 2174 607 2178
rect 611 2174 612 2178
rect 606 2173 612 2174
rect 662 2178 668 2179
rect 662 2174 663 2178
rect 667 2174 668 2178
rect 662 2173 668 2174
rect 726 2178 732 2179
rect 726 2174 727 2178
rect 731 2174 732 2178
rect 726 2173 732 2174
rect 798 2178 804 2179
rect 798 2174 799 2178
rect 803 2174 804 2178
rect 798 2173 804 2174
rect 870 2178 876 2179
rect 870 2174 871 2178
rect 875 2174 876 2178
rect 870 2173 876 2174
rect 942 2178 948 2179
rect 942 2174 943 2178
rect 947 2174 948 2178
rect 942 2173 948 2174
rect 1014 2178 1020 2179
rect 1014 2174 1015 2178
rect 1019 2174 1020 2178
rect 1014 2173 1020 2174
rect 1086 2178 1092 2179
rect 1086 2174 1087 2178
rect 1091 2174 1092 2178
rect 1086 2173 1092 2174
rect 1158 2178 1164 2179
rect 1158 2174 1159 2178
rect 1163 2174 1164 2178
rect 1158 2173 1164 2174
rect 1230 2178 1236 2179
rect 1230 2174 1231 2178
rect 1235 2174 1236 2178
rect 1230 2173 1236 2174
rect 1286 2178 1292 2179
rect 1286 2174 1287 2178
rect 1291 2174 1292 2178
rect 1286 2173 1292 2174
rect 440 2159 442 2173
rect 496 2159 498 2173
rect 552 2159 554 2173
rect 608 2159 610 2173
rect 664 2159 666 2173
rect 728 2159 730 2173
rect 800 2159 802 2173
rect 872 2159 874 2173
rect 944 2159 946 2173
rect 1016 2159 1018 2173
rect 1088 2159 1090 2173
rect 1160 2159 1162 2173
rect 1232 2159 1234 2173
rect 1288 2159 1290 2173
rect 1328 2159 1330 2182
rect 1368 2181 1370 2193
rect 1752 2182 1754 2193
rect 1840 2182 1842 2193
rect 1928 2182 1930 2193
rect 2008 2182 2010 2193
rect 2088 2182 2090 2193
rect 2168 2182 2170 2193
rect 2248 2182 2250 2193
rect 2336 2182 2338 2193
rect 2424 2182 2426 2193
rect 1750 2181 1756 2182
rect 1366 2180 1372 2181
rect 1366 2176 1367 2180
rect 1371 2176 1372 2180
rect 1750 2177 1751 2181
rect 1755 2177 1756 2181
rect 1750 2176 1756 2177
rect 1838 2181 1844 2182
rect 1838 2177 1839 2181
rect 1843 2177 1844 2181
rect 1838 2176 1844 2177
rect 1926 2181 1932 2182
rect 1926 2177 1927 2181
rect 1931 2177 1932 2181
rect 1926 2176 1932 2177
rect 2006 2181 2012 2182
rect 2006 2177 2007 2181
rect 2011 2177 2012 2181
rect 2006 2176 2012 2177
rect 2086 2181 2092 2182
rect 2086 2177 2087 2181
rect 2091 2177 2092 2181
rect 2086 2176 2092 2177
rect 2166 2181 2172 2182
rect 2166 2177 2167 2181
rect 2171 2177 2172 2181
rect 2166 2176 2172 2177
rect 2246 2181 2252 2182
rect 2246 2177 2247 2181
rect 2251 2177 2252 2181
rect 2246 2176 2252 2177
rect 2334 2181 2340 2182
rect 2334 2177 2335 2181
rect 2339 2177 2340 2181
rect 2334 2176 2340 2177
rect 2422 2181 2428 2182
rect 2584 2181 2586 2193
rect 2422 2177 2423 2181
rect 2427 2177 2428 2181
rect 2422 2176 2428 2177
rect 2582 2180 2588 2181
rect 2582 2176 2583 2180
rect 2587 2176 2588 2180
rect 1366 2175 1372 2176
rect 2582 2175 2588 2176
rect 1366 2163 1372 2164
rect 1366 2159 1367 2163
rect 1371 2159 1372 2163
rect 111 2158 115 2159
rect 111 2153 115 2154
rect 199 2158 203 2159
rect 199 2153 203 2154
rect 271 2158 275 2159
rect 271 2153 275 2154
rect 351 2158 355 2159
rect 351 2153 355 2154
rect 439 2158 443 2159
rect 439 2153 443 2154
rect 447 2158 451 2159
rect 447 2153 451 2154
rect 495 2158 499 2159
rect 495 2153 499 2154
rect 551 2158 555 2159
rect 551 2153 555 2154
rect 607 2158 611 2159
rect 607 2153 611 2154
rect 663 2158 667 2159
rect 663 2153 667 2154
rect 727 2158 731 2159
rect 727 2153 731 2154
rect 775 2158 779 2159
rect 775 2153 779 2154
rect 799 2158 803 2159
rect 799 2153 803 2154
rect 871 2158 875 2159
rect 871 2153 875 2154
rect 879 2158 883 2159
rect 879 2153 883 2154
rect 943 2158 947 2159
rect 943 2153 947 2154
rect 983 2158 987 2159
rect 983 2153 987 2154
rect 1015 2158 1019 2159
rect 1015 2153 1019 2154
rect 1079 2158 1083 2159
rect 1079 2153 1083 2154
rect 1087 2158 1091 2159
rect 1087 2153 1091 2154
rect 1159 2158 1163 2159
rect 1159 2153 1163 2154
rect 1183 2158 1187 2159
rect 1183 2153 1187 2154
rect 1231 2158 1235 2159
rect 1231 2153 1235 2154
rect 1287 2158 1291 2159
rect 1287 2153 1291 2154
rect 1327 2158 1331 2159
rect 1366 2158 1372 2159
rect 2582 2163 2588 2164
rect 2582 2159 2583 2163
rect 2587 2159 2588 2163
rect 2582 2158 2588 2159
rect 1327 2153 1331 2154
rect 112 2138 114 2153
rect 200 2147 202 2153
rect 272 2147 274 2153
rect 352 2147 354 2153
rect 448 2147 450 2153
rect 552 2147 554 2153
rect 664 2147 666 2153
rect 776 2147 778 2153
rect 880 2147 882 2153
rect 984 2147 986 2153
rect 1080 2147 1082 2153
rect 1184 2147 1186 2153
rect 1288 2147 1290 2153
rect 198 2146 204 2147
rect 198 2142 199 2146
rect 203 2142 204 2146
rect 198 2141 204 2142
rect 270 2146 276 2147
rect 270 2142 271 2146
rect 275 2142 276 2146
rect 270 2141 276 2142
rect 350 2146 356 2147
rect 350 2142 351 2146
rect 355 2142 356 2146
rect 350 2141 356 2142
rect 446 2146 452 2147
rect 446 2142 447 2146
rect 451 2142 452 2146
rect 446 2141 452 2142
rect 550 2146 556 2147
rect 550 2142 551 2146
rect 555 2142 556 2146
rect 550 2141 556 2142
rect 662 2146 668 2147
rect 662 2142 663 2146
rect 667 2142 668 2146
rect 662 2141 668 2142
rect 774 2146 780 2147
rect 774 2142 775 2146
rect 779 2142 780 2146
rect 774 2141 780 2142
rect 878 2146 884 2147
rect 878 2142 879 2146
rect 883 2142 884 2146
rect 878 2141 884 2142
rect 982 2146 988 2147
rect 982 2142 983 2146
rect 987 2142 988 2146
rect 982 2141 988 2142
rect 1078 2146 1084 2147
rect 1078 2142 1079 2146
rect 1083 2142 1084 2146
rect 1078 2141 1084 2142
rect 1182 2146 1188 2147
rect 1182 2142 1183 2146
rect 1187 2142 1188 2146
rect 1182 2141 1188 2142
rect 1286 2146 1292 2147
rect 1286 2142 1287 2146
rect 1291 2142 1292 2146
rect 1286 2141 1292 2142
rect 1328 2138 1330 2153
rect 1368 2143 1370 2158
rect 1766 2154 1772 2155
rect 1766 2150 1767 2154
rect 1771 2150 1772 2154
rect 1766 2149 1772 2150
rect 1854 2154 1860 2155
rect 1854 2150 1855 2154
rect 1859 2150 1860 2154
rect 1854 2149 1860 2150
rect 1942 2154 1948 2155
rect 1942 2150 1943 2154
rect 1947 2150 1948 2154
rect 1942 2149 1948 2150
rect 2022 2154 2028 2155
rect 2022 2150 2023 2154
rect 2027 2150 2028 2154
rect 2022 2149 2028 2150
rect 2102 2154 2108 2155
rect 2102 2150 2103 2154
rect 2107 2150 2108 2154
rect 2102 2149 2108 2150
rect 2182 2154 2188 2155
rect 2182 2150 2183 2154
rect 2187 2150 2188 2154
rect 2182 2149 2188 2150
rect 2262 2154 2268 2155
rect 2262 2150 2263 2154
rect 2267 2150 2268 2154
rect 2262 2149 2268 2150
rect 2350 2154 2356 2155
rect 2350 2150 2351 2154
rect 2355 2150 2356 2154
rect 2350 2149 2356 2150
rect 2438 2154 2444 2155
rect 2438 2150 2439 2154
rect 2443 2150 2444 2154
rect 2438 2149 2444 2150
rect 1768 2143 1770 2149
rect 1856 2143 1858 2149
rect 1944 2143 1946 2149
rect 2024 2143 2026 2149
rect 2104 2143 2106 2149
rect 2184 2143 2186 2149
rect 2264 2143 2266 2149
rect 2352 2143 2354 2149
rect 2440 2143 2442 2149
rect 2584 2143 2586 2158
rect 1367 2142 1371 2143
rect 110 2137 116 2138
rect 110 2133 111 2137
rect 115 2133 116 2137
rect 110 2132 116 2133
rect 1326 2137 1332 2138
rect 1367 2137 1371 2138
rect 1607 2142 1611 2143
rect 1607 2137 1611 2138
rect 1679 2142 1683 2143
rect 1679 2137 1683 2138
rect 1767 2142 1771 2143
rect 1767 2137 1771 2138
rect 1855 2142 1859 2143
rect 1855 2137 1859 2138
rect 1863 2142 1867 2143
rect 1863 2137 1867 2138
rect 1943 2142 1947 2143
rect 1943 2137 1947 2138
rect 1959 2142 1963 2143
rect 1959 2137 1963 2138
rect 2023 2142 2027 2143
rect 2023 2137 2027 2138
rect 2063 2142 2067 2143
rect 2063 2137 2067 2138
rect 2103 2142 2107 2143
rect 2103 2137 2107 2138
rect 2159 2142 2163 2143
rect 2159 2137 2163 2138
rect 2183 2142 2187 2143
rect 2183 2137 2187 2138
rect 2255 2142 2259 2143
rect 2255 2137 2259 2138
rect 2263 2142 2267 2143
rect 2263 2137 2267 2138
rect 2351 2142 2355 2143
rect 2351 2137 2355 2138
rect 2439 2142 2443 2143
rect 2439 2137 2443 2138
rect 2447 2142 2451 2143
rect 2447 2137 2451 2138
rect 2543 2142 2547 2143
rect 2543 2137 2547 2138
rect 2583 2142 2587 2143
rect 2583 2137 2587 2138
rect 1326 2133 1327 2137
rect 1331 2133 1332 2137
rect 1326 2132 1332 2133
rect 1368 2122 1370 2137
rect 1608 2131 1610 2137
rect 1680 2131 1682 2137
rect 1768 2131 1770 2137
rect 1864 2131 1866 2137
rect 1960 2131 1962 2137
rect 2064 2131 2066 2137
rect 2160 2131 2162 2137
rect 2256 2131 2258 2137
rect 2352 2131 2354 2137
rect 2448 2131 2450 2137
rect 2544 2131 2546 2137
rect 1606 2130 1612 2131
rect 1606 2126 1607 2130
rect 1611 2126 1612 2130
rect 1606 2125 1612 2126
rect 1678 2130 1684 2131
rect 1678 2126 1679 2130
rect 1683 2126 1684 2130
rect 1678 2125 1684 2126
rect 1766 2130 1772 2131
rect 1766 2126 1767 2130
rect 1771 2126 1772 2130
rect 1766 2125 1772 2126
rect 1862 2130 1868 2131
rect 1862 2126 1863 2130
rect 1867 2126 1868 2130
rect 1862 2125 1868 2126
rect 1958 2130 1964 2131
rect 1958 2126 1959 2130
rect 1963 2126 1964 2130
rect 1958 2125 1964 2126
rect 2062 2130 2068 2131
rect 2062 2126 2063 2130
rect 2067 2126 2068 2130
rect 2062 2125 2068 2126
rect 2158 2130 2164 2131
rect 2158 2126 2159 2130
rect 2163 2126 2164 2130
rect 2158 2125 2164 2126
rect 2254 2130 2260 2131
rect 2254 2126 2255 2130
rect 2259 2126 2260 2130
rect 2254 2125 2260 2126
rect 2350 2130 2356 2131
rect 2350 2126 2351 2130
rect 2355 2126 2356 2130
rect 2350 2125 2356 2126
rect 2446 2130 2452 2131
rect 2446 2126 2447 2130
rect 2451 2126 2452 2130
rect 2446 2125 2452 2126
rect 2542 2130 2548 2131
rect 2542 2126 2543 2130
rect 2547 2126 2548 2130
rect 2542 2125 2548 2126
rect 2584 2122 2586 2137
rect 1366 2121 1372 2122
rect 110 2120 116 2121
rect 1326 2120 1332 2121
rect 110 2116 111 2120
rect 115 2116 116 2120
rect 110 2115 116 2116
rect 182 2119 188 2120
rect 182 2115 183 2119
rect 187 2115 188 2119
rect 112 2091 114 2115
rect 182 2114 188 2115
rect 254 2119 260 2120
rect 254 2115 255 2119
rect 259 2115 260 2119
rect 254 2114 260 2115
rect 334 2119 340 2120
rect 334 2115 335 2119
rect 339 2115 340 2119
rect 334 2114 340 2115
rect 430 2119 436 2120
rect 430 2115 431 2119
rect 435 2115 436 2119
rect 430 2114 436 2115
rect 534 2119 540 2120
rect 534 2115 535 2119
rect 539 2115 540 2119
rect 534 2114 540 2115
rect 646 2119 652 2120
rect 646 2115 647 2119
rect 651 2115 652 2119
rect 646 2114 652 2115
rect 758 2119 764 2120
rect 758 2115 759 2119
rect 763 2115 764 2119
rect 758 2114 764 2115
rect 862 2119 868 2120
rect 862 2115 863 2119
rect 867 2115 868 2119
rect 862 2114 868 2115
rect 966 2119 972 2120
rect 966 2115 967 2119
rect 971 2115 972 2119
rect 966 2114 972 2115
rect 1062 2119 1068 2120
rect 1062 2115 1063 2119
rect 1067 2115 1068 2119
rect 1062 2114 1068 2115
rect 1166 2119 1172 2120
rect 1166 2115 1167 2119
rect 1171 2115 1172 2119
rect 1166 2114 1172 2115
rect 1270 2119 1276 2120
rect 1270 2115 1271 2119
rect 1275 2115 1276 2119
rect 1326 2116 1327 2120
rect 1331 2116 1332 2120
rect 1366 2117 1367 2121
rect 1371 2117 1372 2121
rect 1366 2116 1372 2117
rect 2582 2121 2588 2122
rect 2582 2117 2583 2121
rect 2587 2117 2588 2121
rect 2582 2116 2588 2117
rect 1326 2115 1332 2116
rect 1270 2114 1276 2115
rect 184 2091 186 2114
rect 256 2091 258 2114
rect 336 2091 338 2114
rect 432 2091 434 2114
rect 536 2091 538 2114
rect 648 2091 650 2114
rect 760 2091 762 2114
rect 864 2091 866 2114
rect 968 2091 970 2114
rect 1064 2091 1066 2114
rect 1168 2091 1170 2114
rect 1272 2091 1274 2114
rect 1328 2091 1330 2115
rect 1366 2104 1372 2105
rect 2582 2104 2588 2105
rect 1366 2100 1367 2104
rect 1371 2100 1372 2104
rect 1366 2099 1372 2100
rect 1590 2103 1596 2104
rect 1590 2099 1591 2103
rect 1595 2099 1596 2103
rect 111 2090 115 2091
rect 111 2085 115 2086
rect 143 2090 147 2091
rect 143 2085 147 2086
rect 183 2090 187 2091
rect 183 2085 187 2086
rect 199 2090 203 2091
rect 199 2085 203 2086
rect 255 2090 259 2091
rect 255 2085 259 2086
rect 271 2090 275 2091
rect 271 2085 275 2086
rect 335 2090 339 2091
rect 335 2085 339 2086
rect 367 2090 371 2091
rect 367 2085 371 2086
rect 431 2090 435 2091
rect 431 2085 435 2086
rect 463 2090 467 2091
rect 463 2085 467 2086
rect 535 2090 539 2091
rect 535 2085 539 2086
rect 567 2090 571 2091
rect 567 2085 571 2086
rect 647 2090 651 2091
rect 647 2085 651 2086
rect 663 2090 667 2091
rect 663 2085 667 2086
rect 759 2090 763 2091
rect 759 2085 763 2086
rect 847 2090 851 2091
rect 847 2085 851 2086
rect 863 2090 867 2091
rect 863 2085 867 2086
rect 927 2090 931 2091
rect 927 2085 931 2086
rect 967 2090 971 2091
rect 967 2085 971 2086
rect 1007 2090 1011 2091
rect 1007 2085 1011 2086
rect 1063 2090 1067 2091
rect 1063 2085 1067 2086
rect 1095 2090 1099 2091
rect 1095 2085 1099 2086
rect 1167 2090 1171 2091
rect 1167 2085 1171 2086
rect 1183 2090 1187 2091
rect 1183 2085 1187 2086
rect 1271 2090 1275 2091
rect 1271 2085 1275 2086
rect 1327 2090 1331 2091
rect 1368 2087 1370 2099
rect 1590 2098 1596 2099
rect 1662 2103 1668 2104
rect 1662 2099 1663 2103
rect 1667 2099 1668 2103
rect 1662 2098 1668 2099
rect 1750 2103 1756 2104
rect 1750 2099 1751 2103
rect 1755 2099 1756 2103
rect 1750 2098 1756 2099
rect 1846 2103 1852 2104
rect 1846 2099 1847 2103
rect 1851 2099 1852 2103
rect 1846 2098 1852 2099
rect 1942 2103 1948 2104
rect 1942 2099 1943 2103
rect 1947 2099 1948 2103
rect 1942 2098 1948 2099
rect 2046 2103 2052 2104
rect 2046 2099 2047 2103
rect 2051 2099 2052 2103
rect 2046 2098 2052 2099
rect 2142 2103 2148 2104
rect 2142 2099 2143 2103
rect 2147 2099 2148 2103
rect 2142 2098 2148 2099
rect 2238 2103 2244 2104
rect 2238 2099 2239 2103
rect 2243 2099 2244 2103
rect 2238 2098 2244 2099
rect 2334 2103 2340 2104
rect 2334 2099 2335 2103
rect 2339 2099 2340 2103
rect 2334 2098 2340 2099
rect 2430 2103 2436 2104
rect 2430 2099 2431 2103
rect 2435 2099 2436 2103
rect 2430 2098 2436 2099
rect 2526 2103 2532 2104
rect 2526 2099 2527 2103
rect 2531 2099 2532 2103
rect 2582 2100 2583 2104
rect 2587 2100 2588 2104
rect 2582 2099 2588 2100
rect 2526 2098 2532 2099
rect 1592 2087 1594 2098
rect 1664 2087 1666 2098
rect 1752 2087 1754 2098
rect 1848 2087 1850 2098
rect 1944 2087 1946 2098
rect 2048 2087 2050 2098
rect 2144 2087 2146 2098
rect 2240 2087 2242 2098
rect 2336 2087 2338 2098
rect 2432 2087 2434 2098
rect 2528 2087 2530 2098
rect 2584 2087 2586 2099
rect 1327 2085 1331 2086
rect 1367 2086 1371 2087
rect 112 2073 114 2085
rect 144 2074 146 2085
rect 200 2074 202 2085
rect 272 2074 274 2085
rect 368 2074 370 2085
rect 464 2074 466 2085
rect 568 2074 570 2085
rect 664 2074 666 2085
rect 760 2074 762 2085
rect 848 2074 850 2085
rect 928 2074 930 2085
rect 1008 2074 1010 2085
rect 1096 2074 1098 2085
rect 1184 2074 1186 2085
rect 142 2073 148 2074
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 142 2069 143 2073
rect 147 2069 148 2073
rect 142 2068 148 2069
rect 198 2073 204 2074
rect 198 2069 199 2073
rect 203 2069 204 2073
rect 198 2068 204 2069
rect 270 2073 276 2074
rect 270 2069 271 2073
rect 275 2069 276 2073
rect 270 2068 276 2069
rect 366 2073 372 2074
rect 366 2069 367 2073
rect 371 2069 372 2073
rect 366 2068 372 2069
rect 462 2073 468 2074
rect 462 2069 463 2073
rect 467 2069 468 2073
rect 462 2068 468 2069
rect 566 2073 572 2074
rect 566 2069 567 2073
rect 571 2069 572 2073
rect 566 2068 572 2069
rect 662 2073 668 2074
rect 662 2069 663 2073
rect 667 2069 668 2073
rect 662 2068 668 2069
rect 758 2073 764 2074
rect 758 2069 759 2073
rect 763 2069 764 2073
rect 758 2068 764 2069
rect 846 2073 852 2074
rect 846 2069 847 2073
rect 851 2069 852 2073
rect 846 2068 852 2069
rect 926 2073 932 2074
rect 926 2069 927 2073
rect 931 2069 932 2073
rect 926 2068 932 2069
rect 1006 2073 1012 2074
rect 1006 2069 1007 2073
rect 1011 2069 1012 2073
rect 1006 2068 1012 2069
rect 1094 2073 1100 2074
rect 1094 2069 1095 2073
rect 1099 2069 1100 2073
rect 1094 2068 1100 2069
rect 1182 2073 1188 2074
rect 1328 2073 1330 2085
rect 1367 2081 1371 2082
rect 1487 2086 1491 2087
rect 1487 2081 1491 2082
rect 1583 2086 1587 2087
rect 1583 2081 1587 2082
rect 1591 2086 1595 2087
rect 1591 2081 1595 2082
rect 1663 2086 1667 2087
rect 1663 2081 1667 2082
rect 1679 2086 1683 2087
rect 1679 2081 1683 2082
rect 1751 2086 1755 2087
rect 1751 2081 1755 2082
rect 1783 2086 1787 2087
rect 1783 2081 1787 2082
rect 1847 2086 1851 2087
rect 1847 2081 1851 2082
rect 1887 2086 1891 2087
rect 1887 2081 1891 2082
rect 1943 2086 1947 2087
rect 1943 2081 1947 2082
rect 1983 2086 1987 2087
rect 1983 2081 1987 2082
rect 2047 2086 2051 2087
rect 2047 2081 2051 2082
rect 2079 2086 2083 2087
rect 2079 2081 2083 2082
rect 2143 2086 2147 2087
rect 2143 2081 2147 2082
rect 2167 2086 2171 2087
rect 2167 2081 2171 2082
rect 2239 2086 2243 2087
rect 2239 2081 2243 2082
rect 2255 2086 2259 2087
rect 2255 2081 2259 2082
rect 2335 2086 2339 2087
rect 2335 2081 2339 2082
rect 2343 2086 2347 2087
rect 2343 2081 2347 2082
rect 2431 2086 2435 2087
rect 2431 2081 2435 2082
rect 2439 2086 2443 2087
rect 2439 2081 2443 2082
rect 2527 2086 2531 2087
rect 2527 2081 2531 2082
rect 2583 2086 2587 2087
rect 2583 2081 2587 2082
rect 1182 2069 1183 2073
rect 1187 2069 1188 2073
rect 1182 2068 1188 2069
rect 1326 2072 1332 2073
rect 1326 2068 1327 2072
rect 1331 2068 1332 2072
rect 1368 2069 1370 2081
rect 1488 2070 1490 2081
rect 1584 2070 1586 2081
rect 1680 2070 1682 2081
rect 1784 2070 1786 2081
rect 1888 2070 1890 2081
rect 1984 2070 1986 2081
rect 2080 2070 2082 2081
rect 2168 2070 2170 2081
rect 2256 2070 2258 2081
rect 2344 2070 2346 2081
rect 2440 2070 2442 2081
rect 2528 2070 2530 2081
rect 1486 2069 1492 2070
rect 110 2067 116 2068
rect 1326 2067 1332 2068
rect 1366 2068 1372 2069
rect 1366 2064 1367 2068
rect 1371 2064 1372 2068
rect 1486 2065 1487 2069
rect 1491 2065 1492 2069
rect 1486 2064 1492 2065
rect 1582 2069 1588 2070
rect 1582 2065 1583 2069
rect 1587 2065 1588 2069
rect 1582 2064 1588 2065
rect 1678 2069 1684 2070
rect 1678 2065 1679 2069
rect 1683 2065 1684 2069
rect 1678 2064 1684 2065
rect 1782 2069 1788 2070
rect 1782 2065 1783 2069
rect 1787 2065 1788 2069
rect 1782 2064 1788 2065
rect 1886 2069 1892 2070
rect 1886 2065 1887 2069
rect 1891 2065 1892 2069
rect 1886 2064 1892 2065
rect 1982 2069 1988 2070
rect 1982 2065 1983 2069
rect 1987 2065 1988 2069
rect 1982 2064 1988 2065
rect 2078 2069 2084 2070
rect 2078 2065 2079 2069
rect 2083 2065 2084 2069
rect 2078 2064 2084 2065
rect 2166 2069 2172 2070
rect 2166 2065 2167 2069
rect 2171 2065 2172 2069
rect 2166 2064 2172 2065
rect 2254 2069 2260 2070
rect 2254 2065 2255 2069
rect 2259 2065 2260 2069
rect 2254 2064 2260 2065
rect 2342 2069 2348 2070
rect 2342 2065 2343 2069
rect 2347 2065 2348 2069
rect 2342 2064 2348 2065
rect 2438 2069 2444 2070
rect 2438 2065 2439 2069
rect 2443 2065 2444 2069
rect 2438 2064 2444 2065
rect 2526 2069 2532 2070
rect 2584 2069 2586 2081
rect 2526 2065 2527 2069
rect 2531 2065 2532 2069
rect 2526 2064 2532 2065
rect 2582 2068 2588 2069
rect 2582 2064 2583 2068
rect 2587 2064 2588 2068
rect 1366 2063 1372 2064
rect 2582 2063 2588 2064
rect 110 2055 116 2056
rect 110 2051 111 2055
rect 115 2051 116 2055
rect 110 2050 116 2051
rect 1326 2055 1332 2056
rect 1326 2051 1327 2055
rect 1331 2051 1332 2055
rect 1326 2050 1332 2051
rect 1366 2051 1372 2052
rect 112 2027 114 2050
rect 158 2046 164 2047
rect 158 2042 159 2046
rect 163 2042 164 2046
rect 158 2041 164 2042
rect 214 2046 220 2047
rect 214 2042 215 2046
rect 219 2042 220 2046
rect 214 2041 220 2042
rect 286 2046 292 2047
rect 286 2042 287 2046
rect 291 2042 292 2046
rect 286 2041 292 2042
rect 382 2046 388 2047
rect 382 2042 383 2046
rect 387 2042 388 2046
rect 382 2041 388 2042
rect 478 2046 484 2047
rect 478 2042 479 2046
rect 483 2042 484 2046
rect 478 2041 484 2042
rect 582 2046 588 2047
rect 582 2042 583 2046
rect 587 2042 588 2046
rect 582 2041 588 2042
rect 678 2046 684 2047
rect 678 2042 679 2046
rect 683 2042 684 2046
rect 678 2041 684 2042
rect 774 2046 780 2047
rect 774 2042 775 2046
rect 779 2042 780 2046
rect 774 2041 780 2042
rect 862 2046 868 2047
rect 862 2042 863 2046
rect 867 2042 868 2046
rect 862 2041 868 2042
rect 942 2046 948 2047
rect 942 2042 943 2046
rect 947 2042 948 2046
rect 942 2041 948 2042
rect 1022 2046 1028 2047
rect 1022 2042 1023 2046
rect 1027 2042 1028 2046
rect 1022 2041 1028 2042
rect 1110 2046 1116 2047
rect 1110 2042 1111 2046
rect 1115 2042 1116 2046
rect 1110 2041 1116 2042
rect 1198 2046 1204 2047
rect 1198 2042 1199 2046
rect 1203 2042 1204 2046
rect 1198 2041 1204 2042
rect 160 2027 162 2041
rect 216 2027 218 2041
rect 288 2027 290 2041
rect 384 2027 386 2041
rect 480 2027 482 2041
rect 584 2027 586 2041
rect 680 2027 682 2041
rect 776 2027 778 2041
rect 864 2027 866 2041
rect 944 2027 946 2041
rect 1024 2027 1026 2041
rect 1112 2027 1114 2041
rect 1200 2027 1202 2041
rect 1328 2027 1330 2050
rect 1366 2047 1367 2051
rect 1371 2047 1372 2051
rect 1366 2046 1372 2047
rect 2582 2051 2588 2052
rect 2582 2047 2583 2051
rect 2587 2047 2588 2051
rect 2582 2046 2588 2047
rect 1368 2031 1370 2046
rect 1502 2042 1508 2043
rect 1502 2038 1503 2042
rect 1507 2038 1508 2042
rect 1502 2037 1508 2038
rect 1598 2042 1604 2043
rect 1598 2038 1599 2042
rect 1603 2038 1604 2042
rect 1598 2037 1604 2038
rect 1694 2042 1700 2043
rect 1694 2038 1695 2042
rect 1699 2038 1700 2042
rect 1694 2037 1700 2038
rect 1798 2042 1804 2043
rect 1798 2038 1799 2042
rect 1803 2038 1804 2042
rect 1798 2037 1804 2038
rect 1902 2042 1908 2043
rect 1902 2038 1903 2042
rect 1907 2038 1908 2042
rect 1902 2037 1908 2038
rect 1998 2042 2004 2043
rect 1998 2038 1999 2042
rect 2003 2038 2004 2042
rect 1998 2037 2004 2038
rect 2094 2042 2100 2043
rect 2094 2038 2095 2042
rect 2099 2038 2100 2042
rect 2094 2037 2100 2038
rect 2182 2042 2188 2043
rect 2182 2038 2183 2042
rect 2187 2038 2188 2042
rect 2182 2037 2188 2038
rect 2270 2042 2276 2043
rect 2270 2038 2271 2042
rect 2275 2038 2276 2042
rect 2270 2037 2276 2038
rect 2358 2042 2364 2043
rect 2358 2038 2359 2042
rect 2363 2038 2364 2042
rect 2358 2037 2364 2038
rect 2454 2042 2460 2043
rect 2454 2038 2455 2042
rect 2459 2038 2460 2042
rect 2454 2037 2460 2038
rect 2542 2042 2548 2043
rect 2542 2038 2543 2042
rect 2547 2038 2548 2042
rect 2542 2037 2548 2038
rect 1504 2031 1506 2037
rect 1600 2031 1602 2037
rect 1696 2031 1698 2037
rect 1800 2031 1802 2037
rect 1904 2031 1906 2037
rect 2000 2031 2002 2037
rect 2096 2031 2098 2037
rect 2184 2031 2186 2037
rect 2272 2031 2274 2037
rect 2360 2031 2362 2037
rect 2456 2031 2458 2037
rect 2544 2031 2546 2037
rect 2584 2031 2586 2046
rect 1367 2030 1371 2031
rect 111 2026 115 2027
rect 111 2021 115 2022
rect 159 2026 163 2027
rect 159 2021 163 2022
rect 175 2026 179 2027
rect 175 2021 179 2022
rect 215 2026 219 2027
rect 215 2021 219 2022
rect 239 2026 243 2027
rect 239 2021 243 2022
rect 287 2026 291 2027
rect 287 2021 291 2022
rect 311 2026 315 2027
rect 311 2021 315 2022
rect 383 2026 387 2027
rect 383 2021 387 2022
rect 391 2026 395 2027
rect 391 2021 395 2022
rect 471 2026 475 2027
rect 471 2021 475 2022
rect 479 2026 483 2027
rect 479 2021 483 2022
rect 559 2026 563 2027
rect 559 2021 563 2022
rect 583 2026 587 2027
rect 583 2021 587 2022
rect 647 2026 651 2027
rect 647 2021 651 2022
rect 679 2026 683 2027
rect 679 2021 683 2022
rect 735 2026 739 2027
rect 735 2021 739 2022
rect 775 2026 779 2027
rect 775 2021 779 2022
rect 823 2026 827 2027
rect 823 2021 827 2022
rect 863 2026 867 2027
rect 863 2021 867 2022
rect 911 2026 915 2027
rect 911 2021 915 2022
rect 943 2026 947 2027
rect 943 2021 947 2022
rect 1007 2026 1011 2027
rect 1007 2021 1011 2022
rect 1023 2026 1027 2027
rect 1023 2021 1027 2022
rect 1103 2026 1107 2027
rect 1103 2021 1107 2022
rect 1111 2026 1115 2027
rect 1111 2021 1115 2022
rect 1199 2026 1203 2027
rect 1199 2021 1203 2022
rect 1327 2026 1331 2027
rect 1367 2025 1371 2026
rect 1415 2030 1419 2031
rect 1415 2025 1419 2026
rect 1471 2030 1475 2031
rect 1471 2025 1475 2026
rect 1503 2030 1507 2031
rect 1503 2025 1507 2026
rect 1535 2030 1539 2031
rect 1535 2025 1539 2026
rect 1599 2030 1603 2031
rect 1599 2025 1603 2026
rect 1615 2030 1619 2031
rect 1615 2025 1619 2026
rect 1695 2030 1699 2031
rect 1695 2025 1699 2026
rect 1703 2030 1707 2031
rect 1703 2025 1707 2026
rect 1791 2030 1795 2031
rect 1791 2025 1795 2026
rect 1799 2030 1803 2031
rect 1799 2025 1803 2026
rect 1887 2030 1891 2031
rect 1887 2025 1891 2026
rect 1903 2030 1907 2031
rect 1903 2025 1907 2026
rect 1983 2030 1987 2031
rect 1983 2025 1987 2026
rect 1999 2030 2003 2031
rect 1999 2025 2003 2026
rect 2079 2030 2083 2031
rect 2079 2025 2083 2026
rect 2095 2030 2099 2031
rect 2095 2025 2099 2026
rect 2175 2030 2179 2031
rect 2175 2025 2179 2026
rect 2183 2030 2187 2031
rect 2183 2025 2187 2026
rect 2271 2030 2275 2031
rect 2271 2025 2275 2026
rect 2359 2030 2363 2031
rect 2359 2025 2363 2026
rect 2367 2030 2371 2031
rect 2367 2025 2371 2026
rect 2455 2030 2459 2031
rect 2455 2025 2459 2026
rect 2463 2030 2467 2031
rect 2463 2025 2467 2026
rect 2543 2030 2547 2031
rect 2543 2025 2547 2026
rect 2583 2030 2587 2031
rect 2583 2025 2587 2026
rect 1327 2021 1331 2022
rect 112 2006 114 2021
rect 176 2015 178 2021
rect 240 2015 242 2021
rect 312 2015 314 2021
rect 392 2015 394 2021
rect 472 2015 474 2021
rect 560 2015 562 2021
rect 648 2015 650 2021
rect 736 2015 738 2021
rect 824 2015 826 2021
rect 912 2015 914 2021
rect 1008 2015 1010 2021
rect 1104 2015 1106 2021
rect 174 2014 180 2015
rect 174 2010 175 2014
rect 179 2010 180 2014
rect 174 2009 180 2010
rect 238 2014 244 2015
rect 238 2010 239 2014
rect 243 2010 244 2014
rect 238 2009 244 2010
rect 310 2014 316 2015
rect 310 2010 311 2014
rect 315 2010 316 2014
rect 310 2009 316 2010
rect 390 2014 396 2015
rect 390 2010 391 2014
rect 395 2010 396 2014
rect 390 2009 396 2010
rect 470 2014 476 2015
rect 470 2010 471 2014
rect 475 2010 476 2014
rect 470 2009 476 2010
rect 558 2014 564 2015
rect 558 2010 559 2014
rect 563 2010 564 2014
rect 558 2009 564 2010
rect 646 2014 652 2015
rect 646 2010 647 2014
rect 651 2010 652 2014
rect 646 2009 652 2010
rect 734 2014 740 2015
rect 734 2010 735 2014
rect 739 2010 740 2014
rect 734 2009 740 2010
rect 822 2014 828 2015
rect 822 2010 823 2014
rect 827 2010 828 2014
rect 822 2009 828 2010
rect 910 2014 916 2015
rect 910 2010 911 2014
rect 915 2010 916 2014
rect 910 2009 916 2010
rect 1006 2014 1012 2015
rect 1006 2010 1007 2014
rect 1011 2010 1012 2014
rect 1006 2009 1012 2010
rect 1102 2014 1108 2015
rect 1102 2010 1103 2014
rect 1107 2010 1108 2014
rect 1102 2009 1108 2010
rect 1328 2006 1330 2021
rect 1368 2010 1370 2025
rect 1416 2019 1418 2025
rect 1472 2019 1474 2025
rect 1536 2019 1538 2025
rect 1616 2019 1618 2025
rect 1704 2019 1706 2025
rect 1792 2019 1794 2025
rect 1888 2019 1890 2025
rect 1984 2019 1986 2025
rect 2080 2019 2082 2025
rect 2176 2019 2178 2025
rect 2272 2019 2274 2025
rect 2368 2019 2370 2025
rect 2464 2019 2466 2025
rect 2544 2019 2546 2025
rect 1414 2018 1420 2019
rect 1414 2014 1415 2018
rect 1419 2014 1420 2018
rect 1414 2013 1420 2014
rect 1470 2018 1476 2019
rect 1470 2014 1471 2018
rect 1475 2014 1476 2018
rect 1470 2013 1476 2014
rect 1534 2018 1540 2019
rect 1534 2014 1535 2018
rect 1539 2014 1540 2018
rect 1534 2013 1540 2014
rect 1614 2018 1620 2019
rect 1614 2014 1615 2018
rect 1619 2014 1620 2018
rect 1614 2013 1620 2014
rect 1702 2018 1708 2019
rect 1702 2014 1703 2018
rect 1707 2014 1708 2018
rect 1702 2013 1708 2014
rect 1790 2018 1796 2019
rect 1790 2014 1791 2018
rect 1795 2014 1796 2018
rect 1790 2013 1796 2014
rect 1886 2018 1892 2019
rect 1886 2014 1887 2018
rect 1891 2014 1892 2018
rect 1886 2013 1892 2014
rect 1982 2018 1988 2019
rect 1982 2014 1983 2018
rect 1987 2014 1988 2018
rect 1982 2013 1988 2014
rect 2078 2018 2084 2019
rect 2078 2014 2079 2018
rect 2083 2014 2084 2018
rect 2078 2013 2084 2014
rect 2174 2018 2180 2019
rect 2174 2014 2175 2018
rect 2179 2014 2180 2018
rect 2174 2013 2180 2014
rect 2270 2018 2276 2019
rect 2270 2014 2271 2018
rect 2275 2014 2276 2018
rect 2270 2013 2276 2014
rect 2366 2018 2372 2019
rect 2366 2014 2367 2018
rect 2371 2014 2372 2018
rect 2366 2013 2372 2014
rect 2462 2018 2468 2019
rect 2462 2014 2463 2018
rect 2467 2014 2468 2018
rect 2462 2013 2468 2014
rect 2542 2018 2548 2019
rect 2542 2014 2543 2018
rect 2547 2014 2548 2018
rect 2542 2013 2548 2014
rect 2584 2010 2586 2025
rect 1366 2009 1372 2010
rect 110 2005 116 2006
rect 110 2001 111 2005
rect 115 2001 116 2005
rect 110 2000 116 2001
rect 1326 2005 1332 2006
rect 1326 2001 1327 2005
rect 1331 2001 1332 2005
rect 1366 2005 1367 2009
rect 1371 2005 1372 2009
rect 1366 2004 1372 2005
rect 2582 2009 2588 2010
rect 2582 2005 2583 2009
rect 2587 2005 2588 2009
rect 2582 2004 2588 2005
rect 1326 2000 1332 2001
rect 1366 1992 1372 1993
rect 2582 1992 2588 1993
rect 110 1988 116 1989
rect 1326 1988 1332 1989
rect 110 1984 111 1988
rect 115 1984 116 1988
rect 110 1983 116 1984
rect 158 1987 164 1988
rect 158 1983 159 1987
rect 163 1983 164 1987
rect 112 1971 114 1983
rect 158 1982 164 1983
rect 222 1987 228 1988
rect 222 1983 223 1987
rect 227 1983 228 1987
rect 222 1982 228 1983
rect 294 1987 300 1988
rect 294 1983 295 1987
rect 299 1983 300 1987
rect 294 1982 300 1983
rect 374 1987 380 1988
rect 374 1983 375 1987
rect 379 1983 380 1987
rect 374 1982 380 1983
rect 454 1987 460 1988
rect 454 1983 455 1987
rect 459 1983 460 1987
rect 454 1982 460 1983
rect 542 1987 548 1988
rect 542 1983 543 1987
rect 547 1983 548 1987
rect 542 1982 548 1983
rect 630 1987 636 1988
rect 630 1983 631 1987
rect 635 1983 636 1987
rect 630 1982 636 1983
rect 718 1987 724 1988
rect 718 1983 719 1987
rect 723 1983 724 1987
rect 718 1982 724 1983
rect 806 1987 812 1988
rect 806 1983 807 1987
rect 811 1983 812 1987
rect 806 1982 812 1983
rect 894 1987 900 1988
rect 894 1983 895 1987
rect 899 1983 900 1987
rect 894 1982 900 1983
rect 990 1987 996 1988
rect 990 1983 991 1987
rect 995 1983 996 1987
rect 990 1982 996 1983
rect 1086 1987 1092 1988
rect 1086 1983 1087 1987
rect 1091 1983 1092 1987
rect 1326 1984 1327 1988
rect 1331 1984 1332 1988
rect 1366 1988 1367 1992
rect 1371 1988 1372 1992
rect 1366 1987 1372 1988
rect 1398 1991 1404 1992
rect 1398 1987 1399 1991
rect 1403 1987 1404 1991
rect 1326 1983 1332 1984
rect 1086 1982 1092 1983
rect 160 1971 162 1982
rect 224 1971 226 1982
rect 296 1971 298 1982
rect 376 1971 378 1982
rect 456 1971 458 1982
rect 544 1971 546 1982
rect 632 1971 634 1982
rect 720 1971 722 1982
rect 808 1971 810 1982
rect 896 1971 898 1982
rect 992 1971 994 1982
rect 1088 1971 1090 1982
rect 1328 1971 1330 1983
rect 1368 1971 1370 1987
rect 1398 1986 1404 1987
rect 1454 1991 1460 1992
rect 1454 1987 1455 1991
rect 1459 1987 1460 1991
rect 1454 1986 1460 1987
rect 1518 1991 1524 1992
rect 1518 1987 1519 1991
rect 1523 1987 1524 1991
rect 1518 1986 1524 1987
rect 1598 1991 1604 1992
rect 1598 1987 1599 1991
rect 1603 1987 1604 1991
rect 1598 1986 1604 1987
rect 1686 1991 1692 1992
rect 1686 1987 1687 1991
rect 1691 1987 1692 1991
rect 1686 1986 1692 1987
rect 1774 1991 1780 1992
rect 1774 1987 1775 1991
rect 1779 1987 1780 1991
rect 1774 1986 1780 1987
rect 1870 1991 1876 1992
rect 1870 1987 1871 1991
rect 1875 1987 1876 1991
rect 1870 1986 1876 1987
rect 1966 1991 1972 1992
rect 1966 1987 1967 1991
rect 1971 1987 1972 1991
rect 1966 1986 1972 1987
rect 2062 1991 2068 1992
rect 2062 1987 2063 1991
rect 2067 1987 2068 1991
rect 2062 1986 2068 1987
rect 2158 1991 2164 1992
rect 2158 1987 2159 1991
rect 2163 1987 2164 1991
rect 2158 1986 2164 1987
rect 2254 1991 2260 1992
rect 2254 1987 2255 1991
rect 2259 1987 2260 1991
rect 2254 1986 2260 1987
rect 2350 1991 2356 1992
rect 2350 1987 2351 1991
rect 2355 1987 2356 1991
rect 2350 1986 2356 1987
rect 2446 1991 2452 1992
rect 2446 1987 2447 1991
rect 2451 1987 2452 1991
rect 2446 1986 2452 1987
rect 2526 1991 2532 1992
rect 2526 1987 2527 1991
rect 2531 1987 2532 1991
rect 2582 1988 2583 1992
rect 2587 1988 2588 1992
rect 2582 1987 2588 1988
rect 2526 1986 2532 1987
rect 1400 1971 1402 1986
rect 1456 1971 1458 1986
rect 1520 1971 1522 1986
rect 1600 1971 1602 1986
rect 1688 1971 1690 1986
rect 1776 1971 1778 1986
rect 1872 1971 1874 1986
rect 1968 1971 1970 1986
rect 2064 1971 2066 1986
rect 2160 1971 2162 1986
rect 2256 1971 2258 1986
rect 2352 1971 2354 1986
rect 2448 1971 2450 1986
rect 2528 1971 2530 1986
rect 2584 1971 2586 1987
rect 111 1970 115 1971
rect 111 1965 115 1966
rect 159 1970 163 1971
rect 159 1965 163 1966
rect 223 1970 227 1971
rect 223 1965 227 1966
rect 295 1970 299 1971
rect 295 1965 299 1966
rect 375 1970 379 1971
rect 375 1965 379 1966
rect 383 1970 387 1971
rect 383 1965 387 1966
rect 439 1970 443 1971
rect 439 1965 443 1966
rect 455 1970 459 1971
rect 455 1965 459 1966
rect 495 1970 499 1971
rect 495 1965 499 1966
rect 543 1970 547 1971
rect 543 1965 547 1966
rect 551 1970 555 1971
rect 551 1965 555 1966
rect 607 1970 611 1971
rect 607 1965 611 1966
rect 631 1970 635 1971
rect 631 1965 635 1966
rect 671 1970 675 1971
rect 671 1965 675 1966
rect 719 1970 723 1971
rect 719 1965 723 1966
rect 735 1970 739 1971
rect 735 1965 739 1966
rect 807 1970 811 1971
rect 807 1965 811 1966
rect 879 1970 883 1971
rect 879 1965 883 1966
rect 895 1970 899 1971
rect 895 1965 899 1966
rect 951 1970 955 1971
rect 951 1965 955 1966
rect 991 1970 995 1971
rect 991 1965 995 1966
rect 1023 1970 1027 1971
rect 1023 1965 1027 1966
rect 1087 1970 1091 1971
rect 1087 1965 1091 1966
rect 1327 1970 1331 1971
rect 1327 1965 1331 1966
rect 1367 1970 1371 1971
rect 1367 1965 1371 1966
rect 1399 1970 1403 1971
rect 1399 1965 1403 1966
rect 1455 1970 1459 1971
rect 1455 1965 1459 1966
rect 1519 1970 1523 1971
rect 1519 1965 1523 1966
rect 1599 1970 1603 1971
rect 1599 1965 1603 1966
rect 1679 1970 1683 1971
rect 1679 1965 1683 1966
rect 1687 1970 1691 1971
rect 1687 1965 1691 1966
rect 1759 1970 1763 1971
rect 1759 1965 1763 1966
rect 1775 1970 1779 1971
rect 1775 1965 1779 1966
rect 1855 1970 1859 1971
rect 1855 1965 1859 1966
rect 1871 1970 1875 1971
rect 1871 1965 1875 1966
rect 1967 1970 1971 1971
rect 1967 1965 1971 1966
rect 2063 1970 2067 1971
rect 2063 1965 2067 1966
rect 2095 1970 2099 1971
rect 2095 1965 2099 1966
rect 2159 1970 2163 1971
rect 2159 1965 2163 1966
rect 2239 1970 2243 1971
rect 2239 1965 2243 1966
rect 2255 1970 2259 1971
rect 2255 1965 2259 1966
rect 2351 1970 2355 1971
rect 2351 1965 2355 1966
rect 2391 1970 2395 1971
rect 2391 1965 2395 1966
rect 2447 1970 2451 1971
rect 2447 1965 2451 1966
rect 2527 1970 2531 1971
rect 2527 1965 2531 1966
rect 2583 1970 2587 1971
rect 2583 1965 2587 1966
rect 112 1953 114 1965
rect 384 1954 386 1965
rect 440 1954 442 1965
rect 496 1954 498 1965
rect 552 1954 554 1965
rect 608 1954 610 1965
rect 672 1954 674 1965
rect 736 1954 738 1965
rect 808 1954 810 1965
rect 880 1954 882 1965
rect 952 1954 954 1965
rect 1024 1954 1026 1965
rect 382 1953 388 1954
rect 110 1952 116 1953
rect 110 1948 111 1952
rect 115 1948 116 1952
rect 382 1949 383 1953
rect 387 1949 388 1953
rect 382 1948 388 1949
rect 438 1953 444 1954
rect 438 1949 439 1953
rect 443 1949 444 1953
rect 438 1948 444 1949
rect 494 1953 500 1954
rect 494 1949 495 1953
rect 499 1949 500 1953
rect 494 1948 500 1949
rect 550 1953 556 1954
rect 550 1949 551 1953
rect 555 1949 556 1953
rect 550 1948 556 1949
rect 606 1953 612 1954
rect 606 1949 607 1953
rect 611 1949 612 1953
rect 606 1948 612 1949
rect 670 1953 676 1954
rect 670 1949 671 1953
rect 675 1949 676 1953
rect 670 1948 676 1949
rect 734 1953 740 1954
rect 734 1949 735 1953
rect 739 1949 740 1953
rect 734 1948 740 1949
rect 806 1953 812 1954
rect 806 1949 807 1953
rect 811 1949 812 1953
rect 806 1948 812 1949
rect 878 1953 884 1954
rect 878 1949 879 1953
rect 883 1949 884 1953
rect 878 1948 884 1949
rect 950 1953 956 1954
rect 950 1949 951 1953
rect 955 1949 956 1953
rect 950 1948 956 1949
rect 1022 1953 1028 1954
rect 1328 1953 1330 1965
rect 1368 1953 1370 1965
rect 1400 1954 1402 1965
rect 1456 1954 1458 1965
rect 1520 1954 1522 1965
rect 1600 1954 1602 1965
rect 1680 1954 1682 1965
rect 1760 1954 1762 1965
rect 1856 1954 1858 1965
rect 1968 1954 1970 1965
rect 2096 1954 2098 1965
rect 2240 1954 2242 1965
rect 2392 1954 2394 1965
rect 2528 1954 2530 1965
rect 1398 1953 1404 1954
rect 1022 1949 1023 1953
rect 1027 1949 1028 1953
rect 1022 1948 1028 1949
rect 1326 1952 1332 1953
rect 1326 1948 1327 1952
rect 1331 1948 1332 1952
rect 110 1947 116 1948
rect 1326 1947 1332 1948
rect 1366 1952 1372 1953
rect 1366 1948 1367 1952
rect 1371 1948 1372 1952
rect 1398 1949 1399 1953
rect 1403 1949 1404 1953
rect 1398 1948 1404 1949
rect 1454 1953 1460 1954
rect 1454 1949 1455 1953
rect 1459 1949 1460 1953
rect 1454 1948 1460 1949
rect 1518 1953 1524 1954
rect 1518 1949 1519 1953
rect 1523 1949 1524 1953
rect 1518 1948 1524 1949
rect 1598 1953 1604 1954
rect 1598 1949 1599 1953
rect 1603 1949 1604 1953
rect 1598 1948 1604 1949
rect 1678 1953 1684 1954
rect 1678 1949 1679 1953
rect 1683 1949 1684 1953
rect 1678 1948 1684 1949
rect 1758 1953 1764 1954
rect 1758 1949 1759 1953
rect 1763 1949 1764 1953
rect 1758 1948 1764 1949
rect 1854 1953 1860 1954
rect 1854 1949 1855 1953
rect 1859 1949 1860 1953
rect 1854 1948 1860 1949
rect 1966 1953 1972 1954
rect 1966 1949 1967 1953
rect 1971 1949 1972 1953
rect 1966 1948 1972 1949
rect 2094 1953 2100 1954
rect 2094 1949 2095 1953
rect 2099 1949 2100 1953
rect 2094 1948 2100 1949
rect 2238 1953 2244 1954
rect 2238 1949 2239 1953
rect 2243 1949 2244 1953
rect 2238 1948 2244 1949
rect 2390 1953 2396 1954
rect 2390 1949 2391 1953
rect 2395 1949 2396 1953
rect 2390 1948 2396 1949
rect 2526 1953 2532 1954
rect 2584 1953 2586 1965
rect 2526 1949 2527 1953
rect 2531 1949 2532 1953
rect 2526 1948 2532 1949
rect 2582 1952 2588 1953
rect 2582 1948 2583 1952
rect 2587 1948 2588 1952
rect 1366 1947 1372 1948
rect 2582 1947 2588 1948
rect 110 1935 116 1936
rect 110 1931 111 1935
rect 115 1931 116 1935
rect 110 1930 116 1931
rect 1326 1935 1332 1936
rect 1326 1931 1327 1935
rect 1331 1931 1332 1935
rect 1326 1930 1332 1931
rect 1366 1935 1372 1936
rect 1366 1931 1367 1935
rect 1371 1931 1372 1935
rect 1366 1930 1372 1931
rect 2582 1935 2588 1936
rect 2582 1931 2583 1935
rect 2587 1931 2588 1935
rect 2582 1930 2588 1931
rect 112 1915 114 1930
rect 398 1926 404 1927
rect 398 1922 399 1926
rect 403 1922 404 1926
rect 398 1921 404 1922
rect 454 1926 460 1927
rect 454 1922 455 1926
rect 459 1922 460 1926
rect 454 1921 460 1922
rect 510 1926 516 1927
rect 510 1922 511 1926
rect 515 1922 516 1926
rect 510 1921 516 1922
rect 566 1926 572 1927
rect 566 1922 567 1926
rect 571 1922 572 1926
rect 566 1921 572 1922
rect 622 1926 628 1927
rect 622 1922 623 1926
rect 627 1922 628 1926
rect 622 1921 628 1922
rect 686 1926 692 1927
rect 686 1922 687 1926
rect 691 1922 692 1926
rect 686 1921 692 1922
rect 750 1926 756 1927
rect 750 1922 751 1926
rect 755 1922 756 1926
rect 750 1921 756 1922
rect 822 1926 828 1927
rect 822 1922 823 1926
rect 827 1922 828 1926
rect 822 1921 828 1922
rect 894 1926 900 1927
rect 894 1922 895 1926
rect 899 1922 900 1926
rect 894 1921 900 1922
rect 966 1926 972 1927
rect 966 1922 967 1926
rect 971 1922 972 1926
rect 966 1921 972 1922
rect 1038 1926 1044 1927
rect 1038 1922 1039 1926
rect 1043 1922 1044 1926
rect 1038 1921 1044 1922
rect 400 1915 402 1921
rect 456 1915 458 1921
rect 512 1915 514 1921
rect 568 1915 570 1921
rect 624 1915 626 1921
rect 688 1915 690 1921
rect 752 1915 754 1921
rect 824 1915 826 1921
rect 896 1915 898 1921
rect 968 1915 970 1921
rect 1040 1915 1042 1921
rect 1328 1915 1330 1930
rect 1368 1915 1370 1930
rect 1414 1926 1420 1927
rect 1414 1922 1415 1926
rect 1419 1922 1420 1926
rect 1414 1921 1420 1922
rect 1470 1926 1476 1927
rect 1470 1922 1471 1926
rect 1475 1922 1476 1926
rect 1470 1921 1476 1922
rect 1534 1926 1540 1927
rect 1534 1922 1535 1926
rect 1539 1922 1540 1926
rect 1534 1921 1540 1922
rect 1614 1926 1620 1927
rect 1614 1922 1615 1926
rect 1619 1922 1620 1926
rect 1614 1921 1620 1922
rect 1694 1926 1700 1927
rect 1694 1922 1695 1926
rect 1699 1922 1700 1926
rect 1694 1921 1700 1922
rect 1774 1926 1780 1927
rect 1774 1922 1775 1926
rect 1779 1922 1780 1926
rect 1774 1921 1780 1922
rect 1870 1926 1876 1927
rect 1870 1922 1871 1926
rect 1875 1922 1876 1926
rect 1870 1921 1876 1922
rect 1982 1926 1988 1927
rect 1982 1922 1983 1926
rect 1987 1922 1988 1926
rect 1982 1921 1988 1922
rect 2110 1926 2116 1927
rect 2110 1922 2111 1926
rect 2115 1922 2116 1926
rect 2110 1921 2116 1922
rect 2254 1926 2260 1927
rect 2254 1922 2255 1926
rect 2259 1922 2260 1926
rect 2254 1921 2260 1922
rect 2406 1926 2412 1927
rect 2406 1922 2407 1926
rect 2411 1922 2412 1926
rect 2406 1921 2412 1922
rect 2542 1926 2548 1927
rect 2542 1922 2543 1926
rect 2547 1922 2548 1926
rect 2542 1921 2548 1922
rect 1416 1915 1418 1921
rect 1472 1915 1474 1921
rect 1536 1915 1538 1921
rect 1616 1915 1618 1921
rect 1696 1915 1698 1921
rect 1776 1915 1778 1921
rect 1872 1915 1874 1921
rect 1984 1915 1986 1921
rect 2112 1915 2114 1921
rect 2256 1915 2258 1921
rect 2408 1915 2410 1921
rect 2544 1915 2546 1921
rect 2584 1915 2586 1930
rect 111 1914 115 1915
rect 111 1909 115 1910
rect 399 1914 403 1915
rect 399 1909 403 1910
rect 455 1914 459 1915
rect 455 1909 459 1910
rect 511 1914 515 1915
rect 511 1909 515 1910
rect 519 1914 523 1915
rect 519 1909 523 1910
rect 567 1914 571 1915
rect 567 1909 571 1910
rect 575 1914 579 1915
rect 575 1909 579 1910
rect 623 1914 627 1915
rect 623 1909 627 1910
rect 631 1914 635 1915
rect 631 1909 635 1910
rect 687 1914 691 1915
rect 687 1909 691 1910
rect 743 1914 747 1915
rect 743 1909 747 1910
rect 751 1914 755 1915
rect 751 1909 755 1910
rect 807 1914 811 1915
rect 807 1909 811 1910
rect 823 1914 827 1915
rect 823 1909 827 1910
rect 871 1914 875 1915
rect 871 1909 875 1910
rect 895 1914 899 1915
rect 895 1909 899 1910
rect 935 1914 939 1915
rect 935 1909 939 1910
rect 967 1914 971 1915
rect 967 1909 971 1910
rect 999 1914 1003 1915
rect 999 1909 1003 1910
rect 1039 1914 1043 1915
rect 1039 1909 1043 1910
rect 1327 1914 1331 1915
rect 1327 1909 1331 1910
rect 1367 1914 1371 1915
rect 1367 1909 1371 1910
rect 1415 1914 1419 1915
rect 1415 1909 1419 1910
rect 1471 1914 1475 1915
rect 1471 1909 1475 1910
rect 1535 1914 1539 1915
rect 1535 1909 1539 1910
rect 1575 1914 1579 1915
rect 1575 1909 1579 1910
rect 1615 1914 1619 1915
rect 1615 1909 1619 1910
rect 1631 1914 1635 1915
rect 1631 1909 1635 1910
rect 1687 1914 1691 1915
rect 1687 1909 1691 1910
rect 1695 1914 1699 1915
rect 1695 1909 1699 1910
rect 1743 1914 1747 1915
rect 1743 1909 1747 1910
rect 1775 1914 1779 1915
rect 1775 1909 1779 1910
rect 1799 1914 1803 1915
rect 1799 1909 1803 1910
rect 1855 1914 1859 1915
rect 1855 1909 1859 1910
rect 1871 1914 1875 1915
rect 1871 1909 1875 1910
rect 1927 1914 1931 1915
rect 1927 1909 1931 1910
rect 1983 1914 1987 1915
rect 1983 1909 1987 1910
rect 2015 1914 2019 1915
rect 2015 1909 2019 1910
rect 2111 1914 2115 1915
rect 2111 1909 2115 1910
rect 2127 1914 2131 1915
rect 2127 1909 2131 1910
rect 2247 1914 2251 1915
rect 2247 1909 2251 1910
rect 2255 1914 2259 1915
rect 2255 1909 2259 1910
rect 2383 1914 2387 1915
rect 2383 1909 2387 1910
rect 2407 1914 2411 1915
rect 2407 1909 2411 1910
rect 2519 1914 2523 1915
rect 2519 1909 2523 1910
rect 2543 1914 2547 1915
rect 2543 1909 2547 1910
rect 2583 1914 2587 1915
rect 2583 1909 2587 1910
rect 112 1894 114 1909
rect 520 1903 522 1909
rect 576 1903 578 1909
rect 632 1903 634 1909
rect 688 1903 690 1909
rect 744 1903 746 1909
rect 808 1903 810 1909
rect 872 1903 874 1909
rect 936 1903 938 1909
rect 1000 1903 1002 1909
rect 518 1902 524 1903
rect 518 1898 519 1902
rect 523 1898 524 1902
rect 518 1897 524 1898
rect 574 1902 580 1903
rect 574 1898 575 1902
rect 579 1898 580 1902
rect 574 1897 580 1898
rect 630 1902 636 1903
rect 630 1898 631 1902
rect 635 1898 636 1902
rect 630 1897 636 1898
rect 686 1902 692 1903
rect 686 1898 687 1902
rect 691 1898 692 1902
rect 686 1897 692 1898
rect 742 1902 748 1903
rect 742 1898 743 1902
rect 747 1898 748 1902
rect 742 1897 748 1898
rect 806 1902 812 1903
rect 806 1898 807 1902
rect 811 1898 812 1902
rect 806 1897 812 1898
rect 870 1902 876 1903
rect 870 1898 871 1902
rect 875 1898 876 1902
rect 870 1897 876 1898
rect 934 1902 940 1903
rect 934 1898 935 1902
rect 939 1898 940 1902
rect 934 1897 940 1898
rect 998 1902 1004 1903
rect 998 1898 999 1902
rect 1003 1898 1004 1902
rect 998 1897 1004 1898
rect 1328 1894 1330 1909
rect 1368 1894 1370 1909
rect 1576 1903 1578 1909
rect 1632 1903 1634 1909
rect 1688 1903 1690 1909
rect 1744 1903 1746 1909
rect 1800 1903 1802 1909
rect 1856 1903 1858 1909
rect 1928 1903 1930 1909
rect 2016 1903 2018 1909
rect 2128 1903 2130 1909
rect 2248 1903 2250 1909
rect 2384 1903 2386 1909
rect 2520 1903 2522 1909
rect 1574 1902 1580 1903
rect 1574 1898 1575 1902
rect 1579 1898 1580 1902
rect 1574 1897 1580 1898
rect 1630 1902 1636 1903
rect 1630 1898 1631 1902
rect 1635 1898 1636 1902
rect 1630 1897 1636 1898
rect 1686 1902 1692 1903
rect 1686 1898 1687 1902
rect 1691 1898 1692 1902
rect 1686 1897 1692 1898
rect 1742 1902 1748 1903
rect 1742 1898 1743 1902
rect 1747 1898 1748 1902
rect 1742 1897 1748 1898
rect 1798 1902 1804 1903
rect 1798 1898 1799 1902
rect 1803 1898 1804 1902
rect 1798 1897 1804 1898
rect 1854 1902 1860 1903
rect 1854 1898 1855 1902
rect 1859 1898 1860 1902
rect 1854 1897 1860 1898
rect 1926 1902 1932 1903
rect 1926 1898 1927 1902
rect 1931 1898 1932 1902
rect 1926 1897 1932 1898
rect 2014 1902 2020 1903
rect 2014 1898 2015 1902
rect 2019 1898 2020 1902
rect 2014 1897 2020 1898
rect 2126 1902 2132 1903
rect 2126 1898 2127 1902
rect 2131 1898 2132 1902
rect 2126 1897 2132 1898
rect 2246 1902 2252 1903
rect 2246 1898 2247 1902
rect 2251 1898 2252 1902
rect 2246 1897 2252 1898
rect 2382 1902 2388 1903
rect 2382 1898 2383 1902
rect 2387 1898 2388 1902
rect 2382 1897 2388 1898
rect 2518 1902 2524 1903
rect 2518 1898 2519 1902
rect 2523 1898 2524 1902
rect 2518 1897 2524 1898
rect 2584 1894 2586 1909
rect 110 1893 116 1894
rect 110 1889 111 1893
rect 115 1889 116 1893
rect 110 1888 116 1889
rect 1326 1893 1332 1894
rect 1326 1889 1327 1893
rect 1331 1889 1332 1893
rect 1326 1888 1332 1889
rect 1366 1893 1372 1894
rect 1366 1889 1367 1893
rect 1371 1889 1372 1893
rect 1366 1888 1372 1889
rect 2582 1893 2588 1894
rect 2582 1889 2583 1893
rect 2587 1889 2588 1893
rect 2582 1888 2588 1889
rect 110 1876 116 1877
rect 1326 1876 1332 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 502 1875 508 1876
rect 502 1871 503 1875
rect 507 1871 508 1875
rect 112 1855 114 1871
rect 502 1870 508 1871
rect 558 1875 564 1876
rect 558 1871 559 1875
rect 563 1871 564 1875
rect 558 1870 564 1871
rect 614 1875 620 1876
rect 614 1871 615 1875
rect 619 1871 620 1875
rect 614 1870 620 1871
rect 670 1875 676 1876
rect 670 1871 671 1875
rect 675 1871 676 1875
rect 670 1870 676 1871
rect 726 1875 732 1876
rect 726 1871 727 1875
rect 731 1871 732 1875
rect 726 1870 732 1871
rect 790 1875 796 1876
rect 790 1871 791 1875
rect 795 1871 796 1875
rect 790 1870 796 1871
rect 854 1875 860 1876
rect 854 1871 855 1875
rect 859 1871 860 1875
rect 854 1870 860 1871
rect 918 1875 924 1876
rect 918 1871 919 1875
rect 923 1871 924 1875
rect 918 1870 924 1871
rect 982 1875 988 1876
rect 982 1871 983 1875
rect 987 1871 988 1875
rect 1326 1872 1327 1876
rect 1331 1872 1332 1876
rect 1326 1871 1332 1872
rect 1366 1876 1372 1877
rect 2582 1876 2588 1877
rect 1366 1872 1367 1876
rect 1371 1872 1372 1876
rect 1366 1871 1372 1872
rect 1558 1875 1564 1876
rect 1558 1871 1559 1875
rect 1563 1871 1564 1875
rect 982 1870 988 1871
rect 504 1855 506 1870
rect 560 1855 562 1870
rect 616 1855 618 1870
rect 672 1855 674 1870
rect 728 1855 730 1870
rect 792 1855 794 1870
rect 856 1855 858 1870
rect 920 1855 922 1870
rect 984 1855 986 1870
rect 1328 1855 1330 1871
rect 111 1854 115 1855
rect 111 1849 115 1850
rect 143 1854 147 1855
rect 143 1849 147 1850
rect 199 1854 203 1855
rect 199 1849 203 1850
rect 255 1854 259 1855
rect 255 1849 259 1850
rect 311 1854 315 1855
rect 311 1849 315 1850
rect 375 1854 379 1855
rect 375 1849 379 1850
rect 455 1854 459 1855
rect 455 1849 459 1850
rect 503 1854 507 1855
rect 503 1849 507 1850
rect 543 1854 547 1855
rect 543 1849 547 1850
rect 559 1854 563 1855
rect 559 1849 563 1850
rect 615 1854 619 1855
rect 615 1849 619 1850
rect 631 1854 635 1855
rect 631 1849 635 1850
rect 671 1854 675 1855
rect 671 1849 675 1850
rect 719 1854 723 1855
rect 719 1849 723 1850
rect 727 1854 731 1855
rect 727 1849 731 1850
rect 791 1854 795 1855
rect 791 1849 795 1850
rect 799 1854 803 1855
rect 799 1849 803 1850
rect 855 1854 859 1855
rect 855 1849 859 1850
rect 887 1854 891 1855
rect 887 1849 891 1850
rect 919 1854 923 1855
rect 919 1849 923 1850
rect 975 1854 979 1855
rect 975 1849 979 1850
rect 983 1854 987 1855
rect 983 1849 987 1850
rect 1063 1854 1067 1855
rect 1063 1849 1067 1850
rect 1327 1854 1331 1855
rect 1368 1851 1370 1871
rect 1558 1870 1564 1871
rect 1614 1875 1620 1876
rect 1614 1871 1615 1875
rect 1619 1871 1620 1875
rect 1614 1870 1620 1871
rect 1670 1875 1676 1876
rect 1670 1871 1671 1875
rect 1675 1871 1676 1875
rect 1670 1870 1676 1871
rect 1726 1875 1732 1876
rect 1726 1871 1727 1875
rect 1731 1871 1732 1875
rect 1726 1870 1732 1871
rect 1782 1875 1788 1876
rect 1782 1871 1783 1875
rect 1787 1871 1788 1875
rect 1782 1870 1788 1871
rect 1838 1875 1844 1876
rect 1838 1871 1839 1875
rect 1843 1871 1844 1875
rect 1838 1870 1844 1871
rect 1910 1875 1916 1876
rect 1910 1871 1911 1875
rect 1915 1871 1916 1875
rect 1910 1870 1916 1871
rect 1998 1875 2004 1876
rect 1998 1871 1999 1875
rect 2003 1871 2004 1875
rect 1998 1870 2004 1871
rect 2110 1875 2116 1876
rect 2110 1871 2111 1875
rect 2115 1871 2116 1875
rect 2110 1870 2116 1871
rect 2230 1875 2236 1876
rect 2230 1871 2231 1875
rect 2235 1871 2236 1875
rect 2230 1870 2236 1871
rect 2366 1875 2372 1876
rect 2366 1871 2367 1875
rect 2371 1871 2372 1875
rect 2366 1870 2372 1871
rect 2502 1875 2508 1876
rect 2502 1871 2503 1875
rect 2507 1871 2508 1875
rect 2582 1872 2583 1876
rect 2587 1872 2588 1876
rect 2582 1871 2588 1872
rect 2502 1870 2508 1871
rect 1560 1851 1562 1870
rect 1616 1851 1618 1870
rect 1672 1851 1674 1870
rect 1728 1851 1730 1870
rect 1784 1851 1786 1870
rect 1840 1851 1842 1870
rect 1912 1851 1914 1870
rect 2000 1851 2002 1870
rect 2112 1851 2114 1870
rect 2232 1851 2234 1870
rect 2368 1851 2370 1870
rect 2504 1851 2506 1870
rect 2584 1851 2586 1871
rect 1327 1849 1331 1850
rect 1367 1850 1371 1851
rect 112 1837 114 1849
rect 144 1838 146 1849
rect 200 1838 202 1849
rect 256 1838 258 1849
rect 312 1838 314 1849
rect 376 1838 378 1849
rect 456 1838 458 1849
rect 544 1838 546 1849
rect 632 1838 634 1849
rect 720 1838 722 1849
rect 800 1838 802 1849
rect 888 1838 890 1849
rect 976 1838 978 1849
rect 1064 1838 1066 1849
rect 142 1837 148 1838
rect 110 1836 116 1837
rect 110 1832 111 1836
rect 115 1832 116 1836
rect 142 1833 143 1837
rect 147 1833 148 1837
rect 142 1832 148 1833
rect 198 1837 204 1838
rect 198 1833 199 1837
rect 203 1833 204 1837
rect 198 1832 204 1833
rect 254 1837 260 1838
rect 254 1833 255 1837
rect 259 1833 260 1837
rect 254 1832 260 1833
rect 310 1837 316 1838
rect 310 1833 311 1837
rect 315 1833 316 1837
rect 310 1832 316 1833
rect 374 1837 380 1838
rect 374 1833 375 1837
rect 379 1833 380 1837
rect 374 1832 380 1833
rect 454 1837 460 1838
rect 454 1833 455 1837
rect 459 1833 460 1837
rect 454 1832 460 1833
rect 542 1837 548 1838
rect 542 1833 543 1837
rect 547 1833 548 1837
rect 542 1832 548 1833
rect 630 1837 636 1838
rect 630 1833 631 1837
rect 635 1833 636 1837
rect 630 1832 636 1833
rect 718 1837 724 1838
rect 718 1833 719 1837
rect 723 1833 724 1837
rect 718 1832 724 1833
rect 798 1837 804 1838
rect 798 1833 799 1837
rect 803 1833 804 1837
rect 798 1832 804 1833
rect 886 1837 892 1838
rect 886 1833 887 1837
rect 891 1833 892 1837
rect 886 1832 892 1833
rect 974 1837 980 1838
rect 974 1833 975 1837
rect 979 1833 980 1837
rect 974 1832 980 1833
rect 1062 1837 1068 1838
rect 1328 1837 1330 1849
rect 1367 1845 1371 1846
rect 1559 1850 1563 1851
rect 1559 1845 1563 1846
rect 1615 1850 1619 1851
rect 1615 1845 1619 1846
rect 1623 1850 1627 1851
rect 1623 1845 1627 1846
rect 1671 1850 1675 1851
rect 1671 1845 1675 1846
rect 1679 1850 1683 1851
rect 1679 1845 1683 1846
rect 1727 1850 1731 1851
rect 1727 1845 1731 1846
rect 1735 1850 1739 1851
rect 1735 1845 1739 1846
rect 1783 1850 1787 1851
rect 1783 1845 1787 1846
rect 1791 1850 1795 1851
rect 1791 1845 1795 1846
rect 1839 1850 1843 1851
rect 1839 1845 1843 1846
rect 1847 1850 1851 1851
rect 1847 1845 1851 1846
rect 1903 1850 1907 1851
rect 1903 1845 1907 1846
rect 1911 1850 1915 1851
rect 1911 1845 1915 1846
rect 1967 1850 1971 1851
rect 1967 1845 1971 1846
rect 1999 1850 2003 1851
rect 1999 1845 2003 1846
rect 2039 1850 2043 1851
rect 2039 1845 2043 1846
rect 2111 1850 2115 1851
rect 2111 1845 2115 1846
rect 2127 1850 2131 1851
rect 2127 1845 2131 1846
rect 2223 1850 2227 1851
rect 2223 1845 2227 1846
rect 2231 1850 2235 1851
rect 2231 1845 2235 1846
rect 2327 1850 2331 1851
rect 2327 1845 2331 1846
rect 2367 1850 2371 1851
rect 2367 1845 2371 1846
rect 2439 1850 2443 1851
rect 2439 1845 2443 1846
rect 2503 1850 2507 1851
rect 2503 1845 2507 1846
rect 2527 1850 2531 1851
rect 2527 1845 2531 1846
rect 2583 1850 2587 1851
rect 2583 1845 2587 1846
rect 1062 1833 1063 1837
rect 1067 1833 1068 1837
rect 1062 1832 1068 1833
rect 1326 1836 1332 1837
rect 1326 1832 1327 1836
rect 1331 1832 1332 1836
rect 1368 1833 1370 1845
rect 1624 1834 1626 1845
rect 1680 1834 1682 1845
rect 1736 1834 1738 1845
rect 1792 1834 1794 1845
rect 1848 1834 1850 1845
rect 1904 1834 1906 1845
rect 1968 1834 1970 1845
rect 2040 1834 2042 1845
rect 2128 1834 2130 1845
rect 2224 1834 2226 1845
rect 2328 1834 2330 1845
rect 2440 1834 2442 1845
rect 2528 1834 2530 1845
rect 1622 1833 1628 1834
rect 110 1831 116 1832
rect 1326 1831 1332 1832
rect 1366 1832 1372 1833
rect 1366 1828 1367 1832
rect 1371 1828 1372 1832
rect 1622 1829 1623 1833
rect 1627 1829 1628 1833
rect 1622 1828 1628 1829
rect 1678 1833 1684 1834
rect 1678 1829 1679 1833
rect 1683 1829 1684 1833
rect 1678 1828 1684 1829
rect 1734 1833 1740 1834
rect 1734 1829 1735 1833
rect 1739 1829 1740 1833
rect 1734 1828 1740 1829
rect 1790 1833 1796 1834
rect 1790 1829 1791 1833
rect 1795 1829 1796 1833
rect 1790 1828 1796 1829
rect 1846 1833 1852 1834
rect 1846 1829 1847 1833
rect 1851 1829 1852 1833
rect 1846 1828 1852 1829
rect 1902 1833 1908 1834
rect 1902 1829 1903 1833
rect 1907 1829 1908 1833
rect 1902 1828 1908 1829
rect 1966 1833 1972 1834
rect 1966 1829 1967 1833
rect 1971 1829 1972 1833
rect 1966 1828 1972 1829
rect 2038 1833 2044 1834
rect 2038 1829 2039 1833
rect 2043 1829 2044 1833
rect 2038 1828 2044 1829
rect 2126 1833 2132 1834
rect 2126 1829 2127 1833
rect 2131 1829 2132 1833
rect 2126 1828 2132 1829
rect 2222 1833 2228 1834
rect 2222 1829 2223 1833
rect 2227 1829 2228 1833
rect 2222 1828 2228 1829
rect 2326 1833 2332 1834
rect 2326 1829 2327 1833
rect 2331 1829 2332 1833
rect 2326 1828 2332 1829
rect 2438 1833 2444 1834
rect 2438 1829 2439 1833
rect 2443 1829 2444 1833
rect 2438 1828 2444 1829
rect 2526 1833 2532 1834
rect 2584 1833 2586 1845
rect 2526 1829 2527 1833
rect 2531 1829 2532 1833
rect 2526 1828 2532 1829
rect 2582 1832 2588 1833
rect 2582 1828 2583 1832
rect 2587 1828 2588 1832
rect 1366 1827 1372 1828
rect 2582 1827 2588 1828
rect 110 1819 116 1820
rect 110 1815 111 1819
rect 115 1815 116 1819
rect 110 1814 116 1815
rect 1326 1819 1332 1820
rect 1326 1815 1327 1819
rect 1331 1815 1332 1819
rect 1326 1814 1332 1815
rect 1366 1815 1372 1816
rect 112 1791 114 1814
rect 158 1810 164 1811
rect 158 1806 159 1810
rect 163 1806 164 1810
rect 158 1805 164 1806
rect 214 1810 220 1811
rect 214 1806 215 1810
rect 219 1806 220 1810
rect 214 1805 220 1806
rect 270 1810 276 1811
rect 270 1806 271 1810
rect 275 1806 276 1810
rect 270 1805 276 1806
rect 326 1810 332 1811
rect 326 1806 327 1810
rect 331 1806 332 1810
rect 326 1805 332 1806
rect 390 1810 396 1811
rect 390 1806 391 1810
rect 395 1806 396 1810
rect 390 1805 396 1806
rect 470 1810 476 1811
rect 470 1806 471 1810
rect 475 1806 476 1810
rect 470 1805 476 1806
rect 558 1810 564 1811
rect 558 1806 559 1810
rect 563 1806 564 1810
rect 558 1805 564 1806
rect 646 1810 652 1811
rect 646 1806 647 1810
rect 651 1806 652 1810
rect 646 1805 652 1806
rect 734 1810 740 1811
rect 734 1806 735 1810
rect 739 1806 740 1810
rect 734 1805 740 1806
rect 814 1810 820 1811
rect 814 1806 815 1810
rect 819 1806 820 1810
rect 814 1805 820 1806
rect 902 1810 908 1811
rect 902 1806 903 1810
rect 907 1806 908 1810
rect 902 1805 908 1806
rect 990 1810 996 1811
rect 990 1806 991 1810
rect 995 1806 996 1810
rect 990 1805 996 1806
rect 1078 1810 1084 1811
rect 1078 1806 1079 1810
rect 1083 1806 1084 1810
rect 1078 1805 1084 1806
rect 160 1791 162 1805
rect 216 1791 218 1805
rect 272 1791 274 1805
rect 328 1791 330 1805
rect 392 1791 394 1805
rect 472 1791 474 1805
rect 560 1791 562 1805
rect 648 1791 650 1805
rect 736 1791 738 1805
rect 816 1791 818 1805
rect 904 1791 906 1805
rect 992 1791 994 1805
rect 1080 1791 1082 1805
rect 1328 1791 1330 1814
rect 1366 1811 1367 1815
rect 1371 1811 1372 1815
rect 1366 1810 1372 1811
rect 2582 1815 2588 1816
rect 2582 1811 2583 1815
rect 2587 1811 2588 1815
rect 2582 1810 2588 1811
rect 111 1790 115 1791
rect 111 1785 115 1786
rect 159 1790 163 1791
rect 159 1785 163 1786
rect 215 1790 219 1791
rect 215 1785 219 1786
rect 255 1790 259 1791
rect 255 1785 259 1786
rect 271 1790 275 1791
rect 271 1785 275 1786
rect 327 1790 331 1791
rect 327 1785 331 1786
rect 375 1790 379 1791
rect 375 1785 379 1786
rect 391 1790 395 1791
rect 391 1785 395 1786
rect 471 1790 475 1791
rect 471 1785 475 1786
rect 503 1790 507 1791
rect 503 1785 507 1786
rect 559 1790 563 1791
rect 559 1785 563 1786
rect 623 1790 627 1791
rect 623 1785 627 1786
rect 647 1790 651 1791
rect 647 1785 651 1786
rect 735 1790 739 1791
rect 735 1785 739 1786
rect 743 1790 747 1791
rect 743 1785 747 1786
rect 815 1790 819 1791
rect 815 1785 819 1786
rect 855 1790 859 1791
rect 855 1785 859 1786
rect 903 1790 907 1791
rect 903 1785 907 1786
rect 959 1790 963 1791
rect 959 1785 963 1786
rect 991 1790 995 1791
rect 991 1785 995 1786
rect 1055 1790 1059 1791
rect 1055 1785 1059 1786
rect 1079 1790 1083 1791
rect 1079 1785 1083 1786
rect 1151 1790 1155 1791
rect 1151 1785 1155 1786
rect 1247 1790 1251 1791
rect 1247 1785 1251 1786
rect 1327 1790 1331 1791
rect 1368 1787 1370 1810
rect 1638 1806 1644 1807
rect 1638 1802 1639 1806
rect 1643 1802 1644 1806
rect 1638 1801 1644 1802
rect 1694 1806 1700 1807
rect 1694 1802 1695 1806
rect 1699 1802 1700 1806
rect 1694 1801 1700 1802
rect 1750 1806 1756 1807
rect 1750 1802 1751 1806
rect 1755 1802 1756 1806
rect 1750 1801 1756 1802
rect 1806 1806 1812 1807
rect 1806 1802 1807 1806
rect 1811 1802 1812 1806
rect 1806 1801 1812 1802
rect 1862 1806 1868 1807
rect 1862 1802 1863 1806
rect 1867 1802 1868 1806
rect 1862 1801 1868 1802
rect 1918 1806 1924 1807
rect 1918 1802 1919 1806
rect 1923 1802 1924 1806
rect 1918 1801 1924 1802
rect 1982 1806 1988 1807
rect 1982 1802 1983 1806
rect 1987 1802 1988 1806
rect 1982 1801 1988 1802
rect 2054 1806 2060 1807
rect 2054 1802 2055 1806
rect 2059 1802 2060 1806
rect 2054 1801 2060 1802
rect 2142 1806 2148 1807
rect 2142 1802 2143 1806
rect 2147 1802 2148 1806
rect 2142 1801 2148 1802
rect 2238 1806 2244 1807
rect 2238 1802 2239 1806
rect 2243 1802 2244 1806
rect 2238 1801 2244 1802
rect 2342 1806 2348 1807
rect 2342 1802 2343 1806
rect 2347 1802 2348 1806
rect 2342 1801 2348 1802
rect 2454 1806 2460 1807
rect 2454 1802 2455 1806
rect 2459 1802 2460 1806
rect 2454 1801 2460 1802
rect 2542 1806 2548 1807
rect 2542 1802 2543 1806
rect 2547 1802 2548 1806
rect 2542 1801 2548 1802
rect 1640 1787 1642 1801
rect 1696 1787 1698 1801
rect 1752 1787 1754 1801
rect 1808 1787 1810 1801
rect 1864 1787 1866 1801
rect 1920 1787 1922 1801
rect 1984 1787 1986 1801
rect 2056 1787 2058 1801
rect 2144 1787 2146 1801
rect 2240 1787 2242 1801
rect 2344 1787 2346 1801
rect 2456 1787 2458 1801
rect 2544 1787 2546 1801
rect 2584 1787 2586 1810
rect 1327 1785 1331 1786
rect 1367 1786 1371 1787
rect 112 1770 114 1785
rect 160 1779 162 1785
rect 256 1779 258 1785
rect 376 1779 378 1785
rect 504 1779 506 1785
rect 624 1779 626 1785
rect 744 1779 746 1785
rect 856 1779 858 1785
rect 960 1779 962 1785
rect 1056 1779 1058 1785
rect 1152 1779 1154 1785
rect 1248 1779 1250 1785
rect 158 1778 164 1779
rect 158 1774 159 1778
rect 163 1774 164 1778
rect 158 1773 164 1774
rect 254 1778 260 1779
rect 254 1774 255 1778
rect 259 1774 260 1778
rect 254 1773 260 1774
rect 374 1778 380 1779
rect 374 1774 375 1778
rect 379 1774 380 1778
rect 374 1773 380 1774
rect 502 1778 508 1779
rect 502 1774 503 1778
rect 507 1774 508 1778
rect 502 1773 508 1774
rect 622 1778 628 1779
rect 622 1774 623 1778
rect 627 1774 628 1778
rect 622 1773 628 1774
rect 742 1778 748 1779
rect 742 1774 743 1778
rect 747 1774 748 1778
rect 742 1773 748 1774
rect 854 1778 860 1779
rect 854 1774 855 1778
rect 859 1774 860 1778
rect 854 1773 860 1774
rect 958 1778 964 1779
rect 958 1774 959 1778
rect 963 1774 964 1778
rect 958 1773 964 1774
rect 1054 1778 1060 1779
rect 1054 1774 1055 1778
rect 1059 1774 1060 1778
rect 1054 1773 1060 1774
rect 1150 1778 1156 1779
rect 1150 1774 1151 1778
rect 1155 1774 1156 1778
rect 1150 1773 1156 1774
rect 1246 1778 1252 1779
rect 1246 1774 1247 1778
rect 1251 1774 1252 1778
rect 1246 1773 1252 1774
rect 1328 1770 1330 1785
rect 1367 1781 1371 1782
rect 1471 1786 1475 1787
rect 1471 1781 1475 1782
rect 1535 1786 1539 1787
rect 1535 1781 1539 1782
rect 1615 1786 1619 1787
rect 1615 1781 1619 1782
rect 1639 1786 1643 1787
rect 1639 1781 1643 1782
rect 1695 1786 1699 1787
rect 1695 1781 1699 1782
rect 1751 1786 1755 1787
rect 1751 1781 1755 1782
rect 1783 1786 1787 1787
rect 1783 1781 1787 1782
rect 1807 1786 1811 1787
rect 1807 1781 1811 1782
rect 1863 1786 1867 1787
rect 1863 1781 1867 1782
rect 1879 1786 1883 1787
rect 1879 1781 1883 1782
rect 1919 1786 1923 1787
rect 1919 1781 1923 1782
rect 1975 1786 1979 1787
rect 1975 1781 1979 1782
rect 1983 1786 1987 1787
rect 1983 1781 1987 1782
rect 2055 1786 2059 1787
rect 2055 1781 2059 1782
rect 2071 1786 2075 1787
rect 2071 1781 2075 1782
rect 2143 1786 2147 1787
rect 2143 1781 2147 1782
rect 2167 1786 2171 1787
rect 2167 1781 2171 1782
rect 2239 1786 2243 1787
rect 2239 1781 2243 1782
rect 2263 1786 2267 1787
rect 2263 1781 2267 1782
rect 2343 1786 2347 1787
rect 2343 1781 2347 1782
rect 2359 1786 2363 1787
rect 2359 1781 2363 1782
rect 2455 1786 2459 1787
rect 2455 1781 2459 1782
rect 2463 1786 2467 1787
rect 2463 1781 2467 1782
rect 2543 1786 2547 1787
rect 2543 1781 2547 1782
rect 2583 1786 2587 1787
rect 2583 1781 2587 1782
rect 110 1769 116 1770
rect 110 1765 111 1769
rect 115 1765 116 1769
rect 110 1764 116 1765
rect 1326 1769 1332 1770
rect 1326 1765 1327 1769
rect 1331 1765 1332 1769
rect 1368 1766 1370 1781
rect 1472 1775 1474 1781
rect 1536 1775 1538 1781
rect 1616 1775 1618 1781
rect 1696 1775 1698 1781
rect 1784 1775 1786 1781
rect 1880 1775 1882 1781
rect 1976 1775 1978 1781
rect 2072 1775 2074 1781
rect 2168 1775 2170 1781
rect 2264 1775 2266 1781
rect 2360 1775 2362 1781
rect 2464 1775 2466 1781
rect 2544 1775 2546 1781
rect 1470 1774 1476 1775
rect 1470 1770 1471 1774
rect 1475 1770 1476 1774
rect 1470 1769 1476 1770
rect 1534 1774 1540 1775
rect 1534 1770 1535 1774
rect 1539 1770 1540 1774
rect 1534 1769 1540 1770
rect 1614 1774 1620 1775
rect 1614 1770 1615 1774
rect 1619 1770 1620 1774
rect 1614 1769 1620 1770
rect 1694 1774 1700 1775
rect 1694 1770 1695 1774
rect 1699 1770 1700 1774
rect 1694 1769 1700 1770
rect 1782 1774 1788 1775
rect 1782 1770 1783 1774
rect 1787 1770 1788 1774
rect 1782 1769 1788 1770
rect 1878 1774 1884 1775
rect 1878 1770 1879 1774
rect 1883 1770 1884 1774
rect 1878 1769 1884 1770
rect 1974 1774 1980 1775
rect 1974 1770 1975 1774
rect 1979 1770 1980 1774
rect 1974 1769 1980 1770
rect 2070 1774 2076 1775
rect 2070 1770 2071 1774
rect 2075 1770 2076 1774
rect 2070 1769 2076 1770
rect 2166 1774 2172 1775
rect 2166 1770 2167 1774
rect 2171 1770 2172 1774
rect 2166 1769 2172 1770
rect 2262 1774 2268 1775
rect 2262 1770 2263 1774
rect 2267 1770 2268 1774
rect 2262 1769 2268 1770
rect 2358 1774 2364 1775
rect 2358 1770 2359 1774
rect 2363 1770 2364 1774
rect 2358 1769 2364 1770
rect 2462 1774 2468 1775
rect 2462 1770 2463 1774
rect 2467 1770 2468 1774
rect 2462 1769 2468 1770
rect 2542 1774 2548 1775
rect 2542 1770 2543 1774
rect 2547 1770 2548 1774
rect 2542 1769 2548 1770
rect 2584 1766 2586 1781
rect 1326 1764 1332 1765
rect 1366 1765 1372 1766
rect 1366 1761 1367 1765
rect 1371 1761 1372 1765
rect 1366 1760 1372 1761
rect 2582 1765 2588 1766
rect 2582 1761 2583 1765
rect 2587 1761 2588 1765
rect 2582 1760 2588 1761
rect 110 1752 116 1753
rect 1326 1752 1332 1753
rect 110 1748 111 1752
rect 115 1748 116 1752
rect 110 1747 116 1748
rect 142 1751 148 1752
rect 142 1747 143 1751
rect 147 1747 148 1751
rect 112 1735 114 1747
rect 142 1746 148 1747
rect 238 1751 244 1752
rect 238 1747 239 1751
rect 243 1747 244 1751
rect 238 1746 244 1747
rect 358 1751 364 1752
rect 358 1747 359 1751
rect 363 1747 364 1751
rect 358 1746 364 1747
rect 486 1751 492 1752
rect 486 1747 487 1751
rect 491 1747 492 1751
rect 486 1746 492 1747
rect 606 1751 612 1752
rect 606 1747 607 1751
rect 611 1747 612 1751
rect 606 1746 612 1747
rect 726 1751 732 1752
rect 726 1747 727 1751
rect 731 1747 732 1751
rect 726 1746 732 1747
rect 838 1751 844 1752
rect 838 1747 839 1751
rect 843 1747 844 1751
rect 838 1746 844 1747
rect 942 1751 948 1752
rect 942 1747 943 1751
rect 947 1747 948 1751
rect 942 1746 948 1747
rect 1038 1751 1044 1752
rect 1038 1747 1039 1751
rect 1043 1747 1044 1751
rect 1038 1746 1044 1747
rect 1134 1751 1140 1752
rect 1134 1747 1135 1751
rect 1139 1747 1140 1751
rect 1134 1746 1140 1747
rect 1230 1751 1236 1752
rect 1230 1747 1231 1751
rect 1235 1747 1236 1751
rect 1326 1748 1327 1752
rect 1331 1748 1332 1752
rect 1326 1747 1332 1748
rect 1366 1748 1372 1749
rect 2582 1748 2588 1749
rect 1230 1746 1236 1747
rect 144 1735 146 1746
rect 240 1735 242 1746
rect 360 1735 362 1746
rect 488 1735 490 1746
rect 608 1735 610 1746
rect 728 1735 730 1746
rect 840 1735 842 1746
rect 944 1735 946 1746
rect 1040 1735 1042 1746
rect 1136 1735 1138 1746
rect 1232 1735 1234 1746
rect 1328 1735 1330 1747
rect 1366 1744 1367 1748
rect 1371 1744 1372 1748
rect 1366 1743 1372 1744
rect 1454 1747 1460 1748
rect 1454 1743 1455 1747
rect 1459 1743 1460 1747
rect 111 1734 115 1735
rect 111 1729 115 1730
rect 143 1734 147 1735
rect 143 1729 147 1730
rect 239 1734 243 1735
rect 239 1729 243 1730
rect 263 1734 267 1735
rect 263 1729 267 1730
rect 359 1734 363 1735
rect 359 1729 363 1730
rect 415 1734 419 1735
rect 415 1729 419 1730
rect 487 1734 491 1735
rect 487 1729 491 1730
rect 567 1734 571 1735
rect 567 1729 571 1730
rect 607 1734 611 1735
rect 607 1729 611 1730
rect 711 1734 715 1735
rect 711 1729 715 1730
rect 727 1734 731 1735
rect 727 1729 731 1730
rect 839 1734 843 1735
rect 839 1729 843 1730
rect 855 1734 859 1735
rect 855 1729 859 1730
rect 943 1734 947 1735
rect 943 1729 947 1730
rect 999 1734 1003 1735
rect 999 1729 1003 1730
rect 1039 1734 1043 1735
rect 1039 1729 1043 1730
rect 1135 1734 1139 1735
rect 1135 1729 1139 1730
rect 1143 1734 1147 1735
rect 1143 1729 1147 1730
rect 1231 1734 1235 1735
rect 1231 1729 1235 1730
rect 1271 1734 1275 1735
rect 1271 1729 1275 1730
rect 1327 1734 1331 1735
rect 1327 1729 1331 1730
rect 112 1717 114 1729
rect 144 1718 146 1729
rect 264 1718 266 1729
rect 416 1718 418 1729
rect 568 1718 570 1729
rect 712 1718 714 1729
rect 856 1718 858 1729
rect 1000 1718 1002 1729
rect 1144 1718 1146 1729
rect 1272 1718 1274 1729
rect 142 1717 148 1718
rect 110 1716 116 1717
rect 110 1712 111 1716
rect 115 1712 116 1716
rect 142 1713 143 1717
rect 147 1713 148 1717
rect 142 1712 148 1713
rect 262 1717 268 1718
rect 262 1713 263 1717
rect 267 1713 268 1717
rect 262 1712 268 1713
rect 414 1717 420 1718
rect 414 1713 415 1717
rect 419 1713 420 1717
rect 414 1712 420 1713
rect 566 1717 572 1718
rect 566 1713 567 1717
rect 571 1713 572 1717
rect 566 1712 572 1713
rect 710 1717 716 1718
rect 710 1713 711 1717
rect 715 1713 716 1717
rect 710 1712 716 1713
rect 854 1717 860 1718
rect 854 1713 855 1717
rect 859 1713 860 1717
rect 854 1712 860 1713
rect 998 1717 1004 1718
rect 998 1713 999 1717
rect 1003 1713 1004 1717
rect 998 1712 1004 1713
rect 1142 1717 1148 1718
rect 1142 1713 1143 1717
rect 1147 1713 1148 1717
rect 1142 1712 1148 1713
rect 1270 1717 1276 1718
rect 1328 1717 1330 1729
rect 1368 1727 1370 1743
rect 1454 1742 1460 1743
rect 1518 1747 1524 1748
rect 1518 1743 1519 1747
rect 1523 1743 1524 1747
rect 1518 1742 1524 1743
rect 1598 1747 1604 1748
rect 1598 1743 1599 1747
rect 1603 1743 1604 1747
rect 1598 1742 1604 1743
rect 1678 1747 1684 1748
rect 1678 1743 1679 1747
rect 1683 1743 1684 1747
rect 1678 1742 1684 1743
rect 1766 1747 1772 1748
rect 1766 1743 1767 1747
rect 1771 1743 1772 1747
rect 1766 1742 1772 1743
rect 1862 1747 1868 1748
rect 1862 1743 1863 1747
rect 1867 1743 1868 1747
rect 1862 1742 1868 1743
rect 1958 1747 1964 1748
rect 1958 1743 1959 1747
rect 1963 1743 1964 1747
rect 1958 1742 1964 1743
rect 2054 1747 2060 1748
rect 2054 1743 2055 1747
rect 2059 1743 2060 1747
rect 2054 1742 2060 1743
rect 2150 1747 2156 1748
rect 2150 1743 2151 1747
rect 2155 1743 2156 1747
rect 2150 1742 2156 1743
rect 2246 1747 2252 1748
rect 2246 1743 2247 1747
rect 2251 1743 2252 1747
rect 2246 1742 2252 1743
rect 2342 1747 2348 1748
rect 2342 1743 2343 1747
rect 2347 1743 2348 1747
rect 2342 1742 2348 1743
rect 2446 1747 2452 1748
rect 2446 1743 2447 1747
rect 2451 1743 2452 1747
rect 2446 1742 2452 1743
rect 2526 1747 2532 1748
rect 2526 1743 2527 1747
rect 2531 1743 2532 1747
rect 2582 1744 2583 1748
rect 2587 1744 2588 1748
rect 2582 1743 2588 1744
rect 2526 1742 2532 1743
rect 1456 1727 1458 1742
rect 1520 1727 1522 1742
rect 1600 1727 1602 1742
rect 1680 1727 1682 1742
rect 1768 1727 1770 1742
rect 1864 1727 1866 1742
rect 1960 1727 1962 1742
rect 2056 1727 2058 1742
rect 2152 1727 2154 1742
rect 2248 1727 2250 1742
rect 2344 1727 2346 1742
rect 2448 1727 2450 1742
rect 2528 1727 2530 1742
rect 2584 1727 2586 1743
rect 1367 1726 1371 1727
rect 1367 1721 1371 1722
rect 1399 1726 1403 1727
rect 1399 1721 1403 1722
rect 1455 1726 1459 1727
rect 1455 1721 1459 1722
rect 1479 1726 1483 1727
rect 1479 1721 1483 1722
rect 1519 1726 1523 1727
rect 1519 1721 1523 1722
rect 1599 1726 1603 1727
rect 1599 1721 1603 1722
rect 1679 1726 1683 1727
rect 1679 1721 1683 1722
rect 1719 1726 1723 1727
rect 1719 1721 1723 1722
rect 1767 1726 1771 1727
rect 1767 1721 1771 1722
rect 1839 1726 1843 1727
rect 1839 1721 1843 1722
rect 1863 1726 1867 1727
rect 1863 1721 1867 1722
rect 1951 1726 1955 1727
rect 1951 1721 1955 1722
rect 1959 1726 1963 1727
rect 1959 1721 1963 1722
rect 2055 1726 2059 1727
rect 2055 1721 2059 1722
rect 2151 1726 2155 1727
rect 2151 1721 2155 1722
rect 2159 1726 2163 1727
rect 2159 1721 2163 1722
rect 2247 1726 2251 1727
rect 2247 1721 2251 1722
rect 2255 1726 2259 1727
rect 2255 1721 2259 1722
rect 2343 1726 2347 1727
rect 2343 1721 2347 1722
rect 2351 1726 2355 1727
rect 2351 1721 2355 1722
rect 2447 1726 2451 1727
rect 2447 1721 2451 1722
rect 2527 1726 2531 1727
rect 2527 1721 2531 1722
rect 2583 1726 2587 1727
rect 2583 1721 2587 1722
rect 1270 1713 1271 1717
rect 1275 1713 1276 1717
rect 1270 1712 1276 1713
rect 1326 1716 1332 1717
rect 1326 1712 1327 1716
rect 1331 1712 1332 1716
rect 110 1711 116 1712
rect 1326 1711 1332 1712
rect 1368 1709 1370 1721
rect 1400 1710 1402 1721
rect 1480 1710 1482 1721
rect 1600 1710 1602 1721
rect 1720 1710 1722 1721
rect 1840 1710 1842 1721
rect 1952 1710 1954 1721
rect 2056 1710 2058 1721
rect 2160 1710 2162 1721
rect 2256 1710 2258 1721
rect 2352 1710 2354 1721
rect 2448 1710 2450 1721
rect 2528 1710 2530 1721
rect 1398 1709 1404 1710
rect 1366 1708 1372 1709
rect 1366 1704 1367 1708
rect 1371 1704 1372 1708
rect 1398 1705 1399 1709
rect 1403 1705 1404 1709
rect 1398 1704 1404 1705
rect 1478 1709 1484 1710
rect 1478 1705 1479 1709
rect 1483 1705 1484 1709
rect 1478 1704 1484 1705
rect 1598 1709 1604 1710
rect 1598 1705 1599 1709
rect 1603 1705 1604 1709
rect 1598 1704 1604 1705
rect 1718 1709 1724 1710
rect 1718 1705 1719 1709
rect 1723 1705 1724 1709
rect 1718 1704 1724 1705
rect 1838 1709 1844 1710
rect 1838 1705 1839 1709
rect 1843 1705 1844 1709
rect 1838 1704 1844 1705
rect 1950 1709 1956 1710
rect 1950 1705 1951 1709
rect 1955 1705 1956 1709
rect 1950 1704 1956 1705
rect 2054 1709 2060 1710
rect 2054 1705 2055 1709
rect 2059 1705 2060 1709
rect 2054 1704 2060 1705
rect 2158 1709 2164 1710
rect 2158 1705 2159 1709
rect 2163 1705 2164 1709
rect 2158 1704 2164 1705
rect 2254 1709 2260 1710
rect 2254 1705 2255 1709
rect 2259 1705 2260 1709
rect 2254 1704 2260 1705
rect 2350 1709 2356 1710
rect 2350 1705 2351 1709
rect 2355 1705 2356 1709
rect 2350 1704 2356 1705
rect 2446 1709 2452 1710
rect 2446 1705 2447 1709
rect 2451 1705 2452 1709
rect 2446 1704 2452 1705
rect 2526 1709 2532 1710
rect 2584 1709 2586 1721
rect 2526 1705 2527 1709
rect 2531 1705 2532 1709
rect 2526 1704 2532 1705
rect 2582 1708 2588 1709
rect 2582 1704 2583 1708
rect 2587 1704 2588 1708
rect 1366 1703 1372 1704
rect 2582 1703 2588 1704
rect 110 1699 116 1700
rect 110 1695 111 1699
rect 115 1695 116 1699
rect 110 1694 116 1695
rect 1326 1699 1332 1700
rect 1326 1695 1327 1699
rect 1331 1695 1332 1699
rect 1326 1694 1332 1695
rect 112 1675 114 1694
rect 158 1690 164 1691
rect 158 1686 159 1690
rect 163 1686 164 1690
rect 158 1685 164 1686
rect 278 1690 284 1691
rect 278 1686 279 1690
rect 283 1686 284 1690
rect 278 1685 284 1686
rect 430 1690 436 1691
rect 430 1686 431 1690
rect 435 1686 436 1690
rect 430 1685 436 1686
rect 582 1690 588 1691
rect 582 1686 583 1690
rect 587 1686 588 1690
rect 582 1685 588 1686
rect 726 1690 732 1691
rect 726 1686 727 1690
rect 731 1686 732 1690
rect 726 1685 732 1686
rect 870 1690 876 1691
rect 870 1686 871 1690
rect 875 1686 876 1690
rect 870 1685 876 1686
rect 1014 1690 1020 1691
rect 1014 1686 1015 1690
rect 1019 1686 1020 1690
rect 1014 1685 1020 1686
rect 1158 1690 1164 1691
rect 1158 1686 1159 1690
rect 1163 1686 1164 1690
rect 1158 1685 1164 1686
rect 1286 1690 1292 1691
rect 1286 1686 1287 1690
rect 1291 1686 1292 1690
rect 1286 1685 1292 1686
rect 160 1675 162 1685
rect 280 1675 282 1685
rect 432 1675 434 1685
rect 584 1675 586 1685
rect 728 1675 730 1685
rect 872 1675 874 1685
rect 1016 1675 1018 1685
rect 1160 1675 1162 1685
rect 1288 1675 1290 1685
rect 1328 1675 1330 1694
rect 1366 1691 1372 1692
rect 1366 1687 1367 1691
rect 1371 1687 1372 1691
rect 1366 1686 1372 1687
rect 2582 1691 2588 1692
rect 2582 1687 2583 1691
rect 2587 1687 2588 1691
rect 2582 1686 2588 1687
rect 111 1674 115 1675
rect 111 1669 115 1670
rect 159 1674 163 1675
rect 159 1669 163 1670
rect 223 1674 227 1675
rect 223 1669 227 1670
rect 279 1674 283 1675
rect 279 1669 283 1670
rect 303 1674 307 1675
rect 303 1669 307 1670
rect 383 1674 387 1675
rect 383 1669 387 1670
rect 431 1674 435 1675
rect 431 1669 435 1670
rect 463 1674 467 1675
rect 463 1669 467 1670
rect 535 1674 539 1675
rect 535 1669 539 1670
rect 583 1674 587 1675
rect 583 1669 587 1670
rect 607 1674 611 1675
rect 607 1669 611 1670
rect 679 1674 683 1675
rect 679 1669 683 1670
rect 727 1674 731 1675
rect 727 1669 731 1670
rect 767 1674 771 1675
rect 767 1669 771 1670
rect 863 1674 867 1675
rect 863 1669 867 1670
rect 871 1674 875 1675
rect 871 1669 875 1670
rect 967 1674 971 1675
rect 967 1669 971 1670
rect 1015 1674 1019 1675
rect 1015 1669 1019 1670
rect 1079 1674 1083 1675
rect 1079 1669 1083 1670
rect 1159 1674 1163 1675
rect 1159 1669 1163 1670
rect 1191 1674 1195 1675
rect 1191 1669 1195 1670
rect 1287 1674 1291 1675
rect 1287 1669 1291 1670
rect 1327 1674 1331 1675
rect 1368 1671 1370 1686
rect 1414 1682 1420 1683
rect 1414 1678 1415 1682
rect 1419 1678 1420 1682
rect 1414 1677 1420 1678
rect 1494 1682 1500 1683
rect 1494 1678 1495 1682
rect 1499 1678 1500 1682
rect 1494 1677 1500 1678
rect 1614 1682 1620 1683
rect 1614 1678 1615 1682
rect 1619 1678 1620 1682
rect 1614 1677 1620 1678
rect 1734 1682 1740 1683
rect 1734 1678 1735 1682
rect 1739 1678 1740 1682
rect 1734 1677 1740 1678
rect 1854 1682 1860 1683
rect 1854 1678 1855 1682
rect 1859 1678 1860 1682
rect 1854 1677 1860 1678
rect 1966 1682 1972 1683
rect 1966 1678 1967 1682
rect 1971 1678 1972 1682
rect 1966 1677 1972 1678
rect 2070 1682 2076 1683
rect 2070 1678 2071 1682
rect 2075 1678 2076 1682
rect 2070 1677 2076 1678
rect 2174 1682 2180 1683
rect 2174 1678 2175 1682
rect 2179 1678 2180 1682
rect 2174 1677 2180 1678
rect 2270 1682 2276 1683
rect 2270 1678 2271 1682
rect 2275 1678 2276 1682
rect 2270 1677 2276 1678
rect 2366 1682 2372 1683
rect 2366 1678 2367 1682
rect 2371 1678 2372 1682
rect 2366 1677 2372 1678
rect 2462 1682 2468 1683
rect 2462 1678 2463 1682
rect 2467 1678 2468 1682
rect 2462 1677 2468 1678
rect 2542 1682 2548 1683
rect 2542 1678 2543 1682
rect 2547 1678 2548 1682
rect 2542 1677 2548 1678
rect 1416 1671 1418 1677
rect 1496 1671 1498 1677
rect 1616 1671 1618 1677
rect 1736 1671 1738 1677
rect 1856 1671 1858 1677
rect 1968 1671 1970 1677
rect 2072 1671 2074 1677
rect 2176 1671 2178 1677
rect 2272 1671 2274 1677
rect 2368 1671 2370 1677
rect 2464 1671 2466 1677
rect 2544 1671 2546 1677
rect 2584 1671 2586 1686
rect 1327 1669 1331 1670
rect 1367 1670 1371 1671
rect 112 1654 114 1669
rect 160 1663 162 1669
rect 224 1663 226 1669
rect 304 1663 306 1669
rect 384 1663 386 1669
rect 464 1663 466 1669
rect 536 1663 538 1669
rect 608 1663 610 1669
rect 680 1663 682 1669
rect 768 1663 770 1669
rect 864 1663 866 1669
rect 968 1663 970 1669
rect 1080 1663 1082 1669
rect 1192 1663 1194 1669
rect 1288 1663 1290 1669
rect 158 1662 164 1663
rect 158 1658 159 1662
rect 163 1658 164 1662
rect 158 1657 164 1658
rect 222 1662 228 1663
rect 222 1658 223 1662
rect 227 1658 228 1662
rect 222 1657 228 1658
rect 302 1662 308 1663
rect 302 1658 303 1662
rect 307 1658 308 1662
rect 302 1657 308 1658
rect 382 1662 388 1663
rect 382 1658 383 1662
rect 387 1658 388 1662
rect 382 1657 388 1658
rect 462 1662 468 1663
rect 462 1658 463 1662
rect 467 1658 468 1662
rect 462 1657 468 1658
rect 534 1662 540 1663
rect 534 1658 535 1662
rect 539 1658 540 1662
rect 534 1657 540 1658
rect 606 1662 612 1663
rect 606 1658 607 1662
rect 611 1658 612 1662
rect 606 1657 612 1658
rect 678 1662 684 1663
rect 678 1658 679 1662
rect 683 1658 684 1662
rect 678 1657 684 1658
rect 766 1662 772 1663
rect 766 1658 767 1662
rect 771 1658 772 1662
rect 766 1657 772 1658
rect 862 1662 868 1663
rect 862 1658 863 1662
rect 867 1658 868 1662
rect 862 1657 868 1658
rect 966 1662 972 1663
rect 966 1658 967 1662
rect 971 1658 972 1662
rect 966 1657 972 1658
rect 1078 1662 1084 1663
rect 1078 1658 1079 1662
rect 1083 1658 1084 1662
rect 1078 1657 1084 1658
rect 1190 1662 1196 1663
rect 1190 1658 1191 1662
rect 1195 1658 1196 1662
rect 1190 1657 1196 1658
rect 1286 1662 1292 1663
rect 1286 1658 1287 1662
rect 1291 1658 1292 1662
rect 1286 1657 1292 1658
rect 1328 1654 1330 1669
rect 1367 1665 1371 1666
rect 1415 1670 1419 1671
rect 1415 1665 1419 1666
rect 1495 1670 1499 1671
rect 1495 1665 1499 1666
rect 1503 1670 1507 1671
rect 1503 1665 1507 1666
rect 1615 1670 1619 1671
rect 1615 1665 1619 1666
rect 1623 1670 1627 1671
rect 1623 1665 1627 1666
rect 1735 1670 1739 1671
rect 1735 1665 1739 1666
rect 1751 1670 1755 1671
rect 1751 1665 1755 1666
rect 1855 1670 1859 1671
rect 1855 1665 1859 1666
rect 1879 1670 1883 1671
rect 1879 1665 1883 1666
rect 1967 1670 1971 1671
rect 1967 1665 1971 1666
rect 1999 1670 2003 1671
rect 1999 1665 2003 1666
rect 2071 1670 2075 1671
rect 2071 1665 2075 1666
rect 2119 1670 2123 1671
rect 2119 1665 2123 1666
rect 2175 1670 2179 1671
rect 2175 1665 2179 1666
rect 2231 1670 2235 1671
rect 2231 1665 2235 1666
rect 2271 1670 2275 1671
rect 2271 1665 2275 1666
rect 2343 1670 2347 1671
rect 2343 1665 2347 1666
rect 2367 1670 2371 1671
rect 2367 1665 2371 1666
rect 2455 1670 2459 1671
rect 2455 1665 2459 1666
rect 2463 1670 2467 1671
rect 2463 1665 2467 1666
rect 2543 1670 2547 1671
rect 2543 1665 2547 1666
rect 2583 1670 2587 1671
rect 2583 1665 2587 1666
rect 110 1653 116 1654
rect 110 1649 111 1653
rect 115 1649 116 1653
rect 110 1648 116 1649
rect 1326 1653 1332 1654
rect 1326 1649 1327 1653
rect 1331 1649 1332 1653
rect 1368 1650 1370 1665
rect 1416 1659 1418 1665
rect 1504 1659 1506 1665
rect 1624 1659 1626 1665
rect 1752 1659 1754 1665
rect 1880 1659 1882 1665
rect 2000 1659 2002 1665
rect 2120 1659 2122 1665
rect 2232 1659 2234 1665
rect 2344 1659 2346 1665
rect 2456 1659 2458 1665
rect 2544 1659 2546 1665
rect 1414 1658 1420 1659
rect 1414 1654 1415 1658
rect 1419 1654 1420 1658
rect 1414 1653 1420 1654
rect 1502 1658 1508 1659
rect 1502 1654 1503 1658
rect 1507 1654 1508 1658
rect 1502 1653 1508 1654
rect 1622 1658 1628 1659
rect 1622 1654 1623 1658
rect 1627 1654 1628 1658
rect 1622 1653 1628 1654
rect 1750 1658 1756 1659
rect 1750 1654 1751 1658
rect 1755 1654 1756 1658
rect 1750 1653 1756 1654
rect 1878 1658 1884 1659
rect 1878 1654 1879 1658
rect 1883 1654 1884 1658
rect 1878 1653 1884 1654
rect 1998 1658 2004 1659
rect 1998 1654 1999 1658
rect 2003 1654 2004 1658
rect 1998 1653 2004 1654
rect 2118 1658 2124 1659
rect 2118 1654 2119 1658
rect 2123 1654 2124 1658
rect 2118 1653 2124 1654
rect 2230 1658 2236 1659
rect 2230 1654 2231 1658
rect 2235 1654 2236 1658
rect 2230 1653 2236 1654
rect 2342 1658 2348 1659
rect 2342 1654 2343 1658
rect 2347 1654 2348 1658
rect 2342 1653 2348 1654
rect 2454 1658 2460 1659
rect 2454 1654 2455 1658
rect 2459 1654 2460 1658
rect 2454 1653 2460 1654
rect 2542 1658 2548 1659
rect 2542 1654 2543 1658
rect 2547 1654 2548 1658
rect 2542 1653 2548 1654
rect 2584 1650 2586 1665
rect 1326 1648 1332 1649
rect 1366 1649 1372 1650
rect 1366 1645 1367 1649
rect 1371 1645 1372 1649
rect 1366 1644 1372 1645
rect 2582 1649 2588 1650
rect 2582 1645 2583 1649
rect 2587 1645 2588 1649
rect 2582 1644 2588 1645
rect 110 1636 116 1637
rect 1326 1636 1332 1637
rect 110 1632 111 1636
rect 115 1632 116 1636
rect 110 1631 116 1632
rect 142 1635 148 1636
rect 142 1631 143 1635
rect 147 1631 148 1635
rect 112 1619 114 1631
rect 142 1630 148 1631
rect 206 1635 212 1636
rect 206 1631 207 1635
rect 211 1631 212 1635
rect 206 1630 212 1631
rect 286 1635 292 1636
rect 286 1631 287 1635
rect 291 1631 292 1635
rect 286 1630 292 1631
rect 366 1635 372 1636
rect 366 1631 367 1635
rect 371 1631 372 1635
rect 366 1630 372 1631
rect 446 1635 452 1636
rect 446 1631 447 1635
rect 451 1631 452 1635
rect 446 1630 452 1631
rect 518 1635 524 1636
rect 518 1631 519 1635
rect 523 1631 524 1635
rect 518 1630 524 1631
rect 590 1635 596 1636
rect 590 1631 591 1635
rect 595 1631 596 1635
rect 590 1630 596 1631
rect 662 1635 668 1636
rect 662 1631 663 1635
rect 667 1631 668 1635
rect 662 1630 668 1631
rect 750 1635 756 1636
rect 750 1631 751 1635
rect 755 1631 756 1635
rect 750 1630 756 1631
rect 846 1635 852 1636
rect 846 1631 847 1635
rect 851 1631 852 1635
rect 846 1630 852 1631
rect 950 1635 956 1636
rect 950 1631 951 1635
rect 955 1631 956 1635
rect 950 1630 956 1631
rect 1062 1635 1068 1636
rect 1062 1631 1063 1635
rect 1067 1631 1068 1635
rect 1062 1630 1068 1631
rect 1174 1635 1180 1636
rect 1174 1631 1175 1635
rect 1179 1631 1180 1635
rect 1174 1630 1180 1631
rect 1270 1635 1276 1636
rect 1270 1631 1271 1635
rect 1275 1631 1276 1635
rect 1326 1632 1327 1636
rect 1331 1632 1332 1636
rect 1326 1631 1332 1632
rect 1366 1632 1372 1633
rect 2582 1632 2588 1633
rect 1270 1630 1276 1631
rect 144 1619 146 1630
rect 208 1619 210 1630
rect 288 1619 290 1630
rect 368 1619 370 1630
rect 448 1619 450 1630
rect 520 1619 522 1630
rect 592 1619 594 1630
rect 664 1619 666 1630
rect 752 1619 754 1630
rect 848 1619 850 1630
rect 952 1619 954 1630
rect 1064 1619 1066 1630
rect 1176 1619 1178 1630
rect 1272 1619 1274 1630
rect 1328 1619 1330 1631
rect 1366 1628 1367 1632
rect 1371 1628 1372 1632
rect 1366 1627 1372 1628
rect 1398 1631 1404 1632
rect 1398 1627 1399 1631
rect 1403 1627 1404 1631
rect 111 1618 115 1619
rect 111 1613 115 1614
rect 143 1618 147 1619
rect 143 1613 147 1614
rect 207 1618 211 1619
rect 207 1613 211 1614
rect 247 1618 251 1619
rect 247 1613 251 1614
rect 287 1618 291 1619
rect 287 1613 291 1614
rect 367 1618 371 1619
rect 367 1613 371 1614
rect 447 1618 451 1619
rect 447 1613 451 1614
rect 479 1618 483 1619
rect 479 1613 483 1614
rect 519 1618 523 1619
rect 519 1613 523 1614
rect 575 1618 579 1619
rect 575 1613 579 1614
rect 591 1618 595 1619
rect 591 1613 595 1614
rect 663 1618 667 1619
rect 663 1613 667 1614
rect 671 1618 675 1619
rect 671 1613 675 1614
rect 751 1618 755 1619
rect 751 1613 755 1614
rect 767 1618 771 1619
rect 767 1613 771 1614
rect 847 1618 851 1619
rect 847 1613 851 1614
rect 863 1618 867 1619
rect 863 1613 867 1614
rect 951 1618 955 1619
rect 951 1613 955 1614
rect 959 1618 963 1619
rect 959 1613 963 1614
rect 1063 1618 1067 1619
rect 1063 1613 1067 1614
rect 1175 1618 1179 1619
rect 1175 1613 1179 1614
rect 1271 1618 1275 1619
rect 1271 1613 1275 1614
rect 1327 1618 1331 1619
rect 1327 1613 1331 1614
rect 112 1601 114 1613
rect 144 1602 146 1613
rect 248 1602 250 1613
rect 368 1602 370 1613
rect 480 1602 482 1613
rect 576 1602 578 1613
rect 672 1602 674 1613
rect 768 1602 770 1613
rect 864 1602 866 1613
rect 960 1602 962 1613
rect 1064 1602 1066 1613
rect 1176 1602 1178 1613
rect 1272 1602 1274 1613
rect 142 1601 148 1602
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 142 1597 143 1601
rect 147 1597 148 1601
rect 142 1596 148 1597
rect 246 1601 252 1602
rect 246 1597 247 1601
rect 251 1597 252 1601
rect 246 1596 252 1597
rect 366 1601 372 1602
rect 366 1597 367 1601
rect 371 1597 372 1601
rect 366 1596 372 1597
rect 478 1601 484 1602
rect 478 1597 479 1601
rect 483 1597 484 1601
rect 478 1596 484 1597
rect 574 1601 580 1602
rect 574 1597 575 1601
rect 579 1597 580 1601
rect 574 1596 580 1597
rect 670 1601 676 1602
rect 670 1597 671 1601
rect 675 1597 676 1601
rect 670 1596 676 1597
rect 766 1601 772 1602
rect 766 1597 767 1601
rect 771 1597 772 1601
rect 766 1596 772 1597
rect 862 1601 868 1602
rect 862 1597 863 1601
rect 867 1597 868 1601
rect 862 1596 868 1597
rect 958 1601 964 1602
rect 958 1597 959 1601
rect 963 1597 964 1601
rect 958 1596 964 1597
rect 1062 1601 1068 1602
rect 1062 1597 1063 1601
rect 1067 1597 1068 1601
rect 1062 1596 1068 1597
rect 1174 1601 1180 1602
rect 1174 1597 1175 1601
rect 1179 1597 1180 1601
rect 1174 1596 1180 1597
rect 1270 1601 1276 1602
rect 1328 1601 1330 1613
rect 1368 1603 1370 1627
rect 1398 1626 1404 1627
rect 1486 1631 1492 1632
rect 1486 1627 1487 1631
rect 1491 1627 1492 1631
rect 1486 1626 1492 1627
rect 1606 1631 1612 1632
rect 1606 1627 1607 1631
rect 1611 1627 1612 1631
rect 1606 1626 1612 1627
rect 1734 1631 1740 1632
rect 1734 1627 1735 1631
rect 1739 1627 1740 1631
rect 1734 1626 1740 1627
rect 1862 1631 1868 1632
rect 1862 1627 1863 1631
rect 1867 1627 1868 1631
rect 1862 1626 1868 1627
rect 1982 1631 1988 1632
rect 1982 1627 1983 1631
rect 1987 1627 1988 1631
rect 1982 1626 1988 1627
rect 2102 1631 2108 1632
rect 2102 1627 2103 1631
rect 2107 1627 2108 1631
rect 2102 1626 2108 1627
rect 2214 1631 2220 1632
rect 2214 1627 2215 1631
rect 2219 1627 2220 1631
rect 2214 1626 2220 1627
rect 2326 1631 2332 1632
rect 2326 1627 2327 1631
rect 2331 1627 2332 1631
rect 2326 1626 2332 1627
rect 2438 1631 2444 1632
rect 2438 1627 2439 1631
rect 2443 1627 2444 1631
rect 2438 1626 2444 1627
rect 2526 1631 2532 1632
rect 2526 1627 2527 1631
rect 2531 1627 2532 1631
rect 2582 1628 2583 1632
rect 2587 1628 2588 1632
rect 2582 1627 2588 1628
rect 2526 1626 2532 1627
rect 1400 1603 1402 1626
rect 1488 1603 1490 1626
rect 1608 1603 1610 1626
rect 1736 1603 1738 1626
rect 1864 1603 1866 1626
rect 1984 1603 1986 1626
rect 2104 1603 2106 1626
rect 2216 1603 2218 1626
rect 2328 1603 2330 1626
rect 2440 1603 2442 1626
rect 2528 1603 2530 1626
rect 2584 1603 2586 1627
rect 1367 1602 1371 1603
rect 1270 1597 1271 1601
rect 1275 1597 1276 1601
rect 1270 1596 1276 1597
rect 1326 1600 1332 1601
rect 1326 1596 1327 1600
rect 1331 1596 1332 1600
rect 1367 1597 1371 1598
rect 1399 1602 1403 1603
rect 1399 1597 1403 1598
rect 1487 1602 1491 1603
rect 1487 1597 1491 1598
rect 1495 1602 1499 1603
rect 1495 1597 1499 1598
rect 1607 1602 1611 1603
rect 1607 1597 1611 1598
rect 1615 1602 1619 1603
rect 1615 1597 1619 1598
rect 1735 1602 1739 1603
rect 1735 1597 1739 1598
rect 1743 1602 1747 1603
rect 1743 1597 1747 1598
rect 1863 1602 1867 1603
rect 1863 1597 1867 1598
rect 1983 1602 1987 1603
rect 1983 1597 1987 1598
rect 2095 1602 2099 1603
rect 2095 1597 2099 1598
rect 2103 1602 2107 1603
rect 2103 1597 2107 1598
rect 2199 1602 2203 1603
rect 2199 1597 2203 1598
rect 2215 1602 2219 1603
rect 2215 1597 2219 1598
rect 2295 1602 2299 1603
rect 2295 1597 2299 1598
rect 2327 1602 2331 1603
rect 2327 1597 2331 1598
rect 2391 1602 2395 1603
rect 2391 1597 2395 1598
rect 2439 1602 2443 1603
rect 2439 1597 2443 1598
rect 2495 1602 2499 1603
rect 2495 1597 2499 1598
rect 2527 1602 2531 1603
rect 2527 1597 2531 1598
rect 2583 1602 2587 1603
rect 2583 1597 2587 1598
rect 110 1595 116 1596
rect 1326 1595 1332 1596
rect 1368 1585 1370 1597
rect 1400 1586 1402 1597
rect 1496 1586 1498 1597
rect 1616 1586 1618 1597
rect 1744 1586 1746 1597
rect 1864 1586 1866 1597
rect 1984 1586 1986 1597
rect 2096 1586 2098 1597
rect 2200 1586 2202 1597
rect 2296 1586 2298 1597
rect 2392 1586 2394 1597
rect 2496 1586 2498 1597
rect 1398 1585 1404 1586
rect 1366 1584 1372 1585
rect 110 1583 116 1584
rect 110 1579 111 1583
rect 115 1579 116 1583
rect 110 1578 116 1579
rect 1326 1583 1332 1584
rect 1326 1579 1327 1583
rect 1331 1579 1332 1583
rect 1366 1580 1367 1584
rect 1371 1580 1372 1584
rect 1398 1581 1399 1585
rect 1403 1581 1404 1585
rect 1398 1580 1404 1581
rect 1494 1585 1500 1586
rect 1494 1581 1495 1585
rect 1499 1581 1500 1585
rect 1494 1580 1500 1581
rect 1614 1585 1620 1586
rect 1614 1581 1615 1585
rect 1619 1581 1620 1585
rect 1614 1580 1620 1581
rect 1742 1585 1748 1586
rect 1742 1581 1743 1585
rect 1747 1581 1748 1585
rect 1742 1580 1748 1581
rect 1862 1585 1868 1586
rect 1862 1581 1863 1585
rect 1867 1581 1868 1585
rect 1862 1580 1868 1581
rect 1982 1585 1988 1586
rect 1982 1581 1983 1585
rect 1987 1581 1988 1585
rect 1982 1580 1988 1581
rect 2094 1585 2100 1586
rect 2094 1581 2095 1585
rect 2099 1581 2100 1585
rect 2094 1580 2100 1581
rect 2198 1585 2204 1586
rect 2198 1581 2199 1585
rect 2203 1581 2204 1585
rect 2198 1580 2204 1581
rect 2294 1585 2300 1586
rect 2294 1581 2295 1585
rect 2299 1581 2300 1585
rect 2294 1580 2300 1581
rect 2390 1585 2396 1586
rect 2390 1581 2391 1585
rect 2395 1581 2396 1585
rect 2390 1580 2396 1581
rect 2494 1585 2500 1586
rect 2584 1585 2586 1597
rect 2494 1581 2495 1585
rect 2499 1581 2500 1585
rect 2494 1580 2500 1581
rect 2582 1584 2588 1585
rect 2582 1580 2583 1584
rect 2587 1580 2588 1584
rect 1366 1579 1372 1580
rect 2582 1579 2588 1580
rect 1326 1578 1332 1579
rect 112 1559 114 1578
rect 158 1574 164 1575
rect 158 1570 159 1574
rect 163 1570 164 1574
rect 158 1569 164 1570
rect 262 1574 268 1575
rect 262 1570 263 1574
rect 267 1570 268 1574
rect 262 1569 268 1570
rect 382 1574 388 1575
rect 382 1570 383 1574
rect 387 1570 388 1574
rect 382 1569 388 1570
rect 494 1574 500 1575
rect 494 1570 495 1574
rect 499 1570 500 1574
rect 494 1569 500 1570
rect 590 1574 596 1575
rect 590 1570 591 1574
rect 595 1570 596 1574
rect 590 1569 596 1570
rect 686 1574 692 1575
rect 686 1570 687 1574
rect 691 1570 692 1574
rect 686 1569 692 1570
rect 782 1574 788 1575
rect 782 1570 783 1574
rect 787 1570 788 1574
rect 782 1569 788 1570
rect 878 1574 884 1575
rect 878 1570 879 1574
rect 883 1570 884 1574
rect 878 1569 884 1570
rect 974 1574 980 1575
rect 974 1570 975 1574
rect 979 1570 980 1574
rect 974 1569 980 1570
rect 1078 1574 1084 1575
rect 1078 1570 1079 1574
rect 1083 1570 1084 1574
rect 1078 1569 1084 1570
rect 1190 1574 1196 1575
rect 1190 1570 1191 1574
rect 1195 1570 1196 1574
rect 1190 1569 1196 1570
rect 1286 1574 1292 1575
rect 1286 1570 1287 1574
rect 1291 1570 1292 1574
rect 1286 1569 1292 1570
rect 160 1559 162 1569
rect 264 1559 266 1569
rect 384 1559 386 1569
rect 496 1559 498 1569
rect 592 1559 594 1569
rect 688 1559 690 1569
rect 784 1559 786 1569
rect 880 1559 882 1569
rect 976 1559 978 1569
rect 1080 1559 1082 1569
rect 1192 1559 1194 1569
rect 1288 1559 1290 1569
rect 1328 1559 1330 1578
rect 1366 1567 1372 1568
rect 1366 1563 1367 1567
rect 1371 1563 1372 1567
rect 1366 1562 1372 1563
rect 2582 1567 2588 1568
rect 2582 1563 2583 1567
rect 2587 1563 2588 1567
rect 2582 1562 2588 1563
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 159 1558 163 1559
rect 159 1553 163 1554
rect 231 1558 235 1559
rect 231 1553 235 1554
rect 263 1558 267 1559
rect 263 1553 267 1554
rect 335 1558 339 1559
rect 335 1553 339 1554
rect 383 1558 387 1559
rect 383 1553 387 1554
rect 455 1558 459 1559
rect 455 1553 459 1554
rect 495 1558 499 1559
rect 495 1553 499 1554
rect 583 1558 587 1559
rect 583 1553 587 1554
rect 591 1558 595 1559
rect 591 1553 595 1554
rect 687 1558 691 1559
rect 687 1553 691 1554
rect 719 1558 723 1559
rect 719 1553 723 1554
rect 783 1558 787 1559
rect 783 1553 787 1554
rect 863 1558 867 1559
rect 863 1553 867 1554
rect 879 1558 883 1559
rect 879 1553 883 1554
rect 975 1558 979 1559
rect 975 1553 979 1554
rect 1007 1558 1011 1559
rect 1007 1553 1011 1554
rect 1079 1558 1083 1559
rect 1079 1553 1083 1554
rect 1151 1558 1155 1559
rect 1151 1553 1155 1554
rect 1191 1558 1195 1559
rect 1191 1553 1195 1554
rect 1287 1558 1291 1559
rect 1287 1553 1291 1554
rect 1327 1558 1331 1559
rect 1327 1553 1331 1554
rect 112 1538 114 1553
rect 160 1547 162 1553
rect 232 1547 234 1553
rect 336 1547 338 1553
rect 456 1547 458 1553
rect 584 1547 586 1553
rect 720 1547 722 1553
rect 864 1547 866 1553
rect 1008 1547 1010 1553
rect 1152 1547 1154 1553
rect 1288 1547 1290 1553
rect 158 1546 164 1547
rect 158 1542 159 1546
rect 163 1542 164 1546
rect 158 1541 164 1542
rect 230 1546 236 1547
rect 230 1542 231 1546
rect 235 1542 236 1546
rect 230 1541 236 1542
rect 334 1546 340 1547
rect 334 1542 335 1546
rect 339 1542 340 1546
rect 334 1541 340 1542
rect 454 1546 460 1547
rect 454 1542 455 1546
rect 459 1542 460 1546
rect 454 1541 460 1542
rect 582 1546 588 1547
rect 582 1542 583 1546
rect 587 1542 588 1546
rect 582 1541 588 1542
rect 718 1546 724 1547
rect 718 1542 719 1546
rect 723 1542 724 1546
rect 718 1541 724 1542
rect 862 1546 868 1547
rect 862 1542 863 1546
rect 867 1542 868 1546
rect 862 1541 868 1542
rect 1006 1546 1012 1547
rect 1006 1542 1007 1546
rect 1011 1542 1012 1546
rect 1006 1541 1012 1542
rect 1150 1546 1156 1547
rect 1150 1542 1151 1546
rect 1155 1542 1156 1546
rect 1150 1541 1156 1542
rect 1286 1546 1292 1547
rect 1286 1542 1287 1546
rect 1291 1542 1292 1546
rect 1286 1541 1292 1542
rect 1328 1538 1330 1553
rect 1368 1543 1370 1562
rect 1414 1558 1420 1559
rect 1414 1554 1415 1558
rect 1419 1554 1420 1558
rect 1414 1553 1420 1554
rect 1510 1558 1516 1559
rect 1510 1554 1511 1558
rect 1515 1554 1516 1558
rect 1510 1553 1516 1554
rect 1630 1558 1636 1559
rect 1630 1554 1631 1558
rect 1635 1554 1636 1558
rect 1630 1553 1636 1554
rect 1758 1558 1764 1559
rect 1758 1554 1759 1558
rect 1763 1554 1764 1558
rect 1758 1553 1764 1554
rect 1878 1558 1884 1559
rect 1878 1554 1879 1558
rect 1883 1554 1884 1558
rect 1878 1553 1884 1554
rect 1998 1558 2004 1559
rect 1998 1554 1999 1558
rect 2003 1554 2004 1558
rect 1998 1553 2004 1554
rect 2110 1558 2116 1559
rect 2110 1554 2111 1558
rect 2115 1554 2116 1558
rect 2110 1553 2116 1554
rect 2214 1558 2220 1559
rect 2214 1554 2215 1558
rect 2219 1554 2220 1558
rect 2214 1553 2220 1554
rect 2310 1558 2316 1559
rect 2310 1554 2311 1558
rect 2315 1554 2316 1558
rect 2310 1553 2316 1554
rect 2406 1558 2412 1559
rect 2406 1554 2407 1558
rect 2411 1554 2412 1558
rect 2406 1553 2412 1554
rect 2510 1558 2516 1559
rect 2510 1554 2511 1558
rect 2515 1554 2516 1558
rect 2510 1553 2516 1554
rect 1416 1543 1418 1553
rect 1512 1543 1514 1553
rect 1632 1543 1634 1553
rect 1760 1543 1762 1553
rect 1880 1543 1882 1553
rect 2000 1543 2002 1553
rect 2112 1543 2114 1553
rect 2216 1543 2218 1553
rect 2312 1543 2314 1553
rect 2408 1543 2410 1553
rect 2512 1543 2514 1553
rect 2584 1543 2586 1562
rect 1367 1542 1371 1543
rect 110 1537 116 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 110 1532 116 1533
rect 1326 1537 1332 1538
rect 1367 1537 1371 1538
rect 1415 1542 1419 1543
rect 1415 1537 1419 1538
rect 1511 1542 1515 1543
rect 1511 1537 1515 1538
rect 1527 1542 1531 1543
rect 1527 1537 1531 1538
rect 1631 1542 1635 1543
rect 1631 1537 1635 1538
rect 1647 1542 1651 1543
rect 1647 1537 1651 1538
rect 1759 1542 1763 1543
rect 1759 1537 1763 1538
rect 1767 1542 1771 1543
rect 1767 1537 1771 1538
rect 1879 1542 1883 1543
rect 1879 1537 1883 1538
rect 1983 1542 1987 1543
rect 1983 1537 1987 1538
rect 1999 1542 2003 1543
rect 1999 1537 2003 1538
rect 2079 1542 2083 1543
rect 2079 1537 2083 1538
rect 2111 1542 2115 1543
rect 2111 1537 2115 1538
rect 2167 1542 2171 1543
rect 2167 1537 2171 1538
rect 2215 1542 2219 1543
rect 2215 1537 2219 1538
rect 2255 1542 2259 1543
rect 2255 1537 2259 1538
rect 2311 1542 2315 1543
rect 2311 1537 2315 1538
rect 2335 1542 2339 1543
rect 2335 1537 2339 1538
rect 2407 1542 2411 1543
rect 2407 1537 2411 1538
rect 2487 1542 2491 1543
rect 2487 1537 2491 1538
rect 2511 1542 2515 1543
rect 2511 1537 2515 1538
rect 2543 1542 2547 1543
rect 2543 1537 2547 1538
rect 2583 1542 2587 1543
rect 2583 1537 2587 1538
rect 1326 1533 1327 1537
rect 1331 1533 1332 1537
rect 1326 1532 1332 1533
rect 1368 1522 1370 1537
rect 1416 1531 1418 1537
rect 1528 1531 1530 1537
rect 1648 1531 1650 1537
rect 1768 1531 1770 1537
rect 1880 1531 1882 1537
rect 1984 1531 1986 1537
rect 2080 1531 2082 1537
rect 2168 1531 2170 1537
rect 2256 1531 2258 1537
rect 2336 1531 2338 1537
rect 2408 1531 2410 1537
rect 2488 1531 2490 1537
rect 2544 1531 2546 1537
rect 1414 1530 1420 1531
rect 1414 1526 1415 1530
rect 1419 1526 1420 1530
rect 1414 1525 1420 1526
rect 1526 1530 1532 1531
rect 1526 1526 1527 1530
rect 1531 1526 1532 1530
rect 1526 1525 1532 1526
rect 1646 1530 1652 1531
rect 1646 1526 1647 1530
rect 1651 1526 1652 1530
rect 1646 1525 1652 1526
rect 1766 1530 1772 1531
rect 1766 1526 1767 1530
rect 1771 1526 1772 1530
rect 1766 1525 1772 1526
rect 1878 1530 1884 1531
rect 1878 1526 1879 1530
rect 1883 1526 1884 1530
rect 1878 1525 1884 1526
rect 1982 1530 1988 1531
rect 1982 1526 1983 1530
rect 1987 1526 1988 1530
rect 1982 1525 1988 1526
rect 2078 1530 2084 1531
rect 2078 1526 2079 1530
rect 2083 1526 2084 1530
rect 2078 1525 2084 1526
rect 2166 1530 2172 1531
rect 2166 1526 2167 1530
rect 2171 1526 2172 1530
rect 2166 1525 2172 1526
rect 2254 1530 2260 1531
rect 2254 1526 2255 1530
rect 2259 1526 2260 1530
rect 2254 1525 2260 1526
rect 2334 1530 2340 1531
rect 2334 1526 2335 1530
rect 2339 1526 2340 1530
rect 2334 1525 2340 1526
rect 2406 1530 2412 1531
rect 2406 1526 2407 1530
rect 2411 1526 2412 1530
rect 2406 1525 2412 1526
rect 2486 1530 2492 1531
rect 2486 1526 2487 1530
rect 2491 1526 2492 1530
rect 2486 1525 2492 1526
rect 2542 1530 2548 1531
rect 2542 1526 2543 1530
rect 2547 1526 2548 1530
rect 2542 1525 2548 1526
rect 2584 1522 2586 1537
rect 1366 1521 1372 1522
rect 110 1520 116 1521
rect 1326 1520 1332 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 110 1515 116 1516
rect 142 1519 148 1520
rect 142 1515 143 1519
rect 147 1515 148 1519
rect 112 1503 114 1515
rect 142 1514 148 1515
rect 214 1519 220 1520
rect 214 1515 215 1519
rect 219 1515 220 1519
rect 214 1514 220 1515
rect 318 1519 324 1520
rect 318 1515 319 1519
rect 323 1515 324 1519
rect 318 1514 324 1515
rect 438 1519 444 1520
rect 438 1515 439 1519
rect 443 1515 444 1519
rect 438 1514 444 1515
rect 566 1519 572 1520
rect 566 1515 567 1519
rect 571 1515 572 1519
rect 566 1514 572 1515
rect 702 1519 708 1520
rect 702 1515 703 1519
rect 707 1515 708 1519
rect 702 1514 708 1515
rect 846 1519 852 1520
rect 846 1515 847 1519
rect 851 1515 852 1519
rect 846 1514 852 1515
rect 990 1519 996 1520
rect 990 1515 991 1519
rect 995 1515 996 1519
rect 990 1514 996 1515
rect 1134 1519 1140 1520
rect 1134 1515 1135 1519
rect 1139 1515 1140 1519
rect 1134 1514 1140 1515
rect 1270 1519 1276 1520
rect 1270 1515 1271 1519
rect 1275 1515 1276 1519
rect 1326 1516 1327 1520
rect 1331 1516 1332 1520
rect 1366 1517 1367 1521
rect 1371 1517 1372 1521
rect 1366 1516 1372 1517
rect 2582 1521 2588 1522
rect 2582 1517 2583 1521
rect 2587 1517 2588 1521
rect 2582 1516 2588 1517
rect 1326 1515 1332 1516
rect 1270 1514 1276 1515
rect 144 1503 146 1514
rect 216 1503 218 1514
rect 320 1503 322 1514
rect 440 1503 442 1514
rect 568 1503 570 1514
rect 704 1503 706 1514
rect 848 1503 850 1514
rect 992 1503 994 1514
rect 1136 1503 1138 1514
rect 1272 1503 1274 1514
rect 1328 1503 1330 1515
rect 1366 1504 1372 1505
rect 2582 1504 2588 1505
rect 111 1502 115 1503
rect 111 1497 115 1498
rect 143 1502 147 1503
rect 143 1497 147 1498
rect 199 1502 203 1503
rect 199 1497 203 1498
rect 215 1502 219 1503
rect 215 1497 219 1498
rect 271 1502 275 1503
rect 271 1497 275 1498
rect 319 1502 323 1503
rect 319 1497 323 1498
rect 367 1502 371 1503
rect 367 1497 371 1498
rect 439 1502 443 1503
rect 439 1497 443 1498
rect 479 1502 483 1503
rect 479 1497 483 1498
rect 567 1502 571 1503
rect 567 1497 571 1498
rect 591 1502 595 1503
rect 591 1497 595 1498
rect 703 1502 707 1503
rect 703 1497 707 1498
rect 807 1502 811 1503
rect 807 1497 811 1498
rect 847 1502 851 1503
rect 847 1497 851 1498
rect 911 1502 915 1503
rect 911 1497 915 1498
rect 991 1502 995 1503
rect 991 1497 995 1498
rect 1007 1502 1011 1503
rect 1007 1497 1011 1498
rect 1103 1502 1107 1503
rect 1103 1497 1107 1498
rect 1135 1502 1139 1503
rect 1135 1497 1139 1498
rect 1199 1502 1203 1503
rect 1199 1497 1203 1498
rect 1271 1502 1275 1503
rect 1271 1497 1275 1498
rect 1327 1502 1331 1503
rect 1366 1500 1367 1504
rect 1371 1500 1372 1504
rect 1366 1499 1372 1500
rect 1398 1503 1404 1504
rect 1398 1499 1399 1503
rect 1403 1499 1404 1503
rect 1327 1497 1331 1498
rect 112 1485 114 1497
rect 144 1486 146 1497
rect 200 1486 202 1497
rect 272 1486 274 1497
rect 368 1486 370 1497
rect 480 1486 482 1497
rect 592 1486 594 1497
rect 704 1486 706 1497
rect 808 1486 810 1497
rect 912 1486 914 1497
rect 1008 1486 1010 1497
rect 1104 1486 1106 1497
rect 1200 1486 1202 1497
rect 1272 1486 1274 1497
rect 142 1485 148 1486
rect 110 1484 116 1485
rect 110 1480 111 1484
rect 115 1480 116 1484
rect 142 1481 143 1485
rect 147 1481 148 1485
rect 142 1480 148 1481
rect 198 1485 204 1486
rect 198 1481 199 1485
rect 203 1481 204 1485
rect 198 1480 204 1481
rect 270 1485 276 1486
rect 270 1481 271 1485
rect 275 1481 276 1485
rect 270 1480 276 1481
rect 366 1485 372 1486
rect 366 1481 367 1485
rect 371 1481 372 1485
rect 366 1480 372 1481
rect 478 1485 484 1486
rect 478 1481 479 1485
rect 483 1481 484 1485
rect 478 1480 484 1481
rect 590 1485 596 1486
rect 590 1481 591 1485
rect 595 1481 596 1485
rect 590 1480 596 1481
rect 702 1485 708 1486
rect 702 1481 703 1485
rect 707 1481 708 1485
rect 702 1480 708 1481
rect 806 1485 812 1486
rect 806 1481 807 1485
rect 811 1481 812 1485
rect 806 1480 812 1481
rect 910 1485 916 1486
rect 910 1481 911 1485
rect 915 1481 916 1485
rect 910 1480 916 1481
rect 1006 1485 1012 1486
rect 1006 1481 1007 1485
rect 1011 1481 1012 1485
rect 1006 1480 1012 1481
rect 1102 1485 1108 1486
rect 1102 1481 1103 1485
rect 1107 1481 1108 1485
rect 1102 1480 1108 1481
rect 1198 1485 1204 1486
rect 1198 1481 1199 1485
rect 1203 1481 1204 1485
rect 1198 1480 1204 1481
rect 1270 1485 1276 1486
rect 1328 1485 1330 1497
rect 1270 1481 1271 1485
rect 1275 1481 1276 1485
rect 1270 1480 1276 1481
rect 1326 1484 1332 1485
rect 1326 1480 1327 1484
rect 1331 1480 1332 1484
rect 110 1479 116 1480
rect 1326 1479 1332 1480
rect 1368 1479 1370 1499
rect 1398 1498 1404 1499
rect 1510 1503 1516 1504
rect 1510 1499 1511 1503
rect 1515 1499 1516 1503
rect 1510 1498 1516 1499
rect 1630 1503 1636 1504
rect 1630 1499 1631 1503
rect 1635 1499 1636 1503
rect 1630 1498 1636 1499
rect 1750 1503 1756 1504
rect 1750 1499 1751 1503
rect 1755 1499 1756 1503
rect 1750 1498 1756 1499
rect 1862 1503 1868 1504
rect 1862 1499 1863 1503
rect 1867 1499 1868 1503
rect 1862 1498 1868 1499
rect 1966 1503 1972 1504
rect 1966 1499 1967 1503
rect 1971 1499 1972 1503
rect 1966 1498 1972 1499
rect 2062 1503 2068 1504
rect 2062 1499 2063 1503
rect 2067 1499 2068 1503
rect 2062 1498 2068 1499
rect 2150 1503 2156 1504
rect 2150 1499 2151 1503
rect 2155 1499 2156 1503
rect 2150 1498 2156 1499
rect 2238 1503 2244 1504
rect 2238 1499 2239 1503
rect 2243 1499 2244 1503
rect 2238 1498 2244 1499
rect 2318 1503 2324 1504
rect 2318 1499 2319 1503
rect 2323 1499 2324 1503
rect 2318 1498 2324 1499
rect 2390 1503 2396 1504
rect 2390 1499 2391 1503
rect 2395 1499 2396 1503
rect 2390 1498 2396 1499
rect 2470 1503 2476 1504
rect 2470 1499 2471 1503
rect 2475 1499 2476 1503
rect 2470 1498 2476 1499
rect 2526 1503 2532 1504
rect 2526 1499 2527 1503
rect 2531 1499 2532 1503
rect 2582 1500 2583 1504
rect 2587 1500 2588 1504
rect 2582 1499 2588 1500
rect 2526 1498 2532 1499
rect 1400 1479 1402 1498
rect 1512 1479 1514 1498
rect 1632 1479 1634 1498
rect 1752 1479 1754 1498
rect 1864 1479 1866 1498
rect 1968 1479 1970 1498
rect 2064 1479 2066 1498
rect 2152 1479 2154 1498
rect 2240 1479 2242 1498
rect 2320 1479 2322 1498
rect 2392 1479 2394 1498
rect 2472 1479 2474 1498
rect 2528 1479 2530 1498
rect 2584 1479 2586 1499
rect 1367 1478 1371 1479
rect 1367 1473 1371 1474
rect 1399 1478 1403 1479
rect 1399 1473 1403 1474
rect 1503 1478 1507 1479
rect 1503 1473 1507 1474
rect 1511 1478 1515 1479
rect 1511 1473 1515 1474
rect 1631 1478 1635 1479
rect 1631 1473 1635 1474
rect 1751 1478 1755 1479
rect 1751 1473 1755 1474
rect 1863 1478 1867 1479
rect 1863 1473 1867 1474
rect 1871 1478 1875 1479
rect 1871 1473 1875 1474
rect 1967 1478 1971 1479
rect 1967 1473 1971 1474
rect 1983 1478 1987 1479
rect 1983 1473 1987 1474
rect 2063 1478 2067 1479
rect 2063 1473 2067 1474
rect 2087 1478 2091 1479
rect 2087 1473 2091 1474
rect 2151 1478 2155 1479
rect 2151 1473 2155 1474
rect 2183 1478 2187 1479
rect 2183 1473 2187 1474
rect 2239 1478 2243 1479
rect 2239 1473 2243 1474
rect 2271 1478 2275 1479
rect 2271 1473 2275 1474
rect 2319 1478 2323 1479
rect 2319 1473 2323 1474
rect 2359 1478 2363 1479
rect 2359 1473 2363 1474
rect 2391 1478 2395 1479
rect 2391 1473 2395 1474
rect 2455 1478 2459 1479
rect 2455 1473 2459 1474
rect 2471 1478 2475 1479
rect 2471 1473 2475 1474
rect 2527 1478 2531 1479
rect 2527 1473 2531 1474
rect 2583 1478 2587 1479
rect 2583 1473 2587 1474
rect 110 1467 116 1468
rect 110 1463 111 1467
rect 115 1463 116 1467
rect 110 1462 116 1463
rect 1326 1467 1332 1468
rect 1326 1463 1327 1467
rect 1331 1463 1332 1467
rect 1326 1462 1332 1463
rect 112 1443 114 1462
rect 158 1458 164 1459
rect 158 1454 159 1458
rect 163 1454 164 1458
rect 158 1453 164 1454
rect 214 1458 220 1459
rect 214 1454 215 1458
rect 219 1454 220 1458
rect 214 1453 220 1454
rect 286 1458 292 1459
rect 286 1454 287 1458
rect 291 1454 292 1458
rect 286 1453 292 1454
rect 382 1458 388 1459
rect 382 1454 383 1458
rect 387 1454 388 1458
rect 382 1453 388 1454
rect 494 1458 500 1459
rect 494 1454 495 1458
rect 499 1454 500 1458
rect 494 1453 500 1454
rect 606 1458 612 1459
rect 606 1454 607 1458
rect 611 1454 612 1458
rect 606 1453 612 1454
rect 718 1458 724 1459
rect 718 1454 719 1458
rect 723 1454 724 1458
rect 718 1453 724 1454
rect 822 1458 828 1459
rect 822 1454 823 1458
rect 827 1454 828 1458
rect 822 1453 828 1454
rect 926 1458 932 1459
rect 926 1454 927 1458
rect 931 1454 932 1458
rect 926 1453 932 1454
rect 1022 1458 1028 1459
rect 1022 1454 1023 1458
rect 1027 1454 1028 1458
rect 1022 1453 1028 1454
rect 1118 1458 1124 1459
rect 1118 1454 1119 1458
rect 1123 1454 1124 1458
rect 1118 1453 1124 1454
rect 1214 1458 1220 1459
rect 1214 1454 1215 1458
rect 1219 1454 1220 1458
rect 1214 1453 1220 1454
rect 1286 1458 1292 1459
rect 1286 1454 1287 1458
rect 1291 1454 1292 1458
rect 1286 1453 1292 1454
rect 160 1443 162 1453
rect 216 1443 218 1453
rect 288 1443 290 1453
rect 384 1443 386 1453
rect 496 1443 498 1453
rect 608 1443 610 1453
rect 720 1443 722 1453
rect 824 1443 826 1453
rect 928 1443 930 1453
rect 1024 1443 1026 1453
rect 1120 1443 1122 1453
rect 1216 1443 1218 1453
rect 1288 1443 1290 1453
rect 1328 1443 1330 1462
rect 1368 1461 1370 1473
rect 1400 1462 1402 1473
rect 1504 1462 1506 1473
rect 1632 1462 1634 1473
rect 1752 1462 1754 1473
rect 1872 1462 1874 1473
rect 1984 1462 1986 1473
rect 2088 1462 2090 1473
rect 2184 1462 2186 1473
rect 2272 1462 2274 1473
rect 2360 1462 2362 1473
rect 2456 1462 2458 1473
rect 2528 1462 2530 1473
rect 1398 1461 1404 1462
rect 1366 1460 1372 1461
rect 1366 1456 1367 1460
rect 1371 1456 1372 1460
rect 1398 1457 1399 1461
rect 1403 1457 1404 1461
rect 1398 1456 1404 1457
rect 1502 1461 1508 1462
rect 1502 1457 1503 1461
rect 1507 1457 1508 1461
rect 1502 1456 1508 1457
rect 1630 1461 1636 1462
rect 1630 1457 1631 1461
rect 1635 1457 1636 1461
rect 1630 1456 1636 1457
rect 1750 1461 1756 1462
rect 1750 1457 1751 1461
rect 1755 1457 1756 1461
rect 1750 1456 1756 1457
rect 1870 1461 1876 1462
rect 1870 1457 1871 1461
rect 1875 1457 1876 1461
rect 1870 1456 1876 1457
rect 1982 1461 1988 1462
rect 1982 1457 1983 1461
rect 1987 1457 1988 1461
rect 1982 1456 1988 1457
rect 2086 1461 2092 1462
rect 2086 1457 2087 1461
rect 2091 1457 2092 1461
rect 2086 1456 2092 1457
rect 2182 1461 2188 1462
rect 2182 1457 2183 1461
rect 2187 1457 2188 1461
rect 2182 1456 2188 1457
rect 2270 1461 2276 1462
rect 2270 1457 2271 1461
rect 2275 1457 2276 1461
rect 2270 1456 2276 1457
rect 2358 1461 2364 1462
rect 2358 1457 2359 1461
rect 2363 1457 2364 1461
rect 2358 1456 2364 1457
rect 2454 1461 2460 1462
rect 2454 1457 2455 1461
rect 2459 1457 2460 1461
rect 2454 1456 2460 1457
rect 2526 1461 2532 1462
rect 2584 1461 2586 1473
rect 2526 1457 2527 1461
rect 2531 1457 2532 1461
rect 2526 1456 2532 1457
rect 2582 1460 2588 1461
rect 2582 1456 2583 1460
rect 2587 1456 2588 1460
rect 1366 1455 1372 1456
rect 2582 1455 2588 1456
rect 1366 1443 1372 1444
rect 111 1442 115 1443
rect 111 1437 115 1438
rect 159 1442 163 1443
rect 159 1437 163 1438
rect 215 1442 219 1443
rect 215 1437 219 1438
rect 255 1442 259 1443
rect 255 1437 259 1438
rect 287 1442 291 1443
rect 287 1437 291 1438
rect 311 1442 315 1443
rect 311 1437 315 1438
rect 375 1442 379 1443
rect 375 1437 379 1438
rect 383 1442 387 1443
rect 383 1437 387 1438
rect 447 1442 451 1443
rect 447 1437 451 1438
rect 495 1442 499 1443
rect 495 1437 499 1438
rect 527 1442 531 1443
rect 527 1437 531 1438
rect 607 1442 611 1443
rect 607 1437 611 1438
rect 695 1442 699 1443
rect 695 1437 699 1438
rect 719 1442 723 1443
rect 719 1437 723 1438
rect 783 1442 787 1443
rect 783 1437 787 1438
rect 823 1442 827 1443
rect 823 1437 827 1438
rect 871 1442 875 1443
rect 871 1437 875 1438
rect 927 1442 931 1443
rect 927 1437 931 1438
rect 959 1442 963 1443
rect 959 1437 963 1438
rect 1023 1442 1027 1443
rect 1023 1437 1027 1438
rect 1055 1442 1059 1443
rect 1055 1437 1059 1438
rect 1119 1442 1123 1443
rect 1119 1437 1123 1438
rect 1151 1442 1155 1443
rect 1151 1437 1155 1438
rect 1215 1442 1219 1443
rect 1215 1437 1219 1438
rect 1287 1442 1291 1443
rect 1287 1437 1291 1438
rect 1327 1442 1331 1443
rect 1366 1439 1367 1443
rect 1371 1439 1372 1443
rect 1366 1438 1372 1439
rect 2582 1443 2588 1444
rect 2582 1439 2583 1443
rect 2587 1439 2588 1443
rect 2582 1438 2588 1439
rect 1327 1437 1331 1438
rect 112 1422 114 1437
rect 256 1431 258 1437
rect 312 1431 314 1437
rect 376 1431 378 1437
rect 448 1431 450 1437
rect 528 1431 530 1437
rect 608 1431 610 1437
rect 696 1431 698 1437
rect 784 1431 786 1437
rect 872 1431 874 1437
rect 960 1431 962 1437
rect 1056 1431 1058 1437
rect 1152 1431 1154 1437
rect 254 1430 260 1431
rect 254 1426 255 1430
rect 259 1426 260 1430
rect 254 1425 260 1426
rect 310 1430 316 1431
rect 310 1426 311 1430
rect 315 1426 316 1430
rect 310 1425 316 1426
rect 374 1430 380 1431
rect 374 1426 375 1430
rect 379 1426 380 1430
rect 374 1425 380 1426
rect 446 1430 452 1431
rect 446 1426 447 1430
rect 451 1426 452 1430
rect 446 1425 452 1426
rect 526 1430 532 1431
rect 526 1426 527 1430
rect 531 1426 532 1430
rect 526 1425 532 1426
rect 606 1430 612 1431
rect 606 1426 607 1430
rect 611 1426 612 1430
rect 606 1425 612 1426
rect 694 1430 700 1431
rect 694 1426 695 1430
rect 699 1426 700 1430
rect 694 1425 700 1426
rect 782 1430 788 1431
rect 782 1426 783 1430
rect 787 1426 788 1430
rect 782 1425 788 1426
rect 870 1430 876 1431
rect 870 1426 871 1430
rect 875 1426 876 1430
rect 870 1425 876 1426
rect 958 1430 964 1431
rect 958 1426 959 1430
rect 963 1426 964 1430
rect 958 1425 964 1426
rect 1054 1430 1060 1431
rect 1054 1426 1055 1430
rect 1059 1426 1060 1430
rect 1054 1425 1060 1426
rect 1150 1430 1156 1431
rect 1150 1426 1151 1430
rect 1155 1426 1156 1430
rect 1150 1425 1156 1426
rect 1328 1422 1330 1437
rect 110 1421 116 1422
rect 110 1417 111 1421
rect 115 1417 116 1421
rect 110 1416 116 1417
rect 1326 1421 1332 1422
rect 1326 1417 1327 1421
rect 1331 1417 1332 1421
rect 1368 1419 1370 1438
rect 1414 1434 1420 1435
rect 1414 1430 1415 1434
rect 1419 1430 1420 1434
rect 1414 1429 1420 1430
rect 1518 1434 1524 1435
rect 1518 1430 1519 1434
rect 1523 1430 1524 1434
rect 1518 1429 1524 1430
rect 1646 1434 1652 1435
rect 1646 1430 1647 1434
rect 1651 1430 1652 1434
rect 1646 1429 1652 1430
rect 1766 1434 1772 1435
rect 1766 1430 1767 1434
rect 1771 1430 1772 1434
rect 1766 1429 1772 1430
rect 1886 1434 1892 1435
rect 1886 1430 1887 1434
rect 1891 1430 1892 1434
rect 1886 1429 1892 1430
rect 1998 1434 2004 1435
rect 1998 1430 1999 1434
rect 2003 1430 2004 1434
rect 1998 1429 2004 1430
rect 2102 1434 2108 1435
rect 2102 1430 2103 1434
rect 2107 1430 2108 1434
rect 2102 1429 2108 1430
rect 2198 1434 2204 1435
rect 2198 1430 2199 1434
rect 2203 1430 2204 1434
rect 2198 1429 2204 1430
rect 2286 1434 2292 1435
rect 2286 1430 2287 1434
rect 2291 1430 2292 1434
rect 2286 1429 2292 1430
rect 2374 1434 2380 1435
rect 2374 1430 2375 1434
rect 2379 1430 2380 1434
rect 2374 1429 2380 1430
rect 2470 1434 2476 1435
rect 2470 1430 2471 1434
rect 2475 1430 2476 1434
rect 2470 1429 2476 1430
rect 2542 1434 2548 1435
rect 2542 1430 2543 1434
rect 2547 1430 2548 1434
rect 2542 1429 2548 1430
rect 1416 1419 1418 1429
rect 1520 1419 1522 1429
rect 1648 1419 1650 1429
rect 1768 1419 1770 1429
rect 1888 1419 1890 1429
rect 2000 1419 2002 1429
rect 2104 1419 2106 1429
rect 2200 1419 2202 1429
rect 2288 1419 2290 1429
rect 2376 1419 2378 1429
rect 2472 1419 2474 1429
rect 2544 1419 2546 1429
rect 2584 1419 2586 1438
rect 1326 1416 1332 1417
rect 1367 1418 1371 1419
rect 1367 1413 1371 1414
rect 1415 1418 1419 1419
rect 1415 1413 1419 1414
rect 1471 1418 1475 1419
rect 1471 1413 1475 1414
rect 1519 1418 1523 1419
rect 1519 1413 1523 1414
rect 1551 1418 1555 1419
rect 1551 1413 1555 1414
rect 1631 1418 1635 1419
rect 1631 1413 1635 1414
rect 1647 1418 1651 1419
rect 1647 1413 1651 1414
rect 1711 1418 1715 1419
rect 1711 1413 1715 1414
rect 1767 1418 1771 1419
rect 1767 1413 1771 1414
rect 1791 1418 1795 1419
rect 1791 1413 1795 1414
rect 1871 1418 1875 1419
rect 1871 1413 1875 1414
rect 1887 1418 1891 1419
rect 1887 1413 1891 1414
rect 1959 1418 1963 1419
rect 1959 1413 1963 1414
rect 1999 1418 2003 1419
rect 1999 1413 2003 1414
rect 2055 1418 2059 1419
rect 2055 1413 2059 1414
rect 2103 1418 2107 1419
rect 2103 1413 2107 1414
rect 2167 1418 2171 1419
rect 2167 1413 2171 1414
rect 2199 1418 2203 1419
rect 2199 1413 2203 1414
rect 2287 1418 2291 1419
rect 2287 1413 2291 1414
rect 2295 1418 2299 1419
rect 2295 1413 2299 1414
rect 2375 1418 2379 1419
rect 2375 1413 2379 1414
rect 2431 1418 2435 1419
rect 2431 1413 2435 1414
rect 2471 1418 2475 1419
rect 2471 1413 2475 1414
rect 2543 1418 2547 1419
rect 2543 1413 2547 1414
rect 2583 1418 2587 1419
rect 2583 1413 2587 1414
rect 110 1404 116 1405
rect 1326 1404 1332 1405
rect 110 1400 111 1404
rect 115 1400 116 1404
rect 110 1399 116 1400
rect 238 1403 244 1404
rect 238 1399 239 1403
rect 243 1399 244 1403
rect 112 1379 114 1399
rect 238 1398 244 1399
rect 294 1403 300 1404
rect 294 1399 295 1403
rect 299 1399 300 1403
rect 294 1398 300 1399
rect 358 1403 364 1404
rect 358 1399 359 1403
rect 363 1399 364 1403
rect 358 1398 364 1399
rect 430 1403 436 1404
rect 430 1399 431 1403
rect 435 1399 436 1403
rect 430 1398 436 1399
rect 510 1403 516 1404
rect 510 1399 511 1403
rect 515 1399 516 1403
rect 510 1398 516 1399
rect 590 1403 596 1404
rect 590 1399 591 1403
rect 595 1399 596 1403
rect 590 1398 596 1399
rect 678 1403 684 1404
rect 678 1399 679 1403
rect 683 1399 684 1403
rect 678 1398 684 1399
rect 766 1403 772 1404
rect 766 1399 767 1403
rect 771 1399 772 1403
rect 766 1398 772 1399
rect 854 1403 860 1404
rect 854 1399 855 1403
rect 859 1399 860 1403
rect 854 1398 860 1399
rect 942 1403 948 1404
rect 942 1399 943 1403
rect 947 1399 948 1403
rect 942 1398 948 1399
rect 1038 1403 1044 1404
rect 1038 1399 1039 1403
rect 1043 1399 1044 1403
rect 1038 1398 1044 1399
rect 1134 1403 1140 1404
rect 1134 1399 1135 1403
rect 1139 1399 1140 1403
rect 1326 1400 1327 1404
rect 1331 1400 1332 1404
rect 1326 1399 1332 1400
rect 1134 1398 1140 1399
rect 240 1379 242 1398
rect 296 1379 298 1398
rect 360 1379 362 1398
rect 432 1379 434 1398
rect 512 1379 514 1398
rect 592 1379 594 1398
rect 680 1379 682 1398
rect 768 1379 770 1398
rect 856 1379 858 1398
rect 944 1379 946 1398
rect 1040 1379 1042 1398
rect 1136 1379 1138 1398
rect 1328 1379 1330 1399
rect 1368 1398 1370 1413
rect 1416 1407 1418 1413
rect 1472 1407 1474 1413
rect 1552 1407 1554 1413
rect 1632 1407 1634 1413
rect 1712 1407 1714 1413
rect 1792 1407 1794 1413
rect 1872 1407 1874 1413
rect 1960 1407 1962 1413
rect 2056 1407 2058 1413
rect 2168 1407 2170 1413
rect 2296 1407 2298 1413
rect 2432 1407 2434 1413
rect 2544 1407 2546 1413
rect 1414 1406 1420 1407
rect 1414 1402 1415 1406
rect 1419 1402 1420 1406
rect 1414 1401 1420 1402
rect 1470 1406 1476 1407
rect 1470 1402 1471 1406
rect 1475 1402 1476 1406
rect 1470 1401 1476 1402
rect 1550 1406 1556 1407
rect 1550 1402 1551 1406
rect 1555 1402 1556 1406
rect 1550 1401 1556 1402
rect 1630 1406 1636 1407
rect 1630 1402 1631 1406
rect 1635 1402 1636 1406
rect 1630 1401 1636 1402
rect 1710 1406 1716 1407
rect 1710 1402 1711 1406
rect 1715 1402 1716 1406
rect 1710 1401 1716 1402
rect 1790 1406 1796 1407
rect 1790 1402 1791 1406
rect 1795 1402 1796 1406
rect 1790 1401 1796 1402
rect 1870 1406 1876 1407
rect 1870 1402 1871 1406
rect 1875 1402 1876 1406
rect 1870 1401 1876 1402
rect 1958 1406 1964 1407
rect 1958 1402 1959 1406
rect 1963 1402 1964 1406
rect 1958 1401 1964 1402
rect 2054 1406 2060 1407
rect 2054 1402 2055 1406
rect 2059 1402 2060 1406
rect 2054 1401 2060 1402
rect 2166 1406 2172 1407
rect 2166 1402 2167 1406
rect 2171 1402 2172 1406
rect 2166 1401 2172 1402
rect 2294 1406 2300 1407
rect 2294 1402 2295 1406
rect 2299 1402 2300 1406
rect 2294 1401 2300 1402
rect 2430 1406 2436 1407
rect 2430 1402 2431 1406
rect 2435 1402 2436 1406
rect 2430 1401 2436 1402
rect 2542 1406 2548 1407
rect 2542 1402 2543 1406
rect 2547 1402 2548 1406
rect 2542 1401 2548 1402
rect 2584 1398 2586 1413
rect 1366 1397 1372 1398
rect 1366 1393 1367 1397
rect 1371 1393 1372 1397
rect 1366 1392 1372 1393
rect 2582 1397 2588 1398
rect 2582 1393 2583 1397
rect 2587 1393 2588 1397
rect 2582 1392 2588 1393
rect 1366 1380 1372 1381
rect 2582 1380 2588 1381
rect 111 1378 115 1379
rect 111 1373 115 1374
rect 239 1378 243 1379
rect 239 1373 243 1374
rect 295 1378 299 1379
rect 295 1373 299 1374
rect 359 1378 363 1379
rect 359 1373 363 1374
rect 415 1378 419 1379
rect 415 1373 419 1374
rect 431 1378 435 1379
rect 431 1373 435 1374
rect 471 1378 475 1379
rect 471 1373 475 1374
rect 511 1378 515 1379
rect 511 1373 515 1374
rect 527 1378 531 1379
rect 527 1373 531 1374
rect 591 1378 595 1379
rect 591 1373 595 1374
rect 671 1378 675 1379
rect 671 1373 675 1374
rect 679 1378 683 1379
rect 679 1373 683 1374
rect 751 1378 755 1379
rect 751 1373 755 1374
rect 767 1378 771 1379
rect 767 1373 771 1374
rect 839 1378 843 1379
rect 839 1373 843 1374
rect 855 1378 859 1379
rect 855 1373 859 1374
rect 935 1378 939 1379
rect 935 1373 939 1374
rect 943 1378 947 1379
rect 943 1373 947 1374
rect 1031 1378 1035 1379
rect 1031 1373 1035 1374
rect 1039 1378 1043 1379
rect 1039 1373 1043 1374
rect 1127 1378 1131 1379
rect 1127 1373 1131 1374
rect 1135 1378 1139 1379
rect 1135 1373 1139 1374
rect 1231 1378 1235 1379
rect 1231 1373 1235 1374
rect 1327 1378 1331 1379
rect 1366 1376 1367 1380
rect 1371 1376 1372 1380
rect 1366 1375 1372 1376
rect 1398 1379 1404 1380
rect 1398 1375 1399 1379
rect 1403 1375 1404 1379
rect 1327 1373 1331 1374
rect 112 1361 114 1373
rect 360 1362 362 1373
rect 416 1362 418 1373
rect 472 1362 474 1373
rect 528 1362 530 1373
rect 592 1362 594 1373
rect 672 1362 674 1373
rect 752 1362 754 1373
rect 840 1362 842 1373
rect 936 1362 938 1373
rect 1032 1362 1034 1373
rect 1128 1362 1130 1373
rect 1232 1362 1234 1373
rect 358 1361 364 1362
rect 110 1360 116 1361
rect 110 1356 111 1360
rect 115 1356 116 1360
rect 358 1357 359 1361
rect 363 1357 364 1361
rect 358 1356 364 1357
rect 414 1361 420 1362
rect 414 1357 415 1361
rect 419 1357 420 1361
rect 414 1356 420 1357
rect 470 1361 476 1362
rect 470 1357 471 1361
rect 475 1357 476 1361
rect 470 1356 476 1357
rect 526 1361 532 1362
rect 526 1357 527 1361
rect 531 1357 532 1361
rect 526 1356 532 1357
rect 590 1361 596 1362
rect 590 1357 591 1361
rect 595 1357 596 1361
rect 590 1356 596 1357
rect 670 1361 676 1362
rect 670 1357 671 1361
rect 675 1357 676 1361
rect 670 1356 676 1357
rect 750 1361 756 1362
rect 750 1357 751 1361
rect 755 1357 756 1361
rect 750 1356 756 1357
rect 838 1361 844 1362
rect 838 1357 839 1361
rect 843 1357 844 1361
rect 838 1356 844 1357
rect 934 1361 940 1362
rect 934 1357 935 1361
rect 939 1357 940 1361
rect 934 1356 940 1357
rect 1030 1361 1036 1362
rect 1030 1357 1031 1361
rect 1035 1357 1036 1361
rect 1030 1356 1036 1357
rect 1126 1361 1132 1362
rect 1126 1357 1127 1361
rect 1131 1357 1132 1361
rect 1126 1356 1132 1357
rect 1230 1361 1236 1362
rect 1328 1361 1330 1373
rect 1368 1363 1370 1375
rect 1398 1374 1404 1375
rect 1454 1379 1460 1380
rect 1454 1375 1455 1379
rect 1459 1375 1460 1379
rect 1454 1374 1460 1375
rect 1534 1379 1540 1380
rect 1534 1375 1535 1379
rect 1539 1375 1540 1379
rect 1534 1374 1540 1375
rect 1614 1379 1620 1380
rect 1614 1375 1615 1379
rect 1619 1375 1620 1379
rect 1614 1374 1620 1375
rect 1694 1379 1700 1380
rect 1694 1375 1695 1379
rect 1699 1375 1700 1379
rect 1694 1374 1700 1375
rect 1774 1379 1780 1380
rect 1774 1375 1775 1379
rect 1779 1375 1780 1379
rect 1774 1374 1780 1375
rect 1854 1379 1860 1380
rect 1854 1375 1855 1379
rect 1859 1375 1860 1379
rect 1854 1374 1860 1375
rect 1942 1379 1948 1380
rect 1942 1375 1943 1379
rect 1947 1375 1948 1379
rect 1942 1374 1948 1375
rect 2038 1379 2044 1380
rect 2038 1375 2039 1379
rect 2043 1375 2044 1379
rect 2038 1374 2044 1375
rect 2150 1379 2156 1380
rect 2150 1375 2151 1379
rect 2155 1375 2156 1379
rect 2150 1374 2156 1375
rect 2278 1379 2284 1380
rect 2278 1375 2279 1379
rect 2283 1375 2284 1379
rect 2278 1374 2284 1375
rect 2414 1379 2420 1380
rect 2414 1375 2415 1379
rect 2419 1375 2420 1379
rect 2414 1374 2420 1375
rect 2526 1379 2532 1380
rect 2526 1375 2527 1379
rect 2531 1375 2532 1379
rect 2582 1376 2583 1380
rect 2587 1376 2588 1380
rect 2582 1375 2588 1376
rect 2526 1374 2532 1375
rect 1400 1363 1402 1374
rect 1456 1363 1458 1374
rect 1536 1363 1538 1374
rect 1616 1363 1618 1374
rect 1696 1363 1698 1374
rect 1776 1363 1778 1374
rect 1856 1363 1858 1374
rect 1944 1363 1946 1374
rect 2040 1363 2042 1374
rect 2152 1363 2154 1374
rect 2280 1363 2282 1374
rect 2416 1363 2418 1374
rect 2528 1363 2530 1374
rect 2584 1363 2586 1375
rect 1367 1362 1371 1363
rect 1230 1357 1231 1361
rect 1235 1357 1236 1361
rect 1230 1356 1236 1357
rect 1326 1360 1332 1361
rect 1326 1356 1327 1360
rect 1331 1356 1332 1360
rect 1367 1357 1371 1358
rect 1399 1362 1403 1363
rect 1399 1357 1403 1358
rect 1423 1362 1427 1363
rect 1423 1357 1427 1358
rect 1455 1362 1459 1363
rect 1455 1357 1459 1358
rect 1495 1362 1499 1363
rect 1495 1357 1499 1358
rect 1535 1362 1539 1363
rect 1535 1357 1539 1358
rect 1575 1362 1579 1363
rect 1575 1357 1579 1358
rect 1615 1362 1619 1363
rect 1615 1357 1619 1358
rect 1655 1362 1659 1363
rect 1655 1357 1659 1358
rect 1695 1362 1699 1363
rect 1695 1357 1699 1358
rect 1759 1362 1763 1363
rect 1759 1357 1763 1358
rect 1775 1362 1779 1363
rect 1775 1357 1779 1358
rect 1855 1362 1859 1363
rect 1855 1357 1859 1358
rect 1879 1362 1883 1363
rect 1879 1357 1883 1358
rect 1943 1362 1947 1363
rect 1943 1357 1947 1358
rect 2023 1362 2027 1363
rect 2023 1357 2027 1358
rect 2039 1362 2043 1363
rect 2039 1357 2043 1358
rect 2151 1362 2155 1363
rect 2151 1357 2155 1358
rect 2183 1362 2187 1363
rect 2183 1357 2187 1358
rect 2279 1362 2283 1363
rect 2279 1357 2283 1358
rect 2359 1362 2363 1363
rect 2359 1357 2363 1358
rect 2415 1362 2419 1363
rect 2415 1357 2419 1358
rect 2527 1362 2531 1363
rect 2527 1357 2531 1358
rect 2583 1362 2587 1363
rect 2583 1357 2587 1358
rect 110 1355 116 1356
rect 1326 1355 1332 1356
rect 1368 1345 1370 1357
rect 1424 1346 1426 1357
rect 1496 1346 1498 1357
rect 1576 1346 1578 1357
rect 1656 1346 1658 1357
rect 1760 1346 1762 1357
rect 1880 1346 1882 1357
rect 2024 1346 2026 1357
rect 2184 1346 2186 1357
rect 2360 1346 2362 1357
rect 2528 1346 2530 1357
rect 1422 1345 1428 1346
rect 1366 1344 1372 1345
rect 110 1343 116 1344
rect 110 1339 111 1343
rect 115 1339 116 1343
rect 110 1338 116 1339
rect 1326 1343 1332 1344
rect 1326 1339 1327 1343
rect 1331 1339 1332 1343
rect 1366 1340 1367 1344
rect 1371 1340 1372 1344
rect 1422 1341 1423 1345
rect 1427 1341 1428 1345
rect 1422 1340 1428 1341
rect 1494 1345 1500 1346
rect 1494 1341 1495 1345
rect 1499 1341 1500 1345
rect 1494 1340 1500 1341
rect 1574 1345 1580 1346
rect 1574 1341 1575 1345
rect 1579 1341 1580 1345
rect 1574 1340 1580 1341
rect 1654 1345 1660 1346
rect 1654 1341 1655 1345
rect 1659 1341 1660 1345
rect 1654 1340 1660 1341
rect 1758 1345 1764 1346
rect 1758 1341 1759 1345
rect 1763 1341 1764 1345
rect 1758 1340 1764 1341
rect 1878 1345 1884 1346
rect 1878 1341 1879 1345
rect 1883 1341 1884 1345
rect 1878 1340 1884 1341
rect 2022 1345 2028 1346
rect 2022 1341 2023 1345
rect 2027 1341 2028 1345
rect 2022 1340 2028 1341
rect 2182 1345 2188 1346
rect 2182 1341 2183 1345
rect 2187 1341 2188 1345
rect 2182 1340 2188 1341
rect 2358 1345 2364 1346
rect 2358 1341 2359 1345
rect 2363 1341 2364 1345
rect 2358 1340 2364 1341
rect 2526 1345 2532 1346
rect 2584 1345 2586 1357
rect 2526 1341 2527 1345
rect 2531 1341 2532 1345
rect 2526 1340 2532 1341
rect 2582 1344 2588 1345
rect 2582 1340 2583 1344
rect 2587 1340 2588 1344
rect 1366 1339 1372 1340
rect 2582 1339 2588 1340
rect 1326 1338 1332 1339
rect 112 1315 114 1338
rect 374 1334 380 1335
rect 374 1330 375 1334
rect 379 1330 380 1334
rect 374 1329 380 1330
rect 430 1334 436 1335
rect 430 1330 431 1334
rect 435 1330 436 1334
rect 430 1329 436 1330
rect 486 1334 492 1335
rect 486 1330 487 1334
rect 491 1330 492 1334
rect 486 1329 492 1330
rect 542 1334 548 1335
rect 542 1330 543 1334
rect 547 1330 548 1334
rect 542 1329 548 1330
rect 606 1334 612 1335
rect 606 1330 607 1334
rect 611 1330 612 1334
rect 606 1329 612 1330
rect 686 1334 692 1335
rect 686 1330 687 1334
rect 691 1330 692 1334
rect 686 1329 692 1330
rect 766 1334 772 1335
rect 766 1330 767 1334
rect 771 1330 772 1334
rect 766 1329 772 1330
rect 854 1334 860 1335
rect 854 1330 855 1334
rect 859 1330 860 1334
rect 854 1329 860 1330
rect 950 1334 956 1335
rect 950 1330 951 1334
rect 955 1330 956 1334
rect 950 1329 956 1330
rect 1046 1334 1052 1335
rect 1046 1330 1047 1334
rect 1051 1330 1052 1334
rect 1046 1329 1052 1330
rect 1142 1334 1148 1335
rect 1142 1330 1143 1334
rect 1147 1330 1148 1334
rect 1142 1329 1148 1330
rect 1246 1334 1252 1335
rect 1246 1330 1247 1334
rect 1251 1330 1252 1334
rect 1246 1329 1252 1330
rect 376 1315 378 1329
rect 432 1315 434 1329
rect 488 1315 490 1329
rect 544 1315 546 1329
rect 608 1315 610 1329
rect 688 1315 690 1329
rect 768 1315 770 1329
rect 856 1315 858 1329
rect 952 1315 954 1329
rect 1048 1315 1050 1329
rect 1144 1315 1146 1329
rect 1248 1315 1250 1329
rect 1328 1315 1330 1338
rect 1366 1327 1372 1328
rect 1366 1323 1367 1327
rect 1371 1323 1372 1327
rect 1366 1322 1372 1323
rect 2582 1327 2588 1328
rect 2582 1323 2583 1327
rect 2587 1323 2588 1327
rect 2582 1322 2588 1323
rect 111 1314 115 1315
rect 111 1309 115 1310
rect 375 1314 379 1315
rect 375 1309 379 1310
rect 431 1314 435 1315
rect 431 1309 435 1310
rect 471 1314 475 1315
rect 471 1309 475 1310
rect 487 1314 491 1315
rect 487 1309 491 1310
rect 527 1314 531 1315
rect 527 1309 531 1310
rect 543 1314 547 1315
rect 543 1309 547 1310
rect 583 1314 587 1315
rect 583 1309 587 1310
rect 607 1314 611 1315
rect 607 1309 611 1310
rect 647 1314 651 1315
rect 647 1309 651 1310
rect 687 1314 691 1315
rect 687 1309 691 1310
rect 727 1314 731 1315
rect 727 1309 731 1310
rect 767 1314 771 1315
rect 767 1309 771 1310
rect 807 1314 811 1315
rect 807 1309 811 1310
rect 855 1314 859 1315
rect 855 1309 859 1310
rect 895 1314 899 1315
rect 895 1309 899 1310
rect 951 1314 955 1315
rect 951 1309 955 1310
rect 991 1314 995 1315
rect 991 1309 995 1310
rect 1047 1314 1051 1315
rect 1047 1309 1051 1310
rect 1095 1314 1099 1315
rect 1095 1309 1099 1310
rect 1143 1314 1147 1315
rect 1143 1309 1147 1310
rect 1199 1314 1203 1315
rect 1199 1309 1203 1310
rect 1247 1314 1251 1315
rect 1247 1309 1251 1310
rect 1287 1314 1291 1315
rect 1287 1309 1291 1310
rect 1327 1314 1331 1315
rect 1327 1309 1331 1310
rect 112 1294 114 1309
rect 472 1303 474 1309
rect 528 1303 530 1309
rect 584 1303 586 1309
rect 648 1303 650 1309
rect 728 1303 730 1309
rect 808 1303 810 1309
rect 896 1303 898 1309
rect 992 1303 994 1309
rect 1096 1303 1098 1309
rect 1200 1303 1202 1309
rect 1288 1303 1290 1309
rect 470 1302 476 1303
rect 470 1298 471 1302
rect 475 1298 476 1302
rect 470 1297 476 1298
rect 526 1302 532 1303
rect 526 1298 527 1302
rect 531 1298 532 1302
rect 526 1297 532 1298
rect 582 1302 588 1303
rect 582 1298 583 1302
rect 587 1298 588 1302
rect 582 1297 588 1298
rect 646 1302 652 1303
rect 646 1298 647 1302
rect 651 1298 652 1302
rect 646 1297 652 1298
rect 726 1302 732 1303
rect 726 1298 727 1302
rect 731 1298 732 1302
rect 726 1297 732 1298
rect 806 1302 812 1303
rect 806 1298 807 1302
rect 811 1298 812 1302
rect 806 1297 812 1298
rect 894 1302 900 1303
rect 894 1298 895 1302
rect 899 1298 900 1302
rect 894 1297 900 1298
rect 990 1302 996 1303
rect 990 1298 991 1302
rect 995 1298 996 1302
rect 990 1297 996 1298
rect 1094 1302 1100 1303
rect 1094 1298 1095 1302
rect 1099 1298 1100 1302
rect 1094 1297 1100 1298
rect 1198 1302 1204 1303
rect 1198 1298 1199 1302
rect 1203 1298 1204 1302
rect 1198 1297 1204 1298
rect 1286 1302 1292 1303
rect 1286 1298 1287 1302
rect 1291 1298 1292 1302
rect 1286 1297 1292 1298
rect 1328 1294 1330 1309
rect 1368 1307 1370 1322
rect 1438 1318 1444 1319
rect 1438 1314 1439 1318
rect 1443 1314 1444 1318
rect 1438 1313 1444 1314
rect 1510 1318 1516 1319
rect 1510 1314 1511 1318
rect 1515 1314 1516 1318
rect 1510 1313 1516 1314
rect 1590 1318 1596 1319
rect 1590 1314 1591 1318
rect 1595 1314 1596 1318
rect 1590 1313 1596 1314
rect 1670 1318 1676 1319
rect 1670 1314 1671 1318
rect 1675 1314 1676 1318
rect 1670 1313 1676 1314
rect 1774 1318 1780 1319
rect 1774 1314 1775 1318
rect 1779 1314 1780 1318
rect 1774 1313 1780 1314
rect 1894 1318 1900 1319
rect 1894 1314 1895 1318
rect 1899 1314 1900 1318
rect 1894 1313 1900 1314
rect 2038 1318 2044 1319
rect 2038 1314 2039 1318
rect 2043 1314 2044 1318
rect 2038 1313 2044 1314
rect 2198 1318 2204 1319
rect 2198 1314 2199 1318
rect 2203 1314 2204 1318
rect 2198 1313 2204 1314
rect 2374 1318 2380 1319
rect 2374 1314 2375 1318
rect 2379 1314 2380 1318
rect 2374 1313 2380 1314
rect 2542 1318 2548 1319
rect 2542 1314 2543 1318
rect 2547 1314 2548 1318
rect 2542 1313 2548 1314
rect 1440 1307 1442 1313
rect 1512 1307 1514 1313
rect 1592 1307 1594 1313
rect 1672 1307 1674 1313
rect 1776 1307 1778 1313
rect 1896 1307 1898 1313
rect 2040 1307 2042 1313
rect 2200 1307 2202 1313
rect 2376 1307 2378 1313
rect 2544 1307 2546 1313
rect 2584 1307 2586 1322
rect 1367 1306 1371 1307
rect 1367 1301 1371 1302
rect 1431 1306 1435 1307
rect 1431 1301 1435 1302
rect 1439 1306 1443 1307
rect 1439 1301 1443 1302
rect 1495 1306 1499 1307
rect 1495 1301 1499 1302
rect 1511 1306 1515 1307
rect 1511 1301 1515 1302
rect 1559 1306 1563 1307
rect 1559 1301 1563 1302
rect 1591 1306 1595 1307
rect 1591 1301 1595 1302
rect 1631 1306 1635 1307
rect 1631 1301 1635 1302
rect 1671 1306 1675 1307
rect 1671 1301 1675 1302
rect 1703 1306 1707 1307
rect 1703 1301 1707 1302
rect 1775 1306 1779 1307
rect 1775 1301 1779 1302
rect 1855 1306 1859 1307
rect 1855 1301 1859 1302
rect 1895 1306 1899 1307
rect 1895 1301 1899 1302
rect 1943 1306 1947 1307
rect 1943 1301 1947 1302
rect 2039 1306 2043 1307
rect 2039 1301 2043 1302
rect 2047 1306 2051 1307
rect 2047 1301 2051 1302
rect 2159 1306 2163 1307
rect 2159 1301 2163 1302
rect 2199 1306 2203 1307
rect 2199 1301 2203 1302
rect 2287 1306 2291 1307
rect 2287 1301 2291 1302
rect 2375 1306 2379 1307
rect 2375 1301 2379 1302
rect 2423 1306 2427 1307
rect 2423 1301 2427 1302
rect 2543 1306 2547 1307
rect 2543 1301 2547 1302
rect 2583 1306 2587 1307
rect 2583 1301 2587 1302
rect 110 1293 116 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 1326 1293 1332 1294
rect 1326 1289 1327 1293
rect 1331 1289 1332 1293
rect 1326 1288 1332 1289
rect 1368 1286 1370 1301
rect 1432 1295 1434 1301
rect 1496 1295 1498 1301
rect 1560 1295 1562 1301
rect 1632 1295 1634 1301
rect 1704 1295 1706 1301
rect 1776 1295 1778 1301
rect 1856 1295 1858 1301
rect 1944 1295 1946 1301
rect 2048 1295 2050 1301
rect 2160 1295 2162 1301
rect 2288 1295 2290 1301
rect 2424 1295 2426 1301
rect 2544 1295 2546 1301
rect 1430 1294 1436 1295
rect 1430 1290 1431 1294
rect 1435 1290 1436 1294
rect 1430 1289 1436 1290
rect 1494 1294 1500 1295
rect 1494 1290 1495 1294
rect 1499 1290 1500 1294
rect 1494 1289 1500 1290
rect 1558 1294 1564 1295
rect 1558 1290 1559 1294
rect 1563 1290 1564 1294
rect 1558 1289 1564 1290
rect 1630 1294 1636 1295
rect 1630 1290 1631 1294
rect 1635 1290 1636 1294
rect 1630 1289 1636 1290
rect 1702 1294 1708 1295
rect 1702 1290 1703 1294
rect 1707 1290 1708 1294
rect 1702 1289 1708 1290
rect 1774 1294 1780 1295
rect 1774 1290 1775 1294
rect 1779 1290 1780 1294
rect 1774 1289 1780 1290
rect 1854 1294 1860 1295
rect 1854 1290 1855 1294
rect 1859 1290 1860 1294
rect 1854 1289 1860 1290
rect 1942 1294 1948 1295
rect 1942 1290 1943 1294
rect 1947 1290 1948 1294
rect 1942 1289 1948 1290
rect 2046 1294 2052 1295
rect 2046 1290 2047 1294
rect 2051 1290 2052 1294
rect 2046 1289 2052 1290
rect 2158 1294 2164 1295
rect 2158 1290 2159 1294
rect 2163 1290 2164 1294
rect 2158 1289 2164 1290
rect 2286 1294 2292 1295
rect 2286 1290 2287 1294
rect 2291 1290 2292 1294
rect 2286 1289 2292 1290
rect 2422 1294 2428 1295
rect 2422 1290 2423 1294
rect 2427 1290 2428 1294
rect 2422 1289 2428 1290
rect 2542 1294 2548 1295
rect 2542 1290 2543 1294
rect 2547 1290 2548 1294
rect 2542 1289 2548 1290
rect 2584 1286 2586 1301
rect 1366 1285 1372 1286
rect 1366 1281 1367 1285
rect 1371 1281 1372 1285
rect 1366 1280 1372 1281
rect 2582 1285 2588 1286
rect 2582 1281 2583 1285
rect 2587 1281 2588 1285
rect 2582 1280 2588 1281
rect 110 1276 116 1277
rect 1326 1276 1332 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 110 1271 116 1272
rect 454 1275 460 1276
rect 454 1271 455 1275
rect 459 1271 460 1275
rect 112 1255 114 1271
rect 454 1270 460 1271
rect 510 1275 516 1276
rect 510 1271 511 1275
rect 515 1271 516 1275
rect 510 1270 516 1271
rect 566 1275 572 1276
rect 566 1271 567 1275
rect 571 1271 572 1275
rect 566 1270 572 1271
rect 630 1275 636 1276
rect 630 1271 631 1275
rect 635 1271 636 1275
rect 630 1270 636 1271
rect 710 1275 716 1276
rect 710 1271 711 1275
rect 715 1271 716 1275
rect 710 1270 716 1271
rect 790 1275 796 1276
rect 790 1271 791 1275
rect 795 1271 796 1275
rect 790 1270 796 1271
rect 878 1275 884 1276
rect 878 1271 879 1275
rect 883 1271 884 1275
rect 878 1270 884 1271
rect 974 1275 980 1276
rect 974 1271 975 1275
rect 979 1271 980 1275
rect 974 1270 980 1271
rect 1078 1275 1084 1276
rect 1078 1271 1079 1275
rect 1083 1271 1084 1275
rect 1078 1270 1084 1271
rect 1182 1275 1188 1276
rect 1182 1271 1183 1275
rect 1187 1271 1188 1275
rect 1182 1270 1188 1271
rect 1270 1275 1276 1276
rect 1270 1271 1271 1275
rect 1275 1271 1276 1275
rect 1326 1272 1327 1276
rect 1331 1272 1332 1276
rect 1326 1271 1332 1272
rect 1270 1270 1276 1271
rect 456 1255 458 1270
rect 512 1255 514 1270
rect 568 1255 570 1270
rect 632 1255 634 1270
rect 712 1255 714 1270
rect 792 1255 794 1270
rect 880 1255 882 1270
rect 976 1255 978 1270
rect 1080 1255 1082 1270
rect 1184 1255 1186 1270
rect 1272 1255 1274 1270
rect 1328 1255 1330 1271
rect 1366 1268 1372 1269
rect 2582 1268 2588 1269
rect 1366 1264 1367 1268
rect 1371 1264 1372 1268
rect 1366 1263 1372 1264
rect 1414 1267 1420 1268
rect 1414 1263 1415 1267
rect 1419 1263 1420 1267
rect 111 1254 115 1255
rect 111 1249 115 1250
rect 383 1254 387 1255
rect 383 1249 387 1250
rect 439 1254 443 1255
rect 439 1249 443 1250
rect 455 1254 459 1255
rect 455 1249 459 1250
rect 503 1254 507 1255
rect 503 1249 507 1250
rect 511 1254 515 1255
rect 511 1249 515 1250
rect 567 1254 571 1255
rect 567 1249 571 1250
rect 575 1254 579 1255
rect 575 1249 579 1250
rect 631 1254 635 1255
rect 631 1249 635 1250
rect 647 1254 651 1255
rect 647 1249 651 1250
rect 711 1254 715 1255
rect 711 1249 715 1250
rect 727 1254 731 1255
rect 727 1249 731 1250
rect 791 1254 795 1255
rect 791 1249 795 1250
rect 815 1254 819 1255
rect 815 1249 819 1250
rect 879 1254 883 1255
rect 879 1249 883 1250
rect 903 1254 907 1255
rect 903 1249 907 1250
rect 975 1254 979 1255
rect 975 1249 979 1250
rect 991 1254 995 1255
rect 991 1249 995 1250
rect 1079 1254 1083 1255
rect 1079 1249 1083 1250
rect 1175 1254 1179 1255
rect 1175 1249 1179 1250
rect 1183 1254 1187 1255
rect 1183 1249 1187 1250
rect 1271 1254 1275 1255
rect 1271 1249 1275 1250
rect 1327 1254 1331 1255
rect 1327 1249 1331 1250
rect 112 1237 114 1249
rect 384 1238 386 1249
rect 440 1238 442 1249
rect 504 1238 506 1249
rect 576 1238 578 1249
rect 648 1238 650 1249
rect 728 1238 730 1249
rect 816 1238 818 1249
rect 904 1238 906 1249
rect 992 1238 994 1249
rect 1080 1238 1082 1249
rect 1176 1238 1178 1249
rect 1272 1238 1274 1249
rect 382 1237 388 1238
rect 110 1236 116 1237
rect 110 1232 111 1236
rect 115 1232 116 1236
rect 382 1233 383 1237
rect 387 1233 388 1237
rect 382 1232 388 1233
rect 438 1237 444 1238
rect 438 1233 439 1237
rect 443 1233 444 1237
rect 438 1232 444 1233
rect 502 1237 508 1238
rect 502 1233 503 1237
rect 507 1233 508 1237
rect 502 1232 508 1233
rect 574 1237 580 1238
rect 574 1233 575 1237
rect 579 1233 580 1237
rect 574 1232 580 1233
rect 646 1237 652 1238
rect 646 1233 647 1237
rect 651 1233 652 1237
rect 646 1232 652 1233
rect 726 1237 732 1238
rect 726 1233 727 1237
rect 731 1233 732 1237
rect 726 1232 732 1233
rect 814 1237 820 1238
rect 814 1233 815 1237
rect 819 1233 820 1237
rect 814 1232 820 1233
rect 902 1237 908 1238
rect 902 1233 903 1237
rect 907 1233 908 1237
rect 902 1232 908 1233
rect 990 1237 996 1238
rect 990 1233 991 1237
rect 995 1233 996 1237
rect 990 1232 996 1233
rect 1078 1237 1084 1238
rect 1078 1233 1079 1237
rect 1083 1233 1084 1237
rect 1078 1232 1084 1233
rect 1174 1237 1180 1238
rect 1174 1233 1175 1237
rect 1179 1233 1180 1237
rect 1174 1232 1180 1233
rect 1270 1237 1276 1238
rect 1328 1237 1330 1249
rect 1368 1247 1370 1263
rect 1414 1262 1420 1263
rect 1478 1267 1484 1268
rect 1478 1263 1479 1267
rect 1483 1263 1484 1267
rect 1478 1262 1484 1263
rect 1542 1267 1548 1268
rect 1542 1263 1543 1267
rect 1547 1263 1548 1267
rect 1542 1262 1548 1263
rect 1614 1267 1620 1268
rect 1614 1263 1615 1267
rect 1619 1263 1620 1267
rect 1614 1262 1620 1263
rect 1686 1267 1692 1268
rect 1686 1263 1687 1267
rect 1691 1263 1692 1267
rect 1686 1262 1692 1263
rect 1758 1267 1764 1268
rect 1758 1263 1759 1267
rect 1763 1263 1764 1267
rect 1758 1262 1764 1263
rect 1838 1267 1844 1268
rect 1838 1263 1839 1267
rect 1843 1263 1844 1267
rect 1838 1262 1844 1263
rect 1926 1267 1932 1268
rect 1926 1263 1927 1267
rect 1931 1263 1932 1267
rect 1926 1262 1932 1263
rect 2030 1267 2036 1268
rect 2030 1263 2031 1267
rect 2035 1263 2036 1267
rect 2030 1262 2036 1263
rect 2142 1267 2148 1268
rect 2142 1263 2143 1267
rect 2147 1263 2148 1267
rect 2142 1262 2148 1263
rect 2270 1267 2276 1268
rect 2270 1263 2271 1267
rect 2275 1263 2276 1267
rect 2270 1262 2276 1263
rect 2406 1267 2412 1268
rect 2406 1263 2407 1267
rect 2411 1263 2412 1267
rect 2406 1262 2412 1263
rect 2526 1267 2532 1268
rect 2526 1263 2527 1267
rect 2531 1263 2532 1267
rect 2582 1264 2583 1268
rect 2587 1264 2588 1268
rect 2582 1263 2588 1264
rect 2526 1262 2532 1263
rect 1416 1247 1418 1262
rect 1480 1247 1482 1262
rect 1544 1247 1546 1262
rect 1616 1247 1618 1262
rect 1688 1247 1690 1262
rect 1760 1247 1762 1262
rect 1840 1247 1842 1262
rect 1928 1247 1930 1262
rect 2032 1247 2034 1262
rect 2144 1247 2146 1262
rect 2272 1247 2274 1262
rect 2408 1247 2410 1262
rect 2528 1247 2530 1262
rect 2584 1247 2586 1263
rect 1367 1246 1371 1247
rect 1367 1241 1371 1242
rect 1399 1246 1403 1247
rect 1399 1241 1403 1242
rect 1415 1246 1419 1247
rect 1415 1241 1419 1242
rect 1455 1246 1459 1247
rect 1455 1241 1459 1242
rect 1479 1246 1483 1247
rect 1479 1241 1483 1242
rect 1535 1246 1539 1247
rect 1535 1241 1539 1242
rect 1543 1246 1547 1247
rect 1543 1241 1547 1242
rect 1615 1246 1619 1247
rect 1615 1241 1619 1242
rect 1687 1246 1691 1247
rect 1687 1241 1691 1242
rect 1695 1246 1699 1247
rect 1695 1241 1699 1242
rect 1759 1246 1763 1247
rect 1759 1241 1763 1242
rect 1775 1246 1779 1247
rect 1775 1241 1779 1242
rect 1839 1246 1843 1247
rect 1839 1241 1843 1242
rect 1855 1246 1859 1247
rect 1855 1241 1859 1242
rect 1927 1246 1931 1247
rect 1927 1241 1931 1242
rect 1943 1246 1947 1247
rect 1943 1241 1947 1242
rect 2031 1246 2035 1247
rect 2031 1241 2035 1242
rect 2039 1246 2043 1247
rect 2039 1241 2043 1242
rect 2143 1246 2147 1247
rect 2143 1241 2147 1242
rect 2151 1246 2155 1247
rect 2151 1241 2155 1242
rect 2271 1246 2275 1247
rect 2271 1241 2275 1242
rect 2279 1246 2283 1247
rect 2279 1241 2283 1242
rect 2407 1246 2411 1247
rect 2407 1241 2411 1242
rect 2415 1246 2419 1247
rect 2415 1241 2419 1242
rect 2527 1246 2531 1247
rect 2527 1241 2531 1242
rect 2583 1246 2587 1247
rect 2583 1241 2587 1242
rect 1270 1233 1271 1237
rect 1275 1233 1276 1237
rect 1270 1232 1276 1233
rect 1326 1236 1332 1237
rect 1326 1232 1327 1236
rect 1331 1232 1332 1236
rect 110 1231 116 1232
rect 1326 1231 1332 1232
rect 1368 1229 1370 1241
rect 1400 1230 1402 1241
rect 1456 1230 1458 1241
rect 1536 1230 1538 1241
rect 1616 1230 1618 1241
rect 1696 1230 1698 1241
rect 1776 1230 1778 1241
rect 1856 1230 1858 1241
rect 1944 1230 1946 1241
rect 2040 1230 2042 1241
rect 2152 1230 2154 1241
rect 2280 1230 2282 1241
rect 2416 1230 2418 1241
rect 2528 1230 2530 1241
rect 1398 1229 1404 1230
rect 1366 1228 1372 1229
rect 1366 1224 1367 1228
rect 1371 1224 1372 1228
rect 1398 1225 1399 1229
rect 1403 1225 1404 1229
rect 1398 1224 1404 1225
rect 1454 1229 1460 1230
rect 1454 1225 1455 1229
rect 1459 1225 1460 1229
rect 1454 1224 1460 1225
rect 1534 1229 1540 1230
rect 1534 1225 1535 1229
rect 1539 1225 1540 1229
rect 1534 1224 1540 1225
rect 1614 1229 1620 1230
rect 1614 1225 1615 1229
rect 1619 1225 1620 1229
rect 1614 1224 1620 1225
rect 1694 1229 1700 1230
rect 1694 1225 1695 1229
rect 1699 1225 1700 1229
rect 1694 1224 1700 1225
rect 1774 1229 1780 1230
rect 1774 1225 1775 1229
rect 1779 1225 1780 1229
rect 1774 1224 1780 1225
rect 1854 1229 1860 1230
rect 1854 1225 1855 1229
rect 1859 1225 1860 1229
rect 1854 1224 1860 1225
rect 1942 1229 1948 1230
rect 1942 1225 1943 1229
rect 1947 1225 1948 1229
rect 1942 1224 1948 1225
rect 2038 1229 2044 1230
rect 2038 1225 2039 1229
rect 2043 1225 2044 1229
rect 2038 1224 2044 1225
rect 2150 1229 2156 1230
rect 2150 1225 2151 1229
rect 2155 1225 2156 1229
rect 2150 1224 2156 1225
rect 2278 1229 2284 1230
rect 2278 1225 2279 1229
rect 2283 1225 2284 1229
rect 2278 1224 2284 1225
rect 2414 1229 2420 1230
rect 2414 1225 2415 1229
rect 2419 1225 2420 1229
rect 2414 1224 2420 1225
rect 2526 1229 2532 1230
rect 2584 1229 2586 1241
rect 2526 1225 2527 1229
rect 2531 1225 2532 1229
rect 2526 1224 2532 1225
rect 2582 1228 2588 1229
rect 2582 1224 2583 1228
rect 2587 1224 2588 1228
rect 1366 1223 1372 1224
rect 2582 1223 2588 1224
rect 110 1219 116 1220
rect 110 1215 111 1219
rect 115 1215 116 1219
rect 110 1214 116 1215
rect 1326 1219 1332 1220
rect 1326 1215 1327 1219
rect 1331 1215 1332 1219
rect 1326 1214 1332 1215
rect 112 1195 114 1214
rect 398 1210 404 1211
rect 398 1206 399 1210
rect 403 1206 404 1210
rect 398 1205 404 1206
rect 454 1210 460 1211
rect 454 1206 455 1210
rect 459 1206 460 1210
rect 454 1205 460 1206
rect 518 1210 524 1211
rect 518 1206 519 1210
rect 523 1206 524 1210
rect 518 1205 524 1206
rect 590 1210 596 1211
rect 590 1206 591 1210
rect 595 1206 596 1210
rect 590 1205 596 1206
rect 662 1210 668 1211
rect 662 1206 663 1210
rect 667 1206 668 1210
rect 662 1205 668 1206
rect 742 1210 748 1211
rect 742 1206 743 1210
rect 747 1206 748 1210
rect 742 1205 748 1206
rect 830 1210 836 1211
rect 830 1206 831 1210
rect 835 1206 836 1210
rect 830 1205 836 1206
rect 918 1210 924 1211
rect 918 1206 919 1210
rect 923 1206 924 1210
rect 918 1205 924 1206
rect 1006 1210 1012 1211
rect 1006 1206 1007 1210
rect 1011 1206 1012 1210
rect 1006 1205 1012 1206
rect 1094 1210 1100 1211
rect 1094 1206 1095 1210
rect 1099 1206 1100 1210
rect 1094 1205 1100 1206
rect 1190 1210 1196 1211
rect 1190 1206 1191 1210
rect 1195 1206 1196 1210
rect 1190 1205 1196 1206
rect 1286 1210 1292 1211
rect 1286 1206 1287 1210
rect 1291 1206 1292 1210
rect 1286 1205 1292 1206
rect 400 1195 402 1205
rect 456 1195 458 1205
rect 520 1195 522 1205
rect 592 1195 594 1205
rect 664 1195 666 1205
rect 744 1195 746 1205
rect 832 1195 834 1205
rect 920 1195 922 1205
rect 1008 1195 1010 1205
rect 1096 1195 1098 1205
rect 1192 1195 1194 1205
rect 1288 1195 1290 1205
rect 1328 1195 1330 1214
rect 1366 1211 1372 1212
rect 1366 1207 1367 1211
rect 1371 1207 1372 1211
rect 1366 1206 1372 1207
rect 2582 1211 2588 1212
rect 2582 1207 2583 1211
rect 2587 1207 2588 1211
rect 2582 1206 2588 1207
rect 111 1194 115 1195
rect 111 1189 115 1190
rect 279 1194 283 1195
rect 279 1189 283 1190
rect 343 1194 347 1195
rect 343 1189 347 1190
rect 399 1194 403 1195
rect 399 1189 403 1190
rect 415 1194 419 1195
rect 415 1189 419 1190
rect 455 1194 459 1195
rect 455 1189 459 1190
rect 495 1194 499 1195
rect 495 1189 499 1190
rect 519 1194 523 1195
rect 519 1189 523 1190
rect 583 1194 587 1195
rect 583 1189 587 1190
rect 591 1194 595 1195
rect 591 1189 595 1190
rect 663 1194 667 1195
rect 663 1189 667 1190
rect 671 1194 675 1195
rect 671 1189 675 1190
rect 743 1194 747 1195
rect 743 1189 747 1190
rect 759 1194 763 1195
rect 759 1189 763 1190
rect 831 1194 835 1195
rect 831 1189 835 1190
rect 847 1194 851 1195
rect 847 1189 851 1190
rect 919 1194 923 1195
rect 919 1189 923 1190
rect 935 1194 939 1195
rect 935 1189 939 1190
rect 1007 1194 1011 1195
rect 1007 1189 1011 1190
rect 1015 1194 1019 1195
rect 1015 1189 1019 1190
rect 1087 1194 1091 1195
rect 1087 1189 1091 1190
rect 1095 1194 1099 1195
rect 1095 1189 1099 1190
rect 1159 1194 1163 1195
rect 1159 1189 1163 1190
rect 1191 1194 1195 1195
rect 1191 1189 1195 1190
rect 1231 1194 1235 1195
rect 1231 1189 1235 1190
rect 1287 1194 1291 1195
rect 1287 1189 1291 1190
rect 1327 1194 1331 1195
rect 1327 1189 1331 1190
rect 112 1174 114 1189
rect 280 1183 282 1189
rect 344 1183 346 1189
rect 416 1183 418 1189
rect 496 1183 498 1189
rect 584 1183 586 1189
rect 672 1183 674 1189
rect 760 1183 762 1189
rect 848 1183 850 1189
rect 936 1183 938 1189
rect 1016 1183 1018 1189
rect 1088 1183 1090 1189
rect 1160 1183 1162 1189
rect 1232 1183 1234 1189
rect 1288 1183 1290 1189
rect 278 1182 284 1183
rect 278 1178 279 1182
rect 283 1178 284 1182
rect 278 1177 284 1178
rect 342 1182 348 1183
rect 342 1178 343 1182
rect 347 1178 348 1182
rect 342 1177 348 1178
rect 414 1182 420 1183
rect 414 1178 415 1182
rect 419 1178 420 1182
rect 414 1177 420 1178
rect 494 1182 500 1183
rect 494 1178 495 1182
rect 499 1178 500 1182
rect 494 1177 500 1178
rect 582 1182 588 1183
rect 582 1178 583 1182
rect 587 1178 588 1182
rect 582 1177 588 1178
rect 670 1182 676 1183
rect 670 1178 671 1182
rect 675 1178 676 1182
rect 670 1177 676 1178
rect 758 1182 764 1183
rect 758 1178 759 1182
rect 763 1178 764 1182
rect 758 1177 764 1178
rect 846 1182 852 1183
rect 846 1178 847 1182
rect 851 1178 852 1182
rect 846 1177 852 1178
rect 934 1182 940 1183
rect 934 1178 935 1182
rect 939 1178 940 1182
rect 934 1177 940 1178
rect 1014 1182 1020 1183
rect 1014 1178 1015 1182
rect 1019 1178 1020 1182
rect 1014 1177 1020 1178
rect 1086 1182 1092 1183
rect 1086 1178 1087 1182
rect 1091 1178 1092 1182
rect 1086 1177 1092 1178
rect 1158 1182 1164 1183
rect 1158 1178 1159 1182
rect 1163 1178 1164 1182
rect 1158 1177 1164 1178
rect 1230 1182 1236 1183
rect 1230 1178 1231 1182
rect 1235 1178 1236 1182
rect 1230 1177 1236 1178
rect 1286 1182 1292 1183
rect 1286 1178 1287 1182
rect 1291 1178 1292 1182
rect 1286 1177 1292 1178
rect 1328 1174 1330 1189
rect 1368 1183 1370 1206
rect 1414 1202 1420 1203
rect 1414 1198 1415 1202
rect 1419 1198 1420 1202
rect 1414 1197 1420 1198
rect 1470 1202 1476 1203
rect 1470 1198 1471 1202
rect 1475 1198 1476 1202
rect 1470 1197 1476 1198
rect 1550 1202 1556 1203
rect 1550 1198 1551 1202
rect 1555 1198 1556 1202
rect 1550 1197 1556 1198
rect 1630 1202 1636 1203
rect 1630 1198 1631 1202
rect 1635 1198 1636 1202
rect 1630 1197 1636 1198
rect 1710 1202 1716 1203
rect 1710 1198 1711 1202
rect 1715 1198 1716 1202
rect 1710 1197 1716 1198
rect 1790 1202 1796 1203
rect 1790 1198 1791 1202
rect 1795 1198 1796 1202
rect 1790 1197 1796 1198
rect 1870 1202 1876 1203
rect 1870 1198 1871 1202
rect 1875 1198 1876 1202
rect 1870 1197 1876 1198
rect 1958 1202 1964 1203
rect 1958 1198 1959 1202
rect 1963 1198 1964 1202
rect 1958 1197 1964 1198
rect 2054 1202 2060 1203
rect 2054 1198 2055 1202
rect 2059 1198 2060 1202
rect 2054 1197 2060 1198
rect 2166 1202 2172 1203
rect 2166 1198 2167 1202
rect 2171 1198 2172 1202
rect 2166 1197 2172 1198
rect 2294 1202 2300 1203
rect 2294 1198 2295 1202
rect 2299 1198 2300 1202
rect 2294 1197 2300 1198
rect 2430 1202 2436 1203
rect 2430 1198 2431 1202
rect 2435 1198 2436 1202
rect 2430 1197 2436 1198
rect 2542 1202 2548 1203
rect 2542 1198 2543 1202
rect 2547 1198 2548 1202
rect 2542 1197 2548 1198
rect 1416 1183 1418 1197
rect 1472 1183 1474 1197
rect 1552 1183 1554 1197
rect 1632 1183 1634 1197
rect 1712 1183 1714 1197
rect 1792 1183 1794 1197
rect 1872 1183 1874 1197
rect 1960 1183 1962 1197
rect 2056 1183 2058 1197
rect 2168 1183 2170 1197
rect 2296 1183 2298 1197
rect 2432 1183 2434 1197
rect 2544 1183 2546 1197
rect 2584 1183 2586 1206
rect 1367 1182 1371 1183
rect 1367 1177 1371 1178
rect 1415 1182 1419 1183
rect 1415 1177 1419 1178
rect 1471 1182 1475 1183
rect 1471 1177 1475 1178
rect 1551 1182 1555 1183
rect 1551 1177 1555 1178
rect 1631 1182 1635 1183
rect 1631 1177 1635 1178
rect 1695 1182 1699 1183
rect 1695 1177 1699 1178
rect 1711 1182 1715 1183
rect 1711 1177 1715 1178
rect 1767 1182 1771 1183
rect 1767 1177 1771 1178
rect 1791 1182 1795 1183
rect 1791 1177 1795 1178
rect 1847 1182 1851 1183
rect 1847 1177 1851 1178
rect 1871 1182 1875 1183
rect 1871 1177 1875 1178
rect 1919 1182 1923 1183
rect 1919 1177 1923 1178
rect 1959 1182 1963 1183
rect 1959 1177 1963 1178
rect 1991 1182 1995 1183
rect 1991 1177 1995 1178
rect 2055 1182 2059 1183
rect 2055 1177 2059 1178
rect 2063 1182 2067 1183
rect 2063 1177 2067 1178
rect 2135 1182 2139 1183
rect 2135 1177 2139 1178
rect 2167 1182 2171 1183
rect 2167 1177 2171 1178
rect 2207 1182 2211 1183
rect 2207 1177 2211 1178
rect 2287 1182 2291 1183
rect 2287 1177 2291 1178
rect 2295 1182 2299 1183
rect 2295 1177 2299 1178
rect 2367 1182 2371 1183
rect 2367 1177 2371 1178
rect 2431 1182 2435 1183
rect 2431 1177 2435 1178
rect 2543 1182 2547 1183
rect 2543 1177 2547 1178
rect 2583 1182 2587 1183
rect 2583 1177 2587 1178
rect 110 1173 116 1174
rect 110 1169 111 1173
rect 115 1169 116 1173
rect 110 1168 116 1169
rect 1326 1173 1332 1174
rect 1326 1169 1327 1173
rect 1331 1169 1332 1173
rect 1326 1168 1332 1169
rect 1368 1162 1370 1177
rect 1696 1171 1698 1177
rect 1768 1171 1770 1177
rect 1848 1171 1850 1177
rect 1920 1171 1922 1177
rect 1992 1171 1994 1177
rect 2064 1171 2066 1177
rect 2136 1171 2138 1177
rect 2208 1171 2210 1177
rect 2288 1171 2290 1177
rect 2368 1171 2370 1177
rect 1694 1170 1700 1171
rect 1694 1166 1695 1170
rect 1699 1166 1700 1170
rect 1694 1165 1700 1166
rect 1766 1170 1772 1171
rect 1766 1166 1767 1170
rect 1771 1166 1772 1170
rect 1766 1165 1772 1166
rect 1846 1170 1852 1171
rect 1846 1166 1847 1170
rect 1851 1166 1852 1170
rect 1846 1165 1852 1166
rect 1918 1170 1924 1171
rect 1918 1166 1919 1170
rect 1923 1166 1924 1170
rect 1918 1165 1924 1166
rect 1990 1170 1996 1171
rect 1990 1166 1991 1170
rect 1995 1166 1996 1170
rect 1990 1165 1996 1166
rect 2062 1170 2068 1171
rect 2062 1166 2063 1170
rect 2067 1166 2068 1170
rect 2062 1165 2068 1166
rect 2134 1170 2140 1171
rect 2134 1166 2135 1170
rect 2139 1166 2140 1170
rect 2134 1165 2140 1166
rect 2206 1170 2212 1171
rect 2206 1166 2207 1170
rect 2211 1166 2212 1170
rect 2206 1165 2212 1166
rect 2286 1170 2292 1171
rect 2286 1166 2287 1170
rect 2291 1166 2292 1170
rect 2286 1165 2292 1166
rect 2366 1170 2372 1171
rect 2366 1166 2367 1170
rect 2371 1166 2372 1170
rect 2366 1165 2372 1166
rect 2584 1162 2586 1177
rect 1366 1161 1372 1162
rect 1366 1157 1367 1161
rect 1371 1157 1372 1161
rect 110 1156 116 1157
rect 1326 1156 1332 1157
rect 1366 1156 1372 1157
rect 2582 1161 2588 1162
rect 2582 1157 2583 1161
rect 2587 1157 2588 1161
rect 2582 1156 2588 1157
rect 110 1152 111 1156
rect 115 1152 116 1156
rect 110 1151 116 1152
rect 262 1155 268 1156
rect 262 1151 263 1155
rect 267 1151 268 1155
rect 112 1131 114 1151
rect 262 1150 268 1151
rect 326 1155 332 1156
rect 326 1151 327 1155
rect 331 1151 332 1155
rect 326 1150 332 1151
rect 398 1155 404 1156
rect 398 1151 399 1155
rect 403 1151 404 1155
rect 398 1150 404 1151
rect 478 1155 484 1156
rect 478 1151 479 1155
rect 483 1151 484 1155
rect 478 1150 484 1151
rect 566 1155 572 1156
rect 566 1151 567 1155
rect 571 1151 572 1155
rect 566 1150 572 1151
rect 654 1155 660 1156
rect 654 1151 655 1155
rect 659 1151 660 1155
rect 654 1150 660 1151
rect 742 1155 748 1156
rect 742 1151 743 1155
rect 747 1151 748 1155
rect 742 1150 748 1151
rect 830 1155 836 1156
rect 830 1151 831 1155
rect 835 1151 836 1155
rect 830 1150 836 1151
rect 918 1155 924 1156
rect 918 1151 919 1155
rect 923 1151 924 1155
rect 918 1150 924 1151
rect 998 1155 1004 1156
rect 998 1151 999 1155
rect 1003 1151 1004 1155
rect 998 1150 1004 1151
rect 1070 1155 1076 1156
rect 1070 1151 1071 1155
rect 1075 1151 1076 1155
rect 1070 1150 1076 1151
rect 1142 1155 1148 1156
rect 1142 1151 1143 1155
rect 1147 1151 1148 1155
rect 1142 1150 1148 1151
rect 1214 1155 1220 1156
rect 1214 1151 1215 1155
rect 1219 1151 1220 1155
rect 1214 1150 1220 1151
rect 1270 1155 1276 1156
rect 1270 1151 1271 1155
rect 1275 1151 1276 1155
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1326 1151 1332 1152
rect 1270 1150 1276 1151
rect 264 1131 266 1150
rect 328 1131 330 1150
rect 400 1131 402 1150
rect 480 1131 482 1150
rect 568 1131 570 1150
rect 656 1131 658 1150
rect 744 1131 746 1150
rect 832 1131 834 1150
rect 920 1131 922 1150
rect 1000 1131 1002 1150
rect 1072 1131 1074 1150
rect 1144 1131 1146 1150
rect 1216 1131 1218 1150
rect 1272 1131 1274 1150
rect 1328 1131 1330 1151
rect 1366 1144 1372 1145
rect 2582 1144 2588 1145
rect 1366 1140 1367 1144
rect 1371 1140 1372 1144
rect 1366 1139 1372 1140
rect 1678 1143 1684 1144
rect 1678 1139 1679 1143
rect 1683 1139 1684 1143
rect 111 1130 115 1131
rect 111 1125 115 1126
rect 143 1130 147 1131
rect 143 1125 147 1126
rect 207 1130 211 1131
rect 207 1125 211 1126
rect 263 1130 267 1131
rect 263 1125 267 1126
rect 271 1130 275 1131
rect 271 1125 275 1126
rect 327 1130 331 1131
rect 327 1125 331 1126
rect 343 1130 347 1131
rect 343 1125 347 1126
rect 399 1130 403 1131
rect 399 1125 403 1126
rect 423 1130 427 1131
rect 423 1125 427 1126
rect 479 1130 483 1131
rect 479 1125 483 1126
rect 503 1130 507 1131
rect 503 1125 507 1126
rect 567 1130 571 1131
rect 567 1125 571 1126
rect 583 1130 587 1131
rect 583 1125 587 1126
rect 655 1130 659 1131
rect 655 1125 659 1126
rect 663 1130 667 1131
rect 663 1125 667 1126
rect 743 1130 747 1131
rect 743 1125 747 1126
rect 831 1130 835 1131
rect 831 1125 835 1126
rect 919 1130 923 1131
rect 919 1125 923 1126
rect 999 1130 1003 1131
rect 999 1125 1003 1126
rect 1007 1130 1011 1131
rect 1007 1125 1011 1126
rect 1071 1130 1075 1131
rect 1071 1125 1075 1126
rect 1143 1130 1147 1131
rect 1143 1125 1147 1126
rect 1215 1130 1219 1131
rect 1215 1125 1219 1126
rect 1271 1130 1275 1131
rect 1271 1125 1275 1126
rect 1327 1130 1331 1131
rect 1368 1127 1370 1139
rect 1678 1138 1684 1139
rect 1750 1143 1756 1144
rect 1750 1139 1751 1143
rect 1755 1139 1756 1143
rect 1750 1138 1756 1139
rect 1830 1143 1836 1144
rect 1830 1139 1831 1143
rect 1835 1139 1836 1143
rect 1830 1138 1836 1139
rect 1902 1143 1908 1144
rect 1902 1139 1903 1143
rect 1907 1139 1908 1143
rect 1902 1138 1908 1139
rect 1974 1143 1980 1144
rect 1974 1139 1975 1143
rect 1979 1139 1980 1143
rect 1974 1138 1980 1139
rect 2046 1143 2052 1144
rect 2046 1139 2047 1143
rect 2051 1139 2052 1143
rect 2046 1138 2052 1139
rect 2118 1143 2124 1144
rect 2118 1139 2119 1143
rect 2123 1139 2124 1143
rect 2118 1138 2124 1139
rect 2190 1143 2196 1144
rect 2190 1139 2191 1143
rect 2195 1139 2196 1143
rect 2190 1138 2196 1139
rect 2270 1143 2276 1144
rect 2270 1139 2271 1143
rect 2275 1139 2276 1143
rect 2270 1138 2276 1139
rect 2350 1143 2356 1144
rect 2350 1139 2351 1143
rect 2355 1139 2356 1143
rect 2582 1140 2583 1144
rect 2587 1140 2588 1144
rect 2582 1139 2588 1140
rect 2350 1138 2356 1139
rect 1680 1127 1682 1138
rect 1752 1127 1754 1138
rect 1832 1127 1834 1138
rect 1904 1127 1906 1138
rect 1976 1127 1978 1138
rect 2048 1127 2050 1138
rect 2120 1127 2122 1138
rect 2192 1127 2194 1138
rect 2272 1127 2274 1138
rect 2352 1127 2354 1138
rect 2584 1127 2586 1139
rect 1327 1125 1331 1126
rect 1367 1126 1371 1127
rect 112 1113 114 1125
rect 144 1114 146 1125
rect 208 1114 210 1125
rect 272 1114 274 1125
rect 344 1114 346 1125
rect 424 1114 426 1125
rect 504 1114 506 1125
rect 584 1114 586 1125
rect 664 1114 666 1125
rect 744 1114 746 1125
rect 832 1114 834 1125
rect 920 1114 922 1125
rect 1008 1114 1010 1125
rect 142 1113 148 1114
rect 110 1112 116 1113
rect 110 1108 111 1112
rect 115 1108 116 1112
rect 142 1109 143 1113
rect 147 1109 148 1113
rect 142 1108 148 1109
rect 206 1113 212 1114
rect 206 1109 207 1113
rect 211 1109 212 1113
rect 206 1108 212 1109
rect 270 1113 276 1114
rect 270 1109 271 1113
rect 275 1109 276 1113
rect 270 1108 276 1109
rect 342 1113 348 1114
rect 342 1109 343 1113
rect 347 1109 348 1113
rect 342 1108 348 1109
rect 422 1113 428 1114
rect 422 1109 423 1113
rect 427 1109 428 1113
rect 422 1108 428 1109
rect 502 1113 508 1114
rect 502 1109 503 1113
rect 507 1109 508 1113
rect 502 1108 508 1109
rect 582 1113 588 1114
rect 582 1109 583 1113
rect 587 1109 588 1113
rect 582 1108 588 1109
rect 662 1113 668 1114
rect 662 1109 663 1113
rect 667 1109 668 1113
rect 662 1108 668 1109
rect 742 1113 748 1114
rect 742 1109 743 1113
rect 747 1109 748 1113
rect 742 1108 748 1109
rect 830 1113 836 1114
rect 830 1109 831 1113
rect 835 1109 836 1113
rect 830 1108 836 1109
rect 918 1113 924 1114
rect 918 1109 919 1113
rect 923 1109 924 1113
rect 918 1108 924 1109
rect 1006 1113 1012 1114
rect 1328 1113 1330 1125
rect 1367 1121 1371 1122
rect 1399 1126 1403 1127
rect 1399 1121 1403 1122
rect 1479 1126 1483 1127
rect 1479 1121 1483 1122
rect 1583 1126 1587 1127
rect 1583 1121 1587 1122
rect 1679 1126 1683 1127
rect 1679 1121 1683 1122
rect 1687 1126 1691 1127
rect 1687 1121 1691 1122
rect 1751 1126 1755 1127
rect 1751 1121 1755 1122
rect 1783 1126 1787 1127
rect 1783 1121 1787 1122
rect 1831 1126 1835 1127
rect 1831 1121 1835 1122
rect 1879 1126 1883 1127
rect 1879 1121 1883 1122
rect 1903 1126 1907 1127
rect 1903 1121 1907 1122
rect 1975 1126 1979 1127
rect 1975 1121 1979 1122
rect 2047 1126 2051 1127
rect 2047 1121 2051 1122
rect 2063 1126 2067 1127
rect 2063 1121 2067 1122
rect 2119 1126 2123 1127
rect 2119 1121 2123 1122
rect 2151 1126 2155 1127
rect 2151 1121 2155 1122
rect 2191 1126 2195 1127
rect 2191 1121 2195 1122
rect 2239 1126 2243 1127
rect 2239 1121 2243 1122
rect 2271 1126 2275 1127
rect 2271 1121 2275 1122
rect 2327 1126 2331 1127
rect 2327 1121 2331 1122
rect 2351 1126 2355 1127
rect 2351 1121 2355 1122
rect 2415 1126 2419 1127
rect 2415 1121 2419 1122
rect 2583 1126 2587 1127
rect 2583 1121 2587 1122
rect 1006 1109 1007 1113
rect 1011 1109 1012 1113
rect 1006 1108 1012 1109
rect 1326 1112 1332 1113
rect 1326 1108 1327 1112
rect 1331 1108 1332 1112
rect 1368 1109 1370 1121
rect 1400 1110 1402 1121
rect 1480 1110 1482 1121
rect 1584 1110 1586 1121
rect 1688 1110 1690 1121
rect 1784 1110 1786 1121
rect 1880 1110 1882 1121
rect 1976 1110 1978 1121
rect 2064 1110 2066 1121
rect 2152 1110 2154 1121
rect 2240 1110 2242 1121
rect 2328 1110 2330 1121
rect 2416 1110 2418 1121
rect 1398 1109 1404 1110
rect 110 1107 116 1108
rect 1326 1107 1332 1108
rect 1366 1108 1372 1109
rect 1366 1104 1367 1108
rect 1371 1104 1372 1108
rect 1398 1105 1399 1109
rect 1403 1105 1404 1109
rect 1398 1104 1404 1105
rect 1478 1109 1484 1110
rect 1478 1105 1479 1109
rect 1483 1105 1484 1109
rect 1478 1104 1484 1105
rect 1582 1109 1588 1110
rect 1582 1105 1583 1109
rect 1587 1105 1588 1109
rect 1582 1104 1588 1105
rect 1686 1109 1692 1110
rect 1686 1105 1687 1109
rect 1691 1105 1692 1109
rect 1686 1104 1692 1105
rect 1782 1109 1788 1110
rect 1782 1105 1783 1109
rect 1787 1105 1788 1109
rect 1782 1104 1788 1105
rect 1878 1109 1884 1110
rect 1878 1105 1879 1109
rect 1883 1105 1884 1109
rect 1878 1104 1884 1105
rect 1974 1109 1980 1110
rect 1974 1105 1975 1109
rect 1979 1105 1980 1109
rect 1974 1104 1980 1105
rect 2062 1109 2068 1110
rect 2062 1105 2063 1109
rect 2067 1105 2068 1109
rect 2062 1104 2068 1105
rect 2150 1109 2156 1110
rect 2150 1105 2151 1109
rect 2155 1105 2156 1109
rect 2150 1104 2156 1105
rect 2238 1109 2244 1110
rect 2238 1105 2239 1109
rect 2243 1105 2244 1109
rect 2238 1104 2244 1105
rect 2326 1109 2332 1110
rect 2326 1105 2327 1109
rect 2331 1105 2332 1109
rect 2326 1104 2332 1105
rect 2414 1109 2420 1110
rect 2584 1109 2586 1121
rect 2414 1105 2415 1109
rect 2419 1105 2420 1109
rect 2414 1104 2420 1105
rect 2582 1108 2588 1109
rect 2582 1104 2583 1108
rect 2587 1104 2588 1108
rect 1366 1103 1372 1104
rect 2582 1103 2588 1104
rect 110 1095 116 1096
rect 110 1091 111 1095
rect 115 1091 116 1095
rect 110 1090 116 1091
rect 1326 1095 1332 1096
rect 1326 1091 1327 1095
rect 1331 1091 1332 1095
rect 1326 1090 1332 1091
rect 1366 1091 1372 1092
rect 112 1071 114 1090
rect 158 1086 164 1087
rect 158 1082 159 1086
rect 163 1082 164 1086
rect 158 1081 164 1082
rect 222 1086 228 1087
rect 222 1082 223 1086
rect 227 1082 228 1086
rect 222 1081 228 1082
rect 286 1086 292 1087
rect 286 1082 287 1086
rect 291 1082 292 1086
rect 286 1081 292 1082
rect 358 1086 364 1087
rect 358 1082 359 1086
rect 363 1082 364 1086
rect 358 1081 364 1082
rect 438 1086 444 1087
rect 438 1082 439 1086
rect 443 1082 444 1086
rect 438 1081 444 1082
rect 518 1086 524 1087
rect 518 1082 519 1086
rect 523 1082 524 1086
rect 518 1081 524 1082
rect 598 1086 604 1087
rect 598 1082 599 1086
rect 603 1082 604 1086
rect 598 1081 604 1082
rect 678 1086 684 1087
rect 678 1082 679 1086
rect 683 1082 684 1086
rect 678 1081 684 1082
rect 758 1086 764 1087
rect 758 1082 759 1086
rect 763 1082 764 1086
rect 758 1081 764 1082
rect 846 1086 852 1087
rect 846 1082 847 1086
rect 851 1082 852 1086
rect 846 1081 852 1082
rect 934 1086 940 1087
rect 934 1082 935 1086
rect 939 1082 940 1086
rect 934 1081 940 1082
rect 1022 1086 1028 1087
rect 1022 1082 1023 1086
rect 1027 1082 1028 1086
rect 1022 1081 1028 1082
rect 160 1071 162 1081
rect 224 1071 226 1081
rect 288 1071 290 1081
rect 360 1071 362 1081
rect 440 1071 442 1081
rect 520 1071 522 1081
rect 600 1071 602 1081
rect 680 1071 682 1081
rect 760 1071 762 1081
rect 848 1071 850 1081
rect 936 1071 938 1081
rect 1024 1071 1026 1081
rect 1328 1071 1330 1090
rect 1366 1087 1367 1091
rect 1371 1087 1372 1091
rect 1366 1086 1372 1087
rect 2582 1091 2588 1092
rect 2582 1087 2583 1091
rect 2587 1087 2588 1091
rect 2582 1086 2588 1087
rect 1368 1071 1370 1086
rect 1414 1082 1420 1083
rect 1414 1078 1415 1082
rect 1419 1078 1420 1082
rect 1414 1077 1420 1078
rect 1494 1082 1500 1083
rect 1494 1078 1495 1082
rect 1499 1078 1500 1082
rect 1494 1077 1500 1078
rect 1598 1082 1604 1083
rect 1598 1078 1599 1082
rect 1603 1078 1604 1082
rect 1598 1077 1604 1078
rect 1702 1082 1708 1083
rect 1702 1078 1703 1082
rect 1707 1078 1708 1082
rect 1702 1077 1708 1078
rect 1798 1082 1804 1083
rect 1798 1078 1799 1082
rect 1803 1078 1804 1082
rect 1798 1077 1804 1078
rect 1894 1082 1900 1083
rect 1894 1078 1895 1082
rect 1899 1078 1900 1082
rect 1894 1077 1900 1078
rect 1990 1082 1996 1083
rect 1990 1078 1991 1082
rect 1995 1078 1996 1082
rect 1990 1077 1996 1078
rect 2078 1082 2084 1083
rect 2078 1078 2079 1082
rect 2083 1078 2084 1082
rect 2078 1077 2084 1078
rect 2166 1082 2172 1083
rect 2166 1078 2167 1082
rect 2171 1078 2172 1082
rect 2166 1077 2172 1078
rect 2254 1082 2260 1083
rect 2254 1078 2255 1082
rect 2259 1078 2260 1082
rect 2254 1077 2260 1078
rect 2342 1082 2348 1083
rect 2342 1078 2343 1082
rect 2347 1078 2348 1082
rect 2342 1077 2348 1078
rect 2430 1082 2436 1083
rect 2430 1078 2431 1082
rect 2435 1078 2436 1082
rect 2430 1077 2436 1078
rect 1416 1071 1418 1077
rect 1496 1071 1498 1077
rect 1600 1071 1602 1077
rect 1704 1071 1706 1077
rect 1800 1071 1802 1077
rect 1896 1071 1898 1077
rect 1992 1071 1994 1077
rect 2080 1071 2082 1077
rect 2168 1071 2170 1077
rect 2256 1071 2258 1077
rect 2344 1071 2346 1077
rect 2432 1071 2434 1077
rect 2584 1071 2586 1086
rect 111 1070 115 1071
rect 111 1065 115 1066
rect 159 1070 163 1071
rect 159 1065 163 1066
rect 215 1070 219 1071
rect 215 1065 219 1066
rect 223 1070 227 1071
rect 223 1065 227 1066
rect 287 1070 291 1071
rect 287 1065 291 1066
rect 359 1070 363 1071
rect 359 1065 363 1066
rect 383 1070 387 1071
rect 383 1065 387 1066
rect 439 1070 443 1071
rect 439 1065 443 1066
rect 479 1070 483 1071
rect 479 1065 483 1066
rect 519 1070 523 1071
rect 519 1065 523 1066
rect 583 1070 587 1071
rect 583 1065 587 1066
rect 599 1070 603 1071
rect 599 1065 603 1066
rect 679 1070 683 1071
rect 679 1065 683 1066
rect 687 1070 691 1071
rect 687 1065 691 1066
rect 759 1070 763 1071
rect 759 1065 763 1066
rect 783 1070 787 1071
rect 783 1065 787 1066
rect 847 1070 851 1071
rect 847 1065 851 1066
rect 879 1070 883 1071
rect 879 1065 883 1066
rect 935 1070 939 1071
rect 935 1065 939 1066
rect 967 1070 971 1071
rect 967 1065 971 1066
rect 1023 1070 1027 1071
rect 1023 1065 1027 1066
rect 1063 1070 1067 1071
rect 1063 1065 1067 1066
rect 1159 1070 1163 1071
rect 1159 1065 1163 1066
rect 1327 1070 1331 1071
rect 1327 1065 1331 1066
rect 1367 1070 1371 1071
rect 1367 1065 1371 1066
rect 1415 1070 1419 1071
rect 1415 1065 1419 1066
rect 1495 1070 1499 1071
rect 1495 1065 1499 1066
rect 1511 1070 1515 1071
rect 1511 1065 1515 1066
rect 1599 1070 1603 1071
rect 1599 1065 1603 1066
rect 1631 1070 1635 1071
rect 1631 1065 1635 1066
rect 1703 1070 1707 1071
rect 1703 1065 1707 1066
rect 1751 1070 1755 1071
rect 1751 1065 1755 1066
rect 1799 1070 1803 1071
rect 1799 1065 1803 1066
rect 1871 1070 1875 1071
rect 1871 1065 1875 1066
rect 1895 1070 1899 1071
rect 1895 1065 1899 1066
rect 1991 1070 1995 1071
rect 1991 1065 1995 1066
rect 2079 1070 2083 1071
rect 2079 1065 2083 1066
rect 2103 1070 2107 1071
rect 2103 1065 2107 1066
rect 2167 1070 2171 1071
rect 2167 1065 2171 1066
rect 2199 1070 2203 1071
rect 2199 1065 2203 1066
rect 2255 1070 2259 1071
rect 2255 1065 2259 1066
rect 2295 1070 2299 1071
rect 2295 1065 2299 1066
rect 2343 1070 2347 1071
rect 2343 1065 2347 1066
rect 2383 1070 2387 1071
rect 2383 1065 2387 1066
rect 2431 1070 2435 1071
rect 2431 1065 2435 1066
rect 2471 1070 2475 1071
rect 2471 1065 2475 1066
rect 2543 1070 2547 1071
rect 2543 1065 2547 1066
rect 2583 1070 2587 1071
rect 2583 1065 2587 1066
rect 112 1050 114 1065
rect 160 1059 162 1065
rect 216 1059 218 1065
rect 288 1059 290 1065
rect 384 1059 386 1065
rect 480 1059 482 1065
rect 584 1059 586 1065
rect 688 1059 690 1065
rect 784 1059 786 1065
rect 880 1059 882 1065
rect 968 1059 970 1065
rect 1064 1059 1066 1065
rect 1160 1059 1162 1065
rect 158 1058 164 1059
rect 158 1054 159 1058
rect 163 1054 164 1058
rect 158 1053 164 1054
rect 214 1058 220 1059
rect 214 1054 215 1058
rect 219 1054 220 1058
rect 214 1053 220 1054
rect 286 1058 292 1059
rect 286 1054 287 1058
rect 291 1054 292 1058
rect 286 1053 292 1054
rect 382 1058 388 1059
rect 382 1054 383 1058
rect 387 1054 388 1058
rect 382 1053 388 1054
rect 478 1058 484 1059
rect 478 1054 479 1058
rect 483 1054 484 1058
rect 478 1053 484 1054
rect 582 1058 588 1059
rect 582 1054 583 1058
rect 587 1054 588 1058
rect 582 1053 588 1054
rect 686 1058 692 1059
rect 686 1054 687 1058
rect 691 1054 692 1058
rect 686 1053 692 1054
rect 782 1058 788 1059
rect 782 1054 783 1058
rect 787 1054 788 1058
rect 782 1053 788 1054
rect 878 1058 884 1059
rect 878 1054 879 1058
rect 883 1054 884 1058
rect 878 1053 884 1054
rect 966 1058 972 1059
rect 966 1054 967 1058
rect 971 1054 972 1058
rect 966 1053 972 1054
rect 1062 1058 1068 1059
rect 1062 1054 1063 1058
rect 1067 1054 1068 1058
rect 1062 1053 1068 1054
rect 1158 1058 1164 1059
rect 1158 1054 1159 1058
rect 1163 1054 1164 1058
rect 1158 1053 1164 1054
rect 1328 1050 1330 1065
rect 1368 1050 1370 1065
rect 1416 1059 1418 1065
rect 1512 1059 1514 1065
rect 1632 1059 1634 1065
rect 1752 1059 1754 1065
rect 1872 1059 1874 1065
rect 1992 1059 1994 1065
rect 2104 1059 2106 1065
rect 2200 1059 2202 1065
rect 2296 1059 2298 1065
rect 2384 1059 2386 1065
rect 2472 1059 2474 1065
rect 2544 1059 2546 1065
rect 1414 1058 1420 1059
rect 1414 1054 1415 1058
rect 1419 1054 1420 1058
rect 1414 1053 1420 1054
rect 1510 1058 1516 1059
rect 1510 1054 1511 1058
rect 1515 1054 1516 1058
rect 1510 1053 1516 1054
rect 1630 1058 1636 1059
rect 1630 1054 1631 1058
rect 1635 1054 1636 1058
rect 1630 1053 1636 1054
rect 1750 1058 1756 1059
rect 1750 1054 1751 1058
rect 1755 1054 1756 1058
rect 1750 1053 1756 1054
rect 1870 1058 1876 1059
rect 1870 1054 1871 1058
rect 1875 1054 1876 1058
rect 1870 1053 1876 1054
rect 1990 1058 1996 1059
rect 1990 1054 1991 1058
rect 1995 1054 1996 1058
rect 1990 1053 1996 1054
rect 2102 1058 2108 1059
rect 2102 1054 2103 1058
rect 2107 1054 2108 1058
rect 2102 1053 2108 1054
rect 2198 1058 2204 1059
rect 2198 1054 2199 1058
rect 2203 1054 2204 1058
rect 2198 1053 2204 1054
rect 2294 1058 2300 1059
rect 2294 1054 2295 1058
rect 2299 1054 2300 1058
rect 2294 1053 2300 1054
rect 2382 1058 2388 1059
rect 2382 1054 2383 1058
rect 2387 1054 2388 1058
rect 2382 1053 2388 1054
rect 2470 1058 2476 1059
rect 2470 1054 2471 1058
rect 2475 1054 2476 1058
rect 2470 1053 2476 1054
rect 2542 1058 2548 1059
rect 2542 1054 2543 1058
rect 2547 1054 2548 1058
rect 2542 1053 2548 1054
rect 2584 1050 2586 1065
rect 110 1049 116 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 1326 1049 1332 1050
rect 1326 1045 1327 1049
rect 1331 1045 1332 1049
rect 1326 1044 1332 1045
rect 1366 1049 1372 1050
rect 1366 1045 1367 1049
rect 1371 1045 1372 1049
rect 1366 1044 1372 1045
rect 2582 1049 2588 1050
rect 2582 1045 2583 1049
rect 2587 1045 2588 1049
rect 2582 1044 2588 1045
rect 110 1032 116 1033
rect 1326 1032 1332 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 110 1027 116 1028
rect 142 1031 148 1032
rect 142 1027 143 1031
rect 147 1027 148 1031
rect 112 1011 114 1027
rect 142 1026 148 1027
rect 198 1031 204 1032
rect 198 1027 199 1031
rect 203 1027 204 1031
rect 198 1026 204 1027
rect 270 1031 276 1032
rect 270 1027 271 1031
rect 275 1027 276 1031
rect 270 1026 276 1027
rect 366 1031 372 1032
rect 366 1027 367 1031
rect 371 1027 372 1031
rect 366 1026 372 1027
rect 462 1031 468 1032
rect 462 1027 463 1031
rect 467 1027 468 1031
rect 462 1026 468 1027
rect 566 1031 572 1032
rect 566 1027 567 1031
rect 571 1027 572 1031
rect 566 1026 572 1027
rect 670 1031 676 1032
rect 670 1027 671 1031
rect 675 1027 676 1031
rect 670 1026 676 1027
rect 766 1031 772 1032
rect 766 1027 767 1031
rect 771 1027 772 1031
rect 766 1026 772 1027
rect 862 1031 868 1032
rect 862 1027 863 1031
rect 867 1027 868 1031
rect 862 1026 868 1027
rect 950 1031 956 1032
rect 950 1027 951 1031
rect 955 1027 956 1031
rect 950 1026 956 1027
rect 1046 1031 1052 1032
rect 1046 1027 1047 1031
rect 1051 1027 1052 1031
rect 1046 1026 1052 1027
rect 1142 1031 1148 1032
rect 1142 1027 1143 1031
rect 1147 1027 1148 1031
rect 1326 1028 1327 1032
rect 1331 1028 1332 1032
rect 1326 1027 1332 1028
rect 1366 1032 1372 1033
rect 2582 1032 2588 1033
rect 1366 1028 1367 1032
rect 1371 1028 1372 1032
rect 1366 1027 1372 1028
rect 1398 1031 1404 1032
rect 1398 1027 1399 1031
rect 1403 1027 1404 1031
rect 1142 1026 1148 1027
rect 144 1011 146 1026
rect 200 1011 202 1026
rect 272 1011 274 1026
rect 368 1011 370 1026
rect 464 1011 466 1026
rect 568 1011 570 1026
rect 672 1011 674 1026
rect 768 1011 770 1026
rect 864 1011 866 1026
rect 952 1011 954 1026
rect 1048 1011 1050 1026
rect 1144 1011 1146 1026
rect 1328 1011 1330 1027
rect 1368 1011 1370 1027
rect 1398 1026 1404 1027
rect 1494 1031 1500 1032
rect 1494 1027 1495 1031
rect 1499 1027 1500 1031
rect 1494 1026 1500 1027
rect 1614 1031 1620 1032
rect 1614 1027 1615 1031
rect 1619 1027 1620 1031
rect 1614 1026 1620 1027
rect 1734 1031 1740 1032
rect 1734 1027 1735 1031
rect 1739 1027 1740 1031
rect 1734 1026 1740 1027
rect 1854 1031 1860 1032
rect 1854 1027 1855 1031
rect 1859 1027 1860 1031
rect 1854 1026 1860 1027
rect 1974 1031 1980 1032
rect 1974 1027 1975 1031
rect 1979 1027 1980 1031
rect 1974 1026 1980 1027
rect 2086 1031 2092 1032
rect 2086 1027 2087 1031
rect 2091 1027 2092 1031
rect 2086 1026 2092 1027
rect 2182 1031 2188 1032
rect 2182 1027 2183 1031
rect 2187 1027 2188 1031
rect 2182 1026 2188 1027
rect 2278 1031 2284 1032
rect 2278 1027 2279 1031
rect 2283 1027 2284 1031
rect 2278 1026 2284 1027
rect 2366 1031 2372 1032
rect 2366 1027 2367 1031
rect 2371 1027 2372 1031
rect 2366 1026 2372 1027
rect 2454 1031 2460 1032
rect 2454 1027 2455 1031
rect 2459 1027 2460 1031
rect 2454 1026 2460 1027
rect 2526 1031 2532 1032
rect 2526 1027 2527 1031
rect 2531 1027 2532 1031
rect 2582 1028 2583 1032
rect 2587 1028 2588 1032
rect 2582 1027 2588 1028
rect 2526 1026 2532 1027
rect 1400 1011 1402 1026
rect 1496 1011 1498 1026
rect 1616 1011 1618 1026
rect 1736 1011 1738 1026
rect 1856 1011 1858 1026
rect 1976 1011 1978 1026
rect 2088 1011 2090 1026
rect 2184 1011 2186 1026
rect 2280 1011 2282 1026
rect 2368 1011 2370 1026
rect 2456 1011 2458 1026
rect 2528 1011 2530 1026
rect 2584 1011 2586 1027
rect 111 1010 115 1011
rect 111 1005 115 1006
rect 143 1010 147 1011
rect 143 1005 147 1006
rect 199 1010 203 1011
rect 199 1005 203 1006
rect 271 1010 275 1011
rect 271 1005 275 1006
rect 279 1010 283 1011
rect 279 1005 283 1006
rect 367 1010 371 1011
rect 367 1005 371 1006
rect 383 1010 387 1011
rect 383 1005 387 1006
rect 463 1010 467 1011
rect 463 1005 467 1006
rect 495 1010 499 1011
rect 495 1005 499 1006
rect 567 1010 571 1011
rect 567 1005 571 1006
rect 615 1010 619 1011
rect 615 1005 619 1006
rect 671 1010 675 1011
rect 671 1005 675 1006
rect 727 1010 731 1011
rect 727 1005 731 1006
rect 767 1010 771 1011
rect 767 1005 771 1006
rect 839 1010 843 1011
rect 839 1005 843 1006
rect 863 1010 867 1011
rect 863 1005 867 1006
rect 951 1010 955 1011
rect 951 1005 955 1006
rect 1047 1010 1051 1011
rect 1047 1005 1051 1006
rect 1055 1010 1059 1011
rect 1055 1005 1059 1006
rect 1143 1010 1147 1011
rect 1143 1005 1147 1006
rect 1159 1010 1163 1011
rect 1159 1005 1163 1006
rect 1271 1010 1275 1011
rect 1271 1005 1275 1006
rect 1327 1010 1331 1011
rect 1327 1005 1331 1006
rect 1367 1010 1371 1011
rect 1367 1005 1371 1006
rect 1399 1010 1403 1011
rect 1399 1005 1403 1006
rect 1487 1010 1491 1011
rect 1487 1005 1491 1006
rect 1495 1010 1499 1011
rect 1495 1005 1499 1006
rect 1583 1010 1587 1011
rect 1583 1005 1587 1006
rect 1615 1010 1619 1011
rect 1615 1005 1619 1006
rect 1695 1010 1699 1011
rect 1695 1005 1699 1006
rect 1735 1010 1739 1011
rect 1735 1005 1739 1006
rect 1807 1010 1811 1011
rect 1807 1005 1811 1006
rect 1855 1010 1859 1011
rect 1855 1005 1859 1006
rect 1919 1010 1923 1011
rect 1919 1005 1923 1006
rect 1975 1010 1979 1011
rect 1975 1005 1979 1006
rect 2023 1010 2027 1011
rect 2023 1005 2027 1006
rect 2087 1010 2091 1011
rect 2087 1005 2091 1006
rect 2119 1010 2123 1011
rect 2119 1005 2123 1006
rect 2183 1010 2187 1011
rect 2183 1005 2187 1006
rect 2215 1010 2219 1011
rect 2215 1005 2219 1006
rect 2279 1010 2283 1011
rect 2279 1005 2283 1006
rect 2303 1010 2307 1011
rect 2303 1005 2307 1006
rect 2367 1010 2371 1011
rect 2367 1005 2371 1006
rect 2383 1010 2387 1011
rect 2383 1005 2387 1006
rect 2455 1010 2459 1011
rect 2455 1005 2459 1006
rect 2463 1010 2467 1011
rect 2463 1005 2467 1006
rect 2527 1010 2531 1011
rect 2527 1005 2531 1006
rect 2583 1010 2587 1011
rect 2583 1005 2587 1006
rect 112 993 114 1005
rect 144 994 146 1005
rect 200 994 202 1005
rect 280 994 282 1005
rect 384 994 386 1005
rect 496 994 498 1005
rect 616 994 618 1005
rect 728 994 730 1005
rect 840 994 842 1005
rect 952 994 954 1005
rect 1056 994 1058 1005
rect 1160 994 1162 1005
rect 1272 994 1274 1005
rect 142 993 148 994
rect 110 992 116 993
rect 110 988 111 992
rect 115 988 116 992
rect 142 989 143 993
rect 147 989 148 993
rect 142 988 148 989
rect 198 993 204 994
rect 198 989 199 993
rect 203 989 204 993
rect 198 988 204 989
rect 278 993 284 994
rect 278 989 279 993
rect 283 989 284 993
rect 278 988 284 989
rect 382 993 388 994
rect 382 989 383 993
rect 387 989 388 993
rect 382 988 388 989
rect 494 993 500 994
rect 494 989 495 993
rect 499 989 500 993
rect 494 988 500 989
rect 614 993 620 994
rect 614 989 615 993
rect 619 989 620 993
rect 614 988 620 989
rect 726 993 732 994
rect 726 989 727 993
rect 731 989 732 993
rect 726 988 732 989
rect 838 993 844 994
rect 838 989 839 993
rect 843 989 844 993
rect 838 988 844 989
rect 950 993 956 994
rect 950 989 951 993
rect 955 989 956 993
rect 950 988 956 989
rect 1054 993 1060 994
rect 1054 989 1055 993
rect 1059 989 1060 993
rect 1054 988 1060 989
rect 1158 993 1164 994
rect 1158 989 1159 993
rect 1163 989 1164 993
rect 1158 988 1164 989
rect 1270 993 1276 994
rect 1328 993 1330 1005
rect 1368 993 1370 1005
rect 1488 994 1490 1005
rect 1584 994 1586 1005
rect 1696 994 1698 1005
rect 1808 994 1810 1005
rect 1920 994 1922 1005
rect 2024 994 2026 1005
rect 2120 994 2122 1005
rect 2216 994 2218 1005
rect 2304 994 2306 1005
rect 2384 994 2386 1005
rect 2464 994 2466 1005
rect 2528 994 2530 1005
rect 1486 993 1492 994
rect 1270 989 1271 993
rect 1275 989 1276 993
rect 1270 988 1276 989
rect 1326 992 1332 993
rect 1326 988 1327 992
rect 1331 988 1332 992
rect 110 987 116 988
rect 1326 987 1332 988
rect 1366 992 1372 993
rect 1366 988 1367 992
rect 1371 988 1372 992
rect 1486 989 1487 993
rect 1491 989 1492 993
rect 1486 988 1492 989
rect 1582 993 1588 994
rect 1582 989 1583 993
rect 1587 989 1588 993
rect 1582 988 1588 989
rect 1694 993 1700 994
rect 1694 989 1695 993
rect 1699 989 1700 993
rect 1694 988 1700 989
rect 1806 993 1812 994
rect 1806 989 1807 993
rect 1811 989 1812 993
rect 1806 988 1812 989
rect 1918 993 1924 994
rect 1918 989 1919 993
rect 1923 989 1924 993
rect 1918 988 1924 989
rect 2022 993 2028 994
rect 2022 989 2023 993
rect 2027 989 2028 993
rect 2022 988 2028 989
rect 2118 993 2124 994
rect 2118 989 2119 993
rect 2123 989 2124 993
rect 2118 988 2124 989
rect 2214 993 2220 994
rect 2214 989 2215 993
rect 2219 989 2220 993
rect 2214 988 2220 989
rect 2302 993 2308 994
rect 2302 989 2303 993
rect 2307 989 2308 993
rect 2302 988 2308 989
rect 2382 993 2388 994
rect 2382 989 2383 993
rect 2387 989 2388 993
rect 2382 988 2388 989
rect 2462 993 2468 994
rect 2462 989 2463 993
rect 2467 989 2468 993
rect 2462 988 2468 989
rect 2526 993 2532 994
rect 2584 993 2586 1005
rect 2526 989 2527 993
rect 2531 989 2532 993
rect 2526 988 2532 989
rect 2582 992 2588 993
rect 2582 988 2583 992
rect 2587 988 2588 992
rect 1366 987 1372 988
rect 2582 987 2588 988
rect 110 975 116 976
rect 110 971 111 975
rect 115 971 116 975
rect 110 970 116 971
rect 1326 975 1332 976
rect 1326 971 1327 975
rect 1331 971 1332 975
rect 1326 970 1332 971
rect 1366 975 1372 976
rect 1366 971 1367 975
rect 1371 971 1372 975
rect 1366 970 1372 971
rect 2582 975 2588 976
rect 2582 971 2583 975
rect 2587 971 2588 975
rect 2582 970 2588 971
rect 112 947 114 970
rect 158 966 164 967
rect 158 962 159 966
rect 163 962 164 966
rect 158 961 164 962
rect 214 966 220 967
rect 214 962 215 966
rect 219 962 220 966
rect 214 961 220 962
rect 294 966 300 967
rect 294 962 295 966
rect 299 962 300 966
rect 294 961 300 962
rect 398 966 404 967
rect 398 962 399 966
rect 403 962 404 966
rect 398 961 404 962
rect 510 966 516 967
rect 510 962 511 966
rect 515 962 516 966
rect 510 961 516 962
rect 630 966 636 967
rect 630 962 631 966
rect 635 962 636 966
rect 630 961 636 962
rect 742 966 748 967
rect 742 962 743 966
rect 747 962 748 966
rect 742 961 748 962
rect 854 966 860 967
rect 854 962 855 966
rect 859 962 860 966
rect 854 961 860 962
rect 966 966 972 967
rect 966 962 967 966
rect 971 962 972 966
rect 966 961 972 962
rect 1070 966 1076 967
rect 1070 962 1071 966
rect 1075 962 1076 966
rect 1070 961 1076 962
rect 1174 966 1180 967
rect 1174 962 1175 966
rect 1179 962 1180 966
rect 1174 961 1180 962
rect 1286 966 1292 967
rect 1286 962 1287 966
rect 1291 962 1292 966
rect 1286 961 1292 962
rect 160 947 162 961
rect 216 947 218 961
rect 296 947 298 961
rect 400 947 402 961
rect 512 947 514 961
rect 632 947 634 961
rect 744 947 746 961
rect 856 947 858 961
rect 968 947 970 961
rect 1072 947 1074 961
rect 1176 947 1178 961
rect 1288 947 1290 961
rect 1328 947 1330 970
rect 1368 947 1370 970
rect 1502 966 1508 967
rect 1502 962 1503 966
rect 1507 962 1508 966
rect 1502 961 1508 962
rect 1598 966 1604 967
rect 1598 962 1599 966
rect 1603 962 1604 966
rect 1598 961 1604 962
rect 1710 966 1716 967
rect 1710 962 1711 966
rect 1715 962 1716 966
rect 1710 961 1716 962
rect 1822 966 1828 967
rect 1822 962 1823 966
rect 1827 962 1828 966
rect 1822 961 1828 962
rect 1934 966 1940 967
rect 1934 962 1935 966
rect 1939 962 1940 966
rect 1934 961 1940 962
rect 2038 966 2044 967
rect 2038 962 2039 966
rect 2043 962 2044 966
rect 2038 961 2044 962
rect 2134 966 2140 967
rect 2134 962 2135 966
rect 2139 962 2140 966
rect 2134 961 2140 962
rect 2230 966 2236 967
rect 2230 962 2231 966
rect 2235 962 2236 966
rect 2230 961 2236 962
rect 2318 966 2324 967
rect 2318 962 2319 966
rect 2323 962 2324 966
rect 2318 961 2324 962
rect 2398 966 2404 967
rect 2398 962 2399 966
rect 2403 962 2404 966
rect 2398 961 2404 962
rect 2478 966 2484 967
rect 2478 962 2479 966
rect 2483 962 2484 966
rect 2478 961 2484 962
rect 2542 966 2548 967
rect 2542 962 2543 966
rect 2547 962 2548 966
rect 2542 961 2548 962
rect 1504 947 1506 961
rect 1600 947 1602 961
rect 1712 947 1714 961
rect 1824 947 1826 961
rect 1936 947 1938 961
rect 2040 947 2042 961
rect 2136 947 2138 961
rect 2232 947 2234 961
rect 2320 947 2322 961
rect 2400 947 2402 961
rect 2480 947 2482 961
rect 2544 947 2546 961
rect 2584 947 2586 970
rect 111 946 115 947
rect 111 941 115 942
rect 159 946 163 947
rect 159 941 163 942
rect 215 946 219 947
rect 215 941 219 942
rect 287 946 291 947
rect 287 941 291 942
rect 295 946 299 947
rect 295 941 299 942
rect 375 946 379 947
rect 375 941 379 942
rect 399 946 403 947
rect 399 941 403 942
rect 471 946 475 947
rect 471 941 475 942
rect 511 946 515 947
rect 511 941 515 942
rect 567 946 571 947
rect 567 941 571 942
rect 631 946 635 947
rect 631 941 635 942
rect 671 946 675 947
rect 671 941 675 942
rect 743 946 747 947
rect 743 941 747 942
rect 767 946 771 947
rect 767 941 771 942
rect 855 946 859 947
rect 855 941 859 942
rect 863 946 867 947
rect 863 941 867 942
rect 959 946 963 947
rect 959 941 963 942
rect 967 946 971 947
rect 967 941 971 942
rect 1047 946 1051 947
rect 1047 941 1051 942
rect 1071 946 1075 947
rect 1071 941 1075 942
rect 1135 946 1139 947
rect 1135 941 1139 942
rect 1175 946 1179 947
rect 1175 941 1179 942
rect 1223 946 1227 947
rect 1223 941 1227 942
rect 1287 946 1291 947
rect 1287 941 1291 942
rect 1327 946 1331 947
rect 1327 941 1331 942
rect 1367 946 1371 947
rect 1367 941 1371 942
rect 1415 946 1419 947
rect 1415 941 1419 942
rect 1503 946 1507 947
rect 1503 941 1507 942
rect 1535 946 1539 947
rect 1535 941 1539 942
rect 1599 946 1603 947
rect 1599 941 1603 942
rect 1671 946 1675 947
rect 1671 941 1675 942
rect 1711 946 1715 947
rect 1711 941 1715 942
rect 1807 946 1811 947
rect 1807 941 1811 942
rect 1823 946 1827 947
rect 1823 941 1827 942
rect 1935 946 1939 947
rect 1935 941 1939 942
rect 2039 946 2043 947
rect 2039 941 2043 942
rect 2055 946 2059 947
rect 2055 941 2059 942
rect 2135 946 2139 947
rect 2135 941 2139 942
rect 2167 946 2171 947
rect 2167 941 2171 942
rect 2231 946 2235 947
rect 2231 941 2235 942
rect 2271 946 2275 947
rect 2271 941 2275 942
rect 2319 946 2323 947
rect 2319 941 2323 942
rect 2367 946 2371 947
rect 2367 941 2371 942
rect 2399 946 2403 947
rect 2399 941 2403 942
rect 2463 946 2467 947
rect 2463 941 2467 942
rect 2479 946 2483 947
rect 2479 941 2483 942
rect 2543 946 2547 947
rect 2543 941 2547 942
rect 2583 946 2587 947
rect 2583 941 2587 942
rect 112 926 114 941
rect 160 935 162 941
rect 216 935 218 941
rect 288 935 290 941
rect 376 935 378 941
rect 472 935 474 941
rect 568 935 570 941
rect 672 935 674 941
rect 768 935 770 941
rect 864 935 866 941
rect 960 935 962 941
rect 1048 935 1050 941
rect 1136 935 1138 941
rect 1224 935 1226 941
rect 1288 935 1290 941
rect 158 934 164 935
rect 158 930 159 934
rect 163 930 164 934
rect 158 929 164 930
rect 214 934 220 935
rect 214 930 215 934
rect 219 930 220 934
rect 214 929 220 930
rect 286 934 292 935
rect 286 930 287 934
rect 291 930 292 934
rect 286 929 292 930
rect 374 934 380 935
rect 374 930 375 934
rect 379 930 380 934
rect 374 929 380 930
rect 470 934 476 935
rect 470 930 471 934
rect 475 930 476 934
rect 470 929 476 930
rect 566 934 572 935
rect 566 930 567 934
rect 571 930 572 934
rect 566 929 572 930
rect 670 934 676 935
rect 670 930 671 934
rect 675 930 676 934
rect 670 929 676 930
rect 766 934 772 935
rect 766 930 767 934
rect 771 930 772 934
rect 766 929 772 930
rect 862 934 868 935
rect 862 930 863 934
rect 867 930 868 934
rect 862 929 868 930
rect 958 934 964 935
rect 958 930 959 934
rect 963 930 964 934
rect 958 929 964 930
rect 1046 934 1052 935
rect 1046 930 1047 934
rect 1051 930 1052 934
rect 1046 929 1052 930
rect 1134 934 1140 935
rect 1134 930 1135 934
rect 1139 930 1140 934
rect 1134 929 1140 930
rect 1222 934 1228 935
rect 1222 930 1223 934
rect 1227 930 1228 934
rect 1222 929 1228 930
rect 1286 934 1292 935
rect 1286 930 1287 934
rect 1291 930 1292 934
rect 1286 929 1292 930
rect 1328 926 1330 941
rect 1368 926 1370 941
rect 1416 935 1418 941
rect 1536 935 1538 941
rect 1672 935 1674 941
rect 1808 935 1810 941
rect 1936 935 1938 941
rect 2056 935 2058 941
rect 2168 935 2170 941
rect 2272 935 2274 941
rect 2368 935 2370 941
rect 2464 935 2466 941
rect 2544 935 2546 941
rect 1414 934 1420 935
rect 1414 930 1415 934
rect 1419 930 1420 934
rect 1414 929 1420 930
rect 1534 934 1540 935
rect 1534 930 1535 934
rect 1539 930 1540 934
rect 1534 929 1540 930
rect 1670 934 1676 935
rect 1670 930 1671 934
rect 1675 930 1676 934
rect 1670 929 1676 930
rect 1806 934 1812 935
rect 1806 930 1807 934
rect 1811 930 1812 934
rect 1806 929 1812 930
rect 1934 934 1940 935
rect 1934 930 1935 934
rect 1939 930 1940 934
rect 1934 929 1940 930
rect 2054 934 2060 935
rect 2054 930 2055 934
rect 2059 930 2060 934
rect 2054 929 2060 930
rect 2166 934 2172 935
rect 2166 930 2167 934
rect 2171 930 2172 934
rect 2166 929 2172 930
rect 2270 934 2276 935
rect 2270 930 2271 934
rect 2275 930 2276 934
rect 2270 929 2276 930
rect 2366 934 2372 935
rect 2366 930 2367 934
rect 2371 930 2372 934
rect 2366 929 2372 930
rect 2462 934 2468 935
rect 2462 930 2463 934
rect 2467 930 2468 934
rect 2462 929 2468 930
rect 2542 934 2548 935
rect 2542 930 2543 934
rect 2547 930 2548 934
rect 2542 929 2548 930
rect 2584 926 2586 941
rect 110 925 116 926
rect 110 921 111 925
rect 115 921 116 925
rect 110 920 116 921
rect 1326 925 1332 926
rect 1326 921 1327 925
rect 1331 921 1332 925
rect 1326 920 1332 921
rect 1366 925 1372 926
rect 1366 921 1367 925
rect 1371 921 1372 925
rect 1366 920 1372 921
rect 2582 925 2588 926
rect 2582 921 2583 925
rect 2587 921 2588 925
rect 2582 920 2588 921
rect 110 908 116 909
rect 1326 908 1332 909
rect 110 904 111 908
rect 115 904 116 908
rect 110 903 116 904
rect 142 907 148 908
rect 142 903 143 907
rect 147 903 148 907
rect 112 887 114 903
rect 142 902 148 903
rect 198 907 204 908
rect 198 903 199 907
rect 203 903 204 907
rect 198 902 204 903
rect 270 907 276 908
rect 270 903 271 907
rect 275 903 276 907
rect 270 902 276 903
rect 358 907 364 908
rect 358 903 359 907
rect 363 903 364 907
rect 358 902 364 903
rect 454 907 460 908
rect 454 903 455 907
rect 459 903 460 907
rect 454 902 460 903
rect 550 907 556 908
rect 550 903 551 907
rect 555 903 556 907
rect 550 902 556 903
rect 654 907 660 908
rect 654 903 655 907
rect 659 903 660 907
rect 654 902 660 903
rect 750 907 756 908
rect 750 903 751 907
rect 755 903 756 907
rect 750 902 756 903
rect 846 907 852 908
rect 846 903 847 907
rect 851 903 852 907
rect 846 902 852 903
rect 942 907 948 908
rect 942 903 943 907
rect 947 903 948 907
rect 942 902 948 903
rect 1030 907 1036 908
rect 1030 903 1031 907
rect 1035 903 1036 907
rect 1030 902 1036 903
rect 1118 907 1124 908
rect 1118 903 1119 907
rect 1123 903 1124 907
rect 1118 902 1124 903
rect 1206 907 1212 908
rect 1206 903 1207 907
rect 1211 903 1212 907
rect 1206 902 1212 903
rect 1270 907 1276 908
rect 1270 903 1271 907
rect 1275 903 1276 907
rect 1326 904 1327 908
rect 1331 904 1332 908
rect 1326 903 1332 904
rect 1366 908 1372 909
rect 2582 908 2588 909
rect 1366 904 1367 908
rect 1371 904 1372 908
rect 1366 903 1372 904
rect 1398 907 1404 908
rect 1398 903 1399 907
rect 1403 903 1404 907
rect 1270 902 1276 903
rect 144 887 146 902
rect 200 887 202 902
rect 272 887 274 902
rect 360 887 362 902
rect 456 887 458 902
rect 552 887 554 902
rect 656 887 658 902
rect 752 887 754 902
rect 848 887 850 902
rect 944 887 946 902
rect 1032 887 1034 902
rect 1120 887 1122 902
rect 1208 887 1210 902
rect 1272 887 1274 902
rect 1328 887 1330 903
rect 1368 887 1370 903
rect 1398 902 1404 903
rect 1518 907 1524 908
rect 1518 903 1519 907
rect 1523 903 1524 907
rect 1518 902 1524 903
rect 1654 907 1660 908
rect 1654 903 1655 907
rect 1659 903 1660 907
rect 1654 902 1660 903
rect 1790 907 1796 908
rect 1790 903 1791 907
rect 1795 903 1796 907
rect 1790 902 1796 903
rect 1918 907 1924 908
rect 1918 903 1919 907
rect 1923 903 1924 907
rect 1918 902 1924 903
rect 2038 907 2044 908
rect 2038 903 2039 907
rect 2043 903 2044 907
rect 2038 902 2044 903
rect 2150 907 2156 908
rect 2150 903 2151 907
rect 2155 903 2156 907
rect 2150 902 2156 903
rect 2254 907 2260 908
rect 2254 903 2255 907
rect 2259 903 2260 907
rect 2254 902 2260 903
rect 2350 907 2356 908
rect 2350 903 2351 907
rect 2355 903 2356 907
rect 2350 902 2356 903
rect 2446 907 2452 908
rect 2446 903 2447 907
rect 2451 903 2452 907
rect 2446 902 2452 903
rect 2526 907 2532 908
rect 2526 903 2527 907
rect 2531 903 2532 907
rect 2582 904 2583 908
rect 2587 904 2588 908
rect 2582 903 2588 904
rect 2526 902 2532 903
rect 1400 887 1402 902
rect 1520 887 1522 902
rect 1656 887 1658 902
rect 1792 887 1794 902
rect 1920 887 1922 902
rect 2040 887 2042 902
rect 2152 887 2154 902
rect 2256 887 2258 902
rect 2352 887 2354 902
rect 2448 887 2450 902
rect 2528 887 2530 902
rect 2584 887 2586 903
rect 111 886 115 887
rect 111 881 115 882
rect 143 886 147 887
rect 143 881 147 882
rect 183 886 187 887
rect 183 881 187 882
rect 199 886 203 887
rect 199 881 203 882
rect 239 886 243 887
rect 239 881 243 882
rect 271 886 275 887
rect 271 881 275 882
rect 303 886 307 887
rect 303 881 307 882
rect 359 886 363 887
rect 359 881 363 882
rect 375 886 379 887
rect 375 881 379 882
rect 455 886 459 887
rect 455 881 459 882
rect 543 886 547 887
rect 543 881 547 882
rect 551 886 555 887
rect 551 881 555 882
rect 639 886 643 887
rect 639 881 643 882
rect 655 886 659 887
rect 655 881 659 882
rect 743 886 747 887
rect 743 881 747 882
rect 751 886 755 887
rect 751 881 755 882
rect 847 886 851 887
rect 847 881 851 882
rect 855 886 859 887
rect 855 881 859 882
rect 943 886 947 887
rect 943 881 947 882
rect 967 886 971 887
rect 967 881 971 882
rect 1031 886 1035 887
rect 1031 881 1035 882
rect 1087 886 1091 887
rect 1087 881 1091 882
rect 1119 886 1123 887
rect 1119 881 1123 882
rect 1207 886 1211 887
rect 1207 881 1211 882
rect 1215 886 1219 887
rect 1215 881 1219 882
rect 1271 886 1275 887
rect 1271 881 1275 882
rect 1327 886 1331 887
rect 1327 881 1331 882
rect 1367 886 1371 887
rect 1367 881 1371 882
rect 1399 886 1403 887
rect 1399 881 1403 882
rect 1455 886 1459 887
rect 1455 881 1459 882
rect 1519 886 1523 887
rect 1519 881 1523 882
rect 1607 886 1611 887
rect 1607 881 1611 882
rect 1655 886 1659 887
rect 1655 881 1659 882
rect 1695 886 1699 887
rect 1695 881 1699 882
rect 1791 886 1795 887
rect 1791 881 1795 882
rect 1895 886 1899 887
rect 1895 881 1899 882
rect 1919 886 1923 887
rect 1919 881 1923 882
rect 1999 886 2003 887
rect 1999 881 2003 882
rect 2039 886 2043 887
rect 2039 881 2043 882
rect 2103 886 2107 887
rect 2103 881 2107 882
rect 2151 886 2155 887
rect 2151 881 2155 882
rect 2207 886 2211 887
rect 2207 881 2211 882
rect 2255 886 2259 887
rect 2255 881 2259 882
rect 2311 886 2315 887
rect 2311 881 2315 882
rect 2351 886 2355 887
rect 2351 881 2355 882
rect 2423 886 2427 887
rect 2423 881 2427 882
rect 2447 886 2451 887
rect 2447 881 2451 882
rect 2527 886 2531 887
rect 2527 881 2531 882
rect 2583 886 2587 887
rect 2583 881 2587 882
rect 112 869 114 881
rect 184 870 186 881
rect 240 870 242 881
rect 304 870 306 881
rect 376 870 378 881
rect 456 870 458 881
rect 544 870 546 881
rect 640 870 642 881
rect 744 870 746 881
rect 856 870 858 881
rect 968 870 970 881
rect 1088 870 1090 881
rect 1216 870 1218 881
rect 182 869 188 870
rect 110 868 116 869
rect 110 864 111 868
rect 115 864 116 868
rect 182 865 183 869
rect 187 865 188 869
rect 182 864 188 865
rect 238 869 244 870
rect 238 865 239 869
rect 243 865 244 869
rect 238 864 244 865
rect 302 869 308 870
rect 302 865 303 869
rect 307 865 308 869
rect 302 864 308 865
rect 374 869 380 870
rect 374 865 375 869
rect 379 865 380 869
rect 374 864 380 865
rect 454 869 460 870
rect 454 865 455 869
rect 459 865 460 869
rect 454 864 460 865
rect 542 869 548 870
rect 542 865 543 869
rect 547 865 548 869
rect 542 864 548 865
rect 638 869 644 870
rect 638 865 639 869
rect 643 865 644 869
rect 638 864 644 865
rect 742 869 748 870
rect 742 865 743 869
rect 747 865 748 869
rect 742 864 748 865
rect 854 869 860 870
rect 854 865 855 869
rect 859 865 860 869
rect 854 864 860 865
rect 966 869 972 870
rect 966 865 967 869
rect 971 865 972 869
rect 966 864 972 865
rect 1086 869 1092 870
rect 1086 865 1087 869
rect 1091 865 1092 869
rect 1086 864 1092 865
rect 1214 869 1220 870
rect 1328 869 1330 881
rect 1368 869 1370 881
rect 1400 870 1402 881
rect 1456 870 1458 881
rect 1520 870 1522 881
rect 1608 870 1610 881
rect 1696 870 1698 881
rect 1792 870 1794 881
rect 1896 870 1898 881
rect 2000 870 2002 881
rect 2104 870 2106 881
rect 2208 870 2210 881
rect 2312 870 2314 881
rect 2424 870 2426 881
rect 2528 870 2530 881
rect 1398 869 1404 870
rect 1214 865 1215 869
rect 1219 865 1220 869
rect 1214 864 1220 865
rect 1326 868 1332 869
rect 1326 864 1327 868
rect 1331 864 1332 868
rect 110 863 116 864
rect 1326 863 1332 864
rect 1366 868 1372 869
rect 1366 864 1367 868
rect 1371 864 1372 868
rect 1398 865 1399 869
rect 1403 865 1404 869
rect 1398 864 1404 865
rect 1454 869 1460 870
rect 1454 865 1455 869
rect 1459 865 1460 869
rect 1454 864 1460 865
rect 1518 869 1524 870
rect 1518 865 1519 869
rect 1523 865 1524 869
rect 1518 864 1524 865
rect 1606 869 1612 870
rect 1606 865 1607 869
rect 1611 865 1612 869
rect 1606 864 1612 865
rect 1694 869 1700 870
rect 1694 865 1695 869
rect 1699 865 1700 869
rect 1694 864 1700 865
rect 1790 869 1796 870
rect 1790 865 1791 869
rect 1795 865 1796 869
rect 1790 864 1796 865
rect 1894 869 1900 870
rect 1894 865 1895 869
rect 1899 865 1900 869
rect 1894 864 1900 865
rect 1998 869 2004 870
rect 1998 865 1999 869
rect 2003 865 2004 869
rect 1998 864 2004 865
rect 2102 869 2108 870
rect 2102 865 2103 869
rect 2107 865 2108 869
rect 2102 864 2108 865
rect 2206 869 2212 870
rect 2206 865 2207 869
rect 2211 865 2212 869
rect 2206 864 2212 865
rect 2310 869 2316 870
rect 2310 865 2311 869
rect 2315 865 2316 869
rect 2310 864 2316 865
rect 2422 869 2428 870
rect 2422 865 2423 869
rect 2427 865 2428 869
rect 2422 864 2428 865
rect 2526 869 2532 870
rect 2584 869 2586 881
rect 2526 865 2527 869
rect 2531 865 2532 869
rect 2526 864 2532 865
rect 2582 868 2588 869
rect 2582 864 2583 868
rect 2587 864 2588 868
rect 1366 863 1372 864
rect 2582 863 2588 864
rect 110 851 116 852
rect 110 847 111 851
rect 115 847 116 851
rect 110 846 116 847
rect 1326 851 1332 852
rect 1326 847 1327 851
rect 1331 847 1332 851
rect 1326 846 1332 847
rect 1366 851 1372 852
rect 1366 847 1367 851
rect 1371 847 1372 851
rect 1366 846 1372 847
rect 2582 851 2588 852
rect 2582 847 2583 851
rect 2587 847 2588 851
rect 2582 846 2588 847
rect 112 823 114 846
rect 198 842 204 843
rect 198 838 199 842
rect 203 838 204 842
rect 198 837 204 838
rect 254 842 260 843
rect 254 838 255 842
rect 259 838 260 842
rect 254 837 260 838
rect 318 842 324 843
rect 318 838 319 842
rect 323 838 324 842
rect 318 837 324 838
rect 390 842 396 843
rect 390 838 391 842
rect 395 838 396 842
rect 390 837 396 838
rect 470 842 476 843
rect 470 838 471 842
rect 475 838 476 842
rect 470 837 476 838
rect 558 842 564 843
rect 558 838 559 842
rect 563 838 564 842
rect 558 837 564 838
rect 654 842 660 843
rect 654 838 655 842
rect 659 838 660 842
rect 654 837 660 838
rect 758 842 764 843
rect 758 838 759 842
rect 763 838 764 842
rect 758 837 764 838
rect 870 842 876 843
rect 870 838 871 842
rect 875 838 876 842
rect 870 837 876 838
rect 982 842 988 843
rect 982 838 983 842
rect 987 838 988 842
rect 982 837 988 838
rect 1102 842 1108 843
rect 1102 838 1103 842
rect 1107 838 1108 842
rect 1102 837 1108 838
rect 1230 842 1236 843
rect 1230 838 1231 842
rect 1235 838 1236 842
rect 1230 837 1236 838
rect 200 823 202 837
rect 256 823 258 837
rect 320 823 322 837
rect 392 823 394 837
rect 472 823 474 837
rect 560 823 562 837
rect 656 823 658 837
rect 760 823 762 837
rect 872 823 874 837
rect 984 823 986 837
rect 1104 823 1106 837
rect 1232 823 1234 837
rect 1328 823 1330 846
rect 1368 827 1370 846
rect 1414 842 1420 843
rect 1414 838 1415 842
rect 1419 838 1420 842
rect 1414 837 1420 838
rect 1470 842 1476 843
rect 1470 838 1471 842
rect 1475 838 1476 842
rect 1470 837 1476 838
rect 1534 842 1540 843
rect 1534 838 1535 842
rect 1539 838 1540 842
rect 1534 837 1540 838
rect 1622 842 1628 843
rect 1622 838 1623 842
rect 1627 838 1628 842
rect 1622 837 1628 838
rect 1710 842 1716 843
rect 1710 838 1711 842
rect 1715 838 1716 842
rect 1710 837 1716 838
rect 1806 842 1812 843
rect 1806 838 1807 842
rect 1811 838 1812 842
rect 1806 837 1812 838
rect 1910 842 1916 843
rect 1910 838 1911 842
rect 1915 838 1916 842
rect 1910 837 1916 838
rect 2014 842 2020 843
rect 2014 838 2015 842
rect 2019 838 2020 842
rect 2014 837 2020 838
rect 2118 842 2124 843
rect 2118 838 2119 842
rect 2123 838 2124 842
rect 2118 837 2124 838
rect 2222 842 2228 843
rect 2222 838 2223 842
rect 2227 838 2228 842
rect 2222 837 2228 838
rect 2326 842 2332 843
rect 2326 838 2327 842
rect 2331 838 2332 842
rect 2326 837 2332 838
rect 2438 842 2444 843
rect 2438 838 2439 842
rect 2443 838 2444 842
rect 2438 837 2444 838
rect 2542 842 2548 843
rect 2542 838 2543 842
rect 2547 838 2548 842
rect 2542 837 2548 838
rect 1416 827 1418 837
rect 1472 827 1474 837
rect 1536 827 1538 837
rect 1624 827 1626 837
rect 1712 827 1714 837
rect 1808 827 1810 837
rect 1912 827 1914 837
rect 2016 827 2018 837
rect 2120 827 2122 837
rect 2224 827 2226 837
rect 2328 827 2330 837
rect 2440 827 2442 837
rect 2544 827 2546 837
rect 2584 827 2586 846
rect 1367 826 1371 827
rect 111 822 115 823
rect 111 817 115 818
rect 199 822 203 823
rect 199 817 203 818
rect 255 822 259 823
rect 255 817 259 818
rect 319 822 323 823
rect 319 817 323 818
rect 383 822 387 823
rect 383 817 387 818
rect 391 822 395 823
rect 391 817 395 818
rect 439 822 443 823
rect 439 817 443 818
rect 471 822 475 823
rect 471 817 475 818
rect 495 822 499 823
rect 495 817 499 818
rect 559 822 563 823
rect 559 817 563 818
rect 631 822 635 823
rect 631 817 635 818
rect 655 822 659 823
rect 655 817 659 818
rect 703 822 707 823
rect 703 817 707 818
rect 759 822 763 823
rect 759 817 763 818
rect 783 822 787 823
rect 783 817 787 818
rect 871 822 875 823
rect 871 817 875 818
rect 959 822 963 823
rect 959 817 963 818
rect 983 822 987 823
rect 983 817 987 818
rect 1047 822 1051 823
rect 1047 817 1051 818
rect 1103 822 1107 823
rect 1103 817 1107 818
rect 1135 822 1139 823
rect 1135 817 1139 818
rect 1223 822 1227 823
rect 1223 817 1227 818
rect 1231 822 1235 823
rect 1231 817 1235 818
rect 1327 822 1331 823
rect 1367 821 1371 822
rect 1415 826 1419 827
rect 1415 821 1419 822
rect 1471 826 1475 827
rect 1471 821 1475 822
rect 1527 826 1531 827
rect 1527 821 1531 822
rect 1535 826 1539 827
rect 1535 821 1539 822
rect 1583 826 1587 827
rect 1583 821 1587 822
rect 1623 826 1627 827
rect 1623 821 1627 822
rect 1639 826 1643 827
rect 1639 821 1643 822
rect 1695 826 1699 827
rect 1695 821 1699 822
rect 1711 826 1715 827
rect 1711 821 1715 822
rect 1751 826 1755 827
rect 1751 821 1755 822
rect 1807 826 1811 827
rect 1807 821 1811 822
rect 1879 826 1883 827
rect 1879 821 1883 822
rect 1911 826 1915 827
rect 1911 821 1915 822
rect 1959 826 1963 827
rect 1959 821 1963 822
rect 2015 826 2019 827
rect 2015 821 2019 822
rect 2055 826 2059 827
rect 2055 821 2059 822
rect 2119 826 2123 827
rect 2119 821 2123 822
rect 2167 826 2171 827
rect 2167 821 2171 822
rect 2223 826 2227 827
rect 2223 821 2227 822
rect 2295 826 2299 827
rect 2295 821 2299 822
rect 2327 826 2331 827
rect 2327 821 2331 822
rect 2431 826 2435 827
rect 2431 821 2435 822
rect 2439 826 2443 827
rect 2439 821 2443 822
rect 2543 826 2547 827
rect 2543 821 2547 822
rect 2583 826 2587 827
rect 2583 821 2587 822
rect 1327 817 1331 818
rect 112 802 114 817
rect 384 811 386 817
rect 440 811 442 817
rect 496 811 498 817
rect 560 811 562 817
rect 632 811 634 817
rect 704 811 706 817
rect 784 811 786 817
rect 872 811 874 817
rect 960 811 962 817
rect 1048 811 1050 817
rect 1136 811 1138 817
rect 1224 811 1226 817
rect 382 810 388 811
rect 382 806 383 810
rect 387 806 388 810
rect 382 805 388 806
rect 438 810 444 811
rect 438 806 439 810
rect 443 806 444 810
rect 438 805 444 806
rect 494 810 500 811
rect 494 806 495 810
rect 499 806 500 810
rect 494 805 500 806
rect 558 810 564 811
rect 558 806 559 810
rect 563 806 564 810
rect 558 805 564 806
rect 630 810 636 811
rect 630 806 631 810
rect 635 806 636 810
rect 630 805 636 806
rect 702 810 708 811
rect 702 806 703 810
rect 707 806 708 810
rect 702 805 708 806
rect 782 810 788 811
rect 782 806 783 810
rect 787 806 788 810
rect 782 805 788 806
rect 870 810 876 811
rect 870 806 871 810
rect 875 806 876 810
rect 870 805 876 806
rect 958 810 964 811
rect 958 806 959 810
rect 963 806 964 810
rect 958 805 964 806
rect 1046 810 1052 811
rect 1046 806 1047 810
rect 1051 806 1052 810
rect 1046 805 1052 806
rect 1134 810 1140 811
rect 1134 806 1135 810
rect 1139 806 1140 810
rect 1134 805 1140 806
rect 1222 810 1228 811
rect 1222 806 1223 810
rect 1227 806 1228 810
rect 1222 805 1228 806
rect 1328 802 1330 817
rect 1368 806 1370 821
rect 1528 815 1530 821
rect 1584 815 1586 821
rect 1640 815 1642 821
rect 1696 815 1698 821
rect 1752 815 1754 821
rect 1808 815 1810 821
rect 1880 815 1882 821
rect 1960 815 1962 821
rect 2056 815 2058 821
rect 2168 815 2170 821
rect 2296 815 2298 821
rect 2432 815 2434 821
rect 2544 815 2546 821
rect 1526 814 1532 815
rect 1526 810 1527 814
rect 1531 810 1532 814
rect 1526 809 1532 810
rect 1582 814 1588 815
rect 1582 810 1583 814
rect 1587 810 1588 814
rect 1582 809 1588 810
rect 1638 814 1644 815
rect 1638 810 1639 814
rect 1643 810 1644 814
rect 1638 809 1644 810
rect 1694 814 1700 815
rect 1694 810 1695 814
rect 1699 810 1700 814
rect 1694 809 1700 810
rect 1750 814 1756 815
rect 1750 810 1751 814
rect 1755 810 1756 814
rect 1750 809 1756 810
rect 1806 814 1812 815
rect 1806 810 1807 814
rect 1811 810 1812 814
rect 1806 809 1812 810
rect 1878 814 1884 815
rect 1878 810 1879 814
rect 1883 810 1884 814
rect 1878 809 1884 810
rect 1958 814 1964 815
rect 1958 810 1959 814
rect 1963 810 1964 814
rect 1958 809 1964 810
rect 2054 814 2060 815
rect 2054 810 2055 814
rect 2059 810 2060 814
rect 2054 809 2060 810
rect 2166 814 2172 815
rect 2166 810 2167 814
rect 2171 810 2172 814
rect 2166 809 2172 810
rect 2294 814 2300 815
rect 2294 810 2295 814
rect 2299 810 2300 814
rect 2294 809 2300 810
rect 2430 814 2436 815
rect 2430 810 2431 814
rect 2435 810 2436 814
rect 2430 809 2436 810
rect 2542 814 2548 815
rect 2542 810 2543 814
rect 2547 810 2548 814
rect 2542 809 2548 810
rect 2584 806 2586 821
rect 1366 805 1372 806
rect 110 801 116 802
rect 110 797 111 801
rect 115 797 116 801
rect 110 796 116 797
rect 1326 801 1332 802
rect 1326 797 1327 801
rect 1331 797 1332 801
rect 1366 801 1367 805
rect 1371 801 1372 805
rect 1366 800 1372 801
rect 2582 805 2588 806
rect 2582 801 2583 805
rect 2587 801 2588 805
rect 2582 800 2588 801
rect 1326 796 1332 797
rect 1366 788 1372 789
rect 2582 788 2588 789
rect 110 784 116 785
rect 1326 784 1332 785
rect 110 780 111 784
rect 115 780 116 784
rect 110 779 116 780
rect 366 783 372 784
rect 366 779 367 783
rect 371 779 372 783
rect 112 767 114 779
rect 366 778 372 779
rect 422 783 428 784
rect 422 779 423 783
rect 427 779 428 783
rect 422 778 428 779
rect 478 783 484 784
rect 478 779 479 783
rect 483 779 484 783
rect 478 778 484 779
rect 542 783 548 784
rect 542 779 543 783
rect 547 779 548 783
rect 542 778 548 779
rect 614 783 620 784
rect 614 779 615 783
rect 619 779 620 783
rect 614 778 620 779
rect 686 783 692 784
rect 686 779 687 783
rect 691 779 692 783
rect 686 778 692 779
rect 766 783 772 784
rect 766 779 767 783
rect 771 779 772 783
rect 766 778 772 779
rect 854 783 860 784
rect 854 779 855 783
rect 859 779 860 783
rect 854 778 860 779
rect 942 783 948 784
rect 942 779 943 783
rect 947 779 948 783
rect 942 778 948 779
rect 1030 783 1036 784
rect 1030 779 1031 783
rect 1035 779 1036 783
rect 1030 778 1036 779
rect 1118 783 1124 784
rect 1118 779 1119 783
rect 1123 779 1124 783
rect 1118 778 1124 779
rect 1206 783 1212 784
rect 1206 779 1207 783
rect 1211 779 1212 783
rect 1326 780 1327 784
rect 1331 780 1332 784
rect 1366 784 1367 788
rect 1371 784 1372 788
rect 1366 783 1372 784
rect 1510 787 1516 788
rect 1510 783 1511 787
rect 1515 783 1516 787
rect 1326 779 1332 780
rect 1206 778 1212 779
rect 368 767 370 778
rect 424 767 426 778
rect 480 767 482 778
rect 544 767 546 778
rect 616 767 618 778
rect 688 767 690 778
rect 768 767 770 778
rect 856 767 858 778
rect 944 767 946 778
rect 1032 767 1034 778
rect 1120 767 1122 778
rect 1208 767 1210 778
rect 1328 767 1330 779
rect 111 766 115 767
rect 111 761 115 762
rect 367 766 371 767
rect 367 761 371 762
rect 383 766 387 767
rect 383 761 387 762
rect 423 766 427 767
rect 423 761 427 762
rect 439 766 443 767
rect 439 761 443 762
rect 479 766 483 767
rect 479 761 483 762
rect 495 766 499 767
rect 495 761 499 762
rect 543 766 547 767
rect 543 761 547 762
rect 559 766 563 767
rect 559 761 563 762
rect 615 766 619 767
rect 615 761 619 762
rect 631 766 635 767
rect 631 761 635 762
rect 687 766 691 767
rect 687 761 691 762
rect 711 766 715 767
rect 711 761 715 762
rect 767 766 771 767
rect 767 761 771 762
rect 791 766 795 767
rect 791 761 795 762
rect 855 766 859 767
rect 855 761 859 762
rect 871 766 875 767
rect 871 761 875 762
rect 943 766 947 767
rect 943 761 947 762
rect 951 766 955 767
rect 951 761 955 762
rect 1031 766 1035 767
rect 1031 761 1035 762
rect 1039 766 1043 767
rect 1039 761 1043 762
rect 1119 766 1123 767
rect 1119 761 1123 762
rect 1127 766 1131 767
rect 1127 761 1131 762
rect 1207 766 1211 767
rect 1207 761 1211 762
rect 1327 766 1331 767
rect 1368 763 1370 783
rect 1510 782 1516 783
rect 1566 787 1572 788
rect 1566 783 1567 787
rect 1571 783 1572 787
rect 1566 782 1572 783
rect 1622 787 1628 788
rect 1622 783 1623 787
rect 1627 783 1628 787
rect 1622 782 1628 783
rect 1678 787 1684 788
rect 1678 783 1679 787
rect 1683 783 1684 787
rect 1678 782 1684 783
rect 1734 787 1740 788
rect 1734 783 1735 787
rect 1739 783 1740 787
rect 1734 782 1740 783
rect 1790 787 1796 788
rect 1790 783 1791 787
rect 1795 783 1796 787
rect 1790 782 1796 783
rect 1862 787 1868 788
rect 1862 783 1863 787
rect 1867 783 1868 787
rect 1862 782 1868 783
rect 1942 787 1948 788
rect 1942 783 1943 787
rect 1947 783 1948 787
rect 1942 782 1948 783
rect 2038 787 2044 788
rect 2038 783 2039 787
rect 2043 783 2044 787
rect 2038 782 2044 783
rect 2150 787 2156 788
rect 2150 783 2151 787
rect 2155 783 2156 787
rect 2150 782 2156 783
rect 2278 787 2284 788
rect 2278 783 2279 787
rect 2283 783 2284 787
rect 2278 782 2284 783
rect 2414 787 2420 788
rect 2414 783 2415 787
rect 2419 783 2420 787
rect 2414 782 2420 783
rect 2526 787 2532 788
rect 2526 783 2527 787
rect 2531 783 2532 787
rect 2582 784 2583 788
rect 2587 784 2588 788
rect 2582 783 2588 784
rect 2526 782 2532 783
rect 1512 763 1514 782
rect 1568 763 1570 782
rect 1624 763 1626 782
rect 1680 763 1682 782
rect 1736 763 1738 782
rect 1792 763 1794 782
rect 1864 763 1866 782
rect 1944 763 1946 782
rect 2040 763 2042 782
rect 2152 763 2154 782
rect 2280 763 2282 782
rect 2416 763 2418 782
rect 2528 763 2530 782
rect 2584 763 2586 783
rect 1327 761 1331 762
rect 1367 762 1371 763
rect 112 749 114 761
rect 384 750 386 761
rect 440 750 442 761
rect 496 750 498 761
rect 560 750 562 761
rect 632 750 634 761
rect 712 750 714 761
rect 792 750 794 761
rect 872 750 874 761
rect 952 750 954 761
rect 1040 750 1042 761
rect 1128 750 1130 761
rect 382 749 388 750
rect 110 748 116 749
rect 110 744 111 748
rect 115 744 116 748
rect 382 745 383 749
rect 387 745 388 749
rect 382 744 388 745
rect 438 749 444 750
rect 438 745 439 749
rect 443 745 444 749
rect 438 744 444 745
rect 494 749 500 750
rect 494 745 495 749
rect 499 745 500 749
rect 494 744 500 745
rect 558 749 564 750
rect 558 745 559 749
rect 563 745 564 749
rect 558 744 564 745
rect 630 749 636 750
rect 630 745 631 749
rect 635 745 636 749
rect 630 744 636 745
rect 710 749 716 750
rect 710 745 711 749
rect 715 745 716 749
rect 710 744 716 745
rect 790 749 796 750
rect 790 745 791 749
rect 795 745 796 749
rect 790 744 796 745
rect 870 749 876 750
rect 870 745 871 749
rect 875 745 876 749
rect 870 744 876 745
rect 950 749 956 750
rect 950 745 951 749
rect 955 745 956 749
rect 950 744 956 745
rect 1038 749 1044 750
rect 1038 745 1039 749
rect 1043 745 1044 749
rect 1038 744 1044 745
rect 1126 749 1132 750
rect 1328 749 1330 761
rect 1367 757 1371 758
rect 1511 762 1515 763
rect 1511 757 1515 758
rect 1567 762 1571 763
rect 1567 757 1571 758
rect 1623 762 1627 763
rect 1623 757 1627 758
rect 1647 762 1651 763
rect 1647 757 1651 758
rect 1679 762 1683 763
rect 1679 757 1683 758
rect 1703 762 1707 763
rect 1703 757 1707 758
rect 1735 762 1739 763
rect 1735 757 1739 758
rect 1759 762 1763 763
rect 1759 757 1763 758
rect 1791 762 1795 763
rect 1791 757 1795 758
rect 1815 762 1819 763
rect 1815 757 1819 758
rect 1863 762 1867 763
rect 1863 757 1867 758
rect 1871 762 1875 763
rect 1871 757 1875 758
rect 1927 762 1931 763
rect 1927 757 1931 758
rect 1943 762 1947 763
rect 1943 757 1947 758
rect 1991 762 1995 763
rect 1991 757 1995 758
rect 2039 762 2043 763
rect 2039 757 2043 758
rect 2063 762 2067 763
rect 2063 757 2067 758
rect 2143 762 2147 763
rect 2143 757 2147 758
rect 2151 762 2155 763
rect 2151 757 2155 758
rect 2231 762 2235 763
rect 2231 757 2235 758
rect 2279 762 2283 763
rect 2279 757 2283 758
rect 2335 762 2339 763
rect 2335 757 2339 758
rect 2415 762 2419 763
rect 2415 757 2419 758
rect 2439 762 2443 763
rect 2439 757 2443 758
rect 2527 762 2531 763
rect 2527 757 2531 758
rect 2583 762 2587 763
rect 2583 757 2587 758
rect 1126 745 1127 749
rect 1131 745 1132 749
rect 1126 744 1132 745
rect 1326 748 1332 749
rect 1326 744 1327 748
rect 1331 744 1332 748
rect 1368 745 1370 757
rect 1648 746 1650 757
rect 1704 746 1706 757
rect 1760 746 1762 757
rect 1816 746 1818 757
rect 1872 746 1874 757
rect 1928 746 1930 757
rect 1992 746 1994 757
rect 2064 746 2066 757
rect 2144 746 2146 757
rect 2232 746 2234 757
rect 2336 746 2338 757
rect 2440 746 2442 757
rect 2528 746 2530 757
rect 1646 745 1652 746
rect 110 743 116 744
rect 1326 743 1332 744
rect 1366 744 1372 745
rect 1366 740 1367 744
rect 1371 740 1372 744
rect 1646 741 1647 745
rect 1651 741 1652 745
rect 1646 740 1652 741
rect 1702 745 1708 746
rect 1702 741 1703 745
rect 1707 741 1708 745
rect 1702 740 1708 741
rect 1758 745 1764 746
rect 1758 741 1759 745
rect 1763 741 1764 745
rect 1758 740 1764 741
rect 1814 745 1820 746
rect 1814 741 1815 745
rect 1819 741 1820 745
rect 1814 740 1820 741
rect 1870 745 1876 746
rect 1870 741 1871 745
rect 1875 741 1876 745
rect 1870 740 1876 741
rect 1926 745 1932 746
rect 1926 741 1927 745
rect 1931 741 1932 745
rect 1926 740 1932 741
rect 1990 745 1996 746
rect 1990 741 1991 745
rect 1995 741 1996 745
rect 1990 740 1996 741
rect 2062 745 2068 746
rect 2062 741 2063 745
rect 2067 741 2068 745
rect 2062 740 2068 741
rect 2142 745 2148 746
rect 2142 741 2143 745
rect 2147 741 2148 745
rect 2142 740 2148 741
rect 2230 745 2236 746
rect 2230 741 2231 745
rect 2235 741 2236 745
rect 2230 740 2236 741
rect 2334 745 2340 746
rect 2334 741 2335 745
rect 2339 741 2340 745
rect 2334 740 2340 741
rect 2438 745 2444 746
rect 2438 741 2439 745
rect 2443 741 2444 745
rect 2438 740 2444 741
rect 2526 745 2532 746
rect 2584 745 2586 757
rect 2526 741 2527 745
rect 2531 741 2532 745
rect 2526 740 2532 741
rect 2582 744 2588 745
rect 2582 740 2583 744
rect 2587 740 2588 744
rect 1366 739 1372 740
rect 2582 739 2588 740
rect 110 731 116 732
rect 110 727 111 731
rect 115 727 116 731
rect 110 726 116 727
rect 1326 731 1332 732
rect 1326 727 1327 731
rect 1331 727 1332 731
rect 1326 726 1332 727
rect 1366 727 1372 728
rect 112 711 114 726
rect 398 722 404 723
rect 398 718 399 722
rect 403 718 404 722
rect 398 717 404 718
rect 454 722 460 723
rect 454 718 455 722
rect 459 718 460 722
rect 454 717 460 718
rect 510 722 516 723
rect 510 718 511 722
rect 515 718 516 722
rect 510 717 516 718
rect 574 722 580 723
rect 574 718 575 722
rect 579 718 580 722
rect 574 717 580 718
rect 646 722 652 723
rect 646 718 647 722
rect 651 718 652 722
rect 646 717 652 718
rect 726 722 732 723
rect 726 718 727 722
rect 731 718 732 722
rect 726 717 732 718
rect 806 722 812 723
rect 806 718 807 722
rect 811 718 812 722
rect 806 717 812 718
rect 886 722 892 723
rect 886 718 887 722
rect 891 718 892 722
rect 886 717 892 718
rect 966 722 972 723
rect 966 718 967 722
rect 971 718 972 722
rect 966 717 972 718
rect 1054 722 1060 723
rect 1054 718 1055 722
rect 1059 718 1060 722
rect 1054 717 1060 718
rect 1142 722 1148 723
rect 1142 718 1143 722
rect 1147 718 1148 722
rect 1142 717 1148 718
rect 400 711 402 717
rect 456 711 458 717
rect 512 711 514 717
rect 576 711 578 717
rect 648 711 650 717
rect 728 711 730 717
rect 808 711 810 717
rect 888 711 890 717
rect 968 711 970 717
rect 1056 711 1058 717
rect 1144 711 1146 717
rect 1328 711 1330 726
rect 1366 723 1367 727
rect 1371 723 1372 727
rect 1366 722 1372 723
rect 2582 727 2588 728
rect 2582 723 2583 727
rect 2587 723 2588 727
rect 2582 722 2588 723
rect 111 710 115 711
rect 111 705 115 706
rect 343 710 347 711
rect 343 705 347 706
rect 399 710 403 711
rect 399 705 403 706
rect 415 710 419 711
rect 415 705 419 706
rect 455 710 459 711
rect 455 705 459 706
rect 487 710 491 711
rect 487 705 491 706
rect 511 710 515 711
rect 511 705 515 706
rect 559 710 563 711
rect 559 705 563 706
rect 575 710 579 711
rect 575 705 579 706
rect 631 710 635 711
rect 631 705 635 706
rect 647 710 651 711
rect 647 705 651 706
rect 695 710 699 711
rect 695 705 699 706
rect 727 710 731 711
rect 727 705 731 706
rect 759 710 763 711
rect 759 705 763 706
rect 807 710 811 711
rect 807 705 811 706
rect 823 710 827 711
rect 823 705 827 706
rect 887 710 891 711
rect 887 705 891 706
rect 951 710 955 711
rect 951 705 955 706
rect 967 710 971 711
rect 967 705 971 706
rect 1023 710 1027 711
rect 1023 705 1027 706
rect 1055 710 1059 711
rect 1055 705 1059 706
rect 1143 710 1147 711
rect 1143 705 1147 706
rect 1327 710 1331 711
rect 1327 705 1331 706
rect 112 690 114 705
rect 344 699 346 705
rect 416 699 418 705
rect 488 699 490 705
rect 560 699 562 705
rect 632 699 634 705
rect 696 699 698 705
rect 760 699 762 705
rect 824 699 826 705
rect 888 699 890 705
rect 952 699 954 705
rect 1024 699 1026 705
rect 342 698 348 699
rect 342 694 343 698
rect 347 694 348 698
rect 342 693 348 694
rect 414 698 420 699
rect 414 694 415 698
rect 419 694 420 698
rect 414 693 420 694
rect 486 698 492 699
rect 486 694 487 698
rect 491 694 492 698
rect 486 693 492 694
rect 558 698 564 699
rect 558 694 559 698
rect 563 694 564 698
rect 558 693 564 694
rect 630 698 636 699
rect 630 694 631 698
rect 635 694 636 698
rect 630 693 636 694
rect 694 698 700 699
rect 694 694 695 698
rect 699 694 700 698
rect 694 693 700 694
rect 758 698 764 699
rect 758 694 759 698
rect 763 694 764 698
rect 758 693 764 694
rect 822 698 828 699
rect 822 694 823 698
rect 827 694 828 698
rect 822 693 828 694
rect 886 698 892 699
rect 886 694 887 698
rect 891 694 892 698
rect 886 693 892 694
rect 950 698 956 699
rect 950 694 951 698
rect 955 694 956 698
rect 950 693 956 694
rect 1022 698 1028 699
rect 1022 694 1023 698
rect 1027 694 1028 698
rect 1022 693 1028 694
rect 1328 690 1330 705
rect 1368 703 1370 722
rect 1662 718 1668 719
rect 1662 714 1663 718
rect 1667 714 1668 718
rect 1662 713 1668 714
rect 1718 718 1724 719
rect 1718 714 1719 718
rect 1723 714 1724 718
rect 1718 713 1724 714
rect 1774 718 1780 719
rect 1774 714 1775 718
rect 1779 714 1780 718
rect 1774 713 1780 714
rect 1830 718 1836 719
rect 1830 714 1831 718
rect 1835 714 1836 718
rect 1830 713 1836 714
rect 1886 718 1892 719
rect 1886 714 1887 718
rect 1891 714 1892 718
rect 1886 713 1892 714
rect 1942 718 1948 719
rect 1942 714 1943 718
rect 1947 714 1948 718
rect 1942 713 1948 714
rect 2006 718 2012 719
rect 2006 714 2007 718
rect 2011 714 2012 718
rect 2006 713 2012 714
rect 2078 718 2084 719
rect 2078 714 2079 718
rect 2083 714 2084 718
rect 2078 713 2084 714
rect 2158 718 2164 719
rect 2158 714 2159 718
rect 2163 714 2164 718
rect 2158 713 2164 714
rect 2246 718 2252 719
rect 2246 714 2247 718
rect 2251 714 2252 718
rect 2246 713 2252 714
rect 2350 718 2356 719
rect 2350 714 2351 718
rect 2355 714 2356 718
rect 2350 713 2356 714
rect 2454 718 2460 719
rect 2454 714 2455 718
rect 2459 714 2460 718
rect 2454 713 2460 714
rect 2542 718 2548 719
rect 2542 714 2543 718
rect 2547 714 2548 718
rect 2542 713 2548 714
rect 1664 703 1666 713
rect 1720 703 1722 713
rect 1776 703 1778 713
rect 1832 703 1834 713
rect 1888 703 1890 713
rect 1944 703 1946 713
rect 2008 703 2010 713
rect 2080 703 2082 713
rect 2160 703 2162 713
rect 2248 703 2250 713
rect 2352 703 2354 713
rect 2456 703 2458 713
rect 2544 703 2546 713
rect 2584 703 2586 722
rect 1367 702 1371 703
rect 1367 697 1371 698
rect 1663 702 1667 703
rect 1663 697 1667 698
rect 1719 702 1723 703
rect 1719 697 1723 698
rect 1735 702 1739 703
rect 1735 697 1739 698
rect 1775 702 1779 703
rect 1775 697 1779 698
rect 1791 702 1795 703
rect 1791 697 1795 698
rect 1831 702 1835 703
rect 1831 697 1835 698
rect 1855 702 1859 703
rect 1855 697 1859 698
rect 1887 702 1891 703
rect 1887 697 1891 698
rect 1919 702 1923 703
rect 1919 697 1923 698
rect 1943 702 1947 703
rect 1943 697 1947 698
rect 1991 702 1995 703
rect 1991 697 1995 698
rect 2007 702 2011 703
rect 2007 697 2011 698
rect 2063 702 2067 703
rect 2063 697 2067 698
rect 2079 702 2083 703
rect 2079 697 2083 698
rect 2127 702 2131 703
rect 2127 697 2131 698
rect 2159 702 2163 703
rect 2159 697 2163 698
rect 2199 702 2203 703
rect 2199 697 2203 698
rect 2247 702 2251 703
rect 2247 697 2251 698
rect 2271 702 2275 703
rect 2271 697 2275 698
rect 2343 702 2347 703
rect 2343 697 2347 698
rect 2351 702 2355 703
rect 2351 697 2355 698
rect 2415 702 2419 703
rect 2415 697 2419 698
rect 2455 702 2459 703
rect 2455 697 2459 698
rect 2487 702 2491 703
rect 2487 697 2491 698
rect 2543 702 2547 703
rect 2543 697 2547 698
rect 2583 702 2587 703
rect 2583 697 2587 698
rect 110 689 116 690
rect 110 685 111 689
rect 115 685 116 689
rect 110 684 116 685
rect 1326 689 1332 690
rect 1326 685 1327 689
rect 1331 685 1332 689
rect 1326 684 1332 685
rect 1368 682 1370 697
rect 1736 691 1738 697
rect 1792 691 1794 697
rect 1856 691 1858 697
rect 1920 691 1922 697
rect 1992 691 1994 697
rect 2064 691 2066 697
rect 2128 691 2130 697
rect 2200 691 2202 697
rect 2272 691 2274 697
rect 2344 691 2346 697
rect 2416 691 2418 697
rect 2488 691 2490 697
rect 2544 691 2546 697
rect 1734 690 1740 691
rect 1734 686 1735 690
rect 1739 686 1740 690
rect 1734 685 1740 686
rect 1790 690 1796 691
rect 1790 686 1791 690
rect 1795 686 1796 690
rect 1790 685 1796 686
rect 1854 690 1860 691
rect 1854 686 1855 690
rect 1859 686 1860 690
rect 1854 685 1860 686
rect 1918 690 1924 691
rect 1918 686 1919 690
rect 1923 686 1924 690
rect 1918 685 1924 686
rect 1990 690 1996 691
rect 1990 686 1991 690
rect 1995 686 1996 690
rect 1990 685 1996 686
rect 2062 690 2068 691
rect 2062 686 2063 690
rect 2067 686 2068 690
rect 2062 685 2068 686
rect 2126 690 2132 691
rect 2126 686 2127 690
rect 2131 686 2132 690
rect 2126 685 2132 686
rect 2198 690 2204 691
rect 2198 686 2199 690
rect 2203 686 2204 690
rect 2198 685 2204 686
rect 2270 690 2276 691
rect 2270 686 2271 690
rect 2275 686 2276 690
rect 2270 685 2276 686
rect 2342 690 2348 691
rect 2342 686 2343 690
rect 2347 686 2348 690
rect 2342 685 2348 686
rect 2414 690 2420 691
rect 2414 686 2415 690
rect 2419 686 2420 690
rect 2414 685 2420 686
rect 2486 690 2492 691
rect 2486 686 2487 690
rect 2491 686 2492 690
rect 2486 685 2492 686
rect 2542 690 2548 691
rect 2542 686 2543 690
rect 2547 686 2548 690
rect 2542 685 2548 686
rect 2584 682 2586 697
rect 1366 681 1372 682
rect 1366 677 1367 681
rect 1371 677 1372 681
rect 1366 676 1372 677
rect 2582 681 2588 682
rect 2582 677 2583 681
rect 2587 677 2588 681
rect 2582 676 2588 677
rect 110 672 116 673
rect 1326 672 1332 673
rect 110 668 111 672
rect 115 668 116 672
rect 110 667 116 668
rect 326 671 332 672
rect 326 667 327 671
rect 331 667 332 671
rect 112 651 114 667
rect 326 666 332 667
rect 398 671 404 672
rect 398 667 399 671
rect 403 667 404 671
rect 398 666 404 667
rect 470 671 476 672
rect 470 667 471 671
rect 475 667 476 671
rect 470 666 476 667
rect 542 671 548 672
rect 542 667 543 671
rect 547 667 548 671
rect 542 666 548 667
rect 614 671 620 672
rect 614 667 615 671
rect 619 667 620 671
rect 614 666 620 667
rect 678 671 684 672
rect 678 667 679 671
rect 683 667 684 671
rect 678 666 684 667
rect 742 671 748 672
rect 742 667 743 671
rect 747 667 748 671
rect 742 666 748 667
rect 806 671 812 672
rect 806 667 807 671
rect 811 667 812 671
rect 806 666 812 667
rect 870 671 876 672
rect 870 667 871 671
rect 875 667 876 671
rect 870 666 876 667
rect 934 671 940 672
rect 934 667 935 671
rect 939 667 940 671
rect 934 666 940 667
rect 1006 671 1012 672
rect 1006 667 1007 671
rect 1011 667 1012 671
rect 1326 668 1327 672
rect 1331 668 1332 672
rect 1326 667 1332 668
rect 1006 666 1012 667
rect 328 651 330 666
rect 400 651 402 666
rect 472 651 474 666
rect 544 651 546 666
rect 616 651 618 666
rect 680 651 682 666
rect 744 651 746 666
rect 808 651 810 666
rect 872 651 874 666
rect 936 651 938 666
rect 1008 651 1010 666
rect 1328 651 1330 667
rect 1366 664 1372 665
rect 2582 664 2588 665
rect 1366 660 1367 664
rect 1371 660 1372 664
rect 1366 659 1372 660
rect 1718 663 1724 664
rect 1718 659 1719 663
rect 1723 659 1724 663
rect 111 650 115 651
rect 111 645 115 646
rect 231 650 235 651
rect 231 645 235 646
rect 295 650 299 651
rect 295 645 299 646
rect 327 650 331 651
rect 327 645 331 646
rect 359 650 363 651
rect 359 645 363 646
rect 399 650 403 651
rect 399 645 403 646
rect 423 650 427 651
rect 423 645 427 646
rect 471 650 475 651
rect 471 645 475 646
rect 479 650 483 651
rect 479 645 483 646
rect 535 650 539 651
rect 535 645 539 646
rect 543 650 547 651
rect 543 645 547 646
rect 599 650 603 651
rect 599 645 603 646
rect 615 650 619 651
rect 615 645 619 646
rect 663 650 667 651
rect 663 645 667 646
rect 679 650 683 651
rect 679 645 683 646
rect 727 650 731 651
rect 727 645 731 646
rect 743 650 747 651
rect 743 645 747 646
rect 791 650 795 651
rect 791 645 795 646
rect 807 650 811 651
rect 807 645 811 646
rect 855 650 859 651
rect 855 645 859 646
rect 871 650 875 651
rect 871 645 875 646
rect 919 650 923 651
rect 919 645 923 646
rect 935 650 939 651
rect 935 645 939 646
rect 1007 650 1011 651
rect 1007 645 1011 646
rect 1327 650 1331 651
rect 1327 645 1331 646
rect 112 633 114 645
rect 232 634 234 645
rect 296 634 298 645
rect 360 634 362 645
rect 424 634 426 645
rect 480 634 482 645
rect 536 634 538 645
rect 600 634 602 645
rect 664 634 666 645
rect 728 634 730 645
rect 792 634 794 645
rect 856 634 858 645
rect 920 634 922 645
rect 230 633 236 634
rect 110 632 116 633
rect 110 628 111 632
rect 115 628 116 632
rect 230 629 231 633
rect 235 629 236 633
rect 230 628 236 629
rect 294 633 300 634
rect 294 629 295 633
rect 299 629 300 633
rect 294 628 300 629
rect 358 633 364 634
rect 358 629 359 633
rect 363 629 364 633
rect 358 628 364 629
rect 422 633 428 634
rect 422 629 423 633
rect 427 629 428 633
rect 422 628 428 629
rect 478 633 484 634
rect 478 629 479 633
rect 483 629 484 633
rect 478 628 484 629
rect 534 633 540 634
rect 534 629 535 633
rect 539 629 540 633
rect 534 628 540 629
rect 598 633 604 634
rect 598 629 599 633
rect 603 629 604 633
rect 598 628 604 629
rect 662 633 668 634
rect 662 629 663 633
rect 667 629 668 633
rect 662 628 668 629
rect 726 633 732 634
rect 726 629 727 633
rect 731 629 732 633
rect 726 628 732 629
rect 790 633 796 634
rect 790 629 791 633
rect 795 629 796 633
rect 790 628 796 629
rect 854 633 860 634
rect 854 629 855 633
rect 859 629 860 633
rect 854 628 860 629
rect 918 633 924 634
rect 1328 633 1330 645
rect 1368 643 1370 659
rect 1718 658 1724 659
rect 1774 663 1780 664
rect 1774 659 1775 663
rect 1779 659 1780 663
rect 1774 658 1780 659
rect 1838 663 1844 664
rect 1838 659 1839 663
rect 1843 659 1844 663
rect 1838 658 1844 659
rect 1902 663 1908 664
rect 1902 659 1903 663
rect 1907 659 1908 663
rect 1902 658 1908 659
rect 1974 663 1980 664
rect 1974 659 1975 663
rect 1979 659 1980 663
rect 1974 658 1980 659
rect 2046 663 2052 664
rect 2046 659 2047 663
rect 2051 659 2052 663
rect 2046 658 2052 659
rect 2110 663 2116 664
rect 2110 659 2111 663
rect 2115 659 2116 663
rect 2110 658 2116 659
rect 2182 663 2188 664
rect 2182 659 2183 663
rect 2187 659 2188 663
rect 2182 658 2188 659
rect 2254 663 2260 664
rect 2254 659 2255 663
rect 2259 659 2260 663
rect 2254 658 2260 659
rect 2326 663 2332 664
rect 2326 659 2327 663
rect 2331 659 2332 663
rect 2326 658 2332 659
rect 2398 663 2404 664
rect 2398 659 2399 663
rect 2403 659 2404 663
rect 2398 658 2404 659
rect 2470 663 2476 664
rect 2470 659 2471 663
rect 2475 659 2476 663
rect 2470 658 2476 659
rect 2526 663 2532 664
rect 2526 659 2527 663
rect 2531 659 2532 663
rect 2582 660 2583 664
rect 2587 660 2588 664
rect 2582 659 2588 660
rect 2526 658 2532 659
rect 1720 643 1722 658
rect 1776 643 1778 658
rect 1840 643 1842 658
rect 1904 643 1906 658
rect 1976 643 1978 658
rect 2048 643 2050 658
rect 2112 643 2114 658
rect 2184 643 2186 658
rect 2256 643 2258 658
rect 2328 643 2330 658
rect 2400 643 2402 658
rect 2472 643 2474 658
rect 2528 643 2530 658
rect 2584 643 2586 659
rect 1367 642 1371 643
rect 1367 637 1371 638
rect 1615 642 1619 643
rect 1615 637 1619 638
rect 1679 642 1683 643
rect 1679 637 1683 638
rect 1719 642 1723 643
rect 1719 637 1723 638
rect 1759 642 1763 643
rect 1759 637 1763 638
rect 1775 642 1779 643
rect 1775 637 1779 638
rect 1839 642 1843 643
rect 1839 637 1843 638
rect 1903 642 1907 643
rect 1903 637 1907 638
rect 1927 642 1931 643
rect 1927 637 1931 638
rect 1975 642 1979 643
rect 1975 637 1979 638
rect 2015 642 2019 643
rect 2015 637 2019 638
rect 2047 642 2051 643
rect 2047 637 2051 638
rect 2095 642 2099 643
rect 2095 637 2099 638
rect 2111 642 2115 643
rect 2111 637 2115 638
rect 2175 642 2179 643
rect 2175 637 2179 638
rect 2183 642 2187 643
rect 2183 637 2187 638
rect 2255 642 2259 643
rect 2255 637 2259 638
rect 2327 642 2331 643
rect 2327 637 2331 638
rect 2399 642 2403 643
rect 2399 637 2403 638
rect 2471 642 2475 643
rect 2471 637 2475 638
rect 2527 642 2531 643
rect 2527 637 2531 638
rect 2583 642 2587 643
rect 2583 637 2587 638
rect 918 629 919 633
rect 923 629 924 633
rect 918 628 924 629
rect 1326 632 1332 633
rect 1326 628 1327 632
rect 1331 628 1332 632
rect 110 627 116 628
rect 1326 627 1332 628
rect 1368 625 1370 637
rect 1616 626 1618 637
rect 1680 626 1682 637
rect 1760 626 1762 637
rect 1840 626 1842 637
rect 1928 626 1930 637
rect 2016 626 2018 637
rect 2096 626 2098 637
rect 2176 626 2178 637
rect 2256 626 2258 637
rect 2328 626 2330 637
rect 2400 626 2402 637
rect 2472 626 2474 637
rect 2528 626 2530 637
rect 1614 625 1620 626
rect 1366 624 1372 625
rect 1366 620 1367 624
rect 1371 620 1372 624
rect 1614 621 1615 625
rect 1619 621 1620 625
rect 1614 620 1620 621
rect 1678 625 1684 626
rect 1678 621 1679 625
rect 1683 621 1684 625
rect 1678 620 1684 621
rect 1758 625 1764 626
rect 1758 621 1759 625
rect 1763 621 1764 625
rect 1758 620 1764 621
rect 1838 625 1844 626
rect 1838 621 1839 625
rect 1843 621 1844 625
rect 1838 620 1844 621
rect 1926 625 1932 626
rect 1926 621 1927 625
rect 1931 621 1932 625
rect 1926 620 1932 621
rect 2014 625 2020 626
rect 2014 621 2015 625
rect 2019 621 2020 625
rect 2014 620 2020 621
rect 2094 625 2100 626
rect 2094 621 2095 625
rect 2099 621 2100 625
rect 2094 620 2100 621
rect 2174 625 2180 626
rect 2174 621 2175 625
rect 2179 621 2180 625
rect 2174 620 2180 621
rect 2254 625 2260 626
rect 2254 621 2255 625
rect 2259 621 2260 625
rect 2254 620 2260 621
rect 2326 625 2332 626
rect 2326 621 2327 625
rect 2331 621 2332 625
rect 2326 620 2332 621
rect 2398 625 2404 626
rect 2398 621 2399 625
rect 2403 621 2404 625
rect 2398 620 2404 621
rect 2470 625 2476 626
rect 2470 621 2471 625
rect 2475 621 2476 625
rect 2470 620 2476 621
rect 2526 625 2532 626
rect 2584 625 2586 637
rect 2526 621 2527 625
rect 2531 621 2532 625
rect 2526 620 2532 621
rect 2582 624 2588 625
rect 2582 620 2583 624
rect 2587 620 2588 624
rect 1366 619 1372 620
rect 2582 619 2588 620
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 110 610 116 611
rect 1326 615 1332 616
rect 1326 611 1327 615
rect 1331 611 1332 615
rect 1326 610 1332 611
rect 112 587 114 610
rect 246 606 252 607
rect 246 602 247 606
rect 251 602 252 606
rect 246 601 252 602
rect 310 606 316 607
rect 310 602 311 606
rect 315 602 316 606
rect 310 601 316 602
rect 374 606 380 607
rect 374 602 375 606
rect 379 602 380 606
rect 374 601 380 602
rect 438 606 444 607
rect 438 602 439 606
rect 443 602 444 606
rect 438 601 444 602
rect 494 606 500 607
rect 494 602 495 606
rect 499 602 500 606
rect 494 601 500 602
rect 550 606 556 607
rect 550 602 551 606
rect 555 602 556 606
rect 550 601 556 602
rect 614 606 620 607
rect 614 602 615 606
rect 619 602 620 606
rect 614 601 620 602
rect 678 606 684 607
rect 678 602 679 606
rect 683 602 684 606
rect 678 601 684 602
rect 742 606 748 607
rect 742 602 743 606
rect 747 602 748 606
rect 742 601 748 602
rect 806 606 812 607
rect 806 602 807 606
rect 811 602 812 606
rect 806 601 812 602
rect 870 606 876 607
rect 870 602 871 606
rect 875 602 876 606
rect 870 601 876 602
rect 934 606 940 607
rect 934 602 935 606
rect 939 602 940 606
rect 934 601 940 602
rect 248 587 250 601
rect 312 587 314 601
rect 376 587 378 601
rect 440 587 442 601
rect 496 587 498 601
rect 552 587 554 601
rect 616 587 618 601
rect 680 587 682 601
rect 744 587 746 601
rect 808 587 810 601
rect 872 587 874 601
rect 936 587 938 601
rect 1328 587 1330 610
rect 1366 607 1372 608
rect 1366 603 1367 607
rect 1371 603 1372 607
rect 1366 602 1372 603
rect 2582 607 2588 608
rect 2582 603 2583 607
rect 2587 603 2588 607
rect 2582 602 2588 603
rect 111 586 115 587
rect 111 581 115 582
rect 191 586 195 587
rect 191 581 195 582
rect 247 586 251 587
rect 247 581 251 582
rect 279 586 283 587
rect 279 581 283 582
rect 311 586 315 587
rect 311 581 315 582
rect 367 586 371 587
rect 367 581 371 582
rect 375 586 379 587
rect 375 581 379 582
rect 439 586 443 587
rect 439 581 443 582
rect 463 586 467 587
rect 463 581 467 582
rect 495 586 499 587
rect 495 581 499 582
rect 551 586 555 587
rect 551 581 555 582
rect 559 586 563 587
rect 559 581 563 582
rect 615 586 619 587
rect 615 581 619 582
rect 647 586 651 587
rect 647 581 651 582
rect 679 586 683 587
rect 679 581 683 582
rect 735 586 739 587
rect 735 581 739 582
rect 743 586 747 587
rect 743 581 747 582
rect 807 586 811 587
rect 807 581 811 582
rect 815 586 819 587
rect 815 581 819 582
rect 871 586 875 587
rect 871 581 875 582
rect 887 586 891 587
rect 887 581 891 582
rect 935 586 939 587
rect 935 581 939 582
rect 967 586 971 587
rect 967 581 971 582
rect 1047 586 1051 587
rect 1047 581 1051 582
rect 1127 586 1131 587
rect 1127 581 1131 582
rect 1327 586 1331 587
rect 1327 581 1331 582
rect 112 566 114 581
rect 192 575 194 581
rect 280 575 282 581
rect 368 575 370 581
rect 464 575 466 581
rect 560 575 562 581
rect 648 575 650 581
rect 736 575 738 581
rect 816 575 818 581
rect 888 575 890 581
rect 968 575 970 581
rect 1048 575 1050 581
rect 1128 575 1130 581
rect 190 574 196 575
rect 190 570 191 574
rect 195 570 196 574
rect 190 569 196 570
rect 278 574 284 575
rect 278 570 279 574
rect 283 570 284 574
rect 278 569 284 570
rect 366 574 372 575
rect 366 570 367 574
rect 371 570 372 574
rect 366 569 372 570
rect 462 574 468 575
rect 462 570 463 574
rect 467 570 468 574
rect 462 569 468 570
rect 558 574 564 575
rect 558 570 559 574
rect 563 570 564 574
rect 558 569 564 570
rect 646 574 652 575
rect 646 570 647 574
rect 651 570 652 574
rect 646 569 652 570
rect 734 574 740 575
rect 734 570 735 574
rect 739 570 740 574
rect 734 569 740 570
rect 814 574 820 575
rect 814 570 815 574
rect 819 570 820 574
rect 814 569 820 570
rect 886 574 892 575
rect 886 570 887 574
rect 891 570 892 574
rect 886 569 892 570
rect 966 574 972 575
rect 966 570 967 574
rect 971 570 972 574
rect 966 569 972 570
rect 1046 574 1052 575
rect 1046 570 1047 574
rect 1051 570 1052 574
rect 1046 569 1052 570
rect 1126 574 1132 575
rect 1126 570 1127 574
rect 1131 570 1132 574
rect 1126 569 1132 570
rect 1328 566 1330 581
rect 1368 579 1370 602
rect 1630 598 1636 599
rect 1630 594 1631 598
rect 1635 594 1636 598
rect 1630 593 1636 594
rect 1694 598 1700 599
rect 1694 594 1695 598
rect 1699 594 1700 598
rect 1694 593 1700 594
rect 1774 598 1780 599
rect 1774 594 1775 598
rect 1779 594 1780 598
rect 1774 593 1780 594
rect 1854 598 1860 599
rect 1854 594 1855 598
rect 1859 594 1860 598
rect 1854 593 1860 594
rect 1942 598 1948 599
rect 1942 594 1943 598
rect 1947 594 1948 598
rect 1942 593 1948 594
rect 2030 598 2036 599
rect 2030 594 2031 598
rect 2035 594 2036 598
rect 2030 593 2036 594
rect 2110 598 2116 599
rect 2110 594 2111 598
rect 2115 594 2116 598
rect 2110 593 2116 594
rect 2190 598 2196 599
rect 2190 594 2191 598
rect 2195 594 2196 598
rect 2190 593 2196 594
rect 2270 598 2276 599
rect 2270 594 2271 598
rect 2275 594 2276 598
rect 2270 593 2276 594
rect 2342 598 2348 599
rect 2342 594 2343 598
rect 2347 594 2348 598
rect 2342 593 2348 594
rect 2414 598 2420 599
rect 2414 594 2415 598
rect 2419 594 2420 598
rect 2414 593 2420 594
rect 2486 598 2492 599
rect 2486 594 2487 598
rect 2491 594 2492 598
rect 2486 593 2492 594
rect 2542 598 2548 599
rect 2542 594 2543 598
rect 2547 594 2548 598
rect 2542 593 2548 594
rect 1632 579 1634 593
rect 1696 579 1698 593
rect 1776 579 1778 593
rect 1856 579 1858 593
rect 1944 579 1946 593
rect 2032 579 2034 593
rect 2112 579 2114 593
rect 2192 579 2194 593
rect 2272 579 2274 593
rect 2344 579 2346 593
rect 2416 579 2418 593
rect 2488 579 2490 593
rect 2544 579 2546 593
rect 2584 579 2586 602
rect 1367 578 1371 579
rect 1367 573 1371 574
rect 1511 578 1515 579
rect 1511 573 1515 574
rect 1575 578 1579 579
rect 1575 573 1579 574
rect 1631 578 1635 579
rect 1631 573 1635 574
rect 1655 578 1659 579
rect 1655 573 1659 574
rect 1695 578 1699 579
rect 1695 573 1699 574
rect 1735 578 1739 579
rect 1735 573 1739 574
rect 1775 578 1779 579
rect 1775 573 1779 574
rect 1823 578 1827 579
rect 1823 573 1827 574
rect 1855 578 1859 579
rect 1855 573 1859 574
rect 1911 578 1915 579
rect 1911 573 1915 574
rect 1943 578 1947 579
rect 1943 573 1947 574
rect 1999 578 2003 579
rect 1999 573 2003 574
rect 2031 578 2035 579
rect 2031 573 2035 574
rect 2087 578 2091 579
rect 2087 573 2091 574
rect 2111 578 2115 579
rect 2111 573 2115 574
rect 2175 578 2179 579
rect 2175 573 2179 574
rect 2191 578 2195 579
rect 2191 573 2195 574
rect 2271 578 2275 579
rect 2271 573 2275 574
rect 2343 578 2347 579
rect 2343 573 2347 574
rect 2367 578 2371 579
rect 2367 573 2371 574
rect 2415 578 2419 579
rect 2415 573 2419 574
rect 2463 578 2467 579
rect 2463 573 2467 574
rect 2487 578 2491 579
rect 2487 573 2491 574
rect 2543 578 2547 579
rect 2543 573 2547 574
rect 2583 578 2587 579
rect 2583 573 2587 574
rect 110 565 116 566
rect 110 561 111 565
rect 115 561 116 565
rect 110 560 116 561
rect 1326 565 1332 566
rect 1326 561 1327 565
rect 1331 561 1332 565
rect 1326 560 1332 561
rect 1368 558 1370 573
rect 1512 567 1514 573
rect 1576 567 1578 573
rect 1656 567 1658 573
rect 1736 567 1738 573
rect 1824 567 1826 573
rect 1912 567 1914 573
rect 2000 567 2002 573
rect 2088 567 2090 573
rect 2176 567 2178 573
rect 2272 567 2274 573
rect 2368 567 2370 573
rect 2464 567 2466 573
rect 2544 567 2546 573
rect 1510 566 1516 567
rect 1510 562 1511 566
rect 1515 562 1516 566
rect 1510 561 1516 562
rect 1574 566 1580 567
rect 1574 562 1575 566
rect 1579 562 1580 566
rect 1574 561 1580 562
rect 1654 566 1660 567
rect 1654 562 1655 566
rect 1659 562 1660 566
rect 1654 561 1660 562
rect 1734 566 1740 567
rect 1734 562 1735 566
rect 1739 562 1740 566
rect 1734 561 1740 562
rect 1822 566 1828 567
rect 1822 562 1823 566
rect 1827 562 1828 566
rect 1822 561 1828 562
rect 1910 566 1916 567
rect 1910 562 1911 566
rect 1915 562 1916 566
rect 1910 561 1916 562
rect 1998 566 2004 567
rect 1998 562 1999 566
rect 2003 562 2004 566
rect 1998 561 2004 562
rect 2086 566 2092 567
rect 2086 562 2087 566
rect 2091 562 2092 566
rect 2086 561 2092 562
rect 2174 566 2180 567
rect 2174 562 2175 566
rect 2179 562 2180 566
rect 2174 561 2180 562
rect 2270 566 2276 567
rect 2270 562 2271 566
rect 2275 562 2276 566
rect 2270 561 2276 562
rect 2366 566 2372 567
rect 2366 562 2367 566
rect 2371 562 2372 566
rect 2366 561 2372 562
rect 2462 566 2468 567
rect 2462 562 2463 566
rect 2467 562 2468 566
rect 2462 561 2468 562
rect 2542 566 2548 567
rect 2542 562 2543 566
rect 2547 562 2548 566
rect 2542 561 2548 562
rect 2584 558 2586 573
rect 1366 557 1372 558
rect 1366 553 1367 557
rect 1371 553 1372 557
rect 1366 552 1372 553
rect 2582 557 2588 558
rect 2582 553 2583 557
rect 2587 553 2588 557
rect 2582 552 2588 553
rect 110 548 116 549
rect 1326 548 1332 549
rect 110 544 111 548
rect 115 544 116 548
rect 110 543 116 544
rect 174 547 180 548
rect 174 543 175 547
rect 179 543 180 547
rect 112 527 114 543
rect 174 542 180 543
rect 262 547 268 548
rect 262 543 263 547
rect 267 543 268 547
rect 262 542 268 543
rect 350 547 356 548
rect 350 543 351 547
rect 355 543 356 547
rect 350 542 356 543
rect 446 547 452 548
rect 446 543 447 547
rect 451 543 452 547
rect 446 542 452 543
rect 542 547 548 548
rect 542 543 543 547
rect 547 543 548 547
rect 542 542 548 543
rect 630 547 636 548
rect 630 543 631 547
rect 635 543 636 547
rect 630 542 636 543
rect 718 547 724 548
rect 718 543 719 547
rect 723 543 724 547
rect 718 542 724 543
rect 798 547 804 548
rect 798 543 799 547
rect 803 543 804 547
rect 798 542 804 543
rect 870 547 876 548
rect 870 543 871 547
rect 875 543 876 547
rect 870 542 876 543
rect 950 547 956 548
rect 950 543 951 547
rect 955 543 956 547
rect 950 542 956 543
rect 1030 547 1036 548
rect 1030 543 1031 547
rect 1035 543 1036 547
rect 1030 542 1036 543
rect 1110 547 1116 548
rect 1110 543 1111 547
rect 1115 543 1116 547
rect 1326 544 1327 548
rect 1331 544 1332 548
rect 1326 543 1332 544
rect 1110 542 1116 543
rect 176 527 178 542
rect 264 527 266 542
rect 352 527 354 542
rect 448 527 450 542
rect 544 527 546 542
rect 632 527 634 542
rect 720 527 722 542
rect 800 527 802 542
rect 872 527 874 542
rect 952 527 954 542
rect 1032 527 1034 542
rect 1112 527 1114 542
rect 1328 527 1330 543
rect 1366 540 1372 541
rect 2582 540 2588 541
rect 1366 536 1367 540
rect 1371 536 1372 540
rect 1366 535 1372 536
rect 1494 539 1500 540
rect 1494 535 1495 539
rect 1499 535 1500 539
rect 111 526 115 527
rect 111 521 115 522
rect 143 526 147 527
rect 143 521 147 522
rect 175 526 179 527
rect 175 521 179 522
rect 207 526 211 527
rect 207 521 211 522
rect 263 526 267 527
rect 263 521 267 522
rect 311 526 315 527
rect 311 521 315 522
rect 351 526 355 527
rect 351 521 355 522
rect 431 526 435 527
rect 431 521 435 522
rect 447 526 451 527
rect 447 521 451 522
rect 543 526 547 527
rect 543 521 547 522
rect 551 526 555 527
rect 551 521 555 522
rect 631 526 635 527
rect 631 521 635 522
rect 671 526 675 527
rect 671 521 675 522
rect 719 526 723 527
rect 719 521 723 522
rect 791 526 795 527
rect 791 521 795 522
rect 799 526 803 527
rect 799 521 803 522
rect 871 526 875 527
rect 871 521 875 522
rect 903 526 907 527
rect 903 521 907 522
rect 951 526 955 527
rect 951 521 955 522
rect 1007 526 1011 527
rect 1007 521 1011 522
rect 1031 526 1035 527
rect 1031 521 1035 522
rect 1103 526 1107 527
rect 1103 521 1107 522
rect 1111 526 1115 527
rect 1111 521 1115 522
rect 1199 526 1203 527
rect 1199 521 1203 522
rect 1271 526 1275 527
rect 1271 521 1275 522
rect 1327 526 1331 527
rect 1327 521 1331 522
rect 112 509 114 521
rect 144 510 146 521
rect 208 510 210 521
rect 312 510 314 521
rect 432 510 434 521
rect 552 510 554 521
rect 672 510 674 521
rect 792 510 794 521
rect 904 510 906 521
rect 1008 510 1010 521
rect 1104 510 1106 521
rect 1200 510 1202 521
rect 1272 510 1274 521
rect 142 509 148 510
rect 110 508 116 509
rect 110 504 111 508
rect 115 504 116 508
rect 142 505 143 509
rect 147 505 148 509
rect 142 504 148 505
rect 206 509 212 510
rect 206 505 207 509
rect 211 505 212 509
rect 206 504 212 505
rect 310 509 316 510
rect 310 505 311 509
rect 315 505 316 509
rect 310 504 316 505
rect 430 509 436 510
rect 430 505 431 509
rect 435 505 436 509
rect 430 504 436 505
rect 550 509 556 510
rect 550 505 551 509
rect 555 505 556 509
rect 550 504 556 505
rect 670 509 676 510
rect 670 505 671 509
rect 675 505 676 509
rect 670 504 676 505
rect 790 509 796 510
rect 790 505 791 509
rect 795 505 796 509
rect 790 504 796 505
rect 902 509 908 510
rect 902 505 903 509
rect 907 505 908 509
rect 902 504 908 505
rect 1006 509 1012 510
rect 1006 505 1007 509
rect 1011 505 1012 509
rect 1006 504 1012 505
rect 1102 509 1108 510
rect 1102 505 1103 509
rect 1107 505 1108 509
rect 1102 504 1108 505
rect 1198 509 1204 510
rect 1198 505 1199 509
rect 1203 505 1204 509
rect 1198 504 1204 505
rect 1270 509 1276 510
rect 1328 509 1330 521
rect 1368 519 1370 535
rect 1494 534 1500 535
rect 1558 539 1564 540
rect 1558 535 1559 539
rect 1563 535 1564 539
rect 1558 534 1564 535
rect 1638 539 1644 540
rect 1638 535 1639 539
rect 1643 535 1644 539
rect 1638 534 1644 535
rect 1718 539 1724 540
rect 1718 535 1719 539
rect 1723 535 1724 539
rect 1718 534 1724 535
rect 1806 539 1812 540
rect 1806 535 1807 539
rect 1811 535 1812 539
rect 1806 534 1812 535
rect 1894 539 1900 540
rect 1894 535 1895 539
rect 1899 535 1900 539
rect 1894 534 1900 535
rect 1982 539 1988 540
rect 1982 535 1983 539
rect 1987 535 1988 539
rect 1982 534 1988 535
rect 2070 539 2076 540
rect 2070 535 2071 539
rect 2075 535 2076 539
rect 2070 534 2076 535
rect 2158 539 2164 540
rect 2158 535 2159 539
rect 2163 535 2164 539
rect 2158 534 2164 535
rect 2254 539 2260 540
rect 2254 535 2255 539
rect 2259 535 2260 539
rect 2254 534 2260 535
rect 2350 539 2356 540
rect 2350 535 2351 539
rect 2355 535 2356 539
rect 2350 534 2356 535
rect 2446 539 2452 540
rect 2446 535 2447 539
rect 2451 535 2452 539
rect 2446 534 2452 535
rect 2526 539 2532 540
rect 2526 535 2527 539
rect 2531 535 2532 539
rect 2582 536 2583 540
rect 2587 536 2588 540
rect 2582 535 2588 536
rect 2526 534 2532 535
rect 1496 519 1498 534
rect 1560 519 1562 534
rect 1640 519 1642 534
rect 1720 519 1722 534
rect 1808 519 1810 534
rect 1896 519 1898 534
rect 1984 519 1986 534
rect 2072 519 2074 534
rect 2160 519 2162 534
rect 2256 519 2258 534
rect 2352 519 2354 534
rect 2448 519 2450 534
rect 2528 519 2530 534
rect 2584 519 2586 535
rect 1367 518 1371 519
rect 1367 513 1371 514
rect 1399 518 1403 519
rect 1399 513 1403 514
rect 1455 518 1459 519
rect 1455 513 1459 514
rect 1495 518 1499 519
rect 1495 513 1499 514
rect 1519 518 1523 519
rect 1519 513 1523 514
rect 1559 518 1563 519
rect 1559 513 1563 514
rect 1607 518 1611 519
rect 1607 513 1611 514
rect 1639 518 1643 519
rect 1639 513 1643 514
rect 1695 518 1699 519
rect 1695 513 1699 514
rect 1719 518 1723 519
rect 1719 513 1723 514
rect 1791 518 1795 519
rect 1791 513 1795 514
rect 1807 518 1811 519
rect 1807 513 1811 514
rect 1887 518 1891 519
rect 1887 513 1891 514
rect 1895 518 1899 519
rect 1895 513 1899 514
rect 1983 518 1987 519
rect 1983 513 1987 514
rect 2071 518 2075 519
rect 2071 513 2075 514
rect 2087 518 2091 519
rect 2087 513 2091 514
rect 2159 518 2163 519
rect 2159 513 2163 514
rect 2199 518 2203 519
rect 2199 513 2203 514
rect 2255 518 2259 519
rect 2255 513 2259 514
rect 2311 518 2315 519
rect 2311 513 2315 514
rect 2351 518 2355 519
rect 2351 513 2355 514
rect 2431 518 2435 519
rect 2431 513 2435 514
rect 2447 518 2451 519
rect 2447 513 2451 514
rect 2527 518 2531 519
rect 2527 513 2531 514
rect 2583 518 2587 519
rect 2583 513 2587 514
rect 1270 505 1271 509
rect 1275 505 1276 509
rect 1270 504 1276 505
rect 1326 508 1332 509
rect 1326 504 1327 508
rect 1331 504 1332 508
rect 110 503 116 504
rect 1326 503 1332 504
rect 1368 501 1370 513
rect 1400 502 1402 513
rect 1456 502 1458 513
rect 1520 502 1522 513
rect 1608 502 1610 513
rect 1696 502 1698 513
rect 1792 502 1794 513
rect 1888 502 1890 513
rect 1984 502 1986 513
rect 2088 502 2090 513
rect 2200 502 2202 513
rect 2312 502 2314 513
rect 2432 502 2434 513
rect 2528 502 2530 513
rect 1398 501 1404 502
rect 1366 500 1372 501
rect 1366 496 1367 500
rect 1371 496 1372 500
rect 1398 497 1399 501
rect 1403 497 1404 501
rect 1398 496 1404 497
rect 1454 501 1460 502
rect 1454 497 1455 501
rect 1459 497 1460 501
rect 1454 496 1460 497
rect 1518 501 1524 502
rect 1518 497 1519 501
rect 1523 497 1524 501
rect 1518 496 1524 497
rect 1606 501 1612 502
rect 1606 497 1607 501
rect 1611 497 1612 501
rect 1606 496 1612 497
rect 1694 501 1700 502
rect 1694 497 1695 501
rect 1699 497 1700 501
rect 1694 496 1700 497
rect 1790 501 1796 502
rect 1790 497 1791 501
rect 1795 497 1796 501
rect 1790 496 1796 497
rect 1886 501 1892 502
rect 1886 497 1887 501
rect 1891 497 1892 501
rect 1886 496 1892 497
rect 1982 501 1988 502
rect 1982 497 1983 501
rect 1987 497 1988 501
rect 1982 496 1988 497
rect 2086 501 2092 502
rect 2086 497 2087 501
rect 2091 497 2092 501
rect 2086 496 2092 497
rect 2198 501 2204 502
rect 2198 497 2199 501
rect 2203 497 2204 501
rect 2198 496 2204 497
rect 2310 501 2316 502
rect 2310 497 2311 501
rect 2315 497 2316 501
rect 2310 496 2316 497
rect 2430 501 2436 502
rect 2430 497 2431 501
rect 2435 497 2436 501
rect 2430 496 2436 497
rect 2526 501 2532 502
rect 2584 501 2586 513
rect 2526 497 2527 501
rect 2531 497 2532 501
rect 2526 496 2532 497
rect 2582 500 2588 501
rect 2582 496 2583 500
rect 2587 496 2588 500
rect 1366 495 1372 496
rect 2582 495 2588 496
rect 110 491 116 492
rect 110 487 111 491
rect 115 487 116 491
rect 110 486 116 487
rect 1326 491 1332 492
rect 1326 487 1327 491
rect 1331 487 1332 491
rect 1326 486 1332 487
rect 112 467 114 486
rect 158 482 164 483
rect 158 478 159 482
rect 163 478 164 482
rect 158 477 164 478
rect 222 482 228 483
rect 222 478 223 482
rect 227 478 228 482
rect 222 477 228 478
rect 326 482 332 483
rect 326 478 327 482
rect 331 478 332 482
rect 326 477 332 478
rect 446 482 452 483
rect 446 478 447 482
rect 451 478 452 482
rect 446 477 452 478
rect 566 482 572 483
rect 566 478 567 482
rect 571 478 572 482
rect 566 477 572 478
rect 686 482 692 483
rect 686 478 687 482
rect 691 478 692 482
rect 686 477 692 478
rect 806 482 812 483
rect 806 478 807 482
rect 811 478 812 482
rect 806 477 812 478
rect 918 482 924 483
rect 918 478 919 482
rect 923 478 924 482
rect 918 477 924 478
rect 1022 482 1028 483
rect 1022 478 1023 482
rect 1027 478 1028 482
rect 1022 477 1028 478
rect 1118 482 1124 483
rect 1118 478 1119 482
rect 1123 478 1124 482
rect 1118 477 1124 478
rect 1214 482 1220 483
rect 1214 478 1215 482
rect 1219 478 1220 482
rect 1214 477 1220 478
rect 1286 482 1292 483
rect 1286 478 1287 482
rect 1291 478 1292 482
rect 1286 477 1292 478
rect 160 467 162 477
rect 224 467 226 477
rect 328 467 330 477
rect 448 467 450 477
rect 568 467 570 477
rect 688 467 690 477
rect 808 467 810 477
rect 920 467 922 477
rect 1024 467 1026 477
rect 1120 467 1122 477
rect 1216 467 1218 477
rect 1288 467 1290 477
rect 1328 467 1330 486
rect 1366 483 1372 484
rect 1366 479 1367 483
rect 1371 479 1372 483
rect 1366 478 1372 479
rect 2582 483 2588 484
rect 2582 479 2583 483
rect 2587 479 2588 483
rect 2582 478 2588 479
rect 111 466 115 467
rect 111 461 115 462
rect 159 466 163 467
rect 159 461 163 462
rect 223 466 227 467
rect 223 461 227 462
rect 319 466 323 467
rect 319 461 323 462
rect 327 466 331 467
rect 327 461 331 462
rect 423 466 427 467
rect 423 461 427 462
rect 447 466 451 467
rect 447 461 451 462
rect 535 466 539 467
rect 535 461 539 462
rect 567 466 571 467
rect 567 461 571 462
rect 639 466 643 467
rect 639 461 643 462
rect 687 466 691 467
rect 687 461 691 462
rect 743 466 747 467
rect 743 461 747 462
rect 807 466 811 467
rect 807 461 811 462
rect 839 466 843 467
rect 839 461 843 462
rect 919 466 923 467
rect 919 461 923 462
rect 927 466 931 467
rect 927 461 931 462
rect 1007 466 1011 467
rect 1007 461 1011 462
rect 1023 466 1027 467
rect 1023 461 1027 462
rect 1079 466 1083 467
rect 1079 461 1083 462
rect 1119 466 1123 467
rect 1119 461 1123 462
rect 1151 466 1155 467
rect 1151 461 1155 462
rect 1215 466 1219 467
rect 1215 461 1219 462
rect 1231 466 1235 467
rect 1231 461 1235 462
rect 1287 466 1291 467
rect 1287 461 1291 462
rect 1327 466 1331 467
rect 1327 461 1331 462
rect 112 446 114 461
rect 160 455 162 461
rect 224 455 226 461
rect 320 455 322 461
rect 424 455 426 461
rect 536 455 538 461
rect 640 455 642 461
rect 744 455 746 461
rect 840 455 842 461
rect 928 455 930 461
rect 1008 455 1010 461
rect 1080 455 1082 461
rect 1152 455 1154 461
rect 1232 455 1234 461
rect 1288 455 1290 461
rect 158 454 164 455
rect 158 450 159 454
rect 163 450 164 454
rect 158 449 164 450
rect 222 454 228 455
rect 222 450 223 454
rect 227 450 228 454
rect 222 449 228 450
rect 318 454 324 455
rect 318 450 319 454
rect 323 450 324 454
rect 318 449 324 450
rect 422 454 428 455
rect 422 450 423 454
rect 427 450 428 454
rect 422 449 428 450
rect 534 454 540 455
rect 534 450 535 454
rect 539 450 540 454
rect 534 449 540 450
rect 638 454 644 455
rect 638 450 639 454
rect 643 450 644 454
rect 638 449 644 450
rect 742 454 748 455
rect 742 450 743 454
rect 747 450 748 454
rect 742 449 748 450
rect 838 454 844 455
rect 838 450 839 454
rect 843 450 844 454
rect 838 449 844 450
rect 926 454 932 455
rect 926 450 927 454
rect 931 450 932 454
rect 926 449 932 450
rect 1006 454 1012 455
rect 1006 450 1007 454
rect 1011 450 1012 454
rect 1006 449 1012 450
rect 1078 454 1084 455
rect 1078 450 1079 454
rect 1083 450 1084 454
rect 1078 449 1084 450
rect 1150 454 1156 455
rect 1150 450 1151 454
rect 1155 450 1156 454
rect 1150 449 1156 450
rect 1230 454 1236 455
rect 1230 450 1231 454
rect 1235 450 1236 454
rect 1230 449 1236 450
rect 1286 454 1292 455
rect 1286 450 1287 454
rect 1291 450 1292 454
rect 1286 449 1292 450
rect 1328 446 1330 461
rect 1368 455 1370 478
rect 1414 474 1420 475
rect 1414 470 1415 474
rect 1419 470 1420 474
rect 1414 469 1420 470
rect 1470 474 1476 475
rect 1470 470 1471 474
rect 1475 470 1476 474
rect 1470 469 1476 470
rect 1534 474 1540 475
rect 1534 470 1535 474
rect 1539 470 1540 474
rect 1534 469 1540 470
rect 1622 474 1628 475
rect 1622 470 1623 474
rect 1627 470 1628 474
rect 1622 469 1628 470
rect 1710 474 1716 475
rect 1710 470 1711 474
rect 1715 470 1716 474
rect 1710 469 1716 470
rect 1806 474 1812 475
rect 1806 470 1807 474
rect 1811 470 1812 474
rect 1806 469 1812 470
rect 1902 474 1908 475
rect 1902 470 1903 474
rect 1907 470 1908 474
rect 1902 469 1908 470
rect 1998 474 2004 475
rect 1998 470 1999 474
rect 2003 470 2004 474
rect 1998 469 2004 470
rect 2102 474 2108 475
rect 2102 470 2103 474
rect 2107 470 2108 474
rect 2102 469 2108 470
rect 2214 474 2220 475
rect 2214 470 2215 474
rect 2219 470 2220 474
rect 2214 469 2220 470
rect 2326 474 2332 475
rect 2326 470 2327 474
rect 2331 470 2332 474
rect 2326 469 2332 470
rect 2446 474 2452 475
rect 2446 470 2447 474
rect 2451 470 2452 474
rect 2446 469 2452 470
rect 2542 474 2548 475
rect 2542 470 2543 474
rect 2547 470 2548 474
rect 2542 469 2548 470
rect 1416 455 1418 469
rect 1472 455 1474 469
rect 1536 455 1538 469
rect 1624 455 1626 469
rect 1712 455 1714 469
rect 1808 455 1810 469
rect 1904 455 1906 469
rect 2000 455 2002 469
rect 2104 455 2106 469
rect 2216 455 2218 469
rect 2328 455 2330 469
rect 2448 455 2450 469
rect 2544 455 2546 469
rect 2584 455 2586 478
rect 1367 454 1371 455
rect 1367 449 1371 450
rect 1415 454 1419 455
rect 1415 449 1419 450
rect 1471 454 1475 455
rect 1471 449 1475 450
rect 1487 454 1491 455
rect 1487 449 1491 450
rect 1535 454 1539 455
rect 1535 449 1539 450
rect 1575 454 1579 455
rect 1575 449 1579 450
rect 1623 454 1627 455
rect 1623 449 1627 450
rect 1663 454 1667 455
rect 1663 449 1667 450
rect 1711 454 1715 455
rect 1711 449 1715 450
rect 1759 454 1763 455
rect 1759 449 1763 450
rect 1807 454 1811 455
rect 1807 449 1811 450
rect 1863 454 1867 455
rect 1863 449 1867 450
rect 1903 454 1907 455
rect 1903 449 1907 450
rect 1975 454 1979 455
rect 1975 449 1979 450
rect 1999 454 2003 455
rect 1999 449 2003 450
rect 2103 454 2107 455
rect 2103 449 2107 450
rect 2111 454 2115 455
rect 2111 449 2115 450
rect 2215 454 2219 455
rect 2215 449 2219 450
rect 2255 454 2259 455
rect 2255 449 2259 450
rect 2327 454 2331 455
rect 2327 449 2331 450
rect 2407 454 2411 455
rect 2407 449 2411 450
rect 2447 454 2451 455
rect 2447 449 2451 450
rect 2543 454 2547 455
rect 2543 449 2547 450
rect 2583 454 2587 455
rect 2583 449 2587 450
rect 110 445 116 446
rect 110 441 111 445
rect 115 441 116 445
rect 110 440 116 441
rect 1326 445 1332 446
rect 1326 441 1327 445
rect 1331 441 1332 445
rect 1326 440 1332 441
rect 1368 434 1370 449
rect 1416 443 1418 449
rect 1488 443 1490 449
rect 1576 443 1578 449
rect 1664 443 1666 449
rect 1760 443 1762 449
rect 1864 443 1866 449
rect 1976 443 1978 449
rect 2112 443 2114 449
rect 2256 443 2258 449
rect 2408 443 2410 449
rect 2544 443 2546 449
rect 1414 442 1420 443
rect 1414 438 1415 442
rect 1419 438 1420 442
rect 1414 437 1420 438
rect 1486 442 1492 443
rect 1486 438 1487 442
rect 1491 438 1492 442
rect 1486 437 1492 438
rect 1574 442 1580 443
rect 1574 438 1575 442
rect 1579 438 1580 442
rect 1574 437 1580 438
rect 1662 442 1668 443
rect 1662 438 1663 442
rect 1667 438 1668 442
rect 1662 437 1668 438
rect 1758 442 1764 443
rect 1758 438 1759 442
rect 1763 438 1764 442
rect 1758 437 1764 438
rect 1862 442 1868 443
rect 1862 438 1863 442
rect 1867 438 1868 442
rect 1862 437 1868 438
rect 1974 442 1980 443
rect 1974 438 1975 442
rect 1979 438 1980 442
rect 1974 437 1980 438
rect 2110 442 2116 443
rect 2110 438 2111 442
rect 2115 438 2116 442
rect 2110 437 2116 438
rect 2254 442 2260 443
rect 2254 438 2255 442
rect 2259 438 2260 442
rect 2254 437 2260 438
rect 2406 442 2412 443
rect 2406 438 2407 442
rect 2411 438 2412 442
rect 2406 437 2412 438
rect 2542 442 2548 443
rect 2542 438 2543 442
rect 2547 438 2548 442
rect 2542 437 2548 438
rect 2584 434 2586 449
rect 1366 433 1372 434
rect 1366 429 1367 433
rect 1371 429 1372 433
rect 110 428 116 429
rect 1326 428 1332 429
rect 1366 428 1372 429
rect 2582 433 2588 434
rect 2582 429 2583 433
rect 2587 429 2588 433
rect 2582 428 2588 429
rect 110 424 111 428
rect 115 424 116 428
rect 110 423 116 424
rect 142 427 148 428
rect 142 423 143 427
rect 147 423 148 427
rect 112 403 114 423
rect 142 422 148 423
rect 206 427 212 428
rect 206 423 207 427
rect 211 423 212 427
rect 206 422 212 423
rect 302 427 308 428
rect 302 423 303 427
rect 307 423 308 427
rect 302 422 308 423
rect 406 427 412 428
rect 406 423 407 427
rect 411 423 412 427
rect 406 422 412 423
rect 518 427 524 428
rect 518 423 519 427
rect 523 423 524 427
rect 518 422 524 423
rect 622 427 628 428
rect 622 423 623 427
rect 627 423 628 427
rect 622 422 628 423
rect 726 427 732 428
rect 726 423 727 427
rect 731 423 732 427
rect 726 422 732 423
rect 822 427 828 428
rect 822 423 823 427
rect 827 423 828 427
rect 822 422 828 423
rect 910 427 916 428
rect 910 423 911 427
rect 915 423 916 427
rect 910 422 916 423
rect 990 427 996 428
rect 990 423 991 427
rect 995 423 996 427
rect 990 422 996 423
rect 1062 427 1068 428
rect 1062 423 1063 427
rect 1067 423 1068 427
rect 1062 422 1068 423
rect 1134 427 1140 428
rect 1134 423 1135 427
rect 1139 423 1140 427
rect 1134 422 1140 423
rect 1214 427 1220 428
rect 1214 423 1215 427
rect 1219 423 1220 427
rect 1214 422 1220 423
rect 1270 427 1276 428
rect 1270 423 1271 427
rect 1275 423 1276 427
rect 1326 424 1327 428
rect 1331 424 1332 428
rect 1326 423 1332 424
rect 1270 422 1276 423
rect 144 403 146 422
rect 208 403 210 422
rect 304 403 306 422
rect 408 403 410 422
rect 520 403 522 422
rect 624 403 626 422
rect 728 403 730 422
rect 824 403 826 422
rect 912 403 914 422
rect 992 403 994 422
rect 1064 403 1066 422
rect 1136 403 1138 422
rect 1216 403 1218 422
rect 1272 403 1274 422
rect 1328 403 1330 423
rect 1366 416 1372 417
rect 2582 416 2588 417
rect 1366 412 1367 416
rect 1371 412 1372 416
rect 1366 411 1372 412
rect 1398 415 1404 416
rect 1398 411 1399 415
rect 1403 411 1404 415
rect 111 402 115 403
rect 111 397 115 398
rect 143 402 147 403
rect 143 397 147 398
rect 207 402 211 403
rect 207 397 211 398
rect 303 402 307 403
rect 303 397 307 398
rect 399 402 403 403
rect 399 397 403 398
rect 407 402 411 403
rect 407 397 411 398
rect 495 402 499 403
rect 495 397 499 398
rect 519 402 523 403
rect 519 397 523 398
rect 583 402 587 403
rect 583 397 587 398
rect 623 402 627 403
rect 623 397 627 398
rect 671 402 675 403
rect 671 397 675 398
rect 727 402 731 403
rect 727 397 731 398
rect 751 402 755 403
rect 751 397 755 398
rect 823 402 827 403
rect 823 397 827 398
rect 895 402 899 403
rect 895 397 899 398
rect 911 402 915 403
rect 911 397 915 398
rect 967 402 971 403
rect 967 397 971 398
rect 991 402 995 403
rect 991 397 995 398
rect 1047 402 1051 403
rect 1047 397 1051 398
rect 1063 402 1067 403
rect 1063 397 1067 398
rect 1135 402 1139 403
rect 1135 397 1139 398
rect 1215 402 1219 403
rect 1215 397 1219 398
rect 1271 402 1275 403
rect 1271 397 1275 398
rect 1327 402 1331 403
rect 1327 397 1331 398
rect 112 385 114 397
rect 144 386 146 397
rect 208 386 210 397
rect 304 386 306 397
rect 400 386 402 397
rect 496 386 498 397
rect 584 386 586 397
rect 672 386 674 397
rect 752 386 754 397
rect 824 386 826 397
rect 896 386 898 397
rect 968 386 970 397
rect 1048 386 1050 397
rect 142 385 148 386
rect 110 384 116 385
rect 110 380 111 384
rect 115 380 116 384
rect 142 381 143 385
rect 147 381 148 385
rect 142 380 148 381
rect 206 385 212 386
rect 206 381 207 385
rect 211 381 212 385
rect 206 380 212 381
rect 302 385 308 386
rect 302 381 303 385
rect 307 381 308 385
rect 302 380 308 381
rect 398 385 404 386
rect 398 381 399 385
rect 403 381 404 385
rect 398 380 404 381
rect 494 385 500 386
rect 494 381 495 385
rect 499 381 500 385
rect 494 380 500 381
rect 582 385 588 386
rect 582 381 583 385
rect 587 381 588 385
rect 582 380 588 381
rect 670 385 676 386
rect 670 381 671 385
rect 675 381 676 385
rect 670 380 676 381
rect 750 385 756 386
rect 750 381 751 385
rect 755 381 756 385
rect 750 380 756 381
rect 822 385 828 386
rect 822 381 823 385
rect 827 381 828 385
rect 822 380 828 381
rect 894 385 900 386
rect 894 381 895 385
rect 899 381 900 385
rect 894 380 900 381
rect 966 385 972 386
rect 966 381 967 385
rect 971 381 972 385
rect 966 380 972 381
rect 1046 385 1052 386
rect 1328 385 1330 397
rect 1368 395 1370 411
rect 1398 410 1404 411
rect 1470 415 1476 416
rect 1470 411 1471 415
rect 1475 411 1476 415
rect 1470 410 1476 411
rect 1558 415 1564 416
rect 1558 411 1559 415
rect 1563 411 1564 415
rect 1558 410 1564 411
rect 1646 415 1652 416
rect 1646 411 1647 415
rect 1651 411 1652 415
rect 1646 410 1652 411
rect 1742 415 1748 416
rect 1742 411 1743 415
rect 1747 411 1748 415
rect 1742 410 1748 411
rect 1846 415 1852 416
rect 1846 411 1847 415
rect 1851 411 1852 415
rect 1846 410 1852 411
rect 1958 415 1964 416
rect 1958 411 1959 415
rect 1963 411 1964 415
rect 1958 410 1964 411
rect 2094 415 2100 416
rect 2094 411 2095 415
rect 2099 411 2100 415
rect 2094 410 2100 411
rect 2238 415 2244 416
rect 2238 411 2239 415
rect 2243 411 2244 415
rect 2238 410 2244 411
rect 2390 415 2396 416
rect 2390 411 2391 415
rect 2395 411 2396 415
rect 2390 410 2396 411
rect 2526 415 2532 416
rect 2526 411 2527 415
rect 2531 411 2532 415
rect 2582 412 2583 416
rect 2587 412 2588 416
rect 2582 411 2588 412
rect 2526 410 2532 411
rect 1400 395 1402 410
rect 1472 395 1474 410
rect 1560 395 1562 410
rect 1648 395 1650 410
rect 1744 395 1746 410
rect 1848 395 1850 410
rect 1960 395 1962 410
rect 2096 395 2098 410
rect 2240 395 2242 410
rect 2392 395 2394 410
rect 2528 395 2530 410
rect 2584 395 2586 411
rect 1367 394 1371 395
rect 1367 389 1371 390
rect 1399 394 1403 395
rect 1399 389 1403 390
rect 1455 394 1459 395
rect 1455 389 1459 390
rect 1471 394 1475 395
rect 1471 389 1475 390
rect 1511 394 1515 395
rect 1511 389 1515 390
rect 1559 394 1563 395
rect 1559 389 1563 390
rect 1567 394 1571 395
rect 1567 389 1571 390
rect 1631 394 1635 395
rect 1631 389 1635 390
rect 1647 394 1651 395
rect 1647 389 1651 390
rect 1695 394 1699 395
rect 1695 389 1699 390
rect 1743 394 1747 395
rect 1743 389 1747 390
rect 1759 394 1763 395
rect 1759 389 1763 390
rect 1839 394 1843 395
rect 1839 389 1843 390
rect 1847 394 1851 395
rect 1847 389 1851 390
rect 1943 394 1947 395
rect 1943 389 1947 390
rect 1959 394 1963 395
rect 1959 389 1963 390
rect 2071 394 2075 395
rect 2071 389 2075 390
rect 2095 394 2099 395
rect 2095 389 2099 390
rect 2215 394 2219 395
rect 2215 389 2219 390
rect 2239 394 2243 395
rect 2239 389 2243 390
rect 2367 394 2371 395
rect 2367 389 2371 390
rect 2391 394 2395 395
rect 2391 389 2395 390
rect 2527 394 2531 395
rect 2527 389 2531 390
rect 2583 394 2587 395
rect 2583 389 2587 390
rect 1046 381 1047 385
rect 1051 381 1052 385
rect 1046 380 1052 381
rect 1326 384 1332 385
rect 1326 380 1327 384
rect 1331 380 1332 384
rect 110 379 116 380
rect 1326 379 1332 380
rect 1368 377 1370 389
rect 1400 378 1402 389
rect 1456 378 1458 389
rect 1512 378 1514 389
rect 1568 378 1570 389
rect 1632 378 1634 389
rect 1696 378 1698 389
rect 1760 378 1762 389
rect 1840 378 1842 389
rect 1944 378 1946 389
rect 2072 378 2074 389
rect 2216 378 2218 389
rect 2368 378 2370 389
rect 2528 378 2530 389
rect 1398 377 1404 378
rect 1366 376 1372 377
rect 1366 372 1367 376
rect 1371 372 1372 376
rect 1398 373 1399 377
rect 1403 373 1404 377
rect 1398 372 1404 373
rect 1454 377 1460 378
rect 1454 373 1455 377
rect 1459 373 1460 377
rect 1454 372 1460 373
rect 1510 377 1516 378
rect 1510 373 1511 377
rect 1515 373 1516 377
rect 1510 372 1516 373
rect 1566 377 1572 378
rect 1566 373 1567 377
rect 1571 373 1572 377
rect 1566 372 1572 373
rect 1630 377 1636 378
rect 1630 373 1631 377
rect 1635 373 1636 377
rect 1630 372 1636 373
rect 1694 377 1700 378
rect 1694 373 1695 377
rect 1699 373 1700 377
rect 1694 372 1700 373
rect 1758 377 1764 378
rect 1758 373 1759 377
rect 1763 373 1764 377
rect 1758 372 1764 373
rect 1838 377 1844 378
rect 1838 373 1839 377
rect 1843 373 1844 377
rect 1838 372 1844 373
rect 1942 377 1948 378
rect 1942 373 1943 377
rect 1947 373 1948 377
rect 1942 372 1948 373
rect 2070 377 2076 378
rect 2070 373 2071 377
rect 2075 373 2076 377
rect 2070 372 2076 373
rect 2214 377 2220 378
rect 2214 373 2215 377
rect 2219 373 2220 377
rect 2214 372 2220 373
rect 2366 377 2372 378
rect 2366 373 2367 377
rect 2371 373 2372 377
rect 2366 372 2372 373
rect 2526 377 2532 378
rect 2584 377 2586 389
rect 2526 373 2527 377
rect 2531 373 2532 377
rect 2526 372 2532 373
rect 2582 376 2588 377
rect 2582 372 2583 376
rect 2587 372 2588 376
rect 1366 371 1372 372
rect 2582 371 2588 372
rect 110 367 116 368
rect 110 363 111 367
rect 115 363 116 367
rect 110 362 116 363
rect 1326 367 1332 368
rect 1326 363 1327 367
rect 1331 363 1332 367
rect 1326 362 1332 363
rect 112 343 114 362
rect 158 358 164 359
rect 158 354 159 358
rect 163 354 164 358
rect 158 353 164 354
rect 222 358 228 359
rect 222 354 223 358
rect 227 354 228 358
rect 222 353 228 354
rect 318 358 324 359
rect 318 354 319 358
rect 323 354 324 358
rect 318 353 324 354
rect 414 358 420 359
rect 414 354 415 358
rect 419 354 420 358
rect 414 353 420 354
rect 510 358 516 359
rect 510 354 511 358
rect 515 354 516 358
rect 510 353 516 354
rect 598 358 604 359
rect 598 354 599 358
rect 603 354 604 358
rect 598 353 604 354
rect 686 358 692 359
rect 686 354 687 358
rect 691 354 692 358
rect 686 353 692 354
rect 766 358 772 359
rect 766 354 767 358
rect 771 354 772 358
rect 766 353 772 354
rect 838 358 844 359
rect 838 354 839 358
rect 843 354 844 358
rect 838 353 844 354
rect 910 358 916 359
rect 910 354 911 358
rect 915 354 916 358
rect 910 353 916 354
rect 982 358 988 359
rect 982 354 983 358
rect 987 354 988 358
rect 982 353 988 354
rect 1062 358 1068 359
rect 1062 354 1063 358
rect 1067 354 1068 358
rect 1062 353 1068 354
rect 160 343 162 353
rect 224 343 226 353
rect 320 343 322 353
rect 416 343 418 353
rect 512 343 514 353
rect 600 343 602 353
rect 688 343 690 353
rect 768 343 770 353
rect 840 343 842 353
rect 912 343 914 353
rect 984 343 986 353
rect 1064 343 1066 353
rect 1328 343 1330 362
rect 1366 359 1372 360
rect 1366 355 1367 359
rect 1371 355 1372 359
rect 1366 354 1372 355
rect 2582 359 2588 360
rect 2582 355 2583 359
rect 2587 355 2588 359
rect 2582 354 2588 355
rect 111 342 115 343
rect 111 337 115 338
rect 159 342 163 343
rect 159 337 163 338
rect 223 342 227 343
rect 223 337 227 338
rect 311 342 315 343
rect 311 337 315 338
rect 319 342 323 343
rect 319 337 323 338
rect 391 342 395 343
rect 391 337 395 338
rect 415 342 419 343
rect 415 337 419 338
rect 471 342 475 343
rect 471 337 475 338
rect 511 342 515 343
rect 511 337 515 338
rect 543 342 547 343
rect 543 337 547 338
rect 599 342 603 343
rect 599 337 603 338
rect 607 342 611 343
rect 607 337 611 338
rect 671 342 675 343
rect 671 337 675 338
rect 687 342 691 343
rect 687 337 691 338
rect 735 342 739 343
rect 735 337 739 338
rect 767 342 771 343
rect 767 337 771 338
rect 799 342 803 343
rect 799 337 803 338
rect 839 342 843 343
rect 839 337 843 338
rect 863 342 867 343
rect 863 337 867 338
rect 911 342 915 343
rect 911 337 915 338
rect 935 342 939 343
rect 935 337 939 338
rect 983 342 987 343
rect 983 337 987 338
rect 1063 342 1067 343
rect 1063 337 1067 338
rect 1327 342 1331 343
rect 1327 337 1331 338
rect 112 322 114 337
rect 160 331 162 337
rect 224 331 226 337
rect 312 331 314 337
rect 392 331 394 337
rect 472 331 474 337
rect 544 331 546 337
rect 608 331 610 337
rect 672 331 674 337
rect 736 331 738 337
rect 800 331 802 337
rect 864 331 866 337
rect 936 331 938 337
rect 158 330 164 331
rect 158 326 159 330
rect 163 326 164 330
rect 158 325 164 326
rect 222 330 228 331
rect 222 326 223 330
rect 227 326 228 330
rect 222 325 228 326
rect 310 330 316 331
rect 310 326 311 330
rect 315 326 316 330
rect 310 325 316 326
rect 390 330 396 331
rect 390 326 391 330
rect 395 326 396 330
rect 390 325 396 326
rect 470 330 476 331
rect 470 326 471 330
rect 475 326 476 330
rect 470 325 476 326
rect 542 330 548 331
rect 542 326 543 330
rect 547 326 548 330
rect 542 325 548 326
rect 606 330 612 331
rect 606 326 607 330
rect 611 326 612 330
rect 606 325 612 326
rect 670 330 676 331
rect 670 326 671 330
rect 675 326 676 330
rect 670 325 676 326
rect 734 330 740 331
rect 734 326 735 330
rect 739 326 740 330
rect 734 325 740 326
rect 798 330 804 331
rect 798 326 799 330
rect 803 326 804 330
rect 798 325 804 326
rect 862 330 868 331
rect 862 326 863 330
rect 867 326 868 330
rect 862 325 868 326
rect 934 330 940 331
rect 934 326 935 330
rect 939 326 940 330
rect 934 325 940 326
rect 1328 322 1330 337
rect 1368 335 1370 354
rect 1414 350 1420 351
rect 1414 346 1415 350
rect 1419 346 1420 350
rect 1414 345 1420 346
rect 1470 350 1476 351
rect 1470 346 1471 350
rect 1475 346 1476 350
rect 1470 345 1476 346
rect 1526 350 1532 351
rect 1526 346 1527 350
rect 1531 346 1532 350
rect 1526 345 1532 346
rect 1582 350 1588 351
rect 1582 346 1583 350
rect 1587 346 1588 350
rect 1582 345 1588 346
rect 1646 350 1652 351
rect 1646 346 1647 350
rect 1651 346 1652 350
rect 1646 345 1652 346
rect 1710 350 1716 351
rect 1710 346 1711 350
rect 1715 346 1716 350
rect 1710 345 1716 346
rect 1774 350 1780 351
rect 1774 346 1775 350
rect 1779 346 1780 350
rect 1774 345 1780 346
rect 1854 350 1860 351
rect 1854 346 1855 350
rect 1859 346 1860 350
rect 1854 345 1860 346
rect 1958 350 1964 351
rect 1958 346 1959 350
rect 1963 346 1964 350
rect 1958 345 1964 346
rect 2086 350 2092 351
rect 2086 346 2087 350
rect 2091 346 2092 350
rect 2086 345 2092 346
rect 2230 350 2236 351
rect 2230 346 2231 350
rect 2235 346 2236 350
rect 2230 345 2236 346
rect 2382 350 2388 351
rect 2382 346 2383 350
rect 2387 346 2388 350
rect 2382 345 2388 346
rect 2542 350 2548 351
rect 2542 346 2543 350
rect 2547 346 2548 350
rect 2542 345 2548 346
rect 1416 335 1418 345
rect 1472 335 1474 345
rect 1528 335 1530 345
rect 1584 335 1586 345
rect 1648 335 1650 345
rect 1712 335 1714 345
rect 1776 335 1778 345
rect 1856 335 1858 345
rect 1960 335 1962 345
rect 2088 335 2090 345
rect 2232 335 2234 345
rect 2384 335 2386 345
rect 2544 335 2546 345
rect 2584 335 2586 354
rect 1367 334 1371 335
rect 1367 329 1371 330
rect 1415 334 1419 335
rect 1415 329 1419 330
rect 1471 334 1475 335
rect 1471 329 1475 330
rect 1527 334 1531 335
rect 1527 329 1531 330
rect 1583 334 1587 335
rect 1583 329 1587 330
rect 1607 334 1611 335
rect 1607 329 1611 330
rect 1647 334 1651 335
rect 1647 329 1651 330
rect 1663 334 1667 335
rect 1663 329 1667 330
rect 1711 334 1715 335
rect 1711 329 1715 330
rect 1719 334 1723 335
rect 1719 329 1723 330
rect 1775 334 1779 335
rect 1775 329 1779 330
rect 1831 334 1835 335
rect 1831 329 1835 330
rect 1855 334 1859 335
rect 1855 329 1859 330
rect 1887 334 1891 335
rect 1887 329 1891 330
rect 1951 334 1955 335
rect 1951 329 1955 330
rect 1959 334 1963 335
rect 1959 329 1963 330
rect 2031 334 2035 335
rect 2031 329 2035 330
rect 2087 334 2091 335
rect 2087 329 2091 330
rect 2119 334 2123 335
rect 2119 329 2123 330
rect 2223 334 2227 335
rect 2223 329 2227 330
rect 2231 334 2235 335
rect 2231 329 2235 330
rect 2335 334 2339 335
rect 2335 329 2339 330
rect 2383 334 2387 335
rect 2383 329 2387 330
rect 2447 334 2451 335
rect 2447 329 2451 330
rect 2543 334 2547 335
rect 2543 329 2547 330
rect 2583 334 2587 335
rect 2583 329 2587 330
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 110 316 116 317
rect 1326 321 1332 322
rect 1326 317 1327 321
rect 1331 317 1332 321
rect 1326 316 1332 317
rect 1368 314 1370 329
rect 1608 323 1610 329
rect 1664 323 1666 329
rect 1720 323 1722 329
rect 1776 323 1778 329
rect 1832 323 1834 329
rect 1888 323 1890 329
rect 1952 323 1954 329
rect 2032 323 2034 329
rect 2120 323 2122 329
rect 2224 323 2226 329
rect 2336 323 2338 329
rect 2448 323 2450 329
rect 2544 323 2546 329
rect 1606 322 1612 323
rect 1606 318 1607 322
rect 1611 318 1612 322
rect 1606 317 1612 318
rect 1662 322 1668 323
rect 1662 318 1663 322
rect 1667 318 1668 322
rect 1662 317 1668 318
rect 1718 322 1724 323
rect 1718 318 1719 322
rect 1723 318 1724 322
rect 1718 317 1724 318
rect 1774 322 1780 323
rect 1774 318 1775 322
rect 1779 318 1780 322
rect 1774 317 1780 318
rect 1830 322 1836 323
rect 1830 318 1831 322
rect 1835 318 1836 322
rect 1830 317 1836 318
rect 1886 322 1892 323
rect 1886 318 1887 322
rect 1891 318 1892 322
rect 1886 317 1892 318
rect 1950 322 1956 323
rect 1950 318 1951 322
rect 1955 318 1956 322
rect 1950 317 1956 318
rect 2030 322 2036 323
rect 2030 318 2031 322
rect 2035 318 2036 322
rect 2030 317 2036 318
rect 2118 322 2124 323
rect 2118 318 2119 322
rect 2123 318 2124 322
rect 2118 317 2124 318
rect 2222 322 2228 323
rect 2222 318 2223 322
rect 2227 318 2228 322
rect 2222 317 2228 318
rect 2334 322 2340 323
rect 2334 318 2335 322
rect 2339 318 2340 322
rect 2334 317 2340 318
rect 2446 322 2452 323
rect 2446 318 2447 322
rect 2451 318 2452 322
rect 2446 317 2452 318
rect 2542 322 2548 323
rect 2542 318 2543 322
rect 2547 318 2548 322
rect 2542 317 2548 318
rect 2584 314 2586 329
rect 1366 313 1372 314
rect 1366 309 1367 313
rect 1371 309 1372 313
rect 1366 308 1372 309
rect 2582 313 2588 314
rect 2582 309 2583 313
rect 2587 309 2588 313
rect 2582 308 2588 309
rect 110 304 116 305
rect 1326 304 1332 305
rect 110 300 111 304
rect 115 300 116 304
rect 110 299 116 300
rect 142 303 148 304
rect 142 299 143 303
rect 147 299 148 303
rect 112 279 114 299
rect 142 298 148 299
rect 206 303 212 304
rect 206 299 207 303
rect 211 299 212 303
rect 206 298 212 299
rect 294 303 300 304
rect 294 299 295 303
rect 299 299 300 303
rect 294 298 300 299
rect 374 303 380 304
rect 374 299 375 303
rect 379 299 380 303
rect 374 298 380 299
rect 454 303 460 304
rect 454 299 455 303
rect 459 299 460 303
rect 454 298 460 299
rect 526 303 532 304
rect 526 299 527 303
rect 531 299 532 303
rect 526 298 532 299
rect 590 303 596 304
rect 590 299 591 303
rect 595 299 596 303
rect 590 298 596 299
rect 654 303 660 304
rect 654 299 655 303
rect 659 299 660 303
rect 654 298 660 299
rect 718 303 724 304
rect 718 299 719 303
rect 723 299 724 303
rect 718 298 724 299
rect 782 303 788 304
rect 782 299 783 303
rect 787 299 788 303
rect 782 298 788 299
rect 846 303 852 304
rect 846 299 847 303
rect 851 299 852 303
rect 846 298 852 299
rect 918 303 924 304
rect 918 299 919 303
rect 923 299 924 303
rect 1326 300 1327 304
rect 1331 300 1332 304
rect 1326 299 1332 300
rect 918 298 924 299
rect 144 279 146 298
rect 208 279 210 298
rect 296 279 298 298
rect 376 279 378 298
rect 456 279 458 298
rect 528 279 530 298
rect 592 279 594 298
rect 656 279 658 298
rect 720 279 722 298
rect 784 279 786 298
rect 848 279 850 298
rect 920 279 922 298
rect 1328 279 1330 299
rect 1366 296 1372 297
rect 2582 296 2588 297
rect 1366 292 1367 296
rect 1371 292 1372 296
rect 1366 291 1372 292
rect 1590 295 1596 296
rect 1590 291 1591 295
rect 1595 291 1596 295
rect 111 278 115 279
rect 111 273 115 274
rect 143 278 147 279
rect 143 273 147 274
rect 207 278 211 279
rect 207 273 211 274
rect 231 278 235 279
rect 231 273 235 274
rect 295 278 299 279
rect 295 273 299 274
rect 335 278 339 279
rect 335 273 339 274
rect 375 278 379 279
rect 375 273 379 274
rect 431 278 435 279
rect 431 273 435 274
rect 455 278 459 279
rect 455 273 459 274
rect 519 278 523 279
rect 519 273 523 274
rect 527 278 531 279
rect 527 273 531 274
rect 591 278 595 279
rect 591 273 595 274
rect 599 278 603 279
rect 599 273 603 274
rect 655 278 659 279
rect 655 273 659 274
rect 679 278 683 279
rect 679 273 683 274
rect 719 278 723 279
rect 719 273 723 274
rect 751 278 755 279
rect 751 273 755 274
rect 783 278 787 279
rect 783 273 787 274
rect 815 278 819 279
rect 815 273 819 274
rect 847 278 851 279
rect 847 273 851 274
rect 887 278 891 279
rect 887 273 891 274
rect 919 278 923 279
rect 919 273 923 274
rect 959 278 963 279
rect 959 273 963 274
rect 1031 278 1035 279
rect 1031 273 1035 274
rect 1327 278 1331 279
rect 1368 275 1370 291
rect 1590 290 1596 291
rect 1646 295 1652 296
rect 1646 291 1647 295
rect 1651 291 1652 295
rect 1646 290 1652 291
rect 1702 295 1708 296
rect 1702 291 1703 295
rect 1707 291 1708 295
rect 1702 290 1708 291
rect 1758 295 1764 296
rect 1758 291 1759 295
rect 1763 291 1764 295
rect 1758 290 1764 291
rect 1814 295 1820 296
rect 1814 291 1815 295
rect 1819 291 1820 295
rect 1814 290 1820 291
rect 1870 295 1876 296
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 1870 290 1876 291
rect 1934 295 1940 296
rect 1934 291 1935 295
rect 1939 291 1940 295
rect 1934 290 1940 291
rect 2014 295 2020 296
rect 2014 291 2015 295
rect 2019 291 2020 295
rect 2014 290 2020 291
rect 2102 295 2108 296
rect 2102 291 2103 295
rect 2107 291 2108 295
rect 2102 290 2108 291
rect 2206 295 2212 296
rect 2206 291 2207 295
rect 2211 291 2212 295
rect 2206 290 2212 291
rect 2318 295 2324 296
rect 2318 291 2319 295
rect 2323 291 2324 295
rect 2318 290 2324 291
rect 2430 295 2436 296
rect 2430 291 2431 295
rect 2435 291 2436 295
rect 2430 290 2436 291
rect 2526 295 2532 296
rect 2526 291 2527 295
rect 2531 291 2532 295
rect 2582 292 2583 296
rect 2587 292 2588 296
rect 2582 291 2588 292
rect 2526 290 2532 291
rect 1592 275 1594 290
rect 1648 275 1650 290
rect 1704 275 1706 290
rect 1760 275 1762 290
rect 1816 275 1818 290
rect 1872 275 1874 290
rect 1936 275 1938 290
rect 2016 275 2018 290
rect 2104 275 2106 290
rect 2208 275 2210 290
rect 2320 275 2322 290
rect 2432 275 2434 290
rect 2528 275 2530 290
rect 2584 275 2586 291
rect 1327 273 1331 274
rect 1367 274 1371 275
rect 112 261 114 273
rect 144 262 146 273
rect 232 262 234 273
rect 336 262 338 273
rect 432 262 434 273
rect 520 262 522 273
rect 600 262 602 273
rect 680 262 682 273
rect 752 262 754 273
rect 816 262 818 273
rect 888 262 890 273
rect 960 262 962 273
rect 1032 262 1034 273
rect 142 261 148 262
rect 110 260 116 261
rect 110 256 111 260
rect 115 256 116 260
rect 142 257 143 261
rect 147 257 148 261
rect 142 256 148 257
rect 230 261 236 262
rect 230 257 231 261
rect 235 257 236 261
rect 230 256 236 257
rect 334 261 340 262
rect 334 257 335 261
rect 339 257 340 261
rect 334 256 340 257
rect 430 261 436 262
rect 430 257 431 261
rect 435 257 436 261
rect 430 256 436 257
rect 518 261 524 262
rect 518 257 519 261
rect 523 257 524 261
rect 518 256 524 257
rect 598 261 604 262
rect 598 257 599 261
rect 603 257 604 261
rect 598 256 604 257
rect 678 261 684 262
rect 678 257 679 261
rect 683 257 684 261
rect 678 256 684 257
rect 750 261 756 262
rect 750 257 751 261
rect 755 257 756 261
rect 750 256 756 257
rect 814 261 820 262
rect 814 257 815 261
rect 819 257 820 261
rect 814 256 820 257
rect 886 261 892 262
rect 886 257 887 261
rect 891 257 892 261
rect 886 256 892 257
rect 958 261 964 262
rect 958 257 959 261
rect 963 257 964 261
rect 958 256 964 257
rect 1030 261 1036 262
rect 1328 261 1330 273
rect 1367 269 1371 270
rect 1591 274 1595 275
rect 1591 269 1595 270
rect 1647 274 1651 275
rect 1647 269 1651 270
rect 1703 274 1707 275
rect 1703 269 1707 270
rect 1727 274 1731 275
rect 1727 269 1731 270
rect 1759 274 1763 275
rect 1759 269 1763 270
rect 1783 274 1787 275
rect 1783 269 1787 270
rect 1815 274 1819 275
rect 1815 269 1819 270
rect 1839 274 1843 275
rect 1839 269 1843 270
rect 1871 274 1875 275
rect 1871 269 1875 270
rect 1895 274 1899 275
rect 1895 269 1899 270
rect 1935 274 1939 275
rect 1935 269 1939 270
rect 1951 274 1955 275
rect 1951 269 1955 270
rect 2007 274 2011 275
rect 2007 269 2011 270
rect 2015 274 2019 275
rect 2015 269 2019 270
rect 2071 274 2075 275
rect 2071 269 2075 270
rect 2103 274 2107 275
rect 2103 269 2107 270
rect 2143 274 2147 275
rect 2143 269 2147 270
rect 2207 274 2211 275
rect 2207 269 2211 270
rect 2231 274 2235 275
rect 2231 269 2235 270
rect 2319 274 2323 275
rect 2319 269 2323 270
rect 2335 274 2339 275
rect 2335 269 2339 270
rect 2431 274 2435 275
rect 2431 269 2435 270
rect 2439 274 2443 275
rect 2439 269 2443 270
rect 2527 274 2531 275
rect 2527 269 2531 270
rect 2583 274 2587 275
rect 2583 269 2587 270
rect 1030 257 1031 261
rect 1035 257 1036 261
rect 1030 256 1036 257
rect 1326 260 1332 261
rect 1326 256 1327 260
rect 1331 256 1332 260
rect 1368 257 1370 269
rect 1728 258 1730 269
rect 1784 258 1786 269
rect 1840 258 1842 269
rect 1896 258 1898 269
rect 1952 258 1954 269
rect 2008 258 2010 269
rect 2072 258 2074 269
rect 2144 258 2146 269
rect 2232 258 2234 269
rect 2336 258 2338 269
rect 2440 258 2442 269
rect 2528 258 2530 269
rect 1726 257 1732 258
rect 110 255 116 256
rect 1326 255 1332 256
rect 1366 256 1372 257
rect 1366 252 1367 256
rect 1371 252 1372 256
rect 1726 253 1727 257
rect 1731 253 1732 257
rect 1726 252 1732 253
rect 1782 257 1788 258
rect 1782 253 1783 257
rect 1787 253 1788 257
rect 1782 252 1788 253
rect 1838 257 1844 258
rect 1838 253 1839 257
rect 1843 253 1844 257
rect 1838 252 1844 253
rect 1894 257 1900 258
rect 1894 253 1895 257
rect 1899 253 1900 257
rect 1894 252 1900 253
rect 1950 257 1956 258
rect 1950 253 1951 257
rect 1955 253 1956 257
rect 1950 252 1956 253
rect 2006 257 2012 258
rect 2006 253 2007 257
rect 2011 253 2012 257
rect 2006 252 2012 253
rect 2070 257 2076 258
rect 2070 253 2071 257
rect 2075 253 2076 257
rect 2070 252 2076 253
rect 2142 257 2148 258
rect 2142 253 2143 257
rect 2147 253 2148 257
rect 2142 252 2148 253
rect 2230 257 2236 258
rect 2230 253 2231 257
rect 2235 253 2236 257
rect 2230 252 2236 253
rect 2334 257 2340 258
rect 2334 253 2335 257
rect 2339 253 2340 257
rect 2334 252 2340 253
rect 2438 257 2444 258
rect 2438 253 2439 257
rect 2443 253 2444 257
rect 2438 252 2444 253
rect 2526 257 2532 258
rect 2584 257 2586 269
rect 2526 253 2527 257
rect 2531 253 2532 257
rect 2526 252 2532 253
rect 2582 256 2588 257
rect 2582 252 2583 256
rect 2587 252 2588 256
rect 1366 251 1372 252
rect 2582 251 2588 252
rect 110 243 116 244
rect 110 239 111 243
rect 115 239 116 243
rect 110 238 116 239
rect 1326 243 1332 244
rect 1326 239 1327 243
rect 1331 239 1332 243
rect 1326 238 1332 239
rect 1366 239 1372 240
rect 112 219 114 238
rect 158 234 164 235
rect 158 230 159 234
rect 163 230 164 234
rect 158 229 164 230
rect 246 234 252 235
rect 246 230 247 234
rect 251 230 252 234
rect 246 229 252 230
rect 350 234 356 235
rect 350 230 351 234
rect 355 230 356 234
rect 350 229 356 230
rect 446 234 452 235
rect 446 230 447 234
rect 451 230 452 234
rect 446 229 452 230
rect 534 234 540 235
rect 534 230 535 234
rect 539 230 540 234
rect 534 229 540 230
rect 614 234 620 235
rect 614 230 615 234
rect 619 230 620 234
rect 614 229 620 230
rect 694 234 700 235
rect 694 230 695 234
rect 699 230 700 234
rect 694 229 700 230
rect 766 234 772 235
rect 766 230 767 234
rect 771 230 772 234
rect 766 229 772 230
rect 830 234 836 235
rect 830 230 831 234
rect 835 230 836 234
rect 830 229 836 230
rect 902 234 908 235
rect 902 230 903 234
rect 907 230 908 234
rect 902 229 908 230
rect 974 234 980 235
rect 974 230 975 234
rect 979 230 980 234
rect 974 229 980 230
rect 1046 234 1052 235
rect 1046 230 1047 234
rect 1051 230 1052 234
rect 1046 229 1052 230
rect 160 219 162 229
rect 248 219 250 229
rect 352 219 354 229
rect 448 219 450 229
rect 536 219 538 229
rect 616 219 618 229
rect 696 219 698 229
rect 768 219 770 229
rect 832 219 834 229
rect 904 219 906 229
rect 976 219 978 229
rect 1048 219 1050 229
rect 1328 219 1330 238
rect 1366 235 1367 239
rect 1371 235 1372 239
rect 1366 234 1372 235
rect 2582 239 2588 240
rect 2582 235 2583 239
rect 2587 235 2588 239
rect 2582 234 2588 235
rect 1368 219 1370 234
rect 1742 230 1748 231
rect 1742 226 1743 230
rect 1747 226 1748 230
rect 1742 225 1748 226
rect 1798 230 1804 231
rect 1798 226 1799 230
rect 1803 226 1804 230
rect 1798 225 1804 226
rect 1854 230 1860 231
rect 1854 226 1855 230
rect 1859 226 1860 230
rect 1854 225 1860 226
rect 1910 230 1916 231
rect 1910 226 1911 230
rect 1915 226 1916 230
rect 1910 225 1916 226
rect 1966 230 1972 231
rect 1966 226 1967 230
rect 1971 226 1972 230
rect 1966 225 1972 226
rect 2022 230 2028 231
rect 2022 226 2023 230
rect 2027 226 2028 230
rect 2022 225 2028 226
rect 2086 230 2092 231
rect 2086 226 2087 230
rect 2091 226 2092 230
rect 2086 225 2092 226
rect 2158 230 2164 231
rect 2158 226 2159 230
rect 2163 226 2164 230
rect 2158 225 2164 226
rect 2246 230 2252 231
rect 2246 226 2247 230
rect 2251 226 2252 230
rect 2246 225 2252 226
rect 2350 230 2356 231
rect 2350 226 2351 230
rect 2355 226 2356 230
rect 2350 225 2356 226
rect 2454 230 2460 231
rect 2454 226 2455 230
rect 2459 226 2460 230
rect 2454 225 2460 226
rect 2542 230 2548 231
rect 2542 226 2543 230
rect 2547 226 2548 230
rect 2542 225 2548 226
rect 1744 219 1746 225
rect 1800 219 1802 225
rect 1856 219 1858 225
rect 1912 219 1914 225
rect 1968 219 1970 225
rect 2024 219 2026 225
rect 2088 219 2090 225
rect 2160 219 2162 225
rect 2248 219 2250 225
rect 2352 219 2354 225
rect 2456 219 2458 225
rect 2544 219 2546 225
rect 2584 219 2586 234
rect 111 218 115 219
rect 111 213 115 214
rect 159 218 163 219
rect 159 213 163 214
rect 167 218 171 219
rect 167 213 171 214
rect 247 218 251 219
rect 247 213 251 214
rect 255 218 259 219
rect 255 213 259 214
rect 351 218 355 219
rect 351 213 355 214
rect 447 218 451 219
rect 447 213 451 214
rect 535 218 539 219
rect 535 213 539 214
rect 551 218 555 219
rect 551 213 555 214
rect 615 218 619 219
rect 615 213 619 214
rect 655 218 659 219
rect 655 213 659 214
rect 695 218 699 219
rect 695 213 699 214
rect 751 218 755 219
rect 751 213 755 214
rect 767 218 771 219
rect 767 213 771 214
rect 831 218 835 219
rect 831 213 835 214
rect 847 218 851 219
rect 847 213 851 214
rect 903 218 907 219
rect 903 213 907 214
rect 935 218 939 219
rect 935 213 939 214
rect 975 218 979 219
rect 975 213 979 214
rect 1023 218 1027 219
rect 1023 213 1027 214
rect 1047 218 1051 219
rect 1047 213 1051 214
rect 1111 218 1115 219
rect 1111 213 1115 214
rect 1199 218 1203 219
rect 1199 213 1203 214
rect 1327 218 1331 219
rect 1327 213 1331 214
rect 1367 218 1371 219
rect 1367 213 1371 214
rect 1463 218 1467 219
rect 1463 213 1467 214
rect 1535 218 1539 219
rect 1535 213 1539 214
rect 1623 218 1627 219
rect 1623 213 1627 214
rect 1719 218 1723 219
rect 1719 213 1723 214
rect 1743 218 1747 219
rect 1743 213 1747 214
rect 1799 218 1803 219
rect 1799 213 1803 214
rect 1823 218 1827 219
rect 1823 213 1827 214
rect 1855 218 1859 219
rect 1855 213 1859 214
rect 1911 218 1915 219
rect 1911 213 1915 214
rect 1927 218 1931 219
rect 1927 213 1931 214
rect 1967 218 1971 219
rect 1967 213 1971 214
rect 2023 218 2027 219
rect 2023 213 2027 214
rect 2031 218 2035 219
rect 2031 213 2035 214
rect 2087 218 2091 219
rect 2087 213 2091 214
rect 2135 218 2139 219
rect 2135 213 2139 214
rect 2159 218 2163 219
rect 2159 213 2163 214
rect 2239 218 2243 219
rect 2239 213 2243 214
rect 2247 218 2251 219
rect 2247 213 2251 214
rect 2343 218 2347 219
rect 2343 213 2347 214
rect 2351 218 2355 219
rect 2351 213 2355 214
rect 2455 218 2459 219
rect 2455 213 2459 214
rect 2543 218 2547 219
rect 2543 213 2547 214
rect 2583 218 2587 219
rect 2583 213 2587 214
rect 112 198 114 213
rect 168 207 170 213
rect 256 207 258 213
rect 352 207 354 213
rect 448 207 450 213
rect 552 207 554 213
rect 656 207 658 213
rect 752 207 754 213
rect 848 207 850 213
rect 936 207 938 213
rect 1024 207 1026 213
rect 1112 207 1114 213
rect 1200 207 1202 213
rect 166 206 172 207
rect 166 202 167 206
rect 171 202 172 206
rect 166 201 172 202
rect 254 206 260 207
rect 254 202 255 206
rect 259 202 260 206
rect 254 201 260 202
rect 350 206 356 207
rect 350 202 351 206
rect 355 202 356 206
rect 350 201 356 202
rect 446 206 452 207
rect 446 202 447 206
rect 451 202 452 206
rect 446 201 452 202
rect 550 206 556 207
rect 550 202 551 206
rect 555 202 556 206
rect 550 201 556 202
rect 654 206 660 207
rect 654 202 655 206
rect 659 202 660 206
rect 654 201 660 202
rect 750 206 756 207
rect 750 202 751 206
rect 755 202 756 206
rect 750 201 756 202
rect 846 206 852 207
rect 846 202 847 206
rect 851 202 852 206
rect 846 201 852 202
rect 934 206 940 207
rect 934 202 935 206
rect 939 202 940 206
rect 934 201 940 202
rect 1022 206 1028 207
rect 1022 202 1023 206
rect 1027 202 1028 206
rect 1022 201 1028 202
rect 1110 206 1116 207
rect 1110 202 1111 206
rect 1115 202 1116 206
rect 1110 201 1116 202
rect 1198 206 1204 207
rect 1198 202 1199 206
rect 1203 202 1204 206
rect 1198 201 1204 202
rect 1328 198 1330 213
rect 1368 198 1370 213
rect 1464 207 1466 213
rect 1536 207 1538 213
rect 1624 207 1626 213
rect 1720 207 1722 213
rect 1824 207 1826 213
rect 1928 207 1930 213
rect 2032 207 2034 213
rect 2136 207 2138 213
rect 2240 207 2242 213
rect 2344 207 2346 213
rect 2456 207 2458 213
rect 2544 207 2546 213
rect 1462 206 1468 207
rect 1462 202 1463 206
rect 1467 202 1468 206
rect 1462 201 1468 202
rect 1534 206 1540 207
rect 1534 202 1535 206
rect 1539 202 1540 206
rect 1534 201 1540 202
rect 1622 206 1628 207
rect 1622 202 1623 206
rect 1627 202 1628 206
rect 1622 201 1628 202
rect 1718 206 1724 207
rect 1718 202 1719 206
rect 1723 202 1724 206
rect 1718 201 1724 202
rect 1822 206 1828 207
rect 1822 202 1823 206
rect 1827 202 1828 206
rect 1822 201 1828 202
rect 1926 206 1932 207
rect 1926 202 1927 206
rect 1931 202 1932 206
rect 1926 201 1932 202
rect 2030 206 2036 207
rect 2030 202 2031 206
rect 2035 202 2036 206
rect 2030 201 2036 202
rect 2134 206 2140 207
rect 2134 202 2135 206
rect 2139 202 2140 206
rect 2134 201 2140 202
rect 2238 206 2244 207
rect 2238 202 2239 206
rect 2243 202 2244 206
rect 2238 201 2244 202
rect 2342 206 2348 207
rect 2342 202 2343 206
rect 2347 202 2348 206
rect 2342 201 2348 202
rect 2454 206 2460 207
rect 2454 202 2455 206
rect 2459 202 2460 206
rect 2454 201 2460 202
rect 2542 206 2548 207
rect 2542 202 2543 206
rect 2547 202 2548 206
rect 2542 201 2548 202
rect 2584 198 2586 213
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 110 192 116 193
rect 1326 197 1332 198
rect 1326 193 1327 197
rect 1331 193 1332 197
rect 1326 192 1332 193
rect 1366 197 1372 198
rect 1366 193 1367 197
rect 1371 193 1372 197
rect 1366 192 1372 193
rect 2582 197 2588 198
rect 2582 193 2583 197
rect 2587 193 2588 197
rect 2582 192 2588 193
rect 110 180 116 181
rect 1326 180 1332 181
rect 110 176 111 180
rect 115 176 116 180
rect 110 175 116 176
rect 150 179 156 180
rect 150 175 151 179
rect 155 175 156 179
rect 112 139 114 175
rect 150 174 156 175
rect 238 179 244 180
rect 238 175 239 179
rect 243 175 244 179
rect 238 174 244 175
rect 334 179 340 180
rect 334 175 335 179
rect 339 175 340 179
rect 334 174 340 175
rect 430 179 436 180
rect 430 175 431 179
rect 435 175 436 179
rect 430 174 436 175
rect 534 179 540 180
rect 534 175 535 179
rect 539 175 540 179
rect 534 174 540 175
rect 638 179 644 180
rect 638 175 639 179
rect 643 175 644 179
rect 638 174 644 175
rect 734 179 740 180
rect 734 175 735 179
rect 739 175 740 179
rect 734 174 740 175
rect 830 179 836 180
rect 830 175 831 179
rect 835 175 836 179
rect 830 174 836 175
rect 918 179 924 180
rect 918 175 919 179
rect 923 175 924 179
rect 918 174 924 175
rect 1006 179 1012 180
rect 1006 175 1007 179
rect 1011 175 1012 179
rect 1006 174 1012 175
rect 1094 179 1100 180
rect 1094 175 1095 179
rect 1099 175 1100 179
rect 1094 174 1100 175
rect 1182 179 1188 180
rect 1182 175 1183 179
rect 1187 175 1188 179
rect 1326 176 1327 180
rect 1331 176 1332 180
rect 1326 175 1332 176
rect 1366 180 1372 181
rect 2582 180 2588 181
rect 1366 176 1367 180
rect 1371 176 1372 180
rect 1366 175 1372 176
rect 1446 179 1452 180
rect 1446 175 1447 179
rect 1451 175 1452 179
rect 1182 174 1188 175
rect 152 139 154 174
rect 240 139 242 174
rect 336 139 338 174
rect 432 139 434 174
rect 536 139 538 174
rect 640 139 642 174
rect 736 139 738 174
rect 832 139 834 174
rect 920 139 922 174
rect 1008 139 1010 174
rect 1096 139 1098 174
rect 1184 139 1186 174
rect 1328 139 1330 175
rect 1368 147 1370 175
rect 1446 174 1452 175
rect 1518 179 1524 180
rect 1518 175 1519 179
rect 1523 175 1524 179
rect 1518 174 1524 175
rect 1606 179 1612 180
rect 1606 175 1607 179
rect 1611 175 1612 179
rect 1606 174 1612 175
rect 1702 179 1708 180
rect 1702 175 1703 179
rect 1707 175 1708 179
rect 1702 174 1708 175
rect 1806 179 1812 180
rect 1806 175 1807 179
rect 1811 175 1812 179
rect 1806 174 1812 175
rect 1910 179 1916 180
rect 1910 175 1911 179
rect 1915 175 1916 179
rect 1910 174 1916 175
rect 2014 179 2020 180
rect 2014 175 2015 179
rect 2019 175 2020 179
rect 2014 174 2020 175
rect 2118 179 2124 180
rect 2118 175 2119 179
rect 2123 175 2124 179
rect 2118 174 2124 175
rect 2222 179 2228 180
rect 2222 175 2223 179
rect 2227 175 2228 179
rect 2222 174 2228 175
rect 2326 179 2332 180
rect 2326 175 2327 179
rect 2331 175 2332 179
rect 2326 174 2332 175
rect 2438 179 2444 180
rect 2438 175 2439 179
rect 2443 175 2444 179
rect 2438 174 2444 175
rect 2526 179 2532 180
rect 2526 175 2527 179
rect 2531 175 2532 179
rect 2582 176 2583 180
rect 2587 176 2588 180
rect 2582 175 2588 176
rect 2526 174 2532 175
rect 1448 147 1450 174
rect 1520 147 1522 174
rect 1608 147 1610 174
rect 1704 147 1706 174
rect 1808 147 1810 174
rect 1912 147 1914 174
rect 2016 147 2018 174
rect 2120 147 2122 174
rect 2224 147 2226 174
rect 2328 147 2330 174
rect 2440 147 2442 174
rect 2528 147 2530 174
rect 2584 147 2586 175
rect 1367 146 1371 147
rect 1367 141 1371 142
rect 1399 146 1403 147
rect 1399 141 1403 142
rect 1447 146 1451 147
rect 1447 141 1451 142
rect 1455 146 1459 147
rect 1455 141 1459 142
rect 1511 146 1515 147
rect 1511 141 1515 142
rect 1519 146 1523 147
rect 1519 141 1523 142
rect 1567 146 1571 147
rect 1567 141 1571 142
rect 1607 146 1611 147
rect 1607 141 1611 142
rect 1639 146 1643 147
rect 1639 141 1643 142
rect 1703 146 1707 147
rect 1703 141 1707 142
rect 1719 146 1723 147
rect 1719 141 1723 142
rect 1799 146 1803 147
rect 1799 141 1803 142
rect 1807 146 1811 147
rect 1807 141 1811 142
rect 1879 146 1883 147
rect 1879 141 1883 142
rect 1911 146 1915 147
rect 1911 141 1915 142
rect 1959 146 1963 147
rect 1959 141 1963 142
rect 2015 146 2019 147
rect 2015 141 2019 142
rect 2031 146 2035 147
rect 2031 141 2035 142
rect 2103 146 2107 147
rect 2103 141 2107 142
rect 2119 146 2123 147
rect 2119 141 2123 142
rect 2167 146 2171 147
rect 2167 141 2171 142
rect 2223 146 2227 147
rect 2223 141 2227 142
rect 2231 146 2235 147
rect 2231 141 2235 142
rect 2295 146 2299 147
rect 2295 141 2299 142
rect 2327 146 2331 147
rect 2327 141 2331 142
rect 2359 146 2363 147
rect 2359 141 2363 142
rect 2415 146 2419 147
rect 2415 141 2419 142
rect 2439 146 2443 147
rect 2439 141 2443 142
rect 2471 146 2475 147
rect 2471 141 2475 142
rect 2527 146 2531 147
rect 2527 141 2531 142
rect 2583 146 2587 147
rect 2583 141 2587 142
rect 111 138 115 139
rect 111 133 115 134
rect 143 138 147 139
rect 143 133 147 134
rect 151 138 155 139
rect 151 133 155 134
rect 199 138 203 139
rect 199 133 203 134
rect 239 138 243 139
rect 239 133 243 134
rect 255 138 259 139
rect 255 133 259 134
rect 311 138 315 139
rect 311 133 315 134
rect 335 138 339 139
rect 335 133 339 134
rect 367 138 371 139
rect 367 133 371 134
rect 423 138 427 139
rect 423 133 427 134
rect 431 138 435 139
rect 431 133 435 134
rect 479 138 483 139
rect 479 133 483 134
rect 535 138 539 139
rect 535 133 539 134
rect 607 138 611 139
rect 607 133 611 134
rect 639 138 643 139
rect 639 133 643 134
rect 671 138 675 139
rect 671 133 675 134
rect 735 138 739 139
rect 735 133 739 134
rect 799 138 803 139
rect 799 133 803 134
rect 831 138 835 139
rect 831 133 835 134
rect 855 138 859 139
rect 855 133 859 134
rect 911 138 915 139
rect 911 133 915 134
rect 919 138 923 139
rect 919 133 923 134
rect 975 138 979 139
rect 975 133 979 134
rect 1007 138 1011 139
rect 1007 133 1011 134
rect 1039 138 1043 139
rect 1039 133 1043 134
rect 1095 138 1099 139
rect 1095 133 1099 134
rect 1103 138 1107 139
rect 1103 133 1107 134
rect 1159 138 1163 139
rect 1159 133 1163 134
rect 1183 138 1187 139
rect 1183 133 1187 134
rect 1215 138 1219 139
rect 1215 133 1219 134
rect 1271 138 1275 139
rect 1271 133 1275 134
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 112 121 114 133
rect 144 122 146 133
rect 200 122 202 133
rect 256 122 258 133
rect 312 122 314 133
rect 368 122 370 133
rect 424 122 426 133
rect 480 122 482 133
rect 536 122 538 133
rect 608 122 610 133
rect 672 122 674 133
rect 736 122 738 133
rect 800 122 802 133
rect 856 122 858 133
rect 912 122 914 133
rect 976 122 978 133
rect 1040 122 1042 133
rect 1104 122 1106 133
rect 1160 122 1162 133
rect 1216 122 1218 133
rect 1272 122 1274 133
rect 142 121 148 122
rect 110 120 116 121
rect 110 116 111 120
rect 115 116 116 120
rect 142 117 143 121
rect 147 117 148 121
rect 142 116 148 117
rect 198 121 204 122
rect 198 117 199 121
rect 203 117 204 121
rect 198 116 204 117
rect 254 121 260 122
rect 254 117 255 121
rect 259 117 260 121
rect 254 116 260 117
rect 310 121 316 122
rect 310 117 311 121
rect 315 117 316 121
rect 310 116 316 117
rect 366 121 372 122
rect 366 117 367 121
rect 371 117 372 121
rect 366 116 372 117
rect 422 121 428 122
rect 422 117 423 121
rect 427 117 428 121
rect 422 116 428 117
rect 478 121 484 122
rect 478 117 479 121
rect 483 117 484 121
rect 478 116 484 117
rect 534 121 540 122
rect 534 117 535 121
rect 539 117 540 121
rect 534 116 540 117
rect 606 121 612 122
rect 606 117 607 121
rect 611 117 612 121
rect 606 116 612 117
rect 670 121 676 122
rect 670 117 671 121
rect 675 117 676 121
rect 670 116 676 117
rect 734 121 740 122
rect 734 117 735 121
rect 739 117 740 121
rect 734 116 740 117
rect 798 121 804 122
rect 798 117 799 121
rect 803 117 804 121
rect 798 116 804 117
rect 854 121 860 122
rect 854 117 855 121
rect 859 117 860 121
rect 854 116 860 117
rect 910 121 916 122
rect 910 117 911 121
rect 915 117 916 121
rect 910 116 916 117
rect 974 121 980 122
rect 974 117 975 121
rect 979 117 980 121
rect 974 116 980 117
rect 1038 121 1044 122
rect 1038 117 1039 121
rect 1043 117 1044 121
rect 1038 116 1044 117
rect 1102 121 1108 122
rect 1102 117 1103 121
rect 1107 117 1108 121
rect 1102 116 1108 117
rect 1158 121 1164 122
rect 1158 117 1159 121
rect 1163 117 1164 121
rect 1158 116 1164 117
rect 1214 121 1220 122
rect 1214 117 1215 121
rect 1219 117 1220 121
rect 1214 116 1220 117
rect 1270 121 1276 122
rect 1328 121 1330 133
rect 1368 129 1370 141
rect 1400 130 1402 141
rect 1456 130 1458 141
rect 1512 130 1514 141
rect 1568 130 1570 141
rect 1640 130 1642 141
rect 1720 130 1722 141
rect 1800 130 1802 141
rect 1880 130 1882 141
rect 1960 130 1962 141
rect 2032 130 2034 141
rect 2104 130 2106 141
rect 2168 130 2170 141
rect 2232 130 2234 141
rect 2296 130 2298 141
rect 2360 130 2362 141
rect 2416 130 2418 141
rect 2472 130 2474 141
rect 2528 130 2530 141
rect 1398 129 1404 130
rect 1366 128 1372 129
rect 1366 124 1367 128
rect 1371 124 1372 128
rect 1398 125 1399 129
rect 1403 125 1404 129
rect 1398 124 1404 125
rect 1454 129 1460 130
rect 1454 125 1455 129
rect 1459 125 1460 129
rect 1454 124 1460 125
rect 1510 129 1516 130
rect 1510 125 1511 129
rect 1515 125 1516 129
rect 1510 124 1516 125
rect 1566 129 1572 130
rect 1566 125 1567 129
rect 1571 125 1572 129
rect 1566 124 1572 125
rect 1638 129 1644 130
rect 1638 125 1639 129
rect 1643 125 1644 129
rect 1638 124 1644 125
rect 1718 129 1724 130
rect 1718 125 1719 129
rect 1723 125 1724 129
rect 1718 124 1724 125
rect 1798 129 1804 130
rect 1798 125 1799 129
rect 1803 125 1804 129
rect 1798 124 1804 125
rect 1878 129 1884 130
rect 1878 125 1879 129
rect 1883 125 1884 129
rect 1878 124 1884 125
rect 1958 129 1964 130
rect 1958 125 1959 129
rect 1963 125 1964 129
rect 1958 124 1964 125
rect 2030 129 2036 130
rect 2030 125 2031 129
rect 2035 125 2036 129
rect 2030 124 2036 125
rect 2102 129 2108 130
rect 2102 125 2103 129
rect 2107 125 2108 129
rect 2102 124 2108 125
rect 2166 129 2172 130
rect 2166 125 2167 129
rect 2171 125 2172 129
rect 2166 124 2172 125
rect 2230 129 2236 130
rect 2230 125 2231 129
rect 2235 125 2236 129
rect 2230 124 2236 125
rect 2294 129 2300 130
rect 2294 125 2295 129
rect 2299 125 2300 129
rect 2294 124 2300 125
rect 2358 129 2364 130
rect 2358 125 2359 129
rect 2363 125 2364 129
rect 2358 124 2364 125
rect 2414 129 2420 130
rect 2414 125 2415 129
rect 2419 125 2420 129
rect 2414 124 2420 125
rect 2470 129 2476 130
rect 2470 125 2471 129
rect 2475 125 2476 129
rect 2470 124 2476 125
rect 2526 129 2532 130
rect 2584 129 2586 141
rect 2526 125 2527 129
rect 2531 125 2532 129
rect 2526 124 2532 125
rect 2582 128 2588 129
rect 2582 124 2583 128
rect 2587 124 2588 128
rect 1366 123 1372 124
rect 2582 123 2588 124
rect 1270 117 1271 121
rect 1275 117 1276 121
rect 1270 116 1276 117
rect 1326 120 1332 121
rect 1326 116 1327 120
rect 1331 116 1332 120
rect 110 115 116 116
rect 1326 115 1332 116
rect 1366 111 1372 112
rect 1366 107 1367 111
rect 1371 107 1372 111
rect 1366 106 1372 107
rect 2582 111 2588 112
rect 2582 107 2583 111
rect 2587 107 2588 111
rect 2582 106 2588 107
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 110 98 116 99
rect 1326 103 1332 104
rect 1326 99 1327 103
rect 1331 99 1332 103
rect 1326 98 1332 99
rect 112 83 114 98
rect 158 94 164 95
rect 158 90 159 94
rect 163 90 164 94
rect 158 89 164 90
rect 214 94 220 95
rect 214 90 215 94
rect 219 90 220 94
rect 214 89 220 90
rect 270 94 276 95
rect 270 90 271 94
rect 275 90 276 94
rect 270 89 276 90
rect 326 94 332 95
rect 326 90 327 94
rect 331 90 332 94
rect 326 89 332 90
rect 382 94 388 95
rect 382 90 383 94
rect 387 90 388 94
rect 382 89 388 90
rect 438 94 444 95
rect 438 90 439 94
rect 443 90 444 94
rect 438 89 444 90
rect 494 94 500 95
rect 494 90 495 94
rect 499 90 500 94
rect 494 89 500 90
rect 550 94 556 95
rect 550 90 551 94
rect 555 90 556 94
rect 550 89 556 90
rect 622 94 628 95
rect 622 90 623 94
rect 627 90 628 94
rect 622 89 628 90
rect 686 94 692 95
rect 686 90 687 94
rect 691 90 692 94
rect 686 89 692 90
rect 750 94 756 95
rect 750 90 751 94
rect 755 90 756 94
rect 750 89 756 90
rect 814 94 820 95
rect 814 90 815 94
rect 819 90 820 94
rect 814 89 820 90
rect 870 94 876 95
rect 870 90 871 94
rect 875 90 876 94
rect 870 89 876 90
rect 926 94 932 95
rect 926 90 927 94
rect 931 90 932 94
rect 926 89 932 90
rect 990 94 996 95
rect 990 90 991 94
rect 995 90 996 94
rect 990 89 996 90
rect 1054 94 1060 95
rect 1054 90 1055 94
rect 1059 90 1060 94
rect 1054 89 1060 90
rect 1118 94 1124 95
rect 1118 90 1119 94
rect 1123 90 1124 94
rect 1118 89 1124 90
rect 1174 94 1180 95
rect 1174 90 1175 94
rect 1179 90 1180 94
rect 1174 89 1180 90
rect 1230 94 1236 95
rect 1230 90 1231 94
rect 1235 90 1236 94
rect 1230 89 1236 90
rect 1286 94 1292 95
rect 1286 90 1287 94
rect 1291 90 1292 94
rect 1286 89 1292 90
rect 160 83 162 89
rect 216 83 218 89
rect 272 83 274 89
rect 328 83 330 89
rect 384 83 386 89
rect 440 83 442 89
rect 496 83 498 89
rect 552 83 554 89
rect 624 83 626 89
rect 688 83 690 89
rect 752 83 754 89
rect 816 83 818 89
rect 872 83 874 89
rect 928 83 930 89
rect 992 83 994 89
rect 1056 83 1058 89
rect 1120 83 1122 89
rect 1176 83 1178 89
rect 1232 83 1234 89
rect 1288 83 1290 89
rect 1328 83 1330 98
rect 1368 91 1370 106
rect 1414 102 1420 103
rect 1414 98 1415 102
rect 1419 98 1420 102
rect 1414 97 1420 98
rect 1470 102 1476 103
rect 1470 98 1471 102
rect 1475 98 1476 102
rect 1470 97 1476 98
rect 1526 102 1532 103
rect 1526 98 1527 102
rect 1531 98 1532 102
rect 1526 97 1532 98
rect 1582 102 1588 103
rect 1582 98 1583 102
rect 1587 98 1588 102
rect 1582 97 1588 98
rect 1654 102 1660 103
rect 1654 98 1655 102
rect 1659 98 1660 102
rect 1654 97 1660 98
rect 1734 102 1740 103
rect 1734 98 1735 102
rect 1739 98 1740 102
rect 1734 97 1740 98
rect 1814 102 1820 103
rect 1814 98 1815 102
rect 1819 98 1820 102
rect 1814 97 1820 98
rect 1894 102 1900 103
rect 1894 98 1895 102
rect 1899 98 1900 102
rect 1894 97 1900 98
rect 1974 102 1980 103
rect 1974 98 1975 102
rect 1979 98 1980 102
rect 1974 97 1980 98
rect 2046 102 2052 103
rect 2046 98 2047 102
rect 2051 98 2052 102
rect 2046 97 2052 98
rect 2118 102 2124 103
rect 2118 98 2119 102
rect 2123 98 2124 102
rect 2118 97 2124 98
rect 2182 102 2188 103
rect 2182 98 2183 102
rect 2187 98 2188 102
rect 2182 97 2188 98
rect 2246 102 2252 103
rect 2246 98 2247 102
rect 2251 98 2252 102
rect 2246 97 2252 98
rect 2310 102 2316 103
rect 2310 98 2311 102
rect 2315 98 2316 102
rect 2310 97 2316 98
rect 2374 102 2380 103
rect 2374 98 2375 102
rect 2379 98 2380 102
rect 2374 97 2380 98
rect 2430 102 2436 103
rect 2430 98 2431 102
rect 2435 98 2436 102
rect 2430 97 2436 98
rect 2486 102 2492 103
rect 2486 98 2487 102
rect 2491 98 2492 102
rect 2486 97 2492 98
rect 2542 102 2548 103
rect 2542 98 2543 102
rect 2547 98 2548 102
rect 2542 97 2548 98
rect 1416 91 1418 97
rect 1472 91 1474 97
rect 1528 91 1530 97
rect 1584 91 1586 97
rect 1656 91 1658 97
rect 1736 91 1738 97
rect 1816 91 1818 97
rect 1896 91 1898 97
rect 1976 91 1978 97
rect 2048 91 2050 97
rect 2120 91 2122 97
rect 2184 91 2186 97
rect 2248 91 2250 97
rect 2312 91 2314 97
rect 2376 91 2378 97
rect 2432 91 2434 97
rect 2488 91 2490 97
rect 2544 91 2546 97
rect 2584 91 2586 106
rect 1367 90 1371 91
rect 1367 85 1371 86
rect 1415 90 1419 91
rect 1415 85 1419 86
rect 1471 90 1475 91
rect 1471 85 1475 86
rect 1527 90 1531 91
rect 1527 85 1531 86
rect 1583 90 1587 91
rect 1583 85 1587 86
rect 1655 90 1659 91
rect 1655 85 1659 86
rect 1735 90 1739 91
rect 1735 85 1739 86
rect 1815 90 1819 91
rect 1815 85 1819 86
rect 1895 90 1899 91
rect 1895 85 1899 86
rect 1975 90 1979 91
rect 1975 85 1979 86
rect 2047 90 2051 91
rect 2047 85 2051 86
rect 2119 90 2123 91
rect 2119 85 2123 86
rect 2183 90 2187 91
rect 2183 85 2187 86
rect 2247 90 2251 91
rect 2247 85 2251 86
rect 2311 90 2315 91
rect 2311 85 2315 86
rect 2375 90 2379 91
rect 2375 85 2379 86
rect 2431 90 2435 91
rect 2431 85 2435 86
rect 2487 90 2491 91
rect 2487 85 2491 86
rect 2543 90 2547 91
rect 2543 85 2547 86
rect 2583 90 2587 91
rect 2583 85 2587 86
rect 111 82 115 83
rect 111 77 115 78
rect 159 82 163 83
rect 159 77 163 78
rect 215 82 219 83
rect 215 77 219 78
rect 271 82 275 83
rect 271 77 275 78
rect 327 82 331 83
rect 327 77 331 78
rect 383 82 387 83
rect 383 77 387 78
rect 439 82 443 83
rect 439 77 443 78
rect 495 82 499 83
rect 495 77 499 78
rect 551 82 555 83
rect 551 77 555 78
rect 623 82 627 83
rect 623 77 627 78
rect 687 82 691 83
rect 687 77 691 78
rect 751 82 755 83
rect 751 77 755 78
rect 815 82 819 83
rect 815 77 819 78
rect 871 82 875 83
rect 871 77 875 78
rect 927 82 931 83
rect 927 77 931 78
rect 991 82 995 83
rect 991 77 995 78
rect 1055 82 1059 83
rect 1055 77 1059 78
rect 1119 82 1123 83
rect 1119 77 1123 78
rect 1175 82 1179 83
rect 1175 77 1179 78
rect 1231 82 1235 83
rect 1231 77 1235 78
rect 1287 82 1291 83
rect 1287 77 1291 78
rect 1327 82 1331 83
rect 1327 77 1331 78
<< m4c >>
rect 111 2658 115 2662
rect 159 2658 163 2662
rect 215 2658 219 2662
rect 271 2658 275 2662
rect 327 2658 331 2662
rect 1327 2658 1331 2662
rect 111 2602 115 2606
rect 143 2602 147 2606
rect 199 2602 203 2606
rect 255 2602 259 2606
rect 263 2602 267 2606
rect 311 2602 315 2606
rect 343 2602 347 2606
rect 431 2602 435 2606
rect 519 2602 523 2606
rect 607 2602 611 2606
rect 687 2602 691 2606
rect 767 2602 771 2606
rect 839 2602 843 2606
rect 903 2602 907 2606
rect 967 2602 971 2606
rect 1031 2602 1035 2606
rect 1095 2602 1099 2606
rect 1159 2602 1163 2606
rect 1215 2602 1219 2606
rect 1271 2602 1275 2606
rect 1327 2602 1331 2606
rect 1367 2606 1371 2610
rect 1415 2606 1419 2610
rect 1471 2606 1475 2610
rect 1527 2606 1531 2610
rect 1583 2606 1587 2610
rect 1639 2606 1643 2610
rect 1695 2606 1699 2610
rect 2583 2606 2587 2610
rect 1367 2550 1371 2554
rect 1399 2550 1403 2554
rect 1455 2550 1459 2554
rect 1511 2550 1515 2554
rect 1567 2550 1571 2554
rect 1623 2550 1627 2554
rect 1679 2550 1683 2554
rect 1735 2550 1739 2554
rect 2583 2550 2587 2554
rect 111 2534 115 2538
rect 159 2534 163 2538
rect 215 2534 219 2538
rect 279 2534 283 2538
rect 319 2534 323 2538
rect 359 2534 363 2538
rect 431 2534 435 2538
rect 447 2534 451 2538
rect 535 2534 539 2538
rect 551 2534 555 2538
rect 623 2534 627 2538
rect 671 2534 675 2538
rect 703 2534 707 2538
rect 783 2534 787 2538
rect 791 2534 795 2538
rect 855 2534 859 2538
rect 903 2534 907 2538
rect 919 2534 923 2538
rect 983 2534 987 2538
rect 1007 2534 1011 2538
rect 1047 2534 1051 2538
rect 1103 2534 1107 2538
rect 1111 2534 1115 2538
rect 1175 2534 1179 2538
rect 1207 2534 1211 2538
rect 1231 2534 1235 2538
rect 1287 2534 1291 2538
rect 1327 2534 1331 2538
rect 1367 2490 1371 2494
rect 1415 2490 1419 2494
rect 1471 2490 1475 2494
rect 1527 2490 1531 2494
rect 1583 2490 1587 2494
rect 1639 2490 1643 2494
rect 1695 2490 1699 2494
rect 1751 2490 1755 2494
rect 2583 2490 2587 2494
rect 111 2470 115 2474
rect 143 2470 147 2474
rect 199 2470 203 2474
rect 295 2470 299 2474
rect 303 2470 307 2474
rect 407 2470 411 2474
rect 415 2470 419 2474
rect 519 2470 523 2474
rect 535 2470 539 2474
rect 639 2470 643 2474
rect 655 2470 659 2474
rect 751 2470 755 2474
rect 775 2470 779 2474
rect 855 2470 859 2474
rect 887 2470 891 2474
rect 951 2470 955 2474
rect 991 2470 995 2474
rect 1047 2470 1051 2474
rect 1087 2470 1091 2474
rect 1143 2470 1147 2474
rect 1191 2470 1195 2474
rect 1239 2470 1243 2474
rect 1271 2470 1275 2474
rect 1327 2470 1331 2474
rect 1367 2426 1371 2430
rect 1455 2426 1459 2430
rect 1479 2426 1483 2430
rect 1511 2426 1515 2430
rect 1535 2426 1539 2430
rect 1567 2426 1571 2430
rect 1591 2426 1595 2430
rect 1623 2426 1627 2430
rect 1647 2426 1651 2430
rect 1679 2426 1683 2430
rect 1703 2426 1707 2430
rect 1735 2426 1739 2430
rect 1759 2426 1763 2430
rect 2583 2426 2587 2430
rect 111 2406 115 2410
rect 159 2406 163 2410
rect 215 2406 219 2410
rect 223 2406 227 2410
rect 287 2406 291 2410
rect 311 2406 315 2410
rect 367 2406 371 2410
rect 423 2406 427 2410
rect 455 2406 459 2410
rect 535 2406 539 2410
rect 543 2406 547 2410
rect 639 2406 643 2410
rect 655 2406 659 2410
rect 727 2406 731 2410
rect 767 2406 771 2410
rect 815 2406 819 2410
rect 871 2406 875 2410
rect 895 2406 899 2410
rect 967 2406 971 2410
rect 975 2406 979 2410
rect 1055 2406 1059 2410
rect 1063 2406 1067 2410
rect 1143 2406 1147 2410
rect 1159 2406 1163 2410
rect 1255 2406 1259 2410
rect 1327 2406 1331 2410
rect 1367 2366 1371 2370
rect 1471 2366 1475 2370
rect 1495 2366 1499 2370
rect 1527 2366 1531 2370
rect 1551 2366 1555 2370
rect 1583 2366 1587 2370
rect 1607 2366 1611 2370
rect 1639 2366 1643 2370
rect 1663 2366 1667 2370
rect 1695 2366 1699 2370
rect 1719 2366 1723 2370
rect 1775 2366 1779 2370
rect 2583 2366 2587 2370
rect 111 2342 115 2346
rect 207 2342 211 2346
rect 271 2342 275 2346
rect 327 2342 331 2346
rect 351 2342 355 2346
rect 383 2342 387 2346
rect 439 2342 443 2346
rect 503 2342 507 2346
rect 527 2342 531 2346
rect 567 2342 571 2346
rect 623 2342 627 2346
rect 631 2342 635 2346
rect 695 2342 699 2346
rect 711 2342 715 2346
rect 759 2342 763 2346
rect 799 2342 803 2346
rect 823 2342 827 2346
rect 879 2342 883 2346
rect 887 2342 891 2346
rect 951 2342 955 2346
rect 959 2342 963 2346
rect 1015 2342 1019 2346
rect 1039 2342 1043 2346
rect 1127 2342 1131 2346
rect 1327 2342 1331 2346
rect 1367 2310 1371 2314
rect 1399 2310 1403 2314
rect 1455 2310 1459 2314
rect 1511 2310 1515 2314
rect 1567 2310 1571 2314
rect 1623 2310 1627 2314
rect 1679 2310 1683 2314
rect 1735 2310 1739 2314
rect 1791 2310 1795 2314
rect 1847 2310 1851 2314
rect 1903 2310 1907 2314
rect 1959 2310 1963 2314
rect 2015 2310 2019 2314
rect 2071 2310 2075 2314
rect 2127 2310 2131 2314
rect 2183 2310 2187 2314
rect 2247 2310 2251 2314
rect 2311 2310 2315 2314
rect 2375 2310 2379 2314
rect 2439 2310 2443 2314
rect 2583 2310 2587 2314
rect 111 2278 115 2282
rect 343 2278 347 2282
rect 399 2278 403 2282
rect 407 2278 411 2282
rect 455 2278 459 2282
rect 463 2278 467 2282
rect 519 2278 523 2282
rect 575 2278 579 2282
rect 583 2278 587 2282
rect 631 2278 635 2282
rect 647 2278 651 2282
rect 687 2278 691 2282
rect 711 2278 715 2282
rect 743 2278 747 2282
rect 775 2278 779 2282
rect 799 2278 803 2282
rect 839 2278 843 2282
rect 855 2278 859 2282
rect 903 2278 907 2282
rect 911 2278 915 2282
rect 967 2278 971 2282
rect 1031 2278 1035 2282
rect 1327 2278 1331 2282
rect 1367 2254 1371 2258
rect 1415 2254 1419 2258
rect 1471 2254 1475 2258
rect 1511 2254 1515 2258
rect 1527 2254 1531 2258
rect 1583 2254 1587 2258
rect 1623 2254 1627 2258
rect 1639 2254 1643 2258
rect 1695 2254 1699 2258
rect 1727 2254 1731 2258
rect 1751 2254 1755 2258
rect 1807 2254 1811 2258
rect 1823 2254 1827 2258
rect 1863 2254 1867 2258
rect 1903 2254 1907 2258
rect 1919 2254 1923 2258
rect 1975 2254 1979 2258
rect 1983 2254 1987 2258
rect 2031 2254 2035 2258
rect 2055 2254 2059 2258
rect 2087 2254 2091 2258
rect 2119 2254 2123 2258
rect 2143 2254 2147 2258
rect 2191 2254 2195 2258
rect 2199 2254 2203 2258
rect 2263 2254 2267 2258
rect 2327 2254 2331 2258
rect 2335 2254 2339 2258
rect 2391 2254 2395 2258
rect 2455 2254 2459 2258
rect 2583 2254 2587 2258
rect 111 2218 115 2222
rect 391 2218 395 2222
rect 423 2218 427 2222
rect 447 2218 451 2222
rect 479 2218 483 2222
rect 503 2218 507 2222
rect 535 2218 539 2222
rect 559 2218 563 2222
rect 591 2218 595 2222
rect 615 2218 619 2222
rect 647 2218 651 2222
rect 671 2218 675 2222
rect 711 2218 715 2222
rect 727 2218 731 2222
rect 783 2218 787 2222
rect 839 2218 843 2222
rect 855 2218 859 2222
rect 895 2218 899 2222
rect 927 2218 931 2222
rect 951 2218 955 2222
rect 999 2218 1003 2222
rect 1071 2218 1075 2222
rect 1143 2218 1147 2222
rect 1215 2218 1219 2222
rect 1271 2218 1275 2222
rect 1327 2218 1331 2222
rect 1367 2194 1371 2198
rect 1399 2194 1403 2198
rect 1495 2194 1499 2198
rect 1607 2194 1611 2198
rect 1711 2194 1715 2198
rect 1751 2194 1755 2198
rect 1807 2194 1811 2198
rect 1839 2194 1843 2198
rect 1887 2194 1891 2198
rect 1927 2194 1931 2198
rect 1967 2194 1971 2198
rect 2007 2194 2011 2198
rect 2039 2194 2043 2198
rect 2087 2194 2091 2198
rect 2103 2194 2107 2198
rect 2167 2194 2171 2198
rect 2175 2194 2179 2198
rect 2247 2194 2251 2198
rect 2319 2194 2323 2198
rect 2335 2194 2339 2198
rect 2423 2194 2427 2198
rect 2583 2194 2587 2198
rect 111 2154 115 2158
rect 199 2154 203 2158
rect 271 2154 275 2158
rect 351 2154 355 2158
rect 439 2154 443 2158
rect 447 2154 451 2158
rect 495 2154 499 2158
rect 551 2154 555 2158
rect 607 2154 611 2158
rect 663 2154 667 2158
rect 727 2154 731 2158
rect 775 2154 779 2158
rect 799 2154 803 2158
rect 871 2154 875 2158
rect 879 2154 883 2158
rect 943 2154 947 2158
rect 983 2154 987 2158
rect 1015 2154 1019 2158
rect 1079 2154 1083 2158
rect 1087 2154 1091 2158
rect 1159 2154 1163 2158
rect 1183 2154 1187 2158
rect 1231 2154 1235 2158
rect 1287 2154 1291 2158
rect 1327 2154 1331 2158
rect 1367 2138 1371 2142
rect 1607 2138 1611 2142
rect 1679 2138 1683 2142
rect 1767 2138 1771 2142
rect 1855 2138 1859 2142
rect 1863 2138 1867 2142
rect 1943 2138 1947 2142
rect 1959 2138 1963 2142
rect 2023 2138 2027 2142
rect 2063 2138 2067 2142
rect 2103 2138 2107 2142
rect 2159 2138 2163 2142
rect 2183 2138 2187 2142
rect 2255 2138 2259 2142
rect 2263 2138 2267 2142
rect 2351 2138 2355 2142
rect 2439 2138 2443 2142
rect 2447 2138 2451 2142
rect 2543 2138 2547 2142
rect 2583 2138 2587 2142
rect 111 2086 115 2090
rect 143 2086 147 2090
rect 183 2086 187 2090
rect 199 2086 203 2090
rect 255 2086 259 2090
rect 271 2086 275 2090
rect 335 2086 339 2090
rect 367 2086 371 2090
rect 431 2086 435 2090
rect 463 2086 467 2090
rect 535 2086 539 2090
rect 567 2086 571 2090
rect 647 2086 651 2090
rect 663 2086 667 2090
rect 759 2086 763 2090
rect 847 2086 851 2090
rect 863 2086 867 2090
rect 927 2086 931 2090
rect 967 2086 971 2090
rect 1007 2086 1011 2090
rect 1063 2086 1067 2090
rect 1095 2086 1099 2090
rect 1167 2086 1171 2090
rect 1183 2086 1187 2090
rect 1271 2086 1275 2090
rect 1327 2086 1331 2090
rect 1367 2082 1371 2086
rect 1487 2082 1491 2086
rect 1583 2082 1587 2086
rect 1591 2082 1595 2086
rect 1663 2082 1667 2086
rect 1679 2082 1683 2086
rect 1751 2082 1755 2086
rect 1783 2082 1787 2086
rect 1847 2082 1851 2086
rect 1887 2082 1891 2086
rect 1943 2082 1947 2086
rect 1983 2082 1987 2086
rect 2047 2082 2051 2086
rect 2079 2082 2083 2086
rect 2143 2082 2147 2086
rect 2167 2082 2171 2086
rect 2239 2082 2243 2086
rect 2255 2082 2259 2086
rect 2335 2082 2339 2086
rect 2343 2082 2347 2086
rect 2431 2082 2435 2086
rect 2439 2082 2443 2086
rect 2527 2082 2531 2086
rect 2583 2082 2587 2086
rect 111 2022 115 2026
rect 159 2022 163 2026
rect 175 2022 179 2026
rect 215 2022 219 2026
rect 239 2022 243 2026
rect 287 2022 291 2026
rect 311 2022 315 2026
rect 383 2022 387 2026
rect 391 2022 395 2026
rect 471 2022 475 2026
rect 479 2022 483 2026
rect 559 2022 563 2026
rect 583 2022 587 2026
rect 647 2022 651 2026
rect 679 2022 683 2026
rect 735 2022 739 2026
rect 775 2022 779 2026
rect 823 2022 827 2026
rect 863 2022 867 2026
rect 911 2022 915 2026
rect 943 2022 947 2026
rect 1007 2022 1011 2026
rect 1023 2022 1027 2026
rect 1103 2022 1107 2026
rect 1111 2022 1115 2026
rect 1199 2022 1203 2026
rect 1327 2022 1331 2026
rect 1367 2026 1371 2030
rect 1415 2026 1419 2030
rect 1471 2026 1475 2030
rect 1503 2026 1507 2030
rect 1535 2026 1539 2030
rect 1599 2026 1603 2030
rect 1615 2026 1619 2030
rect 1695 2026 1699 2030
rect 1703 2026 1707 2030
rect 1791 2026 1795 2030
rect 1799 2026 1803 2030
rect 1887 2026 1891 2030
rect 1903 2026 1907 2030
rect 1983 2026 1987 2030
rect 1999 2026 2003 2030
rect 2079 2026 2083 2030
rect 2095 2026 2099 2030
rect 2175 2026 2179 2030
rect 2183 2026 2187 2030
rect 2271 2026 2275 2030
rect 2359 2026 2363 2030
rect 2367 2026 2371 2030
rect 2455 2026 2459 2030
rect 2463 2026 2467 2030
rect 2543 2026 2547 2030
rect 2583 2026 2587 2030
rect 111 1966 115 1970
rect 159 1966 163 1970
rect 223 1966 227 1970
rect 295 1966 299 1970
rect 375 1966 379 1970
rect 383 1966 387 1970
rect 439 1966 443 1970
rect 455 1966 459 1970
rect 495 1966 499 1970
rect 543 1966 547 1970
rect 551 1966 555 1970
rect 607 1966 611 1970
rect 631 1966 635 1970
rect 671 1966 675 1970
rect 719 1966 723 1970
rect 735 1966 739 1970
rect 807 1966 811 1970
rect 879 1966 883 1970
rect 895 1966 899 1970
rect 951 1966 955 1970
rect 991 1966 995 1970
rect 1023 1966 1027 1970
rect 1087 1966 1091 1970
rect 1327 1966 1331 1970
rect 1367 1966 1371 1970
rect 1399 1966 1403 1970
rect 1455 1966 1459 1970
rect 1519 1966 1523 1970
rect 1599 1966 1603 1970
rect 1679 1966 1683 1970
rect 1687 1966 1691 1970
rect 1759 1966 1763 1970
rect 1775 1966 1779 1970
rect 1855 1966 1859 1970
rect 1871 1966 1875 1970
rect 1967 1966 1971 1970
rect 2063 1966 2067 1970
rect 2095 1966 2099 1970
rect 2159 1966 2163 1970
rect 2239 1966 2243 1970
rect 2255 1966 2259 1970
rect 2351 1966 2355 1970
rect 2391 1966 2395 1970
rect 2447 1966 2451 1970
rect 2527 1966 2531 1970
rect 2583 1966 2587 1970
rect 111 1910 115 1914
rect 399 1910 403 1914
rect 455 1910 459 1914
rect 511 1910 515 1914
rect 519 1910 523 1914
rect 567 1910 571 1914
rect 575 1910 579 1914
rect 623 1910 627 1914
rect 631 1910 635 1914
rect 687 1910 691 1914
rect 743 1910 747 1914
rect 751 1910 755 1914
rect 807 1910 811 1914
rect 823 1910 827 1914
rect 871 1910 875 1914
rect 895 1910 899 1914
rect 935 1910 939 1914
rect 967 1910 971 1914
rect 999 1910 1003 1914
rect 1039 1910 1043 1914
rect 1327 1910 1331 1914
rect 1367 1910 1371 1914
rect 1415 1910 1419 1914
rect 1471 1910 1475 1914
rect 1535 1910 1539 1914
rect 1575 1910 1579 1914
rect 1615 1910 1619 1914
rect 1631 1910 1635 1914
rect 1687 1910 1691 1914
rect 1695 1910 1699 1914
rect 1743 1910 1747 1914
rect 1775 1910 1779 1914
rect 1799 1910 1803 1914
rect 1855 1910 1859 1914
rect 1871 1910 1875 1914
rect 1927 1910 1931 1914
rect 1983 1910 1987 1914
rect 2015 1910 2019 1914
rect 2111 1910 2115 1914
rect 2127 1910 2131 1914
rect 2247 1910 2251 1914
rect 2255 1910 2259 1914
rect 2383 1910 2387 1914
rect 2407 1910 2411 1914
rect 2519 1910 2523 1914
rect 2543 1910 2547 1914
rect 2583 1910 2587 1914
rect 111 1850 115 1854
rect 143 1850 147 1854
rect 199 1850 203 1854
rect 255 1850 259 1854
rect 311 1850 315 1854
rect 375 1850 379 1854
rect 455 1850 459 1854
rect 503 1850 507 1854
rect 543 1850 547 1854
rect 559 1850 563 1854
rect 615 1850 619 1854
rect 631 1850 635 1854
rect 671 1850 675 1854
rect 719 1850 723 1854
rect 727 1850 731 1854
rect 791 1850 795 1854
rect 799 1850 803 1854
rect 855 1850 859 1854
rect 887 1850 891 1854
rect 919 1850 923 1854
rect 975 1850 979 1854
rect 983 1850 987 1854
rect 1063 1850 1067 1854
rect 1327 1850 1331 1854
rect 1367 1846 1371 1850
rect 1559 1846 1563 1850
rect 1615 1846 1619 1850
rect 1623 1846 1627 1850
rect 1671 1846 1675 1850
rect 1679 1846 1683 1850
rect 1727 1846 1731 1850
rect 1735 1846 1739 1850
rect 1783 1846 1787 1850
rect 1791 1846 1795 1850
rect 1839 1846 1843 1850
rect 1847 1846 1851 1850
rect 1903 1846 1907 1850
rect 1911 1846 1915 1850
rect 1967 1846 1971 1850
rect 1999 1846 2003 1850
rect 2039 1846 2043 1850
rect 2111 1846 2115 1850
rect 2127 1846 2131 1850
rect 2223 1846 2227 1850
rect 2231 1846 2235 1850
rect 2327 1846 2331 1850
rect 2367 1846 2371 1850
rect 2439 1846 2443 1850
rect 2503 1846 2507 1850
rect 2527 1846 2531 1850
rect 2583 1846 2587 1850
rect 111 1786 115 1790
rect 159 1786 163 1790
rect 215 1786 219 1790
rect 255 1786 259 1790
rect 271 1786 275 1790
rect 327 1786 331 1790
rect 375 1786 379 1790
rect 391 1786 395 1790
rect 471 1786 475 1790
rect 503 1786 507 1790
rect 559 1786 563 1790
rect 623 1786 627 1790
rect 647 1786 651 1790
rect 735 1786 739 1790
rect 743 1786 747 1790
rect 815 1786 819 1790
rect 855 1786 859 1790
rect 903 1786 907 1790
rect 959 1786 963 1790
rect 991 1786 995 1790
rect 1055 1786 1059 1790
rect 1079 1786 1083 1790
rect 1151 1786 1155 1790
rect 1247 1786 1251 1790
rect 1327 1786 1331 1790
rect 1367 1782 1371 1786
rect 1471 1782 1475 1786
rect 1535 1782 1539 1786
rect 1615 1782 1619 1786
rect 1639 1782 1643 1786
rect 1695 1782 1699 1786
rect 1751 1782 1755 1786
rect 1783 1782 1787 1786
rect 1807 1782 1811 1786
rect 1863 1782 1867 1786
rect 1879 1782 1883 1786
rect 1919 1782 1923 1786
rect 1975 1782 1979 1786
rect 1983 1782 1987 1786
rect 2055 1782 2059 1786
rect 2071 1782 2075 1786
rect 2143 1782 2147 1786
rect 2167 1782 2171 1786
rect 2239 1782 2243 1786
rect 2263 1782 2267 1786
rect 2343 1782 2347 1786
rect 2359 1782 2363 1786
rect 2455 1782 2459 1786
rect 2463 1782 2467 1786
rect 2543 1782 2547 1786
rect 2583 1782 2587 1786
rect 111 1730 115 1734
rect 143 1730 147 1734
rect 239 1730 243 1734
rect 263 1730 267 1734
rect 359 1730 363 1734
rect 415 1730 419 1734
rect 487 1730 491 1734
rect 567 1730 571 1734
rect 607 1730 611 1734
rect 711 1730 715 1734
rect 727 1730 731 1734
rect 839 1730 843 1734
rect 855 1730 859 1734
rect 943 1730 947 1734
rect 999 1730 1003 1734
rect 1039 1730 1043 1734
rect 1135 1730 1139 1734
rect 1143 1730 1147 1734
rect 1231 1730 1235 1734
rect 1271 1730 1275 1734
rect 1327 1730 1331 1734
rect 1367 1722 1371 1726
rect 1399 1722 1403 1726
rect 1455 1722 1459 1726
rect 1479 1722 1483 1726
rect 1519 1722 1523 1726
rect 1599 1722 1603 1726
rect 1679 1722 1683 1726
rect 1719 1722 1723 1726
rect 1767 1722 1771 1726
rect 1839 1722 1843 1726
rect 1863 1722 1867 1726
rect 1951 1722 1955 1726
rect 1959 1722 1963 1726
rect 2055 1722 2059 1726
rect 2151 1722 2155 1726
rect 2159 1722 2163 1726
rect 2247 1722 2251 1726
rect 2255 1722 2259 1726
rect 2343 1722 2347 1726
rect 2351 1722 2355 1726
rect 2447 1722 2451 1726
rect 2527 1722 2531 1726
rect 2583 1722 2587 1726
rect 111 1670 115 1674
rect 159 1670 163 1674
rect 223 1670 227 1674
rect 279 1670 283 1674
rect 303 1670 307 1674
rect 383 1670 387 1674
rect 431 1670 435 1674
rect 463 1670 467 1674
rect 535 1670 539 1674
rect 583 1670 587 1674
rect 607 1670 611 1674
rect 679 1670 683 1674
rect 727 1670 731 1674
rect 767 1670 771 1674
rect 863 1670 867 1674
rect 871 1670 875 1674
rect 967 1670 971 1674
rect 1015 1670 1019 1674
rect 1079 1670 1083 1674
rect 1159 1670 1163 1674
rect 1191 1670 1195 1674
rect 1287 1670 1291 1674
rect 1327 1670 1331 1674
rect 1367 1666 1371 1670
rect 1415 1666 1419 1670
rect 1495 1666 1499 1670
rect 1503 1666 1507 1670
rect 1615 1666 1619 1670
rect 1623 1666 1627 1670
rect 1735 1666 1739 1670
rect 1751 1666 1755 1670
rect 1855 1666 1859 1670
rect 1879 1666 1883 1670
rect 1967 1666 1971 1670
rect 1999 1666 2003 1670
rect 2071 1666 2075 1670
rect 2119 1666 2123 1670
rect 2175 1666 2179 1670
rect 2231 1666 2235 1670
rect 2271 1666 2275 1670
rect 2343 1666 2347 1670
rect 2367 1666 2371 1670
rect 2455 1666 2459 1670
rect 2463 1666 2467 1670
rect 2543 1666 2547 1670
rect 2583 1666 2587 1670
rect 111 1614 115 1618
rect 143 1614 147 1618
rect 207 1614 211 1618
rect 247 1614 251 1618
rect 287 1614 291 1618
rect 367 1614 371 1618
rect 447 1614 451 1618
rect 479 1614 483 1618
rect 519 1614 523 1618
rect 575 1614 579 1618
rect 591 1614 595 1618
rect 663 1614 667 1618
rect 671 1614 675 1618
rect 751 1614 755 1618
rect 767 1614 771 1618
rect 847 1614 851 1618
rect 863 1614 867 1618
rect 951 1614 955 1618
rect 959 1614 963 1618
rect 1063 1614 1067 1618
rect 1175 1614 1179 1618
rect 1271 1614 1275 1618
rect 1327 1614 1331 1618
rect 1367 1598 1371 1602
rect 1399 1598 1403 1602
rect 1487 1598 1491 1602
rect 1495 1598 1499 1602
rect 1607 1598 1611 1602
rect 1615 1598 1619 1602
rect 1735 1598 1739 1602
rect 1743 1598 1747 1602
rect 1863 1598 1867 1602
rect 1983 1598 1987 1602
rect 2095 1598 2099 1602
rect 2103 1598 2107 1602
rect 2199 1598 2203 1602
rect 2215 1598 2219 1602
rect 2295 1598 2299 1602
rect 2327 1598 2331 1602
rect 2391 1598 2395 1602
rect 2439 1598 2443 1602
rect 2495 1598 2499 1602
rect 2527 1598 2531 1602
rect 2583 1598 2587 1602
rect 111 1554 115 1558
rect 159 1554 163 1558
rect 231 1554 235 1558
rect 263 1554 267 1558
rect 335 1554 339 1558
rect 383 1554 387 1558
rect 455 1554 459 1558
rect 495 1554 499 1558
rect 583 1554 587 1558
rect 591 1554 595 1558
rect 687 1554 691 1558
rect 719 1554 723 1558
rect 783 1554 787 1558
rect 863 1554 867 1558
rect 879 1554 883 1558
rect 975 1554 979 1558
rect 1007 1554 1011 1558
rect 1079 1554 1083 1558
rect 1151 1554 1155 1558
rect 1191 1554 1195 1558
rect 1287 1554 1291 1558
rect 1327 1554 1331 1558
rect 1367 1538 1371 1542
rect 1415 1538 1419 1542
rect 1511 1538 1515 1542
rect 1527 1538 1531 1542
rect 1631 1538 1635 1542
rect 1647 1538 1651 1542
rect 1759 1538 1763 1542
rect 1767 1538 1771 1542
rect 1879 1538 1883 1542
rect 1983 1538 1987 1542
rect 1999 1538 2003 1542
rect 2079 1538 2083 1542
rect 2111 1538 2115 1542
rect 2167 1538 2171 1542
rect 2215 1538 2219 1542
rect 2255 1538 2259 1542
rect 2311 1538 2315 1542
rect 2335 1538 2339 1542
rect 2407 1538 2411 1542
rect 2487 1538 2491 1542
rect 2511 1538 2515 1542
rect 2543 1538 2547 1542
rect 2583 1538 2587 1542
rect 111 1498 115 1502
rect 143 1498 147 1502
rect 199 1498 203 1502
rect 215 1498 219 1502
rect 271 1498 275 1502
rect 319 1498 323 1502
rect 367 1498 371 1502
rect 439 1498 443 1502
rect 479 1498 483 1502
rect 567 1498 571 1502
rect 591 1498 595 1502
rect 703 1498 707 1502
rect 807 1498 811 1502
rect 847 1498 851 1502
rect 911 1498 915 1502
rect 991 1498 995 1502
rect 1007 1498 1011 1502
rect 1103 1498 1107 1502
rect 1135 1498 1139 1502
rect 1199 1498 1203 1502
rect 1271 1498 1275 1502
rect 1327 1498 1331 1502
rect 1367 1474 1371 1478
rect 1399 1474 1403 1478
rect 1503 1474 1507 1478
rect 1511 1474 1515 1478
rect 1631 1474 1635 1478
rect 1751 1474 1755 1478
rect 1863 1474 1867 1478
rect 1871 1474 1875 1478
rect 1967 1474 1971 1478
rect 1983 1474 1987 1478
rect 2063 1474 2067 1478
rect 2087 1474 2091 1478
rect 2151 1474 2155 1478
rect 2183 1474 2187 1478
rect 2239 1474 2243 1478
rect 2271 1474 2275 1478
rect 2319 1474 2323 1478
rect 2359 1474 2363 1478
rect 2391 1474 2395 1478
rect 2455 1474 2459 1478
rect 2471 1474 2475 1478
rect 2527 1474 2531 1478
rect 2583 1474 2587 1478
rect 111 1438 115 1442
rect 159 1438 163 1442
rect 215 1438 219 1442
rect 255 1438 259 1442
rect 287 1438 291 1442
rect 311 1438 315 1442
rect 375 1438 379 1442
rect 383 1438 387 1442
rect 447 1438 451 1442
rect 495 1438 499 1442
rect 527 1438 531 1442
rect 607 1438 611 1442
rect 695 1438 699 1442
rect 719 1438 723 1442
rect 783 1438 787 1442
rect 823 1438 827 1442
rect 871 1438 875 1442
rect 927 1438 931 1442
rect 959 1438 963 1442
rect 1023 1438 1027 1442
rect 1055 1438 1059 1442
rect 1119 1438 1123 1442
rect 1151 1438 1155 1442
rect 1215 1438 1219 1442
rect 1287 1438 1291 1442
rect 1327 1438 1331 1442
rect 1367 1414 1371 1418
rect 1415 1414 1419 1418
rect 1471 1414 1475 1418
rect 1519 1414 1523 1418
rect 1551 1414 1555 1418
rect 1631 1414 1635 1418
rect 1647 1414 1651 1418
rect 1711 1414 1715 1418
rect 1767 1414 1771 1418
rect 1791 1414 1795 1418
rect 1871 1414 1875 1418
rect 1887 1414 1891 1418
rect 1959 1414 1963 1418
rect 1999 1414 2003 1418
rect 2055 1414 2059 1418
rect 2103 1414 2107 1418
rect 2167 1414 2171 1418
rect 2199 1414 2203 1418
rect 2287 1414 2291 1418
rect 2295 1414 2299 1418
rect 2375 1414 2379 1418
rect 2431 1414 2435 1418
rect 2471 1414 2475 1418
rect 2543 1414 2547 1418
rect 2583 1414 2587 1418
rect 111 1374 115 1378
rect 239 1374 243 1378
rect 295 1374 299 1378
rect 359 1374 363 1378
rect 415 1374 419 1378
rect 431 1374 435 1378
rect 471 1374 475 1378
rect 511 1374 515 1378
rect 527 1374 531 1378
rect 591 1374 595 1378
rect 671 1374 675 1378
rect 679 1374 683 1378
rect 751 1374 755 1378
rect 767 1374 771 1378
rect 839 1374 843 1378
rect 855 1374 859 1378
rect 935 1374 939 1378
rect 943 1374 947 1378
rect 1031 1374 1035 1378
rect 1039 1374 1043 1378
rect 1127 1374 1131 1378
rect 1135 1374 1139 1378
rect 1231 1374 1235 1378
rect 1327 1374 1331 1378
rect 1367 1358 1371 1362
rect 1399 1358 1403 1362
rect 1423 1358 1427 1362
rect 1455 1358 1459 1362
rect 1495 1358 1499 1362
rect 1535 1358 1539 1362
rect 1575 1358 1579 1362
rect 1615 1358 1619 1362
rect 1655 1358 1659 1362
rect 1695 1358 1699 1362
rect 1759 1358 1763 1362
rect 1775 1358 1779 1362
rect 1855 1358 1859 1362
rect 1879 1358 1883 1362
rect 1943 1358 1947 1362
rect 2023 1358 2027 1362
rect 2039 1358 2043 1362
rect 2151 1358 2155 1362
rect 2183 1358 2187 1362
rect 2279 1358 2283 1362
rect 2359 1358 2363 1362
rect 2415 1358 2419 1362
rect 2527 1358 2531 1362
rect 2583 1358 2587 1362
rect 111 1310 115 1314
rect 375 1310 379 1314
rect 431 1310 435 1314
rect 471 1310 475 1314
rect 487 1310 491 1314
rect 527 1310 531 1314
rect 543 1310 547 1314
rect 583 1310 587 1314
rect 607 1310 611 1314
rect 647 1310 651 1314
rect 687 1310 691 1314
rect 727 1310 731 1314
rect 767 1310 771 1314
rect 807 1310 811 1314
rect 855 1310 859 1314
rect 895 1310 899 1314
rect 951 1310 955 1314
rect 991 1310 995 1314
rect 1047 1310 1051 1314
rect 1095 1310 1099 1314
rect 1143 1310 1147 1314
rect 1199 1310 1203 1314
rect 1247 1310 1251 1314
rect 1287 1310 1291 1314
rect 1327 1310 1331 1314
rect 1367 1302 1371 1306
rect 1431 1302 1435 1306
rect 1439 1302 1443 1306
rect 1495 1302 1499 1306
rect 1511 1302 1515 1306
rect 1559 1302 1563 1306
rect 1591 1302 1595 1306
rect 1631 1302 1635 1306
rect 1671 1302 1675 1306
rect 1703 1302 1707 1306
rect 1775 1302 1779 1306
rect 1855 1302 1859 1306
rect 1895 1302 1899 1306
rect 1943 1302 1947 1306
rect 2039 1302 2043 1306
rect 2047 1302 2051 1306
rect 2159 1302 2163 1306
rect 2199 1302 2203 1306
rect 2287 1302 2291 1306
rect 2375 1302 2379 1306
rect 2423 1302 2427 1306
rect 2543 1302 2547 1306
rect 2583 1302 2587 1306
rect 111 1250 115 1254
rect 383 1250 387 1254
rect 439 1250 443 1254
rect 455 1250 459 1254
rect 503 1250 507 1254
rect 511 1250 515 1254
rect 567 1250 571 1254
rect 575 1250 579 1254
rect 631 1250 635 1254
rect 647 1250 651 1254
rect 711 1250 715 1254
rect 727 1250 731 1254
rect 791 1250 795 1254
rect 815 1250 819 1254
rect 879 1250 883 1254
rect 903 1250 907 1254
rect 975 1250 979 1254
rect 991 1250 995 1254
rect 1079 1250 1083 1254
rect 1175 1250 1179 1254
rect 1183 1250 1187 1254
rect 1271 1250 1275 1254
rect 1327 1250 1331 1254
rect 1367 1242 1371 1246
rect 1399 1242 1403 1246
rect 1415 1242 1419 1246
rect 1455 1242 1459 1246
rect 1479 1242 1483 1246
rect 1535 1242 1539 1246
rect 1543 1242 1547 1246
rect 1615 1242 1619 1246
rect 1687 1242 1691 1246
rect 1695 1242 1699 1246
rect 1759 1242 1763 1246
rect 1775 1242 1779 1246
rect 1839 1242 1843 1246
rect 1855 1242 1859 1246
rect 1927 1242 1931 1246
rect 1943 1242 1947 1246
rect 2031 1242 2035 1246
rect 2039 1242 2043 1246
rect 2143 1242 2147 1246
rect 2151 1242 2155 1246
rect 2271 1242 2275 1246
rect 2279 1242 2283 1246
rect 2407 1242 2411 1246
rect 2415 1242 2419 1246
rect 2527 1242 2531 1246
rect 2583 1242 2587 1246
rect 111 1190 115 1194
rect 279 1190 283 1194
rect 343 1190 347 1194
rect 399 1190 403 1194
rect 415 1190 419 1194
rect 455 1190 459 1194
rect 495 1190 499 1194
rect 519 1190 523 1194
rect 583 1190 587 1194
rect 591 1190 595 1194
rect 663 1190 667 1194
rect 671 1190 675 1194
rect 743 1190 747 1194
rect 759 1190 763 1194
rect 831 1190 835 1194
rect 847 1190 851 1194
rect 919 1190 923 1194
rect 935 1190 939 1194
rect 1007 1190 1011 1194
rect 1015 1190 1019 1194
rect 1087 1190 1091 1194
rect 1095 1190 1099 1194
rect 1159 1190 1163 1194
rect 1191 1190 1195 1194
rect 1231 1190 1235 1194
rect 1287 1190 1291 1194
rect 1327 1190 1331 1194
rect 1367 1178 1371 1182
rect 1415 1178 1419 1182
rect 1471 1178 1475 1182
rect 1551 1178 1555 1182
rect 1631 1178 1635 1182
rect 1695 1178 1699 1182
rect 1711 1178 1715 1182
rect 1767 1178 1771 1182
rect 1791 1178 1795 1182
rect 1847 1178 1851 1182
rect 1871 1178 1875 1182
rect 1919 1178 1923 1182
rect 1959 1178 1963 1182
rect 1991 1178 1995 1182
rect 2055 1178 2059 1182
rect 2063 1178 2067 1182
rect 2135 1178 2139 1182
rect 2167 1178 2171 1182
rect 2207 1178 2211 1182
rect 2287 1178 2291 1182
rect 2295 1178 2299 1182
rect 2367 1178 2371 1182
rect 2431 1178 2435 1182
rect 2543 1178 2547 1182
rect 2583 1178 2587 1182
rect 111 1126 115 1130
rect 143 1126 147 1130
rect 207 1126 211 1130
rect 263 1126 267 1130
rect 271 1126 275 1130
rect 327 1126 331 1130
rect 343 1126 347 1130
rect 399 1126 403 1130
rect 423 1126 427 1130
rect 479 1126 483 1130
rect 503 1126 507 1130
rect 567 1126 571 1130
rect 583 1126 587 1130
rect 655 1126 659 1130
rect 663 1126 667 1130
rect 743 1126 747 1130
rect 831 1126 835 1130
rect 919 1126 923 1130
rect 999 1126 1003 1130
rect 1007 1126 1011 1130
rect 1071 1126 1075 1130
rect 1143 1126 1147 1130
rect 1215 1126 1219 1130
rect 1271 1126 1275 1130
rect 1327 1126 1331 1130
rect 1367 1122 1371 1126
rect 1399 1122 1403 1126
rect 1479 1122 1483 1126
rect 1583 1122 1587 1126
rect 1679 1122 1683 1126
rect 1687 1122 1691 1126
rect 1751 1122 1755 1126
rect 1783 1122 1787 1126
rect 1831 1122 1835 1126
rect 1879 1122 1883 1126
rect 1903 1122 1907 1126
rect 1975 1122 1979 1126
rect 2047 1122 2051 1126
rect 2063 1122 2067 1126
rect 2119 1122 2123 1126
rect 2151 1122 2155 1126
rect 2191 1122 2195 1126
rect 2239 1122 2243 1126
rect 2271 1122 2275 1126
rect 2327 1122 2331 1126
rect 2351 1122 2355 1126
rect 2415 1122 2419 1126
rect 2583 1122 2587 1126
rect 111 1066 115 1070
rect 159 1066 163 1070
rect 215 1066 219 1070
rect 223 1066 227 1070
rect 287 1066 291 1070
rect 359 1066 363 1070
rect 383 1066 387 1070
rect 439 1066 443 1070
rect 479 1066 483 1070
rect 519 1066 523 1070
rect 583 1066 587 1070
rect 599 1066 603 1070
rect 679 1066 683 1070
rect 687 1066 691 1070
rect 759 1066 763 1070
rect 783 1066 787 1070
rect 847 1066 851 1070
rect 879 1066 883 1070
rect 935 1066 939 1070
rect 967 1066 971 1070
rect 1023 1066 1027 1070
rect 1063 1066 1067 1070
rect 1159 1066 1163 1070
rect 1327 1066 1331 1070
rect 1367 1066 1371 1070
rect 1415 1066 1419 1070
rect 1495 1066 1499 1070
rect 1511 1066 1515 1070
rect 1599 1066 1603 1070
rect 1631 1066 1635 1070
rect 1703 1066 1707 1070
rect 1751 1066 1755 1070
rect 1799 1066 1803 1070
rect 1871 1066 1875 1070
rect 1895 1066 1899 1070
rect 1991 1066 1995 1070
rect 2079 1066 2083 1070
rect 2103 1066 2107 1070
rect 2167 1066 2171 1070
rect 2199 1066 2203 1070
rect 2255 1066 2259 1070
rect 2295 1066 2299 1070
rect 2343 1066 2347 1070
rect 2383 1066 2387 1070
rect 2431 1066 2435 1070
rect 2471 1066 2475 1070
rect 2543 1066 2547 1070
rect 2583 1066 2587 1070
rect 111 1006 115 1010
rect 143 1006 147 1010
rect 199 1006 203 1010
rect 271 1006 275 1010
rect 279 1006 283 1010
rect 367 1006 371 1010
rect 383 1006 387 1010
rect 463 1006 467 1010
rect 495 1006 499 1010
rect 567 1006 571 1010
rect 615 1006 619 1010
rect 671 1006 675 1010
rect 727 1006 731 1010
rect 767 1006 771 1010
rect 839 1006 843 1010
rect 863 1006 867 1010
rect 951 1006 955 1010
rect 1047 1006 1051 1010
rect 1055 1006 1059 1010
rect 1143 1006 1147 1010
rect 1159 1006 1163 1010
rect 1271 1006 1275 1010
rect 1327 1006 1331 1010
rect 1367 1006 1371 1010
rect 1399 1006 1403 1010
rect 1487 1006 1491 1010
rect 1495 1006 1499 1010
rect 1583 1006 1587 1010
rect 1615 1006 1619 1010
rect 1695 1006 1699 1010
rect 1735 1006 1739 1010
rect 1807 1006 1811 1010
rect 1855 1006 1859 1010
rect 1919 1006 1923 1010
rect 1975 1006 1979 1010
rect 2023 1006 2027 1010
rect 2087 1006 2091 1010
rect 2119 1006 2123 1010
rect 2183 1006 2187 1010
rect 2215 1006 2219 1010
rect 2279 1006 2283 1010
rect 2303 1006 2307 1010
rect 2367 1006 2371 1010
rect 2383 1006 2387 1010
rect 2455 1006 2459 1010
rect 2463 1006 2467 1010
rect 2527 1006 2531 1010
rect 2583 1006 2587 1010
rect 111 942 115 946
rect 159 942 163 946
rect 215 942 219 946
rect 287 942 291 946
rect 295 942 299 946
rect 375 942 379 946
rect 399 942 403 946
rect 471 942 475 946
rect 511 942 515 946
rect 567 942 571 946
rect 631 942 635 946
rect 671 942 675 946
rect 743 942 747 946
rect 767 942 771 946
rect 855 942 859 946
rect 863 942 867 946
rect 959 942 963 946
rect 967 942 971 946
rect 1047 942 1051 946
rect 1071 942 1075 946
rect 1135 942 1139 946
rect 1175 942 1179 946
rect 1223 942 1227 946
rect 1287 942 1291 946
rect 1327 942 1331 946
rect 1367 942 1371 946
rect 1415 942 1419 946
rect 1503 942 1507 946
rect 1535 942 1539 946
rect 1599 942 1603 946
rect 1671 942 1675 946
rect 1711 942 1715 946
rect 1807 942 1811 946
rect 1823 942 1827 946
rect 1935 942 1939 946
rect 2039 942 2043 946
rect 2055 942 2059 946
rect 2135 942 2139 946
rect 2167 942 2171 946
rect 2231 942 2235 946
rect 2271 942 2275 946
rect 2319 942 2323 946
rect 2367 942 2371 946
rect 2399 942 2403 946
rect 2463 942 2467 946
rect 2479 942 2483 946
rect 2543 942 2547 946
rect 2583 942 2587 946
rect 111 882 115 886
rect 143 882 147 886
rect 183 882 187 886
rect 199 882 203 886
rect 239 882 243 886
rect 271 882 275 886
rect 303 882 307 886
rect 359 882 363 886
rect 375 882 379 886
rect 455 882 459 886
rect 543 882 547 886
rect 551 882 555 886
rect 639 882 643 886
rect 655 882 659 886
rect 743 882 747 886
rect 751 882 755 886
rect 847 882 851 886
rect 855 882 859 886
rect 943 882 947 886
rect 967 882 971 886
rect 1031 882 1035 886
rect 1087 882 1091 886
rect 1119 882 1123 886
rect 1207 882 1211 886
rect 1215 882 1219 886
rect 1271 882 1275 886
rect 1327 882 1331 886
rect 1367 882 1371 886
rect 1399 882 1403 886
rect 1455 882 1459 886
rect 1519 882 1523 886
rect 1607 882 1611 886
rect 1655 882 1659 886
rect 1695 882 1699 886
rect 1791 882 1795 886
rect 1895 882 1899 886
rect 1919 882 1923 886
rect 1999 882 2003 886
rect 2039 882 2043 886
rect 2103 882 2107 886
rect 2151 882 2155 886
rect 2207 882 2211 886
rect 2255 882 2259 886
rect 2311 882 2315 886
rect 2351 882 2355 886
rect 2423 882 2427 886
rect 2447 882 2451 886
rect 2527 882 2531 886
rect 2583 882 2587 886
rect 111 818 115 822
rect 199 818 203 822
rect 255 818 259 822
rect 319 818 323 822
rect 383 818 387 822
rect 391 818 395 822
rect 439 818 443 822
rect 471 818 475 822
rect 495 818 499 822
rect 559 818 563 822
rect 631 818 635 822
rect 655 818 659 822
rect 703 818 707 822
rect 759 818 763 822
rect 783 818 787 822
rect 871 818 875 822
rect 959 818 963 822
rect 983 818 987 822
rect 1047 818 1051 822
rect 1103 818 1107 822
rect 1135 818 1139 822
rect 1223 818 1227 822
rect 1231 818 1235 822
rect 1327 818 1331 822
rect 1367 822 1371 826
rect 1415 822 1419 826
rect 1471 822 1475 826
rect 1527 822 1531 826
rect 1535 822 1539 826
rect 1583 822 1587 826
rect 1623 822 1627 826
rect 1639 822 1643 826
rect 1695 822 1699 826
rect 1711 822 1715 826
rect 1751 822 1755 826
rect 1807 822 1811 826
rect 1879 822 1883 826
rect 1911 822 1915 826
rect 1959 822 1963 826
rect 2015 822 2019 826
rect 2055 822 2059 826
rect 2119 822 2123 826
rect 2167 822 2171 826
rect 2223 822 2227 826
rect 2295 822 2299 826
rect 2327 822 2331 826
rect 2431 822 2435 826
rect 2439 822 2443 826
rect 2543 822 2547 826
rect 2583 822 2587 826
rect 111 762 115 766
rect 367 762 371 766
rect 383 762 387 766
rect 423 762 427 766
rect 439 762 443 766
rect 479 762 483 766
rect 495 762 499 766
rect 543 762 547 766
rect 559 762 563 766
rect 615 762 619 766
rect 631 762 635 766
rect 687 762 691 766
rect 711 762 715 766
rect 767 762 771 766
rect 791 762 795 766
rect 855 762 859 766
rect 871 762 875 766
rect 943 762 947 766
rect 951 762 955 766
rect 1031 762 1035 766
rect 1039 762 1043 766
rect 1119 762 1123 766
rect 1127 762 1131 766
rect 1207 762 1211 766
rect 1327 762 1331 766
rect 1367 758 1371 762
rect 1511 758 1515 762
rect 1567 758 1571 762
rect 1623 758 1627 762
rect 1647 758 1651 762
rect 1679 758 1683 762
rect 1703 758 1707 762
rect 1735 758 1739 762
rect 1759 758 1763 762
rect 1791 758 1795 762
rect 1815 758 1819 762
rect 1863 758 1867 762
rect 1871 758 1875 762
rect 1927 758 1931 762
rect 1943 758 1947 762
rect 1991 758 1995 762
rect 2039 758 2043 762
rect 2063 758 2067 762
rect 2143 758 2147 762
rect 2151 758 2155 762
rect 2231 758 2235 762
rect 2279 758 2283 762
rect 2335 758 2339 762
rect 2415 758 2419 762
rect 2439 758 2443 762
rect 2527 758 2531 762
rect 2583 758 2587 762
rect 111 706 115 710
rect 343 706 347 710
rect 399 706 403 710
rect 415 706 419 710
rect 455 706 459 710
rect 487 706 491 710
rect 511 706 515 710
rect 559 706 563 710
rect 575 706 579 710
rect 631 706 635 710
rect 647 706 651 710
rect 695 706 699 710
rect 727 706 731 710
rect 759 706 763 710
rect 807 706 811 710
rect 823 706 827 710
rect 887 706 891 710
rect 951 706 955 710
rect 967 706 971 710
rect 1023 706 1027 710
rect 1055 706 1059 710
rect 1143 706 1147 710
rect 1327 706 1331 710
rect 1367 698 1371 702
rect 1663 698 1667 702
rect 1719 698 1723 702
rect 1735 698 1739 702
rect 1775 698 1779 702
rect 1791 698 1795 702
rect 1831 698 1835 702
rect 1855 698 1859 702
rect 1887 698 1891 702
rect 1919 698 1923 702
rect 1943 698 1947 702
rect 1991 698 1995 702
rect 2007 698 2011 702
rect 2063 698 2067 702
rect 2079 698 2083 702
rect 2127 698 2131 702
rect 2159 698 2163 702
rect 2199 698 2203 702
rect 2247 698 2251 702
rect 2271 698 2275 702
rect 2343 698 2347 702
rect 2351 698 2355 702
rect 2415 698 2419 702
rect 2455 698 2459 702
rect 2487 698 2491 702
rect 2543 698 2547 702
rect 2583 698 2587 702
rect 111 646 115 650
rect 231 646 235 650
rect 295 646 299 650
rect 327 646 331 650
rect 359 646 363 650
rect 399 646 403 650
rect 423 646 427 650
rect 471 646 475 650
rect 479 646 483 650
rect 535 646 539 650
rect 543 646 547 650
rect 599 646 603 650
rect 615 646 619 650
rect 663 646 667 650
rect 679 646 683 650
rect 727 646 731 650
rect 743 646 747 650
rect 791 646 795 650
rect 807 646 811 650
rect 855 646 859 650
rect 871 646 875 650
rect 919 646 923 650
rect 935 646 939 650
rect 1007 646 1011 650
rect 1327 646 1331 650
rect 1367 638 1371 642
rect 1615 638 1619 642
rect 1679 638 1683 642
rect 1719 638 1723 642
rect 1759 638 1763 642
rect 1775 638 1779 642
rect 1839 638 1843 642
rect 1903 638 1907 642
rect 1927 638 1931 642
rect 1975 638 1979 642
rect 2015 638 2019 642
rect 2047 638 2051 642
rect 2095 638 2099 642
rect 2111 638 2115 642
rect 2175 638 2179 642
rect 2183 638 2187 642
rect 2255 638 2259 642
rect 2327 638 2331 642
rect 2399 638 2403 642
rect 2471 638 2475 642
rect 2527 638 2531 642
rect 2583 638 2587 642
rect 111 582 115 586
rect 191 582 195 586
rect 247 582 251 586
rect 279 582 283 586
rect 311 582 315 586
rect 367 582 371 586
rect 375 582 379 586
rect 439 582 443 586
rect 463 582 467 586
rect 495 582 499 586
rect 551 582 555 586
rect 559 582 563 586
rect 615 582 619 586
rect 647 582 651 586
rect 679 582 683 586
rect 735 582 739 586
rect 743 582 747 586
rect 807 582 811 586
rect 815 582 819 586
rect 871 582 875 586
rect 887 582 891 586
rect 935 582 939 586
rect 967 582 971 586
rect 1047 582 1051 586
rect 1127 582 1131 586
rect 1327 582 1331 586
rect 1367 574 1371 578
rect 1511 574 1515 578
rect 1575 574 1579 578
rect 1631 574 1635 578
rect 1655 574 1659 578
rect 1695 574 1699 578
rect 1735 574 1739 578
rect 1775 574 1779 578
rect 1823 574 1827 578
rect 1855 574 1859 578
rect 1911 574 1915 578
rect 1943 574 1947 578
rect 1999 574 2003 578
rect 2031 574 2035 578
rect 2087 574 2091 578
rect 2111 574 2115 578
rect 2175 574 2179 578
rect 2191 574 2195 578
rect 2271 574 2275 578
rect 2343 574 2347 578
rect 2367 574 2371 578
rect 2415 574 2419 578
rect 2463 574 2467 578
rect 2487 574 2491 578
rect 2543 574 2547 578
rect 2583 574 2587 578
rect 111 522 115 526
rect 143 522 147 526
rect 175 522 179 526
rect 207 522 211 526
rect 263 522 267 526
rect 311 522 315 526
rect 351 522 355 526
rect 431 522 435 526
rect 447 522 451 526
rect 543 522 547 526
rect 551 522 555 526
rect 631 522 635 526
rect 671 522 675 526
rect 719 522 723 526
rect 791 522 795 526
rect 799 522 803 526
rect 871 522 875 526
rect 903 522 907 526
rect 951 522 955 526
rect 1007 522 1011 526
rect 1031 522 1035 526
rect 1103 522 1107 526
rect 1111 522 1115 526
rect 1199 522 1203 526
rect 1271 522 1275 526
rect 1327 522 1331 526
rect 1367 514 1371 518
rect 1399 514 1403 518
rect 1455 514 1459 518
rect 1495 514 1499 518
rect 1519 514 1523 518
rect 1559 514 1563 518
rect 1607 514 1611 518
rect 1639 514 1643 518
rect 1695 514 1699 518
rect 1719 514 1723 518
rect 1791 514 1795 518
rect 1807 514 1811 518
rect 1887 514 1891 518
rect 1895 514 1899 518
rect 1983 514 1987 518
rect 2071 514 2075 518
rect 2087 514 2091 518
rect 2159 514 2163 518
rect 2199 514 2203 518
rect 2255 514 2259 518
rect 2311 514 2315 518
rect 2351 514 2355 518
rect 2431 514 2435 518
rect 2447 514 2451 518
rect 2527 514 2531 518
rect 2583 514 2587 518
rect 111 462 115 466
rect 159 462 163 466
rect 223 462 227 466
rect 319 462 323 466
rect 327 462 331 466
rect 423 462 427 466
rect 447 462 451 466
rect 535 462 539 466
rect 567 462 571 466
rect 639 462 643 466
rect 687 462 691 466
rect 743 462 747 466
rect 807 462 811 466
rect 839 462 843 466
rect 919 462 923 466
rect 927 462 931 466
rect 1007 462 1011 466
rect 1023 462 1027 466
rect 1079 462 1083 466
rect 1119 462 1123 466
rect 1151 462 1155 466
rect 1215 462 1219 466
rect 1231 462 1235 466
rect 1287 462 1291 466
rect 1327 462 1331 466
rect 1367 450 1371 454
rect 1415 450 1419 454
rect 1471 450 1475 454
rect 1487 450 1491 454
rect 1535 450 1539 454
rect 1575 450 1579 454
rect 1623 450 1627 454
rect 1663 450 1667 454
rect 1711 450 1715 454
rect 1759 450 1763 454
rect 1807 450 1811 454
rect 1863 450 1867 454
rect 1903 450 1907 454
rect 1975 450 1979 454
rect 1999 450 2003 454
rect 2103 450 2107 454
rect 2111 450 2115 454
rect 2215 450 2219 454
rect 2255 450 2259 454
rect 2327 450 2331 454
rect 2407 450 2411 454
rect 2447 450 2451 454
rect 2543 450 2547 454
rect 2583 450 2587 454
rect 111 398 115 402
rect 143 398 147 402
rect 207 398 211 402
rect 303 398 307 402
rect 399 398 403 402
rect 407 398 411 402
rect 495 398 499 402
rect 519 398 523 402
rect 583 398 587 402
rect 623 398 627 402
rect 671 398 675 402
rect 727 398 731 402
rect 751 398 755 402
rect 823 398 827 402
rect 895 398 899 402
rect 911 398 915 402
rect 967 398 971 402
rect 991 398 995 402
rect 1047 398 1051 402
rect 1063 398 1067 402
rect 1135 398 1139 402
rect 1215 398 1219 402
rect 1271 398 1275 402
rect 1327 398 1331 402
rect 1367 390 1371 394
rect 1399 390 1403 394
rect 1455 390 1459 394
rect 1471 390 1475 394
rect 1511 390 1515 394
rect 1559 390 1563 394
rect 1567 390 1571 394
rect 1631 390 1635 394
rect 1647 390 1651 394
rect 1695 390 1699 394
rect 1743 390 1747 394
rect 1759 390 1763 394
rect 1839 390 1843 394
rect 1847 390 1851 394
rect 1943 390 1947 394
rect 1959 390 1963 394
rect 2071 390 2075 394
rect 2095 390 2099 394
rect 2215 390 2219 394
rect 2239 390 2243 394
rect 2367 390 2371 394
rect 2391 390 2395 394
rect 2527 390 2531 394
rect 2583 390 2587 394
rect 111 338 115 342
rect 159 338 163 342
rect 223 338 227 342
rect 311 338 315 342
rect 319 338 323 342
rect 391 338 395 342
rect 415 338 419 342
rect 471 338 475 342
rect 511 338 515 342
rect 543 338 547 342
rect 599 338 603 342
rect 607 338 611 342
rect 671 338 675 342
rect 687 338 691 342
rect 735 338 739 342
rect 767 338 771 342
rect 799 338 803 342
rect 839 338 843 342
rect 863 338 867 342
rect 911 338 915 342
rect 935 338 939 342
rect 983 338 987 342
rect 1063 338 1067 342
rect 1327 338 1331 342
rect 1367 330 1371 334
rect 1415 330 1419 334
rect 1471 330 1475 334
rect 1527 330 1531 334
rect 1583 330 1587 334
rect 1607 330 1611 334
rect 1647 330 1651 334
rect 1663 330 1667 334
rect 1711 330 1715 334
rect 1719 330 1723 334
rect 1775 330 1779 334
rect 1831 330 1835 334
rect 1855 330 1859 334
rect 1887 330 1891 334
rect 1951 330 1955 334
rect 1959 330 1963 334
rect 2031 330 2035 334
rect 2087 330 2091 334
rect 2119 330 2123 334
rect 2223 330 2227 334
rect 2231 330 2235 334
rect 2335 330 2339 334
rect 2383 330 2387 334
rect 2447 330 2451 334
rect 2543 330 2547 334
rect 2583 330 2587 334
rect 111 274 115 278
rect 143 274 147 278
rect 207 274 211 278
rect 231 274 235 278
rect 295 274 299 278
rect 335 274 339 278
rect 375 274 379 278
rect 431 274 435 278
rect 455 274 459 278
rect 519 274 523 278
rect 527 274 531 278
rect 591 274 595 278
rect 599 274 603 278
rect 655 274 659 278
rect 679 274 683 278
rect 719 274 723 278
rect 751 274 755 278
rect 783 274 787 278
rect 815 274 819 278
rect 847 274 851 278
rect 887 274 891 278
rect 919 274 923 278
rect 959 274 963 278
rect 1031 274 1035 278
rect 1327 274 1331 278
rect 1367 270 1371 274
rect 1591 270 1595 274
rect 1647 270 1651 274
rect 1703 270 1707 274
rect 1727 270 1731 274
rect 1759 270 1763 274
rect 1783 270 1787 274
rect 1815 270 1819 274
rect 1839 270 1843 274
rect 1871 270 1875 274
rect 1895 270 1899 274
rect 1935 270 1939 274
rect 1951 270 1955 274
rect 2007 270 2011 274
rect 2015 270 2019 274
rect 2071 270 2075 274
rect 2103 270 2107 274
rect 2143 270 2147 274
rect 2207 270 2211 274
rect 2231 270 2235 274
rect 2319 270 2323 274
rect 2335 270 2339 274
rect 2431 270 2435 274
rect 2439 270 2443 274
rect 2527 270 2531 274
rect 2583 270 2587 274
rect 111 214 115 218
rect 159 214 163 218
rect 167 214 171 218
rect 247 214 251 218
rect 255 214 259 218
rect 351 214 355 218
rect 447 214 451 218
rect 535 214 539 218
rect 551 214 555 218
rect 615 214 619 218
rect 655 214 659 218
rect 695 214 699 218
rect 751 214 755 218
rect 767 214 771 218
rect 831 214 835 218
rect 847 214 851 218
rect 903 214 907 218
rect 935 214 939 218
rect 975 214 979 218
rect 1023 214 1027 218
rect 1047 214 1051 218
rect 1111 214 1115 218
rect 1199 214 1203 218
rect 1327 214 1331 218
rect 1367 214 1371 218
rect 1463 214 1467 218
rect 1535 214 1539 218
rect 1623 214 1627 218
rect 1719 214 1723 218
rect 1743 214 1747 218
rect 1799 214 1803 218
rect 1823 214 1827 218
rect 1855 214 1859 218
rect 1911 214 1915 218
rect 1927 214 1931 218
rect 1967 214 1971 218
rect 2023 214 2027 218
rect 2031 214 2035 218
rect 2087 214 2091 218
rect 2135 214 2139 218
rect 2159 214 2163 218
rect 2239 214 2243 218
rect 2247 214 2251 218
rect 2343 214 2347 218
rect 2351 214 2355 218
rect 2455 214 2459 218
rect 2543 214 2547 218
rect 2583 214 2587 218
rect 1367 142 1371 146
rect 1399 142 1403 146
rect 1447 142 1451 146
rect 1455 142 1459 146
rect 1511 142 1515 146
rect 1519 142 1523 146
rect 1567 142 1571 146
rect 1607 142 1611 146
rect 1639 142 1643 146
rect 1703 142 1707 146
rect 1719 142 1723 146
rect 1799 142 1803 146
rect 1807 142 1811 146
rect 1879 142 1883 146
rect 1911 142 1915 146
rect 1959 142 1963 146
rect 2015 142 2019 146
rect 2031 142 2035 146
rect 2103 142 2107 146
rect 2119 142 2123 146
rect 2167 142 2171 146
rect 2223 142 2227 146
rect 2231 142 2235 146
rect 2295 142 2299 146
rect 2327 142 2331 146
rect 2359 142 2363 146
rect 2415 142 2419 146
rect 2439 142 2443 146
rect 2471 142 2475 146
rect 2527 142 2531 146
rect 2583 142 2587 146
rect 111 134 115 138
rect 143 134 147 138
rect 151 134 155 138
rect 199 134 203 138
rect 239 134 243 138
rect 255 134 259 138
rect 311 134 315 138
rect 335 134 339 138
rect 367 134 371 138
rect 423 134 427 138
rect 431 134 435 138
rect 479 134 483 138
rect 535 134 539 138
rect 607 134 611 138
rect 639 134 643 138
rect 671 134 675 138
rect 735 134 739 138
rect 799 134 803 138
rect 831 134 835 138
rect 855 134 859 138
rect 911 134 915 138
rect 919 134 923 138
rect 975 134 979 138
rect 1007 134 1011 138
rect 1039 134 1043 138
rect 1095 134 1099 138
rect 1103 134 1107 138
rect 1159 134 1163 138
rect 1183 134 1187 138
rect 1215 134 1219 138
rect 1271 134 1275 138
rect 1327 134 1331 138
rect 1367 86 1371 90
rect 1415 86 1419 90
rect 1471 86 1475 90
rect 1527 86 1531 90
rect 1583 86 1587 90
rect 1655 86 1659 90
rect 1735 86 1739 90
rect 1815 86 1819 90
rect 1895 86 1899 90
rect 1975 86 1979 90
rect 2047 86 2051 90
rect 2119 86 2123 90
rect 2183 86 2187 90
rect 2247 86 2251 90
rect 2311 86 2315 90
rect 2375 86 2379 90
rect 2431 86 2435 90
rect 2487 86 2491 90
rect 2543 86 2547 90
rect 2583 86 2587 90
rect 111 78 115 82
rect 159 78 163 82
rect 215 78 219 82
rect 271 78 275 82
rect 327 78 331 82
rect 383 78 387 82
rect 439 78 443 82
rect 495 78 499 82
rect 551 78 555 82
rect 623 78 627 82
rect 687 78 691 82
rect 751 78 755 82
rect 815 78 819 82
rect 871 78 875 82
rect 927 78 931 82
rect 991 78 995 82
rect 1055 78 1059 82
rect 1119 78 1123 82
rect 1175 78 1179 82
rect 1231 78 1235 82
rect 1287 78 1291 82
rect 1327 78 1331 82
<< m4 >>
rect 84 2657 85 2663
rect 91 2662 1339 2663
rect 91 2658 111 2662
rect 115 2658 159 2662
rect 163 2658 215 2662
rect 219 2658 271 2662
rect 275 2658 327 2662
rect 331 2658 1327 2662
rect 1331 2658 1339 2662
rect 91 2657 1339 2658
rect 1345 2657 1346 2663
rect 1338 2611 1339 2617
rect 1345 2611 1370 2617
rect 1364 2610 2611 2611
rect 96 2601 97 2607
rect 103 2606 1351 2607
rect 103 2602 111 2606
rect 115 2602 143 2606
rect 147 2602 199 2606
rect 203 2602 255 2606
rect 259 2602 263 2606
rect 267 2602 311 2606
rect 315 2602 343 2606
rect 347 2602 431 2606
rect 435 2602 519 2606
rect 523 2602 607 2606
rect 611 2602 687 2606
rect 691 2602 767 2606
rect 771 2602 839 2606
rect 843 2602 903 2606
rect 907 2602 967 2606
rect 971 2602 1031 2606
rect 1035 2602 1095 2606
rect 1099 2602 1159 2606
rect 1163 2602 1215 2606
rect 1219 2602 1271 2606
rect 1275 2602 1327 2606
rect 1331 2602 1351 2606
rect 103 2601 1351 2602
rect 1357 2601 1358 2607
rect 1364 2606 1367 2610
rect 1371 2606 1415 2610
rect 1419 2606 1471 2610
rect 1475 2606 1527 2610
rect 1531 2606 1583 2610
rect 1587 2606 1639 2610
rect 1643 2606 1695 2610
rect 1699 2606 2583 2610
rect 2587 2606 2611 2610
rect 1364 2605 2611 2606
rect 2617 2605 2618 2611
rect 1350 2549 1351 2555
rect 1357 2554 2623 2555
rect 1357 2550 1367 2554
rect 1371 2550 1399 2554
rect 1403 2550 1455 2554
rect 1459 2550 1511 2554
rect 1515 2550 1567 2554
rect 1571 2550 1623 2554
rect 1627 2550 1679 2554
rect 1683 2550 1735 2554
rect 1739 2550 2583 2554
rect 2587 2550 2623 2554
rect 1357 2549 2623 2550
rect 2629 2549 2630 2555
rect 84 2533 85 2539
rect 91 2538 1339 2539
rect 91 2534 111 2538
rect 115 2534 159 2538
rect 163 2534 215 2538
rect 219 2534 279 2538
rect 283 2534 319 2538
rect 323 2534 359 2538
rect 363 2534 431 2538
rect 435 2534 447 2538
rect 451 2534 535 2538
rect 539 2534 551 2538
rect 555 2534 623 2538
rect 627 2534 671 2538
rect 675 2534 703 2538
rect 707 2534 783 2538
rect 787 2534 791 2538
rect 795 2534 855 2538
rect 859 2534 903 2538
rect 907 2534 919 2538
rect 923 2534 983 2538
rect 987 2534 1007 2538
rect 1011 2534 1047 2538
rect 1051 2534 1103 2538
rect 1107 2534 1111 2538
rect 1115 2534 1175 2538
rect 1179 2534 1207 2538
rect 1211 2534 1231 2538
rect 1235 2534 1287 2538
rect 1291 2534 1327 2538
rect 1331 2534 1339 2538
rect 91 2533 1339 2534
rect 1345 2533 1346 2539
rect 1338 2489 1339 2495
rect 1345 2494 2611 2495
rect 1345 2490 1367 2494
rect 1371 2490 1415 2494
rect 1419 2490 1471 2494
rect 1475 2490 1527 2494
rect 1531 2490 1583 2494
rect 1587 2490 1639 2494
rect 1643 2490 1695 2494
rect 1699 2490 1751 2494
rect 1755 2490 2583 2494
rect 2587 2490 2611 2494
rect 1345 2489 2611 2490
rect 2617 2489 2618 2495
rect 96 2469 97 2475
rect 103 2474 1351 2475
rect 103 2470 111 2474
rect 115 2470 143 2474
rect 147 2470 199 2474
rect 203 2470 295 2474
rect 299 2470 303 2474
rect 307 2470 407 2474
rect 411 2470 415 2474
rect 419 2470 519 2474
rect 523 2470 535 2474
rect 539 2470 639 2474
rect 643 2470 655 2474
rect 659 2470 751 2474
rect 755 2470 775 2474
rect 779 2470 855 2474
rect 859 2470 887 2474
rect 891 2470 951 2474
rect 955 2470 991 2474
rect 995 2470 1047 2474
rect 1051 2470 1087 2474
rect 1091 2470 1143 2474
rect 1147 2470 1191 2474
rect 1195 2470 1239 2474
rect 1243 2470 1271 2474
rect 1275 2470 1327 2474
rect 1331 2470 1351 2474
rect 103 2469 1351 2470
rect 1357 2469 1358 2475
rect 1350 2425 1351 2431
rect 1357 2430 2623 2431
rect 1357 2426 1367 2430
rect 1371 2426 1455 2430
rect 1459 2426 1479 2430
rect 1483 2426 1511 2430
rect 1515 2426 1535 2430
rect 1539 2426 1567 2430
rect 1571 2426 1591 2430
rect 1595 2426 1623 2430
rect 1627 2426 1647 2430
rect 1651 2426 1679 2430
rect 1683 2426 1703 2430
rect 1707 2426 1735 2430
rect 1739 2426 1759 2430
rect 1763 2426 2583 2430
rect 2587 2426 2623 2430
rect 1357 2425 2623 2426
rect 2629 2425 2630 2431
rect 84 2405 85 2411
rect 91 2410 1339 2411
rect 91 2406 111 2410
rect 115 2406 159 2410
rect 163 2406 215 2410
rect 219 2406 223 2410
rect 227 2406 287 2410
rect 291 2406 311 2410
rect 315 2406 367 2410
rect 371 2406 423 2410
rect 427 2406 455 2410
rect 459 2406 535 2410
rect 539 2406 543 2410
rect 547 2406 639 2410
rect 643 2406 655 2410
rect 659 2406 727 2410
rect 731 2406 767 2410
rect 771 2406 815 2410
rect 819 2406 871 2410
rect 875 2406 895 2410
rect 899 2406 967 2410
rect 971 2406 975 2410
rect 979 2406 1055 2410
rect 1059 2406 1063 2410
rect 1067 2406 1143 2410
rect 1147 2406 1159 2410
rect 1163 2406 1255 2410
rect 1259 2406 1327 2410
rect 1331 2406 1339 2410
rect 91 2405 1339 2406
rect 1345 2405 1346 2411
rect 1338 2365 1339 2371
rect 1345 2370 2611 2371
rect 1345 2366 1367 2370
rect 1371 2366 1471 2370
rect 1475 2366 1495 2370
rect 1499 2366 1527 2370
rect 1531 2366 1551 2370
rect 1555 2366 1583 2370
rect 1587 2366 1607 2370
rect 1611 2366 1639 2370
rect 1643 2366 1663 2370
rect 1667 2366 1695 2370
rect 1699 2366 1719 2370
rect 1723 2366 1775 2370
rect 1779 2366 2583 2370
rect 2587 2366 2611 2370
rect 1345 2365 2611 2366
rect 2617 2365 2618 2371
rect 96 2341 97 2347
rect 103 2346 1351 2347
rect 103 2342 111 2346
rect 115 2342 207 2346
rect 211 2342 271 2346
rect 275 2342 327 2346
rect 331 2342 351 2346
rect 355 2342 383 2346
rect 387 2342 439 2346
rect 443 2342 503 2346
rect 507 2342 527 2346
rect 531 2342 567 2346
rect 571 2342 623 2346
rect 627 2342 631 2346
rect 635 2342 695 2346
rect 699 2342 711 2346
rect 715 2342 759 2346
rect 763 2342 799 2346
rect 803 2342 823 2346
rect 827 2342 879 2346
rect 883 2342 887 2346
rect 891 2342 951 2346
rect 955 2342 959 2346
rect 963 2342 1015 2346
rect 1019 2342 1039 2346
rect 1043 2342 1127 2346
rect 1131 2342 1327 2346
rect 1331 2342 1351 2346
rect 103 2341 1351 2342
rect 1357 2341 1358 2347
rect 1350 2309 1351 2315
rect 1357 2314 2623 2315
rect 1357 2310 1367 2314
rect 1371 2310 1399 2314
rect 1403 2310 1455 2314
rect 1459 2310 1511 2314
rect 1515 2310 1567 2314
rect 1571 2310 1623 2314
rect 1627 2310 1679 2314
rect 1683 2310 1735 2314
rect 1739 2310 1791 2314
rect 1795 2310 1847 2314
rect 1851 2310 1903 2314
rect 1907 2310 1959 2314
rect 1963 2310 2015 2314
rect 2019 2310 2071 2314
rect 2075 2310 2127 2314
rect 2131 2310 2183 2314
rect 2187 2310 2247 2314
rect 2251 2310 2311 2314
rect 2315 2310 2375 2314
rect 2379 2310 2439 2314
rect 2443 2310 2583 2314
rect 2587 2310 2623 2314
rect 1357 2309 2623 2310
rect 2629 2309 2630 2315
rect 84 2277 85 2283
rect 91 2282 1339 2283
rect 91 2278 111 2282
rect 115 2278 343 2282
rect 347 2278 399 2282
rect 403 2278 407 2282
rect 411 2278 455 2282
rect 459 2278 463 2282
rect 467 2278 519 2282
rect 523 2278 575 2282
rect 579 2278 583 2282
rect 587 2278 631 2282
rect 635 2278 647 2282
rect 651 2278 687 2282
rect 691 2278 711 2282
rect 715 2278 743 2282
rect 747 2278 775 2282
rect 779 2278 799 2282
rect 803 2278 839 2282
rect 843 2278 855 2282
rect 859 2278 903 2282
rect 907 2278 911 2282
rect 915 2278 967 2282
rect 971 2278 1031 2282
rect 1035 2278 1327 2282
rect 1331 2278 1339 2282
rect 91 2277 1339 2278
rect 1345 2277 1346 2283
rect 1338 2253 1339 2259
rect 1345 2258 2611 2259
rect 1345 2254 1367 2258
rect 1371 2254 1415 2258
rect 1419 2254 1471 2258
rect 1475 2254 1511 2258
rect 1515 2254 1527 2258
rect 1531 2254 1583 2258
rect 1587 2254 1623 2258
rect 1627 2254 1639 2258
rect 1643 2254 1695 2258
rect 1699 2254 1727 2258
rect 1731 2254 1751 2258
rect 1755 2254 1807 2258
rect 1811 2254 1823 2258
rect 1827 2254 1863 2258
rect 1867 2254 1903 2258
rect 1907 2254 1919 2258
rect 1923 2254 1975 2258
rect 1979 2254 1983 2258
rect 1987 2254 2031 2258
rect 2035 2254 2055 2258
rect 2059 2254 2087 2258
rect 2091 2254 2119 2258
rect 2123 2254 2143 2258
rect 2147 2254 2191 2258
rect 2195 2254 2199 2258
rect 2203 2254 2263 2258
rect 2267 2254 2327 2258
rect 2331 2254 2335 2258
rect 2339 2254 2391 2258
rect 2395 2254 2455 2258
rect 2459 2254 2583 2258
rect 2587 2254 2611 2258
rect 1345 2253 2611 2254
rect 2617 2253 2618 2259
rect 96 2217 97 2223
rect 103 2222 1351 2223
rect 103 2218 111 2222
rect 115 2218 391 2222
rect 395 2218 423 2222
rect 427 2218 447 2222
rect 451 2218 479 2222
rect 483 2218 503 2222
rect 507 2218 535 2222
rect 539 2218 559 2222
rect 563 2218 591 2222
rect 595 2218 615 2222
rect 619 2218 647 2222
rect 651 2218 671 2222
rect 675 2218 711 2222
rect 715 2218 727 2222
rect 731 2218 783 2222
rect 787 2218 839 2222
rect 843 2218 855 2222
rect 859 2218 895 2222
rect 899 2218 927 2222
rect 931 2218 951 2222
rect 955 2218 999 2222
rect 1003 2218 1071 2222
rect 1075 2218 1143 2222
rect 1147 2218 1215 2222
rect 1219 2218 1271 2222
rect 1275 2218 1327 2222
rect 1331 2218 1351 2222
rect 103 2217 1351 2218
rect 1357 2217 1358 2223
rect 1350 2193 1351 2199
rect 1357 2198 2623 2199
rect 1357 2194 1367 2198
rect 1371 2194 1399 2198
rect 1403 2194 1495 2198
rect 1499 2194 1607 2198
rect 1611 2194 1711 2198
rect 1715 2194 1751 2198
rect 1755 2194 1807 2198
rect 1811 2194 1839 2198
rect 1843 2194 1887 2198
rect 1891 2194 1927 2198
rect 1931 2194 1967 2198
rect 1971 2194 2007 2198
rect 2011 2194 2039 2198
rect 2043 2194 2087 2198
rect 2091 2194 2103 2198
rect 2107 2194 2167 2198
rect 2171 2194 2175 2198
rect 2179 2194 2247 2198
rect 2251 2194 2319 2198
rect 2323 2194 2335 2198
rect 2339 2194 2423 2198
rect 2427 2194 2583 2198
rect 2587 2194 2623 2198
rect 1357 2193 2623 2194
rect 2629 2193 2630 2199
rect 84 2153 85 2159
rect 91 2158 1339 2159
rect 91 2154 111 2158
rect 115 2154 199 2158
rect 203 2154 271 2158
rect 275 2154 351 2158
rect 355 2154 439 2158
rect 443 2154 447 2158
rect 451 2154 495 2158
rect 499 2154 551 2158
rect 555 2154 607 2158
rect 611 2154 663 2158
rect 667 2154 727 2158
rect 731 2154 775 2158
rect 779 2154 799 2158
rect 803 2154 871 2158
rect 875 2154 879 2158
rect 883 2154 943 2158
rect 947 2154 983 2158
rect 987 2154 1015 2158
rect 1019 2154 1079 2158
rect 1083 2154 1087 2158
rect 1091 2154 1159 2158
rect 1163 2154 1183 2158
rect 1187 2154 1231 2158
rect 1235 2154 1287 2158
rect 1291 2154 1327 2158
rect 1331 2154 1339 2158
rect 91 2153 1339 2154
rect 1345 2153 1346 2159
rect 1338 2137 1339 2143
rect 1345 2142 2611 2143
rect 1345 2138 1367 2142
rect 1371 2138 1607 2142
rect 1611 2138 1679 2142
rect 1683 2138 1767 2142
rect 1771 2138 1855 2142
rect 1859 2138 1863 2142
rect 1867 2138 1943 2142
rect 1947 2138 1959 2142
rect 1963 2138 2023 2142
rect 2027 2138 2063 2142
rect 2067 2138 2103 2142
rect 2107 2138 2159 2142
rect 2163 2138 2183 2142
rect 2187 2138 2255 2142
rect 2259 2138 2263 2142
rect 2267 2138 2351 2142
rect 2355 2138 2439 2142
rect 2443 2138 2447 2142
rect 2451 2138 2543 2142
rect 2547 2138 2583 2142
rect 2587 2138 2611 2142
rect 1345 2137 2611 2138
rect 2617 2137 2618 2143
rect 96 2085 97 2091
rect 103 2090 1351 2091
rect 103 2086 111 2090
rect 115 2086 143 2090
rect 147 2086 183 2090
rect 187 2086 199 2090
rect 203 2086 255 2090
rect 259 2086 271 2090
rect 275 2086 335 2090
rect 339 2086 367 2090
rect 371 2086 431 2090
rect 435 2086 463 2090
rect 467 2086 535 2090
rect 539 2086 567 2090
rect 571 2086 647 2090
rect 651 2086 663 2090
rect 667 2086 759 2090
rect 763 2086 847 2090
rect 851 2086 863 2090
rect 867 2086 927 2090
rect 931 2086 967 2090
rect 971 2086 1007 2090
rect 1011 2086 1063 2090
rect 1067 2086 1095 2090
rect 1099 2086 1167 2090
rect 1171 2086 1183 2090
rect 1187 2086 1271 2090
rect 1275 2086 1327 2090
rect 1331 2086 1351 2090
rect 103 2085 1351 2086
rect 1357 2087 1358 2091
rect 1357 2086 2630 2087
rect 1357 2085 1367 2086
rect 1350 2082 1367 2085
rect 1371 2082 1487 2086
rect 1491 2082 1583 2086
rect 1587 2082 1591 2086
rect 1595 2082 1663 2086
rect 1667 2082 1679 2086
rect 1683 2082 1751 2086
rect 1755 2082 1783 2086
rect 1787 2082 1847 2086
rect 1851 2082 1887 2086
rect 1891 2082 1943 2086
rect 1947 2082 1983 2086
rect 1987 2082 2047 2086
rect 2051 2082 2079 2086
rect 2083 2082 2143 2086
rect 2147 2082 2167 2086
rect 2171 2082 2239 2086
rect 2243 2082 2255 2086
rect 2259 2082 2335 2086
rect 2339 2082 2343 2086
rect 2347 2082 2431 2086
rect 2435 2082 2439 2086
rect 2443 2082 2527 2086
rect 2531 2082 2583 2086
rect 2587 2082 2630 2086
rect 1350 2081 2630 2082
rect 1338 2030 2618 2031
rect 1338 2027 1367 2030
rect 84 2021 85 2027
rect 91 2026 1339 2027
rect 91 2022 111 2026
rect 115 2022 159 2026
rect 163 2022 175 2026
rect 179 2022 215 2026
rect 219 2022 239 2026
rect 243 2022 287 2026
rect 291 2022 311 2026
rect 315 2022 383 2026
rect 387 2022 391 2026
rect 395 2022 471 2026
rect 475 2022 479 2026
rect 483 2022 559 2026
rect 563 2022 583 2026
rect 587 2022 647 2026
rect 651 2022 679 2026
rect 683 2022 735 2026
rect 739 2022 775 2026
rect 779 2022 823 2026
rect 827 2022 863 2026
rect 867 2022 911 2026
rect 915 2022 943 2026
rect 947 2022 1007 2026
rect 1011 2022 1023 2026
rect 1027 2022 1103 2026
rect 1107 2022 1111 2026
rect 1115 2022 1199 2026
rect 1203 2022 1327 2026
rect 1331 2022 1339 2026
rect 91 2021 1339 2022
rect 1345 2026 1367 2027
rect 1371 2026 1415 2030
rect 1419 2026 1471 2030
rect 1475 2026 1503 2030
rect 1507 2026 1535 2030
rect 1539 2026 1599 2030
rect 1603 2026 1615 2030
rect 1619 2026 1695 2030
rect 1699 2026 1703 2030
rect 1707 2026 1791 2030
rect 1795 2026 1799 2030
rect 1803 2026 1887 2030
rect 1891 2026 1903 2030
rect 1907 2026 1983 2030
rect 1987 2026 1999 2030
rect 2003 2026 2079 2030
rect 2083 2026 2095 2030
rect 2099 2026 2175 2030
rect 2179 2026 2183 2030
rect 2187 2026 2271 2030
rect 2275 2026 2359 2030
rect 2363 2026 2367 2030
rect 2371 2026 2455 2030
rect 2459 2026 2463 2030
rect 2467 2026 2543 2030
rect 2547 2026 2583 2030
rect 2587 2026 2618 2030
rect 1345 2025 2618 2026
rect 1345 2021 1346 2025
rect 96 1965 97 1971
rect 103 1970 1351 1971
rect 103 1966 111 1970
rect 115 1966 159 1970
rect 163 1966 223 1970
rect 227 1966 295 1970
rect 299 1966 375 1970
rect 379 1966 383 1970
rect 387 1966 439 1970
rect 443 1966 455 1970
rect 459 1966 495 1970
rect 499 1966 543 1970
rect 547 1966 551 1970
rect 555 1966 607 1970
rect 611 1966 631 1970
rect 635 1966 671 1970
rect 675 1966 719 1970
rect 723 1966 735 1970
rect 739 1966 807 1970
rect 811 1966 879 1970
rect 883 1966 895 1970
rect 899 1966 951 1970
rect 955 1966 991 1970
rect 995 1966 1023 1970
rect 1027 1966 1087 1970
rect 1091 1966 1327 1970
rect 1331 1966 1351 1970
rect 103 1965 1351 1966
rect 1357 1970 2630 1971
rect 1357 1966 1367 1970
rect 1371 1966 1399 1970
rect 1403 1966 1455 1970
rect 1459 1966 1519 1970
rect 1523 1966 1599 1970
rect 1603 1966 1679 1970
rect 1683 1966 1687 1970
rect 1691 1966 1759 1970
rect 1763 1966 1775 1970
rect 1779 1966 1855 1970
rect 1859 1966 1871 1970
rect 1875 1966 1967 1970
rect 1971 1966 2063 1970
rect 2067 1966 2095 1970
rect 2099 1966 2159 1970
rect 2163 1966 2239 1970
rect 2243 1966 2255 1970
rect 2259 1966 2351 1970
rect 2355 1966 2391 1970
rect 2395 1966 2447 1970
rect 2451 1966 2527 1970
rect 2531 1966 2583 1970
rect 2587 1966 2630 1970
rect 1357 1965 2630 1966
rect 84 1909 85 1915
rect 91 1914 1339 1915
rect 91 1910 111 1914
rect 115 1910 399 1914
rect 403 1910 455 1914
rect 459 1910 511 1914
rect 515 1910 519 1914
rect 523 1910 567 1914
rect 571 1910 575 1914
rect 579 1910 623 1914
rect 627 1910 631 1914
rect 635 1910 687 1914
rect 691 1910 743 1914
rect 747 1910 751 1914
rect 755 1910 807 1914
rect 811 1910 823 1914
rect 827 1910 871 1914
rect 875 1910 895 1914
rect 899 1910 935 1914
rect 939 1910 967 1914
rect 971 1910 999 1914
rect 1003 1910 1039 1914
rect 1043 1910 1327 1914
rect 1331 1910 1339 1914
rect 91 1909 1339 1910
rect 1345 1914 2618 1915
rect 1345 1910 1367 1914
rect 1371 1910 1415 1914
rect 1419 1910 1471 1914
rect 1475 1910 1535 1914
rect 1539 1910 1575 1914
rect 1579 1910 1615 1914
rect 1619 1910 1631 1914
rect 1635 1910 1687 1914
rect 1691 1910 1695 1914
rect 1699 1910 1743 1914
rect 1747 1910 1775 1914
rect 1779 1910 1799 1914
rect 1803 1910 1855 1914
rect 1859 1910 1871 1914
rect 1875 1910 1927 1914
rect 1931 1910 1983 1914
rect 1987 1910 2015 1914
rect 2019 1910 2111 1914
rect 2115 1910 2127 1914
rect 2131 1910 2247 1914
rect 2251 1910 2255 1914
rect 2259 1910 2383 1914
rect 2387 1910 2407 1914
rect 2411 1910 2519 1914
rect 2523 1910 2543 1914
rect 2547 1910 2583 1914
rect 2587 1910 2618 1914
rect 1345 1909 2618 1910
rect 96 1849 97 1855
rect 103 1854 1351 1855
rect 103 1850 111 1854
rect 115 1850 143 1854
rect 147 1850 199 1854
rect 203 1850 255 1854
rect 259 1850 311 1854
rect 315 1850 375 1854
rect 379 1850 455 1854
rect 459 1850 503 1854
rect 507 1850 543 1854
rect 547 1850 559 1854
rect 563 1850 615 1854
rect 619 1850 631 1854
rect 635 1850 671 1854
rect 675 1850 719 1854
rect 723 1850 727 1854
rect 731 1850 791 1854
rect 795 1850 799 1854
rect 803 1850 855 1854
rect 859 1850 887 1854
rect 891 1850 919 1854
rect 923 1850 975 1854
rect 979 1850 983 1854
rect 987 1850 1063 1854
rect 1067 1850 1327 1854
rect 1331 1850 1351 1854
rect 103 1849 1351 1850
rect 1357 1851 1358 1855
rect 1357 1850 2630 1851
rect 1357 1849 1367 1850
rect 1350 1846 1367 1849
rect 1371 1846 1559 1850
rect 1563 1846 1615 1850
rect 1619 1846 1623 1850
rect 1627 1846 1671 1850
rect 1675 1846 1679 1850
rect 1683 1846 1727 1850
rect 1731 1846 1735 1850
rect 1739 1846 1783 1850
rect 1787 1846 1791 1850
rect 1795 1846 1839 1850
rect 1843 1846 1847 1850
rect 1851 1846 1903 1850
rect 1907 1846 1911 1850
rect 1915 1846 1967 1850
rect 1971 1846 1999 1850
rect 2003 1846 2039 1850
rect 2043 1846 2111 1850
rect 2115 1846 2127 1850
rect 2131 1846 2223 1850
rect 2227 1846 2231 1850
rect 2235 1846 2327 1850
rect 2331 1846 2367 1850
rect 2371 1846 2439 1850
rect 2443 1846 2503 1850
rect 2507 1846 2527 1850
rect 2531 1846 2583 1850
rect 2587 1846 2630 1850
rect 1350 1845 2630 1846
rect 84 1785 85 1791
rect 91 1790 1339 1791
rect 91 1786 111 1790
rect 115 1786 159 1790
rect 163 1786 215 1790
rect 219 1786 255 1790
rect 259 1786 271 1790
rect 275 1786 327 1790
rect 331 1786 375 1790
rect 379 1786 391 1790
rect 395 1786 471 1790
rect 475 1786 503 1790
rect 507 1786 559 1790
rect 563 1786 623 1790
rect 627 1786 647 1790
rect 651 1786 735 1790
rect 739 1786 743 1790
rect 747 1786 815 1790
rect 819 1786 855 1790
rect 859 1786 903 1790
rect 907 1786 959 1790
rect 963 1786 991 1790
rect 995 1786 1055 1790
rect 1059 1786 1079 1790
rect 1083 1786 1151 1790
rect 1155 1786 1247 1790
rect 1251 1786 1327 1790
rect 1331 1786 1339 1790
rect 91 1785 1339 1786
rect 1345 1787 1346 1791
rect 1345 1786 2618 1787
rect 1345 1785 1367 1786
rect 1338 1782 1367 1785
rect 1371 1782 1471 1786
rect 1475 1782 1535 1786
rect 1539 1782 1615 1786
rect 1619 1782 1639 1786
rect 1643 1782 1695 1786
rect 1699 1782 1751 1786
rect 1755 1782 1783 1786
rect 1787 1782 1807 1786
rect 1811 1782 1863 1786
rect 1867 1782 1879 1786
rect 1883 1782 1919 1786
rect 1923 1782 1975 1786
rect 1979 1782 1983 1786
rect 1987 1782 2055 1786
rect 2059 1782 2071 1786
rect 2075 1782 2143 1786
rect 2147 1782 2167 1786
rect 2171 1782 2239 1786
rect 2243 1782 2263 1786
rect 2267 1782 2343 1786
rect 2347 1782 2359 1786
rect 2363 1782 2455 1786
rect 2459 1782 2463 1786
rect 2467 1782 2543 1786
rect 2547 1782 2583 1786
rect 2587 1782 2618 1786
rect 1338 1781 2618 1782
rect 96 1729 97 1735
rect 103 1734 1351 1735
rect 103 1730 111 1734
rect 115 1730 143 1734
rect 147 1730 239 1734
rect 243 1730 263 1734
rect 267 1730 359 1734
rect 363 1730 415 1734
rect 419 1730 487 1734
rect 491 1730 567 1734
rect 571 1730 607 1734
rect 611 1730 711 1734
rect 715 1730 727 1734
rect 731 1730 839 1734
rect 843 1730 855 1734
rect 859 1730 943 1734
rect 947 1730 999 1734
rect 1003 1730 1039 1734
rect 1043 1730 1135 1734
rect 1139 1730 1143 1734
rect 1147 1730 1231 1734
rect 1235 1730 1271 1734
rect 1275 1730 1327 1734
rect 1331 1730 1351 1734
rect 103 1729 1351 1730
rect 1357 1729 1358 1735
rect 1350 1727 1358 1729
rect 1350 1721 1351 1727
rect 1357 1726 2623 1727
rect 1357 1722 1367 1726
rect 1371 1722 1399 1726
rect 1403 1722 1455 1726
rect 1459 1722 1479 1726
rect 1483 1722 1519 1726
rect 1523 1722 1599 1726
rect 1603 1722 1679 1726
rect 1683 1722 1719 1726
rect 1723 1722 1767 1726
rect 1771 1722 1839 1726
rect 1843 1722 1863 1726
rect 1867 1722 1951 1726
rect 1955 1722 1959 1726
rect 1963 1722 2055 1726
rect 2059 1722 2151 1726
rect 2155 1722 2159 1726
rect 2163 1722 2247 1726
rect 2251 1722 2255 1726
rect 2259 1722 2343 1726
rect 2347 1722 2351 1726
rect 2355 1722 2447 1726
rect 2451 1722 2527 1726
rect 2531 1722 2583 1726
rect 2587 1722 2623 1726
rect 1357 1721 2623 1722
rect 2629 1721 2630 1727
rect 84 1669 85 1675
rect 91 1674 1339 1675
rect 91 1670 111 1674
rect 115 1670 159 1674
rect 163 1670 223 1674
rect 227 1670 279 1674
rect 283 1670 303 1674
rect 307 1670 383 1674
rect 387 1670 431 1674
rect 435 1670 463 1674
rect 467 1670 535 1674
rect 539 1670 583 1674
rect 587 1670 607 1674
rect 611 1670 679 1674
rect 683 1670 727 1674
rect 731 1670 767 1674
rect 771 1670 863 1674
rect 867 1670 871 1674
rect 875 1670 967 1674
rect 971 1670 1015 1674
rect 1019 1670 1079 1674
rect 1083 1670 1159 1674
rect 1163 1670 1191 1674
rect 1195 1670 1287 1674
rect 1291 1670 1327 1674
rect 1331 1670 1339 1674
rect 91 1669 1339 1670
rect 1345 1671 1346 1675
rect 1345 1670 2618 1671
rect 1345 1669 1367 1670
rect 1338 1666 1367 1669
rect 1371 1666 1415 1670
rect 1419 1666 1495 1670
rect 1499 1666 1503 1670
rect 1507 1666 1615 1670
rect 1619 1666 1623 1670
rect 1627 1666 1735 1670
rect 1739 1666 1751 1670
rect 1755 1666 1855 1670
rect 1859 1666 1879 1670
rect 1883 1666 1967 1670
rect 1971 1666 1999 1670
rect 2003 1666 2071 1670
rect 2075 1666 2119 1670
rect 2123 1666 2175 1670
rect 2179 1666 2231 1670
rect 2235 1666 2271 1670
rect 2275 1666 2343 1670
rect 2347 1666 2367 1670
rect 2371 1666 2455 1670
rect 2459 1666 2463 1670
rect 2467 1666 2543 1670
rect 2547 1666 2583 1670
rect 2587 1666 2618 1670
rect 1338 1665 2618 1666
rect 96 1613 97 1619
rect 103 1618 1351 1619
rect 103 1614 111 1618
rect 115 1614 143 1618
rect 147 1614 207 1618
rect 211 1614 247 1618
rect 251 1614 287 1618
rect 291 1614 367 1618
rect 371 1614 447 1618
rect 451 1614 479 1618
rect 483 1614 519 1618
rect 523 1614 575 1618
rect 579 1614 591 1618
rect 595 1614 663 1618
rect 667 1614 671 1618
rect 675 1614 751 1618
rect 755 1614 767 1618
rect 771 1614 847 1618
rect 851 1614 863 1618
rect 867 1614 951 1618
rect 955 1614 959 1618
rect 963 1614 1063 1618
rect 1067 1614 1175 1618
rect 1179 1614 1271 1618
rect 1275 1614 1327 1618
rect 1331 1614 1351 1618
rect 103 1613 1351 1614
rect 1357 1613 1358 1619
rect 1350 1597 1351 1603
rect 1357 1602 2623 1603
rect 1357 1598 1367 1602
rect 1371 1598 1399 1602
rect 1403 1598 1487 1602
rect 1491 1598 1495 1602
rect 1499 1598 1607 1602
rect 1611 1598 1615 1602
rect 1619 1598 1735 1602
rect 1739 1598 1743 1602
rect 1747 1598 1863 1602
rect 1867 1598 1983 1602
rect 1987 1598 2095 1602
rect 2099 1598 2103 1602
rect 2107 1598 2199 1602
rect 2203 1598 2215 1602
rect 2219 1598 2295 1602
rect 2299 1598 2327 1602
rect 2331 1598 2391 1602
rect 2395 1598 2439 1602
rect 2443 1598 2495 1602
rect 2499 1598 2527 1602
rect 2531 1598 2583 1602
rect 2587 1598 2623 1602
rect 1357 1597 2623 1598
rect 2629 1597 2630 1603
rect 84 1553 85 1559
rect 91 1558 1339 1559
rect 91 1554 111 1558
rect 115 1554 159 1558
rect 163 1554 231 1558
rect 235 1554 263 1558
rect 267 1554 335 1558
rect 339 1554 383 1558
rect 387 1554 455 1558
rect 459 1554 495 1558
rect 499 1554 583 1558
rect 587 1554 591 1558
rect 595 1554 687 1558
rect 691 1554 719 1558
rect 723 1554 783 1558
rect 787 1554 863 1558
rect 867 1554 879 1558
rect 883 1554 975 1558
rect 979 1554 1007 1558
rect 1011 1554 1079 1558
rect 1083 1554 1151 1558
rect 1155 1554 1191 1558
rect 1195 1554 1287 1558
rect 1291 1554 1327 1558
rect 1331 1554 1339 1558
rect 91 1553 1339 1554
rect 1345 1553 1346 1559
rect 1338 1537 1339 1543
rect 1345 1542 2611 1543
rect 1345 1538 1367 1542
rect 1371 1538 1415 1542
rect 1419 1538 1511 1542
rect 1515 1538 1527 1542
rect 1531 1538 1631 1542
rect 1635 1538 1647 1542
rect 1651 1538 1759 1542
rect 1763 1538 1767 1542
rect 1771 1538 1879 1542
rect 1883 1538 1983 1542
rect 1987 1538 1999 1542
rect 2003 1538 2079 1542
rect 2083 1538 2111 1542
rect 2115 1538 2167 1542
rect 2171 1538 2215 1542
rect 2219 1538 2255 1542
rect 2259 1538 2311 1542
rect 2315 1538 2335 1542
rect 2339 1538 2407 1542
rect 2411 1538 2487 1542
rect 2491 1538 2511 1542
rect 2515 1538 2543 1542
rect 2547 1538 2583 1542
rect 2587 1538 2611 1542
rect 1345 1537 2611 1538
rect 2617 1537 2618 1543
rect 96 1497 97 1503
rect 103 1502 1351 1503
rect 103 1498 111 1502
rect 115 1498 143 1502
rect 147 1498 199 1502
rect 203 1498 215 1502
rect 219 1498 271 1502
rect 275 1498 319 1502
rect 323 1498 367 1502
rect 371 1498 439 1502
rect 443 1498 479 1502
rect 483 1498 567 1502
rect 571 1498 591 1502
rect 595 1498 703 1502
rect 707 1498 807 1502
rect 811 1498 847 1502
rect 851 1498 911 1502
rect 915 1498 991 1502
rect 995 1498 1007 1502
rect 1011 1498 1103 1502
rect 1107 1498 1135 1502
rect 1139 1498 1199 1502
rect 1203 1498 1271 1502
rect 1275 1498 1327 1502
rect 1331 1498 1351 1502
rect 103 1497 1351 1498
rect 1357 1497 1358 1503
rect 1350 1473 1351 1479
rect 1357 1478 2623 1479
rect 1357 1474 1367 1478
rect 1371 1474 1399 1478
rect 1403 1474 1503 1478
rect 1507 1474 1511 1478
rect 1515 1474 1631 1478
rect 1635 1474 1751 1478
rect 1755 1474 1863 1478
rect 1867 1474 1871 1478
rect 1875 1474 1967 1478
rect 1971 1474 1983 1478
rect 1987 1474 2063 1478
rect 2067 1474 2087 1478
rect 2091 1474 2151 1478
rect 2155 1474 2183 1478
rect 2187 1474 2239 1478
rect 2243 1474 2271 1478
rect 2275 1474 2319 1478
rect 2323 1474 2359 1478
rect 2363 1474 2391 1478
rect 2395 1474 2455 1478
rect 2459 1474 2471 1478
rect 2475 1474 2527 1478
rect 2531 1474 2583 1478
rect 2587 1474 2623 1478
rect 1357 1473 2623 1474
rect 2629 1473 2630 1479
rect 84 1437 85 1443
rect 91 1442 1339 1443
rect 91 1438 111 1442
rect 115 1438 159 1442
rect 163 1438 215 1442
rect 219 1438 255 1442
rect 259 1438 287 1442
rect 291 1438 311 1442
rect 315 1438 375 1442
rect 379 1438 383 1442
rect 387 1438 447 1442
rect 451 1438 495 1442
rect 499 1438 527 1442
rect 531 1438 607 1442
rect 611 1438 695 1442
rect 699 1438 719 1442
rect 723 1438 783 1442
rect 787 1438 823 1442
rect 827 1438 871 1442
rect 875 1438 927 1442
rect 931 1438 959 1442
rect 963 1438 1023 1442
rect 1027 1438 1055 1442
rect 1059 1438 1119 1442
rect 1123 1438 1151 1442
rect 1155 1438 1215 1442
rect 1219 1438 1287 1442
rect 1291 1438 1327 1442
rect 1331 1438 1339 1442
rect 91 1437 1339 1438
rect 1345 1437 1346 1443
rect 1338 1413 1339 1419
rect 1345 1418 2611 1419
rect 1345 1414 1367 1418
rect 1371 1414 1415 1418
rect 1419 1414 1471 1418
rect 1475 1414 1519 1418
rect 1523 1414 1551 1418
rect 1555 1414 1631 1418
rect 1635 1414 1647 1418
rect 1651 1414 1711 1418
rect 1715 1414 1767 1418
rect 1771 1414 1791 1418
rect 1795 1414 1871 1418
rect 1875 1414 1887 1418
rect 1891 1414 1959 1418
rect 1963 1414 1999 1418
rect 2003 1414 2055 1418
rect 2059 1414 2103 1418
rect 2107 1414 2167 1418
rect 2171 1414 2199 1418
rect 2203 1414 2287 1418
rect 2291 1414 2295 1418
rect 2299 1414 2375 1418
rect 2379 1414 2431 1418
rect 2435 1414 2471 1418
rect 2475 1414 2543 1418
rect 2547 1414 2583 1418
rect 2587 1414 2611 1418
rect 1345 1413 2611 1414
rect 2617 1413 2618 1419
rect 96 1373 97 1379
rect 103 1378 1351 1379
rect 103 1374 111 1378
rect 115 1374 239 1378
rect 243 1374 295 1378
rect 299 1374 359 1378
rect 363 1374 415 1378
rect 419 1374 431 1378
rect 435 1374 471 1378
rect 475 1374 511 1378
rect 515 1374 527 1378
rect 531 1374 591 1378
rect 595 1374 671 1378
rect 675 1374 679 1378
rect 683 1374 751 1378
rect 755 1374 767 1378
rect 771 1374 839 1378
rect 843 1374 855 1378
rect 859 1374 935 1378
rect 939 1374 943 1378
rect 947 1374 1031 1378
rect 1035 1374 1039 1378
rect 1043 1374 1127 1378
rect 1131 1374 1135 1378
rect 1139 1374 1231 1378
rect 1235 1374 1327 1378
rect 1331 1374 1351 1378
rect 103 1373 1351 1374
rect 1357 1373 1358 1379
rect 1350 1357 1351 1363
rect 1357 1362 2623 1363
rect 1357 1358 1367 1362
rect 1371 1358 1399 1362
rect 1403 1358 1423 1362
rect 1427 1358 1455 1362
rect 1459 1358 1495 1362
rect 1499 1358 1535 1362
rect 1539 1358 1575 1362
rect 1579 1358 1615 1362
rect 1619 1358 1655 1362
rect 1659 1358 1695 1362
rect 1699 1358 1759 1362
rect 1763 1358 1775 1362
rect 1779 1358 1855 1362
rect 1859 1358 1879 1362
rect 1883 1358 1943 1362
rect 1947 1358 2023 1362
rect 2027 1358 2039 1362
rect 2043 1358 2151 1362
rect 2155 1358 2183 1362
rect 2187 1358 2279 1362
rect 2283 1358 2359 1362
rect 2363 1358 2415 1362
rect 2419 1358 2527 1362
rect 2531 1358 2583 1362
rect 2587 1358 2623 1362
rect 1357 1357 2623 1358
rect 2629 1357 2630 1363
rect 84 1309 85 1315
rect 91 1314 1339 1315
rect 91 1310 111 1314
rect 115 1310 375 1314
rect 379 1310 431 1314
rect 435 1310 471 1314
rect 475 1310 487 1314
rect 491 1310 527 1314
rect 531 1310 543 1314
rect 547 1310 583 1314
rect 587 1310 607 1314
rect 611 1310 647 1314
rect 651 1310 687 1314
rect 691 1310 727 1314
rect 731 1310 767 1314
rect 771 1310 807 1314
rect 811 1310 855 1314
rect 859 1310 895 1314
rect 899 1310 951 1314
rect 955 1310 991 1314
rect 995 1310 1047 1314
rect 1051 1310 1095 1314
rect 1099 1310 1143 1314
rect 1147 1310 1199 1314
rect 1203 1310 1247 1314
rect 1251 1310 1287 1314
rect 1291 1310 1327 1314
rect 1331 1310 1339 1314
rect 91 1309 1339 1310
rect 1345 1309 1346 1315
rect 1338 1307 1346 1309
rect 1338 1301 1339 1307
rect 1345 1306 2611 1307
rect 1345 1302 1367 1306
rect 1371 1302 1431 1306
rect 1435 1302 1439 1306
rect 1443 1302 1495 1306
rect 1499 1302 1511 1306
rect 1515 1302 1559 1306
rect 1563 1302 1591 1306
rect 1595 1302 1631 1306
rect 1635 1302 1671 1306
rect 1675 1302 1703 1306
rect 1707 1302 1775 1306
rect 1779 1302 1855 1306
rect 1859 1302 1895 1306
rect 1899 1302 1943 1306
rect 1947 1302 2039 1306
rect 2043 1302 2047 1306
rect 2051 1302 2159 1306
rect 2163 1302 2199 1306
rect 2203 1302 2287 1306
rect 2291 1302 2375 1306
rect 2379 1302 2423 1306
rect 2427 1302 2543 1306
rect 2547 1302 2583 1306
rect 2587 1302 2611 1306
rect 1345 1301 2611 1302
rect 2617 1301 2618 1307
rect 96 1249 97 1255
rect 103 1254 1351 1255
rect 103 1250 111 1254
rect 115 1250 383 1254
rect 387 1250 439 1254
rect 443 1250 455 1254
rect 459 1250 503 1254
rect 507 1250 511 1254
rect 515 1250 567 1254
rect 571 1250 575 1254
rect 579 1250 631 1254
rect 635 1250 647 1254
rect 651 1250 711 1254
rect 715 1250 727 1254
rect 731 1250 791 1254
rect 795 1250 815 1254
rect 819 1250 879 1254
rect 883 1250 903 1254
rect 907 1250 975 1254
rect 979 1250 991 1254
rect 995 1250 1079 1254
rect 1083 1250 1175 1254
rect 1179 1250 1183 1254
rect 1187 1250 1271 1254
rect 1275 1250 1327 1254
rect 1331 1250 1351 1254
rect 103 1249 1351 1250
rect 1357 1249 1358 1255
rect 1350 1247 1358 1249
rect 1350 1241 1351 1247
rect 1357 1246 2623 1247
rect 1357 1242 1367 1246
rect 1371 1242 1399 1246
rect 1403 1242 1415 1246
rect 1419 1242 1455 1246
rect 1459 1242 1479 1246
rect 1483 1242 1535 1246
rect 1539 1242 1543 1246
rect 1547 1242 1615 1246
rect 1619 1242 1687 1246
rect 1691 1242 1695 1246
rect 1699 1242 1759 1246
rect 1763 1242 1775 1246
rect 1779 1242 1839 1246
rect 1843 1242 1855 1246
rect 1859 1242 1927 1246
rect 1931 1242 1943 1246
rect 1947 1242 2031 1246
rect 2035 1242 2039 1246
rect 2043 1242 2143 1246
rect 2147 1242 2151 1246
rect 2155 1242 2271 1246
rect 2275 1242 2279 1246
rect 2283 1242 2407 1246
rect 2411 1242 2415 1246
rect 2419 1242 2527 1246
rect 2531 1242 2583 1246
rect 2587 1242 2623 1246
rect 1357 1241 2623 1242
rect 2629 1241 2630 1247
rect 84 1189 85 1195
rect 91 1194 1339 1195
rect 91 1190 111 1194
rect 115 1190 279 1194
rect 283 1190 343 1194
rect 347 1190 399 1194
rect 403 1190 415 1194
rect 419 1190 455 1194
rect 459 1190 495 1194
rect 499 1190 519 1194
rect 523 1190 583 1194
rect 587 1190 591 1194
rect 595 1190 663 1194
rect 667 1190 671 1194
rect 675 1190 743 1194
rect 747 1190 759 1194
rect 763 1190 831 1194
rect 835 1190 847 1194
rect 851 1190 919 1194
rect 923 1190 935 1194
rect 939 1190 1007 1194
rect 1011 1190 1015 1194
rect 1019 1190 1087 1194
rect 1091 1190 1095 1194
rect 1099 1190 1159 1194
rect 1163 1190 1191 1194
rect 1195 1190 1231 1194
rect 1235 1190 1287 1194
rect 1291 1190 1327 1194
rect 1331 1190 1339 1194
rect 91 1189 1339 1190
rect 1345 1189 1346 1195
rect 1338 1177 1339 1183
rect 1345 1182 2611 1183
rect 1345 1178 1367 1182
rect 1371 1178 1415 1182
rect 1419 1178 1471 1182
rect 1475 1178 1551 1182
rect 1555 1178 1631 1182
rect 1635 1178 1695 1182
rect 1699 1178 1711 1182
rect 1715 1178 1767 1182
rect 1771 1178 1791 1182
rect 1795 1178 1847 1182
rect 1851 1178 1871 1182
rect 1875 1178 1919 1182
rect 1923 1178 1959 1182
rect 1963 1178 1991 1182
rect 1995 1178 2055 1182
rect 2059 1178 2063 1182
rect 2067 1178 2135 1182
rect 2139 1178 2167 1182
rect 2171 1178 2207 1182
rect 2211 1178 2287 1182
rect 2291 1178 2295 1182
rect 2299 1178 2367 1182
rect 2371 1178 2431 1182
rect 2435 1178 2543 1182
rect 2547 1178 2583 1182
rect 2587 1178 2611 1182
rect 1345 1177 2611 1178
rect 2617 1177 2618 1183
rect 96 1125 97 1131
rect 103 1130 1351 1131
rect 103 1126 111 1130
rect 115 1126 143 1130
rect 147 1126 207 1130
rect 211 1126 263 1130
rect 267 1126 271 1130
rect 275 1126 327 1130
rect 331 1126 343 1130
rect 347 1126 399 1130
rect 403 1126 423 1130
rect 427 1126 479 1130
rect 483 1126 503 1130
rect 507 1126 567 1130
rect 571 1126 583 1130
rect 587 1126 655 1130
rect 659 1126 663 1130
rect 667 1126 743 1130
rect 747 1126 831 1130
rect 835 1126 919 1130
rect 923 1126 999 1130
rect 1003 1126 1007 1130
rect 1011 1126 1071 1130
rect 1075 1126 1143 1130
rect 1147 1126 1215 1130
rect 1219 1126 1271 1130
rect 1275 1126 1327 1130
rect 1331 1126 1351 1130
rect 103 1125 1351 1126
rect 1357 1127 1358 1131
rect 1357 1126 2630 1127
rect 1357 1125 1367 1126
rect 1350 1122 1367 1125
rect 1371 1122 1399 1126
rect 1403 1122 1479 1126
rect 1483 1122 1583 1126
rect 1587 1122 1679 1126
rect 1683 1122 1687 1126
rect 1691 1122 1751 1126
rect 1755 1122 1783 1126
rect 1787 1122 1831 1126
rect 1835 1122 1879 1126
rect 1883 1122 1903 1126
rect 1907 1122 1975 1126
rect 1979 1122 2047 1126
rect 2051 1122 2063 1126
rect 2067 1122 2119 1126
rect 2123 1122 2151 1126
rect 2155 1122 2191 1126
rect 2195 1122 2239 1126
rect 2243 1122 2271 1126
rect 2275 1122 2327 1126
rect 2331 1122 2351 1126
rect 2355 1122 2415 1126
rect 2419 1122 2583 1126
rect 2587 1122 2630 1126
rect 1350 1121 2630 1122
rect 84 1065 85 1071
rect 91 1070 1339 1071
rect 91 1066 111 1070
rect 115 1066 159 1070
rect 163 1066 215 1070
rect 219 1066 223 1070
rect 227 1066 287 1070
rect 291 1066 359 1070
rect 363 1066 383 1070
rect 387 1066 439 1070
rect 443 1066 479 1070
rect 483 1066 519 1070
rect 523 1066 583 1070
rect 587 1066 599 1070
rect 603 1066 679 1070
rect 683 1066 687 1070
rect 691 1066 759 1070
rect 763 1066 783 1070
rect 787 1066 847 1070
rect 851 1066 879 1070
rect 883 1066 935 1070
rect 939 1066 967 1070
rect 971 1066 1023 1070
rect 1027 1066 1063 1070
rect 1067 1066 1159 1070
rect 1163 1066 1327 1070
rect 1331 1066 1339 1070
rect 91 1065 1339 1066
rect 1345 1070 2618 1071
rect 1345 1066 1367 1070
rect 1371 1066 1415 1070
rect 1419 1066 1495 1070
rect 1499 1066 1511 1070
rect 1515 1066 1599 1070
rect 1603 1066 1631 1070
rect 1635 1066 1703 1070
rect 1707 1066 1751 1070
rect 1755 1066 1799 1070
rect 1803 1066 1871 1070
rect 1875 1066 1895 1070
rect 1899 1066 1991 1070
rect 1995 1066 2079 1070
rect 2083 1066 2103 1070
rect 2107 1066 2167 1070
rect 2171 1066 2199 1070
rect 2203 1066 2255 1070
rect 2259 1066 2295 1070
rect 2299 1066 2343 1070
rect 2347 1066 2383 1070
rect 2387 1066 2431 1070
rect 2435 1066 2471 1070
rect 2475 1066 2543 1070
rect 2547 1066 2583 1070
rect 2587 1066 2618 1070
rect 1345 1065 2618 1066
rect 96 1005 97 1011
rect 103 1010 1351 1011
rect 103 1006 111 1010
rect 115 1006 143 1010
rect 147 1006 199 1010
rect 203 1006 271 1010
rect 275 1006 279 1010
rect 283 1006 367 1010
rect 371 1006 383 1010
rect 387 1006 463 1010
rect 467 1006 495 1010
rect 499 1006 567 1010
rect 571 1006 615 1010
rect 619 1006 671 1010
rect 675 1006 727 1010
rect 731 1006 767 1010
rect 771 1006 839 1010
rect 843 1006 863 1010
rect 867 1006 951 1010
rect 955 1006 1047 1010
rect 1051 1006 1055 1010
rect 1059 1006 1143 1010
rect 1147 1006 1159 1010
rect 1163 1006 1271 1010
rect 1275 1006 1327 1010
rect 1331 1006 1351 1010
rect 103 1005 1351 1006
rect 1357 1010 2630 1011
rect 1357 1006 1367 1010
rect 1371 1006 1399 1010
rect 1403 1006 1487 1010
rect 1491 1006 1495 1010
rect 1499 1006 1583 1010
rect 1587 1006 1615 1010
rect 1619 1006 1695 1010
rect 1699 1006 1735 1010
rect 1739 1006 1807 1010
rect 1811 1006 1855 1010
rect 1859 1006 1919 1010
rect 1923 1006 1975 1010
rect 1979 1006 2023 1010
rect 2027 1006 2087 1010
rect 2091 1006 2119 1010
rect 2123 1006 2183 1010
rect 2187 1006 2215 1010
rect 2219 1006 2279 1010
rect 2283 1006 2303 1010
rect 2307 1006 2367 1010
rect 2371 1006 2383 1010
rect 2387 1006 2455 1010
rect 2459 1006 2463 1010
rect 2467 1006 2527 1010
rect 2531 1006 2583 1010
rect 2587 1006 2630 1010
rect 1357 1005 2630 1006
rect 84 941 85 947
rect 91 946 1339 947
rect 91 942 111 946
rect 115 942 159 946
rect 163 942 215 946
rect 219 942 287 946
rect 291 942 295 946
rect 299 942 375 946
rect 379 942 399 946
rect 403 942 471 946
rect 475 942 511 946
rect 515 942 567 946
rect 571 942 631 946
rect 635 942 671 946
rect 675 942 743 946
rect 747 942 767 946
rect 771 942 855 946
rect 859 942 863 946
rect 867 942 959 946
rect 963 942 967 946
rect 971 942 1047 946
rect 1051 942 1071 946
rect 1075 942 1135 946
rect 1139 942 1175 946
rect 1179 942 1223 946
rect 1227 942 1287 946
rect 1291 942 1327 946
rect 1331 942 1339 946
rect 91 941 1339 942
rect 1345 946 2618 947
rect 1345 942 1367 946
rect 1371 942 1415 946
rect 1419 942 1503 946
rect 1507 942 1535 946
rect 1539 942 1599 946
rect 1603 942 1671 946
rect 1675 942 1711 946
rect 1715 942 1807 946
rect 1811 942 1823 946
rect 1827 942 1935 946
rect 1939 942 2039 946
rect 2043 942 2055 946
rect 2059 942 2135 946
rect 2139 942 2167 946
rect 2171 942 2231 946
rect 2235 942 2271 946
rect 2275 942 2319 946
rect 2323 942 2367 946
rect 2371 942 2399 946
rect 2403 942 2463 946
rect 2467 942 2479 946
rect 2483 942 2543 946
rect 2547 942 2583 946
rect 2587 942 2618 946
rect 1345 941 2618 942
rect 96 881 97 887
rect 103 886 1351 887
rect 103 882 111 886
rect 115 882 143 886
rect 147 882 183 886
rect 187 882 199 886
rect 203 882 239 886
rect 243 882 271 886
rect 275 882 303 886
rect 307 882 359 886
rect 363 882 375 886
rect 379 882 455 886
rect 459 882 543 886
rect 547 882 551 886
rect 555 882 639 886
rect 643 882 655 886
rect 659 882 743 886
rect 747 882 751 886
rect 755 882 847 886
rect 851 882 855 886
rect 859 882 943 886
rect 947 882 967 886
rect 971 882 1031 886
rect 1035 882 1087 886
rect 1091 882 1119 886
rect 1123 882 1207 886
rect 1211 882 1215 886
rect 1219 882 1271 886
rect 1275 882 1327 886
rect 1331 882 1351 886
rect 103 881 1351 882
rect 1357 886 2630 887
rect 1357 882 1367 886
rect 1371 882 1399 886
rect 1403 882 1455 886
rect 1459 882 1519 886
rect 1523 882 1607 886
rect 1611 882 1655 886
rect 1659 882 1695 886
rect 1699 882 1791 886
rect 1795 882 1895 886
rect 1899 882 1919 886
rect 1923 882 1999 886
rect 2003 882 2039 886
rect 2043 882 2103 886
rect 2107 882 2151 886
rect 2155 882 2207 886
rect 2211 882 2255 886
rect 2259 882 2311 886
rect 2315 882 2351 886
rect 2355 882 2423 886
rect 2427 882 2447 886
rect 2451 882 2527 886
rect 2531 882 2583 886
rect 2587 882 2630 886
rect 1357 881 2630 882
rect 1338 826 2618 827
rect 1338 823 1367 826
rect 84 817 85 823
rect 91 822 1339 823
rect 91 818 111 822
rect 115 818 199 822
rect 203 818 255 822
rect 259 818 319 822
rect 323 818 383 822
rect 387 818 391 822
rect 395 818 439 822
rect 443 818 471 822
rect 475 818 495 822
rect 499 818 559 822
rect 563 818 631 822
rect 635 818 655 822
rect 659 818 703 822
rect 707 818 759 822
rect 763 818 783 822
rect 787 818 871 822
rect 875 818 959 822
rect 963 818 983 822
rect 987 818 1047 822
rect 1051 818 1103 822
rect 1107 818 1135 822
rect 1139 818 1223 822
rect 1227 818 1231 822
rect 1235 818 1327 822
rect 1331 818 1339 822
rect 91 817 1339 818
rect 1345 822 1367 823
rect 1371 822 1415 826
rect 1419 822 1471 826
rect 1475 822 1527 826
rect 1531 822 1535 826
rect 1539 822 1583 826
rect 1587 822 1623 826
rect 1627 822 1639 826
rect 1643 822 1695 826
rect 1699 822 1711 826
rect 1715 822 1751 826
rect 1755 822 1807 826
rect 1811 822 1879 826
rect 1883 822 1911 826
rect 1915 822 1959 826
rect 1963 822 2015 826
rect 2019 822 2055 826
rect 2059 822 2119 826
rect 2123 822 2167 826
rect 2171 822 2223 826
rect 2227 822 2295 826
rect 2299 822 2327 826
rect 2331 822 2431 826
rect 2435 822 2439 826
rect 2443 822 2543 826
rect 2547 822 2583 826
rect 2587 822 2618 826
rect 1345 821 2618 822
rect 1345 817 1346 821
rect 96 761 97 767
rect 103 766 1351 767
rect 103 762 111 766
rect 115 762 367 766
rect 371 762 383 766
rect 387 762 423 766
rect 427 762 439 766
rect 443 762 479 766
rect 483 762 495 766
rect 499 762 543 766
rect 547 762 559 766
rect 563 762 615 766
rect 619 762 631 766
rect 635 762 687 766
rect 691 762 711 766
rect 715 762 767 766
rect 771 762 791 766
rect 795 762 855 766
rect 859 762 871 766
rect 875 762 943 766
rect 947 762 951 766
rect 955 762 1031 766
rect 1035 762 1039 766
rect 1043 762 1119 766
rect 1123 762 1127 766
rect 1131 762 1207 766
rect 1211 762 1327 766
rect 1331 762 1351 766
rect 103 761 1351 762
rect 1357 763 1358 767
rect 1357 762 2630 763
rect 1357 761 1367 762
rect 1350 758 1367 761
rect 1371 758 1511 762
rect 1515 758 1567 762
rect 1571 758 1623 762
rect 1627 758 1647 762
rect 1651 758 1679 762
rect 1683 758 1703 762
rect 1707 758 1735 762
rect 1739 758 1759 762
rect 1763 758 1791 762
rect 1795 758 1815 762
rect 1819 758 1863 762
rect 1867 758 1871 762
rect 1875 758 1927 762
rect 1931 758 1943 762
rect 1947 758 1991 762
rect 1995 758 2039 762
rect 2043 758 2063 762
rect 2067 758 2143 762
rect 2147 758 2151 762
rect 2155 758 2231 762
rect 2235 758 2279 762
rect 2283 758 2335 762
rect 2339 758 2415 762
rect 2419 758 2439 762
rect 2443 758 2527 762
rect 2531 758 2583 762
rect 2587 758 2630 762
rect 1350 757 2630 758
rect 84 705 85 711
rect 91 710 1339 711
rect 91 706 111 710
rect 115 706 343 710
rect 347 706 399 710
rect 403 706 415 710
rect 419 706 455 710
rect 459 706 487 710
rect 491 706 511 710
rect 515 706 559 710
rect 563 706 575 710
rect 579 706 631 710
rect 635 706 647 710
rect 651 706 695 710
rect 699 706 727 710
rect 731 706 759 710
rect 763 706 807 710
rect 811 706 823 710
rect 827 706 887 710
rect 891 706 951 710
rect 955 706 967 710
rect 971 706 1023 710
rect 1027 706 1055 710
rect 1059 706 1143 710
rect 1147 706 1327 710
rect 1331 706 1339 710
rect 91 705 1339 706
rect 1345 705 1346 711
rect 1338 703 1346 705
rect 1338 697 1339 703
rect 1345 702 2611 703
rect 1345 698 1367 702
rect 1371 698 1663 702
rect 1667 698 1719 702
rect 1723 698 1735 702
rect 1739 698 1775 702
rect 1779 698 1791 702
rect 1795 698 1831 702
rect 1835 698 1855 702
rect 1859 698 1887 702
rect 1891 698 1919 702
rect 1923 698 1943 702
rect 1947 698 1991 702
rect 1995 698 2007 702
rect 2011 698 2063 702
rect 2067 698 2079 702
rect 2083 698 2127 702
rect 2131 698 2159 702
rect 2163 698 2199 702
rect 2203 698 2247 702
rect 2251 698 2271 702
rect 2275 698 2343 702
rect 2347 698 2351 702
rect 2355 698 2415 702
rect 2419 698 2455 702
rect 2459 698 2487 702
rect 2491 698 2543 702
rect 2547 698 2583 702
rect 2587 698 2611 702
rect 1345 697 2611 698
rect 2617 697 2618 703
rect 96 645 97 651
rect 103 650 1351 651
rect 103 646 111 650
rect 115 646 231 650
rect 235 646 295 650
rect 299 646 327 650
rect 331 646 359 650
rect 363 646 399 650
rect 403 646 423 650
rect 427 646 471 650
rect 475 646 479 650
rect 483 646 535 650
rect 539 646 543 650
rect 547 646 599 650
rect 603 646 615 650
rect 619 646 663 650
rect 667 646 679 650
rect 683 646 727 650
rect 731 646 743 650
rect 747 646 791 650
rect 795 646 807 650
rect 811 646 855 650
rect 859 646 871 650
rect 875 646 919 650
rect 923 646 935 650
rect 939 646 1007 650
rect 1011 646 1327 650
rect 1331 646 1351 650
rect 103 645 1351 646
rect 1357 645 1358 651
rect 1350 643 1358 645
rect 1350 637 1351 643
rect 1357 642 2623 643
rect 1357 638 1367 642
rect 1371 638 1615 642
rect 1619 638 1679 642
rect 1683 638 1719 642
rect 1723 638 1759 642
rect 1763 638 1775 642
rect 1779 638 1839 642
rect 1843 638 1903 642
rect 1907 638 1927 642
rect 1931 638 1975 642
rect 1979 638 2015 642
rect 2019 638 2047 642
rect 2051 638 2095 642
rect 2099 638 2111 642
rect 2115 638 2175 642
rect 2179 638 2183 642
rect 2187 638 2255 642
rect 2259 638 2327 642
rect 2331 638 2399 642
rect 2403 638 2471 642
rect 2475 638 2527 642
rect 2531 638 2583 642
rect 2587 638 2623 642
rect 1357 637 2623 638
rect 2629 637 2630 643
rect 84 581 85 587
rect 91 586 1339 587
rect 91 582 111 586
rect 115 582 191 586
rect 195 582 247 586
rect 251 582 279 586
rect 283 582 311 586
rect 315 582 367 586
rect 371 582 375 586
rect 379 582 439 586
rect 443 582 463 586
rect 467 582 495 586
rect 499 582 551 586
rect 555 582 559 586
rect 563 582 615 586
rect 619 582 647 586
rect 651 582 679 586
rect 683 582 735 586
rect 739 582 743 586
rect 747 582 807 586
rect 811 582 815 586
rect 819 582 871 586
rect 875 582 887 586
rect 891 582 935 586
rect 939 582 967 586
rect 971 582 1047 586
rect 1051 582 1127 586
rect 1131 582 1327 586
rect 1331 582 1339 586
rect 91 581 1339 582
rect 1345 581 1346 587
rect 1338 579 1346 581
rect 1338 573 1339 579
rect 1345 578 2611 579
rect 1345 574 1367 578
rect 1371 574 1511 578
rect 1515 574 1575 578
rect 1579 574 1631 578
rect 1635 574 1655 578
rect 1659 574 1695 578
rect 1699 574 1735 578
rect 1739 574 1775 578
rect 1779 574 1823 578
rect 1827 574 1855 578
rect 1859 574 1911 578
rect 1915 574 1943 578
rect 1947 574 1999 578
rect 2003 574 2031 578
rect 2035 574 2087 578
rect 2091 574 2111 578
rect 2115 574 2175 578
rect 2179 574 2191 578
rect 2195 574 2271 578
rect 2275 574 2343 578
rect 2347 574 2367 578
rect 2371 574 2415 578
rect 2419 574 2463 578
rect 2467 574 2487 578
rect 2491 574 2543 578
rect 2547 574 2583 578
rect 2587 574 2611 578
rect 1345 573 2611 574
rect 2617 573 2618 579
rect 96 521 97 527
rect 103 526 1351 527
rect 103 522 111 526
rect 115 522 143 526
rect 147 522 175 526
rect 179 522 207 526
rect 211 522 263 526
rect 267 522 311 526
rect 315 522 351 526
rect 355 522 431 526
rect 435 522 447 526
rect 451 522 543 526
rect 547 522 551 526
rect 555 522 631 526
rect 635 522 671 526
rect 675 522 719 526
rect 723 522 791 526
rect 795 522 799 526
rect 803 522 871 526
rect 875 522 903 526
rect 907 522 951 526
rect 955 522 1007 526
rect 1011 522 1031 526
rect 1035 522 1103 526
rect 1107 522 1111 526
rect 1115 522 1199 526
rect 1203 522 1271 526
rect 1275 522 1327 526
rect 1331 522 1351 526
rect 103 521 1351 522
rect 1357 521 1358 527
rect 1350 519 1358 521
rect 1350 513 1351 519
rect 1357 518 2623 519
rect 1357 514 1367 518
rect 1371 514 1399 518
rect 1403 514 1455 518
rect 1459 514 1495 518
rect 1499 514 1519 518
rect 1523 514 1559 518
rect 1563 514 1607 518
rect 1611 514 1639 518
rect 1643 514 1695 518
rect 1699 514 1719 518
rect 1723 514 1791 518
rect 1795 514 1807 518
rect 1811 514 1887 518
rect 1891 514 1895 518
rect 1899 514 1983 518
rect 1987 514 2071 518
rect 2075 514 2087 518
rect 2091 514 2159 518
rect 2163 514 2199 518
rect 2203 514 2255 518
rect 2259 514 2311 518
rect 2315 514 2351 518
rect 2355 514 2431 518
rect 2435 514 2447 518
rect 2451 514 2527 518
rect 2531 514 2583 518
rect 2587 514 2623 518
rect 1357 513 2623 514
rect 2629 513 2630 519
rect 84 461 85 467
rect 91 466 1339 467
rect 91 462 111 466
rect 115 462 159 466
rect 163 462 223 466
rect 227 462 319 466
rect 323 462 327 466
rect 331 462 423 466
rect 427 462 447 466
rect 451 462 535 466
rect 539 462 567 466
rect 571 462 639 466
rect 643 462 687 466
rect 691 462 743 466
rect 747 462 807 466
rect 811 462 839 466
rect 843 462 919 466
rect 923 462 927 466
rect 931 462 1007 466
rect 1011 462 1023 466
rect 1027 462 1079 466
rect 1083 462 1119 466
rect 1123 462 1151 466
rect 1155 462 1215 466
rect 1219 462 1231 466
rect 1235 462 1287 466
rect 1291 462 1327 466
rect 1331 462 1339 466
rect 91 461 1339 462
rect 1345 461 1346 467
rect 1338 449 1339 455
rect 1345 454 2611 455
rect 1345 450 1367 454
rect 1371 450 1415 454
rect 1419 450 1471 454
rect 1475 450 1487 454
rect 1491 450 1535 454
rect 1539 450 1575 454
rect 1579 450 1623 454
rect 1627 450 1663 454
rect 1667 450 1711 454
rect 1715 450 1759 454
rect 1763 450 1807 454
rect 1811 450 1863 454
rect 1867 450 1903 454
rect 1907 450 1975 454
rect 1979 450 1999 454
rect 2003 450 2103 454
rect 2107 450 2111 454
rect 2115 450 2215 454
rect 2219 450 2255 454
rect 2259 450 2327 454
rect 2331 450 2407 454
rect 2411 450 2447 454
rect 2451 450 2543 454
rect 2547 450 2583 454
rect 2587 450 2611 454
rect 1345 449 2611 450
rect 2617 449 2618 455
rect 96 397 97 403
rect 103 402 1351 403
rect 103 398 111 402
rect 115 398 143 402
rect 147 398 207 402
rect 211 398 303 402
rect 307 398 399 402
rect 403 398 407 402
rect 411 398 495 402
rect 499 398 519 402
rect 523 398 583 402
rect 587 398 623 402
rect 627 398 671 402
rect 675 398 727 402
rect 731 398 751 402
rect 755 398 823 402
rect 827 398 895 402
rect 899 398 911 402
rect 915 398 967 402
rect 971 398 991 402
rect 995 398 1047 402
rect 1051 398 1063 402
rect 1067 398 1135 402
rect 1139 398 1215 402
rect 1219 398 1271 402
rect 1275 398 1327 402
rect 1331 398 1351 402
rect 103 397 1351 398
rect 1357 397 1358 403
rect 1350 395 1358 397
rect 1350 389 1351 395
rect 1357 394 2623 395
rect 1357 390 1367 394
rect 1371 390 1399 394
rect 1403 390 1455 394
rect 1459 390 1471 394
rect 1475 390 1511 394
rect 1515 390 1559 394
rect 1563 390 1567 394
rect 1571 390 1631 394
rect 1635 390 1647 394
rect 1651 390 1695 394
rect 1699 390 1743 394
rect 1747 390 1759 394
rect 1763 390 1839 394
rect 1843 390 1847 394
rect 1851 390 1943 394
rect 1947 390 1959 394
rect 1963 390 2071 394
rect 2075 390 2095 394
rect 2099 390 2215 394
rect 2219 390 2239 394
rect 2243 390 2367 394
rect 2371 390 2391 394
rect 2395 390 2527 394
rect 2531 390 2583 394
rect 2587 390 2623 394
rect 1357 389 2623 390
rect 2629 389 2630 395
rect 84 337 85 343
rect 91 342 1339 343
rect 91 338 111 342
rect 115 338 159 342
rect 163 338 223 342
rect 227 338 311 342
rect 315 338 319 342
rect 323 338 391 342
rect 395 338 415 342
rect 419 338 471 342
rect 475 338 511 342
rect 515 338 543 342
rect 547 338 599 342
rect 603 338 607 342
rect 611 338 671 342
rect 675 338 687 342
rect 691 338 735 342
rect 739 338 767 342
rect 771 338 799 342
rect 803 338 839 342
rect 843 338 863 342
rect 867 338 911 342
rect 915 338 935 342
rect 939 338 983 342
rect 987 338 1063 342
rect 1067 338 1327 342
rect 1331 338 1339 342
rect 91 337 1339 338
rect 1345 337 1346 343
rect 1338 335 1346 337
rect 1338 329 1339 335
rect 1345 334 2611 335
rect 1345 330 1367 334
rect 1371 330 1415 334
rect 1419 330 1471 334
rect 1475 330 1527 334
rect 1531 330 1583 334
rect 1587 330 1607 334
rect 1611 330 1647 334
rect 1651 330 1663 334
rect 1667 330 1711 334
rect 1715 330 1719 334
rect 1723 330 1775 334
rect 1779 330 1831 334
rect 1835 330 1855 334
rect 1859 330 1887 334
rect 1891 330 1951 334
rect 1955 330 1959 334
rect 1963 330 2031 334
rect 2035 330 2087 334
rect 2091 330 2119 334
rect 2123 330 2223 334
rect 2227 330 2231 334
rect 2235 330 2335 334
rect 2339 330 2383 334
rect 2387 330 2447 334
rect 2451 330 2543 334
rect 2547 330 2583 334
rect 2587 330 2611 334
rect 1345 329 2611 330
rect 2617 329 2618 335
rect 96 273 97 279
rect 103 278 1351 279
rect 103 274 111 278
rect 115 274 143 278
rect 147 274 207 278
rect 211 274 231 278
rect 235 274 295 278
rect 299 274 335 278
rect 339 274 375 278
rect 379 274 431 278
rect 435 274 455 278
rect 459 274 519 278
rect 523 274 527 278
rect 531 274 591 278
rect 595 274 599 278
rect 603 274 655 278
rect 659 274 679 278
rect 683 274 719 278
rect 723 274 751 278
rect 755 274 783 278
rect 787 274 815 278
rect 819 274 847 278
rect 851 274 887 278
rect 891 274 919 278
rect 923 274 959 278
rect 963 274 1031 278
rect 1035 274 1327 278
rect 1331 274 1351 278
rect 103 273 1351 274
rect 1357 275 1358 279
rect 1357 274 2630 275
rect 1357 273 1367 274
rect 1350 270 1367 273
rect 1371 270 1591 274
rect 1595 270 1647 274
rect 1651 270 1703 274
rect 1707 270 1727 274
rect 1731 270 1759 274
rect 1763 270 1783 274
rect 1787 270 1815 274
rect 1819 270 1839 274
rect 1843 270 1871 274
rect 1875 270 1895 274
rect 1899 270 1935 274
rect 1939 270 1951 274
rect 1955 270 2007 274
rect 2011 270 2015 274
rect 2019 270 2071 274
rect 2075 270 2103 274
rect 2107 270 2143 274
rect 2147 270 2207 274
rect 2211 270 2231 274
rect 2235 270 2319 274
rect 2323 270 2335 274
rect 2339 270 2431 274
rect 2435 270 2439 274
rect 2443 270 2527 274
rect 2531 270 2583 274
rect 2587 270 2630 274
rect 1350 269 2630 270
rect 84 213 85 219
rect 91 218 1339 219
rect 91 214 111 218
rect 115 214 159 218
rect 163 214 167 218
rect 171 214 247 218
rect 251 214 255 218
rect 259 214 351 218
rect 355 214 447 218
rect 451 214 535 218
rect 539 214 551 218
rect 555 214 615 218
rect 619 214 655 218
rect 659 214 695 218
rect 699 214 751 218
rect 755 214 767 218
rect 771 214 831 218
rect 835 214 847 218
rect 851 214 903 218
rect 907 214 935 218
rect 939 214 975 218
rect 979 214 1023 218
rect 1027 214 1047 218
rect 1051 214 1111 218
rect 1115 214 1199 218
rect 1203 214 1327 218
rect 1331 214 1339 218
rect 91 213 1339 214
rect 1345 218 2618 219
rect 1345 214 1367 218
rect 1371 214 1463 218
rect 1467 214 1535 218
rect 1539 214 1623 218
rect 1627 214 1719 218
rect 1723 214 1743 218
rect 1747 214 1799 218
rect 1803 214 1823 218
rect 1827 214 1855 218
rect 1859 214 1911 218
rect 1915 214 1927 218
rect 1931 214 1967 218
rect 1971 214 2023 218
rect 2027 214 2031 218
rect 2035 214 2087 218
rect 2091 214 2135 218
rect 2139 214 2159 218
rect 2163 214 2239 218
rect 2243 214 2247 218
rect 2251 214 2343 218
rect 2347 214 2351 218
rect 2355 214 2455 218
rect 2459 214 2543 218
rect 2547 214 2583 218
rect 2587 214 2618 218
rect 1345 213 2618 214
rect 1350 141 1351 147
rect 1357 146 2623 147
rect 1357 142 1367 146
rect 1371 142 1399 146
rect 1403 142 1447 146
rect 1451 142 1455 146
rect 1459 142 1511 146
rect 1515 142 1519 146
rect 1523 142 1567 146
rect 1571 142 1607 146
rect 1611 142 1639 146
rect 1643 142 1703 146
rect 1707 142 1719 146
rect 1723 142 1799 146
rect 1803 142 1807 146
rect 1811 142 1879 146
rect 1883 142 1911 146
rect 1915 142 1959 146
rect 1963 142 2015 146
rect 2019 142 2031 146
rect 2035 142 2103 146
rect 2107 142 2119 146
rect 2123 142 2167 146
rect 2171 142 2223 146
rect 2227 142 2231 146
rect 2235 142 2295 146
rect 2299 142 2327 146
rect 2331 142 2359 146
rect 2363 142 2415 146
rect 2419 142 2439 146
rect 2443 142 2471 146
rect 2475 142 2527 146
rect 2531 142 2583 146
rect 2587 142 2623 146
rect 1357 141 2623 142
rect 2629 141 2630 147
rect 1350 139 1358 141
rect 96 133 97 139
rect 103 138 1351 139
rect 103 134 111 138
rect 115 134 143 138
rect 147 134 151 138
rect 155 134 199 138
rect 203 134 239 138
rect 243 134 255 138
rect 259 134 311 138
rect 315 134 335 138
rect 339 134 367 138
rect 371 134 423 138
rect 427 134 431 138
rect 435 134 479 138
rect 483 134 535 138
rect 539 134 607 138
rect 611 134 639 138
rect 643 134 671 138
rect 675 134 735 138
rect 739 134 799 138
rect 803 134 831 138
rect 835 134 855 138
rect 859 134 911 138
rect 915 134 919 138
rect 923 134 975 138
rect 979 134 1007 138
rect 1011 134 1039 138
rect 1043 134 1095 138
rect 1099 134 1103 138
rect 1107 134 1159 138
rect 1163 134 1183 138
rect 1187 134 1215 138
rect 1219 134 1271 138
rect 1275 134 1327 138
rect 1331 134 1351 138
rect 103 133 1351 134
rect 1357 133 1358 139
rect 1338 85 1339 91
rect 1345 90 2611 91
rect 1345 86 1367 90
rect 1371 86 1415 90
rect 1419 86 1471 90
rect 1475 86 1527 90
rect 1531 86 1583 90
rect 1587 86 1655 90
rect 1659 86 1735 90
rect 1739 86 1815 90
rect 1819 86 1895 90
rect 1899 86 1975 90
rect 1979 86 2047 90
rect 2051 86 2119 90
rect 2123 86 2183 90
rect 2187 86 2247 90
rect 2251 86 2311 90
rect 2315 86 2375 90
rect 2379 86 2431 90
rect 2435 86 2487 90
rect 2491 86 2543 90
rect 2547 86 2583 90
rect 2587 86 2611 90
rect 1345 85 2611 86
rect 2617 85 2618 91
rect 1338 83 1346 85
rect 84 77 85 83
rect 91 82 1339 83
rect 91 78 111 82
rect 115 78 159 82
rect 163 78 215 82
rect 219 78 271 82
rect 275 78 327 82
rect 331 78 383 82
rect 387 78 439 82
rect 443 78 495 82
rect 499 78 551 82
rect 555 78 623 82
rect 627 78 687 82
rect 691 78 751 82
rect 755 78 815 82
rect 819 78 871 82
rect 875 78 927 82
rect 931 78 991 82
rect 995 78 1055 82
rect 1059 78 1119 82
rect 1123 78 1175 82
rect 1179 78 1231 82
rect 1235 78 1287 82
rect 1291 78 1327 82
rect 1331 78 1339 82
rect 91 77 1339 78
rect 1345 77 1346 83
<< m5c >>
rect 85 2657 91 2663
rect 1339 2657 1345 2663
rect 1339 2611 1345 2617
rect 97 2601 103 2607
rect 1351 2601 1357 2607
rect 2611 2605 2617 2611
rect 1351 2549 1357 2555
rect 2623 2549 2629 2555
rect 85 2533 91 2539
rect 1339 2533 1345 2539
rect 1339 2489 1345 2495
rect 2611 2489 2617 2495
rect 97 2469 103 2475
rect 1351 2469 1357 2475
rect 1351 2425 1357 2431
rect 2623 2425 2629 2431
rect 85 2405 91 2411
rect 1339 2405 1345 2411
rect 1339 2365 1345 2371
rect 2611 2365 2617 2371
rect 97 2341 103 2347
rect 1351 2341 1357 2347
rect 1351 2309 1357 2315
rect 2623 2309 2629 2315
rect 85 2277 91 2283
rect 1339 2277 1345 2283
rect 1339 2253 1345 2259
rect 2611 2253 2617 2259
rect 97 2217 103 2223
rect 1351 2217 1357 2223
rect 1351 2193 1357 2199
rect 2623 2193 2629 2199
rect 85 2153 91 2159
rect 1339 2153 1345 2159
rect 1339 2137 1345 2143
rect 2611 2137 2617 2143
rect 97 2085 103 2091
rect 1351 2085 1357 2091
rect 85 2021 91 2027
rect 1339 2021 1345 2027
rect 97 1965 103 1971
rect 1351 1965 1357 1971
rect 85 1909 91 1915
rect 1339 1909 1345 1915
rect 97 1849 103 1855
rect 1351 1849 1357 1855
rect 85 1785 91 1791
rect 1339 1785 1345 1791
rect 97 1729 103 1735
rect 1351 1729 1357 1735
rect 1351 1721 1357 1727
rect 2623 1721 2629 1727
rect 85 1669 91 1675
rect 1339 1669 1345 1675
rect 97 1613 103 1619
rect 1351 1613 1357 1619
rect 1351 1597 1357 1603
rect 2623 1597 2629 1603
rect 85 1553 91 1559
rect 1339 1553 1345 1559
rect 1339 1537 1345 1543
rect 2611 1537 2617 1543
rect 97 1497 103 1503
rect 1351 1497 1357 1503
rect 1351 1473 1357 1479
rect 2623 1473 2629 1479
rect 85 1437 91 1443
rect 1339 1437 1345 1443
rect 1339 1413 1345 1419
rect 2611 1413 2617 1419
rect 97 1373 103 1379
rect 1351 1373 1357 1379
rect 1351 1357 1357 1363
rect 2623 1357 2629 1363
rect 85 1309 91 1315
rect 1339 1309 1345 1315
rect 1339 1301 1345 1307
rect 2611 1301 2617 1307
rect 97 1249 103 1255
rect 1351 1249 1357 1255
rect 1351 1241 1357 1247
rect 2623 1241 2629 1247
rect 85 1189 91 1195
rect 1339 1189 1345 1195
rect 1339 1177 1345 1183
rect 2611 1177 2617 1183
rect 97 1125 103 1131
rect 1351 1125 1357 1131
rect 85 1065 91 1071
rect 1339 1065 1345 1071
rect 97 1005 103 1011
rect 1351 1005 1357 1011
rect 85 941 91 947
rect 1339 941 1345 947
rect 97 881 103 887
rect 1351 881 1357 887
rect 85 817 91 823
rect 1339 817 1345 823
rect 97 761 103 767
rect 1351 761 1357 767
rect 85 705 91 711
rect 1339 705 1345 711
rect 1339 697 1345 703
rect 2611 697 2617 703
rect 97 645 103 651
rect 1351 645 1357 651
rect 1351 637 1357 643
rect 2623 637 2629 643
rect 85 581 91 587
rect 1339 581 1345 587
rect 1339 573 1345 579
rect 2611 573 2617 579
rect 97 521 103 527
rect 1351 521 1357 527
rect 1351 513 1357 519
rect 2623 513 2629 519
rect 85 461 91 467
rect 1339 461 1345 467
rect 1339 449 1345 455
rect 2611 449 2617 455
rect 97 397 103 403
rect 1351 397 1357 403
rect 1351 389 1357 395
rect 2623 389 2629 395
rect 85 337 91 343
rect 1339 337 1345 343
rect 1339 329 1345 335
rect 2611 329 2617 335
rect 97 273 103 279
rect 1351 273 1357 279
rect 85 213 91 219
rect 1339 213 1345 219
rect 1351 141 1357 147
rect 2623 141 2629 147
rect 97 133 103 139
rect 1351 133 1357 139
rect 1339 85 1345 91
rect 2611 85 2617 91
rect 85 77 91 83
rect 1339 77 1345 83
<< m5 >>
rect 84 2663 92 2664
rect 84 2657 85 2663
rect 91 2657 92 2663
rect 84 2539 92 2657
rect 84 2533 85 2539
rect 91 2533 92 2539
rect 84 2411 92 2533
rect 84 2405 85 2411
rect 91 2405 92 2411
rect 84 2283 92 2405
rect 84 2277 85 2283
rect 91 2277 92 2283
rect 84 2159 92 2277
rect 84 2153 85 2159
rect 91 2153 92 2159
rect 84 2027 92 2153
rect 84 2021 85 2027
rect 91 2021 92 2027
rect 84 1915 92 2021
rect 84 1909 85 1915
rect 91 1909 92 1915
rect 84 1791 92 1909
rect 84 1785 85 1791
rect 91 1785 92 1791
rect 84 1675 92 1785
rect 84 1669 85 1675
rect 91 1669 92 1675
rect 84 1559 92 1669
rect 84 1553 85 1559
rect 91 1553 92 1559
rect 84 1443 92 1553
rect 84 1437 85 1443
rect 91 1437 92 1443
rect 84 1315 92 1437
rect 84 1309 85 1315
rect 91 1309 92 1315
rect 84 1195 92 1309
rect 84 1189 85 1195
rect 91 1189 92 1195
rect 84 1071 92 1189
rect 84 1065 85 1071
rect 91 1065 92 1071
rect 84 947 92 1065
rect 84 941 85 947
rect 91 941 92 947
rect 84 823 92 941
rect 84 817 85 823
rect 91 817 92 823
rect 84 711 92 817
rect 84 705 85 711
rect 91 705 92 711
rect 84 587 92 705
rect 84 581 85 587
rect 91 581 92 587
rect 84 467 92 581
rect 84 461 85 467
rect 91 461 92 467
rect 84 343 92 461
rect 84 337 85 343
rect 91 337 92 343
rect 84 219 92 337
rect 84 213 85 219
rect 91 213 92 219
rect 84 83 92 213
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 2607 104 2664
rect 96 2601 97 2607
rect 103 2601 104 2607
rect 96 2475 104 2601
rect 96 2469 97 2475
rect 103 2469 104 2475
rect 96 2347 104 2469
rect 96 2341 97 2347
rect 103 2341 104 2347
rect 96 2223 104 2341
rect 96 2217 97 2223
rect 103 2217 104 2223
rect 96 2091 104 2217
rect 96 2085 97 2091
rect 103 2085 104 2091
rect 96 1971 104 2085
rect 96 1965 97 1971
rect 103 1965 104 1971
rect 96 1855 104 1965
rect 96 1849 97 1855
rect 103 1849 104 1855
rect 96 1735 104 1849
rect 96 1729 97 1735
rect 103 1729 104 1735
rect 96 1619 104 1729
rect 96 1613 97 1619
rect 103 1613 104 1619
rect 96 1503 104 1613
rect 96 1497 97 1503
rect 103 1497 104 1503
rect 96 1379 104 1497
rect 96 1373 97 1379
rect 103 1373 104 1379
rect 96 1255 104 1373
rect 96 1249 97 1255
rect 103 1249 104 1255
rect 96 1131 104 1249
rect 96 1125 97 1131
rect 103 1125 104 1131
rect 96 1011 104 1125
rect 96 1005 97 1011
rect 103 1005 104 1011
rect 96 887 104 1005
rect 96 881 97 887
rect 103 881 104 887
rect 96 767 104 881
rect 96 761 97 767
rect 103 761 104 767
rect 96 651 104 761
rect 96 645 97 651
rect 103 645 104 651
rect 96 527 104 645
rect 96 521 97 527
rect 103 521 104 527
rect 96 403 104 521
rect 96 397 97 403
rect 103 397 104 403
rect 96 279 104 397
rect 96 273 97 279
rect 103 273 104 279
rect 96 139 104 273
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1338 2663 1346 2664
rect 1338 2657 1339 2663
rect 1345 2657 1346 2663
rect 1338 2617 1346 2657
rect 1338 2611 1339 2617
rect 1345 2611 1346 2617
rect 1338 2539 1346 2611
rect 1338 2533 1339 2539
rect 1345 2533 1346 2539
rect 1338 2495 1346 2533
rect 1338 2489 1339 2495
rect 1345 2489 1346 2495
rect 1338 2411 1346 2489
rect 1338 2405 1339 2411
rect 1345 2405 1346 2411
rect 1338 2371 1346 2405
rect 1338 2365 1339 2371
rect 1345 2365 1346 2371
rect 1338 2283 1346 2365
rect 1338 2277 1339 2283
rect 1345 2277 1346 2283
rect 1338 2259 1346 2277
rect 1338 2253 1339 2259
rect 1345 2253 1346 2259
rect 1338 2159 1346 2253
rect 1338 2153 1339 2159
rect 1345 2153 1346 2159
rect 1338 2143 1346 2153
rect 1338 2137 1339 2143
rect 1345 2137 1346 2143
rect 1338 2027 1346 2137
rect 1338 2021 1339 2027
rect 1345 2021 1346 2027
rect 1338 1915 1346 2021
rect 1338 1909 1339 1915
rect 1345 1909 1346 1915
rect 1338 1791 1346 1909
rect 1338 1785 1339 1791
rect 1345 1785 1346 1791
rect 1338 1675 1346 1785
rect 1338 1669 1339 1675
rect 1345 1669 1346 1675
rect 1338 1559 1346 1669
rect 1338 1553 1339 1559
rect 1345 1553 1346 1559
rect 1338 1543 1346 1553
rect 1338 1537 1339 1543
rect 1345 1537 1346 1543
rect 1338 1443 1346 1537
rect 1338 1437 1339 1443
rect 1345 1437 1346 1443
rect 1338 1419 1346 1437
rect 1338 1413 1339 1419
rect 1345 1413 1346 1419
rect 1338 1315 1346 1413
rect 1338 1309 1339 1315
rect 1345 1309 1346 1315
rect 1338 1307 1346 1309
rect 1338 1301 1339 1307
rect 1345 1301 1346 1307
rect 1338 1195 1346 1301
rect 1338 1189 1339 1195
rect 1345 1189 1346 1195
rect 1338 1183 1346 1189
rect 1338 1177 1339 1183
rect 1345 1177 1346 1183
rect 1338 1071 1346 1177
rect 1338 1065 1339 1071
rect 1345 1065 1346 1071
rect 1338 947 1346 1065
rect 1338 941 1339 947
rect 1345 941 1346 947
rect 1338 823 1346 941
rect 1338 817 1339 823
rect 1345 817 1346 823
rect 1338 711 1346 817
rect 1338 705 1339 711
rect 1345 705 1346 711
rect 1338 703 1346 705
rect 1338 697 1339 703
rect 1345 697 1346 703
rect 1338 587 1346 697
rect 1338 581 1339 587
rect 1345 581 1346 587
rect 1338 579 1346 581
rect 1338 573 1339 579
rect 1345 573 1346 579
rect 1338 467 1346 573
rect 1338 461 1339 467
rect 1345 461 1346 467
rect 1338 455 1346 461
rect 1338 449 1339 455
rect 1345 449 1346 455
rect 1338 343 1346 449
rect 1338 337 1339 343
rect 1345 337 1346 343
rect 1338 335 1346 337
rect 1338 329 1339 335
rect 1345 329 1346 335
rect 1338 219 1346 329
rect 1338 213 1339 219
rect 1345 213 1346 219
rect 1338 91 1346 213
rect 1338 85 1339 91
rect 1345 85 1346 91
rect 1338 83 1346 85
rect 1338 77 1339 83
rect 1345 77 1346 83
rect 1338 72 1346 77
rect 1350 2607 1358 2664
rect 1350 2601 1351 2607
rect 1357 2601 1358 2607
rect 1350 2555 1358 2601
rect 1350 2549 1351 2555
rect 1357 2549 1358 2555
rect 1350 2475 1358 2549
rect 1350 2469 1351 2475
rect 1357 2469 1358 2475
rect 1350 2431 1358 2469
rect 1350 2425 1351 2431
rect 1357 2425 1358 2431
rect 1350 2347 1358 2425
rect 1350 2341 1351 2347
rect 1357 2341 1358 2347
rect 1350 2315 1358 2341
rect 1350 2309 1351 2315
rect 1357 2309 1358 2315
rect 1350 2223 1358 2309
rect 1350 2217 1351 2223
rect 1357 2217 1358 2223
rect 1350 2199 1358 2217
rect 1350 2193 1351 2199
rect 1357 2193 1358 2199
rect 1350 2091 1358 2193
rect 1350 2085 1351 2091
rect 1357 2085 1358 2091
rect 1350 1971 1358 2085
rect 1350 1965 1351 1971
rect 1357 1965 1358 1971
rect 1350 1855 1358 1965
rect 1350 1849 1351 1855
rect 1357 1849 1358 1855
rect 1350 1735 1358 1849
rect 1350 1729 1351 1735
rect 1357 1729 1358 1735
rect 1350 1727 1358 1729
rect 1350 1721 1351 1727
rect 1357 1721 1358 1727
rect 1350 1619 1358 1721
rect 1350 1613 1351 1619
rect 1357 1613 1358 1619
rect 1350 1603 1358 1613
rect 1350 1597 1351 1603
rect 1357 1597 1358 1603
rect 1350 1503 1358 1597
rect 1350 1497 1351 1503
rect 1357 1497 1358 1503
rect 1350 1479 1358 1497
rect 1350 1473 1351 1479
rect 1357 1473 1358 1479
rect 1350 1379 1358 1473
rect 1350 1373 1351 1379
rect 1357 1373 1358 1379
rect 1350 1363 1358 1373
rect 1350 1357 1351 1363
rect 1357 1357 1358 1363
rect 1350 1255 1358 1357
rect 1350 1249 1351 1255
rect 1357 1249 1358 1255
rect 1350 1247 1358 1249
rect 1350 1241 1351 1247
rect 1357 1241 1358 1247
rect 1350 1131 1358 1241
rect 1350 1125 1351 1131
rect 1357 1125 1358 1131
rect 1350 1011 1358 1125
rect 1350 1005 1351 1011
rect 1357 1005 1358 1011
rect 1350 887 1358 1005
rect 1350 881 1351 887
rect 1357 881 1358 887
rect 1350 767 1358 881
rect 1350 761 1351 767
rect 1357 761 1358 767
rect 1350 651 1358 761
rect 1350 645 1351 651
rect 1357 645 1358 651
rect 1350 643 1358 645
rect 1350 637 1351 643
rect 1357 637 1358 643
rect 1350 527 1358 637
rect 1350 521 1351 527
rect 1357 521 1358 527
rect 1350 519 1358 521
rect 1350 513 1351 519
rect 1357 513 1358 519
rect 1350 403 1358 513
rect 1350 397 1351 403
rect 1357 397 1358 403
rect 1350 395 1358 397
rect 1350 389 1351 395
rect 1357 389 1358 395
rect 1350 279 1358 389
rect 1350 273 1351 279
rect 1357 273 1358 279
rect 1350 147 1358 273
rect 1350 141 1351 147
rect 1357 141 1358 147
rect 1350 139 1358 141
rect 1350 133 1351 139
rect 1357 133 1358 139
rect 1350 72 1358 133
rect 2610 2611 2618 2664
rect 2610 2605 2611 2611
rect 2617 2605 2618 2611
rect 2610 2495 2618 2605
rect 2610 2489 2611 2495
rect 2617 2489 2618 2495
rect 2610 2371 2618 2489
rect 2610 2365 2611 2371
rect 2617 2365 2618 2371
rect 2610 2259 2618 2365
rect 2610 2253 2611 2259
rect 2617 2253 2618 2259
rect 2610 2143 2618 2253
rect 2610 2137 2611 2143
rect 2617 2137 2618 2143
rect 2610 1543 2618 2137
rect 2610 1537 2611 1543
rect 2617 1537 2618 1543
rect 2610 1419 2618 1537
rect 2610 1413 2611 1419
rect 2617 1413 2618 1419
rect 2610 1307 2618 1413
rect 2610 1301 2611 1307
rect 2617 1301 2618 1307
rect 2610 1183 2618 1301
rect 2610 1177 2611 1183
rect 2617 1177 2618 1183
rect 2610 703 2618 1177
rect 2610 697 2611 703
rect 2617 697 2618 703
rect 2610 579 2618 697
rect 2610 573 2611 579
rect 2617 573 2618 579
rect 2610 455 2618 573
rect 2610 449 2611 455
rect 2617 449 2618 455
rect 2610 335 2618 449
rect 2610 329 2611 335
rect 2617 329 2618 335
rect 2610 91 2618 329
rect 2610 85 2611 91
rect 2617 85 2618 91
rect 2610 72 2618 85
rect 2622 2555 2630 2664
rect 2622 2549 2623 2555
rect 2629 2549 2630 2555
rect 2622 2431 2630 2549
rect 2622 2425 2623 2431
rect 2629 2425 2630 2431
rect 2622 2315 2630 2425
rect 2622 2309 2623 2315
rect 2629 2309 2630 2315
rect 2622 2199 2630 2309
rect 2622 2193 2623 2199
rect 2629 2193 2630 2199
rect 2622 1727 2630 2193
rect 2622 1721 2623 1727
rect 2629 1721 2630 1727
rect 2622 1603 2630 1721
rect 2622 1597 2623 1603
rect 2629 1597 2630 1603
rect 2622 1479 2630 1597
rect 2622 1473 2623 1479
rect 2629 1473 2630 1479
rect 2622 1363 2630 1473
rect 2622 1357 2623 1363
rect 2629 1357 2630 1363
rect 2622 1247 2630 1357
rect 2622 1241 2623 1247
rect 2629 1241 2630 1247
rect 2622 643 2630 1241
rect 2622 637 2623 643
rect 2629 637 2630 643
rect 2622 519 2630 637
rect 2622 513 2623 519
rect 2629 513 2630 519
rect 2622 395 2630 513
rect 2622 389 2623 395
rect 2629 389 2630 395
rect 2622 147 2630 389
rect 2622 141 2623 147
rect 2629 141 2630 147
rect 2622 72 2630 141
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__167
timestamp 1731220379
transform 1 0 2576 0 -1 2592
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220379
transform 1 0 1360 0 -1 2592
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220379
transform 1 0 2576 0 1 2512
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220379
transform 1 0 1360 0 1 2512
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220379
transform 1 0 2576 0 -1 2476
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220379
transform 1 0 1360 0 -1 2476
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220379
transform 1 0 2576 0 1 2388
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220379
transform 1 0 1360 0 1 2388
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220379
transform 1 0 2576 0 -1 2352
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220379
transform 1 0 1360 0 -1 2352
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220379
transform 1 0 2576 0 1 2272
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220379
transform 1 0 1360 0 1 2272
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220379
transform 1 0 2576 0 -1 2240
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220379
transform 1 0 1360 0 -1 2240
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220379
transform 1 0 2576 0 1 2156
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220379
transform 1 0 1360 0 1 2156
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220379
transform 1 0 2576 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220379
transform 1 0 1360 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220379
transform 1 0 2576 0 1 2044
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220379
transform 1 0 1360 0 1 2044
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220379
transform 1 0 2576 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220379
transform 1 0 1360 0 -1 2012
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220379
transform 1 0 2576 0 1 1928
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220379
transform 1 0 1360 0 1 1928
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220379
transform 1 0 2576 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220379
transform 1 0 1360 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220379
transform 1 0 2576 0 1 1808
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220379
transform 1 0 1360 0 1 1808
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220379
transform 1 0 2576 0 -1 1768
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220379
transform 1 0 1360 0 -1 1768
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220379
transform 1 0 2576 0 1 1684
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220379
transform 1 0 1360 0 1 1684
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220379
transform 1 0 2576 0 -1 1652
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220379
transform 1 0 1360 0 -1 1652
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220379
transform 1 0 2576 0 1 1560
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220379
transform 1 0 1360 0 1 1560
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220379
transform 1 0 2576 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220379
transform 1 0 1360 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220379
transform 1 0 2576 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220379
transform 1 0 1360 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220379
transform 1 0 2576 0 -1 1400
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220379
transform 1 0 1360 0 -1 1400
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220379
transform 1 0 2576 0 1 1320
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220379
transform 1 0 1360 0 1 1320
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220379
transform 1 0 2576 0 -1 1288
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220379
transform 1 0 1360 0 -1 1288
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220379
transform 1 0 2576 0 1 1204
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220379
transform 1 0 1360 0 1 1204
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220379
transform 1 0 2576 0 -1 1164
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220379
transform 1 0 1360 0 -1 1164
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220379
transform 1 0 2576 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220379
transform 1 0 1360 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220379
transform 1 0 2576 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220379
transform 1 0 1360 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220379
transform 1 0 2576 0 1 968
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220379
transform 1 0 1360 0 1 968
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220379
transform 1 0 2576 0 -1 928
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220379
transform 1 0 1360 0 -1 928
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220379
transform 1 0 2576 0 1 844
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220379
transform 1 0 1360 0 1 844
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220379
transform 1 0 2576 0 -1 808
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220379
transform 1 0 1360 0 -1 808
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220379
transform 1 0 2576 0 1 720
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220379
transform 1 0 1360 0 1 720
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220379
transform 1 0 2576 0 -1 684
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220379
transform 1 0 1360 0 -1 684
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220379
transform 1 0 2576 0 1 600
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220379
transform 1 0 1360 0 1 600
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220379
transform 1 0 2576 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220379
transform 1 0 1360 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220379
transform 1 0 2576 0 1 476
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220379
transform 1 0 1360 0 1 476
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220379
transform 1 0 2576 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220379
transform 1 0 1360 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220379
transform 1 0 2576 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220379
transform 1 0 1360 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220379
transform 1 0 2576 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220379
transform 1 0 1360 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220379
transform 1 0 2576 0 1 232
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220379
transform 1 0 1360 0 1 232
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220379
transform 1 0 2576 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220379
transform 1 0 1360 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220379
transform 1 0 2576 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220379
transform 1 0 1360 0 1 104
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220379
transform 1 0 1320 0 -1 2644
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220379
transform 1 0 104 0 -1 2644
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220379
transform 1 0 1320 0 1 2564
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220379
transform 1 0 104 0 1 2564
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220379
transform 1 0 1320 0 -1 2520
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220379
transform 1 0 104 0 -1 2520
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220379
transform 1 0 1320 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220379
transform 1 0 104 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220379
transform 1 0 1320 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220379
transform 1 0 104 0 -1 2392
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220379
transform 1 0 1320 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220379
transform 1 0 104 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220379
transform 1 0 1320 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220379
transform 1 0 104 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220379
transform 1 0 1320 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220379
transform 1 0 104 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220379
transform 1 0 1320 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220379
transform 1 0 104 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220379
transform 1 0 1320 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220379
transform 1 0 104 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220379
transform 1 0 1320 0 -1 2008
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220379
transform 1 0 104 0 -1 2008
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220379
transform 1 0 1320 0 1 1928
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220379
transform 1 0 104 0 1 1928
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220379
transform 1 0 1320 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220379
transform 1 0 104 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220379
transform 1 0 1320 0 1 1812
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220379
transform 1 0 104 0 1 1812
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220379
transform 1 0 1320 0 -1 1772
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220379
transform 1 0 104 0 -1 1772
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220379
transform 1 0 1320 0 1 1692
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220379
transform 1 0 104 0 1 1692
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220379
transform 1 0 1320 0 -1 1656
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220379
transform 1 0 104 0 -1 1656
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220379
transform 1 0 1320 0 1 1576
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220379
transform 1 0 104 0 1 1576
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220379
transform 1 0 1320 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220379
transform 1 0 104 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220379
transform 1 0 1320 0 1 1460
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220379
transform 1 0 104 0 1 1460
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220379
transform 1 0 1320 0 -1 1424
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220379
transform 1 0 104 0 -1 1424
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220379
transform 1 0 1320 0 1 1336
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220379
transform 1 0 104 0 1 1336
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220379
transform 1 0 1320 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220379
transform 1 0 104 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220379
transform 1 0 1320 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220379
transform 1 0 104 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220379
transform 1 0 1320 0 -1 1176
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220379
transform 1 0 104 0 -1 1176
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220379
transform 1 0 1320 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220379
transform 1 0 104 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220379
transform 1 0 1320 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220379
transform 1 0 104 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220379
transform 1 0 1320 0 1 968
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220379
transform 1 0 104 0 1 968
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220379
transform 1 0 1320 0 -1 928
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220379
transform 1 0 104 0 -1 928
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220379
transform 1 0 1320 0 1 844
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220379
transform 1 0 104 0 1 844
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220379
transform 1 0 1320 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220379
transform 1 0 104 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220379
transform 1 0 1320 0 1 724
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220379
transform 1 0 104 0 1 724
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220379
transform 1 0 1320 0 -1 692
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220379
transform 1 0 104 0 -1 692
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220379
transform 1 0 1320 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220379
transform 1 0 104 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220379
transform 1 0 1320 0 -1 568
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220379
transform 1 0 104 0 -1 568
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220379
transform 1 0 1320 0 1 484
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220379
transform 1 0 104 0 1 484
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220379
transform 1 0 1320 0 -1 448
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220379
transform 1 0 104 0 -1 448
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220379
transform 1 0 1320 0 1 360
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220379
transform 1 0 104 0 1 360
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220379
transform 1 0 1320 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220379
transform 1 0 104 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220379
transform 1 0 1320 0 1 236
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220379
transform 1 0 104 0 1 236
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220379
transform 1 0 1320 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220379
transform 1 0 104 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220379
transform 1 0 1320 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220379
transform 1 0 104 0 1 96
box 7 3 12 24
use _0_0std_0_0cells_0_0AND2X1  tst_5999_6
timestamp 1731220379
transform 1 0 2456 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5998_6
timestamp 1731220379
transform 1 0 2512 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5997_6
timestamp 1731220379
transform 1 0 2512 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5996_6
timestamp 1731220379
transform 1 0 2512 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5995_6
timestamp 1731220379
transform 1 0 2512 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5994_6
timestamp 1731220379
transform 1 0 2424 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5993_6
timestamp 1731220379
transform 1 0 2400 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5992_6
timestamp 1731220379
transform 1 0 2344 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5991_6
timestamp 1731220379
transform 1 0 2280 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5990_6
timestamp 1731220379
transform 1 0 2216 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5989_6
timestamp 1731220379
transform 1 0 2152 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5988_6
timestamp 1731220379
transform 1 0 2088 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5987_6
timestamp 1731220379
transform 1 0 2016 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5986_6
timestamp 1731220379
transform 1 0 1944 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5985_6
timestamp 1731220379
transform 1 0 1864 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5984_6
timestamp 1731220379
transform 1 0 2312 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5983_6
timestamp 1731220379
transform 1 0 2208 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5982_6
timestamp 1731220379
transform 1 0 2104 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5981_6
timestamp 1731220379
transform 1 0 2000 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5980_6
timestamp 1731220379
transform 1 0 2424 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5979_6
timestamp 1731220379
transform 1 0 2320 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5978_6
timestamp 1731220379
transform 1 0 2216 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5977_6
timestamp 1731220379
transform 1 0 2128 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5976_6
timestamp 1731220379
transform 1 0 2056 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5975_6
timestamp 1731220379
transform 1 0 1992 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5974_6
timestamp 1731220379
transform 1 0 2304 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5973_6
timestamp 1731220379
transform 1 0 2192 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5972_6
timestamp 1731220379
transform 1 0 2088 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5971_6
timestamp 1731220379
transform 1 0 2000 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5970_6
timestamp 1731220379
transform 1 0 1920 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5969_6
timestamp 1731220379
transform 1 0 2352 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5968_6
timestamp 1731220379
transform 1 0 2200 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5967_6
timestamp 1731220379
transform 1 0 2056 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5966_6
timestamp 1731220379
transform 1 0 1928 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5965_6
timestamp 1731220379
transform 1 0 1824 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5964_6
timestamp 1731220379
transform 1 0 1744 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5963_6
timestamp 1731220379
transform 1 0 1728 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5962_6
timestamp 1731220379
transform 1 0 1832 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5961_6
timestamp 1731220379
transform 1 0 1944 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5960_6
timestamp 1731220379
transform 1 0 2376 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5959_6
timestamp 1731220379
transform 1 0 2224 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5958_6
timestamp 1731220379
transform 1 0 2080 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5957_6
timestamp 1731220379
transform 1 0 2072 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5956_6
timestamp 1731220379
transform 1 0 1968 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5955_6
timestamp 1731220379
transform 1 0 1872 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5954_6
timestamp 1731220379
transform 1 0 2296 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5953_6
timestamp 1731220379
transform 1 0 2184 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5952_6
timestamp 1731220379
transform 1 0 2144 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5951_6
timestamp 1731220379
transform 1 0 2056 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5950_6
timestamp 1731220379
transform 1 0 1968 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5949_6
timestamp 1731220379
transform 1 0 2432 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5948_6
timestamp 1731220379
transform 1 0 2336 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5947_6
timestamp 1731220379
transform 1 0 2240 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5946_6
timestamp 1731220379
transform 1 0 2160 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5945_6
timestamp 1731220379
transform 1 0 2080 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5944_6
timestamp 1731220379
transform 1 0 2312 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5943_6
timestamp 1731220379
transform 1 0 2384 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5942_6
timestamp 1731220379
transform 1 0 2456 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5941_6
timestamp 1731220379
transform 1 0 2416 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5940_6
timestamp 1731220379
transform 1 0 2416 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5939_6
timestamp 1731220379
transform 1 0 2512 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5938_6
timestamp 1731220379
transform 1 0 2512 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5937_6
timestamp 1731220379
transform 1 0 2512 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5936_6
timestamp 1731220379
transform 1 0 2512 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5935_6
timestamp 1731220379
transform 1 0 2512 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5934_6
timestamp 1731220379
transform 1 0 2512 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5933_6
timestamp 1731220379
transform 1 0 2512 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5932_6
timestamp 1731220379
transform 1 0 2512 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5931_6
timestamp 1731220379
transform 1 0 2512 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5930_6
timestamp 1731220379
transform 1 0 2512 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5929_6
timestamp 1731220379
transform 1 0 2512 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5928_6
timestamp 1731220379
transform 1 0 2512 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5927_6
timestamp 1731220379
transform 1 0 2440 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5926_6
timestamp 1731220379
transform 1 0 2352 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5925_6
timestamp 1731220379
transform 1 0 2432 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5924_6
timestamp 1731220379
transform 1 0 2408 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5923_6
timestamp 1731220379
transform 1 0 2400 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5922_6
timestamp 1731220379
transform 1 0 2424 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5921_6
timestamp 1731220379
transform 1 0 2456 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5920_6
timestamp 1731220379
transform 1 0 2384 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5919_6
timestamp 1731220379
transform 1 0 2312 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5918_6
timestamp 1731220379
transform 1 0 2240 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5917_6
timestamp 1731220379
transform 1 0 2240 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5916_6
timestamp 1731220379
transform 1 0 2168 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5915_6
timestamp 1731220379
transform 1 0 2096 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5914_6
timestamp 1731220379
transform 1 0 2320 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5913_6
timestamp 1731220379
transform 1 0 2216 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5912_6
timestamp 1731220379
transform 1 0 2128 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5911_6
timestamp 1731220379
transform 1 0 2048 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5910_6
timestamp 1731220379
transform 1 0 1976 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5909_6
timestamp 1731220379
transform 1 0 2136 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5908_6
timestamp 1731220379
transform 1 0 2024 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5907_6
timestamp 1731220379
transform 1 0 1928 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5906_6
timestamp 1731220379
transform 1 0 1848 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5905_6
timestamp 1731220379
transform 1 0 2264 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5904_6
timestamp 1731220379
transform 1 0 2296 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5903_6
timestamp 1731220379
transform 1 0 2192 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5902_6
timestamp 1731220379
transform 1 0 2088 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5901_6
timestamp 1731220379
transform 1 0 1984 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5900_6
timestamp 1731220379
transform 1 0 1880 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5899_6
timestamp 1731220379
transform 1 0 1904 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5898_6
timestamp 1731220379
transform 1 0 2024 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5897_6
timestamp 1731220379
transform 1 0 2136 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5896_6
timestamp 1731220379
transform 1 0 2336 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5895_6
timestamp 1731220379
transform 1 0 2240 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5894_6
timestamp 1731220379
transform 1 0 2200 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5893_6
timestamp 1731220379
transform 1 0 2104 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5892_6
timestamp 1731220379
transform 1 0 2008 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5891_6
timestamp 1731220379
transform 1 0 2448 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5890_6
timestamp 1731220379
transform 1 0 2368 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5889_6
timestamp 1731220379
transform 1 0 2288 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5888_6
timestamp 1731220379
transform 1 0 2264 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5887_6
timestamp 1731220379
transform 1 0 2168 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5886_6
timestamp 1731220379
transform 1 0 2072 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5885_6
timestamp 1731220379
transform 1 0 1960 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5884_6
timestamp 1731220379
transform 1 0 2400 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5883_6
timestamp 1731220379
transform 1 0 2312 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5882_6
timestamp 1731220379
transform 1 0 2224 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5881_6
timestamp 1731220379
transform 1 0 2136 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5880_6
timestamp 1731220379
transform 1 0 2336 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5879_6
timestamp 1731220379
transform 1 0 2256 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5878_6
timestamp 1731220379
transform 1 0 2176 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5877_6
timestamp 1731220379
transform 1 0 2104 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5876_6
timestamp 1731220379
transform 1 0 2032 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5875_6
timestamp 1731220379
transform 1 0 2136 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5874_6
timestamp 1731220379
transform 1 0 2264 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5873_6
timestamp 1731220379
transform 1 0 2400 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5872_6
timestamp 1731220379
transform 1 0 2392 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5871_6
timestamp 1731220379
transform 1 0 2256 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5870_6
timestamp 1731220379
transform 1 0 2128 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5869_6
timestamp 1731220379
transform 1 0 2008 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5868_6
timestamp 1731220379
transform 1 0 1912 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5867_6
timestamp 1731220379
transform 1 0 2016 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5866_6
timestamp 1731220379
transform 1 0 2024 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5865_6
timestamp 1731220379
transform 1 0 1960 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5864_6
timestamp 1731220379
transform 1 0 2048 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5863_6
timestamp 1731220379
transform 1 0 1960 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5862_6
timestamp 1731220379
transform 1 0 1864 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5861_6
timestamp 1731220379
transform 1 0 1768 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5860_6
timestamp 1731220379
transform 1 0 1672 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5859_6
timestamp 1731220379
transform 1 0 1568 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5858_6
timestamp 1731220379
transform 1 0 1664 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5857_6
timestamp 1731220379
transform 1 0 1736 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5856_6
timestamp 1731220379
transform 1 0 1816 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5855_6
timestamp 1731220379
transform 1 0 1888 0 -1 1180
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5854_6
timestamp 1731220379
transform 1 0 1928 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5853_6
timestamp 1731220379
transform 1 0 1840 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5852_6
timestamp 1731220379
transform 1 0 1760 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5851_6
timestamp 1731220379
transform 1 0 1824 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5850_6
timestamp 1731220379
transform 1 0 1864 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5849_6
timestamp 1731220379
transform 1 0 2344 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5848_6
timestamp 1731220379
transform 1 0 2168 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5847_6
timestamp 1731220379
transform 1 0 2024 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5846_6
timestamp 1731220379
transform 1 0 1928 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5845_6
timestamp 1731220379
transform 1 0 1840 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5844_6
timestamp 1731220379
transform 1 0 2136 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5843_6
timestamp 1731220379
transform 1 0 2400 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5842_6
timestamp 1731220379
transform 1 0 2264 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5841_6
timestamp 1731220379
transform 1 0 2168 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5840_6
timestamp 1731220379
transform 1 0 2072 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5839_6
timestamp 1731220379
transform 1 0 1968 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5838_6
timestamp 1731220379
transform 1 0 2256 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5837_6
timestamp 1731220379
transform 1 0 2224 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5836_6
timestamp 1731220379
transform 1 0 2136 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5835_6
timestamp 1731220379
transform 1 0 2048 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5834_6
timestamp 1731220379
transform 1 0 1968 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5833_6
timestamp 1731220379
transform 1 0 2080 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5832_6
timestamp 1731220379
transform 1 0 2184 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5831_6
timestamp 1731220379
transform 1 0 2280 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5830_6
timestamp 1731220379
transform 1 0 2376 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5829_6
timestamp 1731220379
transform 1 0 2480 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5828_6
timestamp 1731220379
transform 1 0 2456 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5827_6
timestamp 1731220379
transform 1 0 2376 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5826_6
timestamp 1731220379
transform 1 0 2304 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5825_6
timestamp 1731220379
transform 1 0 2344 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5824_6
timestamp 1731220379
transform 1 0 2440 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5823_6
timestamp 1731220379
transform 1 0 2512 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5822_6
timestamp 1731220379
transform 1 0 2512 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5821_6
timestamp 1731220379
transform 1 0 2512 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5820_6
timestamp 1731220379
transform 1 0 2512 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5819_6
timestamp 1731220379
transform 1 0 2512 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5818_6
timestamp 1731220379
transform 1 0 2512 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5817_6
timestamp 1731220379
transform 1 0 2512 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5816_6
timestamp 1731220379
transform 1 0 2512 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5815_6
timestamp 1731220379
transform 1 0 2512 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5814_6
timestamp 1731220379
transform 1 0 2512 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5813_6
timestamp 1731220379
transform 1 0 2512 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5812_6
timestamp 1731220379
transform 1 0 2432 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5811_6
timestamp 1731220379
transform 1 0 2336 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5810_6
timestamp 1731220379
transform 1 0 2512 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5809_6
timestamp 1731220379
transform 1 0 2512 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5808_6
timestamp 1731220379
transform 1 0 2488 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5807_6
timestamp 1731220379
transform 1 0 2424 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5806_6
timestamp 1731220379
transform 1 0 2432 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5805_6
timestamp 1731220379
transform 1 0 2328 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5804_6
timestamp 1731220379
transform 1 0 2336 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5803_6
timestamp 1731220379
transform 1 0 2432 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5802_6
timestamp 1731220379
transform 1 0 2424 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5801_6
timestamp 1731220379
transform 1 0 2312 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5800_6
timestamp 1731220379
transform 1 0 2200 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5799_6
timestamp 1731220379
transform 1 0 2088 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5798_6
timestamp 1731220379
transform 1 0 1968 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5797_6
timestamp 1731220379
transform 1 0 2240 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5796_6
timestamp 1731220379
transform 1 0 2144 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5795_6
timestamp 1731220379
transform 1 0 2040 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5794_6
timestamp 1731220379
transform 1 0 1936 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5793_6
timestamp 1731220379
transform 1 0 2232 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5792_6
timestamp 1731220379
transform 1 0 2136 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5791_6
timestamp 1731220379
transform 1 0 2040 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5790_6
timestamp 1731220379
transform 1 0 1944 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5789_6
timestamp 1731220379
transform 1 0 2312 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5788_6
timestamp 1731220379
transform 1 0 2208 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5787_6
timestamp 1731220379
transform 1 0 2112 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5786_6
timestamp 1731220379
transform 1 0 2024 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5785_6
timestamp 1731220379
transform 1 0 1952 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5784_6
timestamp 1731220379
transform 1 0 2352 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5783_6
timestamp 1731220379
transform 1 0 2216 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5782_6
timestamp 1731220379
transform 1 0 2096 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5781_6
timestamp 1731220379
transform 1 0 1984 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5780_6
timestamp 1731220379
transform 1 0 1896 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5779_6
timestamp 1731220379
transform 1 0 1840 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5778_6
timestamp 1731220379
transform 1 0 1744 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5777_6
timestamp 1731220379
transform 1 0 1952 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5776_6
timestamp 1731220379
transform 1 0 2376 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5775_6
timestamp 1731220379
transform 1 0 2224 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5774_6
timestamp 1731220379
transform 1 0 2080 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5773_6
timestamp 1731220379
transform 1 0 2048 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5772_6
timestamp 1731220379
transform 1 0 1952 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5771_6
timestamp 1731220379
transform 1 0 1856 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5770_6
timestamp 1731220379
transform 1 0 2144 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5769_6
timestamp 1731220379
transform 1 0 2240 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5768_6
timestamp 1731220379
transform 1 0 2152 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5767_6
timestamp 1731220379
transform 1 0 2064 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5766_6
timestamp 1731220379
transform 1 0 1968 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5765_6
timestamp 1731220379
transform 1 0 2240 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5764_6
timestamp 1731220379
transform 1 0 2328 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5763_6
timestamp 1731220379
transform 1 0 2424 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5762_6
timestamp 1731220379
transform 1 0 2512 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5761_6
timestamp 1731220379
transform 1 0 2416 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5760_6
timestamp 1731220379
transform 1 0 2320 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5759_6
timestamp 1731220379
transform 1 0 2224 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5758_6
timestamp 1731220379
transform 1 0 2128 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5757_6
timestamp 1731220379
transform 1 0 2408 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5756_6
timestamp 1731220379
transform 1 0 2320 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5755_6
timestamp 1731220379
transform 1 0 2232 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5754_6
timestamp 1731220379
transform 1 0 2152 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5753_6
timestamp 1731220379
transform 1 0 2072 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5752_6
timestamp 1731220379
transform 1 0 2304 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5751_6
timestamp 1731220379
transform 1 0 2232 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5750_6
timestamp 1731220379
transform 1 0 2160 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5749_6
timestamp 1731220379
transform 1 0 2088 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5748_6
timestamp 1731220379
transform 1 0 2024 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5747_6
timestamp 1731220379
transform 1 0 2424 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5746_6
timestamp 1731220379
transform 1 0 2360 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5745_6
timestamp 1731220379
transform 1 0 2296 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5744_6
timestamp 1731220379
transform 1 0 2232 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5743_6
timestamp 1731220379
transform 1 0 2168 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5742_6
timestamp 1731220379
transform 1 0 2112 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5741_6
timestamp 1731220379
transform 1 0 2056 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5740_6
timestamp 1731220379
transform 1 0 2000 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5739_6
timestamp 1731220379
transform 1 0 1944 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5738_6
timestamp 1731220379
transform 1 0 1888 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5737_6
timestamp 1731220379
transform 1 0 1832 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5736_6
timestamp 1731220379
transform 1 0 1776 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5735_6
timestamp 1731220379
transform 1 0 1720 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5734_6
timestamp 1731220379
transform 1 0 1664 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5733_6
timestamp 1731220379
transform 1 0 1952 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5732_6
timestamp 1731220379
transform 1 0 1872 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5731_6
timestamp 1731220379
transform 1 0 1792 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5730_6
timestamp 1731220379
transform 1 0 1696 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5729_6
timestamp 1731220379
transform 1 0 1592 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5728_6
timestamp 1731220379
transform 1 0 1992 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5727_6
timestamp 1731220379
transform 1 0 1912 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5726_6
timestamp 1731220379
transform 1 0 1824 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5725_6
timestamp 1731220379
transform 1 0 1736 0 1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5724_6
timestamp 1731220379
transform 1 0 2032 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5723_6
timestamp 1731220379
transform 1 0 1928 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5722_6
timestamp 1731220379
transform 1 0 1832 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5721_6
timestamp 1731220379
transform 1 0 1736 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5720_6
timestamp 1731220379
transform 1 0 1648 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5719_6
timestamp 1731220379
transform 1 0 1576 0 -1 2140
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5718_6
timestamp 1731220379
transform 1 0 1872 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5717_6
timestamp 1731220379
transform 1 0 1768 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5716_6
timestamp 1731220379
transform 1 0 1664 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5715_6
timestamp 1731220379
transform 1 0 1568 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5714_6
timestamp 1731220379
transform 1 0 1472 0 1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5713_6
timestamp 1731220379
transform 1 0 1760 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5712_6
timestamp 1731220379
transform 1 0 1672 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5711_6
timestamp 1731220379
transform 1 0 1584 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5710_6
timestamp 1731220379
transform 1 0 1504 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5709_6
timestamp 1731220379
transform 1 0 1440 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5708_6
timestamp 1731220379
transform 1 0 1384 0 -1 2028
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5707_6
timestamp 1731220379
transform 1 0 1384 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5706_6
timestamp 1731220379
transform 1 0 1440 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5705_6
timestamp 1731220379
transform 1 0 1504 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5704_6
timestamp 1731220379
transform 1 0 1584 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5703_6
timestamp 1731220379
transform 1 0 1664 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5702_6
timestamp 1731220379
transform 1 0 1656 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5701_6
timestamp 1731220379
transform 1 0 1600 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5700_6
timestamp 1731220379
transform 1 0 1544 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5699_6
timestamp 1731220379
transform 1 0 1712 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5698_6
timestamp 1731220379
transform 1 0 1768 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5697_6
timestamp 1731220379
transform 1 0 1824 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5696_6
timestamp 1731220379
transform 1 0 1888 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5695_6
timestamp 1731220379
transform 1 0 1832 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5694_6
timestamp 1731220379
transform 1 0 1776 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5693_6
timestamp 1731220379
transform 1 0 1720 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5692_6
timestamp 1731220379
transform 1 0 1664 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5691_6
timestamp 1731220379
transform 1 0 1608 0 1 1792
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5690_6
timestamp 1731220379
transform 1 0 1848 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5689_6
timestamp 1731220379
transform 1 0 1752 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5688_6
timestamp 1731220379
transform 1 0 1664 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5687_6
timestamp 1731220379
transform 1 0 1584 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5686_6
timestamp 1731220379
transform 1 0 1504 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5685_6
timestamp 1731220379
transform 1 0 1440 0 -1 1784
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5684_6
timestamp 1731220379
transform 1 0 1824 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5683_6
timestamp 1731220379
transform 1 0 1704 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5682_6
timestamp 1731220379
transform 1 0 1584 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5681_6
timestamp 1731220379
transform 1 0 1464 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5680_6
timestamp 1731220379
transform 1 0 1384 0 1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5679_6
timestamp 1731220379
transform 1 0 1384 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5678_6
timestamp 1731220379
transform 1 0 1472 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5677_6
timestamp 1731220379
transform 1 0 1592 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5676_6
timestamp 1731220379
transform 1 0 1848 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5675_6
timestamp 1731220379
transform 1 0 1720 0 -1 1668
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5674_6
timestamp 1731220379
transform 1 0 1600 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5673_6
timestamp 1731220379
transform 1 0 1480 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5672_6
timestamp 1731220379
transform 1 0 1848 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5671_6
timestamp 1731220379
transform 1 0 1728 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5670_6
timestamp 1731220379
transform 1 0 1616 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5669_6
timestamp 1731220379
transform 1 0 1496 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5668_6
timestamp 1731220379
transform 1 0 1736 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5667_6
timestamp 1731220379
transform 1 0 1848 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5666_6
timestamp 1731220379
transform 1 0 1952 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5665_6
timestamp 1731220379
transform 1 0 1856 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5664_6
timestamp 1731220379
transform 1 0 1736 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5663_6
timestamp 1731220379
transform 1 0 1616 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5662_6
timestamp 1731220379
transform 1 0 1600 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5661_6
timestamp 1731220379
transform 1 0 1680 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5660_6
timestamp 1731220379
transform 1 0 1760 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5659_6
timestamp 1731220379
transform 1 0 1744 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5658_6
timestamp 1731220379
transform 1 0 1640 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5657_6
timestamp 1731220379
transform 1 0 1600 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5656_6
timestamp 1731220379
transform 1 0 1672 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5655_6
timestamp 1731220379
transform 1 0 1744 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5654_6
timestamp 1731220379
transform 1 0 1680 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5653_6
timestamp 1731220379
transform 1 0 1600 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5652_6
timestamp 1731220379
transform 1 0 1520 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5651_6
timestamp 1731220379
transform 1 0 1464 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5650_6
timestamp 1731220379
transform 1 0 1400 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5649_6
timestamp 1731220379
transform 1 0 1408 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5648_6
timestamp 1731220379
transform 1 0 1480 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5647_6
timestamp 1731220379
transform 1 0 1440 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5646_6
timestamp 1731220379
transform 1 0 1384 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5645_6
timestamp 1731220379
transform 1 0 1384 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5644_6
timestamp 1731220379
transform 1 0 1256 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5643_6
timestamp 1731220379
transform 1 0 1256 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5642_6
timestamp 1731220379
transform 1 0 1120 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5641_6
timestamp 1731220379
transform 1 0 1184 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5640_6
timestamp 1731220379
transform 1 0 1088 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5639_6
timestamp 1731220379
transform 1 0 992 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5638_6
timestamp 1731220379
transform 1 0 896 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5637_6
timestamp 1731220379
transform 1 0 928 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5636_6
timestamp 1731220379
transform 1 0 1120 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5635_6
timestamp 1731220379
transform 1 0 1024 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5634_6
timestamp 1731220379
transform 1 0 1016 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5633_6
timestamp 1731220379
transform 1 0 1112 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5632_6
timestamp 1731220379
transform 1 0 1216 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5631_6
timestamp 1731220379
transform 1 0 1168 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5630_6
timestamp 1731220379
transform 1 0 1064 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5629_6
timestamp 1731220379
transform 1 0 1256 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5628_6
timestamp 1731220379
transform 1 0 1256 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5627_6
timestamp 1731220379
transform 1 0 1160 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5626_6
timestamp 1731220379
transform 1 0 1064 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5625_6
timestamp 1731220379
transform 1 0 1128 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5624_6
timestamp 1731220379
transform 1 0 1056 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5623_6
timestamp 1731220379
transform 1 0 984 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5622_6
timestamp 1731220379
transform 1 0 904 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5621_6
timestamp 1731220379
transform 1 0 888 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5620_6
timestamp 1731220379
transform 1 0 800 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5619_6
timestamp 1731220379
transform 1 0 976 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5618_6
timestamp 1731220379
transform 1 0 960 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5617_6
timestamp 1731220379
transform 1 0 864 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5616_6
timestamp 1731220379
transform 1 0 776 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5615_6
timestamp 1731220379
transform 1 0 920 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5614_6
timestamp 1731220379
transform 1 0 824 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5613_6
timestamp 1731220379
transform 1 0 736 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5612_6
timestamp 1731220379
transform 1 0 664 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5611_6
timestamp 1731220379
transform 1 0 752 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5610_6
timestamp 1731220379
transform 1 0 840 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5609_6
timestamp 1731220379
transform 1 0 792 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5608_6
timestamp 1731220379
transform 1 0 688 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5607_6
timestamp 1731220379
transform 1 0 688 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5606_6
timestamp 1731220379
transform 1 0 832 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5605_6
timestamp 1731220379
transform 1 0 976 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5604_6
timestamp 1731220379
transform 1 0 1160 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5603_6
timestamp 1731220379
transform 1 0 1048 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5602_6
timestamp 1731220379
transform 1 0 944 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5601_6
timestamp 1731220379
transform 1 0 848 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5600_6
timestamp 1731220379
transform 1 0 752 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5599_6
timestamp 1731220379
transform 1 0 656 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5598_6
timestamp 1731220379
transform 1 0 1048 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5597_6
timestamp 1731220379
transform 1 0 936 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5596_6
timestamp 1731220379
transform 1 0 832 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5595_6
timestamp 1731220379
transform 1 0 736 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5594_6
timestamp 1731220379
transform 1 0 648 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5593_6
timestamp 1731220379
transform 1 0 576 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5592_6
timestamp 1731220379
transform 1 0 504 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5591_6
timestamp 1731220379
transform 1 0 560 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5590_6
timestamp 1731220379
transform 1 0 464 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5589_6
timestamp 1731220379
transform 1 0 352 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5588_6
timestamp 1731220379
transform 1 0 432 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5587_6
timestamp 1731220379
transform 1 0 352 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5586_6
timestamp 1731220379
transform 1 0 272 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5585_6
timestamp 1731220379
transform 1 0 192 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5584_6
timestamp 1731220379
transform 1 0 400 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5583_6
timestamp 1731220379
transform 1 0 552 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5582_6
timestamp 1731220379
transform 1 0 696 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5581_6
timestamp 1731220379
transform 1 0 592 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5580_6
timestamp 1731220379
transform 1 0 472 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5579_6
timestamp 1731220379
transform 1 0 344 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5578_6
timestamp 1731220379
transform 1 0 616 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5577_6
timestamp 1731220379
transform 1 0 528 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5576_6
timestamp 1731220379
transform 1 0 440 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5575_6
timestamp 1731220379
transform 1 0 360 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5574_6
timestamp 1731220379
transform 1 0 296 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5573_6
timestamp 1731220379
transform 1 0 240 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5572_6
timestamp 1731220379
transform 1 0 184 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5571_6
timestamp 1731220379
transform 1 0 128 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5570_6
timestamp 1731220379
transform 1 0 128 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5569_6
timestamp 1731220379
transform 1 0 224 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5568_6
timestamp 1731220379
transform 1 0 248 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5567_6
timestamp 1731220379
transform 1 0 128 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5566_6
timestamp 1731220379
transform 1 0 128 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5565_6
timestamp 1731220379
transform 1 0 128 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5564_6
timestamp 1731220379
transform 1 0 232 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5563_6
timestamp 1731220379
transform 1 0 200 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5562_6
timestamp 1731220379
transform 1 0 128 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5561_6
timestamp 1731220379
transform 1 0 552 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5560_6
timestamp 1731220379
transform 1 0 424 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5559_6
timestamp 1731220379
transform 1 0 304 0 -1 1556
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5558_6
timestamp 1731220379
transform 1 0 256 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5557_6
timestamp 1731220379
transform 1 0 184 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5556_6
timestamp 1731220379
transform 1 0 128 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5555_6
timestamp 1731220379
transform 1 0 576 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5554_6
timestamp 1731220379
transform 1 0 464 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5553_6
timestamp 1731220379
transform 1 0 352 0 1 1444
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5552_6
timestamp 1731220379
transform 1 0 344 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5551_6
timestamp 1731220379
transform 1 0 280 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5550_6
timestamp 1731220379
transform 1 0 224 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5549_6
timestamp 1731220379
transform 1 0 416 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5548_6
timestamp 1731220379
transform 1 0 576 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5547_6
timestamp 1731220379
transform 1 0 496 0 -1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5546_6
timestamp 1731220379
transform 1 0 456 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5545_6
timestamp 1731220379
transform 1 0 400 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5544_6
timestamp 1731220379
transform 1 0 344 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5543_6
timestamp 1731220379
transform 1 0 512 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5542_6
timestamp 1731220379
transform 1 0 576 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5541_6
timestamp 1731220379
transform 1 0 656 0 1 1320
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5540_6
timestamp 1731220379
transform 1 0 696 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5539_6
timestamp 1731220379
transform 1 0 616 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5538_6
timestamp 1731220379
transform 1 0 552 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5537_6
timestamp 1731220379
transform 1 0 496 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5536_6
timestamp 1731220379
transform 1 0 440 0 -1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5535_6
timestamp 1731220379
transform 1 0 712 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5534_6
timestamp 1731220379
transform 1 0 632 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5533_6
timestamp 1731220379
transform 1 0 560 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5532_6
timestamp 1731220379
transform 1 0 488 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5531_6
timestamp 1731220379
transform 1 0 424 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5530_6
timestamp 1731220379
transform 1 0 368 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5529_6
timestamp 1731220379
transform 1 0 640 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5528_6
timestamp 1731220379
transform 1 0 552 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5527_6
timestamp 1731220379
transform 1 0 464 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5526_6
timestamp 1731220379
transform 1 0 384 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5525_6
timestamp 1731220379
transform 1 0 312 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5524_6
timestamp 1731220379
transform 1 0 248 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5523_6
timestamp 1731220379
transform 1 0 488 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5522_6
timestamp 1731220379
transform 1 0 408 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5521_6
timestamp 1731220379
transform 1 0 328 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5520_6
timestamp 1731220379
transform 1 0 256 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5519_6
timestamp 1731220379
transform 1 0 192 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5518_6
timestamp 1731220379
transform 1 0 128 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5517_6
timestamp 1731220379
transform 1 0 552 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5516_6
timestamp 1731220379
transform 1 0 448 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5515_6
timestamp 1731220379
transform 1 0 352 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5514_6
timestamp 1731220379
transform 1 0 256 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5513_6
timestamp 1731220379
transform 1 0 184 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5512_6
timestamp 1731220379
transform 1 0 128 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5511_6
timestamp 1731220379
transform 1 0 368 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5510_6
timestamp 1731220379
transform 1 0 264 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5509_6
timestamp 1731220379
transform 1 0 184 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5508_6
timestamp 1731220379
transform 1 0 128 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5507_6
timestamp 1731220379
transform 1 0 600 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5506_6
timestamp 1731220379
transform 1 0 480 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5505_6
timestamp 1731220379
transform 1 0 256 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5504_6
timestamp 1731220379
transform 1 0 184 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5503_6
timestamp 1731220379
transform 1 0 128 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5502_6
timestamp 1731220379
transform 1 0 536 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5501_6
timestamp 1731220379
transform 1 0 440 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5500_6
timestamp 1731220379
transform 1 0 344 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5499_6
timestamp 1731220379
transform 1 0 288 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5498_6
timestamp 1731220379
transform 1 0 224 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5497_6
timestamp 1731220379
transform 1 0 168 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5496_6
timestamp 1731220379
transform 1 0 360 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5495_6
timestamp 1731220379
transform 1 0 440 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5494_6
timestamp 1731220379
transform 1 0 528 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5493_6
timestamp 1731220379
transform 1 0 464 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5492_6
timestamp 1731220379
transform 1 0 408 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5491_6
timestamp 1731220379
transform 1 0 352 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5490_6
timestamp 1731220379
transform 1 0 528 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5489_6
timestamp 1731220379
transform 1 0 600 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5488_6
timestamp 1731220379
transform 1 0 672 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5487_6
timestamp 1731220379
transform 1 0 616 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5486_6
timestamp 1731220379
transform 1 0 544 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5485_6
timestamp 1731220379
transform 1 0 480 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5484_6
timestamp 1731220379
transform 1 0 424 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5483_6
timestamp 1731220379
transform 1 0 368 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5482_6
timestamp 1731220379
transform 1 0 384 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5481_6
timestamp 1731220379
transform 1 0 312 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5480_6
timestamp 1731220379
transform 1 0 344 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5479_6
timestamp 1731220379
transform 1 0 280 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5478_6
timestamp 1731220379
transform 1 0 216 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5477_6
timestamp 1731220379
transform 1 0 160 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5476_6
timestamp 1731220379
transform 1 0 248 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5475_6
timestamp 1731220379
transform 1 0 336 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5474_6
timestamp 1731220379
transform 1 0 296 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5473_6
timestamp 1731220379
transform 1 0 192 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5472_6
timestamp 1731220379
transform 1 0 128 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5471_6
timestamp 1731220379
transform 1 0 128 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5470_6
timestamp 1731220379
transform 1 0 192 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5469_6
timestamp 1731220379
transform 1 0 288 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5468_6
timestamp 1731220379
transform 1 0 192 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5467_6
timestamp 1731220379
transform 1 0 128 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5466_6
timestamp 1731220379
transform 1 0 128 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5465_6
timestamp 1731220379
transform 1 0 192 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5464_6
timestamp 1731220379
transform 1 0 280 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5463_6
timestamp 1731220379
transform 1 0 216 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5462_6
timestamp 1731220379
transform 1 0 128 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5461_6
timestamp 1731220379
transform 1 0 136 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5460_6
timestamp 1731220379
transform 1 0 320 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5459_6
timestamp 1731220379
transform 1 0 224 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5458_6
timestamp 1731220379
transform 1 0 240 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5457_6
timestamp 1731220379
transform 1 0 184 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5456_6
timestamp 1731220379
transform 1 0 128 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5455_6
timestamp 1731220379
transform 1 0 296 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5454_6
timestamp 1731220379
transform 1 0 352 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5453_6
timestamp 1731220379
transform 1 0 408 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5452_6
timestamp 1731220379
transform 1 0 592 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5451_6
timestamp 1731220379
transform 1 0 520 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5450_6
timestamp 1731220379
transform 1 0 464 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5449_6
timestamp 1731220379
transform 1 0 416 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5448_6
timestamp 1731220379
transform 1 0 520 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5447_6
timestamp 1731220379
transform 1 0 624 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5446_6
timestamp 1731220379
transform 1 0 584 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5445_6
timestamp 1731220379
transform 1 0 504 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5444_6
timestamp 1731220379
transform 1 0 416 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5443_6
timestamp 1731220379
transform 1 0 320 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5442_6
timestamp 1731220379
transform 1 0 360 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5441_6
timestamp 1731220379
transform 1 0 512 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5440_6
timestamp 1731220379
transform 1 0 440 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5439_6
timestamp 1731220379
transform 1 0 384 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5438_6
timestamp 1731220379
transform 1 0 480 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5437_6
timestamp 1731220379
transform 1 0 568 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5436_6
timestamp 1731220379
transform 1 0 608 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5435_6
timestamp 1731220379
transform 1 0 504 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5434_6
timestamp 1731220379
transform 1 0 392 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5433_6
timestamp 1731220379
transform 1 0 288 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5432_6
timestamp 1731220379
transform 1 0 416 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5431_6
timestamp 1731220379
transform 1 0 536 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5430_6
timestamp 1731220379
transform 1 0 656 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5429_6
timestamp 1731220379
transform 1 0 616 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5428_6
timestamp 1731220379
transform 1 0 528 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5427_6
timestamp 1731220379
transform 1 0 432 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5426_6
timestamp 1731220379
transform 1 0 408 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5425_6
timestamp 1731220379
transform 1 0 464 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5424_6
timestamp 1731220379
transform 1 0 520 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5423_6
timestamp 1731220379
transform 1 0 456 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5422_6
timestamp 1731220379
transform 1 0 528 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5421_6
timestamp 1731220379
transform 1 0 600 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5420_6
timestamp 1731220379
transform 1 0 696 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5419_6
timestamp 1731220379
transform 1 0 776 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5418_6
timestamp 1731220379
transform 1 0 840 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5417_6
timestamp 1731220379
transform 1 0 752 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5416_6
timestamp 1731220379
transform 1 0 728 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5415_6
timestamp 1731220379
transform 1 0 624 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5414_6
timestamp 1731220379
transform 1 0 840 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5413_6
timestamp 1731220379
transform 1 0 952 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5412_6
timestamp 1731220379
transform 1 0 928 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5411_6
timestamp 1731220379
transform 1 0 832 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5410_6
timestamp 1731220379
transform 1 0 736 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5409_6
timestamp 1731220379
transform 1 0 640 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5408_6
timestamp 1731220379
transform 1 0 712 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5407_6
timestamp 1731220379
transform 1 0 824 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5406_6
timestamp 1731220379
transform 1 0 936 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5405_6
timestamp 1731220379
transform 1 0 848 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5404_6
timestamp 1731220379
transform 1 0 752 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5403_6
timestamp 1731220379
transform 1 0 656 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5402_6
timestamp 1731220379
transform 1 0 816 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5401_6
timestamp 1731220379
transform 1 0 728 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5400_6
timestamp 1731220379
transform 1 0 648 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5399_6
timestamp 1731220379
transform 1 0 568 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5398_6
timestamp 1731220379
transform 1 0 728 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5397_6
timestamp 1731220379
transform 1 0 816 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5396_6
timestamp 1731220379
transform 1 0 904 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5395_6
timestamp 1731220379
transform 1 0 992 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5394_6
timestamp 1731220379
transform 1 0 936 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5393_6
timestamp 1731220379
transform 1 0 1032 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5392_6
timestamp 1731220379
transform 1 0 1128 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5391_6
timestamp 1731220379
transform 1 0 1256 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5390_6
timestamp 1731220379
transform 1 0 1144 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5389_6
timestamp 1731220379
transform 1 0 1040 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5388_6
timestamp 1731220379
transform 1 0 1016 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5387_6
timestamp 1731220379
transform 1 0 1104 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5386_6
timestamp 1731220379
transform 1 0 1072 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5385_6
timestamp 1731220379
transform 1 0 1200 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5384_6
timestamp 1731220379
transform 1 0 1192 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5383_6
timestamp 1731220379
transform 1 0 1104 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5382_6
timestamp 1731220379
transform 1 0 1016 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5381_6
timestamp 1731220379
transform 1 0 928 0 -1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5380_6
timestamp 1731220379
transform 1 0 1112 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5379_6
timestamp 1731220379
transform 1 0 1024 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5378_6
timestamp 1731220379
transform 1 0 936 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5377_6
timestamp 1731220379
transform 1 0 856 0 1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5376_6
timestamp 1731220379
transform 1 0 992 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5375_6
timestamp 1731220379
transform 1 0 920 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5374_6
timestamp 1731220379
transform 1 0 856 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5373_6
timestamp 1731220379
transform 1 0 792 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5372_6
timestamp 1731220379
transform 1 0 728 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5371_6
timestamp 1731220379
transform 1 0 664 0 -1 708
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5370_6
timestamp 1731220379
transform 1 0 648 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5369_6
timestamp 1731220379
transform 1 0 584 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5368_6
timestamp 1731220379
transform 1 0 712 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5367_6
timestamp 1731220379
transform 1 0 776 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5366_6
timestamp 1731220379
transform 1 0 904 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5365_6
timestamp 1731220379
transform 1 0 840 0 1 592
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5364_6
timestamp 1731220379
transform 1 0 784 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5363_6
timestamp 1731220379
transform 1 0 704 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5362_6
timestamp 1731220379
transform 1 0 856 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5361_6
timestamp 1731220379
transform 1 0 1096 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5360_6
timestamp 1731220379
transform 1 0 1016 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5359_6
timestamp 1731220379
transform 1 0 936 0 -1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5358_6
timestamp 1731220379
transform 1 0 888 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5357_6
timestamp 1731220379
transform 1 0 776 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5356_6
timestamp 1731220379
transform 1 0 992 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5355_6
timestamp 1731220379
transform 1 0 1256 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5354_6
timestamp 1731220379
transform 1 0 1184 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5353_6
timestamp 1731220379
transform 1 0 1088 0 1 468
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5352_6
timestamp 1731220379
transform 1 0 1048 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5351_6
timestamp 1731220379
transform 1 0 976 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5350_6
timestamp 1731220379
transform 1 0 896 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5349_6
timestamp 1731220379
transform 1 0 808 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5348_6
timestamp 1731220379
transform 1 0 712 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5347_6
timestamp 1731220379
transform 1 0 1032 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5346_6
timestamp 1731220379
transform 1 0 952 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5345_6
timestamp 1731220379
transform 1 0 880 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5344_6
timestamp 1731220379
transform 1 0 808 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5343_6
timestamp 1731220379
transform 1 0 736 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5342_6
timestamp 1731220379
transform 1 0 656 0 1 344
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5341_6
timestamp 1731220379
transform 1 0 904 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5340_6
timestamp 1731220379
transform 1 0 832 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5339_6
timestamp 1731220379
transform 1 0 768 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5338_6
timestamp 1731220379
transform 1 0 704 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5337_6
timestamp 1731220379
transform 1 0 640 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5336_6
timestamp 1731220379
transform 1 0 576 0 -1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5335_6
timestamp 1731220379
transform 1 0 664 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5334_6
timestamp 1731220379
transform 1 0 736 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5333_6
timestamp 1731220379
transform 1 0 800 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5332_6
timestamp 1731220379
transform 1 0 872 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5331_6
timestamp 1731220379
transform 1 0 1016 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5330_6
timestamp 1731220379
transform 1 0 944 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5329_6
timestamp 1731220379
transform 1 0 904 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5328_6
timestamp 1731220379
transform 1 0 816 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5327_6
timestamp 1731220379
transform 1 0 720 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5326_6
timestamp 1731220379
transform 1 0 1168 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5325_6
timestamp 1731220379
transform 1 0 1080 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5324_6
timestamp 1731220379
transform 1 0 992 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5323_6
timestamp 1731220379
transform 1 0 784 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5322_6
timestamp 1731220379
transform 1 0 720 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5321_6
timestamp 1731220379
transform 1 0 656 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5320_6
timestamp 1731220379
transform 1 0 840 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5319_6
timestamp 1731220379
transform 1 0 896 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5318_6
timestamp 1731220379
transform 1 0 960 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5317_6
timestamp 1731220379
transform 1 0 1024 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5316_6
timestamp 1731220379
transform 1 0 1088 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5315_6
timestamp 1731220379
transform 1 0 1144 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5314_6
timestamp 1731220379
transform 1 0 1200 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5313_6
timestamp 1731220379
transform 1 0 1256 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5312_6
timestamp 1731220379
transform 1 0 1384 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5311_6
timestamp 1731220379
transform 1 0 1440 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5310_6
timestamp 1731220379
transform 1 0 1496 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5309_6
timestamp 1731220379
transform 1 0 1552 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5308_6
timestamp 1731220379
transform 1 0 1784 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5307_6
timestamp 1731220379
transform 1 0 1704 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5306_6
timestamp 1731220379
transform 1 0 1624 0 1 88
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5305_6
timestamp 1731220379
transform 1 0 1592 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5304_6
timestamp 1731220379
transform 1 0 1504 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5303_6
timestamp 1731220379
transform 1 0 1432 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5302_6
timestamp 1731220379
transform 1 0 1688 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5301_6
timestamp 1731220379
transform 1 0 1792 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5300_6
timestamp 1731220379
transform 1 0 1896 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5299_6
timestamp 1731220379
transform 1 0 1824 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5298_6
timestamp 1731220379
transform 1 0 1768 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5297_6
timestamp 1731220379
transform 1 0 1712 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5296_6
timestamp 1731220379
transform 1 0 1936 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5295_6
timestamp 1731220379
transform 1 0 1880 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5294_6
timestamp 1731220379
transform 1 0 1856 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5293_6
timestamp 1731220379
transform 1 0 1800 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5292_6
timestamp 1731220379
transform 1 0 1744 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5291_6
timestamp 1731220379
transform 1 0 1688 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5290_6
timestamp 1731220379
transform 1 0 1632 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5289_6
timestamp 1731220379
transform 1 0 1576 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5288_6
timestamp 1731220379
transform 1 0 1680 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5287_6
timestamp 1731220379
transform 1 0 1616 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5286_6
timestamp 1731220379
transform 1 0 1552 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5285_6
timestamp 1731220379
transform 1 0 1496 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5284_6
timestamp 1731220379
transform 1 0 1440 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5283_6
timestamp 1731220379
transform 1 0 1384 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5282_6
timestamp 1731220379
transform 1 0 1632 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5281_6
timestamp 1731220379
transform 1 0 1544 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5280_6
timestamp 1731220379
transform 1 0 1456 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5279_6
timestamp 1731220379
transform 1 0 1256 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5278_6
timestamp 1731220379
transform 1 0 1200 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5277_6
timestamp 1731220379
transform 1 0 1120 0 -1 464
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5276_6
timestamp 1731220379
transform 1 0 1384 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5275_6
timestamp 1731220379
transform 1 0 1384 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5274_6
timestamp 1731220379
transform 1 0 1440 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5273_6
timestamp 1731220379
transform 1 0 1504 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5272_6
timestamp 1731220379
transform 1 0 1776 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5271_6
timestamp 1731220379
transform 1 0 1680 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5270_6
timestamp 1731220379
transform 1 0 1592 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5269_6
timestamp 1731220379
transform 1 0 1544 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5268_6
timestamp 1731220379
transform 1 0 1480 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5267_6
timestamp 1731220379
transform 1 0 1624 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5266_6
timestamp 1731220379
transform 1 0 1880 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5265_6
timestamp 1731220379
transform 1 0 1792 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5264_6
timestamp 1731220379
transform 1 0 1704 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5263_6
timestamp 1731220379
transform 1 0 1664 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5262_6
timestamp 1731220379
transform 1 0 1600 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5261_6
timestamp 1731220379
transform 1 0 1744 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5260_6
timestamp 1731220379
transform 1 0 2000 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5259_6
timestamp 1731220379
transform 1 0 1912 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5258_6
timestamp 1731220379
transform 1 0 1824 0 1 584
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5257_6
timestamp 1731220379
transform 1 0 1824 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5256_6
timestamp 1731220379
transform 1 0 1760 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5255_6
timestamp 1731220379
transform 1 0 1704 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5254_6
timestamp 1731220379
transform 1 0 1888 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5253_6
timestamp 1731220379
transform 1 0 1912 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5252_6
timestamp 1731220379
transform 1 0 2032 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5251_6
timestamp 1731220379
transform 1 0 1960 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5250_6
timestamp 1731220379
transform 1 0 1856 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5249_6
timestamp 1731220379
transform 1 0 1800 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5248_6
timestamp 1731220379
transform 1 0 1744 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5247_6
timestamp 1731220379
transform 1 0 1688 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5246_6
timestamp 1731220379
transform 1 0 1632 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5245_6
timestamp 1731220379
transform 1 0 1776 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5244_6
timestamp 1731220379
transform 1 0 1720 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5243_6
timestamp 1731220379
transform 1 0 1664 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5242_6
timestamp 1731220379
transform 1 0 1608 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5241_6
timestamp 1731220379
transform 1 0 1552 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5240_6
timestamp 1731220379
transform 1 0 1496 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5239_6
timestamp 1731220379
transform 1 0 1776 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5238_6
timestamp 1731220379
transform 1 0 1680 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5237_6
timestamp 1731220379
transform 1 0 1592 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5236_6
timestamp 1731220379
transform 1 0 1504 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5235_6
timestamp 1731220379
transform 1 0 1440 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5234_6
timestamp 1731220379
transform 1 0 1384 0 1 828
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5233_6
timestamp 1731220379
transform 1 0 1256 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5232_6
timestamp 1731220379
transform 1 0 1192 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5231_6
timestamp 1731220379
transform 1 0 1384 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5230_6
timestamp 1731220379
transform 1 0 1504 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5229_6
timestamp 1731220379
transform 1 0 1640 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5228_6
timestamp 1731220379
transform 1 0 1776 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5227_6
timestamp 1731220379
transform 1 0 1792 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5226_6
timestamp 1731220379
transform 1 0 1680 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5225_6
timestamp 1731220379
transform 1 0 1568 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5224_6
timestamp 1731220379
transform 1 0 1472 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5223_6
timestamp 1731220379
transform 1 0 1904 0 1 952
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5222_6
timestamp 1731220379
transform 1 0 1840 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5221_6
timestamp 1731220379
transform 1 0 1720 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5220_6
timestamp 1731220379
transform 1 0 1600 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5219_6
timestamp 1731220379
transform 1 0 1480 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5218_6
timestamp 1731220379
transform 1 0 1384 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5217_6
timestamp 1731220379
transform 1 0 1464 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5216_6
timestamp 1731220379
transform 1 0 1384 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5215_6
timestamp 1731220379
transform 1 0 1256 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5214_6
timestamp 1731220379
transform 1 0 1200 0 -1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5213_6
timestamp 1731220379
transform 1 0 1384 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5212_6
timestamp 1731220379
transform 1 0 1440 0 1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5211_6
timestamp 1731220379
transform 1 0 1528 0 -1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5210_6
timestamp 1731220379
transform 1 0 1560 0 1 1304
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5209_6
timestamp 1731220379
transform 1 0 1520 0 -1 1416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5208_6
timestamp 1731220379
transform 1 0 1488 0 1 1420
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5207_6
timestamp 1731220379
transform 1 0 1384 0 -1 1540
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5206_6
timestamp 1731220379
transform 1 0 1384 0 1 1544
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5205_6
timestamp 1731220379
transform 1 0 1256 0 1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5204_6
timestamp 1731220379
transform 1 0 1256 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5203_6
timestamp 1731220379
transform 1 0 1160 0 -1 1672
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5202_6
timestamp 1731220379
transform 1 0 1256 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5201_6
timestamp 1731220379
transform 1 0 1128 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5200_6
timestamp 1731220379
transform 1 0 984 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5199_6
timestamp 1731220379
transform 1 0 840 0 1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5198_6
timestamp 1731220379
transform 1 0 1216 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5197_6
timestamp 1731220379
transform 1 0 1120 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5196_6
timestamp 1731220379
transform 1 0 1024 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5195_6
timestamp 1731220379
transform 1 0 928 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5194_6
timestamp 1731220379
transform 1 0 824 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5193_6
timestamp 1731220379
transform 1 0 712 0 -1 1788
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5192_6
timestamp 1731220379
transform 1 0 1048 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5191_6
timestamp 1731220379
transform 1 0 960 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5190_6
timestamp 1731220379
transform 1 0 872 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5189_6
timestamp 1731220379
transform 1 0 784 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5188_6
timestamp 1731220379
transform 1 0 704 0 1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5187_6
timestamp 1731220379
transform 1 0 712 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5186_6
timestamp 1731220379
transform 1 0 776 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5185_6
timestamp 1731220379
transform 1 0 840 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5184_6
timestamp 1731220379
transform 1 0 968 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5183_6
timestamp 1731220379
transform 1 0 904 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5182_6
timestamp 1731220379
transform 1 0 864 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5181_6
timestamp 1731220379
transform 1 0 936 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5180_6
timestamp 1731220379
transform 1 0 1008 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5179_6
timestamp 1731220379
transform 1 0 976 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5178_6
timestamp 1731220379
transform 1 0 880 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5177_6
timestamp 1731220379
transform 1 0 1072 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5176_6
timestamp 1731220379
transform 1 0 992 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5175_6
timestamp 1731220379
transform 1 0 912 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5174_6
timestamp 1731220379
transform 1 0 1080 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5173_6
timestamp 1731220379
transform 1 0 1168 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5172_6
timestamp 1731220379
transform 1 0 1256 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5171_6
timestamp 1731220379
transform 1 0 1152 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5170_6
timestamp 1731220379
transform 1 0 1048 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5169_6
timestamp 1731220379
transform 1 0 952 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5168_6
timestamp 1731220379
transform 1 0 984 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5167_6
timestamp 1731220379
transform 1 0 1056 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5166_6
timestamp 1731220379
transform 1 0 1128 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5165_6
timestamp 1731220379
transform 1 0 1200 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5164_6
timestamp 1731220379
transform 1 0 1256 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5163_6
timestamp 1731220379
transform 1 0 1384 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5162_6
timestamp 1731220379
transform 1 0 1480 0 -1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5161_6
timestamp 1731220379
transform 1 0 1608 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5160_6
timestamp 1731220379
transform 1 0 1552 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5159_6
timestamp 1731220379
transform 1 0 1496 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5158_6
timestamp 1731220379
transform 1 0 1440 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5157_6
timestamp 1731220379
transform 1 0 1384 0 1 2256
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5156_6
timestamp 1731220379
transform 1 0 1440 0 -1 2368
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5155_6
timestamp 1731220379
transform 1 0 1496 0 -1 2368
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5154_6
timestamp 1731220379
transform 1 0 1664 0 -1 2368
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5153_6
timestamp 1731220379
transform 1 0 1608 0 -1 2368
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5152_6
timestamp 1731220379
transform 1 0 1552 0 -1 2368
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5151_6
timestamp 1731220379
transform 1 0 1520 0 1 2372
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5150_6
timestamp 1731220379
transform 1 0 1464 0 1 2372
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5149_6
timestamp 1731220379
transform 1 0 1576 0 1 2372
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5148_6
timestamp 1731220379
transform 1 0 1632 0 1 2372
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5147_6
timestamp 1731220379
transform 1 0 1688 0 1 2372
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5146_6
timestamp 1731220379
transform 1 0 1744 0 1 2372
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5145_6
timestamp 1731220379
transform 1 0 1720 0 -1 2492
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5144_6
timestamp 1731220379
transform 1 0 1664 0 -1 2492
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5143_6
timestamp 1731220379
transform 1 0 1608 0 -1 2492
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5142_6
timestamp 1731220379
transform 1 0 1552 0 -1 2492
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5141_6
timestamp 1731220379
transform 1 0 1496 0 -1 2492
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5140_6
timestamp 1731220379
transform 1 0 1440 0 -1 2492
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5139_6
timestamp 1731220379
transform 1 0 1720 0 1 2496
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5138_6
timestamp 1731220379
transform 1 0 1664 0 1 2496
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5137_6
timestamp 1731220379
transform 1 0 1608 0 1 2496
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5136_6
timestamp 1731220379
transform 1 0 1552 0 1 2496
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5135_6
timestamp 1731220379
transform 1 0 1496 0 1 2496
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5134_6
timestamp 1731220379
transform 1 0 1440 0 1 2496
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5133_6
timestamp 1731220379
transform 1 0 1384 0 1 2496
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5132_6
timestamp 1731220379
transform 1 0 1664 0 -1 2608
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5131_6
timestamp 1731220379
transform 1 0 1608 0 -1 2608
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5130_6
timestamp 1731220379
transform 1 0 1552 0 -1 2608
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5129_6
timestamp 1731220379
transform 1 0 1496 0 -1 2608
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5128_6
timestamp 1731220379
transform 1 0 1440 0 -1 2608
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5127_6
timestamp 1731220379
transform 1 0 1384 0 -1 2608
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5126_6
timestamp 1731220379
transform 1 0 1256 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5125_6
timestamp 1731220379
transform 1 0 1200 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5124_6
timestamp 1731220379
transform 1 0 1144 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5123_6
timestamp 1731220379
transform 1 0 1080 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5122_6
timestamp 1731220379
transform 1 0 1016 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5121_6
timestamp 1731220379
transform 1 0 952 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5120_6
timestamp 1731220379
transform 1 0 888 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5119_6
timestamp 1731220379
transform 1 0 824 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5118_6
timestamp 1731220379
transform 1 0 752 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5117_6
timestamp 1731220379
transform 1 0 672 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5116_6
timestamp 1731220379
transform 1 0 592 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5115_6
timestamp 1731220379
transform 1 0 1256 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5114_6
timestamp 1731220379
transform 1 0 1176 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5113_6
timestamp 1731220379
transform 1 0 1072 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5112_6
timestamp 1731220379
transform 1 0 976 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5111_6
timestamp 1731220379
transform 1 0 872 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5110_6
timestamp 1731220379
transform 1 0 760 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5109_6
timestamp 1731220379
transform 1 0 1224 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5108_6
timestamp 1731220379
transform 1 0 1128 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5107_6
timestamp 1731220379
transform 1 0 1032 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5106_6
timestamp 1731220379
transform 1 0 936 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5105_6
timestamp 1731220379
transform 1 0 840 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5104_6
timestamp 1731220379
transform 1 0 736 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5103_6
timestamp 1731220379
transform 1 0 1112 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5102_6
timestamp 1731220379
transform 1 0 1024 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5101_6
timestamp 1731220379
transform 1 0 944 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5100_6
timestamp 1731220379
transform 1 0 864 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_599_6
timestamp 1731220379
transform 1 0 784 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_598_6
timestamp 1731220379
transform 1 0 696 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_597_6
timestamp 1731220379
transform 1 0 1000 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_596_6
timestamp 1731220379
transform 1 0 936 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_595_6
timestamp 1731220379
transform 1 0 872 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_594_6
timestamp 1731220379
transform 1 0 808 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_593_6
timestamp 1731220379
transform 1 0 744 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_592_6
timestamp 1731220379
transform 1 0 680 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_591_6
timestamp 1731220379
transform 1 0 936 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_590_6
timestamp 1731220379
transform 1 0 880 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_589_6
timestamp 1731220379
transform 1 0 824 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_588_6
timestamp 1731220379
transform 1 0 768 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_587_6
timestamp 1731220379
transform 1 0 712 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_586_6
timestamp 1731220379
transform 1 0 912 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_585_6
timestamp 1731220379
transform 1 0 840 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_584_6
timestamp 1731220379
transform 1 0 768 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_583_6
timestamp 1731220379
transform 1 0 744 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_582_6
timestamp 1731220379
transform 1 0 848 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_581_6
timestamp 1731220379
transform 1 0 832 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_580_6
timestamp 1731220379
transform 1 0 744 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_579_6
timestamp 1731220379
transform 1 0 648 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_578_6
timestamp 1731220379
transform 1 0 616 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_577_6
timestamp 1731220379
transform 1 0 704 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_576_6
timestamp 1731220379
transform 1 0 792 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_575_6
timestamp 1731220379
transform 1 0 792 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_574_6
timestamp 1731220379
transform 1 0 720 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_573_6
timestamp 1731220379
transform 1 0 656 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_572_6
timestamp 1731220379
transform 1 0 592 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_571_6
timestamp 1731220379
transform 1 0 656 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_570_6
timestamp 1731220379
transform 1 0 600 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_569_6
timestamp 1731220379
transform 1 0 544 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_568_6
timestamp 1731220379
transform 1 0 488 0 -1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_567_6
timestamp 1731220379
transform 1 0 536 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_566_6
timestamp 1731220379
transform 1 0 480 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_565_6
timestamp 1731220379
transform 1 0 424 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_564_6
timestamp 1731220379
transform 1 0 368 0 1 1912
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_563_6
timestamp 1731220379
transform 1 0 528 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_562_6
timestamp 1731220379
transform 1 0 440 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_561_6
timestamp 1731220379
transform 1 0 360 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_560_6
timestamp 1731220379
transform 1 0 280 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_559_6
timestamp 1731220379
transform 1 0 208 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_558_6
timestamp 1731220379
transform 1 0 144 0 -1 2024
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_557_6
timestamp 1731220379
transform 1 0 552 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_556_6
timestamp 1731220379
transform 1 0 448 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_555_6
timestamp 1731220379
transform 1 0 352 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_554_6
timestamp 1731220379
transform 1 0 256 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_553_6
timestamp 1731220379
transform 1 0 184 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_552_6
timestamp 1731220379
transform 1 0 128 0 1 2032
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_551_6
timestamp 1731220379
transform 1 0 168 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_550_6
timestamp 1731220379
transform 1 0 240 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_549_6
timestamp 1731220379
transform 1 0 320 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_548_6
timestamp 1731220379
transform 1 0 416 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_547_6
timestamp 1731220379
transform 1 0 520 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_546_6
timestamp 1731220379
transform 1 0 632 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_545_6
timestamp 1731220379
transform 1 0 520 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_544_6
timestamp 1731220379
transform 1 0 464 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_543_6
timestamp 1731220379
transform 1 0 408 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_542_6
timestamp 1731220379
transform 1 0 576 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_541_6
timestamp 1731220379
transform 1 0 632 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_540_6
timestamp 1731220379
transform 1 0 696 0 1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_539_6
timestamp 1731220379
transform 1 0 656 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_538_6
timestamp 1731220379
transform 1 0 600 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_537_6
timestamp 1731220379
transform 1 0 544 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_536_6
timestamp 1731220379
transform 1 0 488 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_535_6
timestamp 1731220379
transform 1 0 432 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_534_6
timestamp 1731220379
transform 1 0 376 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_533_6
timestamp 1731220379
transform 1 0 616 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_532_6
timestamp 1731220379
transform 1 0 552 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_531_6
timestamp 1731220379
transform 1 0 488 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_530_6
timestamp 1731220379
transform 1 0 424 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_529_6
timestamp 1731220379
transform 1 0 368 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_528_6
timestamp 1731220379
transform 1 0 312 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_527_6
timestamp 1731220379
transform 1 0 608 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_526_6
timestamp 1731220379
transform 1 0 512 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_525_6
timestamp 1731220379
transform 1 0 424 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_524_6
timestamp 1731220379
transform 1 0 336 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_523_6
timestamp 1731220379
transform 1 0 256 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_522_6
timestamp 1731220379
transform 1 0 192 0 -1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_521_6
timestamp 1731220379
transform 1 0 624 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_520_6
timestamp 1731220379
transform 1 0 504 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_519_6
timestamp 1731220379
transform 1 0 392 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_518_6
timestamp 1731220379
transform 1 0 280 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_517_6
timestamp 1731220379
transform 1 0 184 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_516_6
timestamp 1731220379
transform 1 0 128 0 1 2416
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_515_6
timestamp 1731220379
transform 1 0 640 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_514_6
timestamp 1731220379
transform 1 0 520 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_513_6
timestamp 1731220379
transform 1 0 400 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_512_6
timestamp 1731220379
transform 1 0 288 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_511_6
timestamp 1731220379
transform 1 0 184 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_510_6
timestamp 1731220379
transform 1 0 128 0 -1 2536
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_59_6
timestamp 1731220379
transform 1 0 504 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_58_6
timestamp 1731220379
transform 1 0 416 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_57_6
timestamp 1731220379
transform 1 0 328 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_56_6
timestamp 1731220379
transform 1 0 248 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_55_6
timestamp 1731220379
transform 1 0 184 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_54_6
timestamp 1731220379
transform 1 0 128 0 1 2548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_53_6
timestamp 1731220379
transform 1 0 296 0 -1 2660
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_52_6
timestamp 1731220379
transform 1 0 240 0 -1 2660
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_51_6
timestamp 1731220379
transform 1 0 184 0 -1 2660
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_50_6
timestamp 1731220379
transform 1 0 128 0 -1 2660
box 8 4 52 52
<< end >>
