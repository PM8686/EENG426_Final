magic
tech sky130l
timestamp 1730767165
<< m1 >>
rect 576 1387 580 1435
rect 1024 1319 1028 1351
rect 544 1255 548 1315
rect 448 195 452 219
<< m2c >>
rect 448 1503 452 1507
rect 536 1503 540 1507
rect 624 1503 628 1507
rect 720 1503 724 1507
rect 832 1503 836 1507
rect 952 1503 956 1507
rect 1080 1503 1084 1507
rect 1216 1503 1220 1507
rect 1496 1503 1500 1507
rect 111 1489 115 1493
rect 1567 1489 1571 1493
rect 111 1471 115 1475
rect 1567 1471 1571 1475
rect 576 1435 580 1439
rect 111 1425 115 1429
rect 111 1407 115 1411
rect 472 1391 476 1395
rect 1567 1425 1571 1429
rect 1567 1407 1571 1411
rect 1448 1391 1452 1395
rect 576 1383 580 1387
rect 704 1383 708 1387
rect 944 1383 948 1387
rect 1192 1383 1196 1387
rect 744 1367 748 1371
rect 1440 1367 1444 1371
rect 520 1359 524 1363
rect 968 1359 972 1363
rect 1200 1359 1204 1363
rect 1024 1351 1028 1355
rect 111 1345 115 1349
rect 111 1327 115 1331
rect 1567 1345 1571 1349
rect 1567 1327 1571 1331
rect 544 1315 548 1319
rect 1024 1315 1028 1319
rect 111 1285 115 1289
rect 111 1267 115 1271
rect 1567 1285 1571 1289
rect 1567 1267 1571 1271
rect 544 1251 548 1255
rect 568 1251 572 1255
rect 1256 1251 1260 1255
rect 792 1243 796 1247
rect 1024 1243 1028 1247
rect 1488 1243 1492 1247
rect 1016 1215 1020 1219
rect 1440 1215 1444 1219
rect 616 1207 620 1211
rect 816 1207 820 1211
rect 1224 1207 1228 1211
rect 111 1193 115 1197
rect 1567 1193 1571 1197
rect 111 1175 115 1179
rect 1567 1175 1571 1179
rect 111 1141 115 1145
rect 1567 1141 1571 1145
rect 111 1123 115 1127
rect 1567 1123 1571 1127
rect 752 1107 756 1111
rect 1456 1107 1460 1111
rect 1104 1099 1108 1103
rect 1080 1087 1084 1091
rect 1464 1087 1468 1091
rect 720 1079 724 1083
rect 896 1079 900 1083
rect 1272 1079 1276 1083
rect 111 1065 115 1069
rect 1567 1065 1571 1069
rect 111 1047 115 1051
rect 1567 1047 1571 1051
rect 111 997 115 1001
rect 1567 997 1571 1001
rect 111 979 115 983
rect 1567 979 1571 983
rect 1032 963 1036 967
rect 1456 963 1460 967
rect 624 955 628 959
rect 824 955 828 959
rect 1240 955 1244 959
rect 456 935 460 939
rect 1448 935 1452 939
rect 784 927 788 931
rect 1112 927 1116 931
rect 111 913 115 917
rect 1567 913 1571 917
rect 111 895 115 899
rect 1567 895 1571 899
rect 111 857 115 861
rect 1567 857 1571 861
rect 111 839 115 843
rect 1567 839 1571 843
rect 856 823 860 827
rect 1440 823 1444 827
rect 304 815 308 819
rect 576 815 580 819
rect 1144 815 1148 819
rect 216 783 220 787
rect 1440 783 1444 787
rect 432 775 436 779
rect 672 775 676 779
rect 920 775 924 779
rect 1176 775 1180 779
rect 111 761 115 765
rect 1567 761 1571 765
rect 111 743 115 747
rect 1567 743 1571 747
rect 111 689 115 693
rect 1567 689 1571 693
rect 360 683 364 687
rect 111 671 115 675
rect 1567 671 1571 675
rect 888 655 892 659
rect 1448 655 1452 659
rect 368 647 372 651
rect 624 647 628 651
rect 1168 647 1172 651
rect 1104 623 1108 627
rect 1456 623 1460 627
rect 632 615 636 619
rect 776 615 780 619
rect 936 615 940 619
rect 1280 615 1284 619
rect 111 601 115 605
rect 1567 601 1571 605
rect 111 583 115 587
rect 1567 583 1571 587
rect 111 529 115 533
rect 1567 529 1571 533
rect 111 511 115 515
rect 1567 511 1571 515
rect 808 495 812 499
rect 1376 495 1380 499
rect 912 487 916 491
rect 1024 487 1028 491
rect 1136 487 1140 491
rect 1256 487 1260 491
rect 1496 487 1500 491
rect 1080 463 1084 467
rect 1512 463 1516 467
rect 768 455 772 459
rect 872 455 876 459
rect 976 455 980 459
rect 1184 455 1188 459
rect 1288 455 1292 459
rect 1400 455 1404 459
rect 111 441 115 445
rect 1567 441 1571 445
rect 111 423 115 427
rect 1567 423 1571 427
rect 111 361 115 365
rect 1567 361 1571 365
rect 111 343 115 347
rect 1567 343 1571 347
rect 824 327 828 331
rect 560 319 564 323
rect 648 319 652 323
rect 736 319 740 323
rect 600 299 604 303
rect 424 291 428 295
rect 512 291 516 295
rect 111 277 115 281
rect 1567 277 1571 281
rect 111 259 115 263
rect 1567 259 1571 263
rect 111 225 115 229
rect 1567 225 1571 229
rect 288 219 292 223
rect 448 219 452 223
rect 111 207 115 211
rect 1567 207 1571 211
rect 384 191 388 195
rect 448 191 452 195
rect 472 191 476 195
rect 296 183 300 187
rect 624 143 628 147
rect 184 135 188 139
rect 272 135 276 139
rect 360 135 364 139
rect 448 135 452 139
rect 536 135 540 139
rect 111 121 115 125
rect 1567 121 1571 125
rect 111 103 115 107
rect 1567 103 1571 107
<< m2 >>
rect 398 1510 404 1511
rect 398 1506 399 1510
rect 403 1506 404 1510
rect 486 1510 492 1511
rect 398 1505 404 1506
rect 447 1507 453 1508
rect 447 1503 448 1507
rect 452 1506 453 1507
rect 486 1506 487 1510
rect 491 1506 492 1510
rect 574 1510 580 1511
rect 452 1504 482 1506
rect 486 1505 492 1506
rect 535 1507 541 1508
rect 452 1503 453 1504
rect 447 1502 453 1503
rect 480 1498 482 1504
rect 535 1503 536 1507
rect 540 1506 541 1507
rect 574 1506 575 1510
rect 579 1506 580 1510
rect 670 1510 676 1511
rect 540 1504 570 1506
rect 574 1505 580 1506
rect 623 1507 629 1508
rect 540 1503 541 1504
rect 535 1502 541 1503
rect 502 1499 508 1500
rect 502 1498 503 1499
rect 480 1496 503 1498
rect 502 1495 503 1496
rect 507 1495 508 1499
rect 568 1498 570 1504
rect 623 1503 624 1507
rect 628 1506 629 1507
rect 670 1506 671 1510
rect 675 1506 676 1510
rect 782 1510 788 1511
rect 628 1504 666 1506
rect 670 1505 676 1506
rect 719 1507 725 1508
rect 628 1503 629 1504
rect 623 1502 629 1503
rect 590 1499 596 1500
rect 590 1498 591 1499
rect 568 1496 591 1498
rect 502 1494 508 1495
rect 590 1495 591 1496
rect 595 1495 596 1499
rect 664 1498 666 1504
rect 719 1503 720 1507
rect 724 1506 725 1507
rect 782 1506 783 1510
rect 787 1506 788 1510
rect 902 1510 908 1511
rect 724 1504 762 1506
rect 782 1505 788 1506
rect 831 1507 837 1508
rect 724 1503 725 1504
rect 719 1502 725 1503
rect 686 1499 692 1500
rect 686 1498 687 1499
rect 664 1496 687 1498
rect 590 1494 596 1495
rect 686 1495 687 1496
rect 691 1495 692 1499
rect 760 1498 762 1504
rect 831 1503 832 1507
rect 836 1506 837 1507
rect 902 1506 903 1510
rect 907 1506 908 1510
rect 1030 1510 1036 1511
rect 836 1504 882 1506
rect 902 1505 908 1506
rect 951 1507 957 1508
rect 836 1503 837 1504
rect 831 1502 837 1503
rect 798 1499 804 1500
rect 798 1498 799 1499
rect 760 1496 799 1498
rect 686 1494 692 1495
rect 798 1495 799 1496
rect 803 1495 804 1499
rect 880 1498 882 1504
rect 951 1503 952 1507
rect 956 1506 957 1507
rect 1030 1506 1031 1510
rect 1035 1506 1036 1510
rect 1166 1510 1172 1511
rect 956 1504 1010 1506
rect 1030 1505 1036 1506
rect 1079 1507 1085 1508
rect 956 1503 957 1504
rect 951 1502 957 1503
rect 918 1499 924 1500
rect 918 1498 919 1499
rect 880 1496 919 1498
rect 798 1494 804 1495
rect 918 1495 919 1496
rect 923 1495 924 1499
rect 1008 1498 1010 1504
rect 1079 1503 1080 1507
rect 1084 1506 1085 1507
rect 1166 1506 1167 1510
rect 1171 1506 1172 1510
rect 1302 1510 1308 1511
rect 1084 1504 1150 1506
rect 1166 1505 1172 1506
rect 1210 1507 1221 1508
rect 1084 1503 1085 1504
rect 1079 1502 1085 1503
rect 1046 1499 1052 1500
rect 1046 1498 1047 1499
rect 1008 1496 1047 1498
rect 918 1494 924 1495
rect 1046 1495 1047 1496
rect 1051 1495 1052 1499
rect 1148 1498 1150 1504
rect 1210 1503 1211 1507
rect 1215 1503 1216 1507
rect 1220 1503 1221 1507
rect 1302 1506 1303 1510
rect 1307 1506 1308 1510
rect 1302 1505 1308 1506
rect 1446 1510 1452 1511
rect 1446 1506 1447 1510
rect 1451 1506 1452 1510
rect 1495 1507 1501 1508
rect 1495 1506 1496 1507
rect 1446 1505 1452 1506
rect 1210 1502 1221 1503
rect 1472 1504 1496 1506
rect 1182 1499 1188 1500
rect 1182 1498 1183 1499
rect 1148 1496 1183 1498
rect 1046 1494 1052 1495
rect 1182 1495 1183 1496
rect 1187 1495 1188 1499
rect 1182 1494 1188 1495
rect 1414 1499 1420 1500
rect 1414 1495 1415 1499
rect 1419 1498 1420 1499
rect 1472 1498 1474 1504
rect 1495 1503 1496 1504
rect 1500 1503 1501 1507
rect 1495 1502 1501 1503
rect 1419 1496 1474 1498
rect 1419 1495 1420 1496
rect 1414 1494 1420 1495
rect 110 1493 116 1494
rect 110 1489 111 1493
rect 115 1489 116 1493
rect 110 1488 116 1489
rect 1566 1493 1572 1494
rect 1566 1489 1567 1493
rect 1571 1489 1572 1493
rect 1566 1488 1572 1489
rect 110 1475 116 1476
rect 110 1471 111 1475
rect 115 1471 116 1475
rect 110 1470 116 1471
rect 1566 1475 1572 1476
rect 1566 1471 1567 1475
rect 1571 1471 1572 1475
rect 1566 1470 1572 1471
rect 398 1464 404 1465
rect 486 1464 492 1465
rect 574 1464 580 1465
rect 670 1464 676 1465
rect 782 1464 788 1465
rect 902 1464 908 1465
rect 1030 1464 1036 1465
rect 1166 1464 1172 1465
rect 1302 1464 1308 1465
rect 1446 1464 1452 1465
rect 398 1460 399 1464
rect 403 1460 404 1464
rect 398 1459 404 1460
rect 466 1463 472 1464
rect 466 1459 467 1463
rect 471 1459 472 1463
rect 486 1460 487 1464
rect 491 1460 492 1464
rect 486 1459 492 1460
rect 502 1463 508 1464
rect 502 1459 503 1463
rect 507 1462 508 1463
rect 507 1460 521 1462
rect 574 1460 575 1464
rect 579 1460 580 1464
rect 507 1459 508 1460
rect 574 1459 580 1460
rect 590 1463 596 1464
rect 590 1459 591 1463
rect 595 1462 596 1463
rect 595 1460 609 1462
rect 670 1460 671 1464
rect 675 1460 676 1464
rect 595 1459 596 1460
rect 670 1459 676 1460
rect 686 1463 692 1464
rect 686 1459 687 1463
rect 691 1462 692 1463
rect 691 1460 705 1462
rect 782 1460 783 1464
rect 787 1460 788 1464
rect 691 1459 692 1460
rect 782 1459 788 1460
rect 798 1463 804 1464
rect 798 1459 799 1463
rect 803 1462 804 1463
rect 803 1460 817 1462
rect 902 1460 903 1464
rect 907 1460 908 1464
rect 803 1459 804 1460
rect 902 1459 908 1460
rect 918 1463 924 1464
rect 918 1459 919 1463
rect 923 1462 924 1463
rect 923 1460 937 1462
rect 1030 1460 1031 1464
rect 1035 1460 1036 1464
rect 923 1459 924 1460
rect 1030 1459 1036 1460
rect 1046 1463 1052 1464
rect 1046 1459 1047 1463
rect 1051 1462 1052 1463
rect 1051 1460 1065 1462
rect 1166 1460 1167 1464
rect 1171 1460 1172 1464
rect 1051 1459 1052 1460
rect 1166 1459 1172 1460
rect 1182 1463 1188 1464
rect 1182 1459 1183 1463
rect 1187 1462 1188 1463
rect 1187 1460 1201 1462
rect 1302 1460 1303 1464
rect 1307 1460 1308 1464
rect 1414 1463 1420 1464
rect 1414 1462 1415 1463
rect 1373 1460 1415 1462
rect 1187 1459 1188 1460
rect 1302 1459 1308 1460
rect 1414 1459 1415 1460
rect 1419 1459 1420 1463
rect 1446 1460 1447 1464
rect 1451 1460 1452 1464
rect 1446 1459 1452 1460
rect 1478 1463 1484 1464
rect 1478 1459 1479 1463
rect 1483 1459 1484 1463
rect 466 1458 472 1459
rect 502 1458 508 1459
rect 590 1458 596 1459
rect 686 1458 692 1459
rect 798 1458 804 1459
rect 918 1458 924 1459
rect 1046 1458 1052 1459
rect 1182 1458 1188 1459
rect 1414 1458 1420 1459
rect 1478 1458 1484 1459
rect 422 1440 428 1441
rect 654 1440 660 1441
rect 894 1440 900 1441
rect 1142 1440 1148 1441
rect 1398 1440 1404 1441
rect 422 1436 423 1440
rect 427 1436 428 1440
rect 575 1439 581 1440
rect 575 1438 576 1439
rect 493 1436 576 1438
rect 422 1435 428 1436
rect 575 1435 576 1436
rect 580 1435 581 1439
rect 654 1436 655 1440
rect 659 1436 660 1440
rect 654 1435 660 1436
rect 722 1439 728 1440
rect 722 1435 723 1439
rect 727 1435 728 1439
rect 894 1436 895 1440
rect 899 1436 900 1440
rect 894 1435 900 1436
rect 910 1439 916 1440
rect 910 1435 911 1439
rect 915 1438 916 1439
rect 915 1436 929 1438
rect 1142 1436 1143 1440
rect 1147 1436 1148 1440
rect 915 1435 916 1436
rect 1142 1435 1148 1436
rect 1210 1439 1216 1440
rect 1210 1435 1211 1439
rect 1215 1435 1216 1439
rect 1398 1436 1399 1440
rect 1403 1436 1404 1440
rect 1398 1435 1404 1436
rect 1438 1439 1444 1440
rect 1438 1435 1439 1439
rect 1443 1435 1444 1439
rect 575 1434 581 1435
rect 722 1434 728 1435
rect 910 1434 916 1435
rect 1210 1434 1216 1435
rect 1438 1434 1444 1435
rect 110 1429 116 1430
rect 110 1425 111 1429
rect 115 1425 116 1429
rect 110 1424 116 1425
rect 1566 1429 1572 1430
rect 1566 1425 1567 1429
rect 1571 1425 1572 1429
rect 1566 1424 1572 1425
rect 110 1411 116 1412
rect 110 1407 111 1411
rect 115 1407 116 1411
rect 110 1406 116 1407
rect 1566 1411 1572 1412
rect 1566 1407 1567 1411
rect 1571 1407 1572 1411
rect 1566 1406 1572 1407
rect 466 1395 477 1396
rect 1447 1395 1453 1396
rect 422 1394 428 1395
rect 422 1390 423 1394
rect 427 1390 428 1394
rect 466 1391 467 1395
rect 471 1391 472 1395
rect 476 1391 477 1395
rect 466 1390 477 1391
rect 654 1394 660 1395
rect 654 1390 655 1394
rect 659 1390 660 1394
rect 422 1389 428 1390
rect 654 1389 660 1390
rect 894 1394 900 1395
rect 894 1390 895 1394
rect 899 1390 900 1394
rect 894 1389 900 1390
rect 1142 1394 1148 1395
rect 1142 1390 1143 1394
rect 1147 1390 1148 1394
rect 1142 1389 1148 1390
rect 1398 1394 1404 1395
rect 1398 1390 1399 1394
rect 1403 1390 1404 1394
rect 1447 1391 1448 1395
rect 1452 1394 1453 1395
rect 1478 1395 1484 1396
rect 1478 1394 1479 1395
rect 1452 1392 1479 1394
rect 1452 1391 1453 1392
rect 1447 1390 1453 1391
rect 1478 1391 1479 1392
rect 1483 1391 1484 1395
rect 1478 1390 1484 1391
rect 1398 1389 1404 1390
rect 575 1387 581 1388
rect 575 1383 576 1387
rect 580 1386 581 1387
rect 703 1387 709 1388
rect 703 1386 704 1387
rect 580 1384 704 1386
rect 580 1383 581 1384
rect 575 1382 581 1383
rect 703 1383 704 1384
rect 708 1383 709 1387
rect 703 1382 709 1383
rect 722 1387 728 1388
rect 722 1383 723 1387
rect 727 1386 728 1387
rect 943 1387 949 1388
rect 943 1386 944 1387
rect 727 1384 944 1386
rect 727 1383 728 1384
rect 722 1382 728 1383
rect 943 1383 944 1384
rect 948 1383 949 1387
rect 943 1382 949 1383
rect 1190 1387 1197 1388
rect 1190 1383 1191 1387
rect 1196 1383 1197 1387
rect 1190 1382 1197 1383
rect 743 1371 749 1372
rect 743 1367 744 1371
rect 748 1370 749 1371
rect 910 1371 916 1372
rect 910 1370 911 1371
rect 748 1368 911 1370
rect 748 1367 749 1368
rect 470 1366 476 1367
rect 470 1362 471 1366
rect 475 1362 476 1366
rect 694 1366 700 1367
rect 743 1366 749 1367
rect 910 1367 911 1368
rect 915 1367 916 1371
rect 1438 1371 1445 1372
rect 1438 1367 1439 1371
rect 1444 1367 1445 1371
rect 910 1366 916 1367
rect 918 1366 924 1367
rect 470 1361 476 1362
rect 519 1363 525 1364
rect 519 1359 520 1363
rect 524 1362 525 1363
rect 694 1362 695 1366
rect 699 1362 700 1366
rect 524 1360 626 1362
rect 694 1361 700 1362
rect 918 1362 919 1366
rect 923 1362 924 1366
rect 1150 1366 1156 1367
rect 918 1361 924 1362
rect 967 1363 973 1364
rect 524 1359 525 1360
rect 519 1358 525 1359
rect 624 1354 626 1360
rect 967 1359 968 1363
rect 972 1362 973 1363
rect 1006 1363 1012 1364
rect 1006 1362 1007 1363
rect 972 1360 1007 1362
rect 972 1359 973 1360
rect 967 1358 973 1359
rect 1006 1359 1007 1360
rect 1011 1359 1012 1363
rect 1150 1362 1151 1366
rect 1155 1362 1156 1366
rect 1390 1366 1396 1367
rect 1438 1366 1445 1367
rect 1199 1363 1205 1364
rect 1199 1362 1200 1363
rect 1150 1361 1156 1362
rect 1006 1358 1012 1359
rect 1176 1360 1200 1362
rect 710 1355 716 1356
rect 710 1354 711 1355
rect 624 1352 711 1354
rect 710 1351 711 1352
rect 715 1351 716 1355
rect 710 1350 716 1351
rect 1023 1355 1029 1356
rect 1023 1351 1024 1355
rect 1028 1354 1029 1355
rect 1176 1354 1178 1360
rect 1199 1359 1200 1360
rect 1204 1359 1205 1363
rect 1390 1362 1391 1366
rect 1395 1362 1396 1366
rect 1390 1361 1396 1362
rect 1199 1358 1205 1359
rect 1028 1352 1178 1354
rect 1028 1351 1029 1352
rect 1023 1350 1029 1351
rect 110 1349 116 1350
rect 110 1345 111 1349
rect 115 1345 116 1349
rect 110 1344 116 1345
rect 1566 1349 1572 1350
rect 1566 1345 1567 1349
rect 1571 1345 1572 1349
rect 1566 1344 1572 1345
rect 110 1331 116 1332
rect 110 1327 111 1331
rect 115 1327 116 1331
rect 110 1326 116 1327
rect 1566 1331 1572 1332
rect 1566 1327 1567 1331
rect 1571 1327 1572 1331
rect 1566 1326 1572 1327
rect 470 1320 476 1321
rect 694 1320 700 1321
rect 918 1320 924 1321
rect 1150 1320 1156 1321
rect 1390 1320 1396 1321
rect 470 1316 471 1320
rect 475 1316 476 1320
rect 543 1319 549 1320
rect 543 1318 544 1319
rect 541 1316 544 1318
rect 470 1315 476 1316
rect 543 1315 544 1316
rect 548 1315 549 1319
rect 694 1316 695 1320
rect 699 1316 700 1320
rect 694 1315 700 1316
rect 710 1319 716 1320
rect 710 1315 711 1319
rect 715 1318 716 1319
rect 715 1316 729 1318
rect 918 1316 919 1320
rect 923 1316 924 1320
rect 1023 1319 1029 1320
rect 1023 1318 1024 1319
rect 989 1316 1024 1318
rect 715 1315 716 1316
rect 918 1315 924 1316
rect 1023 1315 1024 1316
rect 1028 1315 1029 1319
rect 1150 1316 1151 1320
rect 1155 1316 1156 1320
rect 1150 1315 1156 1316
rect 1190 1319 1196 1320
rect 1190 1315 1191 1319
rect 1195 1315 1196 1319
rect 1390 1316 1391 1320
rect 1395 1316 1396 1320
rect 1390 1315 1396 1316
rect 1422 1319 1428 1320
rect 1422 1315 1423 1319
rect 1427 1315 1428 1319
rect 543 1314 549 1315
rect 710 1314 716 1315
rect 1023 1314 1029 1315
rect 1190 1314 1196 1315
rect 1422 1314 1428 1315
rect 518 1300 524 1301
rect 742 1300 748 1301
rect 974 1300 980 1301
rect 1206 1300 1212 1301
rect 1438 1300 1444 1301
rect 518 1296 519 1300
rect 523 1296 524 1300
rect 518 1295 524 1296
rect 586 1299 592 1300
rect 586 1295 587 1299
rect 591 1295 592 1299
rect 742 1296 743 1300
rect 747 1296 748 1300
rect 742 1295 748 1296
rect 810 1299 816 1300
rect 810 1295 811 1299
rect 815 1295 816 1299
rect 974 1296 975 1300
rect 979 1296 980 1300
rect 974 1295 980 1296
rect 1006 1299 1012 1300
rect 1006 1295 1007 1299
rect 1011 1295 1012 1299
rect 1206 1296 1207 1300
rect 1211 1296 1212 1300
rect 1206 1295 1212 1296
rect 1274 1299 1280 1300
rect 1274 1295 1275 1299
rect 1279 1295 1280 1299
rect 1438 1296 1439 1300
rect 1443 1296 1444 1300
rect 1438 1295 1444 1296
rect 1470 1299 1476 1300
rect 1470 1295 1471 1299
rect 1475 1295 1476 1299
rect 586 1294 592 1295
rect 810 1294 816 1295
rect 1006 1294 1012 1295
rect 1274 1294 1280 1295
rect 1470 1294 1476 1295
rect 110 1289 116 1290
rect 110 1285 111 1289
rect 115 1285 116 1289
rect 110 1284 116 1285
rect 1566 1289 1572 1290
rect 1566 1285 1567 1289
rect 1571 1285 1572 1289
rect 1566 1284 1572 1285
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 110 1266 116 1267
rect 1566 1271 1572 1272
rect 1566 1267 1567 1271
rect 1571 1267 1572 1271
rect 1566 1266 1572 1267
rect 543 1255 549 1256
rect 518 1254 524 1255
rect 518 1250 519 1254
rect 523 1250 524 1254
rect 543 1251 544 1255
rect 548 1254 549 1255
rect 567 1255 573 1256
rect 1255 1255 1261 1256
rect 567 1254 568 1255
rect 548 1252 568 1254
rect 548 1251 549 1252
rect 543 1250 549 1251
rect 567 1251 568 1252
rect 572 1251 573 1255
rect 567 1250 573 1251
rect 742 1254 748 1255
rect 742 1250 743 1254
rect 747 1250 748 1254
rect 518 1249 524 1250
rect 742 1249 748 1250
rect 974 1254 980 1255
rect 974 1250 975 1254
rect 979 1250 980 1254
rect 974 1249 980 1250
rect 1206 1254 1212 1255
rect 1206 1250 1207 1254
rect 1211 1250 1212 1254
rect 1255 1251 1256 1255
rect 1260 1254 1261 1255
rect 1422 1255 1428 1256
rect 1422 1254 1423 1255
rect 1260 1252 1423 1254
rect 1260 1251 1261 1252
rect 1255 1250 1261 1251
rect 1422 1251 1423 1252
rect 1427 1251 1428 1255
rect 1422 1250 1428 1251
rect 1438 1254 1444 1255
rect 1438 1250 1439 1254
rect 1443 1250 1444 1254
rect 1206 1249 1212 1250
rect 1438 1249 1444 1250
rect 586 1247 592 1248
rect 586 1243 587 1247
rect 591 1246 592 1247
rect 791 1247 797 1248
rect 791 1246 792 1247
rect 591 1244 792 1246
rect 591 1243 592 1244
rect 586 1242 592 1243
rect 791 1243 792 1244
rect 796 1243 797 1247
rect 791 1242 797 1243
rect 1023 1247 1029 1248
rect 1023 1243 1024 1247
rect 1028 1246 1029 1247
rect 1190 1247 1196 1248
rect 1190 1246 1191 1247
rect 1028 1244 1191 1246
rect 1028 1243 1029 1244
rect 1023 1242 1029 1243
rect 1190 1243 1191 1244
rect 1195 1243 1196 1247
rect 1190 1242 1196 1243
rect 1274 1247 1280 1248
rect 1274 1243 1275 1247
rect 1279 1246 1280 1247
rect 1487 1247 1493 1248
rect 1487 1246 1488 1247
rect 1279 1244 1488 1246
rect 1279 1243 1280 1244
rect 1274 1242 1280 1243
rect 1487 1243 1488 1244
rect 1492 1243 1493 1247
rect 1487 1242 1493 1243
rect 810 1223 816 1224
rect 810 1219 811 1223
rect 815 1222 816 1223
rect 815 1220 978 1222
rect 815 1219 816 1220
rect 810 1218 816 1219
rect 976 1218 978 1220
rect 1015 1219 1021 1220
rect 1015 1218 1016 1219
rect 976 1216 1016 1218
rect 1015 1215 1016 1216
rect 1020 1215 1021 1219
rect 1439 1219 1445 1220
rect 1439 1215 1440 1219
rect 1444 1218 1445 1219
rect 1470 1219 1476 1220
rect 1470 1218 1471 1219
rect 1444 1216 1471 1218
rect 1444 1215 1445 1216
rect 566 1214 572 1215
rect 566 1210 567 1214
rect 571 1210 572 1214
rect 766 1214 772 1215
rect 566 1209 572 1210
rect 615 1211 621 1212
rect 615 1207 616 1211
rect 620 1210 621 1211
rect 766 1210 767 1214
rect 771 1210 772 1214
rect 966 1214 972 1215
rect 1015 1214 1021 1215
rect 1174 1214 1180 1215
rect 620 1208 710 1210
rect 766 1209 772 1210
rect 815 1211 821 1212
rect 620 1207 621 1208
rect 615 1206 621 1207
rect 708 1202 710 1208
rect 815 1207 816 1211
rect 820 1210 821 1211
rect 966 1210 967 1214
rect 971 1210 972 1214
rect 820 1208 910 1210
rect 966 1209 972 1210
rect 1174 1210 1175 1214
rect 1179 1210 1180 1214
rect 1390 1214 1396 1215
rect 1439 1214 1445 1215
rect 1470 1215 1471 1216
rect 1475 1215 1476 1219
rect 1470 1214 1476 1215
rect 1174 1209 1180 1210
rect 1223 1211 1229 1212
rect 820 1207 821 1208
rect 815 1206 821 1207
rect 782 1203 788 1204
rect 782 1202 783 1203
rect 708 1200 783 1202
rect 782 1199 783 1200
rect 787 1199 788 1203
rect 908 1202 910 1208
rect 1223 1207 1224 1211
rect 1228 1210 1229 1211
rect 1254 1211 1260 1212
rect 1254 1210 1255 1211
rect 1228 1208 1255 1210
rect 1228 1207 1229 1208
rect 1223 1206 1229 1207
rect 1254 1207 1255 1208
rect 1259 1207 1260 1211
rect 1390 1210 1391 1214
rect 1395 1210 1396 1214
rect 1390 1209 1396 1210
rect 1254 1206 1260 1207
rect 982 1203 988 1204
rect 982 1202 983 1203
rect 908 1200 983 1202
rect 782 1198 788 1199
rect 982 1199 983 1200
rect 987 1199 988 1203
rect 982 1198 988 1199
rect 110 1197 116 1198
rect 110 1193 111 1197
rect 115 1193 116 1197
rect 110 1192 116 1193
rect 1566 1197 1572 1198
rect 1566 1193 1567 1197
rect 1571 1193 1572 1197
rect 1566 1192 1572 1193
rect 110 1179 116 1180
rect 110 1175 111 1179
rect 115 1175 116 1179
rect 110 1174 116 1175
rect 1566 1179 1572 1180
rect 1566 1175 1567 1179
rect 1571 1175 1572 1179
rect 1566 1174 1572 1175
rect 566 1168 572 1169
rect 766 1168 772 1169
rect 966 1168 972 1169
rect 1174 1168 1180 1169
rect 1390 1168 1396 1169
rect 566 1164 567 1168
rect 571 1164 572 1168
rect 726 1167 732 1168
rect 726 1166 727 1167
rect 637 1164 727 1166
rect 566 1163 572 1164
rect 726 1163 727 1164
rect 731 1163 732 1167
rect 766 1164 767 1168
rect 771 1164 772 1168
rect 766 1163 772 1164
rect 782 1167 788 1168
rect 782 1163 783 1167
rect 787 1166 788 1167
rect 787 1164 801 1166
rect 966 1164 967 1168
rect 971 1164 972 1168
rect 787 1163 788 1164
rect 966 1163 972 1164
rect 982 1167 988 1168
rect 982 1163 983 1167
rect 987 1166 988 1167
rect 987 1164 1001 1166
rect 1174 1164 1175 1168
rect 1179 1164 1180 1168
rect 987 1163 988 1164
rect 1174 1163 1180 1164
rect 1190 1167 1196 1168
rect 1190 1163 1191 1167
rect 1195 1166 1196 1167
rect 1195 1164 1209 1166
rect 1390 1164 1391 1168
rect 1395 1164 1396 1168
rect 1195 1163 1196 1164
rect 1390 1163 1396 1164
rect 1454 1167 1460 1168
rect 1454 1163 1455 1167
rect 1459 1163 1460 1167
rect 726 1162 732 1163
rect 782 1162 788 1163
rect 982 1162 988 1163
rect 1190 1162 1196 1163
rect 1454 1162 1460 1163
rect 702 1156 708 1157
rect 1054 1156 1060 1157
rect 1406 1156 1412 1157
rect 702 1152 703 1156
rect 707 1152 708 1156
rect 978 1155 984 1156
rect 978 1154 979 1155
rect 773 1152 979 1154
rect 702 1151 708 1152
rect 978 1151 979 1152
rect 983 1151 984 1155
rect 1054 1152 1055 1156
rect 1059 1152 1060 1156
rect 1054 1151 1060 1152
rect 1078 1155 1084 1156
rect 1078 1151 1079 1155
rect 1083 1154 1084 1155
rect 1083 1152 1089 1154
rect 1406 1152 1407 1156
rect 1411 1152 1412 1156
rect 1083 1151 1084 1152
rect 1406 1151 1412 1152
rect 1462 1155 1468 1156
rect 1462 1151 1463 1155
rect 1467 1151 1468 1155
rect 978 1150 984 1151
rect 1078 1150 1084 1151
rect 1462 1150 1468 1151
rect 110 1145 116 1146
rect 110 1141 111 1145
rect 115 1141 116 1145
rect 110 1140 116 1141
rect 1566 1145 1572 1146
rect 1566 1141 1567 1145
rect 1571 1141 1572 1145
rect 1566 1140 1572 1141
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 110 1122 116 1123
rect 1566 1127 1572 1128
rect 1566 1123 1567 1127
rect 1571 1123 1572 1127
rect 1566 1122 1572 1123
rect 726 1111 732 1112
rect 702 1110 708 1111
rect 702 1106 703 1110
rect 707 1106 708 1110
rect 726 1107 727 1111
rect 731 1110 732 1111
rect 751 1111 757 1112
rect 1454 1111 1461 1112
rect 751 1110 752 1111
rect 731 1108 752 1110
rect 731 1107 732 1108
rect 726 1106 732 1107
rect 751 1107 752 1108
rect 756 1107 757 1111
rect 751 1106 757 1107
rect 1054 1110 1060 1111
rect 1054 1106 1055 1110
rect 1059 1106 1060 1110
rect 702 1105 708 1106
rect 1054 1105 1060 1106
rect 1406 1110 1412 1111
rect 1406 1106 1407 1110
rect 1411 1106 1412 1110
rect 1454 1107 1455 1111
rect 1460 1107 1461 1111
rect 1454 1106 1461 1107
rect 1406 1105 1412 1106
rect 978 1103 984 1104
rect 978 1099 979 1103
rect 983 1102 984 1103
rect 1103 1103 1109 1104
rect 1103 1102 1104 1103
rect 983 1100 1104 1102
rect 983 1099 984 1100
rect 978 1098 984 1099
rect 1103 1099 1104 1100
rect 1108 1099 1109 1103
rect 1103 1098 1109 1099
rect 1078 1091 1085 1092
rect 1078 1087 1079 1091
rect 1084 1087 1085 1091
rect 1462 1091 1469 1092
rect 1462 1087 1463 1091
rect 1468 1087 1469 1091
rect 670 1086 676 1087
rect 670 1082 671 1086
rect 675 1082 676 1086
rect 846 1086 852 1087
rect 670 1081 676 1082
rect 719 1083 725 1084
rect 719 1079 720 1083
rect 724 1082 725 1083
rect 846 1082 847 1086
rect 851 1082 852 1086
rect 1030 1086 1036 1087
rect 1078 1086 1085 1087
rect 1222 1086 1228 1087
rect 724 1080 802 1082
rect 846 1081 852 1082
rect 895 1083 901 1084
rect 724 1079 725 1080
rect 719 1078 725 1079
rect 800 1074 802 1080
rect 895 1079 896 1083
rect 900 1082 901 1083
rect 1030 1082 1031 1086
rect 1035 1082 1036 1086
rect 900 1080 982 1082
rect 1030 1081 1036 1082
rect 1222 1082 1223 1086
rect 1227 1082 1228 1086
rect 1414 1086 1420 1087
rect 1462 1086 1469 1087
rect 1222 1081 1228 1082
rect 1266 1083 1277 1084
rect 900 1079 901 1080
rect 895 1078 901 1079
rect 862 1075 868 1076
rect 862 1074 863 1075
rect 800 1072 863 1074
rect 862 1071 863 1072
rect 867 1071 868 1075
rect 980 1074 982 1080
rect 1266 1079 1267 1083
rect 1271 1079 1272 1083
rect 1276 1079 1277 1083
rect 1414 1082 1415 1086
rect 1419 1082 1420 1086
rect 1414 1081 1420 1082
rect 1266 1078 1277 1079
rect 1046 1075 1052 1076
rect 1046 1074 1047 1075
rect 980 1072 1047 1074
rect 862 1070 868 1071
rect 1046 1071 1047 1072
rect 1051 1071 1052 1075
rect 1046 1070 1052 1071
rect 110 1069 116 1070
rect 110 1065 111 1069
rect 115 1065 116 1069
rect 110 1064 116 1065
rect 1566 1069 1572 1070
rect 1566 1065 1567 1069
rect 1571 1065 1572 1069
rect 1566 1064 1572 1065
rect 110 1051 116 1052
rect 110 1047 111 1051
rect 115 1047 116 1051
rect 110 1046 116 1047
rect 1566 1051 1572 1052
rect 1566 1047 1567 1051
rect 1571 1047 1572 1051
rect 1566 1046 1572 1047
rect 670 1040 676 1041
rect 670 1036 671 1040
rect 675 1036 676 1040
rect 846 1040 852 1041
rect 1030 1040 1036 1041
rect 1222 1040 1228 1041
rect 1414 1040 1420 1041
rect 741 1036 778 1038
rect 670 1035 676 1036
rect 776 1030 778 1036
rect 846 1036 847 1040
rect 851 1036 852 1040
rect 846 1035 852 1036
rect 862 1039 868 1040
rect 862 1035 863 1039
rect 867 1038 868 1039
rect 867 1036 881 1038
rect 1030 1036 1031 1040
rect 1035 1036 1036 1040
rect 867 1035 868 1036
rect 1030 1035 1036 1036
rect 1046 1039 1052 1040
rect 1046 1035 1047 1039
rect 1051 1038 1052 1039
rect 1051 1036 1065 1038
rect 1222 1036 1223 1040
rect 1227 1036 1228 1040
rect 1051 1035 1052 1036
rect 1222 1035 1228 1036
rect 1254 1039 1260 1040
rect 1254 1035 1255 1039
rect 1259 1035 1260 1039
rect 1414 1036 1415 1040
rect 1419 1036 1420 1040
rect 1414 1035 1420 1036
rect 1454 1039 1460 1040
rect 1454 1035 1455 1039
rect 1459 1035 1460 1039
rect 862 1034 868 1035
rect 1046 1034 1052 1035
rect 1254 1034 1260 1035
rect 1454 1034 1460 1035
rect 1006 1031 1012 1032
rect 1006 1030 1007 1031
rect 776 1028 1007 1030
rect 1006 1027 1007 1028
rect 1011 1027 1012 1031
rect 1006 1026 1012 1027
rect 574 1012 580 1013
rect 774 1012 780 1013
rect 982 1012 988 1013
rect 1190 1012 1196 1013
rect 1406 1012 1412 1013
rect 574 1008 575 1012
rect 579 1008 580 1012
rect 574 1007 580 1008
rect 606 1011 612 1012
rect 606 1007 607 1011
rect 611 1007 612 1011
rect 774 1008 775 1012
rect 779 1008 780 1012
rect 774 1007 780 1008
rect 806 1011 812 1012
rect 806 1007 807 1011
rect 811 1007 812 1011
rect 982 1008 983 1012
rect 987 1008 988 1012
rect 982 1007 988 1008
rect 1014 1011 1020 1012
rect 1014 1007 1015 1011
rect 1019 1007 1020 1011
rect 1190 1008 1191 1012
rect 1195 1008 1196 1012
rect 1266 1011 1272 1012
rect 1266 1010 1267 1011
rect 1261 1008 1267 1010
rect 1190 1007 1196 1008
rect 1266 1007 1267 1008
rect 1271 1007 1272 1011
rect 1406 1008 1407 1012
rect 1411 1008 1412 1012
rect 1406 1007 1412 1008
rect 1446 1011 1452 1012
rect 1446 1007 1447 1011
rect 1451 1007 1452 1011
rect 606 1006 612 1007
rect 806 1006 812 1007
rect 1014 1006 1020 1007
rect 1266 1006 1272 1007
rect 1446 1006 1452 1007
rect 110 1001 116 1002
rect 110 997 111 1001
rect 115 997 116 1001
rect 110 996 116 997
rect 1566 1001 1572 1002
rect 1566 997 1567 1001
rect 1571 997 1572 1001
rect 1566 996 1572 997
rect 110 983 116 984
rect 110 979 111 983
rect 115 979 116 983
rect 110 978 116 979
rect 1566 983 1572 984
rect 1566 979 1567 983
rect 1571 979 1572 983
rect 1566 978 1572 979
rect 1006 967 1012 968
rect 574 966 580 967
rect 574 962 575 966
rect 579 962 580 966
rect 574 961 580 962
rect 774 966 780 967
rect 774 962 775 966
rect 779 962 780 966
rect 774 961 780 962
rect 982 966 988 967
rect 982 962 983 966
rect 987 962 988 966
rect 1006 963 1007 967
rect 1011 966 1012 967
rect 1031 967 1037 968
rect 1454 967 1461 968
rect 1031 966 1032 967
rect 1011 964 1032 966
rect 1011 963 1012 964
rect 1006 962 1012 963
rect 1031 963 1032 964
rect 1036 963 1037 967
rect 1031 962 1037 963
rect 1190 966 1196 967
rect 1190 962 1191 966
rect 1195 962 1196 966
rect 982 961 988 962
rect 1190 961 1196 962
rect 1406 966 1412 967
rect 1406 962 1407 966
rect 1411 962 1412 966
rect 1454 963 1455 967
rect 1460 963 1461 967
rect 1454 962 1461 963
rect 1406 961 1412 962
rect 623 959 629 960
rect 623 955 624 959
rect 628 958 629 959
rect 806 959 812 960
rect 806 958 807 959
rect 628 956 807 958
rect 628 955 629 956
rect 623 954 629 955
rect 806 955 807 956
rect 811 955 812 959
rect 806 954 812 955
rect 823 959 829 960
rect 823 955 824 959
rect 828 958 829 959
rect 1014 959 1020 960
rect 1014 958 1015 959
rect 828 956 1015 958
rect 828 955 829 956
rect 823 954 829 955
rect 1014 955 1015 956
rect 1019 955 1020 959
rect 1014 954 1020 955
rect 1162 959 1168 960
rect 1162 955 1163 959
rect 1167 958 1168 959
rect 1239 959 1245 960
rect 1239 958 1240 959
rect 1167 956 1240 958
rect 1167 955 1168 956
rect 1162 954 1168 955
rect 1239 955 1240 956
rect 1244 955 1245 959
rect 1239 954 1245 955
rect 455 939 461 940
rect 455 935 456 939
rect 460 938 461 939
rect 606 939 612 940
rect 606 938 607 939
rect 460 936 607 938
rect 460 935 461 936
rect 406 934 412 935
rect 455 934 461 935
rect 606 935 607 936
rect 611 935 612 939
rect 1446 939 1453 940
rect 1446 935 1447 939
rect 1452 935 1453 939
rect 606 934 612 935
rect 734 934 740 935
rect 406 930 407 934
rect 411 930 412 934
rect 406 929 412 930
rect 734 930 735 934
rect 739 930 740 934
rect 1062 934 1068 935
rect 783 931 789 932
rect 783 930 784 931
rect 734 929 740 930
rect 760 928 784 930
rect 610 923 616 924
rect 610 919 611 923
rect 615 922 616 923
rect 760 922 762 928
rect 783 927 784 928
rect 788 927 789 931
rect 1062 930 1063 934
rect 1067 930 1068 934
rect 1398 934 1404 935
rect 1446 934 1453 935
rect 1111 931 1117 932
rect 1111 930 1112 931
rect 1062 929 1068 930
rect 783 926 789 927
rect 1088 928 1112 930
rect 615 920 762 922
rect 930 923 936 924
rect 615 919 616 920
rect 610 918 616 919
rect 930 919 931 923
rect 935 922 936 923
rect 1088 922 1090 928
rect 1111 927 1112 928
rect 1116 927 1117 931
rect 1398 930 1399 934
rect 1403 930 1404 934
rect 1398 929 1404 930
rect 1111 926 1117 927
rect 935 920 1090 922
rect 935 919 936 920
rect 930 918 936 919
rect 110 917 116 918
rect 110 913 111 917
rect 115 913 116 917
rect 110 912 116 913
rect 1566 917 1572 918
rect 1566 913 1567 917
rect 1571 913 1572 917
rect 1566 912 1572 913
rect 110 899 116 900
rect 110 895 111 899
rect 115 895 116 899
rect 110 894 116 895
rect 1566 899 1572 900
rect 1566 895 1567 899
rect 1571 895 1572 899
rect 1566 894 1572 895
rect 406 888 412 889
rect 734 888 740 889
rect 1062 888 1068 889
rect 1398 888 1404 889
rect 406 884 407 888
rect 411 884 412 888
rect 610 887 616 888
rect 610 886 611 887
rect 477 884 611 886
rect 406 883 412 884
rect 610 883 611 884
rect 615 883 616 887
rect 734 884 735 888
rect 739 884 740 888
rect 930 887 936 888
rect 930 886 931 887
rect 805 884 931 886
rect 734 883 740 884
rect 930 883 931 884
rect 935 883 936 887
rect 1062 884 1063 888
rect 1067 884 1068 888
rect 1062 883 1068 884
rect 1078 887 1084 888
rect 1078 883 1079 887
rect 1083 886 1084 887
rect 1083 884 1097 886
rect 1398 884 1399 888
rect 1403 884 1404 888
rect 1083 883 1084 884
rect 1398 883 1404 884
rect 1438 887 1444 888
rect 1438 883 1439 887
rect 1443 883 1444 887
rect 610 882 616 883
rect 930 882 936 883
rect 1078 882 1084 883
rect 1438 882 1444 883
rect 254 872 260 873
rect 526 872 532 873
rect 806 872 812 873
rect 1094 872 1100 873
rect 1390 872 1396 873
rect 254 868 255 872
rect 259 868 260 872
rect 254 867 260 868
rect 286 871 292 872
rect 286 867 287 871
rect 291 867 292 871
rect 526 868 527 872
rect 531 868 532 872
rect 526 867 532 868
rect 558 871 564 872
rect 558 867 559 871
rect 563 867 564 871
rect 806 868 807 872
rect 811 868 812 872
rect 806 867 812 868
rect 838 871 844 872
rect 838 867 839 871
rect 843 867 844 871
rect 1094 868 1095 872
rect 1099 868 1100 872
rect 1094 867 1100 868
rect 1162 871 1168 872
rect 1162 867 1163 871
rect 1167 867 1168 871
rect 1390 868 1391 872
rect 1395 868 1396 872
rect 1390 867 1396 868
rect 1430 871 1436 872
rect 1430 867 1431 871
rect 1435 867 1436 871
rect 286 866 292 867
rect 558 866 564 867
rect 838 866 844 867
rect 1162 866 1168 867
rect 1430 866 1436 867
rect 110 861 116 862
rect 110 857 111 861
rect 115 857 116 861
rect 110 856 116 857
rect 1566 861 1572 862
rect 1566 857 1567 861
rect 1571 857 1572 861
rect 1566 856 1572 857
rect 110 843 116 844
rect 110 839 111 843
rect 115 839 116 843
rect 110 838 116 839
rect 1566 843 1572 844
rect 1566 839 1567 843
rect 1571 839 1572 843
rect 1566 838 1572 839
rect 855 827 861 828
rect 254 826 260 827
rect 254 822 255 826
rect 259 822 260 826
rect 254 821 260 822
rect 526 826 532 827
rect 526 822 527 826
rect 531 822 532 826
rect 526 821 532 822
rect 806 826 812 827
rect 806 822 807 826
rect 811 822 812 826
rect 855 823 856 827
rect 860 826 861 827
rect 1078 827 1084 828
rect 1438 827 1445 828
rect 1078 826 1079 827
rect 860 824 1079 826
rect 860 823 861 824
rect 855 822 861 823
rect 1078 823 1079 824
rect 1083 823 1084 827
rect 1078 822 1084 823
rect 1094 826 1100 827
rect 1094 822 1095 826
rect 1099 822 1100 826
rect 806 821 812 822
rect 1094 821 1100 822
rect 1390 826 1396 827
rect 1390 822 1391 826
rect 1395 822 1396 826
rect 1438 823 1439 827
rect 1444 823 1445 827
rect 1438 822 1445 823
rect 1390 821 1396 822
rect 303 819 309 820
rect 303 815 304 819
rect 308 818 309 819
rect 558 819 564 820
rect 558 818 559 819
rect 308 816 559 818
rect 308 815 309 816
rect 303 814 309 815
rect 558 815 559 816
rect 563 815 564 819
rect 558 814 564 815
rect 575 819 581 820
rect 575 815 576 819
rect 580 818 581 819
rect 838 819 844 820
rect 838 818 839 819
rect 580 816 839 818
rect 580 815 581 816
rect 575 814 581 815
rect 838 815 839 816
rect 843 815 844 819
rect 838 814 844 815
rect 1143 819 1149 820
rect 1143 815 1144 819
rect 1148 818 1149 819
rect 1158 819 1164 820
rect 1158 818 1159 819
rect 1148 816 1159 818
rect 1148 815 1149 816
rect 1143 814 1149 815
rect 1158 815 1159 816
rect 1163 815 1164 819
rect 1158 814 1164 815
rect 215 787 221 788
rect 215 783 216 787
rect 220 786 221 787
rect 286 787 292 788
rect 286 786 287 787
rect 220 784 287 786
rect 220 783 221 784
rect 166 782 172 783
rect 215 782 221 783
rect 286 783 287 784
rect 291 783 292 787
rect 1430 787 1436 788
rect 1430 783 1431 787
rect 1435 786 1436 787
rect 1439 787 1445 788
rect 1439 786 1440 787
rect 1435 784 1440 786
rect 1435 783 1436 784
rect 286 782 292 783
rect 382 782 388 783
rect 166 778 167 782
rect 171 778 172 782
rect 166 777 172 778
rect 382 778 383 782
rect 387 778 388 782
rect 622 782 628 783
rect 431 779 437 780
rect 431 778 432 779
rect 382 777 388 778
rect 408 776 432 778
rect 318 771 324 772
rect 318 767 319 771
rect 323 770 324 771
rect 408 770 410 776
rect 431 775 432 776
rect 436 775 437 779
rect 622 778 623 782
rect 627 778 628 782
rect 870 782 876 783
rect 671 779 677 780
rect 671 778 672 779
rect 622 777 628 778
rect 431 774 437 775
rect 648 776 672 778
rect 323 768 410 770
rect 542 771 548 772
rect 323 767 324 768
rect 318 766 324 767
rect 542 767 543 771
rect 547 770 548 771
rect 648 770 650 776
rect 671 775 672 776
rect 676 775 677 779
rect 870 778 871 782
rect 875 778 876 782
rect 1126 782 1132 783
rect 919 779 925 780
rect 919 778 920 779
rect 870 777 876 778
rect 671 774 677 775
rect 896 776 920 778
rect 547 768 650 770
rect 786 771 792 772
rect 547 767 548 768
rect 542 766 548 767
rect 786 767 787 771
rect 791 770 792 771
rect 896 770 898 776
rect 919 775 920 776
rect 924 775 925 779
rect 1126 778 1127 782
rect 1131 778 1132 782
rect 1390 782 1396 783
rect 1430 782 1436 783
rect 1439 783 1440 784
rect 1444 783 1445 787
rect 1439 782 1445 783
rect 1126 777 1132 778
rect 1175 779 1181 780
rect 919 774 925 775
rect 1175 775 1176 779
rect 1180 778 1181 779
rect 1262 779 1268 780
rect 1262 778 1263 779
rect 1180 776 1263 778
rect 1180 775 1181 776
rect 1175 774 1181 775
rect 1262 775 1263 776
rect 1267 775 1268 779
rect 1390 778 1391 782
rect 1395 778 1396 782
rect 1390 777 1396 778
rect 1262 774 1268 775
rect 791 768 898 770
rect 791 767 792 768
rect 786 766 792 767
rect 110 765 116 766
rect 110 761 111 765
rect 115 761 116 765
rect 110 760 116 761
rect 1566 765 1572 766
rect 1566 761 1567 765
rect 1571 761 1572 765
rect 1566 760 1572 761
rect 110 747 116 748
rect 110 743 111 747
rect 115 743 116 747
rect 110 742 116 743
rect 1566 747 1572 748
rect 1566 743 1567 747
rect 1571 743 1572 747
rect 1566 742 1572 743
rect 166 736 172 737
rect 382 736 388 737
rect 622 736 628 737
rect 870 736 876 737
rect 1126 736 1132 737
rect 1390 736 1396 737
rect 166 732 167 736
rect 171 732 172 736
rect 318 735 324 736
rect 318 734 319 735
rect 237 732 319 734
rect 166 731 172 732
rect 318 731 319 732
rect 323 731 324 735
rect 382 732 383 736
rect 387 732 388 736
rect 542 735 548 736
rect 542 734 543 735
rect 453 732 543 734
rect 382 731 388 732
rect 542 731 543 732
rect 547 731 548 735
rect 622 732 623 736
rect 627 732 628 736
rect 786 735 792 736
rect 786 734 787 735
rect 693 732 787 734
rect 622 731 628 732
rect 786 731 787 732
rect 791 731 792 735
rect 870 732 871 736
rect 875 732 876 736
rect 870 731 876 732
rect 902 735 908 736
rect 902 731 903 735
rect 907 731 908 735
rect 1126 732 1127 736
rect 1131 732 1132 736
rect 1126 731 1132 732
rect 1158 735 1164 736
rect 1158 731 1159 735
rect 1163 731 1164 735
rect 1390 732 1391 736
rect 1395 732 1396 736
rect 1390 731 1396 732
rect 1446 735 1452 736
rect 1446 731 1447 735
rect 1451 731 1452 735
rect 318 730 324 731
rect 542 730 548 731
rect 786 730 792 731
rect 902 730 908 731
rect 1158 730 1164 731
rect 1446 730 1452 731
rect 318 704 324 705
rect 318 700 319 704
rect 323 700 324 704
rect 318 699 324 700
rect 574 704 580 705
rect 838 704 844 705
rect 1118 704 1124 705
rect 1398 704 1404 705
rect 574 700 575 704
rect 579 700 580 704
rect 574 699 580 700
rect 606 703 612 704
rect 606 699 607 703
rect 611 699 612 703
rect 838 700 839 704
rect 843 700 844 704
rect 838 699 844 700
rect 854 703 860 704
rect 854 699 855 703
rect 859 702 860 703
rect 859 700 873 702
rect 1118 700 1119 704
rect 1123 700 1124 704
rect 859 699 860 700
rect 1118 699 1124 700
rect 1150 703 1156 704
rect 1150 699 1151 703
rect 1155 699 1156 703
rect 1398 700 1399 704
rect 1403 700 1404 704
rect 1398 699 1404 700
rect 1454 703 1460 704
rect 1454 699 1455 703
rect 1459 699 1460 703
rect 606 698 612 699
rect 854 698 860 699
rect 1150 698 1156 699
rect 1454 698 1460 699
rect 110 693 116 694
rect 110 689 111 693
rect 115 689 116 693
rect 110 688 116 689
rect 1566 693 1572 694
rect 1566 689 1567 693
rect 1571 689 1572 693
rect 1566 688 1572 689
rect 359 687 365 688
rect 359 683 360 687
rect 364 686 365 687
rect 978 687 984 688
rect 978 686 979 687
rect 364 684 979 686
rect 364 683 365 684
rect 359 682 365 683
rect 978 683 979 684
rect 983 683 984 687
rect 978 682 984 683
rect 110 675 116 676
rect 110 671 111 675
rect 115 671 116 675
rect 110 670 116 671
rect 1566 675 1572 676
rect 1566 671 1567 675
rect 1571 671 1572 675
rect 1566 670 1572 671
rect 887 659 893 660
rect 318 658 324 659
rect 318 654 319 658
rect 323 654 324 658
rect 318 653 324 654
rect 574 658 580 659
rect 574 654 575 658
rect 579 654 580 658
rect 574 653 580 654
rect 838 658 844 659
rect 838 654 839 658
rect 843 654 844 658
rect 887 655 888 659
rect 892 658 893 659
rect 902 659 908 660
rect 1446 659 1453 660
rect 902 658 903 659
rect 892 656 903 658
rect 892 655 893 656
rect 887 654 893 655
rect 902 655 903 656
rect 907 655 908 659
rect 902 654 908 655
rect 1118 658 1124 659
rect 1118 654 1119 658
rect 1123 654 1124 658
rect 838 653 844 654
rect 1118 653 1124 654
rect 1398 658 1404 659
rect 1398 654 1399 658
rect 1403 654 1404 658
rect 1446 655 1447 659
rect 1452 655 1453 659
rect 1446 654 1453 655
rect 1398 653 1404 654
rect 367 651 373 652
rect 367 647 368 651
rect 372 650 373 651
rect 606 651 612 652
rect 606 650 607 651
rect 372 648 607 650
rect 372 647 373 648
rect 367 646 373 647
rect 606 647 607 648
rect 611 647 612 651
rect 606 646 612 647
rect 623 651 629 652
rect 623 647 624 651
rect 628 650 629 651
rect 854 651 860 652
rect 854 650 855 651
rect 628 648 855 650
rect 628 647 629 648
rect 623 646 629 647
rect 854 647 855 648
rect 859 647 860 651
rect 854 646 860 647
rect 978 651 984 652
rect 978 647 979 651
rect 983 650 984 651
rect 1167 651 1173 652
rect 1167 650 1168 651
rect 983 648 1168 650
rect 983 647 984 648
rect 978 646 984 647
rect 1167 647 1168 648
rect 1172 647 1173 651
rect 1167 646 1173 647
rect 1103 627 1109 628
rect 1103 623 1104 627
rect 1108 626 1109 627
rect 1150 627 1156 628
rect 1150 626 1151 627
rect 1108 624 1151 626
rect 1108 623 1109 624
rect 582 622 588 623
rect 582 618 583 622
rect 587 618 588 622
rect 726 622 732 623
rect 582 617 588 618
rect 631 619 637 620
rect 631 615 632 619
rect 636 618 637 619
rect 726 618 727 622
rect 731 618 732 622
rect 886 622 892 623
rect 636 616 698 618
rect 726 617 732 618
rect 775 619 781 620
rect 636 615 637 616
rect 631 614 637 615
rect 696 610 698 616
rect 775 615 776 619
rect 780 618 781 619
rect 886 618 887 622
rect 891 618 892 622
rect 1054 622 1060 623
rect 1103 622 1109 623
rect 1150 623 1151 624
rect 1155 623 1156 627
rect 1454 627 1461 628
rect 1454 623 1455 627
rect 1460 623 1461 627
rect 1150 622 1156 623
rect 1230 622 1236 623
rect 780 616 850 618
rect 886 617 892 618
rect 935 619 941 620
rect 780 615 781 616
rect 775 614 781 615
rect 742 611 748 612
rect 742 610 743 611
rect 696 608 743 610
rect 742 607 743 608
rect 747 607 748 611
rect 848 610 850 616
rect 935 615 936 619
rect 940 618 941 619
rect 1054 618 1055 622
rect 1059 618 1060 622
rect 940 616 1014 618
rect 1054 617 1060 618
rect 1230 618 1231 622
rect 1235 618 1236 622
rect 1406 622 1412 623
rect 1454 622 1461 623
rect 1230 617 1236 618
rect 1274 619 1285 620
rect 940 615 941 616
rect 935 614 941 615
rect 902 611 908 612
rect 902 610 903 611
rect 848 608 903 610
rect 742 606 748 607
rect 902 607 903 608
rect 907 607 908 611
rect 1012 610 1014 616
rect 1274 615 1275 619
rect 1279 615 1280 619
rect 1284 615 1285 619
rect 1406 618 1407 622
rect 1411 618 1412 622
rect 1406 617 1412 618
rect 1274 614 1285 615
rect 1070 611 1076 612
rect 1070 610 1071 611
rect 1012 608 1071 610
rect 902 606 908 607
rect 1070 607 1071 608
rect 1075 607 1076 611
rect 1070 606 1076 607
rect 110 605 116 606
rect 110 601 111 605
rect 115 601 116 605
rect 110 600 116 601
rect 1566 605 1572 606
rect 1566 601 1567 605
rect 1571 601 1572 605
rect 1566 600 1572 601
rect 110 587 116 588
rect 110 583 111 587
rect 115 583 116 587
rect 110 582 116 583
rect 1566 587 1572 588
rect 1566 583 1567 587
rect 1571 583 1572 587
rect 1566 582 1572 583
rect 582 576 588 577
rect 726 576 732 577
rect 886 576 892 577
rect 1054 576 1060 577
rect 1230 576 1236 577
rect 1406 576 1412 577
rect 582 572 583 576
rect 587 572 588 576
rect 582 571 588 572
rect 650 575 656 576
rect 650 571 651 575
rect 655 571 656 575
rect 726 572 727 576
rect 731 572 732 576
rect 726 571 732 572
rect 742 575 748 576
rect 742 571 743 575
rect 747 574 748 575
rect 747 572 761 574
rect 886 572 887 576
rect 891 572 892 576
rect 747 571 748 572
rect 886 571 892 572
rect 902 575 908 576
rect 902 571 903 575
rect 907 574 908 575
rect 907 572 921 574
rect 1054 572 1055 576
rect 1059 572 1060 576
rect 907 571 908 572
rect 1054 571 1060 572
rect 1070 575 1076 576
rect 1070 571 1071 575
rect 1075 574 1076 575
rect 1075 572 1089 574
rect 1230 572 1231 576
rect 1235 572 1236 576
rect 1075 571 1076 572
rect 1230 571 1236 572
rect 1262 575 1268 576
rect 1262 571 1263 575
rect 1267 571 1268 575
rect 1406 572 1407 576
rect 1411 572 1412 576
rect 1406 571 1412 572
rect 1438 575 1444 576
rect 1438 571 1439 575
rect 1443 571 1444 575
rect 650 570 656 571
rect 742 570 748 571
rect 902 570 908 571
rect 1070 570 1076 571
rect 1262 570 1268 571
rect 1438 570 1444 571
rect 758 544 764 545
rect 862 544 868 545
rect 974 544 980 545
rect 1086 544 1092 545
rect 1206 544 1212 545
rect 1326 544 1332 545
rect 1446 544 1452 545
rect 758 540 759 544
rect 763 540 764 544
rect 758 539 764 540
rect 826 543 832 544
rect 826 539 827 543
rect 831 539 832 543
rect 862 540 863 544
rect 867 540 868 544
rect 862 539 868 540
rect 930 543 936 544
rect 930 539 931 543
rect 935 539 936 543
rect 974 540 975 544
rect 979 540 980 544
rect 974 539 980 540
rect 1042 543 1048 544
rect 1042 539 1043 543
rect 1047 539 1048 543
rect 1086 540 1087 544
rect 1091 540 1092 544
rect 1086 539 1092 540
rect 1118 543 1124 544
rect 1118 539 1119 543
rect 1123 539 1124 543
rect 1206 540 1207 544
rect 1211 540 1212 544
rect 1206 539 1212 540
rect 1274 543 1280 544
rect 1274 539 1275 543
rect 1279 539 1280 543
rect 1326 540 1327 544
rect 1331 540 1332 544
rect 1326 539 1332 540
rect 1394 543 1400 544
rect 1394 539 1395 543
rect 1399 539 1400 543
rect 1446 540 1447 544
rect 1451 540 1452 544
rect 1446 539 1452 540
rect 1510 543 1516 544
rect 1510 539 1511 543
rect 1515 539 1516 543
rect 826 538 832 539
rect 930 538 936 539
rect 1042 538 1048 539
rect 1118 538 1124 539
rect 1274 538 1280 539
rect 1394 538 1400 539
rect 1510 538 1516 539
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 1566 533 1572 534
rect 1566 529 1567 533
rect 1571 529 1572 533
rect 1566 528 1572 529
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 1566 515 1572 516
rect 1566 511 1567 515
rect 1571 511 1572 515
rect 1566 510 1572 511
rect 650 507 656 508
rect 650 503 651 507
rect 655 506 656 507
rect 655 504 786 506
rect 655 503 656 504
rect 650 502 656 503
rect 758 498 764 499
rect 758 494 759 498
rect 763 494 764 498
rect 784 498 786 504
rect 807 499 813 500
rect 1375 499 1381 500
rect 807 498 808 499
rect 784 496 808 498
rect 807 495 808 496
rect 812 495 813 499
rect 807 494 813 495
rect 862 498 868 499
rect 862 494 863 498
rect 867 494 868 498
rect 758 493 764 494
rect 862 493 868 494
rect 974 498 980 499
rect 974 494 975 498
rect 979 494 980 498
rect 974 493 980 494
rect 1086 498 1092 499
rect 1086 494 1087 498
rect 1091 494 1092 498
rect 1086 493 1092 494
rect 1206 498 1212 499
rect 1206 494 1207 498
rect 1211 494 1212 498
rect 1206 493 1212 494
rect 1326 498 1332 499
rect 1326 494 1327 498
rect 1331 494 1332 498
rect 1375 495 1376 499
rect 1380 498 1381 499
rect 1438 499 1444 500
rect 1438 498 1439 499
rect 1380 496 1439 498
rect 1380 495 1381 496
rect 1375 494 1381 495
rect 1438 495 1439 496
rect 1443 495 1444 499
rect 1438 494 1444 495
rect 1446 498 1452 499
rect 1446 494 1447 498
rect 1451 494 1452 498
rect 1326 493 1332 494
rect 1446 493 1452 494
rect 826 491 832 492
rect 826 487 827 491
rect 831 490 832 491
rect 911 491 917 492
rect 911 490 912 491
rect 831 488 912 490
rect 831 487 832 488
rect 826 486 832 487
rect 911 487 912 488
rect 916 487 917 491
rect 911 486 917 487
rect 930 491 936 492
rect 930 487 931 491
rect 935 490 936 491
rect 1023 491 1029 492
rect 1023 490 1024 491
rect 935 488 1024 490
rect 935 487 936 488
rect 930 486 936 487
rect 1023 487 1024 488
rect 1028 487 1029 491
rect 1023 486 1029 487
rect 1042 491 1048 492
rect 1042 487 1043 491
rect 1047 490 1048 491
rect 1135 491 1141 492
rect 1135 490 1136 491
rect 1047 488 1136 490
rect 1047 487 1048 488
rect 1042 486 1048 487
rect 1135 487 1136 488
rect 1140 487 1141 491
rect 1135 486 1141 487
rect 1214 491 1220 492
rect 1214 487 1215 491
rect 1219 490 1220 491
rect 1255 491 1261 492
rect 1255 490 1256 491
rect 1219 488 1256 490
rect 1219 487 1220 488
rect 1214 486 1220 487
rect 1255 487 1256 488
rect 1260 487 1261 491
rect 1255 486 1261 487
rect 1394 491 1400 492
rect 1394 487 1395 491
rect 1399 490 1400 491
rect 1495 491 1501 492
rect 1495 490 1496 491
rect 1399 488 1496 490
rect 1399 487 1400 488
rect 1394 486 1400 487
rect 1495 487 1496 488
rect 1500 487 1501 491
rect 1495 486 1501 487
rect 1079 467 1085 468
rect 1079 463 1080 467
rect 1084 466 1085 467
rect 1118 467 1124 468
rect 1118 466 1119 467
rect 1084 464 1119 466
rect 1084 463 1085 464
rect 718 462 724 463
rect 718 458 719 462
rect 723 458 724 462
rect 822 462 828 463
rect 718 457 724 458
rect 767 459 773 460
rect 767 455 768 459
rect 772 458 773 459
rect 822 458 823 462
rect 827 458 828 462
rect 926 462 932 463
rect 772 456 814 458
rect 822 457 828 458
rect 871 459 877 460
rect 772 455 773 456
rect 767 454 773 455
rect 812 450 814 456
rect 871 455 872 459
rect 876 458 877 459
rect 926 458 927 462
rect 931 458 932 462
rect 1030 462 1036 463
rect 1079 462 1085 463
rect 1118 463 1119 464
rect 1123 463 1124 467
rect 1510 467 1517 468
rect 1510 463 1511 467
rect 1516 463 1517 467
rect 1118 462 1124 463
rect 1134 462 1140 463
rect 876 456 918 458
rect 926 457 932 458
rect 975 459 981 460
rect 876 455 877 456
rect 871 454 877 455
rect 838 451 844 452
rect 838 450 839 451
rect 812 448 839 450
rect 838 447 839 448
rect 843 447 844 451
rect 916 450 918 456
rect 975 455 976 459
rect 980 458 981 459
rect 1030 458 1031 462
rect 1035 458 1036 462
rect 980 456 1022 458
rect 1030 457 1036 458
rect 1134 458 1135 462
rect 1139 458 1140 462
rect 1238 462 1244 463
rect 1134 457 1140 458
rect 1183 459 1189 460
rect 980 455 981 456
rect 975 454 981 455
rect 942 451 948 452
rect 942 450 943 451
rect 916 448 943 450
rect 838 446 844 447
rect 942 447 943 448
rect 947 447 948 451
rect 1020 450 1022 456
rect 1183 455 1184 459
rect 1188 458 1189 459
rect 1238 458 1239 462
rect 1243 458 1244 462
rect 1350 462 1356 463
rect 1188 456 1230 458
rect 1238 457 1244 458
rect 1287 459 1293 460
rect 1188 455 1189 456
rect 1183 454 1189 455
rect 1046 451 1052 452
rect 1046 450 1047 451
rect 1020 448 1047 450
rect 942 446 948 447
rect 1046 447 1047 448
rect 1051 447 1052 451
rect 1228 450 1230 456
rect 1287 455 1288 459
rect 1292 458 1293 459
rect 1350 458 1351 462
rect 1355 458 1356 462
rect 1462 462 1468 463
rect 1510 462 1517 463
rect 1292 456 1338 458
rect 1350 457 1356 458
rect 1399 459 1405 460
rect 1292 455 1293 456
rect 1287 454 1293 455
rect 1254 451 1260 452
rect 1254 450 1255 451
rect 1228 448 1255 450
rect 1046 446 1052 447
rect 1254 447 1255 448
rect 1259 447 1260 451
rect 1336 450 1338 456
rect 1399 455 1400 459
rect 1404 458 1405 459
rect 1462 458 1463 462
rect 1467 458 1468 462
rect 1404 456 1442 458
rect 1462 457 1468 458
rect 1404 455 1405 456
rect 1399 454 1405 455
rect 1366 451 1372 452
rect 1366 450 1367 451
rect 1336 448 1367 450
rect 1254 446 1260 447
rect 1366 447 1367 448
rect 1371 447 1372 451
rect 1440 450 1442 456
rect 1478 451 1484 452
rect 1478 450 1479 451
rect 1440 448 1479 450
rect 1366 446 1372 447
rect 1478 447 1479 448
rect 1483 447 1484 451
rect 1478 446 1484 447
rect 110 445 116 446
rect 110 441 111 445
rect 115 441 116 445
rect 110 440 116 441
rect 1566 445 1572 446
rect 1566 441 1567 445
rect 1571 441 1572 445
rect 1566 440 1572 441
rect 110 427 116 428
rect 110 423 111 427
rect 115 423 116 427
rect 110 422 116 423
rect 1566 427 1572 428
rect 1566 423 1567 427
rect 1571 423 1572 427
rect 1566 422 1572 423
rect 718 416 724 417
rect 822 416 828 417
rect 926 416 932 417
rect 1030 416 1036 417
rect 1134 416 1140 417
rect 1238 416 1244 417
rect 1350 416 1356 417
rect 1462 416 1468 417
rect 718 412 719 416
rect 723 412 724 416
rect 798 415 804 416
rect 798 414 799 415
rect 789 412 799 414
rect 718 411 724 412
rect 798 411 799 412
rect 803 411 804 415
rect 822 412 823 416
rect 827 412 828 416
rect 822 411 828 412
rect 838 415 844 416
rect 838 411 839 415
rect 843 414 844 415
rect 843 412 857 414
rect 926 412 927 416
rect 931 412 932 416
rect 843 411 844 412
rect 926 411 932 412
rect 942 415 948 416
rect 942 411 943 415
rect 947 414 948 415
rect 947 412 961 414
rect 1030 412 1031 416
rect 1035 412 1036 416
rect 947 411 948 412
rect 1030 411 1036 412
rect 1046 415 1052 416
rect 1046 411 1047 415
rect 1051 414 1052 415
rect 1051 412 1065 414
rect 1134 412 1135 416
rect 1139 412 1140 416
rect 1214 415 1220 416
rect 1214 414 1215 415
rect 1205 412 1215 414
rect 1051 411 1052 412
rect 1134 411 1140 412
rect 1214 411 1215 412
rect 1219 411 1220 415
rect 1238 412 1239 416
rect 1243 412 1244 416
rect 1238 411 1244 412
rect 1254 415 1260 416
rect 1254 411 1255 415
rect 1259 414 1260 415
rect 1259 412 1273 414
rect 1350 412 1351 416
rect 1355 412 1356 416
rect 1259 411 1260 412
rect 1350 411 1356 412
rect 1366 415 1372 416
rect 1366 411 1367 415
rect 1371 414 1372 415
rect 1371 412 1385 414
rect 1462 412 1463 416
rect 1467 412 1468 416
rect 1371 411 1372 412
rect 1462 411 1468 412
rect 1478 415 1484 416
rect 1478 411 1479 415
rect 1483 414 1484 415
rect 1483 412 1497 414
rect 1483 411 1484 412
rect 798 410 804 411
rect 838 410 844 411
rect 942 410 948 411
rect 1046 410 1052 411
rect 1214 410 1220 411
rect 1254 410 1260 411
rect 1366 410 1372 411
rect 1478 410 1484 411
rect 510 376 516 377
rect 598 376 604 377
rect 686 376 692 377
rect 774 376 780 377
rect 510 372 511 376
rect 515 372 516 376
rect 510 371 516 372
rect 578 375 584 376
rect 578 371 579 375
rect 583 371 584 375
rect 598 372 599 376
rect 603 372 604 376
rect 598 371 604 372
rect 630 375 636 376
rect 630 371 631 375
rect 635 371 636 375
rect 686 372 687 376
rect 691 372 692 376
rect 686 371 692 372
rect 702 375 708 376
rect 702 371 703 375
rect 707 374 708 375
rect 707 372 721 374
rect 774 372 775 376
rect 779 372 780 376
rect 707 371 708 372
rect 774 371 780 372
rect 806 375 812 376
rect 806 371 807 375
rect 811 371 812 375
rect 578 370 584 371
rect 630 370 636 371
rect 702 370 708 371
rect 806 370 812 371
rect 110 365 116 366
rect 110 361 111 365
rect 115 361 116 365
rect 110 360 116 361
rect 1566 365 1572 366
rect 1566 361 1567 365
rect 1571 361 1572 365
rect 1566 360 1572 361
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 110 342 116 343
rect 1566 347 1572 348
rect 1566 343 1567 347
rect 1571 343 1572 347
rect 1566 342 1572 343
rect 798 331 804 332
rect 510 330 516 331
rect 510 326 511 330
rect 515 326 516 330
rect 510 325 516 326
rect 598 330 604 331
rect 598 326 599 330
rect 603 326 604 330
rect 598 325 604 326
rect 686 330 692 331
rect 686 326 687 330
rect 691 326 692 330
rect 686 325 692 326
rect 774 330 780 331
rect 774 326 775 330
rect 779 326 780 330
rect 798 327 799 331
rect 803 330 804 331
rect 823 331 829 332
rect 823 330 824 331
rect 803 328 824 330
rect 803 327 804 328
rect 798 326 804 327
rect 823 327 824 328
rect 828 327 829 331
rect 823 326 829 327
rect 774 325 780 326
rect 559 323 565 324
rect 559 319 560 323
rect 564 322 565 323
rect 630 323 636 324
rect 630 322 631 323
rect 564 320 631 322
rect 564 319 565 320
rect 559 318 565 319
rect 630 319 631 320
rect 635 319 636 323
rect 630 318 636 319
rect 647 323 653 324
rect 647 319 648 323
rect 652 322 653 323
rect 702 323 708 324
rect 702 322 703 323
rect 652 320 703 322
rect 652 319 653 320
rect 647 318 653 319
rect 702 319 703 320
rect 707 319 708 323
rect 702 318 708 319
rect 735 323 741 324
rect 735 319 736 323
rect 740 322 741 323
rect 806 323 812 324
rect 806 322 807 323
rect 740 320 807 322
rect 740 319 741 320
rect 735 318 741 319
rect 806 319 807 320
rect 811 319 812 323
rect 806 318 812 319
rect 578 303 584 304
rect 578 299 579 303
rect 583 302 584 303
rect 599 303 605 304
rect 599 302 600 303
rect 583 300 600 302
rect 583 299 584 300
rect 374 298 380 299
rect 374 294 375 298
rect 379 294 380 298
rect 462 298 468 299
rect 374 293 380 294
rect 423 295 429 296
rect 423 291 424 295
rect 428 294 429 295
rect 462 294 463 298
rect 467 294 468 298
rect 550 298 556 299
rect 578 298 584 299
rect 599 299 600 300
rect 604 299 605 303
rect 599 298 605 299
rect 428 292 458 294
rect 462 293 468 294
rect 511 295 517 296
rect 428 291 429 292
rect 423 290 429 291
rect 456 286 458 292
rect 511 291 512 295
rect 516 294 517 295
rect 550 294 551 298
rect 555 294 556 298
rect 516 292 546 294
rect 550 293 556 294
rect 516 291 517 292
rect 511 290 517 291
rect 478 287 484 288
rect 478 286 479 287
rect 456 284 479 286
rect 478 283 479 284
rect 483 283 484 287
rect 544 286 546 292
rect 566 287 572 288
rect 566 286 567 287
rect 544 284 567 286
rect 478 282 484 283
rect 566 283 567 284
rect 571 283 572 287
rect 566 282 572 283
rect 110 281 116 282
rect 110 277 111 281
rect 115 277 116 281
rect 110 276 116 277
rect 1566 281 1572 282
rect 1566 277 1567 281
rect 1571 277 1572 281
rect 1566 276 1572 277
rect 110 263 116 264
rect 110 259 111 263
rect 115 259 116 263
rect 110 258 116 259
rect 1566 263 1572 264
rect 1566 259 1567 263
rect 1571 259 1572 263
rect 1566 258 1572 259
rect 374 252 380 253
rect 462 252 468 253
rect 550 252 556 253
rect 374 248 375 252
rect 379 248 380 252
rect 374 247 380 248
rect 406 251 412 252
rect 406 247 407 251
rect 411 247 412 251
rect 462 248 463 252
rect 467 248 468 252
rect 462 247 468 248
rect 478 251 484 252
rect 478 247 479 251
rect 483 250 484 251
rect 483 248 497 250
rect 550 248 551 252
rect 555 248 556 252
rect 483 247 484 248
rect 550 247 556 248
rect 566 251 572 252
rect 566 247 567 251
rect 571 250 572 251
rect 571 248 585 250
rect 571 247 572 248
rect 406 246 412 247
rect 478 246 484 247
rect 566 246 572 247
rect 246 240 252 241
rect 246 236 247 240
rect 251 236 252 240
rect 246 235 252 236
rect 334 240 340 241
rect 422 240 428 241
rect 334 236 335 240
rect 339 236 340 240
rect 334 235 340 236
rect 366 239 372 240
rect 366 235 367 239
rect 371 235 372 239
rect 422 236 423 240
rect 427 236 428 240
rect 582 239 588 240
rect 582 238 583 239
rect 493 236 583 238
rect 422 235 428 236
rect 582 235 583 236
rect 587 235 588 239
rect 366 234 372 235
rect 582 234 588 235
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 1566 229 1572 230
rect 1566 225 1567 229
rect 1571 225 1572 229
rect 1566 224 1572 225
rect 287 223 293 224
rect 287 219 288 223
rect 292 222 293 223
rect 447 223 453 224
rect 447 222 448 223
rect 292 220 448 222
rect 292 219 293 220
rect 287 218 293 219
rect 447 219 448 220
rect 452 219 453 223
rect 447 218 453 219
rect 110 211 116 212
rect 110 207 111 211
rect 115 207 116 211
rect 110 206 116 207
rect 1566 211 1572 212
rect 1566 207 1567 211
rect 1571 207 1572 211
rect 1566 206 1572 207
rect 383 195 389 196
rect 246 194 252 195
rect 246 190 247 194
rect 251 190 252 194
rect 246 189 252 190
rect 334 194 340 195
rect 334 190 335 194
rect 339 190 340 194
rect 383 191 384 195
rect 388 194 389 195
rect 406 195 412 196
rect 447 195 453 196
rect 406 194 407 195
rect 388 192 407 194
rect 388 191 389 192
rect 383 190 389 191
rect 406 191 407 192
rect 411 191 412 195
rect 406 190 412 191
rect 422 194 428 195
rect 422 190 423 194
rect 427 190 428 194
rect 447 191 448 195
rect 452 194 453 195
rect 471 195 477 196
rect 471 194 472 195
rect 452 192 472 194
rect 452 191 453 192
rect 447 190 453 191
rect 471 191 472 192
rect 476 191 477 195
rect 471 190 477 191
rect 334 189 340 190
rect 422 189 428 190
rect 295 187 301 188
rect 295 183 296 187
rect 300 186 301 187
rect 366 187 372 188
rect 366 186 367 187
rect 300 184 367 186
rect 300 183 301 184
rect 295 182 301 183
rect 366 183 367 184
rect 371 183 372 187
rect 366 182 372 183
rect 582 147 588 148
rect 582 143 583 147
rect 587 146 588 147
rect 623 147 629 148
rect 623 146 624 147
rect 587 144 624 146
rect 587 143 588 144
rect 134 142 140 143
rect 134 138 135 142
rect 139 138 140 142
rect 222 142 228 143
rect 134 137 140 138
rect 183 139 189 140
rect 183 135 184 139
rect 188 138 189 139
rect 222 138 223 142
rect 227 138 228 142
rect 310 142 316 143
rect 188 136 218 138
rect 222 137 228 138
rect 271 139 277 140
rect 188 135 189 136
rect 183 134 189 135
rect 216 130 218 136
rect 271 135 272 139
rect 276 138 277 139
rect 310 138 311 142
rect 315 138 316 142
rect 398 142 404 143
rect 276 136 306 138
rect 310 137 316 138
rect 359 139 365 140
rect 276 135 277 136
rect 271 134 277 135
rect 238 131 244 132
rect 238 130 239 131
rect 216 128 239 130
rect 238 127 239 128
rect 243 127 244 131
rect 304 130 306 136
rect 359 135 360 139
rect 364 138 365 139
rect 398 138 399 142
rect 403 138 404 142
rect 486 142 492 143
rect 364 136 394 138
rect 398 137 404 138
rect 447 139 453 140
rect 364 135 365 136
rect 359 134 365 135
rect 326 131 332 132
rect 326 130 327 131
rect 304 128 327 130
rect 238 126 244 127
rect 326 127 327 128
rect 331 127 332 131
rect 392 130 394 136
rect 447 135 448 139
rect 452 138 453 139
rect 486 138 487 142
rect 491 138 492 142
rect 574 142 580 143
rect 582 142 588 143
rect 623 143 624 144
rect 628 143 629 147
rect 623 142 629 143
rect 452 136 482 138
rect 486 137 492 138
rect 535 139 541 140
rect 452 135 453 136
rect 447 134 453 135
rect 414 131 420 132
rect 414 130 415 131
rect 392 128 415 130
rect 326 126 332 127
rect 414 127 415 128
rect 419 127 420 131
rect 480 130 482 136
rect 535 135 536 139
rect 540 138 541 139
rect 574 138 575 142
rect 579 138 580 142
rect 540 136 563 138
rect 574 137 580 138
rect 540 135 541 136
rect 535 134 541 135
rect 502 131 508 132
rect 502 130 503 131
rect 480 128 503 130
rect 414 126 420 127
rect 502 127 503 128
rect 507 127 508 131
rect 561 130 563 136
rect 590 131 596 132
rect 590 130 591 131
rect 561 128 591 130
rect 502 126 508 127
rect 590 127 591 128
rect 595 127 596 131
rect 590 126 596 127
rect 110 125 116 126
rect 110 121 111 125
rect 115 121 116 125
rect 110 120 116 121
rect 1566 125 1572 126
rect 1566 121 1567 125
rect 1571 121 1572 125
rect 1566 120 1572 121
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 110 102 116 103
rect 1566 107 1572 108
rect 1566 103 1567 107
rect 1571 103 1572 107
rect 1566 102 1572 103
rect 134 96 140 97
rect 134 92 135 96
rect 139 92 140 96
rect 134 91 140 92
rect 222 96 228 97
rect 310 96 316 97
rect 398 96 404 97
rect 486 96 492 97
rect 574 96 580 97
rect 222 92 223 96
rect 227 92 228 96
rect 222 91 228 92
rect 238 95 244 96
rect 238 91 239 95
rect 243 94 244 95
rect 243 92 257 94
rect 310 92 311 96
rect 315 92 316 96
rect 243 91 244 92
rect 310 91 316 92
rect 326 95 332 96
rect 326 91 327 95
rect 331 94 332 95
rect 331 92 345 94
rect 398 92 399 96
rect 403 92 404 96
rect 331 91 332 92
rect 398 91 404 92
rect 414 95 420 96
rect 414 91 415 95
rect 419 94 420 95
rect 419 92 433 94
rect 486 92 487 96
rect 491 92 492 96
rect 419 91 420 92
rect 486 91 492 92
rect 502 95 508 96
rect 502 91 503 95
rect 507 94 508 95
rect 507 92 521 94
rect 574 92 575 96
rect 579 92 580 96
rect 507 91 508 92
rect 574 91 580 92
rect 590 95 596 96
rect 590 91 591 95
rect 595 94 596 95
rect 595 92 609 94
rect 595 91 596 92
rect 238 90 244 91
rect 326 90 332 91
rect 414 90 420 91
rect 502 90 508 91
rect 590 90 596 91
<< m3c >>
rect 399 1506 403 1510
rect 487 1506 491 1510
rect 575 1506 579 1510
rect 503 1495 507 1499
rect 671 1506 675 1510
rect 591 1495 595 1499
rect 783 1506 787 1510
rect 687 1495 691 1499
rect 903 1506 907 1510
rect 799 1495 803 1499
rect 1031 1506 1035 1510
rect 919 1495 923 1499
rect 1167 1506 1171 1510
rect 1047 1495 1051 1499
rect 1211 1503 1215 1507
rect 1303 1506 1307 1510
rect 1447 1506 1451 1510
rect 1183 1495 1187 1499
rect 1415 1495 1419 1499
rect 111 1489 115 1493
rect 1567 1489 1571 1493
rect 111 1471 115 1475
rect 1567 1471 1571 1475
rect 399 1460 403 1464
rect 467 1459 471 1463
rect 487 1460 491 1464
rect 503 1459 507 1463
rect 575 1460 579 1464
rect 591 1459 595 1463
rect 671 1460 675 1464
rect 687 1459 691 1463
rect 783 1460 787 1464
rect 799 1459 803 1463
rect 903 1460 907 1464
rect 919 1459 923 1463
rect 1031 1460 1035 1464
rect 1047 1459 1051 1463
rect 1167 1460 1171 1464
rect 1183 1459 1187 1463
rect 1303 1460 1307 1464
rect 1415 1459 1419 1463
rect 1447 1460 1451 1464
rect 1479 1459 1483 1463
rect 423 1436 427 1440
rect 655 1436 659 1440
rect 723 1435 727 1439
rect 895 1436 899 1440
rect 911 1435 915 1439
rect 1143 1436 1147 1440
rect 1211 1435 1215 1439
rect 1399 1436 1403 1440
rect 1439 1435 1443 1439
rect 111 1425 115 1429
rect 1567 1425 1571 1429
rect 111 1407 115 1411
rect 1567 1407 1571 1411
rect 423 1390 427 1394
rect 467 1391 471 1395
rect 655 1390 659 1394
rect 895 1390 899 1394
rect 1143 1390 1147 1394
rect 1399 1390 1403 1394
rect 1479 1391 1483 1395
rect 723 1383 727 1387
rect 1191 1383 1192 1387
rect 1192 1383 1195 1387
rect 471 1362 475 1366
rect 911 1367 915 1371
rect 1439 1367 1440 1371
rect 1440 1367 1443 1371
rect 695 1362 699 1366
rect 919 1362 923 1366
rect 1007 1359 1011 1363
rect 1151 1362 1155 1366
rect 711 1351 715 1355
rect 1391 1362 1395 1366
rect 111 1345 115 1349
rect 1567 1345 1571 1349
rect 111 1327 115 1331
rect 1567 1327 1571 1331
rect 471 1316 475 1320
rect 695 1316 699 1320
rect 711 1315 715 1319
rect 919 1316 923 1320
rect 1151 1316 1155 1320
rect 1191 1315 1195 1319
rect 1391 1316 1395 1320
rect 1423 1315 1427 1319
rect 519 1296 523 1300
rect 587 1295 591 1299
rect 743 1296 747 1300
rect 811 1295 815 1299
rect 975 1296 979 1300
rect 1007 1295 1011 1299
rect 1207 1296 1211 1300
rect 1275 1295 1279 1299
rect 1439 1296 1443 1300
rect 1471 1295 1475 1299
rect 111 1285 115 1289
rect 1567 1285 1571 1289
rect 111 1267 115 1271
rect 1567 1267 1571 1271
rect 519 1250 523 1254
rect 743 1250 747 1254
rect 975 1250 979 1254
rect 1207 1250 1211 1254
rect 1423 1251 1427 1255
rect 1439 1250 1443 1254
rect 587 1243 591 1247
rect 1191 1243 1195 1247
rect 1275 1243 1279 1247
rect 811 1219 815 1223
rect 567 1210 571 1214
rect 767 1210 771 1214
rect 967 1210 971 1214
rect 1175 1210 1179 1214
rect 1471 1215 1475 1219
rect 783 1199 787 1203
rect 1255 1207 1259 1211
rect 1391 1210 1395 1214
rect 983 1199 987 1203
rect 111 1193 115 1197
rect 1567 1193 1571 1197
rect 111 1175 115 1179
rect 1567 1175 1571 1179
rect 567 1164 571 1168
rect 727 1163 731 1167
rect 767 1164 771 1168
rect 783 1163 787 1167
rect 967 1164 971 1168
rect 983 1163 987 1167
rect 1175 1164 1179 1168
rect 1191 1163 1195 1167
rect 1391 1164 1395 1168
rect 1455 1163 1459 1167
rect 703 1152 707 1156
rect 979 1151 983 1155
rect 1055 1152 1059 1156
rect 1079 1151 1083 1155
rect 1407 1152 1411 1156
rect 1463 1151 1467 1155
rect 111 1141 115 1145
rect 1567 1141 1571 1145
rect 111 1123 115 1127
rect 1567 1123 1571 1127
rect 703 1106 707 1110
rect 727 1107 731 1111
rect 1055 1106 1059 1110
rect 1407 1106 1411 1110
rect 1455 1107 1456 1111
rect 1456 1107 1459 1111
rect 979 1099 983 1103
rect 1079 1087 1080 1091
rect 1080 1087 1083 1091
rect 1463 1087 1464 1091
rect 1464 1087 1467 1091
rect 671 1082 675 1086
rect 847 1082 851 1086
rect 1031 1082 1035 1086
rect 1223 1082 1227 1086
rect 863 1071 867 1075
rect 1267 1079 1271 1083
rect 1415 1082 1419 1086
rect 1047 1071 1051 1075
rect 111 1065 115 1069
rect 1567 1065 1571 1069
rect 111 1047 115 1051
rect 1567 1047 1571 1051
rect 671 1036 675 1040
rect 847 1036 851 1040
rect 863 1035 867 1039
rect 1031 1036 1035 1040
rect 1047 1035 1051 1039
rect 1223 1036 1227 1040
rect 1255 1035 1259 1039
rect 1415 1036 1419 1040
rect 1455 1035 1459 1039
rect 1007 1027 1011 1031
rect 575 1008 579 1012
rect 607 1007 611 1011
rect 775 1008 779 1012
rect 807 1007 811 1011
rect 983 1008 987 1012
rect 1015 1007 1019 1011
rect 1191 1008 1195 1012
rect 1267 1007 1271 1011
rect 1407 1008 1411 1012
rect 1447 1007 1451 1011
rect 111 997 115 1001
rect 1567 997 1571 1001
rect 111 979 115 983
rect 1567 979 1571 983
rect 575 962 579 966
rect 775 962 779 966
rect 983 962 987 966
rect 1007 963 1011 967
rect 1191 962 1195 966
rect 1407 962 1411 966
rect 1455 963 1456 967
rect 1456 963 1459 967
rect 807 955 811 959
rect 1015 955 1019 959
rect 1163 955 1167 959
rect 607 935 611 939
rect 1447 935 1448 939
rect 1448 935 1451 939
rect 407 930 411 934
rect 735 930 739 934
rect 611 919 615 923
rect 1063 930 1067 934
rect 931 919 935 923
rect 1399 930 1403 934
rect 111 913 115 917
rect 1567 913 1571 917
rect 111 895 115 899
rect 1567 895 1571 899
rect 407 884 411 888
rect 611 883 615 887
rect 735 884 739 888
rect 931 883 935 887
rect 1063 884 1067 888
rect 1079 883 1083 887
rect 1399 884 1403 888
rect 1439 883 1443 887
rect 255 868 259 872
rect 287 867 291 871
rect 527 868 531 872
rect 559 867 563 871
rect 807 868 811 872
rect 839 867 843 871
rect 1095 868 1099 872
rect 1163 867 1167 871
rect 1391 868 1395 872
rect 1431 867 1435 871
rect 111 857 115 861
rect 1567 857 1571 861
rect 111 839 115 843
rect 1567 839 1571 843
rect 255 822 259 826
rect 527 822 531 826
rect 807 822 811 826
rect 1079 823 1083 827
rect 1095 822 1099 826
rect 1391 822 1395 826
rect 1439 823 1440 827
rect 1440 823 1443 827
rect 559 815 563 819
rect 839 815 843 819
rect 1159 815 1163 819
rect 287 783 291 787
rect 1431 783 1435 787
rect 167 778 171 782
rect 383 778 387 782
rect 319 767 323 771
rect 623 778 627 782
rect 543 767 547 771
rect 871 778 875 782
rect 787 767 791 771
rect 1127 778 1131 782
rect 1263 775 1267 779
rect 1391 778 1395 782
rect 111 761 115 765
rect 1567 761 1571 765
rect 111 743 115 747
rect 1567 743 1571 747
rect 167 732 171 736
rect 319 731 323 735
rect 383 732 387 736
rect 543 731 547 735
rect 623 732 627 736
rect 787 731 791 735
rect 871 732 875 736
rect 903 731 907 735
rect 1127 732 1131 736
rect 1159 731 1163 735
rect 1391 732 1395 736
rect 1447 731 1451 735
rect 319 700 323 704
rect 575 700 579 704
rect 607 699 611 703
rect 839 700 843 704
rect 855 699 859 703
rect 1119 700 1123 704
rect 1151 699 1155 703
rect 1399 700 1403 704
rect 1455 699 1459 703
rect 111 689 115 693
rect 1567 689 1571 693
rect 979 683 983 687
rect 111 671 115 675
rect 1567 671 1571 675
rect 319 654 323 658
rect 575 654 579 658
rect 839 654 843 658
rect 903 655 907 659
rect 1119 654 1123 658
rect 1399 654 1403 658
rect 1447 655 1448 659
rect 1448 655 1451 659
rect 607 647 611 651
rect 855 647 859 651
rect 979 647 983 651
rect 583 618 587 622
rect 727 618 731 622
rect 887 618 891 622
rect 1151 623 1155 627
rect 1455 623 1456 627
rect 1456 623 1459 627
rect 743 607 747 611
rect 1055 618 1059 622
rect 1231 618 1235 622
rect 903 607 907 611
rect 1275 615 1279 619
rect 1407 618 1411 622
rect 1071 607 1075 611
rect 111 601 115 605
rect 1567 601 1571 605
rect 111 583 115 587
rect 1567 583 1571 587
rect 583 572 587 576
rect 651 571 655 575
rect 727 572 731 576
rect 743 571 747 575
rect 887 572 891 576
rect 903 571 907 575
rect 1055 572 1059 576
rect 1071 571 1075 575
rect 1231 572 1235 576
rect 1263 571 1267 575
rect 1407 572 1411 576
rect 1439 571 1443 575
rect 759 540 763 544
rect 827 539 831 543
rect 863 540 867 544
rect 931 539 935 543
rect 975 540 979 544
rect 1043 539 1047 543
rect 1087 540 1091 544
rect 1119 539 1123 543
rect 1207 540 1211 544
rect 1275 539 1279 543
rect 1327 540 1331 544
rect 1395 539 1399 543
rect 1447 540 1451 544
rect 1511 539 1515 543
rect 111 529 115 533
rect 1567 529 1571 533
rect 111 511 115 515
rect 1567 511 1571 515
rect 651 503 655 507
rect 759 494 763 498
rect 863 494 867 498
rect 975 494 979 498
rect 1087 494 1091 498
rect 1207 494 1211 498
rect 1327 494 1331 498
rect 1439 495 1443 499
rect 1447 494 1451 498
rect 827 487 831 491
rect 931 487 935 491
rect 1043 487 1047 491
rect 1215 487 1219 491
rect 1395 487 1399 491
rect 719 458 723 462
rect 823 458 827 462
rect 927 458 931 462
rect 1119 463 1123 467
rect 1511 463 1512 467
rect 1512 463 1515 467
rect 839 447 843 451
rect 1031 458 1035 462
rect 1135 458 1139 462
rect 943 447 947 451
rect 1239 458 1243 462
rect 1047 447 1051 451
rect 1351 458 1355 462
rect 1255 447 1259 451
rect 1463 458 1467 462
rect 1367 447 1371 451
rect 1479 447 1483 451
rect 111 441 115 445
rect 1567 441 1571 445
rect 111 423 115 427
rect 1567 423 1571 427
rect 719 412 723 416
rect 799 411 803 415
rect 823 412 827 416
rect 839 411 843 415
rect 927 412 931 416
rect 943 411 947 415
rect 1031 412 1035 416
rect 1047 411 1051 415
rect 1135 412 1139 416
rect 1215 411 1219 415
rect 1239 412 1243 416
rect 1255 411 1259 415
rect 1351 412 1355 416
rect 1367 411 1371 415
rect 1463 412 1467 416
rect 1479 411 1483 415
rect 511 372 515 376
rect 579 371 583 375
rect 599 372 603 376
rect 631 371 635 375
rect 687 372 691 376
rect 703 371 707 375
rect 775 372 779 376
rect 807 371 811 375
rect 111 361 115 365
rect 1567 361 1571 365
rect 111 343 115 347
rect 1567 343 1571 347
rect 511 326 515 330
rect 599 326 603 330
rect 687 326 691 330
rect 775 326 779 330
rect 799 327 803 331
rect 631 319 635 323
rect 703 319 707 323
rect 807 319 811 323
rect 579 299 583 303
rect 375 294 379 298
rect 463 294 467 298
rect 551 294 555 298
rect 479 283 483 287
rect 567 283 571 287
rect 111 277 115 281
rect 1567 277 1571 281
rect 111 259 115 263
rect 1567 259 1571 263
rect 375 248 379 252
rect 407 247 411 251
rect 463 248 467 252
rect 479 247 483 251
rect 551 248 555 252
rect 567 247 571 251
rect 247 236 251 240
rect 335 236 339 240
rect 367 235 371 239
rect 423 236 427 240
rect 583 235 587 239
rect 111 225 115 229
rect 1567 225 1571 229
rect 111 207 115 211
rect 1567 207 1571 211
rect 247 190 251 194
rect 335 190 339 194
rect 407 191 411 195
rect 423 190 427 194
rect 367 183 371 187
rect 583 143 587 147
rect 135 138 139 142
rect 223 138 227 142
rect 311 138 315 142
rect 239 127 243 131
rect 399 138 403 142
rect 327 127 331 131
rect 487 138 491 142
rect 415 127 419 131
rect 575 138 579 142
rect 503 127 507 131
rect 591 127 595 131
rect 111 121 115 125
rect 1567 121 1571 125
rect 111 103 115 107
rect 1567 103 1571 107
rect 135 92 139 96
rect 223 92 227 96
rect 239 91 243 95
rect 311 92 315 96
rect 327 91 331 95
rect 399 92 403 96
rect 415 91 419 95
rect 487 92 491 96
rect 503 91 507 95
rect 575 92 579 96
rect 591 91 595 95
<< m3 >>
rect 111 1522 115 1523
rect 111 1517 115 1518
rect 399 1522 403 1523
rect 399 1517 403 1518
rect 487 1522 491 1523
rect 487 1517 491 1518
rect 575 1522 579 1523
rect 575 1517 579 1518
rect 671 1522 675 1523
rect 671 1517 675 1518
rect 783 1522 787 1523
rect 783 1517 787 1518
rect 903 1522 907 1523
rect 903 1517 907 1518
rect 1031 1522 1035 1523
rect 1031 1517 1035 1518
rect 1167 1522 1171 1523
rect 1167 1517 1171 1518
rect 1303 1522 1307 1523
rect 1303 1517 1307 1518
rect 1447 1522 1451 1523
rect 1447 1517 1451 1518
rect 1567 1522 1571 1523
rect 1567 1517 1571 1518
rect 112 1494 114 1517
rect 400 1511 402 1517
rect 488 1511 490 1517
rect 576 1511 578 1517
rect 672 1511 674 1517
rect 784 1511 786 1517
rect 904 1511 906 1517
rect 1032 1511 1034 1517
rect 1168 1511 1170 1517
rect 1304 1511 1306 1517
rect 1448 1511 1450 1517
rect 398 1510 404 1511
rect 398 1506 399 1510
rect 403 1506 404 1510
rect 398 1505 404 1506
rect 486 1510 492 1511
rect 486 1506 487 1510
rect 491 1506 492 1510
rect 486 1505 492 1506
rect 574 1510 580 1511
rect 574 1506 575 1510
rect 579 1506 580 1510
rect 574 1505 580 1506
rect 670 1510 676 1511
rect 670 1506 671 1510
rect 675 1506 676 1510
rect 670 1505 676 1506
rect 782 1510 788 1511
rect 782 1506 783 1510
rect 787 1506 788 1510
rect 782 1505 788 1506
rect 902 1510 908 1511
rect 902 1506 903 1510
rect 907 1506 908 1510
rect 902 1505 908 1506
rect 1030 1510 1036 1511
rect 1030 1506 1031 1510
rect 1035 1506 1036 1510
rect 1030 1505 1036 1506
rect 1166 1510 1172 1511
rect 1166 1506 1167 1510
rect 1171 1506 1172 1510
rect 1302 1510 1308 1511
rect 1166 1505 1172 1506
rect 1210 1507 1216 1508
rect 1210 1503 1211 1507
rect 1215 1503 1216 1507
rect 1302 1506 1303 1510
rect 1307 1506 1308 1510
rect 1302 1505 1308 1506
rect 1446 1510 1452 1511
rect 1446 1506 1447 1510
rect 1451 1506 1452 1510
rect 1446 1505 1452 1506
rect 1210 1502 1216 1503
rect 502 1499 508 1500
rect 502 1495 503 1499
rect 507 1495 508 1499
rect 502 1494 508 1495
rect 590 1499 596 1500
rect 590 1495 591 1499
rect 595 1495 596 1499
rect 590 1494 596 1495
rect 686 1499 692 1500
rect 686 1495 687 1499
rect 691 1495 692 1499
rect 686 1494 692 1495
rect 798 1499 804 1500
rect 798 1495 799 1499
rect 803 1495 804 1499
rect 798 1494 804 1495
rect 918 1499 924 1500
rect 918 1495 919 1499
rect 923 1495 924 1499
rect 918 1494 924 1495
rect 1046 1499 1052 1500
rect 1046 1495 1047 1499
rect 1051 1495 1052 1499
rect 1046 1494 1052 1495
rect 1182 1499 1188 1500
rect 1182 1495 1183 1499
rect 1187 1495 1188 1499
rect 1182 1494 1188 1495
rect 110 1493 116 1494
rect 110 1489 111 1493
rect 115 1489 116 1493
rect 110 1488 116 1489
rect 110 1475 116 1476
rect 110 1471 111 1475
rect 115 1471 116 1475
rect 110 1470 116 1471
rect 112 1447 114 1470
rect 398 1464 404 1465
rect 486 1464 492 1465
rect 504 1464 506 1494
rect 574 1464 580 1465
rect 592 1464 594 1494
rect 670 1464 676 1465
rect 688 1464 690 1494
rect 782 1464 788 1465
rect 800 1464 802 1494
rect 902 1464 908 1465
rect 920 1464 922 1494
rect 1030 1464 1036 1465
rect 1048 1464 1050 1494
rect 1166 1464 1172 1465
rect 1184 1464 1186 1494
rect 398 1460 399 1464
rect 403 1460 404 1464
rect 398 1459 404 1460
rect 466 1463 472 1464
rect 466 1459 467 1463
rect 471 1459 472 1463
rect 486 1460 487 1464
rect 491 1460 492 1464
rect 486 1459 492 1460
rect 502 1463 508 1464
rect 502 1459 503 1463
rect 507 1459 508 1463
rect 574 1460 575 1464
rect 579 1460 580 1464
rect 574 1459 580 1460
rect 590 1463 596 1464
rect 590 1459 591 1463
rect 595 1459 596 1463
rect 670 1460 671 1464
rect 675 1460 676 1464
rect 670 1459 676 1460
rect 686 1463 692 1464
rect 686 1459 687 1463
rect 691 1459 692 1463
rect 782 1460 783 1464
rect 787 1460 788 1464
rect 782 1459 788 1460
rect 798 1463 804 1464
rect 798 1459 799 1463
rect 803 1459 804 1463
rect 902 1460 903 1464
rect 907 1460 908 1464
rect 902 1459 908 1460
rect 918 1463 924 1464
rect 918 1459 919 1463
rect 923 1459 924 1463
rect 1030 1460 1031 1464
rect 1035 1460 1036 1464
rect 1030 1459 1036 1460
rect 1046 1463 1052 1464
rect 1046 1459 1047 1463
rect 1051 1459 1052 1463
rect 1166 1460 1167 1464
rect 1171 1460 1172 1464
rect 1166 1459 1172 1460
rect 1182 1463 1188 1464
rect 1182 1459 1183 1463
rect 1187 1459 1188 1463
rect 400 1447 402 1459
rect 466 1458 472 1459
rect 111 1446 115 1447
rect 111 1441 115 1442
rect 399 1446 403 1447
rect 399 1441 403 1442
rect 423 1446 427 1447
rect 423 1441 427 1442
rect 112 1430 114 1441
rect 422 1440 428 1441
rect 422 1436 423 1440
rect 427 1436 428 1440
rect 422 1435 428 1436
rect 110 1429 116 1430
rect 110 1425 111 1429
rect 115 1425 116 1429
rect 110 1424 116 1425
rect 110 1411 116 1412
rect 110 1407 111 1411
rect 115 1407 116 1411
rect 110 1406 116 1407
rect 112 1379 114 1406
rect 468 1396 470 1458
rect 488 1447 490 1459
rect 502 1458 508 1459
rect 576 1447 578 1459
rect 590 1458 596 1459
rect 672 1447 674 1459
rect 686 1458 692 1459
rect 784 1447 786 1459
rect 798 1458 804 1459
rect 904 1447 906 1459
rect 918 1458 924 1459
rect 1032 1447 1034 1459
rect 1046 1458 1052 1459
rect 1168 1447 1170 1459
rect 1182 1458 1188 1459
rect 487 1446 491 1447
rect 487 1441 491 1442
rect 575 1446 579 1447
rect 575 1441 579 1442
rect 655 1446 659 1447
rect 655 1441 659 1442
rect 671 1446 675 1447
rect 671 1441 675 1442
rect 783 1446 787 1447
rect 783 1441 787 1442
rect 895 1446 899 1447
rect 895 1441 899 1442
rect 903 1446 907 1447
rect 903 1441 907 1442
rect 1031 1446 1035 1447
rect 1031 1441 1035 1442
rect 1143 1446 1147 1447
rect 1143 1441 1147 1442
rect 1167 1446 1171 1447
rect 1167 1441 1171 1442
rect 654 1440 660 1441
rect 894 1440 900 1441
rect 1142 1440 1148 1441
rect 1212 1440 1214 1502
rect 1414 1499 1420 1500
rect 1414 1495 1415 1499
rect 1419 1495 1420 1499
rect 1414 1494 1420 1495
rect 1568 1494 1570 1517
rect 1302 1464 1308 1465
rect 1416 1464 1418 1494
rect 1566 1493 1572 1494
rect 1566 1489 1567 1493
rect 1571 1489 1572 1493
rect 1566 1488 1572 1489
rect 1566 1475 1572 1476
rect 1566 1471 1567 1475
rect 1571 1471 1572 1475
rect 1566 1470 1572 1471
rect 1446 1464 1452 1465
rect 1302 1460 1303 1464
rect 1307 1460 1308 1464
rect 1302 1459 1308 1460
rect 1414 1463 1420 1464
rect 1414 1459 1415 1463
rect 1419 1459 1420 1463
rect 1446 1460 1447 1464
rect 1451 1460 1452 1464
rect 1446 1459 1452 1460
rect 1478 1463 1484 1464
rect 1478 1459 1479 1463
rect 1483 1459 1484 1463
rect 1304 1447 1306 1459
rect 1414 1458 1420 1459
rect 1448 1447 1450 1459
rect 1478 1458 1484 1459
rect 1303 1446 1307 1447
rect 1303 1441 1307 1442
rect 1399 1446 1403 1447
rect 1399 1441 1403 1442
rect 1447 1446 1451 1447
rect 1447 1441 1451 1442
rect 1398 1440 1404 1441
rect 654 1436 655 1440
rect 659 1436 660 1440
rect 654 1435 660 1436
rect 722 1439 728 1440
rect 722 1435 723 1439
rect 727 1435 728 1439
rect 894 1436 895 1440
rect 899 1436 900 1440
rect 894 1435 900 1436
rect 910 1439 916 1440
rect 910 1435 911 1439
rect 915 1435 916 1439
rect 1142 1436 1143 1440
rect 1147 1436 1148 1440
rect 1142 1435 1148 1436
rect 1210 1439 1216 1440
rect 1210 1435 1211 1439
rect 1215 1435 1216 1439
rect 1398 1436 1399 1440
rect 1403 1436 1404 1440
rect 1398 1435 1404 1436
rect 1438 1439 1444 1440
rect 1438 1435 1439 1439
rect 1443 1435 1444 1439
rect 722 1434 728 1435
rect 910 1434 916 1435
rect 1210 1434 1216 1435
rect 1438 1434 1444 1435
rect 466 1395 472 1396
rect 422 1394 428 1395
rect 422 1390 423 1394
rect 427 1390 428 1394
rect 466 1391 467 1395
rect 471 1391 472 1395
rect 466 1390 472 1391
rect 654 1394 660 1395
rect 654 1390 655 1394
rect 659 1390 660 1394
rect 422 1389 428 1390
rect 654 1389 660 1390
rect 424 1379 426 1389
rect 656 1379 658 1389
rect 724 1388 726 1434
rect 894 1394 900 1395
rect 894 1390 895 1394
rect 899 1390 900 1394
rect 894 1389 900 1390
rect 722 1387 728 1388
rect 722 1383 723 1387
rect 727 1383 728 1387
rect 722 1382 728 1383
rect 896 1379 898 1389
rect 111 1378 115 1379
rect 111 1373 115 1374
rect 423 1378 427 1379
rect 423 1373 427 1374
rect 471 1378 475 1379
rect 471 1373 475 1374
rect 655 1378 659 1379
rect 655 1373 659 1374
rect 695 1378 699 1379
rect 695 1373 699 1374
rect 895 1378 899 1379
rect 895 1373 899 1374
rect 112 1350 114 1373
rect 472 1367 474 1373
rect 696 1367 698 1373
rect 912 1372 914 1434
rect 1142 1394 1148 1395
rect 1142 1390 1143 1394
rect 1147 1390 1148 1394
rect 1142 1389 1148 1390
rect 1398 1394 1404 1395
rect 1398 1390 1399 1394
rect 1403 1390 1404 1394
rect 1398 1389 1404 1390
rect 1144 1379 1146 1389
rect 1190 1387 1196 1388
rect 1190 1383 1191 1387
rect 1195 1383 1196 1387
rect 1190 1382 1196 1383
rect 919 1378 923 1379
rect 919 1373 923 1374
rect 1143 1378 1147 1379
rect 1143 1373 1147 1374
rect 1151 1378 1155 1379
rect 1151 1373 1155 1374
rect 910 1371 916 1372
rect 910 1367 911 1371
rect 915 1367 916 1371
rect 920 1367 922 1373
rect 1152 1367 1154 1373
rect 470 1366 476 1367
rect 470 1362 471 1366
rect 475 1362 476 1366
rect 470 1361 476 1362
rect 694 1366 700 1367
rect 910 1366 916 1367
rect 918 1366 924 1367
rect 694 1362 695 1366
rect 699 1362 700 1366
rect 694 1361 700 1362
rect 918 1362 919 1366
rect 923 1362 924 1366
rect 1150 1366 1156 1367
rect 918 1361 924 1362
rect 1006 1363 1012 1364
rect 1006 1359 1007 1363
rect 1011 1359 1012 1363
rect 1150 1362 1151 1366
rect 1155 1362 1156 1366
rect 1150 1361 1156 1362
rect 1006 1358 1012 1359
rect 710 1355 716 1356
rect 710 1351 711 1355
rect 715 1351 716 1355
rect 710 1350 716 1351
rect 110 1349 116 1350
rect 110 1345 111 1349
rect 115 1345 116 1349
rect 110 1344 116 1345
rect 110 1331 116 1332
rect 110 1327 111 1331
rect 115 1327 116 1331
rect 110 1326 116 1327
rect 112 1307 114 1326
rect 470 1320 476 1321
rect 470 1316 471 1320
rect 475 1316 476 1320
rect 470 1315 476 1316
rect 694 1320 700 1321
rect 712 1320 714 1350
rect 918 1320 924 1321
rect 694 1316 695 1320
rect 699 1316 700 1320
rect 694 1315 700 1316
rect 710 1319 716 1320
rect 710 1315 711 1319
rect 715 1315 716 1319
rect 918 1316 919 1320
rect 923 1316 924 1320
rect 918 1315 924 1316
rect 472 1307 474 1315
rect 696 1307 698 1315
rect 710 1314 716 1315
rect 920 1307 922 1315
rect 111 1306 115 1307
rect 111 1301 115 1302
rect 471 1306 475 1307
rect 471 1301 475 1302
rect 519 1306 523 1307
rect 519 1301 523 1302
rect 695 1306 699 1307
rect 695 1301 699 1302
rect 743 1306 747 1307
rect 743 1301 747 1302
rect 919 1306 923 1307
rect 919 1301 923 1302
rect 975 1306 979 1307
rect 975 1301 979 1302
rect 112 1290 114 1301
rect 518 1300 524 1301
rect 742 1300 748 1301
rect 974 1300 980 1301
rect 1008 1300 1010 1358
rect 1150 1320 1156 1321
rect 1192 1320 1194 1382
rect 1400 1379 1402 1389
rect 1391 1378 1395 1379
rect 1391 1373 1395 1374
rect 1399 1378 1403 1379
rect 1399 1373 1403 1374
rect 1392 1367 1394 1373
rect 1440 1372 1442 1434
rect 1480 1396 1482 1458
rect 1568 1447 1570 1470
rect 1567 1446 1571 1447
rect 1567 1441 1571 1442
rect 1568 1430 1570 1441
rect 1566 1429 1572 1430
rect 1566 1425 1567 1429
rect 1571 1425 1572 1429
rect 1566 1424 1572 1425
rect 1566 1411 1572 1412
rect 1566 1407 1567 1411
rect 1571 1407 1572 1411
rect 1566 1406 1572 1407
rect 1478 1395 1484 1396
rect 1478 1391 1479 1395
rect 1483 1391 1484 1395
rect 1478 1390 1484 1391
rect 1568 1379 1570 1406
rect 1567 1378 1571 1379
rect 1567 1373 1571 1374
rect 1438 1371 1444 1372
rect 1438 1367 1439 1371
rect 1443 1367 1444 1371
rect 1390 1366 1396 1367
rect 1438 1366 1444 1367
rect 1390 1362 1391 1366
rect 1395 1362 1396 1366
rect 1390 1361 1396 1362
rect 1568 1350 1570 1373
rect 1566 1349 1572 1350
rect 1566 1345 1567 1349
rect 1571 1345 1572 1349
rect 1566 1344 1572 1345
rect 1566 1331 1572 1332
rect 1566 1327 1567 1331
rect 1571 1327 1572 1331
rect 1566 1326 1572 1327
rect 1390 1320 1396 1321
rect 1150 1316 1151 1320
rect 1155 1316 1156 1320
rect 1150 1315 1156 1316
rect 1190 1319 1196 1320
rect 1190 1315 1191 1319
rect 1195 1315 1196 1319
rect 1390 1316 1391 1320
rect 1395 1316 1396 1320
rect 1390 1315 1396 1316
rect 1422 1319 1428 1320
rect 1422 1315 1423 1319
rect 1427 1315 1428 1319
rect 1152 1307 1154 1315
rect 1190 1314 1196 1315
rect 1392 1307 1394 1315
rect 1422 1314 1428 1315
rect 1151 1306 1155 1307
rect 1151 1301 1155 1302
rect 1207 1306 1211 1307
rect 1207 1301 1211 1302
rect 1391 1306 1395 1307
rect 1391 1301 1395 1302
rect 1206 1300 1212 1301
rect 518 1296 519 1300
rect 523 1296 524 1300
rect 518 1295 524 1296
rect 586 1299 592 1300
rect 586 1295 587 1299
rect 591 1295 592 1299
rect 742 1296 743 1300
rect 747 1296 748 1300
rect 742 1295 748 1296
rect 810 1299 816 1300
rect 810 1295 811 1299
rect 815 1295 816 1299
rect 974 1296 975 1300
rect 979 1296 980 1300
rect 974 1295 980 1296
rect 1006 1299 1012 1300
rect 1006 1295 1007 1299
rect 1011 1295 1012 1299
rect 1206 1296 1207 1300
rect 1211 1296 1212 1300
rect 1206 1295 1212 1296
rect 1274 1299 1280 1300
rect 1274 1295 1275 1299
rect 1279 1295 1280 1299
rect 586 1294 592 1295
rect 810 1294 816 1295
rect 1006 1294 1012 1295
rect 1274 1294 1280 1295
rect 110 1289 116 1290
rect 110 1285 111 1289
rect 115 1285 116 1289
rect 110 1284 116 1285
rect 110 1271 116 1272
rect 110 1267 111 1271
rect 115 1267 116 1271
rect 110 1266 116 1267
rect 112 1227 114 1266
rect 518 1254 524 1255
rect 518 1250 519 1254
rect 523 1250 524 1254
rect 518 1249 524 1250
rect 520 1227 522 1249
rect 588 1248 590 1294
rect 742 1254 748 1255
rect 742 1250 743 1254
rect 747 1250 748 1254
rect 742 1249 748 1250
rect 586 1247 592 1248
rect 586 1243 587 1247
rect 591 1243 592 1247
rect 586 1242 592 1243
rect 744 1227 746 1249
rect 111 1226 115 1227
rect 111 1221 115 1222
rect 519 1226 523 1227
rect 519 1221 523 1222
rect 567 1226 571 1227
rect 567 1221 571 1222
rect 743 1226 747 1227
rect 743 1221 747 1222
rect 767 1226 771 1227
rect 812 1224 814 1294
rect 974 1254 980 1255
rect 974 1250 975 1254
rect 979 1250 980 1254
rect 974 1249 980 1250
rect 1206 1254 1212 1255
rect 1206 1250 1207 1254
rect 1211 1250 1212 1254
rect 1206 1249 1212 1250
rect 976 1227 978 1249
rect 1190 1247 1196 1248
rect 1190 1243 1191 1247
rect 1195 1243 1196 1247
rect 1190 1242 1196 1243
rect 967 1226 971 1227
rect 767 1221 771 1222
rect 810 1223 816 1224
rect 112 1198 114 1221
rect 568 1215 570 1221
rect 768 1215 770 1221
rect 810 1219 811 1223
rect 815 1219 816 1223
rect 967 1221 971 1222
rect 975 1226 979 1227
rect 975 1221 979 1222
rect 1175 1226 1179 1227
rect 1175 1221 1179 1222
rect 810 1218 816 1219
rect 968 1215 970 1221
rect 1176 1215 1178 1221
rect 566 1214 572 1215
rect 566 1210 567 1214
rect 571 1210 572 1214
rect 566 1209 572 1210
rect 766 1214 772 1215
rect 766 1210 767 1214
rect 771 1210 772 1214
rect 766 1209 772 1210
rect 966 1214 972 1215
rect 966 1210 967 1214
rect 971 1210 972 1214
rect 966 1209 972 1210
rect 1174 1214 1180 1215
rect 1174 1210 1175 1214
rect 1179 1210 1180 1214
rect 1174 1209 1180 1210
rect 782 1203 788 1204
rect 782 1199 783 1203
rect 787 1199 788 1203
rect 782 1198 788 1199
rect 982 1203 988 1204
rect 982 1199 983 1203
rect 987 1199 988 1203
rect 982 1198 988 1199
rect 110 1197 116 1198
rect 110 1193 111 1197
rect 115 1193 116 1197
rect 110 1192 116 1193
rect 110 1179 116 1180
rect 110 1175 111 1179
rect 115 1175 116 1179
rect 110 1174 116 1175
rect 112 1163 114 1174
rect 566 1168 572 1169
rect 766 1168 772 1169
rect 784 1168 786 1198
rect 966 1168 972 1169
rect 984 1168 986 1198
rect 1174 1168 1180 1169
rect 1192 1168 1194 1242
rect 1208 1227 1210 1249
rect 1276 1248 1278 1294
rect 1424 1256 1426 1314
rect 1568 1307 1570 1326
rect 1439 1306 1443 1307
rect 1439 1301 1443 1302
rect 1567 1306 1571 1307
rect 1567 1301 1571 1302
rect 1438 1300 1444 1301
rect 1438 1296 1439 1300
rect 1443 1296 1444 1300
rect 1438 1295 1444 1296
rect 1470 1299 1476 1300
rect 1470 1295 1471 1299
rect 1475 1295 1476 1299
rect 1470 1294 1476 1295
rect 1422 1255 1428 1256
rect 1422 1251 1423 1255
rect 1427 1251 1428 1255
rect 1422 1250 1428 1251
rect 1438 1254 1444 1255
rect 1438 1250 1439 1254
rect 1443 1250 1444 1254
rect 1438 1249 1444 1250
rect 1274 1247 1280 1248
rect 1274 1243 1275 1247
rect 1279 1243 1280 1247
rect 1274 1242 1280 1243
rect 1440 1227 1442 1249
rect 1207 1226 1211 1227
rect 1207 1221 1211 1222
rect 1391 1226 1395 1227
rect 1391 1221 1395 1222
rect 1439 1226 1443 1227
rect 1439 1221 1443 1222
rect 1392 1215 1394 1221
rect 1472 1220 1474 1294
rect 1568 1290 1570 1301
rect 1566 1289 1572 1290
rect 1566 1285 1567 1289
rect 1571 1285 1572 1289
rect 1566 1284 1572 1285
rect 1566 1271 1572 1272
rect 1566 1267 1567 1271
rect 1571 1267 1572 1271
rect 1566 1266 1572 1267
rect 1568 1227 1570 1266
rect 1567 1226 1571 1227
rect 1567 1221 1571 1222
rect 1470 1219 1476 1220
rect 1470 1215 1471 1219
rect 1475 1215 1476 1219
rect 1390 1214 1396 1215
rect 1470 1214 1476 1215
rect 1254 1211 1260 1212
rect 1254 1207 1255 1211
rect 1259 1207 1260 1211
rect 1390 1210 1391 1214
rect 1395 1210 1396 1214
rect 1390 1209 1396 1210
rect 1254 1206 1260 1207
rect 566 1164 567 1168
rect 571 1164 572 1168
rect 566 1163 572 1164
rect 726 1167 732 1168
rect 726 1163 727 1167
rect 731 1163 732 1167
rect 766 1164 767 1168
rect 771 1164 772 1168
rect 766 1163 772 1164
rect 782 1167 788 1168
rect 782 1163 783 1167
rect 787 1163 788 1167
rect 966 1164 967 1168
rect 971 1164 972 1168
rect 966 1163 972 1164
rect 982 1167 988 1168
rect 982 1163 983 1167
rect 987 1163 988 1167
rect 1174 1164 1175 1168
rect 1179 1164 1180 1168
rect 1174 1163 1180 1164
rect 1190 1167 1196 1168
rect 1190 1163 1191 1167
rect 1195 1163 1196 1167
rect 111 1162 115 1163
rect 111 1157 115 1158
rect 567 1162 571 1163
rect 567 1157 571 1158
rect 703 1162 707 1163
rect 726 1162 732 1163
rect 767 1162 771 1163
rect 782 1162 788 1163
rect 967 1162 971 1163
rect 982 1162 988 1163
rect 1055 1162 1059 1163
rect 703 1157 707 1158
rect 112 1146 114 1157
rect 702 1156 708 1157
rect 702 1152 703 1156
rect 707 1152 708 1156
rect 702 1151 708 1152
rect 110 1145 116 1146
rect 110 1141 111 1145
rect 115 1141 116 1145
rect 110 1140 116 1141
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 110 1122 116 1123
rect 112 1099 114 1122
rect 728 1112 730 1162
rect 767 1157 771 1158
rect 967 1157 971 1158
rect 1055 1157 1059 1158
rect 1175 1162 1179 1163
rect 1190 1162 1196 1163
rect 1175 1157 1179 1158
rect 1054 1156 1060 1157
rect 978 1155 984 1156
rect 978 1151 979 1155
rect 983 1151 984 1155
rect 1054 1152 1055 1156
rect 1059 1152 1060 1156
rect 1054 1151 1060 1152
rect 1078 1155 1084 1156
rect 1078 1151 1079 1155
rect 1083 1151 1084 1155
rect 978 1150 984 1151
rect 1078 1150 1084 1151
rect 726 1111 732 1112
rect 702 1110 708 1111
rect 702 1106 703 1110
rect 707 1106 708 1110
rect 726 1107 727 1111
rect 731 1107 732 1111
rect 726 1106 732 1107
rect 702 1105 708 1106
rect 704 1099 706 1105
rect 980 1104 982 1150
rect 1054 1110 1060 1111
rect 1054 1106 1055 1110
rect 1059 1106 1060 1110
rect 1054 1105 1060 1106
rect 978 1103 984 1104
rect 978 1099 979 1103
rect 983 1099 984 1103
rect 1056 1099 1058 1105
rect 111 1098 115 1099
rect 111 1093 115 1094
rect 671 1098 675 1099
rect 671 1093 675 1094
rect 703 1098 707 1099
rect 703 1093 707 1094
rect 847 1098 851 1099
rect 978 1098 984 1099
rect 1031 1098 1035 1099
rect 847 1093 851 1094
rect 1031 1093 1035 1094
rect 1055 1098 1059 1099
rect 1055 1093 1059 1094
rect 112 1070 114 1093
rect 672 1087 674 1093
rect 848 1087 850 1093
rect 1032 1087 1034 1093
rect 1080 1092 1082 1150
rect 1223 1098 1227 1099
rect 1223 1093 1227 1094
rect 1078 1091 1084 1092
rect 1078 1087 1079 1091
rect 1083 1087 1084 1091
rect 1224 1087 1226 1093
rect 670 1086 676 1087
rect 670 1082 671 1086
rect 675 1082 676 1086
rect 670 1081 676 1082
rect 846 1086 852 1087
rect 846 1082 847 1086
rect 851 1082 852 1086
rect 846 1081 852 1082
rect 1030 1086 1036 1087
rect 1078 1086 1084 1087
rect 1222 1086 1228 1087
rect 1030 1082 1031 1086
rect 1035 1082 1036 1086
rect 1030 1081 1036 1082
rect 1222 1082 1223 1086
rect 1227 1082 1228 1086
rect 1222 1081 1228 1082
rect 862 1075 868 1076
rect 862 1071 863 1075
rect 867 1071 868 1075
rect 862 1070 868 1071
rect 1046 1075 1052 1076
rect 1046 1071 1047 1075
rect 1051 1071 1052 1075
rect 1046 1070 1052 1071
rect 110 1069 116 1070
rect 110 1065 111 1069
rect 115 1065 116 1069
rect 110 1064 116 1065
rect 110 1051 116 1052
rect 110 1047 111 1051
rect 115 1047 116 1051
rect 110 1046 116 1047
rect 112 1019 114 1046
rect 670 1040 676 1041
rect 670 1036 671 1040
rect 675 1036 676 1040
rect 670 1035 676 1036
rect 846 1040 852 1041
rect 864 1040 866 1070
rect 1030 1040 1036 1041
rect 1048 1040 1050 1070
rect 1222 1040 1228 1041
rect 1256 1040 1258 1206
rect 1568 1198 1570 1221
rect 1566 1197 1572 1198
rect 1566 1193 1567 1197
rect 1571 1193 1572 1197
rect 1566 1192 1572 1193
rect 1566 1179 1572 1180
rect 1566 1175 1567 1179
rect 1571 1175 1572 1179
rect 1566 1174 1572 1175
rect 1390 1168 1396 1169
rect 1390 1164 1391 1168
rect 1395 1164 1396 1168
rect 1390 1163 1396 1164
rect 1454 1167 1460 1168
rect 1454 1163 1455 1167
rect 1459 1163 1460 1167
rect 1568 1163 1570 1174
rect 1391 1162 1395 1163
rect 1391 1157 1395 1158
rect 1407 1162 1411 1163
rect 1454 1162 1460 1163
rect 1567 1162 1571 1163
rect 1407 1157 1411 1158
rect 1406 1156 1412 1157
rect 1406 1152 1407 1156
rect 1411 1152 1412 1156
rect 1406 1151 1412 1152
rect 1456 1112 1458 1162
rect 1567 1157 1571 1158
rect 1462 1155 1468 1156
rect 1462 1151 1463 1155
rect 1467 1151 1468 1155
rect 1462 1150 1468 1151
rect 1454 1111 1460 1112
rect 1406 1110 1412 1111
rect 1406 1106 1407 1110
rect 1411 1106 1412 1110
rect 1454 1107 1455 1111
rect 1459 1107 1460 1111
rect 1454 1106 1460 1107
rect 1406 1105 1412 1106
rect 1408 1099 1410 1105
rect 1407 1098 1411 1099
rect 1407 1093 1411 1094
rect 1415 1098 1419 1099
rect 1415 1093 1419 1094
rect 1416 1087 1418 1093
rect 1464 1092 1466 1150
rect 1568 1146 1570 1157
rect 1566 1145 1572 1146
rect 1566 1141 1567 1145
rect 1571 1141 1572 1145
rect 1566 1140 1572 1141
rect 1566 1127 1572 1128
rect 1566 1123 1567 1127
rect 1571 1123 1572 1127
rect 1566 1122 1572 1123
rect 1568 1099 1570 1122
rect 1567 1098 1571 1099
rect 1567 1093 1571 1094
rect 1462 1091 1468 1092
rect 1462 1087 1463 1091
rect 1467 1087 1468 1091
rect 1414 1086 1420 1087
rect 1462 1086 1468 1087
rect 1266 1083 1272 1084
rect 1266 1079 1267 1083
rect 1271 1079 1272 1083
rect 1414 1082 1415 1086
rect 1419 1082 1420 1086
rect 1414 1081 1420 1082
rect 1266 1078 1272 1079
rect 846 1036 847 1040
rect 851 1036 852 1040
rect 846 1035 852 1036
rect 862 1039 868 1040
rect 862 1035 863 1039
rect 867 1035 868 1039
rect 1030 1036 1031 1040
rect 1035 1036 1036 1040
rect 1030 1035 1036 1036
rect 1046 1039 1052 1040
rect 1046 1035 1047 1039
rect 1051 1035 1052 1039
rect 1222 1036 1223 1040
rect 1227 1036 1228 1040
rect 1222 1035 1228 1036
rect 1254 1039 1260 1040
rect 1254 1035 1255 1039
rect 1259 1035 1260 1039
rect 672 1019 674 1035
rect 848 1019 850 1035
rect 862 1034 868 1035
rect 1006 1031 1012 1032
rect 1006 1027 1007 1031
rect 1011 1027 1012 1031
rect 1006 1026 1012 1027
rect 111 1018 115 1019
rect 111 1013 115 1014
rect 575 1018 579 1019
rect 575 1013 579 1014
rect 671 1018 675 1019
rect 671 1013 675 1014
rect 775 1018 779 1019
rect 775 1013 779 1014
rect 847 1018 851 1019
rect 847 1013 851 1014
rect 983 1018 987 1019
rect 983 1013 987 1014
rect 112 1002 114 1013
rect 574 1012 580 1013
rect 774 1012 780 1013
rect 982 1012 988 1013
rect 574 1008 575 1012
rect 579 1008 580 1012
rect 574 1007 580 1008
rect 606 1011 612 1012
rect 606 1007 607 1011
rect 611 1007 612 1011
rect 774 1008 775 1012
rect 779 1008 780 1012
rect 774 1007 780 1008
rect 806 1011 812 1012
rect 806 1007 807 1011
rect 811 1007 812 1011
rect 982 1008 983 1012
rect 987 1008 988 1012
rect 982 1007 988 1008
rect 606 1006 612 1007
rect 806 1006 812 1007
rect 110 1001 116 1002
rect 110 997 111 1001
rect 115 997 116 1001
rect 110 996 116 997
rect 110 983 116 984
rect 110 979 111 983
rect 115 979 116 983
rect 110 978 116 979
rect 112 947 114 978
rect 574 966 580 967
rect 574 962 575 966
rect 579 962 580 966
rect 574 961 580 962
rect 576 947 578 961
rect 111 946 115 947
rect 111 941 115 942
rect 407 946 411 947
rect 407 941 411 942
rect 575 946 579 947
rect 575 941 579 942
rect 112 918 114 941
rect 408 935 410 941
rect 608 940 610 1006
rect 774 966 780 967
rect 774 962 775 966
rect 779 962 780 966
rect 774 961 780 962
rect 776 947 778 961
rect 808 960 810 1006
rect 1008 968 1010 1026
rect 1032 1019 1034 1035
rect 1046 1034 1052 1035
rect 1224 1019 1226 1035
rect 1254 1034 1260 1035
rect 1031 1018 1035 1019
rect 1031 1013 1035 1014
rect 1191 1018 1195 1019
rect 1191 1013 1195 1014
rect 1223 1018 1227 1019
rect 1223 1013 1227 1014
rect 1190 1012 1196 1013
rect 1268 1012 1270 1078
rect 1568 1070 1570 1093
rect 1566 1069 1572 1070
rect 1566 1065 1567 1069
rect 1571 1065 1572 1069
rect 1566 1064 1572 1065
rect 1566 1051 1572 1052
rect 1566 1047 1567 1051
rect 1571 1047 1572 1051
rect 1566 1046 1572 1047
rect 1414 1040 1420 1041
rect 1414 1036 1415 1040
rect 1419 1036 1420 1040
rect 1414 1035 1420 1036
rect 1454 1039 1460 1040
rect 1454 1035 1455 1039
rect 1459 1035 1460 1039
rect 1416 1019 1418 1035
rect 1454 1034 1460 1035
rect 1407 1018 1411 1019
rect 1407 1013 1411 1014
rect 1415 1018 1419 1019
rect 1415 1013 1419 1014
rect 1406 1012 1412 1013
rect 1014 1011 1020 1012
rect 1014 1007 1015 1011
rect 1019 1007 1020 1011
rect 1190 1008 1191 1012
rect 1195 1008 1196 1012
rect 1190 1007 1196 1008
rect 1266 1011 1272 1012
rect 1266 1007 1267 1011
rect 1271 1007 1272 1011
rect 1406 1008 1407 1012
rect 1411 1008 1412 1012
rect 1406 1007 1412 1008
rect 1446 1011 1452 1012
rect 1446 1007 1447 1011
rect 1451 1007 1452 1011
rect 1014 1006 1020 1007
rect 1266 1006 1272 1007
rect 1446 1006 1452 1007
rect 1006 967 1012 968
rect 982 966 988 967
rect 982 962 983 966
rect 987 962 988 966
rect 1006 963 1007 967
rect 1011 963 1012 967
rect 1006 962 1012 963
rect 982 961 988 962
rect 806 959 812 960
rect 806 955 807 959
rect 811 955 812 959
rect 806 954 812 955
rect 984 947 986 961
rect 1016 960 1018 1006
rect 1190 966 1196 967
rect 1190 962 1191 966
rect 1195 962 1196 966
rect 1190 961 1196 962
rect 1406 966 1412 967
rect 1406 962 1407 966
rect 1411 962 1412 966
rect 1406 961 1412 962
rect 1014 959 1020 960
rect 1014 955 1015 959
rect 1019 955 1020 959
rect 1014 954 1020 955
rect 1162 959 1168 960
rect 1162 955 1163 959
rect 1167 955 1168 959
rect 1162 954 1168 955
rect 735 946 739 947
rect 735 941 739 942
rect 775 946 779 947
rect 775 941 779 942
rect 983 946 987 947
rect 983 941 987 942
rect 1063 946 1067 947
rect 1063 941 1067 942
rect 606 939 612 940
rect 606 935 607 939
rect 611 935 612 939
rect 736 935 738 941
rect 1064 935 1066 941
rect 406 934 412 935
rect 606 934 612 935
rect 734 934 740 935
rect 406 930 407 934
rect 411 930 412 934
rect 406 929 412 930
rect 734 930 735 934
rect 739 930 740 934
rect 734 929 740 930
rect 1062 934 1068 935
rect 1062 930 1063 934
rect 1067 930 1068 934
rect 1062 929 1068 930
rect 610 923 616 924
rect 610 919 611 923
rect 615 919 616 923
rect 610 918 616 919
rect 930 923 936 924
rect 930 919 931 923
rect 935 919 936 923
rect 930 918 936 919
rect 110 917 116 918
rect 110 913 111 917
rect 115 913 116 917
rect 110 912 116 913
rect 110 899 116 900
rect 110 895 111 899
rect 115 895 116 899
rect 110 894 116 895
rect 112 879 114 894
rect 406 888 412 889
rect 612 888 614 918
rect 734 888 740 889
rect 932 888 934 918
rect 1062 888 1068 889
rect 406 884 407 888
rect 411 884 412 888
rect 406 883 412 884
rect 610 887 616 888
rect 610 883 611 887
rect 615 883 616 887
rect 734 884 735 888
rect 739 884 740 888
rect 734 883 740 884
rect 930 887 936 888
rect 930 883 931 887
rect 935 883 936 887
rect 1062 884 1063 888
rect 1067 884 1068 888
rect 1062 883 1068 884
rect 1078 887 1084 888
rect 1078 883 1079 887
rect 1083 883 1084 887
rect 408 879 410 883
rect 610 882 616 883
rect 736 879 738 883
rect 930 882 936 883
rect 1064 879 1066 883
rect 1078 882 1084 883
rect 111 878 115 879
rect 111 873 115 874
rect 255 878 259 879
rect 255 873 259 874
rect 407 878 411 879
rect 407 873 411 874
rect 527 878 531 879
rect 527 873 531 874
rect 735 878 739 879
rect 735 873 739 874
rect 807 878 811 879
rect 807 873 811 874
rect 1063 878 1067 879
rect 1063 873 1067 874
rect 112 862 114 873
rect 254 872 260 873
rect 526 872 532 873
rect 806 872 812 873
rect 254 868 255 872
rect 259 868 260 872
rect 254 867 260 868
rect 286 871 292 872
rect 286 867 287 871
rect 291 867 292 871
rect 526 868 527 872
rect 531 868 532 872
rect 526 867 532 868
rect 558 871 564 872
rect 558 867 559 871
rect 563 867 564 871
rect 806 868 807 872
rect 811 868 812 872
rect 806 867 812 868
rect 838 871 844 872
rect 838 867 839 871
rect 843 867 844 871
rect 286 866 292 867
rect 558 866 564 867
rect 838 866 844 867
rect 110 861 116 862
rect 110 857 111 861
rect 115 857 116 861
rect 110 856 116 857
rect 110 843 116 844
rect 110 839 111 843
rect 115 839 116 843
rect 110 838 116 839
rect 112 795 114 838
rect 254 826 260 827
rect 254 822 255 826
rect 259 822 260 826
rect 254 821 260 822
rect 256 795 258 821
rect 111 794 115 795
rect 111 789 115 790
rect 167 794 171 795
rect 167 789 171 790
rect 255 794 259 795
rect 255 789 259 790
rect 112 766 114 789
rect 168 783 170 789
rect 288 788 290 866
rect 526 826 532 827
rect 526 822 527 826
rect 531 822 532 826
rect 526 821 532 822
rect 528 795 530 821
rect 560 820 562 866
rect 806 826 812 827
rect 806 822 807 826
rect 811 822 812 826
rect 806 821 812 822
rect 558 819 564 820
rect 558 815 559 819
rect 563 815 564 819
rect 558 814 564 815
rect 808 795 810 821
rect 840 820 842 866
rect 1080 828 1082 882
rect 1095 878 1099 879
rect 1095 873 1099 874
rect 1094 872 1100 873
rect 1164 872 1166 954
rect 1192 947 1194 961
rect 1408 947 1410 961
rect 1191 946 1195 947
rect 1191 941 1195 942
rect 1399 946 1403 947
rect 1399 941 1403 942
rect 1407 946 1411 947
rect 1407 941 1411 942
rect 1400 935 1402 941
rect 1448 940 1450 1006
rect 1456 968 1458 1034
rect 1568 1019 1570 1046
rect 1567 1018 1571 1019
rect 1567 1013 1571 1014
rect 1568 1002 1570 1013
rect 1566 1001 1572 1002
rect 1566 997 1567 1001
rect 1571 997 1572 1001
rect 1566 996 1572 997
rect 1566 983 1572 984
rect 1566 979 1567 983
rect 1571 979 1572 983
rect 1566 978 1572 979
rect 1454 967 1460 968
rect 1454 963 1455 967
rect 1459 963 1460 967
rect 1454 962 1460 963
rect 1568 947 1570 978
rect 1567 946 1571 947
rect 1567 941 1571 942
rect 1446 939 1452 940
rect 1446 935 1447 939
rect 1451 935 1452 939
rect 1398 934 1404 935
rect 1446 934 1452 935
rect 1398 930 1399 934
rect 1403 930 1404 934
rect 1398 929 1404 930
rect 1568 918 1570 941
rect 1566 917 1572 918
rect 1566 913 1567 917
rect 1571 913 1572 917
rect 1566 912 1572 913
rect 1566 899 1572 900
rect 1566 895 1567 899
rect 1571 895 1572 899
rect 1566 894 1572 895
rect 1398 888 1404 889
rect 1398 884 1399 888
rect 1403 884 1404 888
rect 1398 883 1404 884
rect 1438 887 1444 888
rect 1438 883 1439 887
rect 1443 883 1444 887
rect 1400 879 1402 883
rect 1438 882 1444 883
rect 1391 878 1395 879
rect 1391 873 1395 874
rect 1399 878 1403 879
rect 1399 873 1403 874
rect 1390 872 1396 873
rect 1094 868 1095 872
rect 1099 868 1100 872
rect 1094 867 1100 868
rect 1162 871 1168 872
rect 1162 867 1163 871
rect 1167 867 1168 871
rect 1390 868 1391 872
rect 1395 868 1396 872
rect 1390 867 1396 868
rect 1430 871 1436 872
rect 1430 867 1431 871
rect 1435 867 1436 871
rect 1162 866 1168 867
rect 1430 866 1436 867
rect 1078 827 1084 828
rect 1078 823 1079 827
rect 1083 823 1084 827
rect 1078 822 1084 823
rect 1094 826 1100 827
rect 1094 822 1095 826
rect 1099 822 1100 826
rect 1094 821 1100 822
rect 1390 826 1396 827
rect 1390 822 1391 826
rect 1395 822 1396 826
rect 1390 821 1396 822
rect 838 819 844 820
rect 838 815 839 819
rect 843 815 844 819
rect 838 814 844 815
rect 1096 795 1098 821
rect 1158 819 1164 820
rect 1158 815 1159 819
rect 1163 815 1164 819
rect 1158 814 1164 815
rect 383 794 387 795
rect 383 789 387 790
rect 527 794 531 795
rect 527 789 531 790
rect 623 794 627 795
rect 623 789 627 790
rect 807 794 811 795
rect 807 789 811 790
rect 871 794 875 795
rect 871 789 875 790
rect 1095 794 1099 795
rect 1095 789 1099 790
rect 1127 794 1131 795
rect 1127 789 1131 790
rect 286 787 292 788
rect 286 783 287 787
rect 291 783 292 787
rect 384 783 386 789
rect 624 783 626 789
rect 872 783 874 789
rect 1128 783 1130 789
rect 166 782 172 783
rect 286 782 292 783
rect 382 782 388 783
rect 166 778 167 782
rect 171 778 172 782
rect 166 777 172 778
rect 382 778 383 782
rect 387 778 388 782
rect 382 777 388 778
rect 622 782 628 783
rect 622 778 623 782
rect 627 778 628 782
rect 622 777 628 778
rect 870 782 876 783
rect 870 778 871 782
rect 875 778 876 782
rect 870 777 876 778
rect 1126 782 1132 783
rect 1126 778 1127 782
rect 1131 778 1132 782
rect 1126 777 1132 778
rect 318 771 324 772
rect 318 767 319 771
rect 323 767 324 771
rect 318 766 324 767
rect 542 771 548 772
rect 542 767 543 771
rect 547 767 548 771
rect 542 766 548 767
rect 786 771 792 772
rect 786 767 787 771
rect 791 767 792 771
rect 786 766 792 767
rect 110 765 116 766
rect 110 761 111 765
rect 115 761 116 765
rect 110 760 116 761
rect 110 747 116 748
rect 110 743 111 747
rect 115 743 116 747
rect 110 742 116 743
rect 112 711 114 742
rect 166 736 172 737
rect 320 736 322 766
rect 382 736 388 737
rect 544 736 546 766
rect 622 736 628 737
rect 788 736 790 766
rect 870 736 876 737
rect 1126 736 1132 737
rect 1160 736 1162 814
rect 1392 795 1394 821
rect 1391 794 1395 795
rect 1391 789 1395 790
rect 1392 783 1394 789
rect 1432 788 1434 866
rect 1440 828 1442 882
rect 1568 879 1570 894
rect 1567 878 1571 879
rect 1567 873 1571 874
rect 1568 862 1570 873
rect 1566 861 1572 862
rect 1566 857 1567 861
rect 1571 857 1572 861
rect 1566 856 1572 857
rect 1566 843 1572 844
rect 1566 839 1567 843
rect 1571 839 1572 843
rect 1566 838 1572 839
rect 1438 827 1444 828
rect 1438 823 1439 827
rect 1443 823 1444 827
rect 1438 822 1444 823
rect 1568 795 1570 838
rect 1567 794 1571 795
rect 1567 789 1571 790
rect 1430 787 1436 788
rect 1430 783 1431 787
rect 1435 783 1436 787
rect 1390 782 1396 783
rect 1430 782 1436 783
rect 1262 779 1268 780
rect 1262 775 1263 779
rect 1267 775 1268 779
rect 1390 778 1391 782
rect 1395 778 1396 782
rect 1390 777 1396 778
rect 1262 774 1268 775
rect 166 732 167 736
rect 171 732 172 736
rect 166 731 172 732
rect 318 735 324 736
rect 318 731 319 735
rect 323 731 324 735
rect 382 732 383 736
rect 387 732 388 736
rect 382 731 388 732
rect 542 735 548 736
rect 542 731 543 735
rect 547 731 548 735
rect 622 732 623 736
rect 627 732 628 736
rect 622 731 628 732
rect 786 735 792 736
rect 786 731 787 735
rect 791 731 792 735
rect 870 732 871 736
rect 875 732 876 736
rect 870 731 876 732
rect 902 735 908 736
rect 902 731 903 735
rect 907 731 908 735
rect 1126 732 1127 736
rect 1131 732 1132 736
rect 1126 731 1132 732
rect 1158 735 1164 736
rect 1158 731 1159 735
rect 1163 731 1164 735
rect 168 711 170 731
rect 318 730 324 731
rect 384 711 386 731
rect 542 730 548 731
rect 624 711 626 731
rect 786 730 792 731
rect 872 711 874 731
rect 902 730 908 731
rect 111 710 115 711
rect 111 705 115 706
rect 167 710 171 711
rect 167 705 171 706
rect 319 710 323 711
rect 319 705 323 706
rect 383 710 387 711
rect 383 705 387 706
rect 575 710 579 711
rect 575 705 579 706
rect 623 710 627 711
rect 623 705 627 706
rect 839 710 843 711
rect 839 705 843 706
rect 871 710 875 711
rect 871 705 875 706
rect 112 694 114 705
rect 318 704 324 705
rect 318 700 319 704
rect 323 700 324 704
rect 318 699 324 700
rect 574 704 580 705
rect 838 704 844 705
rect 574 700 575 704
rect 579 700 580 704
rect 574 699 580 700
rect 606 703 612 704
rect 606 699 607 703
rect 611 699 612 703
rect 838 700 839 704
rect 843 700 844 704
rect 838 699 844 700
rect 854 703 860 704
rect 854 699 855 703
rect 859 699 860 703
rect 606 698 612 699
rect 854 698 860 699
rect 110 693 116 694
rect 110 689 111 693
rect 115 689 116 693
rect 110 688 116 689
rect 110 675 116 676
rect 110 671 111 675
rect 115 671 116 675
rect 110 670 116 671
rect 112 635 114 670
rect 318 658 324 659
rect 318 654 319 658
rect 323 654 324 658
rect 318 653 324 654
rect 574 658 580 659
rect 574 654 575 658
rect 579 654 580 658
rect 574 653 580 654
rect 320 635 322 653
rect 576 635 578 653
rect 608 652 610 698
rect 838 658 844 659
rect 838 654 839 658
rect 843 654 844 658
rect 838 653 844 654
rect 606 651 612 652
rect 606 647 607 651
rect 611 647 612 651
rect 606 646 612 647
rect 840 635 842 653
rect 856 652 858 698
rect 904 660 906 730
rect 1128 711 1130 731
rect 1158 730 1164 731
rect 1119 710 1123 711
rect 1119 705 1123 706
rect 1127 710 1131 711
rect 1127 705 1131 706
rect 1118 704 1124 705
rect 1118 700 1119 704
rect 1123 700 1124 704
rect 1118 699 1124 700
rect 1150 703 1156 704
rect 1150 699 1151 703
rect 1155 699 1156 703
rect 1150 698 1156 699
rect 978 687 984 688
rect 978 683 979 687
rect 983 683 984 687
rect 978 682 984 683
rect 902 659 908 660
rect 902 655 903 659
rect 907 655 908 659
rect 902 654 908 655
rect 980 652 982 682
rect 1118 658 1124 659
rect 1118 654 1119 658
rect 1123 654 1124 658
rect 1118 653 1124 654
rect 854 651 860 652
rect 854 647 855 651
rect 859 647 860 651
rect 854 646 860 647
rect 978 651 984 652
rect 978 647 979 651
rect 983 647 984 651
rect 978 646 984 647
rect 1120 635 1122 653
rect 111 634 115 635
rect 111 629 115 630
rect 319 634 323 635
rect 319 629 323 630
rect 575 634 579 635
rect 575 629 579 630
rect 583 634 587 635
rect 583 629 587 630
rect 727 634 731 635
rect 727 629 731 630
rect 839 634 843 635
rect 839 629 843 630
rect 887 634 891 635
rect 887 629 891 630
rect 1055 634 1059 635
rect 1055 629 1059 630
rect 1119 634 1123 635
rect 1119 629 1123 630
rect 112 606 114 629
rect 584 623 586 629
rect 728 623 730 629
rect 888 623 890 629
rect 1056 623 1058 629
rect 1152 628 1154 698
rect 1231 634 1235 635
rect 1231 629 1235 630
rect 1150 627 1156 628
rect 1150 623 1151 627
rect 1155 623 1156 627
rect 1232 623 1234 629
rect 582 622 588 623
rect 582 618 583 622
rect 587 618 588 622
rect 582 617 588 618
rect 726 622 732 623
rect 726 618 727 622
rect 731 618 732 622
rect 726 617 732 618
rect 886 622 892 623
rect 886 618 887 622
rect 891 618 892 622
rect 886 617 892 618
rect 1054 622 1060 623
rect 1150 622 1156 623
rect 1230 622 1236 623
rect 1054 618 1055 622
rect 1059 618 1060 622
rect 1054 617 1060 618
rect 1230 618 1231 622
rect 1235 618 1236 622
rect 1230 617 1236 618
rect 742 611 748 612
rect 742 607 743 611
rect 747 607 748 611
rect 742 606 748 607
rect 902 611 908 612
rect 902 607 903 611
rect 907 607 908 611
rect 902 606 908 607
rect 1070 611 1076 612
rect 1070 607 1071 611
rect 1075 607 1076 611
rect 1070 606 1076 607
rect 110 605 116 606
rect 110 601 111 605
rect 115 601 116 605
rect 110 600 116 601
rect 110 587 116 588
rect 110 583 111 587
rect 115 583 116 587
rect 110 582 116 583
rect 112 551 114 582
rect 582 576 588 577
rect 726 576 732 577
rect 744 576 746 606
rect 886 576 892 577
rect 904 576 906 606
rect 1054 576 1060 577
rect 1072 576 1074 606
rect 1230 576 1236 577
rect 1264 576 1266 774
rect 1568 766 1570 789
rect 1566 765 1572 766
rect 1566 761 1567 765
rect 1571 761 1572 765
rect 1566 760 1572 761
rect 1566 747 1572 748
rect 1566 743 1567 747
rect 1571 743 1572 747
rect 1566 742 1572 743
rect 1390 736 1396 737
rect 1390 732 1391 736
rect 1395 732 1396 736
rect 1390 731 1396 732
rect 1446 735 1452 736
rect 1446 731 1447 735
rect 1451 731 1452 735
rect 1392 711 1394 731
rect 1446 730 1452 731
rect 1391 710 1395 711
rect 1391 705 1395 706
rect 1399 710 1403 711
rect 1399 705 1403 706
rect 1398 704 1404 705
rect 1398 700 1399 704
rect 1403 700 1404 704
rect 1398 699 1404 700
rect 1448 660 1450 730
rect 1568 711 1570 742
rect 1567 710 1571 711
rect 1567 705 1571 706
rect 1454 703 1460 704
rect 1454 699 1455 703
rect 1459 699 1460 703
rect 1454 698 1460 699
rect 1446 659 1452 660
rect 1398 658 1404 659
rect 1398 654 1399 658
rect 1403 654 1404 658
rect 1446 655 1447 659
rect 1451 655 1452 659
rect 1446 654 1452 655
rect 1398 653 1404 654
rect 1400 635 1402 653
rect 1399 634 1403 635
rect 1399 629 1403 630
rect 1407 634 1411 635
rect 1407 629 1411 630
rect 1408 623 1410 629
rect 1456 628 1458 698
rect 1568 694 1570 705
rect 1566 693 1572 694
rect 1566 689 1567 693
rect 1571 689 1572 693
rect 1566 688 1572 689
rect 1566 675 1572 676
rect 1566 671 1567 675
rect 1571 671 1572 675
rect 1566 670 1572 671
rect 1568 635 1570 670
rect 1567 634 1571 635
rect 1567 629 1571 630
rect 1454 627 1460 628
rect 1454 623 1455 627
rect 1459 623 1460 627
rect 1406 622 1412 623
rect 1454 622 1460 623
rect 1274 619 1280 620
rect 1274 615 1275 619
rect 1279 615 1280 619
rect 1406 618 1407 622
rect 1411 618 1412 622
rect 1406 617 1412 618
rect 1274 614 1280 615
rect 582 572 583 576
rect 587 572 588 576
rect 582 571 588 572
rect 650 575 656 576
rect 650 571 651 575
rect 655 571 656 575
rect 726 572 727 576
rect 731 572 732 576
rect 726 571 732 572
rect 742 575 748 576
rect 742 571 743 575
rect 747 571 748 575
rect 886 572 887 576
rect 891 572 892 576
rect 886 571 892 572
rect 902 575 908 576
rect 902 571 903 575
rect 907 571 908 575
rect 1054 572 1055 576
rect 1059 572 1060 576
rect 1054 571 1060 572
rect 1070 575 1076 576
rect 1070 571 1071 575
rect 1075 571 1076 575
rect 1230 572 1231 576
rect 1235 572 1236 576
rect 1230 571 1236 572
rect 1262 575 1268 576
rect 1262 571 1263 575
rect 1267 571 1268 575
rect 584 551 586 571
rect 650 570 656 571
rect 111 550 115 551
rect 111 545 115 546
rect 583 550 587 551
rect 583 545 587 546
rect 112 534 114 545
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 112 475 114 510
rect 652 508 654 570
rect 728 551 730 571
rect 742 570 748 571
rect 888 551 890 571
rect 902 570 908 571
rect 1056 551 1058 571
rect 1070 570 1076 571
rect 1232 551 1234 571
rect 1262 570 1268 571
rect 727 550 731 551
rect 727 545 731 546
rect 759 550 763 551
rect 759 545 763 546
rect 863 550 867 551
rect 863 545 867 546
rect 887 550 891 551
rect 887 545 891 546
rect 975 550 979 551
rect 975 545 979 546
rect 1055 550 1059 551
rect 1055 545 1059 546
rect 1087 550 1091 551
rect 1087 545 1091 546
rect 1207 550 1211 551
rect 1207 545 1211 546
rect 1231 550 1235 551
rect 1231 545 1235 546
rect 758 544 764 545
rect 862 544 868 545
rect 974 544 980 545
rect 1086 544 1092 545
rect 1206 544 1212 545
rect 1276 544 1278 614
rect 1568 606 1570 629
rect 1566 605 1572 606
rect 1566 601 1567 605
rect 1571 601 1572 605
rect 1566 600 1572 601
rect 1566 587 1572 588
rect 1566 583 1567 587
rect 1571 583 1572 587
rect 1566 582 1572 583
rect 1406 576 1412 577
rect 1406 572 1407 576
rect 1411 572 1412 576
rect 1406 571 1412 572
rect 1438 575 1444 576
rect 1438 571 1439 575
rect 1443 571 1444 575
rect 1408 551 1410 571
rect 1438 570 1444 571
rect 1327 550 1331 551
rect 1327 545 1331 546
rect 1407 550 1411 551
rect 1407 545 1411 546
rect 1326 544 1332 545
rect 758 540 759 544
rect 763 540 764 544
rect 758 539 764 540
rect 826 543 832 544
rect 826 539 827 543
rect 831 539 832 543
rect 862 540 863 544
rect 867 540 868 544
rect 862 539 868 540
rect 930 543 936 544
rect 930 539 931 543
rect 935 539 936 543
rect 974 540 975 544
rect 979 540 980 544
rect 974 539 980 540
rect 1042 543 1048 544
rect 1042 539 1043 543
rect 1047 539 1048 543
rect 1086 540 1087 544
rect 1091 540 1092 544
rect 1086 539 1092 540
rect 1118 543 1124 544
rect 1118 539 1119 543
rect 1123 539 1124 543
rect 1206 540 1207 544
rect 1211 540 1212 544
rect 1206 539 1212 540
rect 1274 543 1280 544
rect 1274 539 1275 543
rect 1279 539 1280 543
rect 1326 540 1327 544
rect 1331 540 1332 544
rect 1326 539 1332 540
rect 1394 543 1400 544
rect 1394 539 1395 543
rect 1399 539 1400 543
rect 826 538 832 539
rect 930 538 936 539
rect 1042 538 1048 539
rect 1118 538 1124 539
rect 1274 538 1280 539
rect 1394 538 1400 539
rect 650 507 656 508
rect 650 503 651 507
rect 655 503 656 507
rect 650 502 656 503
rect 758 498 764 499
rect 758 494 759 498
rect 763 494 764 498
rect 758 493 764 494
rect 760 475 762 493
rect 828 492 830 538
rect 862 498 868 499
rect 862 494 863 498
rect 867 494 868 498
rect 862 493 868 494
rect 826 491 832 492
rect 826 487 827 491
rect 831 487 832 491
rect 826 486 832 487
rect 864 475 866 493
rect 932 492 934 538
rect 974 498 980 499
rect 974 494 975 498
rect 979 494 980 498
rect 974 493 980 494
rect 930 491 936 492
rect 930 487 931 491
rect 935 487 936 491
rect 930 486 936 487
rect 976 475 978 493
rect 1044 492 1046 538
rect 1086 498 1092 499
rect 1086 494 1087 498
rect 1091 494 1092 498
rect 1086 493 1092 494
rect 1042 491 1048 492
rect 1042 487 1043 491
rect 1047 487 1048 491
rect 1042 486 1048 487
rect 1088 475 1090 493
rect 111 474 115 475
rect 111 469 115 470
rect 719 474 723 475
rect 719 469 723 470
rect 759 474 763 475
rect 759 469 763 470
rect 823 474 827 475
rect 823 469 827 470
rect 863 474 867 475
rect 863 469 867 470
rect 927 474 931 475
rect 927 469 931 470
rect 975 474 979 475
rect 975 469 979 470
rect 1031 474 1035 475
rect 1031 469 1035 470
rect 1087 474 1091 475
rect 1087 469 1091 470
rect 112 446 114 469
rect 720 463 722 469
rect 824 463 826 469
rect 928 463 930 469
rect 1032 463 1034 469
rect 1120 468 1122 538
rect 1206 498 1212 499
rect 1206 494 1207 498
rect 1211 494 1212 498
rect 1206 493 1212 494
rect 1326 498 1332 499
rect 1326 494 1327 498
rect 1331 494 1332 498
rect 1326 493 1332 494
rect 1208 475 1210 493
rect 1214 491 1220 492
rect 1214 487 1215 491
rect 1219 487 1220 491
rect 1214 486 1220 487
rect 1135 474 1139 475
rect 1135 469 1139 470
rect 1207 474 1211 475
rect 1207 469 1211 470
rect 1118 467 1124 468
rect 1118 463 1119 467
rect 1123 463 1124 467
rect 1136 463 1138 469
rect 718 462 724 463
rect 718 458 719 462
rect 723 458 724 462
rect 718 457 724 458
rect 822 462 828 463
rect 822 458 823 462
rect 827 458 828 462
rect 822 457 828 458
rect 926 462 932 463
rect 926 458 927 462
rect 931 458 932 462
rect 926 457 932 458
rect 1030 462 1036 463
rect 1118 462 1124 463
rect 1134 462 1140 463
rect 1030 458 1031 462
rect 1035 458 1036 462
rect 1030 457 1036 458
rect 1134 458 1135 462
rect 1139 458 1140 462
rect 1134 457 1140 458
rect 838 451 844 452
rect 838 447 839 451
rect 843 447 844 451
rect 838 446 844 447
rect 942 451 948 452
rect 942 447 943 451
rect 947 447 948 451
rect 942 446 948 447
rect 1046 451 1052 452
rect 1046 447 1047 451
rect 1051 447 1052 451
rect 1046 446 1052 447
rect 110 445 116 446
rect 110 441 111 445
rect 115 441 116 445
rect 110 440 116 441
rect 110 427 116 428
rect 110 423 111 427
rect 115 423 116 427
rect 110 422 116 423
rect 112 383 114 422
rect 718 416 724 417
rect 822 416 828 417
rect 840 416 842 446
rect 926 416 932 417
rect 944 416 946 446
rect 1030 416 1036 417
rect 1048 416 1050 446
rect 1134 416 1140 417
rect 1216 416 1218 486
rect 1328 475 1330 493
rect 1396 492 1398 538
rect 1440 500 1442 570
rect 1568 551 1570 582
rect 1447 550 1451 551
rect 1447 545 1451 546
rect 1567 550 1571 551
rect 1567 545 1571 546
rect 1446 544 1452 545
rect 1446 540 1447 544
rect 1451 540 1452 544
rect 1446 539 1452 540
rect 1510 543 1516 544
rect 1510 539 1511 543
rect 1515 539 1516 543
rect 1510 538 1516 539
rect 1438 499 1444 500
rect 1438 495 1439 499
rect 1443 495 1444 499
rect 1438 494 1444 495
rect 1446 498 1452 499
rect 1446 494 1447 498
rect 1451 494 1452 498
rect 1446 493 1452 494
rect 1394 491 1400 492
rect 1394 487 1395 491
rect 1399 487 1400 491
rect 1394 486 1400 487
rect 1448 475 1450 493
rect 1239 474 1243 475
rect 1239 469 1243 470
rect 1327 474 1331 475
rect 1327 469 1331 470
rect 1351 474 1355 475
rect 1351 469 1355 470
rect 1447 474 1451 475
rect 1447 469 1451 470
rect 1463 474 1467 475
rect 1463 469 1467 470
rect 1240 463 1242 469
rect 1352 463 1354 469
rect 1464 463 1466 469
rect 1512 468 1514 538
rect 1568 534 1570 545
rect 1566 533 1572 534
rect 1566 529 1567 533
rect 1571 529 1572 533
rect 1566 528 1572 529
rect 1566 515 1572 516
rect 1566 511 1567 515
rect 1571 511 1572 515
rect 1566 510 1572 511
rect 1568 475 1570 510
rect 1567 474 1571 475
rect 1567 469 1571 470
rect 1510 467 1516 468
rect 1510 463 1511 467
rect 1515 463 1516 467
rect 1238 462 1244 463
rect 1238 458 1239 462
rect 1243 458 1244 462
rect 1238 457 1244 458
rect 1350 462 1356 463
rect 1350 458 1351 462
rect 1355 458 1356 462
rect 1350 457 1356 458
rect 1462 462 1468 463
rect 1510 462 1516 463
rect 1462 458 1463 462
rect 1467 458 1468 462
rect 1462 457 1468 458
rect 1254 451 1260 452
rect 1254 447 1255 451
rect 1259 447 1260 451
rect 1254 446 1260 447
rect 1366 451 1372 452
rect 1366 447 1367 451
rect 1371 447 1372 451
rect 1366 446 1372 447
rect 1478 451 1484 452
rect 1478 447 1479 451
rect 1483 447 1484 451
rect 1478 446 1484 447
rect 1568 446 1570 469
rect 1238 416 1244 417
rect 1256 416 1258 446
rect 1350 416 1356 417
rect 1368 416 1370 446
rect 1462 416 1468 417
rect 1480 416 1482 446
rect 1566 445 1572 446
rect 1566 441 1567 445
rect 1571 441 1572 445
rect 1566 440 1572 441
rect 1566 427 1572 428
rect 1566 423 1567 427
rect 1571 423 1572 427
rect 1566 422 1572 423
rect 718 412 719 416
rect 723 412 724 416
rect 718 411 724 412
rect 798 415 804 416
rect 798 411 799 415
rect 803 411 804 415
rect 822 412 823 416
rect 827 412 828 416
rect 822 411 828 412
rect 838 415 844 416
rect 838 411 839 415
rect 843 411 844 415
rect 926 412 927 416
rect 931 412 932 416
rect 926 411 932 412
rect 942 415 948 416
rect 942 411 943 415
rect 947 411 948 415
rect 1030 412 1031 416
rect 1035 412 1036 416
rect 1030 411 1036 412
rect 1046 415 1052 416
rect 1046 411 1047 415
rect 1051 411 1052 415
rect 1134 412 1135 416
rect 1139 412 1140 416
rect 1134 411 1140 412
rect 1214 415 1220 416
rect 1214 411 1215 415
rect 1219 411 1220 415
rect 1238 412 1239 416
rect 1243 412 1244 416
rect 1238 411 1244 412
rect 1254 415 1260 416
rect 1254 411 1255 415
rect 1259 411 1260 415
rect 1350 412 1351 416
rect 1355 412 1356 416
rect 1350 411 1356 412
rect 1366 415 1372 416
rect 1366 411 1367 415
rect 1371 411 1372 415
rect 1462 412 1463 416
rect 1467 412 1468 416
rect 1462 411 1468 412
rect 1478 415 1484 416
rect 1478 411 1479 415
rect 1483 411 1484 415
rect 720 383 722 411
rect 798 410 804 411
rect 111 382 115 383
rect 111 377 115 378
rect 511 382 515 383
rect 511 377 515 378
rect 599 382 603 383
rect 599 377 603 378
rect 687 382 691 383
rect 687 377 691 378
rect 719 382 723 383
rect 719 377 723 378
rect 775 382 779 383
rect 775 377 779 378
rect 112 366 114 377
rect 510 376 516 377
rect 598 376 604 377
rect 686 376 692 377
rect 774 376 780 377
rect 510 372 511 376
rect 515 372 516 376
rect 510 371 516 372
rect 578 375 584 376
rect 578 371 579 375
rect 583 371 584 375
rect 598 372 599 376
rect 603 372 604 376
rect 598 371 604 372
rect 630 375 636 376
rect 630 371 631 375
rect 635 371 636 375
rect 686 372 687 376
rect 691 372 692 376
rect 686 371 692 372
rect 702 375 708 376
rect 702 371 703 375
rect 707 371 708 375
rect 774 372 775 376
rect 779 372 780 376
rect 774 371 780 372
rect 578 370 584 371
rect 630 370 636 371
rect 702 370 708 371
rect 110 365 116 366
rect 110 361 111 365
rect 115 361 116 365
rect 110 360 116 361
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 110 342 116 343
rect 112 311 114 342
rect 510 330 516 331
rect 510 326 511 330
rect 515 326 516 330
rect 510 325 516 326
rect 512 311 514 325
rect 111 310 115 311
rect 111 305 115 306
rect 375 310 379 311
rect 375 305 379 306
rect 463 310 467 311
rect 463 305 467 306
rect 511 310 515 311
rect 511 305 515 306
rect 551 310 555 311
rect 551 305 555 306
rect 112 282 114 305
rect 376 299 378 305
rect 464 299 466 305
rect 552 299 554 305
rect 580 304 582 370
rect 598 330 604 331
rect 598 326 599 330
rect 603 326 604 330
rect 598 325 604 326
rect 600 311 602 325
rect 632 324 634 370
rect 686 330 692 331
rect 686 326 687 330
rect 691 326 692 330
rect 686 325 692 326
rect 630 323 636 324
rect 630 319 631 323
rect 635 319 636 323
rect 630 318 636 319
rect 688 311 690 325
rect 704 324 706 370
rect 800 332 802 410
rect 824 383 826 411
rect 838 410 844 411
rect 928 383 930 411
rect 942 410 948 411
rect 1032 383 1034 411
rect 1046 410 1052 411
rect 1136 383 1138 411
rect 1214 410 1220 411
rect 1240 383 1242 411
rect 1254 410 1260 411
rect 1352 383 1354 411
rect 1366 410 1372 411
rect 1464 383 1466 411
rect 1478 410 1484 411
rect 1568 383 1570 422
rect 823 382 827 383
rect 823 377 827 378
rect 927 382 931 383
rect 927 377 931 378
rect 1031 382 1035 383
rect 1031 377 1035 378
rect 1135 382 1139 383
rect 1135 377 1139 378
rect 1239 382 1243 383
rect 1239 377 1243 378
rect 1351 382 1355 383
rect 1351 377 1355 378
rect 1463 382 1467 383
rect 1463 377 1467 378
rect 1567 382 1571 383
rect 1567 377 1571 378
rect 806 375 812 376
rect 806 371 807 375
rect 811 371 812 375
rect 806 370 812 371
rect 798 331 804 332
rect 774 330 780 331
rect 774 326 775 330
rect 779 326 780 330
rect 798 327 799 331
rect 803 327 804 331
rect 798 326 804 327
rect 774 325 780 326
rect 702 323 708 324
rect 702 319 703 323
rect 707 319 708 323
rect 702 318 708 319
rect 776 311 778 325
rect 808 324 810 370
rect 1568 366 1570 377
rect 1566 365 1572 366
rect 1566 361 1567 365
rect 1571 361 1572 365
rect 1566 360 1572 361
rect 1566 347 1572 348
rect 1566 343 1567 347
rect 1571 343 1572 347
rect 1566 342 1572 343
rect 806 323 812 324
rect 806 319 807 323
rect 811 319 812 323
rect 806 318 812 319
rect 1568 311 1570 342
rect 599 310 603 311
rect 599 305 603 306
rect 687 310 691 311
rect 687 305 691 306
rect 775 310 779 311
rect 775 305 779 306
rect 1567 310 1571 311
rect 1567 305 1571 306
rect 578 303 584 304
rect 578 299 579 303
rect 583 299 584 303
rect 374 298 380 299
rect 374 294 375 298
rect 379 294 380 298
rect 374 293 380 294
rect 462 298 468 299
rect 462 294 463 298
rect 467 294 468 298
rect 462 293 468 294
rect 550 298 556 299
rect 578 298 584 299
rect 550 294 551 298
rect 555 294 556 298
rect 550 293 556 294
rect 478 287 484 288
rect 478 283 479 287
rect 483 283 484 287
rect 478 282 484 283
rect 566 287 572 288
rect 566 283 567 287
rect 571 283 572 287
rect 566 282 572 283
rect 1568 282 1570 305
rect 110 281 116 282
rect 110 277 111 281
rect 115 277 116 281
rect 110 276 116 277
rect 110 263 116 264
rect 110 259 111 263
rect 115 259 116 263
rect 110 258 116 259
rect 112 247 114 258
rect 374 252 380 253
rect 462 252 468 253
rect 480 252 482 282
rect 550 252 556 253
rect 568 252 570 282
rect 1566 281 1572 282
rect 1566 277 1567 281
rect 1571 277 1572 281
rect 1566 276 1572 277
rect 1566 263 1572 264
rect 1566 259 1567 263
rect 1571 259 1572 263
rect 1566 258 1572 259
rect 374 248 375 252
rect 379 248 380 252
rect 374 247 380 248
rect 406 251 412 252
rect 406 247 407 251
rect 411 247 412 251
rect 462 248 463 252
rect 467 248 468 252
rect 462 247 468 248
rect 478 251 484 252
rect 478 247 479 251
rect 483 247 484 251
rect 550 248 551 252
rect 555 248 556 252
rect 550 247 556 248
rect 566 251 572 252
rect 566 247 567 251
rect 571 247 572 251
rect 1568 247 1570 258
rect 111 246 115 247
rect 111 241 115 242
rect 247 246 251 247
rect 247 241 251 242
rect 335 246 339 247
rect 335 241 339 242
rect 375 246 379 247
rect 406 246 412 247
rect 423 246 427 247
rect 375 241 379 242
rect 112 230 114 241
rect 246 240 252 241
rect 246 236 247 240
rect 251 236 252 240
rect 246 235 252 236
rect 334 240 340 241
rect 334 236 335 240
rect 339 236 340 240
rect 334 235 340 236
rect 366 239 372 240
rect 366 235 367 239
rect 371 235 372 239
rect 366 234 372 235
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 110 211 116 212
rect 110 207 111 211
rect 115 207 116 211
rect 110 206 116 207
rect 112 155 114 206
rect 246 194 252 195
rect 246 190 247 194
rect 251 190 252 194
rect 246 189 252 190
rect 334 194 340 195
rect 334 190 335 194
rect 339 190 340 194
rect 334 189 340 190
rect 248 155 250 189
rect 336 155 338 189
rect 368 188 370 234
rect 408 196 410 246
rect 423 241 427 242
rect 463 246 467 247
rect 478 246 484 247
rect 551 246 555 247
rect 566 246 572 247
rect 1567 246 1571 247
rect 463 241 467 242
rect 551 241 555 242
rect 1567 241 1571 242
rect 422 240 428 241
rect 422 236 423 240
rect 427 236 428 240
rect 422 235 428 236
rect 582 239 588 240
rect 582 235 583 239
rect 587 235 588 239
rect 582 234 588 235
rect 406 195 412 196
rect 406 191 407 195
rect 411 191 412 195
rect 406 190 412 191
rect 422 194 428 195
rect 422 190 423 194
rect 427 190 428 194
rect 422 189 428 190
rect 366 187 372 188
rect 366 183 367 187
rect 371 183 372 187
rect 366 182 372 183
rect 424 155 426 189
rect 111 154 115 155
rect 111 149 115 150
rect 135 154 139 155
rect 135 149 139 150
rect 223 154 227 155
rect 223 149 227 150
rect 247 154 251 155
rect 247 149 251 150
rect 311 154 315 155
rect 311 149 315 150
rect 335 154 339 155
rect 335 149 339 150
rect 399 154 403 155
rect 399 149 403 150
rect 423 154 427 155
rect 423 149 427 150
rect 487 154 491 155
rect 487 149 491 150
rect 575 154 579 155
rect 575 149 579 150
rect 112 126 114 149
rect 136 143 138 149
rect 224 143 226 149
rect 312 143 314 149
rect 400 143 402 149
rect 488 143 490 149
rect 576 143 578 149
rect 584 148 586 234
rect 1568 230 1570 241
rect 1566 229 1572 230
rect 1566 225 1567 229
rect 1571 225 1572 229
rect 1566 224 1572 225
rect 1566 211 1572 212
rect 1566 207 1567 211
rect 1571 207 1572 211
rect 1566 206 1572 207
rect 1568 155 1570 206
rect 1567 154 1571 155
rect 1567 149 1571 150
rect 582 147 588 148
rect 582 143 583 147
rect 587 143 588 147
rect 134 142 140 143
rect 134 138 135 142
rect 139 138 140 142
rect 134 137 140 138
rect 222 142 228 143
rect 222 138 223 142
rect 227 138 228 142
rect 222 137 228 138
rect 310 142 316 143
rect 310 138 311 142
rect 315 138 316 142
rect 310 137 316 138
rect 398 142 404 143
rect 398 138 399 142
rect 403 138 404 142
rect 398 137 404 138
rect 486 142 492 143
rect 486 138 487 142
rect 491 138 492 142
rect 486 137 492 138
rect 574 142 580 143
rect 582 142 588 143
rect 574 138 575 142
rect 579 138 580 142
rect 574 137 580 138
rect 238 131 244 132
rect 238 127 239 131
rect 243 127 244 131
rect 238 126 244 127
rect 326 131 332 132
rect 326 127 327 131
rect 331 127 332 131
rect 326 126 332 127
rect 414 131 420 132
rect 414 127 415 131
rect 419 127 420 131
rect 414 126 420 127
rect 502 131 508 132
rect 502 127 503 131
rect 507 127 508 131
rect 502 126 508 127
rect 590 131 596 132
rect 590 127 591 131
rect 595 127 596 131
rect 590 126 596 127
rect 1568 126 1570 149
rect 110 125 116 126
rect 110 121 111 125
rect 115 121 116 125
rect 110 120 116 121
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 110 102 116 103
rect 112 91 114 102
rect 134 96 140 97
rect 134 92 135 96
rect 139 92 140 96
rect 134 91 140 92
rect 222 96 228 97
rect 240 96 242 126
rect 310 96 316 97
rect 328 96 330 126
rect 398 96 404 97
rect 416 96 418 126
rect 486 96 492 97
rect 504 96 506 126
rect 574 96 580 97
rect 592 96 594 126
rect 1566 125 1572 126
rect 1566 121 1567 125
rect 1571 121 1572 125
rect 1566 120 1572 121
rect 1566 107 1572 108
rect 1566 103 1567 107
rect 1571 103 1572 107
rect 1566 102 1572 103
rect 222 92 223 96
rect 227 92 228 96
rect 222 91 228 92
rect 238 95 244 96
rect 238 91 239 95
rect 243 91 244 95
rect 310 92 311 96
rect 315 92 316 96
rect 310 91 316 92
rect 326 95 332 96
rect 326 91 327 95
rect 331 91 332 95
rect 398 92 399 96
rect 403 92 404 96
rect 398 91 404 92
rect 414 95 420 96
rect 414 91 415 95
rect 419 91 420 95
rect 486 92 487 96
rect 491 92 492 96
rect 486 91 492 92
rect 502 95 508 96
rect 502 91 503 95
rect 507 91 508 95
rect 574 92 575 96
rect 579 92 580 96
rect 574 91 580 92
rect 590 95 596 96
rect 590 91 591 95
rect 595 91 596 95
rect 1568 91 1570 102
rect 111 90 115 91
rect 111 85 115 86
rect 135 90 139 91
rect 135 85 139 86
rect 223 90 227 91
rect 238 90 244 91
rect 311 90 315 91
rect 326 90 332 91
rect 399 90 403 91
rect 414 90 420 91
rect 487 90 491 91
rect 502 90 508 91
rect 575 90 579 91
rect 590 90 596 91
rect 1567 90 1571 91
rect 223 85 227 86
rect 311 85 315 86
rect 399 85 403 86
rect 487 85 491 86
rect 575 85 579 86
rect 1567 85 1571 86
<< m4c >>
rect 111 1518 115 1522
rect 399 1518 403 1522
rect 487 1518 491 1522
rect 575 1518 579 1522
rect 671 1518 675 1522
rect 783 1518 787 1522
rect 903 1518 907 1522
rect 1031 1518 1035 1522
rect 1167 1518 1171 1522
rect 1303 1518 1307 1522
rect 1447 1518 1451 1522
rect 1567 1518 1571 1522
rect 111 1442 115 1446
rect 399 1442 403 1446
rect 423 1442 427 1446
rect 487 1442 491 1446
rect 575 1442 579 1446
rect 655 1442 659 1446
rect 671 1442 675 1446
rect 783 1442 787 1446
rect 895 1442 899 1446
rect 903 1442 907 1446
rect 1031 1442 1035 1446
rect 1143 1442 1147 1446
rect 1167 1442 1171 1446
rect 1303 1442 1307 1446
rect 1399 1442 1403 1446
rect 1447 1442 1451 1446
rect 111 1374 115 1378
rect 423 1374 427 1378
rect 471 1374 475 1378
rect 655 1374 659 1378
rect 695 1374 699 1378
rect 895 1374 899 1378
rect 919 1374 923 1378
rect 1143 1374 1147 1378
rect 1151 1374 1155 1378
rect 111 1302 115 1306
rect 471 1302 475 1306
rect 519 1302 523 1306
rect 695 1302 699 1306
rect 743 1302 747 1306
rect 919 1302 923 1306
rect 975 1302 979 1306
rect 1391 1374 1395 1378
rect 1399 1374 1403 1378
rect 1567 1442 1571 1446
rect 1567 1374 1571 1378
rect 1151 1302 1155 1306
rect 1207 1302 1211 1306
rect 1391 1302 1395 1306
rect 111 1222 115 1226
rect 519 1222 523 1226
rect 567 1222 571 1226
rect 743 1222 747 1226
rect 767 1222 771 1226
rect 967 1222 971 1226
rect 975 1222 979 1226
rect 1175 1222 1179 1226
rect 1439 1302 1443 1306
rect 1567 1302 1571 1306
rect 1207 1222 1211 1226
rect 1391 1222 1395 1226
rect 1439 1222 1443 1226
rect 1567 1222 1571 1226
rect 111 1158 115 1162
rect 567 1158 571 1162
rect 703 1158 707 1162
rect 767 1158 771 1162
rect 967 1158 971 1162
rect 1055 1158 1059 1162
rect 1175 1158 1179 1162
rect 111 1094 115 1098
rect 671 1094 675 1098
rect 703 1094 707 1098
rect 847 1094 851 1098
rect 1031 1094 1035 1098
rect 1055 1094 1059 1098
rect 1223 1094 1227 1098
rect 1391 1158 1395 1162
rect 1407 1158 1411 1162
rect 1567 1158 1571 1162
rect 1407 1094 1411 1098
rect 1415 1094 1419 1098
rect 1567 1094 1571 1098
rect 111 1014 115 1018
rect 575 1014 579 1018
rect 671 1014 675 1018
rect 775 1014 779 1018
rect 847 1014 851 1018
rect 983 1014 987 1018
rect 111 942 115 946
rect 407 942 411 946
rect 575 942 579 946
rect 1031 1014 1035 1018
rect 1191 1014 1195 1018
rect 1223 1014 1227 1018
rect 1407 1014 1411 1018
rect 1415 1014 1419 1018
rect 735 942 739 946
rect 775 942 779 946
rect 983 942 987 946
rect 1063 942 1067 946
rect 111 874 115 878
rect 255 874 259 878
rect 407 874 411 878
rect 527 874 531 878
rect 735 874 739 878
rect 807 874 811 878
rect 1063 874 1067 878
rect 111 790 115 794
rect 167 790 171 794
rect 255 790 259 794
rect 1095 874 1099 878
rect 1191 942 1195 946
rect 1399 942 1403 946
rect 1407 942 1411 946
rect 1567 1014 1571 1018
rect 1567 942 1571 946
rect 1391 874 1395 878
rect 1399 874 1403 878
rect 383 790 387 794
rect 527 790 531 794
rect 623 790 627 794
rect 807 790 811 794
rect 871 790 875 794
rect 1095 790 1099 794
rect 1127 790 1131 794
rect 1391 790 1395 794
rect 1567 874 1571 878
rect 1567 790 1571 794
rect 111 706 115 710
rect 167 706 171 710
rect 319 706 323 710
rect 383 706 387 710
rect 575 706 579 710
rect 623 706 627 710
rect 839 706 843 710
rect 871 706 875 710
rect 1119 706 1123 710
rect 1127 706 1131 710
rect 111 630 115 634
rect 319 630 323 634
rect 575 630 579 634
rect 583 630 587 634
rect 727 630 731 634
rect 839 630 843 634
rect 887 630 891 634
rect 1055 630 1059 634
rect 1119 630 1123 634
rect 1231 630 1235 634
rect 1391 706 1395 710
rect 1399 706 1403 710
rect 1567 706 1571 710
rect 1399 630 1403 634
rect 1407 630 1411 634
rect 1567 630 1571 634
rect 111 546 115 550
rect 583 546 587 550
rect 727 546 731 550
rect 759 546 763 550
rect 863 546 867 550
rect 887 546 891 550
rect 975 546 979 550
rect 1055 546 1059 550
rect 1087 546 1091 550
rect 1207 546 1211 550
rect 1231 546 1235 550
rect 1327 546 1331 550
rect 1407 546 1411 550
rect 111 470 115 474
rect 719 470 723 474
rect 759 470 763 474
rect 823 470 827 474
rect 863 470 867 474
rect 927 470 931 474
rect 975 470 979 474
rect 1031 470 1035 474
rect 1087 470 1091 474
rect 1135 470 1139 474
rect 1207 470 1211 474
rect 1447 546 1451 550
rect 1567 546 1571 550
rect 1239 470 1243 474
rect 1327 470 1331 474
rect 1351 470 1355 474
rect 1447 470 1451 474
rect 1463 470 1467 474
rect 1567 470 1571 474
rect 111 378 115 382
rect 511 378 515 382
rect 599 378 603 382
rect 687 378 691 382
rect 719 378 723 382
rect 775 378 779 382
rect 111 306 115 310
rect 375 306 379 310
rect 463 306 467 310
rect 511 306 515 310
rect 551 306 555 310
rect 823 378 827 382
rect 927 378 931 382
rect 1031 378 1035 382
rect 1135 378 1139 382
rect 1239 378 1243 382
rect 1351 378 1355 382
rect 1463 378 1467 382
rect 1567 378 1571 382
rect 599 306 603 310
rect 687 306 691 310
rect 775 306 779 310
rect 1567 306 1571 310
rect 111 242 115 246
rect 247 242 251 246
rect 335 242 339 246
rect 375 242 379 246
rect 423 242 427 246
rect 463 242 467 246
rect 551 242 555 246
rect 1567 242 1571 246
rect 111 150 115 154
rect 135 150 139 154
rect 223 150 227 154
rect 247 150 251 154
rect 311 150 315 154
rect 335 150 339 154
rect 399 150 403 154
rect 423 150 427 154
rect 487 150 491 154
rect 575 150 579 154
rect 1567 150 1571 154
rect 111 86 115 90
rect 135 86 139 90
rect 223 86 227 90
rect 311 86 315 90
rect 399 86 403 90
rect 487 86 491 90
rect 575 86 579 90
rect 1567 86 1571 90
<< m4 >>
rect 96 1517 97 1523
rect 103 1522 1603 1523
rect 103 1518 111 1522
rect 115 1518 399 1522
rect 403 1518 487 1522
rect 491 1518 575 1522
rect 579 1518 671 1522
rect 675 1518 783 1522
rect 787 1518 903 1522
rect 907 1518 1031 1522
rect 1035 1518 1167 1522
rect 1171 1518 1303 1522
rect 1307 1518 1447 1522
rect 1451 1518 1567 1522
rect 1571 1518 1603 1522
rect 103 1517 1603 1518
rect 1609 1517 1610 1523
rect 84 1441 85 1447
rect 91 1446 1591 1447
rect 91 1442 111 1446
rect 115 1442 399 1446
rect 403 1442 423 1446
rect 427 1442 487 1446
rect 491 1442 575 1446
rect 579 1442 655 1446
rect 659 1442 671 1446
rect 675 1442 783 1446
rect 787 1442 895 1446
rect 899 1442 903 1446
rect 907 1442 1031 1446
rect 1035 1442 1143 1446
rect 1147 1442 1167 1446
rect 1171 1442 1303 1446
rect 1307 1442 1399 1446
rect 1403 1442 1447 1446
rect 1451 1442 1567 1446
rect 1571 1442 1591 1446
rect 91 1441 1591 1442
rect 1597 1441 1598 1447
rect 96 1373 97 1379
rect 103 1378 1603 1379
rect 103 1374 111 1378
rect 115 1374 423 1378
rect 427 1374 471 1378
rect 475 1374 655 1378
rect 659 1374 695 1378
rect 699 1374 895 1378
rect 899 1374 919 1378
rect 923 1374 1143 1378
rect 1147 1374 1151 1378
rect 1155 1374 1391 1378
rect 1395 1374 1399 1378
rect 1403 1374 1567 1378
rect 1571 1374 1603 1378
rect 103 1373 1603 1374
rect 1609 1373 1610 1379
rect 84 1301 85 1307
rect 91 1306 1591 1307
rect 91 1302 111 1306
rect 115 1302 471 1306
rect 475 1302 519 1306
rect 523 1302 695 1306
rect 699 1302 743 1306
rect 747 1302 919 1306
rect 923 1302 975 1306
rect 979 1302 1151 1306
rect 1155 1302 1207 1306
rect 1211 1302 1391 1306
rect 1395 1302 1439 1306
rect 1443 1302 1567 1306
rect 1571 1302 1591 1306
rect 91 1301 1591 1302
rect 1597 1301 1598 1307
rect 96 1221 97 1227
rect 103 1226 1603 1227
rect 103 1222 111 1226
rect 115 1222 519 1226
rect 523 1222 567 1226
rect 571 1222 743 1226
rect 747 1222 767 1226
rect 771 1222 967 1226
rect 971 1222 975 1226
rect 979 1222 1175 1226
rect 1179 1222 1207 1226
rect 1211 1222 1391 1226
rect 1395 1222 1439 1226
rect 1443 1222 1567 1226
rect 1571 1222 1603 1226
rect 103 1221 1603 1222
rect 1609 1221 1610 1227
rect 84 1157 85 1163
rect 91 1162 1591 1163
rect 91 1158 111 1162
rect 115 1158 567 1162
rect 571 1158 703 1162
rect 707 1158 767 1162
rect 771 1158 967 1162
rect 971 1158 1055 1162
rect 1059 1158 1175 1162
rect 1179 1158 1391 1162
rect 1395 1158 1407 1162
rect 1411 1158 1567 1162
rect 1571 1158 1591 1162
rect 91 1157 1591 1158
rect 1597 1157 1598 1163
rect 96 1093 97 1099
rect 103 1098 1603 1099
rect 103 1094 111 1098
rect 115 1094 671 1098
rect 675 1094 703 1098
rect 707 1094 847 1098
rect 851 1094 1031 1098
rect 1035 1094 1055 1098
rect 1059 1094 1223 1098
rect 1227 1094 1407 1098
rect 1411 1094 1415 1098
rect 1419 1094 1567 1098
rect 1571 1094 1603 1098
rect 103 1093 1603 1094
rect 1609 1093 1610 1099
rect 84 1013 85 1019
rect 91 1018 1591 1019
rect 91 1014 111 1018
rect 115 1014 575 1018
rect 579 1014 671 1018
rect 675 1014 775 1018
rect 779 1014 847 1018
rect 851 1014 983 1018
rect 987 1014 1031 1018
rect 1035 1014 1191 1018
rect 1195 1014 1223 1018
rect 1227 1014 1407 1018
rect 1411 1014 1415 1018
rect 1419 1014 1567 1018
rect 1571 1014 1591 1018
rect 91 1013 1591 1014
rect 1597 1013 1598 1019
rect 96 941 97 947
rect 103 946 1603 947
rect 103 942 111 946
rect 115 942 407 946
rect 411 942 575 946
rect 579 942 735 946
rect 739 942 775 946
rect 779 942 983 946
rect 987 942 1063 946
rect 1067 942 1191 946
rect 1195 942 1399 946
rect 1403 942 1407 946
rect 1411 942 1567 946
rect 1571 942 1603 946
rect 103 941 1603 942
rect 1609 941 1610 947
rect 84 873 85 879
rect 91 878 1591 879
rect 91 874 111 878
rect 115 874 255 878
rect 259 874 407 878
rect 411 874 527 878
rect 531 874 735 878
rect 739 874 807 878
rect 811 874 1063 878
rect 1067 874 1095 878
rect 1099 874 1391 878
rect 1395 874 1399 878
rect 1403 874 1567 878
rect 1571 874 1591 878
rect 91 873 1591 874
rect 1597 873 1598 879
rect 96 789 97 795
rect 103 794 1603 795
rect 103 790 111 794
rect 115 790 167 794
rect 171 790 255 794
rect 259 790 383 794
rect 387 790 527 794
rect 531 790 623 794
rect 627 790 807 794
rect 811 790 871 794
rect 875 790 1095 794
rect 1099 790 1127 794
rect 1131 790 1391 794
rect 1395 790 1567 794
rect 1571 790 1603 794
rect 103 789 1603 790
rect 1609 789 1610 795
rect 84 705 85 711
rect 91 710 1591 711
rect 91 706 111 710
rect 115 706 167 710
rect 171 706 319 710
rect 323 706 383 710
rect 387 706 575 710
rect 579 706 623 710
rect 627 706 839 710
rect 843 706 871 710
rect 875 706 1119 710
rect 1123 706 1127 710
rect 1131 706 1391 710
rect 1395 706 1399 710
rect 1403 706 1567 710
rect 1571 706 1591 710
rect 91 705 1591 706
rect 1597 705 1598 711
rect 96 629 97 635
rect 103 634 1603 635
rect 103 630 111 634
rect 115 630 319 634
rect 323 630 575 634
rect 579 630 583 634
rect 587 630 727 634
rect 731 630 839 634
rect 843 630 887 634
rect 891 630 1055 634
rect 1059 630 1119 634
rect 1123 630 1231 634
rect 1235 630 1399 634
rect 1403 630 1407 634
rect 1411 630 1567 634
rect 1571 630 1603 634
rect 103 629 1603 630
rect 1609 629 1610 635
rect 84 545 85 551
rect 91 550 1591 551
rect 91 546 111 550
rect 115 546 583 550
rect 587 546 727 550
rect 731 546 759 550
rect 763 546 863 550
rect 867 546 887 550
rect 891 546 975 550
rect 979 546 1055 550
rect 1059 546 1087 550
rect 1091 546 1207 550
rect 1211 546 1231 550
rect 1235 546 1327 550
rect 1331 546 1407 550
rect 1411 546 1447 550
rect 1451 546 1567 550
rect 1571 546 1591 550
rect 91 545 1591 546
rect 1597 545 1598 551
rect 96 469 97 475
rect 103 474 1603 475
rect 103 470 111 474
rect 115 470 719 474
rect 723 470 759 474
rect 763 470 823 474
rect 827 470 863 474
rect 867 470 927 474
rect 931 470 975 474
rect 979 470 1031 474
rect 1035 470 1087 474
rect 1091 470 1135 474
rect 1139 470 1207 474
rect 1211 470 1239 474
rect 1243 470 1327 474
rect 1331 470 1351 474
rect 1355 470 1447 474
rect 1451 470 1463 474
rect 1467 470 1567 474
rect 1571 470 1603 474
rect 103 469 1603 470
rect 1609 469 1610 475
rect 84 377 85 383
rect 91 382 1591 383
rect 91 378 111 382
rect 115 378 511 382
rect 515 378 599 382
rect 603 378 687 382
rect 691 378 719 382
rect 723 378 775 382
rect 779 378 823 382
rect 827 378 927 382
rect 931 378 1031 382
rect 1035 378 1135 382
rect 1139 378 1239 382
rect 1243 378 1351 382
rect 1355 378 1463 382
rect 1467 378 1567 382
rect 1571 378 1591 382
rect 91 377 1591 378
rect 1597 377 1598 383
rect 96 305 97 311
rect 103 310 1603 311
rect 103 306 111 310
rect 115 306 375 310
rect 379 306 463 310
rect 467 306 511 310
rect 515 306 551 310
rect 555 306 599 310
rect 603 306 687 310
rect 691 306 775 310
rect 779 306 1567 310
rect 1571 306 1603 310
rect 103 305 1603 306
rect 1609 305 1610 311
rect 84 241 85 247
rect 91 246 1591 247
rect 91 242 111 246
rect 115 242 247 246
rect 251 242 335 246
rect 339 242 375 246
rect 379 242 423 246
rect 427 242 463 246
rect 467 242 551 246
rect 555 242 1567 246
rect 1571 242 1591 246
rect 91 241 1591 242
rect 1597 241 1598 247
rect 96 149 97 155
rect 103 154 1603 155
rect 103 150 111 154
rect 115 150 135 154
rect 139 150 223 154
rect 227 150 247 154
rect 251 150 311 154
rect 315 150 335 154
rect 339 150 399 154
rect 403 150 423 154
rect 427 150 487 154
rect 491 150 575 154
rect 579 150 1567 154
rect 1571 150 1603 154
rect 103 149 1603 150
rect 1609 149 1610 155
rect 84 85 85 91
rect 91 90 1591 91
rect 91 86 111 90
rect 115 86 135 90
rect 139 86 223 90
rect 227 86 311 90
rect 315 86 399 90
rect 403 86 487 90
rect 491 86 575 90
rect 579 86 1567 90
rect 1571 86 1591 90
rect 91 85 1591 86
rect 1597 85 1598 91
<< m5c >>
rect 97 1517 103 1523
rect 1603 1517 1609 1523
rect 85 1441 91 1447
rect 1591 1441 1597 1447
rect 97 1373 103 1379
rect 1603 1373 1609 1379
rect 85 1301 91 1307
rect 1591 1301 1597 1307
rect 97 1221 103 1227
rect 1603 1221 1609 1227
rect 85 1157 91 1163
rect 1591 1157 1597 1163
rect 97 1093 103 1099
rect 1603 1093 1609 1099
rect 85 1013 91 1019
rect 1591 1013 1597 1019
rect 97 941 103 947
rect 1603 941 1609 947
rect 85 873 91 879
rect 1591 873 1597 879
rect 97 789 103 795
rect 1603 789 1609 795
rect 85 705 91 711
rect 1591 705 1597 711
rect 97 629 103 635
rect 1603 629 1609 635
rect 85 545 91 551
rect 1591 545 1597 551
rect 97 469 103 475
rect 1603 469 1609 475
rect 85 377 91 383
rect 1591 377 1597 383
rect 97 305 103 311
rect 1603 305 1609 311
rect 85 241 91 247
rect 1591 241 1597 247
rect 97 149 103 155
rect 1603 149 1609 155
rect 85 85 91 91
rect 1591 85 1597 91
<< m5 >>
rect 84 1447 92 1656
rect 84 1441 85 1447
rect 91 1441 92 1447
rect 84 1307 92 1441
rect 84 1301 85 1307
rect 91 1301 92 1307
rect 84 1163 92 1301
rect 84 1157 85 1163
rect 91 1157 92 1163
rect 84 1019 92 1157
rect 84 1013 85 1019
rect 91 1013 92 1019
rect 84 879 92 1013
rect 84 873 85 879
rect 91 873 92 879
rect 84 711 92 873
rect 84 705 85 711
rect 91 705 92 711
rect 84 551 92 705
rect 84 545 85 551
rect 91 545 92 551
rect 84 383 92 545
rect 84 377 85 383
rect 91 377 92 383
rect 84 247 92 377
rect 84 241 85 247
rect 91 241 92 247
rect 84 91 92 241
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 1523 104 1656
rect 96 1517 97 1523
rect 103 1517 104 1523
rect 96 1379 104 1517
rect 96 1373 97 1379
rect 103 1373 104 1379
rect 96 1227 104 1373
rect 96 1221 97 1227
rect 103 1221 104 1227
rect 96 1099 104 1221
rect 96 1093 97 1099
rect 103 1093 104 1099
rect 96 947 104 1093
rect 96 941 97 947
rect 103 941 104 947
rect 96 795 104 941
rect 96 789 97 795
rect 103 789 104 795
rect 96 635 104 789
rect 96 629 97 635
rect 103 629 104 635
rect 96 475 104 629
rect 96 469 97 475
rect 103 469 104 475
rect 96 311 104 469
rect 96 305 97 311
rect 103 305 104 311
rect 96 155 104 305
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 1590 1447 1598 1656
rect 1590 1441 1591 1447
rect 1597 1441 1598 1447
rect 1590 1307 1598 1441
rect 1590 1301 1591 1307
rect 1597 1301 1598 1307
rect 1590 1163 1598 1301
rect 1590 1157 1591 1163
rect 1597 1157 1598 1163
rect 1590 1019 1598 1157
rect 1590 1013 1591 1019
rect 1597 1013 1598 1019
rect 1590 879 1598 1013
rect 1590 873 1591 879
rect 1597 873 1598 879
rect 1590 711 1598 873
rect 1590 705 1591 711
rect 1597 705 1598 711
rect 1590 551 1598 705
rect 1590 545 1591 551
rect 1597 545 1598 551
rect 1590 383 1598 545
rect 1590 377 1591 383
rect 1597 377 1598 383
rect 1590 247 1598 377
rect 1590 241 1591 247
rect 1597 241 1598 247
rect 1590 91 1598 241
rect 1590 85 1591 91
rect 1597 85 1598 91
rect 1590 72 1598 85
rect 1602 1523 1610 1656
rect 1602 1517 1603 1523
rect 1609 1517 1610 1523
rect 1602 1379 1610 1517
rect 1602 1373 1603 1379
rect 1609 1373 1610 1379
rect 1602 1227 1610 1373
rect 1602 1221 1603 1227
rect 1609 1221 1610 1227
rect 1602 1099 1610 1221
rect 1602 1093 1603 1099
rect 1609 1093 1610 1099
rect 1602 947 1610 1093
rect 1602 941 1603 947
rect 1609 941 1610 947
rect 1602 795 1610 941
rect 1602 789 1603 795
rect 1609 789 1610 795
rect 1602 635 1610 789
rect 1602 629 1603 635
rect 1609 629 1610 635
rect 1602 475 1610 629
rect 1602 469 1603 475
rect 1609 469 1610 475
rect 1602 311 1610 469
rect 1602 305 1603 311
rect 1609 305 1610 311
rect 1602 155 1610 305
rect 1602 149 1603 155
rect 1609 149 1610 155
rect 1602 72 1610 149
use _0_0cell_0_0gcelem3x0  celem_599_6_acx0
timestamp 1730767165
transform 1 0 128 0 1 88
box 8 4 79 60
use welltap_svt  __well_tap__0
timestamp 1730767165
transform 1 0 104 0 1 100
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0cell_0_0gcelem3x0  celem_599_6_acx0
timestamp 1730767165
transform 1 0 128 0 1 88
box 8 4 79 60
use welltap_svt  __well_tap__0
timestamp 1730767165
transform 1 0 104 0 1 100
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0cell_0_0gcelem3x0  celem_598_6_acx0
timestamp 1730767165
transform 1 0 216 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_598_6_acx0
timestamp 1730767165
transform 1 0 216 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_597_6_acx0
timestamp 1730767165
transform 1 0 304 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_597_6_acx0
timestamp 1730767165
transform 1 0 304 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_596_6_acx0
timestamp 1730767165
transform 1 0 392 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_596_6_acx0
timestamp 1730767165
transform 1 0 392 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_595_6_acx0
timestamp 1730767165
transform 1 0 480 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_595_6_acx0
timestamp 1730767165
transform 1 0 480 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_594_6_acx0
timestamp 1730767165
transform 1 0 568 0 1 88
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_594_6_acx0
timestamp 1730767165
transform 1 0 568 0 1 88
box 8 4 79 60
use welltap_svt  __well_tap__1
timestamp 1730767165
transform 1 0 1560 0 1 100
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730767165
transform 1 0 1560 0 1 100
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730767165
transform 1 0 104 0 -1 232
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730767165
transform 1 0 104 0 -1 232
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_592_6_acx0
timestamp 1730767165
transform 1 0 240 0 -1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_592_6_acx0
timestamp 1730767165
transform 1 0 240 0 -1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_591_6_acx0
timestamp 1730767165
transform 1 0 328 0 -1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_591_6_acx0
timestamp 1730767165
transform 1 0 328 0 -1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_593_6_acx0
timestamp 1730767165
transform 1 0 416 0 -1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_593_6_acx0
timestamp 1730767165
transform 1 0 416 0 -1 244
box 8 4 79 60
use welltap_svt  __well_tap__3
timestamp 1730767165
transform 1 0 1560 0 -1 232
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730767165
transform 1 0 1560 0 -1 232
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730767165
transform 1 0 104 0 1 256
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730767165
transform 1 0 104 0 1 256
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_590_6_acx0
timestamp 1730767165
transform 1 0 368 0 1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_590_6_acx0
timestamp 1730767165
transform 1 0 368 0 1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_587_6_acx0
timestamp 1730767165
transform 1 0 504 0 -1 380
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_589_6_acx0
timestamp 1730767165
transform 1 0 456 0 1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_587_6_acx0
timestamp 1730767165
transform 1 0 504 0 -1 380
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_589_6_acx0
timestamp 1730767165
transform 1 0 456 0 1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_586_6_acx0
timestamp 1730767165
transform 1 0 592 0 -1 380
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_588_6_acx0
timestamp 1730767165
transform 1 0 544 0 1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_586_6_acx0
timestamp 1730767165
transform 1 0 592 0 -1 380
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_588_6_acx0
timestamp 1730767165
transform 1 0 544 0 1 244
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_585_6_acx0
timestamp 1730767165
transform 1 0 680 0 -1 380
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_585_6_acx0
timestamp 1730767165
transform 1 0 680 0 -1 380
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_584_6_acx0
timestamp 1730767165
transform 1 0 768 0 -1 380
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_584_6_acx0
timestamp 1730767165
transform 1 0 768 0 -1 380
box 8 4 79 60
use welltap_svt  __well_tap__5
timestamp 1730767165
transform 1 0 1560 0 1 256
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730767165
transform 1 0 1560 0 1 256
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730767165
transform 1 0 104 0 -1 368
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730767165
transform 1 0 104 0 -1 368
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_583_6_acx0
timestamp 1730767165
transform 1 0 712 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_583_6_acx0
timestamp 1730767165
transform 1 0 712 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_582_6_acx0
timestamp 1730767165
transform 1 0 816 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_582_6_acx0
timestamp 1730767165
transform 1 0 816 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_581_6_acx0
timestamp 1730767165
transform 1 0 920 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_581_6_acx0
timestamp 1730767165
transform 1 0 920 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_580_6_acx0
timestamp 1730767165
transform 1 0 1024 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_580_6_acx0
timestamp 1730767165
transform 1 0 1024 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_520_6_acx0
timestamp 1730767165
transform 1 0 1128 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_520_6_acx0
timestamp 1730767165
transform 1 0 1128 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_519_6_acx0
timestamp 1730767165
transform 1 0 1232 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_519_6_acx0
timestamp 1730767165
transform 1 0 1232 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_518_6_acx0
timestamp 1730767165
transform 1 0 1344 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_518_6_acx0
timestamp 1730767165
transform 1 0 1344 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_517_6_acx0
timestamp 1730767165
transform 1 0 1456 0 1 408
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_517_6_acx0
timestamp 1730767165
transform 1 0 1456 0 1 408
box 8 4 79 60
use welltap_svt  __well_tap__7
timestamp 1730767165
transform 1 0 1560 0 -1 368
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730767165
transform 1 0 1560 0 -1 368
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730767165
transform 1 0 104 0 1 420
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730767165
transform 1 0 104 0 1 420
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_576_6_acx0
timestamp 1730767165
transform 1 0 752 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_576_6_acx0
timestamp 1730767165
transform 1 0 752 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_577_6_acx0
timestamp 1730767165
transform 1 0 856 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_577_6_acx0
timestamp 1730767165
transform 1 0 856 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_578_6_acx0
timestamp 1730767165
transform 1 0 968 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_578_6_acx0
timestamp 1730767165
transform 1 0 968 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_579_6_acx0
timestamp 1730767165
transform 1 0 1080 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_579_6_acx0
timestamp 1730767165
transform 1 0 1080 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_521_6_acx0
timestamp 1730767165
transform 1 0 1200 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_521_6_acx0
timestamp 1730767165
transform 1 0 1200 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_515_6_acx0
timestamp 1730767165
transform 1 0 1320 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_515_6_acx0
timestamp 1730767165
transform 1 0 1320 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_516_6_acx0
timestamp 1730767165
transform 1 0 1440 0 -1 548
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_516_6_acx0
timestamp 1730767165
transform 1 0 1440 0 -1 548
box 8 4 79 60
use welltap_svt  __well_tap__9
timestamp 1730767165
transform 1 0 1560 0 1 420
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730767165
transform 1 0 1560 0 1 420
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730767165
transform 1 0 104 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730767165
transform 1 0 104 0 1 580
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730767165
transform 1 0 104 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730767165
transform 1 0 104 0 1 580
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_575_6_acx0
timestamp 1730767165
transform 1 0 576 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_575_6_acx0
timestamp 1730767165
transform 1 0 576 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_574_6_acx0
timestamp 1730767165
transform 1 0 720 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_574_6_acx0
timestamp 1730767165
transform 1 0 720 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_573_6_acx0
timestamp 1730767165
transform 1 0 880 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_573_6_acx0
timestamp 1730767165
transform 1 0 880 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_572_6_acx0
timestamp 1730767165
transform 1 0 1048 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_572_6_acx0
timestamp 1730767165
transform 1 0 1048 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_522_6_acx0
timestamp 1730767165
transform 1 0 1224 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_522_6_acx0
timestamp 1730767165
transform 1 0 1224 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_514_6_acx0
timestamp 1730767165
transform 1 0 1400 0 1 568
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_514_6_acx0
timestamp 1730767165
transform 1 0 1400 0 1 568
box 8 4 79 60
use welltap_svt  __well_tap__11
timestamp 1730767165
transform 1 0 1560 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730767165
transform 1 0 1560 0 1 580
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730767165
transform 1 0 1560 0 -1 536
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730767165
transform 1 0 1560 0 1 580
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730767165
transform 1 0 104 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730767165
transform 1 0 104 0 -1 696
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_570_6_acx0
timestamp 1730767165
transform 1 0 312 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_570_6_acx0
timestamp 1730767165
transform 1 0 312 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_569_6_acx0
timestamp 1730767165
transform 1 0 568 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_569_6_acx0
timestamp 1730767165
transform 1 0 568 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_568_6_acx0
timestamp 1730767165
transform 1 0 832 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_568_6_acx0
timestamp 1730767165
transform 1 0 832 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_571_6_acx0
timestamp 1730767165
transform 1 0 1112 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_571_6_acx0
timestamp 1730767165
transform 1 0 1112 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_513_6_acx0
timestamp 1730767165
transform 1 0 1392 0 -1 708
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_513_6_acx0
timestamp 1730767165
transform 1 0 1392 0 -1 708
box 8 4 79 60
use welltap_svt  __well_tap__15
timestamp 1730767165
transform 1 0 1560 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730767165
transform 1 0 1560 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730767165
transform 1 0 104 0 1 740
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730767165
transform 1 0 104 0 1 740
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_564_6_acx0
timestamp 1730767165
transform 1 0 160 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_564_6_acx0
timestamp 1730767165
transform 1 0 160 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_565_6_acx0
timestamp 1730767165
transform 1 0 376 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_565_6_acx0
timestamp 1730767165
transform 1 0 376 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_566_6_acx0
timestamp 1730767165
transform 1 0 616 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_566_6_acx0
timestamp 1730767165
transform 1 0 616 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_567_6_acx0
timestamp 1730767165
transform 1 0 864 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_567_6_acx0
timestamp 1730767165
transform 1 0 864 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_523_6_acx0
timestamp 1730767165
transform 1 0 1120 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_523_6_acx0
timestamp 1730767165
transform 1 0 1120 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_512_6_acx0
timestamp 1730767165
transform 1 0 1384 0 1 728
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_512_6_acx0
timestamp 1730767165
transform 1 0 1384 0 1 728
box 8 4 79 60
use welltap_svt  __well_tap__17
timestamp 1730767165
transform 1 0 1560 0 1 740
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730767165
transform 1 0 1560 0 1 740
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730767165
transform 1 0 104 0 -1 864
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730767165
transform 1 0 104 0 -1 864
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_563_6_acx0
timestamp 1730767165
transform 1 0 248 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_563_6_acx0
timestamp 1730767165
transform 1 0 248 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_562_6_acx0
timestamp 1730767165
transform 1 0 520 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_562_6_acx0
timestamp 1730767165
transform 1 0 520 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_561_6_acx0
timestamp 1730767165
transform 1 0 800 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_561_6_acx0
timestamp 1730767165
transform 1 0 800 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_524_6_acx0
timestamp 1730767165
transform 1 0 1088 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_524_6_acx0
timestamp 1730767165
transform 1 0 1088 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_511_6_acx0
timestamp 1730767165
transform 1 0 1384 0 -1 876
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_511_6_acx0
timestamp 1730767165
transform 1 0 1384 0 -1 876
box 8 4 79 60
use welltap_svt  __well_tap__19
timestamp 1730767165
transform 1 0 1560 0 -1 864
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730767165
transform 1 0 1560 0 -1 864
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730767165
transform 1 0 104 0 1 892
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730767165
transform 1 0 104 0 1 892
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_558_6_acx0
timestamp 1730767165
transform 1 0 400 0 1 880
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_558_6_acx0
timestamp 1730767165
transform 1 0 400 0 1 880
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_559_6_acx0
timestamp 1730767165
transform 1 0 728 0 1 880
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_559_6_acx0
timestamp 1730767165
transform 1 0 728 0 1 880
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_560_6_acx0
timestamp 1730767165
transform 1 0 1056 0 1 880
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_560_6_acx0
timestamp 1730767165
transform 1 0 1056 0 1 880
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_510_6_acx0
timestamp 1730767165
transform 1 0 1392 0 1 880
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_510_6_acx0
timestamp 1730767165
transform 1 0 1392 0 1 880
box 8 4 79 60
use welltap_svt  __well_tap__21
timestamp 1730767165
transform 1 0 1560 0 1 892
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730767165
transform 1 0 1560 0 1 892
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730767165
transform 1 0 104 0 -1 1004
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730767165
transform 1 0 104 0 -1 1004
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_557_6_acx0
timestamp 1730767165
transform 1 0 568 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_557_6_acx0
timestamp 1730767165
transform 1 0 568 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_556_6_acx0
timestamp 1730767165
transform 1 0 768 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_556_6_acx0
timestamp 1730767165
transform 1 0 768 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_555_6_acx0
timestamp 1730767165
transform 1 0 976 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_555_6_acx0
timestamp 1730767165
transform 1 0 976 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_525_6_acx0
timestamp 1730767165
transform 1 0 1184 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_525_6_acx0
timestamp 1730767165
transform 1 0 1184 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_59_6_acx0
timestamp 1730767165
transform 1 0 1400 0 -1 1016
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_59_6_acx0
timestamp 1730767165
transform 1 0 1400 0 -1 1016
box 8 4 79 60
use welltap_svt  __well_tap__23
timestamp 1730767165
transform 1 0 1560 0 -1 1004
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730767165
transform 1 0 1560 0 -1 1004
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730767165
transform 1 0 104 0 1 1044
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730767165
transform 1 0 104 0 1 1044
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_554_6_acx0
timestamp 1730767165
transform 1 0 664 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_554_6_acx0
timestamp 1730767165
transform 1 0 664 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_550_6_acx0
timestamp 1730767165
transform 1 0 696 0 -1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_550_6_acx0
timestamp 1730767165
transform 1 0 696 0 -1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_553_6_acx0
timestamp 1730767165
transform 1 0 840 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_553_6_acx0
timestamp 1730767165
transform 1 0 840 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_552_6_acx0
timestamp 1730767165
transform 1 0 1024 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_552_6_acx0
timestamp 1730767165
transform 1 0 1024 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_551_6_acx0
timestamp 1730767165
transform 1 0 1048 0 -1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_551_6_acx0
timestamp 1730767165
transform 1 0 1048 0 -1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_526_6_acx0
timestamp 1730767165
transform 1 0 1216 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_526_6_acx0
timestamp 1730767165
transform 1 0 1216 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_57_6_acx0
timestamp 1730767165
transform 1 0 1400 0 -1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_58_6_acx0
timestamp 1730767165
transform 1 0 1408 0 1 1032
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_57_6_acx0
timestamp 1730767165
transform 1 0 1400 0 -1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_58_6_acx0
timestamp 1730767165
transform 1 0 1408 0 1 1032
box 8 4 79 60
use welltap_svt  __well_tap__25
timestamp 1730767165
transform 1 0 1560 0 1 1044
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730767165
transform 1 0 1560 0 1 1044
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730767165
transform 1 0 104 0 -1 1148
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730767165
transform 1 0 104 0 1 1172
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730767165
transform 1 0 104 0 -1 1148
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730767165
transform 1 0 104 0 1 1172
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_549_6_acx0
timestamp 1730767165
transform 1 0 560 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_549_6_acx0
timestamp 1730767165
transform 1 0 560 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_548_6_acx0
timestamp 1730767165
transform 1 0 760 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_548_6_acx0
timestamp 1730767165
transform 1 0 760 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_547_6_acx0
timestamp 1730767165
transform 1 0 960 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_547_6_acx0
timestamp 1730767165
transform 1 0 960 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_527_6_acx0
timestamp 1730767165
transform 1 0 1168 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_527_6_acx0
timestamp 1730767165
transform 1 0 1168 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_56_6_acx0
timestamp 1730767165
transform 1 0 1384 0 1 1160
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_56_6_acx0
timestamp 1730767165
transform 1 0 1384 0 1 1160
box 8 4 79 60
use welltap_svt  __well_tap__27
timestamp 1730767165
transform 1 0 1560 0 -1 1148
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730767165
transform 1 0 1560 0 1 1172
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730767165
transform 1 0 1560 0 -1 1148
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730767165
transform 1 0 1560 0 1 1172
box 8 4 12 24
use welltap_svt  __well_tap__30
timestamp 1730767165
transform 1 0 104 0 -1 1292
box 8 4 12 24
use welltap_svt  __well_tap__30
timestamp 1730767165
transform 1 0 104 0 -1 1292
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_545_6_acx0
timestamp 1730767165
transform 1 0 512 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_545_6_acx0
timestamp 1730767165
transform 1 0 512 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_546_6_acx0
timestamp 1730767165
transform 1 0 736 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_546_6_acx0
timestamp 1730767165
transform 1 0 736 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_528_6_acx0
timestamp 1730767165
transform 1 0 968 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_528_6_acx0
timestamp 1730767165
transform 1 0 968 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_54_6_acx0
timestamp 1730767165
transform 1 0 1200 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_54_6_acx0
timestamp 1730767165
transform 1 0 1200 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_55_6_acx0
timestamp 1730767165
transform 1 0 1432 0 -1 1304
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_55_6_acx0
timestamp 1730767165
transform 1 0 1432 0 -1 1304
box 8 4 79 60
use welltap_svt  __well_tap__31
timestamp 1730767165
transform 1 0 1560 0 -1 1292
box 8 4 12 24
use welltap_svt  __well_tap__31
timestamp 1730767165
transform 1 0 1560 0 -1 1292
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730767165
transform 1 0 104 0 1 1324
box 8 4 12 24
use welltap_svt  __well_tap__32
timestamp 1730767165
transform 1 0 104 0 1 1324
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_544_6_acx0
timestamp 1730767165
transform 1 0 464 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_544_6_acx0
timestamp 1730767165
transform 1 0 464 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_543_6_acx0
timestamp 1730767165
transform 1 0 688 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_543_6_acx0
timestamp 1730767165
transform 1 0 688 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_529_6_acx0
timestamp 1730767165
transform 1 0 912 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_529_6_acx0
timestamp 1730767165
transform 1 0 912 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_530_6_acx0
timestamp 1730767165
transform 1 0 1144 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_530_6_acx0
timestamp 1730767165
transform 1 0 1144 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_53_6_acx0
timestamp 1730767165
transform 1 0 1384 0 1 1312
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_53_6_acx0
timestamp 1730767165
transform 1 0 1384 0 1 1312
box 8 4 79 60
use welltap_svt  __well_tap__33
timestamp 1730767165
transform 1 0 1560 0 1 1324
box 8 4 12 24
use welltap_svt  __well_tap__33
timestamp 1730767165
transform 1 0 1560 0 1 1324
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730767165
transform 1 0 104 0 -1 1432
box 8 4 12 24
use welltap_svt  __well_tap__34
timestamp 1730767165
transform 1 0 104 0 -1 1432
box 8 4 12 24
use _0_0cell_0_0gcelem3x0  celem_539_6_acx0
timestamp 1730767165
transform 1 0 392 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_540_6_acx0
timestamp 1730767165
transform 1 0 416 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_539_6_acx0
timestamp 1730767165
transform 1 0 392 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_540_6_acx0
timestamp 1730767165
transform 1 0 416 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_538_6_acx0
timestamp 1730767165
transform 1 0 480 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_538_6_acx0
timestamp 1730767165
transform 1 0 480 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_537_6_acx0
timestamp 1730767165
transform 1 0 568 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_537_6_acx0
timestamp 1730767165
transform 1 0 568 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_536_6_acx0
timestamp 1730767165
transform 1 0 664 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_541_6_acx0
timestamp 1730767165
transform 1 0 648 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_536_6_acx0
timestamp 1730767165
transform 1 0 664 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_541_6_acx0
timestamp 1730767165
transform 1 0 648 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_535_6_acx0
timestamp 1730767165
transform 1 0 776 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_535_6_acx0
timestamp 1730767165
transform 1 0 776 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_534_6_acx0
timestamp 1730767165
transform 1 0 896 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_542_6_acx0
timestamp 1730767165
transform 1 0 888 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_534_6_acx0
timestamp 1730767165
transform 1 0 896 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_542_6_acx0
timestamp 1730767165
transform 1 0 888 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_533_6_acx0
timestamp 1730767165
transform 1 0 1024 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_533_6_acx0
timestamp 1730767165
transform 1 0 1024 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_531_6_acx0
timestamp 1730767165
transform 1 0 1136 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_532_6_acx0
timestamp 1730767165
transform 1 0 1160 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_531_6_acx0
timestamp 1730767165
transform 1 0 1136 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_532_6_acx0
timestamp 1730767165
transform 1 0 1160 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_50_6_acx0
timestamp 1730767165
transform 1 0 1296 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_50_6_acx0
timestamp 1730767165
transform 1 0 1296 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_51_6_acx0
timestamp 1730767165
transform 1 0 1440 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_52_6_acx0
timestamp 1730767165
transform 1 0 1392 0 -1 1444
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_51_6_acx0
timestamp 1730767165
transform 1 0 1440 0 1 1456
box 8 4 79 60
use _0_0cell_0_0gcelem3x0  celem_52_6_acx0
timestamp 1730767165
transform 1 0 1392 0 -1 1444
box 8 4 79 60
use welltap_svt  __well_tap__35
timestamp 1730767165
transform 1 0 1560 0 -1 1432
box 8 4 12 24
use welltap_svt  __well_tap__35
timestamp 1730767165
transform 1 0 1560 0 -1 1432
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730767165
transform 1 0 104 0 1 1468
box 8 4 12 24
use welltap_svt  __well_tap__36
timestamp 1730767165
transform 1 0 104 0 1 1468
box 8 4 12 24
use welltap_svt  __well_tap__37
timestamp 1730767165
transform 1 0 1560 0 1 1468
box 8 4 12 24
use welltap_svt  __well_tap__37
timestamp 1730767165
transform 1 0 1560 0 1 1468
box 8 4 12 24
<< end >>
