magic
tech sky130l
timestamp 1729431977
<< ndiffusion >>
rect 8 12 13 16
rect 8 9 9 12
rect 12 9 13 12
rect 8 6 13 9
rect 15 6 20 16
rect 22 14 27 16
rect 22 11 23 14
rect 26 11 27 14
rect 22 10 27 11
rect 29 15 34 16
rect 29 12 30 15
rect 33 12 34 15
rect 29 10 34 12
rect 22 6 26 10
<< ndc >>
rect 9 9 12 12
rect 23 11 26 14
rect 30 12 33 15
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 27 10 29 16
<< pdiffusion >>
rect 8 28 13 31
rect 8 25 9 28
rect 12 25 13 28
rect 8 23 13 25
rect 15 23 20 31
rect 22 28 27 31
rect 22 25 23 28
rect 26 25 27 28
rect 22 23 27 25
rect 29 28 34 31
rect 29 25 30 28
rect 33 25 34 28
rect 29 23 34 25
<< pdc >>
rect 9 25 12 28
rect 23 25 26 28
rect 30 25 33 28
<< ptransistor >>
rect 13 23 15 31
rect 20 23 22 31
rect 27 23 29 31
<< polysilicon >>
rect 13 40 19 41
rect 13 37 15 40
rect 18 37 19 40
rect 13 36 19 37
rect 13 31 15 36
rect 20 31 22 33
rect 27 31 29 33
rect 13 16 15 23
rect 20 16 22 23
rect 27 16 29 23
rect 27 8 29 10
rect 27 7 36 8
rect 13 4 15 6
rect 20 1 22 6
rect 27 4 32 7
rect 35 4 36 7
rect 31 3 36 4
rect 16 0 22 1
rect 16 -3 17 0
rect 20 -3 22 0
rect 16 -4 22 -3
<< pc >>
rect 15 37 18 40
rect 32 4 35 7
rect 17 -3 20 0
<< m1 >>
rect 15 40 20 41
rect 18 37 20 40
rect 15 36 20 37
rect 8 28 12 36
rect 16 32 20 36
rect 32 29 36 36
rect 8 25 9 28
rect 8 24 12 25
rect 22 28 26 29
rect 22 25 23 28
rect 22 24 26 25
rect 30 28 36 29
rect 33 25 36 28
rect 30 24 36 25
rect 32 16 36 24
rect 30 15 36 16
rect 23 14 27 15
rect 8 12 12 13
rect 8 9 9 12
rect 26 11 27 14
rect 33 12 36 15
rect 30 11 36 12
rect 23 10 27 11
rect 8 7 12 9
rect 24 8 27 10
rect 8 4 9 7
rect 16 0 20 8
rect 24 4 28 8
rect 32 7 36 8
rect 35 4 36 7
rect 32 3 36 4
rect 16 -3 17 0
rect 16 -4 20 -3
<< m2c >>
rect 9 25 12 28
rect 23 25 26 28
rect 9 4 12 7
rect 32 4 35 7
<< m2 >>
rect 8 28 27 29
rect 8 25 9 28
rect 12 25 23 28
rect 26 25 27 28
rect 8 24 27 25
rect 8 7 36 8
rect 8 4 9 7
rect 12 4 32 7
rect 35 4 36 7
rect 8 3 36 4
<< labels >>
rlabel ndiffusion 30 11 30 11 3 Y
rlabel polysilicon 28 22 28 22 3 _Y
rlabel pdiffusion 30 24 30 24 3 Y
rlabel pdiffusion 23 24 23 24 3 Vdd
rlabel polysilicon 21 17 21 17 3 A
rlabel polysilicon 21 22 21 22 3 A
rlabel pdiffusion 16 24 16 24 3 _Y
rlabel polysilicon 14 17 14 17 3 B
rlabel polysilicon 14 22 14 22 3 B
rlabel ndiffusion 9 7 9 7 3 _Y
rlabel m1 17 33 17 33 3 B
port 3 e
rlabel m1 9 33 9 33 4 Vdd
rlabel m1 34 33 34 33 6 Y
rlabel m1 18 2 18 2 1 A
rlabel m1 25 9 25 9 1 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel polysilicon 28 17 28 17 3 _Y
<< end >>
