magic
tech sky130l
timestamp 1731220447
<< m2 >>
rect 1974 5729 1980 5730
rect 3798 5729 3804 5730
rect 1974 5725 1975 5729
rect 1979 5725 1980 5729
rect 1974 5724 1980 5725
rect 2374 5728 2380 5729
rect 2374 5724 2375 5728
rect 2379 5724 2380 5728
rect 2374 5723 2380 5724
rect 2510 5728 2516 5729
rect 2510 5724 2511 5728
rect 2515 5724 2516 5728
rect 2510 5723 2516 5724
rect 2654 5728 2660 5729
rect 2654 5724 2655 5728
rect 2659 5724 2660 5728
rect 2654 5723 2660 5724
rect 2806 5728 2812 5729
rect 2806 5724 2807 5728
rect 2811 5724 2812 5728
rect 2806 5723 2812 5724
rect 2958 5728 2964 5729
rect 2958 5724 2959 5728
rect 2963 5724 2964 5728
rect 2958 5723 2964 5724
rect 3118 5728 3124 5729
rect 3118 5724 3119 5728
rect 3123 5724 3124 5728
rect 3798 5725 3799 5729
rect 3803 5725 3804 5729
rect 3798 5724 3804 5725
rect 3118 5723 3124 5724
rect 2346 5713 2352 5714
rect 1974 5712 1980 5713
rect 1974 5708 1975 5712
rect 1979 5708 1980 5712
rect 2346 5709 2347 5713
rect 2351 5709 2352 5713
rect 2346 5708 2352 5709
rect 2482 5713 2488 5714
rect 2482 5709 2483 5713
rect 2487 5709 2488 5713
rect 2482 5708 2488 5709
rect 2626 5713 2632 5714
rect 2626 5709 2627 5713
rect 2631 5709 2632 5713
rect 2626 5708 2632 5709
rect 2778 5713 2784 5714
rect 2778 5709 2779 5713
rect 2783 5709 2784 5713
rect 2778 5708 2784 5709
rect 2930 5713 2936 5714
rect 2930 5709 2931 5713
rect 2935 5709 2936 5713
rect 2930 5708 2936 5709
rect 3090 5713 3096 5714
rect 3090 5709 3091 5713
rect 3095 5709 3096 5713
rect 3090 5708 3096 5709
rect 3798 5712 3804 5713
rect 3798 5708 3799 5712
rect 3803 5708 3804 5712
rect 1974 5707 1980 5708
rect 3798 5707 3804 5708
rect 110 5689 116 5690
rect 1934 5689 1940 5690
rect 110 5685 111 5689
rect 115 5685 116 5689
rect 110 5684 116 5685
rect 158 5688 164 5689
rect 158 5684 159 5688
rect 163 5684 164 5688
rect 158 5683 164 5684
rect 294 5688 300 5689
rect 294 5684 295 5688
rect 299 5684 300 5688
rect 294 5683 300 5684
rect 430 5688 436 5689
rect 430 5684 431 5688
rect 435 5684 436 5688
rect 430 5683 436 5684
rect 566 5688 572 5689
rect 566 5684 567 5688
rect 571 5684 572 5688
rect 566 5683 572 5684
rect 702 5688 708 5689
rect 702 5684 703 5688
rect 707 5684 708 5688
rect 702 5683 708 5684
rect 838 5688 844 5689
rect 838 5684 839 5688
rect 843 5684 844 5688
rect 838 5683 844 5684
rect 974 5688 980 5689
rect 974 5684 975 5688
rect 979 5684 980 5688
rect 1934 5685 1935 5689
rect 1939 5685 1940 5689
rect 1934 5684 1940 5685
rect 974 5683 980 5684
rect 130 5673 136 5674
rect 110 5672 116 5673
rect 110 5668 111 5672
rect 115 5668 116 5672
rect 130 5669 131 5673
rect 135 5669 136 5673
rect 130 5668 136 5669
rect 266 5673 272 5674
rect 266 5669 267 5673
rect 271 5669 272 5673
rect 266 5668 272 5669
rect 402 5673 408 5674
rect 402 5669 403 5673
rect 407 5669 408 5673
rect 402 5668 408 5669
rect 538 5673 544 5674
rect 538 5669 539 5673
rect 543 5669 544 5673
rect 538 5668 544 5669
rect 674 5673 680 5674
rect 674 5669 675 5673
rect 679 5669 680 5673
rect 674 5668 680 5669
rect 810 5673 816 5674
rect 810 5669 811 5673
rect 815 5669 816 5673
rect 810 5668 816 5669
rect 946 5673 952 5674
rect 946 5669 947 5673
rect 951 5669 952 5673
rect 946 5668 952 5669
rect 1934 5672 1940 5673
rect 1934 5668 1935 5672
rect 1939 5668 1940 5672
rect 110 5667 116 5668
rect 1934 5667 1940 5668
rect 3838 5653 3844 5654
rect 5662 5653 5668 5654
rect 3838 5649 3839 5653
rect 3843 5649 3844 5653
rect 3838 5648 3844 5649
rect 4334 5652 4340 5653
rect 4334 5648 4335 5652
rect 4339 5648 4340 5652
rect 4334 5647 4340 5648
rect 4470 5652 4476 5653
rect 4470 5648 4471 5652
rect 4475 5648 4476 5652
rect 4470 5647 4476 5648
rect 4606 5652 4612 5653
rect 4606 5648 4607 5652
rect 4611 5648 4612 5652
rect 4606 5647 4612 5648
rect 4742 5652 4748 5653
rect 4742 5648 4743 5652
rect 4747 5648 4748 5652
rect 4742 5647 4748 5648
rect 4878 5652 4884 5653
rect 4878 5648 4879 5652
rect 4883 5648 4884 5652
rect 4878 5647 4884 5648
rect 5014 5652 5020 5653
rect 5014 5648 5015 5652
rect 5019 5648 5020 5652
rect 5662 5649 5663 5653
rect 5667 5649 5668 5653
rect 5662 5648 5668 5649
rect 5014 5647 5020 5648
rect 4306 5637 4312 5638
rect 3838 5636 3844 5637
rect 3838 5632 3839 5636
rect 3843 5632 3844 5636
rect 4306 5633 4307 5637
rect 4311 5633 4312 5637
rect 4306 5632 4312 5633
rect 4442 5637 4448 5638
rect 4442 5633 4443 5637
rect 4447 5633 4448 5637
rect 4442 5632 4448 5633
rect 4578 5637 4584 5638
rect 4578 5633 4579 5637
rect 4583 5633 4584 5637
rect 4578 5632 4584 5633
rect 4714 5637 4720 5638
rect 4714 5633 4715 5637
rect 4719 5633 4720 5637
rect 4714 5632 4720 5633
rect 4850 5637 4856 5638
rect 4850 5633 4851 5637
rect 4855 5633 4856 5637
rect 4850 5632 4856 5633
rect 4986 5637 4992 5638
rect 4986 5633 4987 5637
rect 4991 5633 4992 5637
rect 4986 5632 4992 5633
rect 5662 5636 5668 5637
rect 5662 5632 5663 5636
rect 5667 5632 5668 5636
rect 3838 5631 3844 5632
rect 5662 5631 5668 5632
rect 1974 5580 1980 5581
rect 3798 5580 3804 5581
rect 1974 5576 1975 5580
rect 1979 5576 1980 5580
rect 1974 5575 1980 5576
rect 1994 5579 2000 5580
rect 1994 5575 1995 5579
rect 1999 5575 2000 5579
rect 1994 5574 2000 5575
rect 2202 5579 2208 5580
rect 2202 5575 2203 5579
rect 2207 5575 2208 5579
rect 2202 5574 2208 5575
rect 2426 5579 2432 5580
rect 2426 5575 2427 5579
rect 2431 5575 2432 5579
rect 2426 5574 2432 5575
rect 2650 5579 2656 5580
rect 2650 5575 2651 5579
rect 2655 5575 2656 5579
rect 2650 5574 2656 5575
rect 2866 5579 2872 5580
rect 2866 5575 2867 5579
rect 2871 5575 2872 5579
rect 2866 5574 2872 5575
rect 3074 5579 3080 5580
rect 3074 5575 3075 5579
rect 3079 5575 3080 5579
rect 3074 5574 3080 5575
rect 3274 5579 3280 5580
rect 3274 5575 3275 5579
rect 3279 5575 3280 5579
rect 3274 5574 3280 5575
rect 3474 5579 3480 5580
rect 3474 5575 3475 5579
rect 3479 5575 3480 5579
rect 3474 5574 3480 5575
rect 3650 5579 3656 5580
rect 3650 5575 3651 5579
rect 3655 5575 3656 5579
rect 3798 5576 3799 5580
rect 3803 5576 3804 5580
rect 3798 5575 3804 5576
rect 3650 5574 3656 5575
rect 2022 5564 2028 5565
rect 1974 5563 1980 5564
rect 1974 5559 1975 5563
rect 1979 5559 1980 5563
rect 2022 5560 2023 5564
rect 2027 5560 2028 5564
rect 2022 5559 2028 5560
rect 2230 5564 2236 5565
rect 2230 5560 2231 5564
rect 2235 5560 2236 5564
rect 2230 5559 2236 5560
rect 2454 5564 2460 5565
rect 2454 5560 2455 5564
rect 2459 5560 2460 5564
rect 2454 5559 2460 5560
rect 2678 5564 2684 5565
rect 2678 5560 2679 5564
rect 2683 5560 2684 5564
rect 2678 5559 2684 5560
rect 2894 5564 2900 5565
rect 2894 5560 2895 5564
rect 2899 5560 2900 5564
rect 2894 5559 2900 5560
rect 3102 5564 3108 5565
rect 3102 5560 3103 5564
rect 3107 5560 3108 5564
rect 3102 5559 3108 5560
rect 3302 5564 3308 5565
rect 3302 5560 3303 5564
rect 3307 5560 3308 5564
rect 3302 5559 3308 5560
rect 3502 5564 3508 5565
rect 3502 5560 3503 5564
rect 3507 5560 3508 5564
rect 3502 5559 3508 5560
rect 3678 5564 3684 5565
rect 3678 5560 3679 5564
rect 3683 5560 3684 5564
rect 3678 5559 3684 5560
rect 3798 5563 3804 5564
rect 3798 5559 3799 5563
rect 3803 5559 3804 5563
rect 1974 5558 1980 5559
rect 3798 5558 3804 5559
rect 110 5512 116 5513
rect 1934 5512 1940 5513
rect 110 5508 111 5512
rect 115 5508 116 5512
rect 110 5507 116 5508
rect 618 5511 624 5512
rect 618 5507 619 5511
rect 623 5507 624 5511
rect 618 5506 624 5507
rect 754 5511 760 5512
rect 754 5507 755 5511
rect 759 5507 760 5511
rect 754 5506 760 5507
rect 898 5511 904 5512
rect 898 5507 899 5511
rect 903 5507 904 5511
rect 898 5506 904 5507
rect 1050 5511 1056 5512
rect 1050 5507 1051 5511
rect 1055 5507 1056 5511
rect 1050 5506 1056 5507
rect 1202 5511 1208 5512
rect 1202 5507 1203 5511
rect 1207 5507 1208 5511
rect 1202 5506 1208 5507
rect 1354 5511 1360 5512
rect 1354 5507 1355 5511
rect 1359 5507 1360 5511
rect 1354 5506 1360 5507
rect 1506 5511 1512 5512
rect 1506 5507 1507 5511
rect 1511 5507 1512 5511
rect 1506 5506 1512 5507
rect 1650 5511 1656 5512
rect 1650 5507 1651 5511
rect 1655 5507 1656 5511
rect 1650 5506 1656 5507
rect 1786 5511 1792 5512
rect 1786 5507 1787 5511
rect 1791 5507 1792 5511
rect 1934 5508 1935 5512
rect 1939 5508 1940 5512
rect 1934 5507 1940 5508
rect 1786 5506 1792 5507
rect 1974 5505 1980 5506
rect 3798 5505 3804 5506
rect 1974 5501 1975 5505
rect 1979 5501 1980 5505
rect 1974 5500 1980 5501
rect 2950 5504 2956 5505
rect 2950 5500 2951 5504
rect 2955 5500 2956 5504
rect 2950 5499 2956 5500
rect 3102 5504 3108 5505
rect 3102 5500 3103 5504
rect 3107 5500 3108 5504
rect 3102 5499 3108 5500
rect 3254 5504 3260 5505
rect 3254 5500 3255 5504
rect 3259 5500 3260 5504
rect 3254 5499 3260 5500
rect 3414 5504 3420 5505
rect 3414 5500 3415 5504
rect 3419 5500 3420 5504
rect 3798 5501 3799 5505
rect 3803 5501 3804 5505
rect 3798 5500 3804 5501
rect 3838 5504 3844 5505
rect 5662 5504 5668 5505
rect 3838 5500 3839 5504
rect 3843 5500 3844 5504
rect 3414 5499 3420 5500
rect 3838 5499 3844 5500
rect 4210 5503 4216 5504
rect 4210 5499 4211 5503
rect 4215 5499 4216 5503
rect 4210 5498 4216 5499
rect 4402 5503 4408 5504
rect 4402 5499 4403 5503
rect 4407 5499 4408 5503
rect 4402 5498 4408 5499
rect 4594 5503 4600 5504
rect 4594 5499 4595 5503
rect 4599 5499 4600 5503
rect 4594 5498 4600 5499
rect 4794 5503 4800 5504
rect 4794 5499 4795 5503
rect 4799 5499 4800 5503
rect 4794 5498 4800 5499
rect 4994 5503 5000 5504
rect 4994 5499 4995 5503
rect 4999 5499 5000 5503
rect 4994 5498 5000 5499
rect 5194 5503 5200 5504
rect 5194 5499 5195 5503
rect 5199 5499 5200 5503
rect 5662 5500 5663 5504
rect 5667 5500 5668 5504
rect 5662 5499 5668 5500
rect 5194 5498 5200 5499
rect 646 5496 652 5497
rect 110 5495 116 5496
rect 110 5491 111 5495
rect 115 5491 116 5495
rect 646 5492 647 5496
rect 651 5492 652 5496
rect 646 5491 652 5492
rect 782 5496 788 5497
rect 782 5492 783 5496
rect 787 5492 788 5496
rect 782 5491 788 5492
rect 926 5496 932 5497
rect 926 5492 927 5496
rect 931 5492 932 5496
rect 926 5491 932 5492
rect 1078 5496 1084 5497
rect 1078 5492 1079 5496
rect 1083 5492 1084 5496
rect 1078 5491 1084 5492
rect 1230 5496 1236 5497
rect 1230 5492 1231 5496
rect 1235 5492 1236 5496
rect 1230 5491 1236 5492
rect 1382 5496 1388 5497
rect 1382 5492 1383 5496
rect 1387 5492 1388 5496
rect 1382 5491 1388 5492
rect 1534 5496 1540 5497
rect 1534 5492 1535 5496
rect 1539 5492 1540 5496
rect 1534 5491 1540 5492
rect 1678 5496 1684 5497
rect 1678 5492 1679 5496
rect 1683 5492 1684 5496
rect 1678 5491 1684 5492
rect 1814 5496 1820 5497
rect 1814 5492 1815 5496
rect 1819 5492 1820 5496
rect 1814 5491 1820 5492
rect 1934 5495 1940 5496
rect 1934 5491 1935 5495
rect 1939 5491 1940 5495
rect 110 5490 116 5491
rect 1934 5490 1940 5491
rect 2922 5489 2928 5490
rect 1974 5488 1980 5489
rect 1974 5484 1975 5488
rect 1979 5484 1980 5488
rect 2922 5485 2923 5489
rect 2927 5485 2928 5489
rect 2922 5484 2928 5485
rect 3074 5489 3080 5490
rect 3074 5485 3075 5489
rect 3079 5485 3080 5489
rect 3074 5484 3080 5485
rect 3226 5489 3232 5490
rect 3226 5485 3227 5489
rect 3231 5485 3232 5489
rect 3226 5484 3232 5485
rect 3386 5489 3392 5490
rect 3386 5485 3387 5489
rect 3391 5485 3392 5489
rect 3386 5484 3392 5485
rect 3798 5488 3804 5489
rect 4238 5488 4244 5489
rect 3798 5484 3799 5488
rect 3803 5484 3804 5488
rect 1974 5483 1980 5484
rect 3798 5483 3804 5484
rect 3838 5487 3844 5488
rect 3838 5483 3839 5487
rect 3843 5483 3844 5487
rect 4238 5484 4239 5488
rect 4243 5484 4244 5488
rect 4238 5483 4244 5484
rect 4430 5488 4436 5489
rect 4430 5484 4431 5488
rect 4435 5484 4436 5488
rect 4430 5483 4436 5484
rect 4622 5488 4628 5489
rect 4622 5484 4623 5488
rect 4627 5484 4628 5488
rect 4622 5483 4628 5484
rect 4822 5488 4828 5489
rect 4822 5484 4823 5488
rect 4827 5484 4828 5488
rect 4822 5483 4828 5484
rect 5022 5488 5028 5489
rect 5022 5484 5023 5488
rect 5027 5484 5028 5488
rect 5022 5483 5028 5484
rect 5222 5488 5228 5489
rect 5222 5484 5223 5488
rect 5227 5484 5228 5488
rect 5222 5483 5228 5484
rect 5662 5487 5668 5488
rect 5662 5483 5663 5487
rect 5667 5483 5668 5487
rect 3838 5482 3844 5483
rect 5662 5482 5668 5483
rect 110 5429 116 5430
rect 1934 5429 1940 5430
rect 110 5425 111 5429
rect 115 5425 116 5429
rect 110 5424 116 5425
rect 590 5428 596 5429
rect 590 5424 591 5428
rect 595 5424 596 5428
rect 590 5423 596 5424
rect 726 5428 732 5429
rect 726 5424 727 5428
rect 731 5424 732 5428
rect 726 5423 732 5424
rect 862 5428 868 5429
rect 862 5424 863 5428
rect 867 5424 868 5428
rect 862 5423 868 5424
rect 998 5428 1004 5429
rect 998 5424 999 5428
rect 1003 5424 1004 5428
rect 998 5423 1004 5424
rect 1134 5428 1140 5429
rect 1134 5424 1135 5428
rect 1139 5424 1140 5428
rect 1134 5423 1140 5424
rect 1270 5428 1276 5429
rect 1270 5424 1271 5428
rect 1275 5424 1276 5428
rect 1270 5423 1276 5424
rect 1406 5428 1412 5429
rect 1406 5424 1407 5428
rect 1411 5424 1412 5428
rect 1406 5423 1412 5424
rect 1542 5428 1548 5429
rect 1542 5424 1543 5428
rect 1547 5424 1548 5428
rect 1542 5423 1548 5424
rect 1678 5428 1684 5429
rect 1678 5424 1679 5428
rect 1683 5424 1684 5428
rect 1678 5423 1684 5424
rect 1814 5428 1820 5429
rect 1814 5424 1815 5428
rect 1819 5424 1820 5428
rect 1934 5425 1935 5429
rect 1939 5425 1940 5429
rect 1934 5424 1940 5425
rect 1814 5423 1820 5424
rect 562 5413 568 5414
rect 110 5412 116 5413
rect 110 5408 111 5412
rect 115 5408 116 5412
rect 562 5409 563 5413
rect 567 5409 568 5413
rect 562 5408 568 5409
rect 698 5413 704 5414
rect 698 5409 699 5413
rect 703 5409 704 5413
rect 698 5408 704 5409
rect 834 5413 840 5414
rect 834 5409 835 5413
rect 839 5409 840 5413
rect 834 5408 840 5409
rect 970 5413 976 5414
rect 970 5409 971 5413
rect 975 5409 976 5413
rect 970 5408 976 5409
rect 1106 5413 1112 5414
rect 1106 5409 1107 5413
rect 1111 5409 1112 5413
rect 1106 5408 1112 5409
rect 1242 5413 1248 5414
rect 1242 5409 1243 5413
rect 1247 5409 1248 5413
rect 1242 5408 1248 5409
rect 1378 5413 1384 5414
rect 1378 5409 1379 5413
rect 1383 5409 1384 5413
rect 1378 5408 1384 5409
rect 1514 5413 1520 5414
rect 1514 5409 1515 5413
rect 1519 5409 1520 5413
rect 1514 5408 1520 5409
rect 1650 5413 1656 5414
rect 1650 5409 1651 5413
rect 1655 5409 1656 5413
rect 1650 5408 1656 5409
rect 1786 5413 1792 5414
rect 1786 5409 1787 5413
rect 1791 5409 1792 5413
rect 1786 5408 1792 5409
rect 1934 5412 1940 5413
rect 1934 5408 1935 5412
rect 1939 5408 1940 5412
rect 110 5407 116 5408
rect 1934 5407 1940 5408
rect 3838 5393 3844 5394
rect 5662 5393 5668 5394
rect 3838 5389 3839 5393
rect 3843 5389 3844 5393
rect 3838 5388 3844 5389
rect 4302 5392 4308 5393
rect 4302 5388 4303 5392
rect 4307 5388 4308 5392
rect 4302 5387 4308 5388
rect 4518 5392 4524 5393
rect 4518 5388 4519 5392
rect 4523 5388 4524 5392
rect 4518 5387 4524 5388
rect 4734 5392 4740 5393
rect 4734 5388 4735 5392
rect 4739 5388 4740 5392
rect 4734 5387 4740 5388
rect 4950 5392 4956 5393
rect 4950 5388 4951 5392
rect 4955 5388 4956 5392
rect 4950 5387 4956 5388
rect 5174 5392 5180 5393
rect 5174 5388 5175 5392
rect 5179 5388 5180 5392
rect 5174 5387 5180 5388
rect 5398 5392 5404 5393
rect 5398 5388 5399 5392
rect 5403 5388 5404 5392
rect 5662 5389 5663 5393
rect 5667 5389 5668 5393
rect 5662 5388 5668 5389
rect 5398 5387 5404 5388
rect 4274 5377 4280 5378
rect 3838 5376 3844 5377
rect 3838 5372 3839 5376
rect 3843 5372 3844 5376
rect 4274 5373 4275 5377
rect 4279 5373 4280 5377
rect 4274 5372 4280 5373
rect 4490 5377 4496 5378
rect 4490 5373 4491 5377
rect 4495 5373 4496 5377
rect 4490 5372 4496 5373
rect 4706 5377 4712 5378
rect 4706 5373 4707 5377
rect 4711 5373 4712 5377
rect 4706 5372 4712 5373
rect 4922 5377 4928 5378
rect 4922 5373 4923 5377
rect 4927 5373 4928 5377
rect 4922 5372 4928 5373
rect 5146 5377 5152 5378
rect 5146 5373 5147 5377
rect 5151 5373 5152 5377
rect 5146 5372 5152 5373
rect 5370 5377 5376 5378
rect 5370 5373 5371 5377
rect 5375 5373 5376 5377
rect 5370 5372 5376 5373
rect 5662 5376 5668 5377
rect 5662 5372 5663 5376
rect 5667 5372 5668 5376
rect 3838 5371 3844 5372
rect 5662 5371 5668 5372
rect 1974 5308 1980 5309
rect 3798 5308 3804 5309
rect 1974 5304 1975 5308
rect 1979 5304 1980 5308
rect 1974 5303 1980 5304
rect 2642 5307 2648 5308
rect 2642 5303 2643 5307
rect 2647 5303 2648 5307
rect 2642 5302 2648 5303
rect 2810 5307 2816 5308
rect 2810 5303 2811 5307
rect 2815 5303 2816 5307
rect 2810 5302 2816 5303
rect 2978 5307 2984 5308
rect 2978 5303 2979 5307
rect 2983 5303 2984 5307
rect 2978 5302 2984 5303
rect 3138 5307 3144 5308
rect 3138 5303 3139 5307
rect 3143 5303 3144 5307
rect 3138 5302 3144 5303
rect 3306 5307 3312 5308
rect 3306 5303 3307 5307
rect 3311 5303 3312 5307
rect 3306 5302 3312 5303
rect 3474 5307 3480 5308
rect 3474 5303 3475 5307
rect 3479 5303 3480 5307
rect 3474 5302 3480 5303
rect 3642 5307 3648 5308
rect 3642 5303 3643 5307
rect 3647 5303 3648 5307
rect 3798 5304 3799 5308
rect 3803 5304 3804 5308
rect 3798 5303 3804 5304
rect 3642 5302 3648 5303
rect 2670 5292 2676 5293
rect 1974 5291 1980 5292
rect 1974 5287 1975 5291
rect 1979 5287 1980 5291
rect 2670 5288 2671 5292
rect 2675 5288 2676 5292
rect 2670 5287 2676 5288
rect 2838 5292 2844 5293
rect 2838 5288 2839 5292
rect 2843 5288 2844 5292
rect 2838 5287 2844 5288
rect 3006 5292 3012 5293
rect 3006 5288 3007 5292
rect 3011 5288 3012 5292
rect 3006 5287 3012 5288
rect 3166 5292 3172 5293
rect 3166 5288 3167 5292
rect 3171 5288 3172 5292
rect 3166 5287 3172 5288
rect 3334 5292 3340 5293
rect 3334 5288 3335 5292
rect 3339 5288 3340 5292
rect 3334 5287 3340 5288
rect 3502 5292 3508 5293
rect 3502 5288 3503 5292
rect 3507 5288 3508 5292
rect 3502 5287 3508 5288
rect 3670 5292 3676 5293
rect 3670 5288 3671 5292
rect 3675 5288 3676 5292
rect 3670 5287 3676 5288
rect 3798 5291 3804 5292
rect 3798 5287 3799 5291
rect 3803 5287 3804 5291
rect 1974 5286 1980 5287
rect 3798 5286 3804 5287
rect 110 5256 116 5257
rect 1934 5256 1940 5257
rect 110 5252 111 5256
rect 115 5252 116 5256
rect 110 5251 116 5252
rect 410 5255 416 5256
rect 410 5251 411 5255
rect 415 5251 416 5255
rect 410 5250 416 5251
rect 586 5255 592 5256
rect 586 5251 587 5255
rect 591 5251 592 5255
rect 586 5250 592 5251
rect 762 5255 768 5256
rect 762 5251 763 5255
rect 767 5251 768 5255
rect 762 5250 768 5251
rect 938 5255 944 5256
rect 938 5251 939 5255
rect 943 5251 944 5255
rect 938 5250 944 5251
rect 1106 5255 1112 5256
rect 1106 5251 1107 5255
rect 1111 5251 1112 5255
rect 1106 5250 1112 5251
rect 1274 5255 1280 5256
rect 1274 5251 1275 5255
rect 1279 5251 1280 5255
rect 1274 5250 1280 5251
rect 1442 5255 1448 5256
rect 1442 5251 1443 5255
rect 1447 5251 1448 5255
rect 1442 5250 1448 5251
rect 1610 5255 1616 5256
rect 1610 5251 1611 5255
rect 1615 5251 1616 5255
rect 1610 5250 1616 5251
rect 1786 5255 1792 5256
rect 1786 5251 1787 5255
rect 1791 5251 1792 5255
rect 1934 5252 1935 5256
rect 1939 5252 1940 5256
rect 1934 5251 1940 5252
rect 1786 5250 1792 5251
rect 438 5240 444 5241
rect 110 5239 116 5240
rect 110 5235 111 5239
rect 115 5235 116 5239
rect 438 5236 439 5240
rect 443 5236 444 5240
rect 438 5235 444 5236
rect 614 5240 620 5241
rect 614 5236 615 5240
rect 619 5236 620 5240
rect 614 5235 620 5236
rect 790 5240 796 5241
rect 790 5236 791 5240
rect 795 5236 796 5240
rect 790 5235 796 5236
rect 966 5240 972 5241
rect 966 5236 967 5240
rect 971 5236 972 5240
rect 966 5235 972 5236
rect 1134 5240 1140 5241
rect 1134 5236 1135 5240
rect 1139 5236 1140 5240
rect 1134 5235 1140 5236
rect 1302 5240 1308 5241
rect 1302 5236 1303 5240
rect 1307 5236 1308 5240
rect 1302 5235 1308 5236
rect 1470 5240 1476 5241
rect 1470 5236 1471 5240
rect 1475 5236 1476 5240
rect 1470 5235 1476 5236
rect 1638 5240 1644 5241
rect 1638 5236 1639 5240
rect 1643 5236 1644 5240
rect 1638 5235 1644 5236
rect 1814 5240 1820 5241
rect 1814 5236 1815 5240
rect 1819 5236 1820 5240
rect 1814 5235 1820 5236
rect 1934 5239 1940 5240
rect 1934 5235 1935 5239
rect 1939 5235 1940 5239
rect 110 5234 116 5235
rect 1934 5234 1940 5235
rect 1974 5233 1980 5234
rect 3798 5233 3804 5234
rect 1974 5229 1975 5233
rect 1979 5229 1980 5233
rect 1974 5228 1980 5229
rect 2510 5232 2516 5233
rect 2510 5228 2511 5232
rect 2515 5228 2516 5232
rect 2510 5227 2516 5228
rect 2686 5232 2692 5233
rect 2686 5228 2687 5232
rect 2691 5228 2692 5232
rect 2686 5227 2692 5228
rect 2862 5232 2868 5233
rect 2862 5228 2863 5232
rect 2867 5228 2868 5232
rect 2862 5227 2868 5228
rect 3038 5232 3044 5233
rect 3038 5228 3039 5232
rect 3043 5228 3044 5232
rect 3038 5227 3044 5228
rect 3206 5232 3212 5233
rect 3206 5228 3207 5232
rect 3211 5228 3212 5232
rect 3206 5227 3212 5228
rect 3366 5232 3372 5233
rect 3366 5228 3367 5232
rect 3371 5228 3372 5232
rect 3366 5227 3372 5228
rect 3534 5232 3540 5233
rect 3534 5228 3535 5232
rect 3539 5228 3540 5232
rect 3534 5227 3540 5228
rect 3678 5232 3684 5233
rect 3678 5228 3679 5232
rect 3683 5228 3684 5232
rect 3798 5229 3799 5233
rect 3803 5229 3804 5233
rect 3798 5228 3804 5229
rect 3678 5227 3684 5228
rect 2482 5217 2488 5218
rect 1974 5216 1980 5217
rect 1974 5212 1975 5216
rect 1979 5212 1980 5216
rect 2482 5213 2483 5217
rect 2487 5213 2488 5217
rect 2482 5212 2488 5213
rect 2658 5217 2664 5218
rect 2658 5213 2659 5217
rect 2663 5213 2664 5217
rect 2658 5212 2664 5213
rect 2834 5217 2840 5218
rect 2834 5213 2835 5217
rect 2839 5213 2840 5217
rect 2834 5212 2840 5213
rect 3010 5217 3016 5218
rect 3010 5213 3011 5217
rect 3015 5213 3016 5217
rect 3010 5212 3016 5213
rect 3178 5217 3184 5218
rect 3178 5213 3179 5217
rect 3183 5213 3184 5217
rect 3178 5212 3184 5213
rect 3338 5217 3344 5218
rect 3338 5213 3339 5217
rect 3343 5213 3344 5217
rect 3338 5212 3344 5213
rect 3506 5217 3512 5218
rect 3506 5213 3507 5217
rect 3511 5213 3512 5217
rect 3506 5212 3512 5213
rect 3650 5217 3656 5218
rect 3650 5213 3651 5217
rect 3655 5213 3656 5217
rect 3650 5212 3656 5213
rect 3798 5216 3804 5217
rect 3798 5212 3799 5216
rect 3803 5212 3804 5216
rect 1974 5211 1980 5212
rect 3798 5211 3804 5212
rect 3838 5212 3844 5213
rect 5662 5212 5668 5213
rect 3838 5208 3839 5212
rect 3843 5208 3844 5212
rect 3838 5207 3844 5208
rect 4370 5211 4376 5212
rect 4370 5207 4371 5211
rect 4375 5207 4376 5211
rect 4370 5206 4376 5207
rect 4562 5211 4568 5212
rect 4562 5207 4563 5211
rect 4567 5207 4568 5211
rect 4562 5206 4568 5207
rect 4770 5211 4776 5212
rect 4770 5207 4771 5211
rect 4775 5207 4776 5211
rect 4770 5206 4776 5207
rect 4978 5211 4984 5212
rect 4978 5207 4979 5211
rect 4983 5207 4984 5211
rect 4978 5206 4984 5207
rect 5194 5211 5200 5212
rect 5194 5207 5195 5211
rect 5199 5207 5200 5211
rect 5194 5206 5200 5207
rect 5418 5211 5424 5212
rect 5418 5207 5419 5211
rect 5423 5207 5424 5211
rect 5662 5208 5663 5212
rect 5667 5208 5668 5212
rect 5662 5207 5668 5208
rect 5418 5206 5424 5207
rect 4398 5196 4404 5197
rect 3838 5195 3844 5196
rect 3838 5191 3839 5195
rect 3843 5191 3844 5195
rect 4398 5192 4399 5196
rect 4403 5192 4404 5196
rect 4398 5191 4404 5192
rect 4590 5196 4596 5197
rect 4590 5192 4591 5196
rect 4595 5192 4596 5196
rect 4590 5191 4596 5192
rect 4798 5196 4804 5197
rect 4798 5192 4799 5196
rect 4803 5192 4804 5196
rect 4798 5191 4804 5192
rect 5006 5196 5012 5197
rect 5006 5192 5007 5196
rect 5011 5192 5012 5196
rect 5006 5191 5012 5192
rect 5222 5196 5228 5197
rect 5222 5192 5223 5196
rect 5227 5192 5228 5196
rect 5222 5191 5228 5192
rect 5446 5196 5452 5197
rect 5446 5192 5447 5196
rect 5451 5192 5452 5196
rect 5446 5191 5452 5192
rect 5662 5195 5668 5196
rect 5662 5191 5663 5195
rect 5667 5191 5668 5195
rect 3838 5190 3844 5191
rect 5662 5190 5668 5191
rect 110 5173 116 5174
rect 1934 5173 1940 5174
rect 110 5169 111 5173
rect 115 5169 116 5173
rect 110 5168 116 5169
rect 206 5172 212 5173
rect 206 5168 207 5172
rect 211 5168 212 5172
rect 206 5167 212 5168
rect 342 5172 348 5173
rect 342 5168 343 5172
rect 347 5168 348 5172
rect 342 5167 348 5168
rect 478 5172 484 5173
rect 478 5168 479 5172
rect 483 5168 484 5172
rect 478 5167 484 5168
rect 614 5172 620 5173
rect 614 5168 615 5172
rect 619 5168 620 5172
rect 614 5167 620 5168
rect 750 5172 756 5173
rect 750 5168 751 5172
rect 755 5168 756 5172
rect 750 5167 756 5168
rect 886 5172 892 5173
rect 886 5168 887 5172
rect 891 5168 892 5172
rect 886 5167 892 5168
rect 1022 5172 1028 5173
rect 1022 5168 1023 5172
rect 1027 5168 1028 5172
rect 1934 5169 1935 5173
rect 1939 5169 1940 5173
rect 1934 5168 1940 5169
rect 1022 5167 1028 5168
rect 178 5157 184 5158
rect 110 5156 116 5157
rect 110 5152 111 5156
rect 115 5152 116 5156
rect 178 5153 179 5157
rect 183 5153 184 5157
rect 178 5152 184 5153
rect 314 5157 320 5158
rect 314 5153 315 5157
rect 319 5153 320 5157
rect 314 5152 320 5153
rect 450 5157 456 5158
rect 450 5153 451 5157
rect 455 5153 456 5157
rect 450 5152 456 5153
rect 586 5157 592 5158
rect 586 5153 587 5157
rect 591 5153 592 5157
rect 586 5152 592 5153
rect 722 5157 728 5158
rect 722 5153 723 5157
rect 727 5153 728 5157
rect 722 5152 728 5153
rect 858 5157 864 5158
rect 858 5153 859 5157
rect 863 5153 864 5157
rect 858 5152 864 5153
rect 994 5157 1000 5158
rect 994 5153 995 5157
rect 999 5153 1000 5157
rect 994 5152 1000 5153
rect 1934 5156 1940 5157
rect 1934 5152 1935 5156
rect 1939 5152 1940 5156
rect 110 5151 116 5152
rect 1934 5151 1940 5152
rect 3838 5113 3844 5114
rect 5662 5113 5668 5114
rect 3838 5109 3839 5113
rect 3843 5109 3844 5113
rect 3838 5108 3844 5109
rect 3886 5112 3892 5113
rect 3886 5108 3887 5112
rect 3891 5108 3892 5112
rect 3886 5107 3892 5108
rect 4086 5112 4092 5113
rect 4086 5108 4087 5112
rect 4091 5108 4092 5112
rect 4086 5107 4092 5108
rect 4310 5112 4316 5113
rect 4310 5108 4311 5112
rect 4315 5108 4316 5112
rect 4310 5107 4316 5108
rect 4534 5112 4540 5113
rect 4534 5108 4535 5112
rect 4539 5108 4540 5112
rect 4534 5107 4540 5108
rect 4758 5112 4764 5113
rect 4758 5108 4759 5112
rect 4763 5108 4764 5112
rect 4758 5107 4764 5108
rect 4982 5112 4988 5113
rect 4982 5108 4983 5112
rect 4987 5108 4988 5112
rect 4982 5107 4988 5108
rect 5206 5112 5212 5113
rect 5206 5108 5207 5112
rect 5211 5108 5212 5112
rect 5206 5107 5212 5108
rect 5438 5112 5444 5113
rect 5438 5108 5439 5112
rect 5443 5108 5444 5112
rect 5662 5109 5663 5113
rect 5667 5109 5668 5113
rect 5662 5108 5668 5109
rect 5438 5107 5444 5108
rect 3858 5097 3864 5098
rect 3838 5096 3844 5097
rect 3838 5092 3839 5096
rect 3843 5092 3844 5096
rect 3858 5093 3859 5097
rect 3863 5093 3864 5097
rect 3858 5092 3864 5093
rect 4058 5097 4064 5098
rect 4058 5093 4059 5097
rect 4063 5093 4064 5097
rect 4058 5092 4064 5093
rect 4282 5097 4288 5098
rect 4282 5093 4283 5097
rect 4287 5093 4288 5097
rect 4282 5092 4288 5093
rect 4506 5097 4512 5098
rect 4506 5093 4507 5097
rect 4511 5093 4512 5097
rect 4506 5092 4512 5093
rect 4730 5097 4736 5098
rect 4730 5093 4731 5097
rect 4735 5093 4736 5097
rect 4730 5092 4736 5093
rect 4954 5097 4960 5098
rect 4954 5093 4955 5097
rect 4959 5093 4960 5097
rect 4954 5092 4960 5093
rect 5178 5097 5184 5098
rect 5178 5093 5179 5097
rect 5183 5093 5184 5097
rect 5178 5092 5184 5093
rect 5410 5097 5416 5098
rect 5410 5093 5411 5097
rect 5415 5093 5416 5097
rect 5410 5092 5416 5093
rect 5662 5096 5668 5097
rect 5662 5092 5663 5096
rect 5667 5092 5668 5096
rect 3838 5091 3844 5092
rect 5662 5091 5668 5092
rect 1974 5076 1980 5077
rect 3798 5076 3804 5077
rect 1974 5072 1975 5076
rect 1979 5072 1980 5076
rect 1974 5071 1980 5072
rect 2138 5075 2144 5076
rect 2138 5071 2139 5075
rect 2143 5071 2144 5075
rect 2138 5070 2144 5071
rect 2306 5075 2312 5076
rect 2306 5071 2307 5075
rect 2311 5071 2312 5075
rect 2306 5070 2312 5071
rect 2490 5075 2496 5076
rect 2490 5071 2491 5075
rect 2495 5071 2496 5075
rect 2490 5070 2496 5071
rect 2690 5075 2696 5076
rect 2690 5071 2691 5075
rect 2695 5071 2696 5075
rect 2690 5070 2696 5071
rect 2914 5075 2920 5076
rect 2914 5071 2915 5075
rect 2919 5071 2920 5075
rect 2914 5070 2920 5071
rect 3162 5075 3168 5076
rect 3162 5071 3163 5075
rect 3167 5071 3168 5075
rect 3162 5070 3168 5071
rect 3418 5075 3424 5076
rect 3418 5071 3419 5075
rect 3423 5071 3424 5075
rect 3418 5070 3424 5071
rect 3650 5075 3656 5076
rect 3650 5071 3651 5075
rect 3655 5071 3656 5075
rect 3798 5072 3799 5076
rect 3803 5072 3804 5076
rect 3798 5071 3804 5072
rect 3650 5070 3656 5071
rect 2166 5060 2172 5061
rect 1974 5059 1980 5060
rect 1974 5055 1975 5059
rect 1979 5055 1980 5059
rect 2166 5056 2167 5060
rect 2171 5056 2172 5060
rect 2166 5055 2172 5056
rect 2334 5060 2340 5061
rect 2334 5056 2335 5060
rect 2339 5056 2340 5060
rect 2334 5055 2340 5056
rect 2518 5060 2524 5061
rect 2518 5056 2519 5060
rect 2523 5056 2524 5060
rect 2518 5055 2524 5056
rect 2718 5060 2724 5061
rect 2718 5056 2719 5060
rect 2723 5056 2724 5060
rect 2718 5055 2724 5056
rect 2942 5060 2948 5061
rect 2942 5056 2943 5060
rect 2947 5056 2948 5060
rect 2942 5055 2948 5056
rect 3190 5060 3196 5061
rect 3190 5056 3191 5060
rect 3195 5056 3196 5060
rect 3190 5055 3196 5056
rect 3446 5060 3452 5061
rect 3446 5056 3447 5060
rect 3451 5056 3452 5060
rect 3446 5055 3452 5056
rect 3678 5060 3684 5061
rect 3678 5056 3679 5060
rect 3683 5056 3684 5060
rect 3678 5055 3684 5056
rect 3798 5059 3804 5060
rect 3798 5055 3799 5059
rect 3803 5055 3804 5059
rect 1974 5054 1980 5055
rect 3798 5054 3804 5055
rect 110 5004 116 5005
rect 1934 5004 1940 5005
rect 110 5000 111 5004
rect 115 5000 116 5004
rect 110 4999 116 5000
rect 146 5003 152 5004
rect 146 4999 147 5003
rect 151 4999 152 5003
rect 146 4998 152 4999
rect 338 5003 344 5004
rect 338 4999 339 5003
rect 343 4999 344 5003
rect 338 4998 344 4999
rect 530 5003 536 5004
rect 530 4999 531 5003
rect 535 4999 536 5003
rect 530 4998 536 4999
rect 730 5003 736 5004
rect 730 4999 731 5003
rect 735 4999 736 5003
rect 730 4998 736 4999
rect 930 5003 936 5004
rect 930 4999 931 5003
rect 935 4999 936 5003
rect 930 4998 936 4999
rect 1130 5003 1136 5004
rect 1130 4999 1131 5003
rect 1135 4999 1136 5003
rect 1934 5000 1935 5004
rect 1939 5000 1940 5004
rect 1934 4999 1940 5000
rect 1130 4998 1136 4999
rect 174 4988 180 4989
rect 110 4987 116 4988
rect 110 4983 111 4987
rect 115 4983 116 4987
rect 174 4984 175 4988
rect 179 4984 180 4988
rect 174 4983 180 4984
rect 366 4988 372 4989
rect 366 4984 367 4988
rect 371 4984 372 4988
rect 366 4983 372 4984
rect 558 4988 564 4989
rect 558 4984 559 4988
rect 563 4984 564 4988
rect 558 4983 564 4984
rect 758 4988 764 4989
rect 758 4984 759 4988
rect 763 4984 764 4988
rect 758 4983 764 4984
rect 958 4988 964 4989
rect 958 4984 959 4988
rect 963 4984 964 4988
rect 958 4983 964 4984
rect 1158 4988 1164 4989
rect 1158 4984 1159 4988
rect 1163 4984 1164 4988
rect 1158 4983 1164 4984
rect 1934 4987 1940 4988
rect 1934 4983 1935 4987
rect 1939 4983 1940 4987
rect 110 4982 116 4983
rect 1934 4982 1940 4983
rect 1974 4977 1980 4978
rect 3798 4977 3804 4978
rect 1974 4973 1975 4977
rect 1979 4973 1980 4977
rect 1974 4972 1980 4973
rect 2022 4976 2028 4977
rect 2022 4972 2023 4976
rect 2027 4972 2028 4976
rect 2022 4971 2028 4972
rect 2166 4976 2172 4977
rect 2166 4972 2167 4976
rect 2171 4972 2172 4976
rect 2166 4971 2172 4972
rect 2350 4976 2356 4977
rect 2350 4972 2351 4976
rect 2355 4972 2356 4976
rect 2350 4971 2356 4972
rect 2542 4976 2548 4977
rect 2542 4972 2543 4976
rect 2547 4972 2548 4976
rect 2542 4971 2548 4972
rect 2750 4976 2756 4977
rect 2750 4972 2751 4976
rect 2755 4972 2756 4976
rect 2750 4971 2756 4972
rect 2966 4976 2972 4977
rect 2966 4972 2967 4976
rect 2971 4972 2972 4976
rect 2966 4971 2972 4972
rect 3182 4976 3188 4977
rect 3182 4972 3183 4976
rect 3187 4972 3188 4976
rect 3798 4973 3799 4977
rect 3803 4973 3804 4977
rect 3798 4972 3804 4973
rect 3182 4971 3188 4972
rect 1994 4961 2000 4962
rect 1974 4960 1980 4961
rect 1974 4956 1975 4960
rect 1979 4956 1980 4960
rect 1994 4957 1995 4961
rect 1999 4957 2000 4961
rect 1994 4956 2000 4957
rect 2138 4961 2144 4962
rect 2138 4957 2139 4961
rect 2143 4957 2144 4961
rect 2138 4956 2144 4957
rect 2322 4961 2328 4962
rect 2322 4957 2323 4961
rect 2327 4957 2328 4961
rect 2322 4956 2328 4957
rect 2514 4961 2520 4962
rect 2514 4957 2515 4961
rect 2519 4957 2520 4961
rect 2514 4956 2520 4957
rect 2722 4961 2728 4962
rect 2722 4957 2723 4961
rect 2727 4957 2728 4961
rect 2722 4956 2728 4957
rect 2938 4961 2944 4962
rect 2938 4957 2939 4961
rect 2943 4957 2944 4961
rect 2938 4956 2944 4957
rect 3154 4961 3160 4962
rect 3154 4957 3155 4961
rect 3159 4957 3160 4961
rect 3154 4956 3160 4957
rect 3798 4960 3804 4961
rect 3798 4956 3799 4960
rect 3803 4956 3804 4960
rect 1974 4955 1980 4956
rect 3798 4955 3804 4956
rect 3838 4948 3844 4949
rect 5662 4948 5668 4949
rect 3838 4944 3839 4948
rect 3843 4944 3844 4948
rect 3838 4943 3844 4944
rect 3858 4947 3864 4948
rect 3858 4943 3859 4947
rect 3863 4943 3864 4947
rect 3858 4942 3864 4943
rect 3994 4947 4000 4948
rect 3994 4943 3995 4947
rect 3999 4943 4000 4947
rect 3994 4942 4000 4943
rect 4130 4947 4136 4948
rect 4130 4943 4131 4947
rect 4135 4943 4136 4947
rect 4130 4942 4136 4943
rect 4282 4947 4288 4948
rect 4282 4943 4283 4947
rect 4287 4943 4288 4947
rect 4282 4942 4288 4943
rect 4442 4947 4448 4948
rect 4442 4943 4443 4947
rect 4447 4943 4448 4947
rect 4442 4942 4448 4943
rect 4610 4947 4616 4948
rect 4610 4943 4611 4947
rect 4615 4943 4616 4947
rect 4610 4942 4616 4943
rect 4786 4947 4792 4948
rect 4786 4943 4787 4947
rect 4791 4943 4792 4947
rect 4786 4942 4792 4943
rect 4970 4947 4976 4948
rect 4970 4943 4971 4947
rect 4975 4943 4976 4947
rect 4970 4942 4976 4943
rect 5154 4947 5160 4948
rect 5154 4943 5155 4947
rect 5159 4943 5160 4947
rect 5154 4942 5160 4943
rect 5338 4947 5344 4948
rect 5338 4943 5339 4947
rect 5343 4943 5344 4947
rect 5338 4942 5344 4943
rect 5514 4947 5520 4948
rect 5514 4943 5515 4947
rect 5519 4943 5520 4947
rect 5662 4944 5663 4948
rect 5667 4944 5668 4948
rect 5662 4943 5668 4944
rect 5514 4942 5520 4943
rect 3886 4932 3892 4933
rect 3838 4931 3844 4932
rect 3838 4927 3839 4931
rect 3843 4927 3844 4931
rect 3886 4928 3887 4932
rect 3891 4928 3892 4932
rect 3886 4927 3892 4928
rect 4022 4932 4028 4933
rect 4022 4928 4023 4932
rect 4027 4928 4028 4932
rect 4022 4927 4028 4928
rect 4158 4932 4164 4933
rect 4158 4928 4159 4932
rect 4163 4928 4164 4932
rect 4158 4927 4164 4928
rect 4310 4932 4316 4933
rect 4310 4928 4311 4932
rect 4315 4928 4316 4932
rect 4310 4927 4316 4928
rect 4470 4932 4476 4933
rect 4470 4928 4471 4932
rect 4475 4928 4476 4932
rect 4470 4927 4476 4928
rect 4638 4932 4644 4933
rect 4638 4928 4639 4932
rect 4643 4928 4644 4932
rect 4638 4927 4644 4928
rect 4814 4932 4820 4933
rect 4814 4928 4815 4932
rect 4819 4928 4820 4932
rect 4814 4927 4820 4928
rect 4998 4932 5004 4933
rect 4998 4928 4999 4932
rect 5003 4928 5004 4932
rect 4998 4927 5004 4928
rect 5182 4932 5188 4933
rect 5182 4928 5183 4932
rect 5187 4928 5188 4932
rect 5182 4927 5188 4928
rect 5366 4932 5372 4933
rect 5366 4928 5367 4932
rect 5371 4928 5372 4932
rect 5366 4927 5372 4928
rect 5542 4932 5548 4933
rect 5542 4928 5543 4932
rect 5547 4928 5548 4932
rect 5542 4927 5548 4928
rect 5662 4931 5668 4932
rect 5662 4927 5663 4931
rect 5667 4927 5668 4931
rect 3838 4926 3844 4927
rect 5662 4926 5668 4927
rect 110 4917 116 4918
rect 1934 4917 1940 4918
rect 110 4913 111 4917
rect 115 4913 116 4917
rect 110 4912 116 4913
rect 158 4916 164 4917
rect 158 4912 159 4916
rect 163 4912 164 4916
rect 158 4911 164 4912
rect 390 4916 396 4917
rect 390 4912 391 4916
rect 395 4912 396 4916
rect 390 4911 396 4912
rect 646 4916 652 4917
rect 646 4912 647 4916
rect 651 4912 652 4916
rect 646 4911 652 4912
rect 894 4916 900 4917
rect 894 4912 895 4916
rect 899 4912 900 4916
rect 894 4911 900 4912
rect 1134 4916 1140 4917
rect 1134 4912 1135 4916
rect 1139 4912 1140 4916
rect 1134 4911 1140 4912
rect 1366 4916 1372 4917
rect 1366 4912 1367 4916
rect 1371 4912 1372 4916
rect 1366 4911 1372 4912
rect 1598 4916 1604 4917
rect 1598 4912 1599 4916
rect 1603 4912 1604 4916
rect 1598 4911 1604 4912
rect 1814 4916 1820 4917
rect 1814 4912 1815 4916
rect 1819 4912 1820 4916
rect 1934 4913 1935 4917
rect 1939 4913 1940 4917
rect 1934 4912 1940 4913
rect 1814 4911 1820 4912
rect 130 4901 136 4902
rect 110 4900 116 4901
rect 110 4896 111 4900
rect 115 4896 116 4900
rect 130 4897 131 4901
rect 135 4897 136 4901
rect 130 4896 136 4897
rect 362 4901 368 4902
rect 362 4897 363 4901
rect 367 4897 368 4901
rect 362 4896 368 4897
rect 618 4901 624 4902
rect 618 4897 619 4901
rect 623 4897 624 4901
rect 618 4896 624 4897
rect 866 4901 872 4902
rect 866 4897 867 4901
rect 871 4897 872 4901
rect 866 4896 872 4897
rect 1106 4901 1112 4902
rect 1106 4897 1107 4901
rect 1111 4897 1112 4901
rect 1106 4896 1112 4897
rect 1338 4901 1344 4902
rect 1338 4897 1339 4901
rect 1343 4897 1344 4901
rect 1338 4896 1344 4897
rect 1570 4901 1576 4902
rect 1570 4897 1571 4901
rect 1575 4897 1576 4901
rect 1570 4896 1576 4897
rect 1786 4901 1792 4902
rect 1786 4897 1787 4901
rect 1791 4897 1792 4901
rect 1786 4896 1792 4897
rect 1934 4900 1940 4901
rect 1934 4896 1935 4900
rect 1939 4896 1940 4900
rect 110 4895 116 4896
rect 1934 4895 1940 4896
rect 3838 4857 3844 4858
rect 5662 4857 5668 4858
rect 3838 4853 3839 4857
rect 3843 4853 3844 4857
rect 3838 4852 3844 4853
rect 3942 4856 3948 4857
rect 3942 4852 3943 4856
rect 3947 4852 3948 4856
rect 3942 4851 3948 4852
rect 4182 4856 4188 4857
rect 4182 4852 4183 4856
rect 4187 4852 4188 4856
rect 4182 4851 4188 4852
rect 4430 4856 4436 4857
rect 4430 4852 4431 4856
rect 4435 4852 4436 4856
rect 4430 4851 4436 4852
rect 4686 4856 4692 4857
rect 4686 4852 4687 4856
rect 4691 4852 4692 4856
rect 4686 4851 4692 4852
rect 4958 4856 4964 4857
rect 4958 4852 4959 4856
rect 4963 4852 4964 4856
rect 4958 4851 4964 4852
rect 5238 4856 5244 4857
rect 5238 4852 5239 4856
rect 5243 4852 5244 4856
rect 5238 4851 5244 4852
rect 5518 4856 5524 4857
rect 5518 4852 5519 4856
rect 5523 4852 5524 4856
rect 5662 4853 5663 4857
rect 5667 4853 5668 4857
rect 5662 4852 5668 4853
rect 5518 4851 5524 4852
rect 3914 4841 3920 4842
rect 3838 4840 3844 4841
rect 3838 4836 3839 4840
rect 3843 4836 3844 4840
rect 3914 4837 3915 4841
rect 3919 4837 3920 4841
rect 3914 4836 3920 4837
rect 4154 4841 4160 4842
rect 4154 4837 4155 4841
rect 4159 4837 4160 4841
rect 4154 4836 4160 4837
rect 4402 4841 4408 4842
rect 4402 4837 4403 4841
rect 4407 4837 4408 4841
rect 4402 4836 4408 4837
rect 4658 4841 4664 4842
rect 4658 4837 4659 4841
rect 4663 4837 4664 4841
rect 4658 4836 4664 4837
rect 4930 4841 4936 4842
rect 4930 4837 4931 4841
rect 4935 4837 4936 4841
rect 4930 4836 4936 4837
rect 5210 4841 5216 4842
rect 5210 4837 5211 4841
rect 5215 4837 5216 4841
rect 5210 4836 5216 4837
rect 5490 4841 5496 4842
rect 5490 4837 5491 4841
rect 5495 4837 5496 4841
rect 5490 4836 5496 4837
rect 5662 4840 5668 4841
rect 5662 4836 5663 4840
rect 5667 4836 5668 4840
rect 3838 4835 3844 4836
rect 5662 4835 5668 4836
rect 1974 4820 1980 4821
rect 3798 4820 3804 4821
rect 1974 4816 1975 4820
rect 1979 4816 1980 4820
rect 1974 4815 1980 4816
rect 1994 4819 2000 4820
rect 1994 4815 1995 4819
rect 1999 4815 2000 4819
rect 1994 4814 2000 4815
rect 2322 4819 2328 4820
rect 2322 4815 2323 4819
rect 2327 4815 2328 4819
rect 2322 4814 2328 4815
rect 2666 4819 2672 4820
rect 2666 4815 2667 4819
rect 2671 4815 2672 4819
rect 2666 4814 2672 4815
rect 3018 4819 3024 4820
rect 3018 4815 3019 4819
rect 3023 4815 3024 4819
rect 3018 4814 3024 4815
rect 3370 4819 3376 4820
rect 3370 4815 3371 4819
rect 3375 4815 3376 4819
rect 3798 4816 3799 4820
rect 3803 4816 3804 4820
rect 3798 4815 3804 4816
rect 3370 4814 3376 4815
rect 2022 4804 2028 4805
rect 1974 4803 1980 4804
rect 1974 4799 1975 4803
rect 1979 4799 1980 4803
rect 2022 4800 2023 4804
rect 2027 4800 2028 4804
rect 2022 4799 2028 4800
rect 2350 4804 2356 4805
rect 2350 4800 2351 4804
rect 2355 4800 2356 4804
rect 2350 4799 2356 4800
rect 2694 4804 2700 4805
rect 2694 4800 2695 4804
rect 2699 4800 2700 4804
rect 2694 4799 2700 4800
rect 3046 4804 3052 4805
rect 3046 4800 3047 4804
rect 3051 4800 3052 4804
rect 3046 4799 3052 4800
rect 3398 4804 3404 4805
rect 3398 4800 3399 4804
rect 3403 4800 3404 4804
rect 3398 4799 3404 4800
rect 3798 4803 3804 4804
rect 3798 4799 3799 4803
rect 3803 4799 3804 4803
rect 1974 4798 1980 4799
rect 3798 4798 3804 4799
rect 110 4768 116 4769
rect 1934 4768 1940 4769
rect 110 4764 111 4768
rect 115 4764 116 4768
rect 110 4763 116 4764
rect 130 4767 136 4768
rect 130 4763 131 4767
rect 135 4763 136 4767
rect 130 4762 136 4763
rect 474 4767 480 4768
rect 474 4763 475 4767
rect 479 4763 480 4767
rect 474 4762 480 4763
rect 858 4767 864 4768
rect 858 4763 859 4767
rect 863 4763 864 4767
rect 858 4762 864 4763
rect 1250 4767 1256 4768
rect 1250 4763 1251 4767
rect 1255 4763 1256 4767
rect 1250 4762 1256 4763
rect 1642 4767 1648 4768
rect 1642 4763 1643 4767
rect 1647 4763 1648 4767
rect 1934 4764 1935 4768
rect 1939 4764 1940 4768
rect 1934 4763 1940 4764
rect 1642 4762 1648 4763
rect 158 4752 164 4753
rect 110 4751 116 4752
rect 110 4747 111 4751
rect 115 4747 116 4751
rect 158 4748 159 4752
rect 163 4748 164 4752
rect 158 4747 164 4748
rect 502 4752 508 4753
rect 502 4748 503 4752
rect 507 4748 508 4752
rect 502 4747 508 4748
rect 886 4752 892 4753
rect 886 4748 887 4752
rect 891 4748 892 4752
rect 886 4747 892 4748
rect 1278 4752 1284 4753
rect 1278 4748 1279 4752
rect 1283 4748 1284 4752
rect 1278 4747 1284 4748
rect 1670 4752 1676 4753
rect 1670 4748 1671 4752
rect 1675 4748 1676 4752
rect 1670 4747 1676 4748
rect 1934 4751 1940 4752
rect 1934 4747 1935 4751
rect 1939 4747 1940 4751
rect 110 4746 116 4747
rect 1934 4746 1940 4747
rect 3838 4700 3844 4701
rect 5662 4700 5668 4701
rect 1974 4697 1980 4698
rect 3798 4697 3804 4698
rect 1974 4693 1975 4697
rect 1979 4693 1980 4697
rect 1974 4692 1980 4693
rect 2078 4696 2084 4697
rect 2078 4692 2079 4696
rect 2083 4692 2084 4696
rect 2078 4691 2084 4692
rect 2230 4696 2236 4697
rect 2230 4692 2231 4696
rect 2235 4692 2236 4696
rect 2230 4691 2236 4692
rect 2390 4696 2396 4697
rect 2390 4692 2391 4696
rect 2395 4692 2396 4696
rect 2390 4691 2396 4692
rect 2558 4696 2564 4697
rect 2558 4692 2559 4696
rect 2563 4692 2564 4696
rect 2558 4691 2564 4692
rect 2726 4696 2732 4697
rect 2726 4692 2727 4696
rect 2731 4692 2732 4696
rect 2726 4691 2732 4692
rect 2902 4696 2908 4697
rect 2902 4692 2903 4696
rect 2907 4692 2908 4696
rect 2902 4691 2908 4692
rect 3078 4696 3084 4697
rect 3078 4692 3079 4696
rect 3083 4692 3084 4696
rect 3078 4691 3084 4692
rect 3254 4696 3260 4697
rect 3254 4692 3255 4696
rect 3259 4692 3260 4696
rect 3254 4691 3260 4692
rect 3438 4696 3444 4697
rect 3438 4692 3439 4696
rect 3443 4692 3444 4696
rect 3438 4691 3444 4692
rect 3622 4696 3628 4697
rect 3622 4692 3623 4696
rect 3627 4692 3628 4696
rect 3798 4693 3799 4697
rect 3803 4693 3804 4697
rect 3838 4696 3839 4700
rect 3843 4696 3844 4700
rect 3838 4695 3844 4696
rect 3938 4699 3944 4700
rect 3938 4695 3939 4699
rect 3943 4695 3944 4699
rect 3938 4694 3944 4695
rect 4178 4699 4184 4700
rect 4178 4695 4179 4699
rect 4183 4695 4184 4699
rect 4178 4694 4184 4695
rect 4434 4699 4440 4700
rect 4434 4695 4435 4699
rect 4439 4695 4440 4699
rect 4434 4694 4440 4695
rect 4690 4699 4696 4700
rect 4690 4695 4691 4699
rect 4695 4695 4696 4699
rect 4690 4694 4696 4695
rect 4954 4699 4960 4700
rect 4954 4695 4955 4699
rect 4959 4695 4960 4699
rect 4954 4694 4960 4695
rect 5226 4699 5232 4700
rect 5226 4695 5227 4699
rect 5231 4695 5232 4699
rect 5226 4694 5232 4695
rect 5506 4699 5512 4700
rect 5506 4695 5507 4699
rect 5511 4695 5512 4699
rect 5662 4696 5663 4700
rect 5667 4696 5668 4700
rect 5662 4695 5668 4696
rect 5506 4694 5512 4695
rect 3798 4692 3804 4693
rect 3622 4691 3628 4692
rect 3966 4684 3972 4685
rect 3838 4683 3844 4684
rect 2050 4681 2056 4682
rect 1974 4680 1980 4681
rect 1974 4676 1975 4680
rect 1979 4676 1980 4680
rect 2050 4677 2051 4681
rect 2055 4677 2056 4681
rect 2050 4676 2056 4677
rect 2202 4681 2208 4682
rect 2202 4677 2203 4681
rect 2207 4677 2208 4681
rect 2202 4676 2208 4677
rect 2362 4681 2368 4682
rect 2362 4677 2363 4681
rect 2367 4677 2368 4681
rect 2362 4676 2368 4677
rect 2530 4681 2536 4682
rect 2530 4677 2531 4681
rect 2535 4677 2536 4681
rect 2530 4676 2536 4677
rect 2698 4681 2704 4682
rect 2698 4677 2699 4681
rect 2703 4677 2704 4681
rect 2698 4676 2704 4677
rect 2874 4681 2880 4682
rect 2874 4677 2875 4681
rect 2879 4677 2880 4681
rect 2874 4676 2880 4677
rect 3050 4681 3056 4682
rect 3050 4677 3051 4681
rect 3055 4677 3056 4681
rect 3050 4676 3056 4677
rect 3226 4681 3232 4682
rect 3226 4677 3227 4681
rect 3231 4677 3232 4681
rect 3226 4676 3232 4677
rect 3410 4681 3416 4682
rect 3410 4677 3411 4681
rect 3415 4677 3416 4681
rect 3410 4676 3416 4677
rect 3594 4681 3600 4682
rect 3594 4677 3595 4681
rect 3599 4677 3600 4681
rect 3594 4676 3600 4677
rect 3798 4680 3804 4681
rect 3798 4676 3799 4680
rect 3803 4676 3804 4680
rect 3838 4679 3839 4683
rect 3843 4679 3844 4683
rect 3966 4680 3967 4684
rect 3971 4680 3972 4684
rect 3966 4679 3972 4680
rect 4206 4684 4212 4685
rect 4206 4680 4207 4684
rect 4211 4680 4212 4684
rect 4206 4679 4212 4680
rect 4462 4684 4468 4685
rect 4462 4680 4463 4684
rect 4467 4680 4468 4684
rect 4462 4679 4468 4680
rect 4718 4684 4724 4685
rect 4718 4680 4719 4684
rect 4723 4680 4724 4684
rect 4718 4679 4724 4680
rect 4982 4684 4988 4685
rect 4982 4680 4983 4684
rect 4987 4680 4988 4684
rect 4982 4679 4988 4680
rect 5254 4684 5260 4685
rect 5254 4680 5255 4684
rect 5259 4680 5260 4684
rect 5254 4679 5260 4680
rect 5534 4684 5540 4685
rect 5534 4680 5535 4684
rect 5539 4680 5540 4684
rect 5534 4679 5540 4680
rect 5662 4683 5668 4684
rect 5662 4679 5663 4683
rect 5667 4679 5668 4683
rect 3838 4678 3844 4679
rect 5662 4678 5668 4679
rect 1974 4675 1980 4676
rect 3798 4675 3804 4676
rect 110 4673 116 4674
rect 1934 4673 1940 4674
rect 110 4669 111 4673
rect 115 4669 116 4673
rect 110 4668 116 4669
rect 158 4672 164 4673
rect 158 4668 159 4672
rect 163 4668 164 4672
rect 158 4667 164 4668
rect 294 4672 300 4673
rect 294 4668 295 4672
rect 299 4668 300 4672
rect 294 4667 300 4668
rect 430 4672 436 4673
rect 430 4668 431 4672
rect 435 4668 436 4672
rect 430 4667 436 4668
rect 566 4672 572 4673
rect 566 4668 567 4672
rect 571 4668 572 4672
rect 566 4667 572 4668
rect 702 4672 708 4673
rect 702 4668 703 4672
rect 707 4668 708 4672
rect 1934 4669 1935 4673
rect 1939 4669 1940 4673
rect 1934 4668 1940 4669
rect 702 4667 708 4668
rect 130 4657 136 4658
rect 110 4656 116 4657
rect 110 4652 111 4656
rect 115 4652 116 4656
rect 130 4653 131 4657
rect 135 4653 136 4657
rect 130 4652 136 4653
rect 266 4657 272 4658
rect 266 4653 267 4657
rect 271 4653 272 4657
rect 266 4652 272 4653
rect 402 4657 408 4658
rect 402 4653 403 4657
rect 407 4653 408 4657
rect 402 4652 408 4653
rect 538 4657 544 4658
rect 538 4653 539 4657
rect 543 4653 544 4657
rect 538 4652 544 4653
rect 674 4657 680 4658
rect 674 4653 675 4657
rect 679 4653 680 4657
rect 674 4652 680 4653
rect 1934 4656 1940 4657
rect 1934 4652 1935 4656
rect 1939 4652 1940 4656
rect 110 4651 116 4652
rect 1934 4651 1940 4652
rect 3838 4621 3844 4622
rect 5662 4621 5668 4622
rect 3838 4617 3839 4621
rect 3843 4617 3844 4621
rect 3838 4616 3844 4617
rect 4174 4620 4180 4621
rect 4174 4616 4175 4620
rect 4179 4616 4180 4620
rect 4174 4615 4180 4616
rect 4454 4620 4460 4621
rect 4454 4616 4455 4620
rect 4459 4616 4460 4620
rect 4454 4615 4460 4616
rect 4734 4620 4740 4621
rect 4734 4616 4735 4620
rect 4739 4616 4740 4620
rect 4734 4615 4740 4616
rect 5014 4620 5020 4621
rect 5014 4616 5015 4620
rect 5019 4616 5020 4620
rect 5014 4615 5020 4616
rect 5302 4620 5308 4621
rect 5302 4616 5303 4620
rect 5307 4616 5308 4620
rect 5662 4617 5663 4621
rect 5667 4617 5668 4621
rect 5662 4616 5668 4617
rect 5302 4615 5308 4616
rect 4146 4605 4152 4606
rect 3838 4604 3844 4605
rect 3838 4600 3839 4604
rect 3843 4600 3844 4604
rect 4146 4601 4147 4605
rect 4151 4601 4152 4605
rect 4146 4600 4152 4601
rect 4426 4605 4432 4606
rect 4426 4601 4427 4605
rect 4431 4601 4432 4605
rect 4426 4600 4432 4601
rect 4706 4605 4712 4606
rect 4706 4601 4707 4605
rect 4711 4601 4712 4605
rect 4706 4600 4712 4601
rect 4986 4605 4992 4606
rect 4986 4601 4987 4605
rect 4991 4601 4992 4605
rect 4986 4600 4992 4601
rect 5274 4605 5280 4606
rect 5274 4601 5275 4605
rect 5279 4601 5280 4605
rect 5274 4600 5280 4601
rect 5662 4604 5668 4605
rect 5662 4600 5663 4604
rect 5667 4600 5668 4604
rect 3838 4599 3844 4600
rect 5662 4599 5668 4600
rect 1974 4544 1980 4545
rect 3798 4544 3804 4545
rect 1974 4540 1975 4544
rect 1979 4540 1980 4544
rect 1974 4539 1980 4540
rect 2122 4543 2128 4544
rect 2122 4539 2123 4543
rect 2127 4539 2128 4543
rect 2122 4538 2128 4539
rect 2274 4543 2280 4544
rect 2274 4539 2275 4543
rect 2279 4539 2280 4543
rect 2274 4538 2280 4539
rect 2442 4543 2448 4544
rect 2442 4539 2443 4543
rect 2447 4539 2448 4543
rect 2442 4538 2448 4539
rect 2610 4543 2616 4544
rect 2610 4539 2611 4543
rect 2615 4539 2616 4543
rect 2610 4538 2616 4539
rect 2786 4543 2792 4544
rect 2786 4539 2787 4543
rect 2791 4539 2792 4543
rect 2786 4538 2792 4539
rect 2962 4543 2968 4544
rect 2962 4539 2963 4543
rect 2967 4539 2968 4543
rect 2962 4538 2968 4539
rect 3138 4543 3144 4544
rect 3138 4539 3139 4543
rect 3143 4539 3144 4543
rect 3138 4538 3144 4539
rect 3314 4543 3320 4544
rect 3314 4539 3315 4543
rect 3319 4539 3320 4543
rect 3314 4538 3320 4539
rect 3490 4543 3496 4544
rect 3490 4539 3491 4543
rect 3495 4539 3496 4543
rect 3490 4538 3496 4539
rect 3650 4543 3656 4544
rect 3650 4539 3651 4543
rect 3655 4539 3656 4543
rect 3798 4540 3799 4544
rect 3803 4540 3804 4544
rect 3798 4539 3804 4540
rect 3650 4538 3656 4539
rect 2150 4528 2156 4529
rect 1974 4527 1980 4528
rect 1974 4523 1975 4527
rect 1979 4523 1980 4527
rect 2150 4524 2151 4528
rect 2155 4524 2156 4528
rect 2150 4523 2156 4524
rect 2302 4528 2308 4529
rect 2302 4524 2303 4528
rect 2307 4524 2308 4528
rect 2302 4523 2308 4524
rect 2470 4528 2476 4529
rect 2470 4524 2471 4528
rect 2475 4524 2476 4528
rect 2470 4523 2476 4524
rect 2638 4528 2644 4529
rect 2638 4524 2639 4528
rect 2643 4524 2644 4528
rect 2638 4523 2644 4524
rect 2814 4528 2820 4529
rect 2814 4524 2815 4528
rect 2819 4524 2820 4528
rect 2814 4523 2820 4524
rect 2990 4528 2996 4529
rect 2990 4524 2991 4528
rect 2995 4524 2996 4528
rect 2990 4523 2996 4524
rect 3166 4528 3172 4529
rect 3166 4524 3167 4528
rect 3171 4524 3172 4528
rect 3166 4523 3172 4524
rect 3342 4528 3348 4529
rect 3342 4524 3343 4528
rect 3347 4524 3348 4528
rect 3342 4523 3348 4524
rect 3518 4528 3524 4529
rect 3518 4524 3519 4528
rect 3523 4524 3524 4528
rect 3518 4523 3524 4524
rect 3678 4528 3684 4529
rect 3678 4524 3679 4528
rect 3683 4524 3684 4528
rect 3678 4523 3684 4524
rect 3798 4527 3804 4528
rect 3798 4523 3799 4527
rect 3803 4523 3804 4527
rect 1974 4522 1980 4523
rect 3798 4522 3804 4523
rect 110 4508 116 4509
rect 1934 4508 1940 4509
rect 110 4504 111 4508
rect 115 4504 116 4508
rect 110 4503 116 4504
rect 290 4507 296 4508
rect 290 4503 291 4507
rect 295 4503 296 4507
rect 290 4502 296 4503
rect 426 4507 432 4508
rect 426 4503 427 4507
rect 431 4503 432 4507
rect 426 4502 432 4503
rect 562 4507 568 4508
rect 562 4503 563 4507
rect 567 4503 568 4507
rect 562 4502 568 4503
rect 698 4507 704 4508
rect 698 4503 699 4507
rect 703 4503 704 4507
rect 698 4502 704 4503
rect 834 4507 840 4508
rect 834 4503 835 4507
rect 839 4503 840 4507
rect 1934 4504 1935 4508
rect 1939 4504 1940 4508
rect 1934 4503 1940 4504
rect 834 4502 840 4503
rect 318 4492 324 4493
rect 110 4491 116 4492
rect 110 4487 111 4491
rect 115 4487 116 4491
rect 318 4488 319 4492
rect 323 4488 324 4492
rect 318 4487 324 4488
rect 454 4492 460 4493
rect 454 4488 455 4492
rect 459 4488 460 4492
rect 454 4487 460 4488
rect 590 4492 596 4493
rect 590 4488 591 4492
rect 595 4488 596 4492
rect 590 4487 596 4488
rect 726 4492 732 4493
rect 726 4488 727 4492
rect 731 4488 732 4492
rect 726 4487 732 4488
rect 862 4492 868 4493
rect 862 4488 863 4492
rect 867 4488 868 4492
rect 862 4487 868 4488
rect 1934 4491 1940 4492
rect 1934 4487 1935 4491
rect 1939 4487 1940 4491
rect 110 4486 116 4487
rect 1934 4486 1940 4487
rect 3838 4468 3844 4469
rect 5662 4468 5668 4469
rect 3838 4464 3839 4468
rect 3843 4464 3844 4468
rect 3838 4463 3844 4464
rect 3858 4467 3864 4468
rect 3858 4463 3859 4467
rect 3863 4463 3864 4467
rect 3858 4462 3864 4463
rect 4154 4467 4160 4468
rect 4154 4463 4155 4467
rect 4159 4463 4160 4467
rect 4154 4462 4160 4463
rect 4482 4467 4488 4468
rect 4482 4463 4483 4467
rect 4487 4463 4488 4467
rect 4482 4462 4488 4463
rect 4818 4467 4824 4468
rect 4818 4463 4819 4467
rect 4823 4463 4824 4467
rect 4818 4462 4824 4463
rect 5162 4467 5168 4468
rect 5162 4463 5163 4467
rect 5167 4463 5168 4467
rect 5162 4462 5168 4463
rect 5514 4467 5520 4468
rect 5514 4463 5515 4467
rect 5519 4463 5520 4467
rect 5662 4464 5663 4468
rect 5667 4464 5668 4468
rect 5662 4463 5668 4464
rect 5514 4462 5520 4463
rect 1974 4461 1980 4462
rect 3798 4461 3804 4462
rect 1974 4457 1975 4461
rect 1979 4457 1980 4461
rect 1974 4456 1980 4457
rect 2022 4460 2028 4461
rect 2022 4456 2023 4460
rect 2027 4456 2028 4460
rect 2022 4455 2028 4456
rect 2158 4460 2164 4461
rect 2158 4456 2159 4460
rect 2163 4456 2164 4460
rect 2158 4455 2164 4456
rect 2294 4460 2300 4461
rect 2294 4456 2295 4460
rect 2299 4456 2300 4460
rect 2294 4455 2300 4456
rect 2430 4460 2436 4461
rect 2430 4456 2431 4460
rect 2435 4456 2436 4460
rect 2430 4455 2436 4456
rect 2566 4460 2572 4461
rect 2566 4456 2567 4460
rect 2571 4456 2572 4460
rect 2566 4455 2572 4456
rect 2702 4460 2708 4461
rect 2702 4456 2703 4460
rect 2707 4456 2708 4460
rect 2702 4455 2708 4456
rect 2838 4460 2844 4461
rect 2838 4456 2839 4460
rect 2843 4456 2844 4460
rect 2838 4455 2844 4456
rect 2974 4460 2980 4461
rect 2974 4456 2975 4460
rect 2979 4456 2980 4460
rect 3798 4457 3799 4461
rect 3803 4457 3804 4461
rect 3798 4456 3804 4457
rect 2974 4455 2980 4456
rect 3886 4452 3892 4453
rect 3838 4451 3844 4452
rect 3838 4447 3839 4451
rect 3843 4447 3844 4451
rect 3886 4448 3887 4452
rect 3891 4448 3892 4452
rect 3886 4447 3892 4448
rect 4182 4452 4188 4453
rect 4182 4448 4183 4452
rect 4187 4448 4188 4452
rect 4182 4447 4188 4448
rect 4510 4452 4516 4453
rect 4510 4448 4511 4452
rect 4515 4448 4516 4452
rect 4510 4447 4516 4448
rect 4846 4452 4852 4453
rect 4846 4448 4847 4452
rect 4851 4448 4852 4452
rect 4846 4447 4852 4448
rect 5190 4452 5196 4453
rect 5190 4448 5191 4452
rect 5195 4448 5196 4452
rect 5190 4447 5196 4448
rect 5542 4452 5548 4453
rect 5542 4448 5543 4452
rect 5547 4448 5548 4452
rect 5542 4447 5548 4448
rect 5662 4451 5668 4452
rect 5662 4447 5663 4451
rect 5667 4447 5668 4451
rect 3838 4446 3844 4447
rect 5662 4446 5668 4447
rect 1994 4445 2000 4446
rect 1974 4444 1980 4445
rect 1974 4440 1975 4444
rect 1979 4440 1980 4444
rect 1994 4441 1995 4445
rect 1999 4441 2000 4445
rect 1994 4440 2000 4441
rect 2130 4445 2136 4446
rect 2130 4441 2131 4445
rect 2135 4441 2136 4445
rect 2130 4440 2136 4441
rect 2266 4445 2272 4446
rect 2266 4441 2267 4445
rect 2271 4441 2272 4445
rect 2266 4440 2272 4441
rect 2402 4445 2408 4446
rect 2402 4441 2403 4445
rect 2407 4441 2408 4445
rect 2402 4440 2408 4441
rect 2538 4445 2544 4446
rect 2538 4441 2539 4445
rect 2543 4441 2544 4445
rect 2538 4440 2544 4441
rect 2674 4445 2680 4446
rect 2674 4441 2675 4445
rect 2679 4441 2680 4445
rect 2674 4440 2680 4441
rect 2810 4445 2816 4446
rect 2810 4441 2811 4445
rect 2815 4441 2816 4445
rect 2810 4440 2816 4441
rect 2946 4445 2952 4446
rect 2946 4441 2947 4445
rect 2951 4441 2952 4445
rect 2946 4440 2952 4441
rect 3798 4444 3804 4445
rect 3798 4440 3799 4444
rect 3803 4440 3804 4444
rect 1974 4439 1980 4440
rect 3798 4439 3804 4440
rect 110 4417 116 4418
rect 1934 4417 1940 4418
rect 110 4413 111 4417
rect 115 4413 116 4417
rect 110 4412 116 4413
rect 518 4416 524 4417
rect 518 4412 519 4416
rect 523 4412 524 4416
rect 518 4411 524 4412
rect 742 4416 748 4417
rect 742 4412 743 4416
rect 747 4412 748 4416
rect 742 4411 748 4412
rect 990 4416 996 4417
rect 990 4412 991 4416
rect 995 4412 996 4416
rect 990 4411 996 4412
rect 1262 4416 1268 4417
rect 1262 4412 1263 4416
rect 1267 4412 1268 4416
rect 1262 4411 1268 4412
rect 1550 4416 1556 4417
rect 1550 4412 1551 4416
rect 1555 4412 1556 4416
rect 1550 4411 1556 4412
rect 1814 4416 1820 4417
rect 1814 4412 1815 4416
rect 1819 4412 1820 4416
rect 1934 4413 1935 4417
rect 1939 4413 1940 4417
rect 1934 4412 1940 4413
rect 1814 4411 1820 4412
rect 490 4401 496 4402
rect 110 4400 116 4401
rect 110 4396 111 4400
rect 115 4396 116 4400
rect 490 4397 491 4401
rect 495 4397 496 4401
rect 490 4396 496 4397
rect 714 4401 720 4402
rect 714 4397 715 4401
rect 719 4397 720 4401
rect 714 4396 720 4397
rect 962 4401 968 4402
rect 962 4397 963 4401
rect 967 4397 968 4401
rect 962 4396 968 4397
rect 1234 4401 1240 4402
rect 1234 4397 1235 4401
rect 1239 4397 1240 4401
rect 1234 4396 1240 4397
rect 1522 4401 1528 4402
rect 1522 4397 1523 4401
rect 1527 4397 1528 4401
rect 1522 4396 1528 4397
rect 1786 4401 1792 4402
rect 1786 4397 1787 4401
rect 1791 4397 1792 4401
rect 1786 4396 1792 4397
rect 1934 4400 1940 4401
rect 1934 4396 1935 4400
rect 1939 4396 1940 4400
rect 110 4395 116 4396
rect 1934 4395 1940 4396
rect 3838 4393 3844 4394
rect 5662 4393 5668 4394
rect 3838 4389 3839 4393
rect 3843 4389 3844 4393
rect 3838 4388 3844 4389
rect 3886 4392 3892 4393
rect 3886 4388 3887 4392
rect 3891 4388 3892 4392
rect 3886 4387 3892 4388
rect 4142 4392 4148 4393
rect 4142 4388 4143 4392
rect 4147 4388 4148 4392
rect 4142 4387 4148 4388
rect 4422 4392 4428 4393
rect 4422 4388 4423 4392
rect 4427 4388 4428 4392
rect 4422 4387 4428 4388
rect 4702 4392 4708 4393
rect 4702 4388 4703 4392
rect 4707 4388 4708 4392
rect 4702 4387 4708 4388
rect 4982 4392 4988 4393
rect 4982 4388 4983 4392
rect 4987 4388 4988 4392
rect 4982 4387 4988 4388
rect 5262 4392 5268 4393
rect 5262 4388 5263 4392
rect 5267 4388 5268 4392
rect 5262 4387 5268 4388
rect 5542 4392 5548 4393
rect 5542 4388 5543 4392
rect 5547 4388 5548 4392
rect 5662 4389 5663 4393
rect 5667 4389 5668 4393
rect 5662 4388 5668 4389
rect 5542 4387 5548 4388
rect 3858 4377 3864 4378
rect 3838 4376 3844 4377
rect 3838 4372 3839 4376
rect 3843 4372 3844 4376
rect 3858 4373 3859 4377
rect 3863 4373 3864 4377
rect 3858 4372 3864 4373
rect 4114 4377 4120 4378
rect 4114 4373 4115 4377
rect 4119 4373 4120 4377
rect 4114 4372 4120 4373
rect 4394 4377 4400 4378
rect 4394 4373 4395 4377
rect 4399 4373 4400 4377
rect 4394 4372 4400 4373
rect 4674 4377 4680 4378
rect 4674 4373 4675 4377
rect 4679 4373 4680 4377
rect 4674 4372 4680 4373
rect 4954 4377 4960 4378
rect 4954 4373 4955 4377
rect 4959 4373 4960 4377
rect 4954 4372 4960 4373
rect 5234 4377 5240 4378
rect 5234 4373 5235 4377
rect 5239 4373 5240 4377
rect 5234 4372 5240 4373
rect 5514 4377 5520 4378
rect 5514 4373 5515 4377
rect 5519 4373 5520 4377
rect 5514 4372 5520 4373
rect 5662 4376 5668 4377
rect 5662 4372 5663 4376
rect 5667 4372 5668 4376
rect 3838 4371 3844 4372
rect 5662 4371 5668 4372
rect 1974 4296 1980 4297
rect 3798 4296 3804 4297
rect 1974 4292 1975 4296
rect 1979 4292 1980 4296
rect 1974 4291 1980 4292
rect 2778 4295 2784 4296
rect 2778 4291 2779 4295
rect 2783 4291 2784 4295
rect 2778 4290 2784 4291
rect 2994 4295 3000 4296
rect 2994 4291 2995 4295
rect 2999 4291 3000 4295
rect 2994 4290 3000 4291
rect 3218 4295 3224 4296
rect 3218 4291 3219 4295
rect 3223 4291 3224 4295
rect 3218 4290 3224 4291
rect 3442 4295 3448 4296
rect 3442 4291 3443 4295
rect 3447 4291 3448 4295
rect 3442 4290 3448 4291
rect 3650 4295 3656 4296
rect 3650 4291 3651 4295
rect 3655 4291 3656 4295
rect 3798 4292 3799 4296
rect 3803 4292 3804 4296
rect 3798 4291 3804 4292
rect 3650 4290 3656 4291
rect 2806 4280 2812 4281
rect 1974 4279 1980 4280
rect 1974 4275 1975 4279
rect 1979 4275 1980 4279
rect 2806 4276 2807 4280
rect 2811 4276 2812 4280
rect 2806 4275 2812 4276
rect 3022 4280 3028 4281
rect 3022 4276 3023 4280
rect 3027 4276 3028 4280
rect 3022 4275 3028 4276
rect 3246 4280 3252 4281
rect 3246 4276 3247 4280
rect 3251 4276 3252 4280
rect 3246 4275 3252 4276
rect 3470 4280 3476 4281
rect 3470 4276 3471 4280
rect 3475 4276 3476 4280
rect 3470 4275 3476 4276
rect 3678 4280 3684 4281
rect 3678 4276 3679 4280
rect 3683 4276 3684 4280
rect 3678 4275 3684 4276
rect 3798 4279 3804 4280
rect 3798 4275 3799 4279
rect 3803 4275 3804 4279
rect 1974 4274 1980 4275
rect 3798 4274 3804 4275
rect 110 4268 116 4269
rect 1934 4268 1940 4269
rect 110 4264 111 4268
rect 115 4264 116 4268
rect 110 4263 116 4264
rect 562 4267 568 4268
rect 562 4263 563 4267
rect 567 4263 568 4267
rect 562 4262 568 4263
rect 698 4267 704 4268
rect 698 4263 699 4267
rect 703 4263 704 4267
rect 698 4262 704 4263
rect 834 4267 840 4268
rect 834 4263 835 4267
rect 839 4263 840 4267
rect 834 4262 840 4263
rect 970 4267 976 4268
rect 970 4263 971 4267
rect 975 4263 976 4267
rect 970 4262 976 4263
rect 1106 4267 1112 4268
rect 1106 4263 1107 4267
rect 1111 4263 1112 4267
rect 1106 4262 1112 4263
rect 1242 4267 1248 4268
rect 1242 4263 1243 4267
rect 1247 4263 1248 4267
rect 1242 4262 1248 4263
rect 1378 4267 1384 4268
rect 1378 4263 1379 4267
rect 1383 4263 1384 4267
rect 1378 4262 1384 4263
rect 1514 4267 1520 4268
rect 1514 4263 1515 4267
rect 1519 4263 1520 4267
rect 1514 4262 1520 4263
rect 1650 4267 1656 4268
rect 1650 4263 1651 4267
rect 1655 4263 1656 4267
rect 1650 4262 1656 4263
rect 1786 4267 1792 4268
rect 1786 4263 1787 4267
rect 1791 4263 1792 4267
rect 1934 4264 1935 4268
rect 1939 4264 1940 4268
rect 1934 4263 1940 4264
rect 1786 4262 1792 4263
rect 590 4252 596 4253
rect 110 4251 116 4252
rect 110 4247 111 4251
rect 115 4247 116 4251
rect 590 4248 591 4252
rect 595 4248 596 4252
rect 590 4247 596 4248
rect 726 4252 732 4253
rect 726 4248 727 4252
rect 731 4248 732 4252
rect 726 4247 732 4248
rect 862 4252 868 4253
rect 862 4248 863 4252
rect 867 4248 868 4252
rect 862 4247 868 4248
rect 998 4252 1004 4253
rect 998 4248 999 4252
rect 1003 4248 1004 4252
rect 998 4247 1004 4248
rect 1134 4252 1140 4253
rect 1134 4248 1135 4252
rect 1139 4248 1140 4252
rect 1134 4247 1140 4248
rect 1270 4252 1276 4253
rect 1270 4248 1271 4252
rect 1275 4248 1276 4252
rect 1270 4247 1276 4248
rect 1406 4252 1412 4253
rect 1406 4248 1407 4252
rect 1411 4248 1412 4252
rect 1406 4247 1412 4248
rect 1542 4252 1548 4253
rect 1542 4248 1543 4252
rect 1547 4248 1548 4252
rect 1542 4247 1548 4248
rect 1678 4252 1684 4253
rect 1678 4248 1679 4252
rect 1683 4248 1684 4252
rect 1678 4247 1684 4248
rect 1814 4252 1820 4253
rect 1814 4248 1815 4252
rect 1819 4248 1820 4252
rect 1814 4247 1820 4248
rect 1934 4251 1940 4252
rect 1934 4247 1935 4251
rect 1939 4247 1940 4251
rect 110 4246 116 4247
rect 1934 4246 1940 4247
rect 3838 4232 3844 4233
rect 5662 4232 5668 4233
rect 3838 4228 3839 4232
rect 3843 4228 3844 4232
rect 3838 4227 3844 4228
rect 4570 4231 4576 4232
rect 4570 4227 4571 4231
rect 4575 4227 4576 4231
rect 4570 4226 4576 4227
rect 4738 4231 4744 4232
rect 4738 4227 4739 4231
rect 4743 4227 4744 4231
rect 4738 4226 4744 4227
rect 4914 4231 4920 4232
rect 4914 4227 4915 4231
rect 4919 4227 4920 4231
rect 4914 4226 4920 4227
rect 5106 4231 5112 4232
rect 5106 4227 5107 4231
rect 5111 4227 5112 4231
rect 5106 4226 5112 4227
rect 5306 4231 5312 4232
rect 5306 4227 5307 4231
rect 5311 4227 5312 4231
rect 5306 4226 5312 4227
rect 5514 4231 5520 4232
rect 5514 4227 5515 4231
rect 5519 4227 5520 4231
rect 5662 4228 5663 4232
rect 5667 4228 5668 4232
rect 5662 4227 5668 4228
rect 5514 4226 5520 4227
rect 4598 4216 4604 4217
rect 3838 4215 3844 4216
rect 3838 4211 3839 4215
rect 3843 4211 3844 4215
rect 4598 4212 4599 4216
rect 4603 4212 4604 4216
rect 4598 4211 4604 4212
rect 4766 4216 4772 4217
rect 4766 4212 4767 4216
rect 4771 4212 4772 4216
rect 4766 4211 4772 4212
rect 4942 4216 4948 4217
rect 4942 4212 4943 4216
rect 4947 4212 4948 4216
rect 4942 4211 4948 4212
rect 5134 4216 5140 4217
rect 5134 4212 5135 4216
rect 5139 4212 5140 4216
rect 5134 4211 5140 4212
rect 5334 4216 5340 4217
rect 5334 4212 5335 4216
rect 5339 4212 5340 4216
rect 5334 4211 5340 4212
rect 5542 4216 5548 4217
rect 5542 4212 5543 4216
rect 5547 4212 5548 4216
rect 5542 4211 5548 4212
rect 5662 4215 5668 4216
rect 5662 4211 5663 4215
rect 5667 4211 5668 4215
rect 3838 4210 3844 4211
rect 5662 4210 5668 4211
rect 1974 4193 1980 4194
rect 3798 4193 3804 4194
rect 1974 4189 1975 4193
rect 1979 4189 1980 4193
rect 1974 4188 1980 4189
rect 2950 4192 2956 4193
rect 2950 4188 2951 4192
rect 2955 4188 2956 4192
rect 2950 4187 2956 4188
rect 3094 4192 3100 4193
rect 3094 4188 3095 4192
rect 3099 4188 3100 4192
rect 3094 4187 3100 4188
rect 3238 4192 3244 4193
rect 3238 4188 3239 4192
rect 3243 4188 3244 4192
rect 3238 4187 3244 4188
rect 3390 4192 3396 4193
rect 3390 4188 3391 4192
rect 3395 4188 3396 4192
rect 3390 4187 3396 4188
rect 3542 4192 3548 4193
rect 3542 4188 3543 4192
rect 3547 4188 3548 4192
rect 3542 4187 3548 4188
rect 3678 4192 3684 4193
rect 3678 4188 3679 4192
rect 3683 4188 3684 4192
rect 3798 4189 3799 4193
rect 3803 4189 3804 4193
rect 3798 4188 3804 4189
rect 3678 4187 3684 4188
rect 110 4181 116 4182
rect 1934 4181 1940 4182
rect 110 4177 111 4181
rect 115 4177 116 4181
rect 110 4176 116 4177
rect 590 4180 596 4181
rect 590 4176 591 4180
rect 595 4176 596 4180
rect 590 4175 596 4176
rect 726 4180 732 4181
rect 726 4176 727 4180
rect 731 4176 732 4180
rect 726 4175 732 4176
rect 862 4180 868 4181
rect 862 4176 863 4180
rect 867 4176 868 4180
rect 862 4175 868 4176
rect 998 4180 1004 4181
rect 998 4176 999 4180
rect 1003 4176 1004 4180
rect 998 4175 1004 4176
rect 1134 4180 1140 4181
rect 1134 4176 1135 4180
rect 1139 4176 1140 4180
rect 1134 4175 1140 4176
rect 1270 4180 1276 4181
rect 1270 4176 1271 4180
rect 1275 4176 1276 4180
rect 1270 4175 1276 4176
rect 1406 4180 1412 4181
rect 1406 4176 1407 4180
rect 1411 4176 1412 4180
rect 1406 4175 1412 4176
rect 1542 4180 1548 4181
rect 1542 4176 1543 4180
rect 1547 4176 1548 4180
rect 1542 4175 1548 4176
rect 1678 4180 1684 4181
rect 1678 4176 1679 4180
rect 1683 4176 1684 4180
rect 1678 4175 1684 4176
rect 1814 4180 1820 4181
rect 1814 4176 1815 4180
rect 1819 4176 1820 4180
rect 1934 4177 1935 4181
rect 1939 4177 1940 4181
rect 2922 4177 2928 4178
rect 1934 4176 1940 4177
rect 1974 4176 1980 4177
rect 1814 4175 1820 4176
rect 1974 4172 1975 4176
rect 1979 4172 1980 4176
rect 2922 4173 2923 4177
rect 2927 4173 2928 4177
rect 2922 4172 2928 4173
rect 3066 4177 3072 4178
rect 3066 4173 3067 4177
rect 3071 4173 3072 4177
rect 3066 4172 3072 4173
rect 3210 4177 3216 4178
rect 3210 4173 3211 4177
rect 3215 4173 3216 4177
rect 3210 4172 3216 4173
rect 3362 4177 3368 4178
rect 3362 4173 3363 4177
rect 3367 4173 3368 4177
rect 3362 4172 3368 4173
rect 3514 4177 3520 4178
rect 3514 4173 3515 4177
rect 3519 4173 3520 4177
rect 3514 4172 3520 4173
rect 3650 4177 3656 4178
rect 3650 4173 3651 4177
rect 3655 4173 3656 4177
rect 3650 4172 3656 4173
rect 3798 4176 3804 4177
rect 3798 4172 3799 4176
rect 3803 4172 3804 4176
rect 1974 4171 1980 4172
rect 3798 4171 3804 4172
rect 562 4165 568 4166
rect 110 4164 116 4165
rect 110 4160 111 4164
rect 115 4160 116 4164
rect 562 4161 563 4165
rect 567 4161 568 4165
rect 562 4160 568 4161
rect 698 4165 704 4166
rect 698 4161 699 4165
rect 703 4161 704 4165
rect 698 4160 704 4161
rect 834 4165 840 4166
rect 834 4161 835 4165
rect 839 4161 840 4165
rect 834 4160 840 4161
rect 970 4165 976 4166
rect 970 4161 971 4165
rect 975 4161 976 4165
rect 970 4160 976 4161
rect 1106 4165 1112 4166
rect 1106 4161 1107 4165
rect 1111 4161 1112 4165
rect 1106 4160 1112 4161
rect 1242 4165 1248 4166
rect 1242 4161 1243 4165
rect 1247 4161 1248 4165
rect 1242 4160 1248 4161
rect 1378 4165 1384 4166
rect 1378 4161 1379 4165
rect 1383 4161 1384 4165
rect 1378 4160 1384 4161
rect 1514 4165 1520 4166
rect 1514 4161 1515 4165
rect 1519 4161 1520 4165
rect 1514 4160 1520 4161
rect 1650 4165 1656 4166
rect 1650 4161 1651 4165
rect 1655 4161 1656 4165
rect 1650 4160 1656 4161
rect 1786 4165 1792 4166
rect 1786 4161 1787 4165
rect 1791 4161 1792 4165
rect 1786 4160 1792 4161
rect 1934 4164 1940 4165
rect 1934 4160 1935 4164
rect 1939 4160 1940 4164
rect 110 4159 116 4160
rect 1934 4159 1940 4160
rect 3838 4157 3844 4158
rect 5662 4157 5668 4158
rect 3838 4153 3839 4157
rect 3843 4153 3844 4157
rect 3838 4152 3844 4153
rect 4654 4156 4660 4157
rect 4654 4152 4655 4156
rect 4659 4152 4660 4156
rect 4654 4151 4660 4152
rect 4814 4156 4820 4157
rect 4814 4152 4815 4156
rect 4819 4152 4820 4156
rect 4814 4151 4820 4152
rect 4982 4156 4988 4157
rect 4982 4152 4983 4156
rect 4987 4152 4988 4156
rect 4982 4151 4988 4152
rect 5166 4156 5172 4157
rect 5166 4152 5167 4156
rect 5171 4152 5172 4156
rect 5166 4151 5172 4152
rect 5358 4156 5364 4157
rect 5358 4152 5359 4156
rect 5363 4152 5364 4156
rect 5358 4151 5364 4152
rect 5542 4156 5548 4157
rect 5542 4152 5543 4156
rect 5547 4152 5548 4156
rect 5662 4153 5663 4157
rect 5667 4153 5668 4157
rect 5662 4152 5668 4153
rect 5542 4151 5548 4152
rect 4626 4141 4632 4142
rect 3838 4140 3844 4141
rect 3838 4136 3839 4140
rect 3843 4136 3844 4140
rect 4626 4137 4627 4141
rect 4631 4137 4632 4141
rect 4626 4136 4632 4137
rect 4786 4141 4792 4142
rect 4786 4137 4787 4141
rect 4791 4137 4792 4141
rect 4786 4136 4792 4137
rect 4954 4141 4960 4142
rect 4954 4137 4955 4141
rect 4959 4137 4960 4141
rect 4954 4136 4960 4137
rect 5138 4141 5144 4142
rect 5138 4137 5139 4141
rect 5143 4137 5144 4141
rect 5138 4136 5144 4137
rect 5330 4141 5336 4142
rect 5330 4137 5331 4141
rect 5335 4137 5336 4141
rect 5330 4136 5336 4137
rect 5514 4141 5520 4142
rect 5514 4137 5515 4141
rect 5519 4137 5520 4141
rect 5514 4136 5520 4137
rect 5662 4140 5668 4141
rect 5662 4136 5663 4140
rect 5667 4136 5668 4140
rect 3838 4135 3844 4136
rect 5662 4135 5668 4136
rect 110 4032 116 4033
rect 1934 4032 1940 4033
rect 110 4028 111 4032
rect 115 4028 116 4032
rect 110 4027 116 4028
rect 698 4031 704 4032
rect 698 4027 699 4031
rect 703 4027 704 4031
rect 698 4026 704 4027
rect 834 4031 840 4032
rect 834 4027 835 4031
rect 839 4027 840 4031
rect 834 4026 840 4027
rect 970 4031 976 4032
rect 970 4027 971 4031
rect 975 4027 976 4031
rect 970 4026 976 4027
rect 1106 4031 1112 4032
rect 1106 4027 1107 4031
rect 1111 4027 1112 4031
rect 1106 4026 1112 4027
rect 1242 4031 1248 4032
rect 1242 4027 1243 4031
rect 1247 4027 1248 4031
rect 1242 4026 1248 4027
rect 1378 4031 1384 4032
rect 1378 4027 1379 4031
rect 1383 4027 1384 4031
rect 1378 4026 1384 4027
rect 1514 4031 1520 4032
rect 1514 4027 1515 4031
rect 1519 4027 1520 4031
rect 1514 4026 1520 4027
rect 1650 4031 1656 4032
rect 1650 4027 1651 4031
rect 1655 4027 1656 4031
rect 1650 4026 1656 4027
rect 1786 4031 1792 4032
rect 1786 4027 1787 4031
rect 1791 4027 1792 4031
rect 1934 4028 1935 4032
rect 1939 4028 1940 4032
rect 1934 4027 1940 4028
rect 1786 4026 1792 4027
rect 726 4016 732 4017
rect 110 4015 116 4016
rect 110 4011 111 4015
rect 115 4011 116 4015
rect 726 4012 727 4016
rect 731 4012 732 4016
rect 726 4011 732 4012
rect 862 4016 868 4017
rect 862 4012 863 4016
rect 867 4012 868 4016
rect 862 4011 868 4012
rect 998 4016 1004 4017
rect 998 4012 999 4016
rect 1003 4012 1004 4016
rect 998 4011 1004 4012
rect 1134 4016 1140 4017
rect 1134 4012 1135 4016
rect 1139 4012 1140 4016
rect 1134 4011 1140 4012
rect 1270 4016 1276 4017
rect 1270 4012 1271 4016
rect 1275 4012 1276 4016
rect 1270 4011 1276 4012
rect 1406 4016 1412 4017
rect 1406 4012 1407 4016
rect 1411 4012 1412 4016
rect 1406 4011 1412 4012
rect 1542 4016 1548 4017
rect 1542 4012 1543 4016
rect 1547 4012 1548 4016
rect 1542 4011 1548 4012
rect 1678 4016 1684 4017
rect 1678 4012 1679 4016
rect 1683 4012 1684 4016
rect 1678 4011 1684 4012
rect 1814 4016 1820 4017
rect 1814 4012 1815 4016
rect 1819 4012 1820 4016
rect 1814 4011 1820 4012
rect 1934 4015 1940 4016
rect 1934 4011 1935 4015
rect 1939 4011 1940 4015
rect 110 4010 116 4011
rect 1934 4010 1940 4011
rect 1974 4008 1980 4009
rect 3798 4008 3804 4009
rect 1974 4004 1975 4008
rect 1979 4004 1980 4008
rect 1974 4003 1980 4004
rect 2898 4007 2904 4008
rect 2898 4003 2899 4007
rect 2903 4003 2904 4007
rect 2898 4002 2904 4003
rect 3042 4007 3048 4008
rect 3042 4003 3043 4007
rect 3047 4003 3048 4007
rect 3042 4002 3048 4003
rect 3186 4007 3192 4008
rect 3186 4003 3187 4007
rect 3191 4003 3192 4007
rect 3186 4002 3192 4003
rect 3338 4007 3344 4008
rect 3338 4003 3339 4007
rect 3343 4003 3344 4007
rect 3338 4002 3344 4003
rect 3490 4007 3496 4008
rect 3490 4003 3491 4007
rect 3495 4003 3496 4007
rect 3490 4002 3496 4003
rect 3642 4007 3648 4008
rect 3642 4003 3643 4007
rect 3647 4003 3648 4007
rect 3798 4004 3799 4008
rect 3803 4004 3804 4008
rect 3798 4003 3804 4004
rect 3642 4002 3648 4003
rect 2926 3992 2932 3993
rect 1974 3991 1980 3992
rect 1974 3987 1975 3991
rect 1979 3987 1980 3991
rect 2926 3988 2927 3992
rect 2931 3988 2932 3992
rect 2926 3987 2932 3988
rect 3070 3992 3076 3993
rect 3070 3988 3071 3992
rect 3075 3988 3076 3992
rect 3070 3987 3076 3988
rect 3214 3992 3220 3993
rect 3214 3988 3215 3992
rect 3219 3988 3220 3992
rect 3214 3987 3220 3988
rect 3366 3992 3372 3993
rect 3366 3988 3367 3992
rect 3371 3988 3372 3992
rect 3366 3987 3372 3988
rect 3518 3992 3524 3993
rect 3518 3988 3519 3992
rect 3523 3988 3524 3992
rect 3518 3987 3524 3988
rect 3670 3992 3676 3993
rect 3670 3988 3671 3992
rect 3675 3988 3676 3992
rect 3670 3987 3676 3988
rect 3798 3991 3804 3992
rect 3798 3987 3799 3991
rect 3803 3987 3804 3991
rect 1974 3986 1980 3987
rect 3798 3986 3804 3987
rect 3838 3972 3844 3973
rect 5662 3972 5668 3973
rect 3838 3968 3839 3972
rect 3843 3968 3844 3972
rect 3838 3967 3844 3968
rect 4938 3971 4944 3972
rect 4938 3967 4939 3971
rect 4943 3967 4944 3971
rect 4938 3966 4944 3967
rect 5074 3971 5080 3972
rect 5074 3967 5075 3971
rect 5079 3967 5080 3971
rect 5074 3966 5080 3967
rect 5210 3971 5216 3972
rect 5210 3967 5211 3971
rect 5215 3967 5216 3971
rect 5210 3966 5216 3967
rect 5346 3971 5352 3972
rect 5346 3967 5347 3971
rect 5351 3967 5352 3971
rect 5662 3968 5663 3972
rect 5667 3968 5668 3972
rect 5662 3967 5668 3968
rect 5346 3966 5352 3967
rect 4966 3956 4972 3957
rect 3838 3955 3844 3956
rect 110 3953 116 3954
rect 1934 3953 1940 3954
rect 110 3949 111 3953
rect 115 3949 116 3953
rect 110 3948 116 3949
rect 694 3952 700 3953
rect 694 3948 695 3952
rect 699 3948 700 3952
rect 694 3947 700 3948
rect 830 3952 836 3953
rect 830 3948 831 3952
rect 835 3948 836 3952
rect 830 3947 836 3948
rect 966 3952 972 3953
rect 966 3948 967 3952
rect 971 3948 972 3952
rect 966 3947 972 3948
rect 1110 3952 1116 3953
rect 1110 3948 1111 3952
rect 1115 3948 1116 3952
rect 1110 3947 1116 3948
rect 1254 3952 1260 3953
rect 1254 3948 1255 3952
rect 1259 3948 1260 3952
rect 1254 3947 1260 3948
rect 1398 3952 1404 3953
rect 1398 3948 1399 3952
rect 1403 3948 1404 3952
rect 1398 3947 1404 3948
rect 1542 3952 1548 3953
rect 1542 3948 1543 3952
rect 1547 3948 1548 3952
rect 1542 3947 1548 3948
rect 1678 3952 1684 3953
rect 1678 3948 1679 3952
rect 1683 3948 1684 3952
rect 1678 3947 1684 3948
rect 1814 3952 1820 3953
rect 1814 3948 1815 3952
rect 1819 3948 1820 3952
rect 1934 3949 1935 3953
rect 1939 3949 1940 3953
rect 3838 3951 3839 3955
rect 3843 3951 3844 3955
rect 4966 3952 4967 3956
rect 4971 3952 4972 3956
rect 4966 3951 4972 3952
rect 5102 3956 5108 3957
rect 5102 3952 5103 3956
rect 5107 3952 5108 3956
rect 5102 3951 5108 3952
rect 5238 3956 5244 3957
rect 5238 3952 5239 3956
rect 5243 3952 5244 3956
rect 5238 3951 5244 3952
rect 5374 3956 5380 3957
rect 5374 3952 5375 3956
rect 5379 3952 5380 3956
rect 5374 3951 5380 3952
rect 5662 3955 5668 3956
rect 5662 3951 5663 3955
rect 5667 3951 5668 3955
rect 3838 3950 3844 3951
rect 5662 3950 5668 3951
rect 1934 3948 1940 3949
rect 1814 3947 1820 3948
rect 666 3937 672 3938
rect 110 3936 116 3937
rect 110 3932 111 3936
rect 115 3932 116 3936
rect 666 3933 667 3937
rect 671 3933 672 3937
rect 666 3932 672 3933
rect 802 3937 808 3938
rect 802 3933 803 3937
rect 807 3933 808 3937
rect 802 3932 808 3933
rect 938 3937 944 3938
rect 938 3933 939 3937
rect 943 3933 944 3937
rect 938 3932 944 3933
rect 1082 3937 1088 3938
rect 1082 3933 1083 3937
rect 1087 3933 1088 3937
rect 1082 3932 1088 3933
rect 1226 3937 1232 3938
rect 1226 3933 1227 3937
rect 1231 3933 1232 3937
rect 1226 3932 1232 3933
rect 1370 3937 1376 3938
rect 1370 3933 1371 3937
rect 1375 3933 1376 3937
rect 1370 3932 1376 3933
rect 1514 3937 1520 3938
rect 1514 3933 1515 3937
rect 1519 3933 1520 3937
rect 1514 3932 1520 3933
rect 1650 3937 1656 3938
rect 1650 3933 1651 3937
rect 1655 3933 1656 3937
rect 1650 3932 1656 3933
rect 1786 3937 1792 3938
rect 1786 3933 1787 3937
rect 1791 3933 1792 3937
rect 1786 3932 1792 3933
rect 1934 3936 1940 3937
rect 1934 3932 1935 3936
rect 1939 3932 1940 3936
rect 110 3931 116 3932
rect 1934 3931 1940 3932
rect 1974 3905 1980 3906
rect 3798 3905 3804 3906
rect 1974 3901 1975 3905
rect 1979 3901 1980 3905
rect 1974 3900 1980 3901
rect 2758 3904 2764 3905
rect 2758 3900 2759 3904
rect 2763 3900 2764 3904
rect 2758 3899 2764 3900
rect 2910 3904 2916 3905
rect 2910 3900 2911 3904
rect 2915 3900 2916 3904
rect 2910 3899 2916 3900
rect 3070 3904 3076 3905
rect 3070 3900 3071 3904
rect 3075 3900 3076 3904
rect 3070 3899 3076 3900
rect 3238 3904 3244 3905
rect 3238 3900 3239 3904
rect 3243 3900 3244 3904
rect 3238 3899 3244 3900
rect 3414 3904 3420 3905
rect 3414 3900 3415 3904
rect 3419 3900 3420 3904
rect 3414 3899 3420 3900
rect 3590 3904 3596 3905
rect 3590 3900 3591 3904
rect 3595 3900 3596 3904
rect 3798 3901 3799 3905
rect 3803 3901 3804 3905
rect 3798 3900 3804 3901
rect 3590 3899 3596 3900
rect 3838 3897 3844 3898
rect 5662 3897 5668 3898
rect 3838 3893 3839 3897
rect 3843 3893 3844 3897
rect 3838 3892 3844 3893
rect 4686 3896 4692 3897
rect 4686 3892 4687 3896
rect 4691 3892 4692 3896
rect 4686 3891 4692 3892
rect 4846 3896 4852 3897
rect 4846 3892 4847 3896
rect 4851 3892 4852 3896
rect 4846 3891 4852 3892
rect 5014 3896 5020 3897
rect 5014 3892 5015 3896
rect 5019 3892 5020 3896
rect 5014 3891 5020 3892
rect 5190 3896 5196 3897
rect 5190 3892 5191 3896
rect 5195 3892 5196 3896
rect 5190 3891 5196 3892
rect 5374 3896 5380 3897
rect 5374 3892 5375 3896
rect 5379 3892 5380 3896
rect 5374 3891 5380 3892
rect 5542 3896 5548 3897
rect 5542 3892 5543 3896
rect 5547 3892 5548 3896
rect 5662 3893 5663 3897
rect 5667 3893 5668 3897
rect 5662 3892 5668 3893
rect 5542 3891 5548 3892
rect 2730 3889 2736 3890
rect 1974 3888 1980 3889
rect 1974 3884 1975 3888
rect 1979 3884 1980 3888
rect 2730 3885 2731 3889
rect 2735 3885 2736 3889
rect 2730 3884 2736 3885
rect 2882 3889 2888 3890
rect 2882 3885 2883 3889
rect 2887 3885 2888 3889
rect 2882 3884 2888 3885
rect 3042 3889 3048 3890
rect 3042 3885 3043 3889
rect 3047 3885 3048 3889
rect 3042 3884 3048 3885
rect 3210 3889 3216 3890
rect 3210 3885 3211 3889
rect 3215 3885 3216 3889
rect 3210 3884 3216 3885
rect 3386 3889 3392 3890
rect 3386 3885 3387 3889
rect 3391 3885 3392 3889
rect 3386 3884 3392 3885
rect 3562 3889 3568 3890
rect 3562 3885 3563 3889
rect 3567 3885 3568 3889
rect 3562 3884 3568 3885
rect 3798 3888 3804 3889
rect 3798 3884 3799 3888
rect 3803 3884 3804 3888
rect 1974 3883 1980 3884
rect 3798 3883 3804 3884
rect 4658 3881 4664 3882
rect 3838 3880 3844 3881
rect 3838 3876 3839 3880
rect 3843 3876 3844 3880
rect 4658 3877 4659 3881
rect 4663 3877 4664 3881
rect 4658 3876 4664 3877
rect 4818 3881 4824 3882
rect 4818 3877 4819 3881
rect 4823 3877 4824 3881
rect 4818 3876 4824 3877
rect 4986 3881 4992 3882
rect 4986 3877 4987 3881
rect 4991 3877 4992 3881
rect 4986 3876 4992 3877
rect 5162 3881 5168 3882
rect 5162 3877 5163 3881
rect 5167 3877 5168 3881
rect 5162 3876 5168 3877
rect 5346 3881 5352 3882
rect 5346 3877 5347 3881
rect 5351 3877 5352 3881
rect 5346 3876 5352 3877
rect 5514 3881 5520 3882
rect 5514 3877 5515 3881
rect 5519 3877 5520 3881
rect 5514 3876 5520 3877
rect 5662 3880 5668 3881
rect 5662 3876 5663 3880
rect 5667 3876 5668 3880
rect 3838 3875 3844 3876
rect 5662 3875 5668 3876
rect 110 3800 116 3801
rect 1934 3800 1940 3801
rect 110 3796 111 3800
rect 115 3796 116 3800
rect 110 3795 116 3796
rect 434 3799 440 3800
rect 434 3795 435 3799
rect 439 3795 440 3799
rect 434 3794 440 3795
rect 618 3799 624 3800
rect 618 3795 619 3799
rect 623 3795 624 3799
rect 618 3794 624 3795
rect 818 3799 824 3800
rect 818 3795 819 3799
rect 823 3795 824 3799
rect 818 3794 824 3795
rect 1026 3799 1032 3800
rect 1026 3795 1027 3799
rect 1031 3795 1032 3799
rect 1026 3794 1032 3795
rect 1250 3799 1256 3800
rect 1250 3795 1251 3799
rect 1255 3795 1256 3799
rect 1250 3794 1256 3795
rect 1482 3799 1488 3800
rect 1482 3795 1483 3799
rect 1487 3795 1488 3799
rect 1482 3794 1488 3795
rect 1722 3799 1728 3800
rect 1722 3795 1723 3799
rect 1727 3795 1728 3799
rect 1934 3796 1935 3800
rect 1939 3796 1940 3800
rect 1934 3795 1940 3796
rect 1722 3794 1728 3795
rect 462 3784 468 3785
rect 110 3783 116 3784
rect 110 3779 111 3783
rect 115 3779 116 3783
rect 462 3780 463 3784
rect 467 3780 468 3784
rect 462 3779 468 3780
rect 646 3784 652 3785
rect 646 3780 647 3784
rect 651 3780 652 3784
rect 646 3779 652 3780
rect 846 3784 852 3785
rect 846 3780 847 3784
rect 851 3780 852 3784
rect 846 3779 852 3780
rect 1054 3784 1060 3785
rect 1054 3780 1055 3784
rect 1059 3780 1060 3784
rect 1054 3779 1060 3780
rect 1278 3784 1284 3785
rect 1278 3780 1279 3784
rect 1283 3780 1284 3784
rect 1278 3779 1284 3780
rect 1510 3784 1516 3785
rect 1510 3780 1511 3784
rect 1515 3780 1516 3784
rect 1510 3779 1516 3780
rect 1750 3784 1756 3785
rect 1750 3780 1751 3784
rect 1755 3780 1756 3784
rect 1750 3779 1756 3780
rect 1934 3783 1940 3784
rect 1934 3779 1935 3783
rect 1939 3779 1940 3783
rect 110 3778 116 3779
rect 1934 3778 1940 3779
rect 1974 3748 1980 3749
rect 3798 3748 3804 3749
rect 1974 3744 1975 3748
rect 1979 3744 1980 3748
rect 1974 3743 1980 3744
rect 2114 3747 2120 3748
rect 2114 3743 2115 3747
rect 2119 3743 2120 3747
rect 2114 3742 2120 3743
rect 2250 3747 2256 3748
rect 2250 3743 2251 3747
rect 2255 3743 2256 3747
rect 2250 3742 2256 3743
rect 2386 3747 2392 3748
rect 2386 3743 2387 3747
rect 2391 3743 2392 3747
rect 2386 3742 2392 3743
rect 2522 3747 2528 3748
rect 2522 3743 2523 3747
rect 2527 3743 2528 3747
rect 2522 3742 2528 3743
rect 2658 3747 2664 3748
rect 2658 3743 2659 3747
rect 2663 3743 2664 3747
rect 2658 3742 2664 3743
rect 2794 3747 2800 3748
rect 2794 3743 2795 3747
rect 2799 3743 2800 3747
rect 2794 3742 2800 3743
rect 2938 3747 2944 3748
rect 2938 3743 2939 3747
rect 2943 3743 2944 3747
rect 2938 3742 2944 3743
rect 3082 3747 3088 3748
rect 3082 3743 3083 3747
rect 3087 3743 3088 3747
rect 3082 3742 3088 3743
rect 3234 3747 3240 3748
rect 3234 3743 3235 3747
rect 3239 3743 3240 3747
rect 3234 3742 3240 3743
rect 3394 3747 3400 3748
rect 3394 3743 3395 3747
rect 3399 3743 3400 3747
rect 3394 3742 3400 3743
rect 3554 3747 3560 3748
rect 3554 3743 3555 3747
rect 3559 3743 3560 3747
rect 3798 3744 3799 3748
rect 3803 3744 3804 3748
rect 3798 3743 3804 3744
rect 3838 3748 3844 3749
rect 5662 3748 5668 3749
rect 3838 3744 3839 3748
rect 3843 3744 3844 3748
rect 3838 3743 3844 3744
rect 4410 3747 4416 3748
rect 4410 3743 4411 3747
rect 4415 3743 4416 3747
rect 3554 3742 3560 3743
rect 4410 3742 4416 3743
rect 4618 3747 4624 3748
rect 4618 3743 4619 3747
rect 4623 3743 4624 3747
rect 4618 3742 4624 3743
rect 4834 3747 4840 3748
rect 4834 3743 4835 3747
rect 4839 3743 4840 3747
rect 4834 3742 4840 3743
rect 5066 3747 5072 3748
rect 5066 3743 5067 3747
rect 5071 3743 5072 3747
rect 5066 3742 5072 3743
rect 5298 3747 5304 3748
rect 5298 3743 5299 3747
rect 5303 3743 5304 3747
rect 5298 3742 5304 3743
rect 5514 3747 5520 3748
rect 5514 3743 5515 3747
rect 5519 3743 5520 3747
rect 5662 3744 5663 3748
rect 5667 3744 5668 3748
rect 5662 3743 5668 3744
rect 5514 3742 5520 3743
rect 2142 3732 2148 3733
rect 1974 3731 1980 3732
rect 1974 3727 1975 3731
rect 1979 3727 1980 3731
rect 2142 3728 2143 3732
rect 2147 3728 2148 3732
rect 2142 3727 2148 3728
rect 2278 3732 2284 3733
rect 2278 3728 2279 3732
rect 2283 3728 2284 3732
rect 2278 3727 2284 3728
rect 2414 3732 2420 3733
rect 2414 3728 2415 3732
rect 2419 3728 2420 3732
rect 2414 3727 2420 3728
rect 2550 3732 2556 3733
rect 2550 3728 2551 3732
rect 2555 3728 2556 3732
rect 2550 3727 2556 3728
rect 2686 3732 2692 3733
rect 2686 3728 2687 3732
rect 2691 3728 2692 3732
rect 2686 3727 2692 3728
rect 2822 3732 2828 3733
rect 2822 3728 2823 3732
rect 2827 3728 2828 3732
rect 2822 3727 2828 3728
rect 2966 3732 2972 3733
rect 2966 3728 2967 3732
rect 2971 3728 2972 3732
rect 2966 3727 2972 3728
rect 3110 3732 3116 3733
rect 3110 3728 3111 3732
rect 3115 3728 3116 3732
rect 3110 3727 3116 3728
rect 3262 3732 3268 3733
rect 3262 3728 3263 3732
rect 3267 3728 3268 3732
rect 3262 3727 3268 3728
rect 3422 3732 3428 3733
rect 3422 3728 3423 3732
rect 3427 3728 3428 3732
rect 3422 3727 3428 3728
rect 3582 3732 3588 3733
rect 4438 3732 4444 3733
rect 3582 3728 3583 3732
rect 3587 3728 3588 3732
rect 3582 3727 3588 3728
rect 3798 3731 3804 3732
rect 3798 3727 3799 3731
rect 3803 3727 3804 3731
rect 1974 3726 1980 3727
rect 3798 3726 3804 3727
rect 3838 3731 3844 3732
rect 3838 3727 3839 3731
rect 3843 3727 3844 3731
rect 4438 3728 4439 3732
rect 4443 3728 4444 3732
rect 4438 3727 4444 3728
rect 4646 3732 4652 3733
rect 4646 3728 4647 3732
rect 4651 3728 4652 3732
rect 4646 3727 4652 3728
rect 4862 3732 4868 3733
rect 4862 3728 4863 3732
rect 4867 3728 4868 3732
rect 4862 3727 4868 3728
rect 5094 3732 5100 3733
rect 5094 3728 5095 3732
rect 5099 3728 5100 3732
rect 5094 3727 5100 3728
rect 5326 3732 5332 3733
rect 5326 3728 5327 3732
rect 5331 3728 5332 3732
rect 5326 3727 5332 3728
rect 5542 3732 5548 3733
rect 5542 3728 5543 3732
rect 5547 3728 5548 3732
rect 5542 3727 5548 3728
rect 5662 3731 5668 3732
rect 5662 3727 5663 3731
rect 5667 3727 5668 3731
rect 3838 3726 3844 3727
rect 5662 3726 5668 3727
rect 110 3721 116 3722
rect 1934 3721 1940 3722
rect 110 3717 111 3721
rect 115 3717 116 3721
rect 110 3716 116 3717
rect 230 3720 236 3721
rect 230 3716 231 3720
rect 235 3716 236 3720
rect 230 3715 236 3716
rect 430 3720 436 3721
rect 430 3716 431 3720
rect 435 3716 436 3720
rect 430 3715 436 3716
rect 654 3720 660 3721
rect 654 3716 655 3720
rect 659 3716 660 3720
rect 654 3715 660 3716
rect 894 3720 900 3721
rect 894 3716 895 3720
rect 899 3716 900 3720
rect 894 3715 900 3716
rect 1150 3720 1156 3721
rect 1150 3716 1151 3720
rect 1155 3716 1156 3720
rect 1150 3715 1156 3716
rect 1414 3720 1420 3721
rect 1414 3716 1415 3720
rect 1419 3716 1420 3720
rect 1414 3715 1420 3716
rect 1678 3720 1684 3721
rect 1678 3716 1679 3720
rect 1683 3716 1684 3720
rect 1934 3717 1935 3721
rect 1939 3717 1940 3721
rect 1934 3716 1940 3717
rect 1678 3715 1684 3716
rect 202 3705 208 3706
rect 110 3704 116 3705
rect 110 3700 111 3704
rect 115 3700 116 3704
rect 202 3701 203 3705
rect 207 3701 208 3705
rect 202 3700 208 3701
rect 402 3705 408 3706
rect 402 3701 403 3705
rect 407 3701 408 3705
rect 402 3700 408 3701
rect 626 3705 632 3706
rect 626 3701 627 3705
rect 631 3701 632 3705
rect 626 3700 632 3701
rect 866 3705 872 3706
rect 866 3701 867 3705
rect 871 3701 872 3705
rect 866 3700 872 3701
rect 1122 3705 1128 3706
rect 1122 3701 1123 3705
rect 1127 3701 1128 3705
rect 1122 3700 1128 3701
rect 1386 3705 1392 3706
rect 1386 3701 1387 3705
rect 1391 3701 1392 3705
rect 1386 3700 1392 3701
rect 1650 3705 1656 3706
rect 1650 3701 1651 3705
rect 1655 3701 1656 3705
rect 1650 3700 1656 3701
rect 1934 3704 1940 3705
rect 1934 3700 1935 3704
rect 1939 3700 1940 3704
rect 110 3699 116 3700
rect 1934 3699 1940 3700
rect 1974 3665 1980 3666
rect 3798 3665 3804 3666
rect 1974 3661 1975 3665
rect 1979 3661 1980 3665
rect 1974 3660 1980 3661
rect 2230 3664 2236 3665
rect 2230 3660 2231 3664
rect 2235 3660 2236 3664
rect 2230 3659 2236 3660
rect 2446 3664 2452 3665
rect 2446 3660 2447 3664
rect 2451 3660 2452 3664
rect 2446 3659 2452 3660
rect 2662 3664 2668 3665
rect 2662 3660 2663 3664
rect 2667 3660 2668 3664
rect 2662 3659 2668 3660
rect 2870 3664 2876 3665
rect 2870 3660 2871 3664
rect 2875 3660 2876 3664
rect 2870 3659 2876 3660
rect 3078 3664 3084 3665
rect 3078 3660 3079 3664
rect 3083 3660 3084 3664
rect 3078 3659 3084 3660
rect 3286 3664 3292 3665
rect 3286 3660 3287 3664
rect 3291 3660 3292 3664
rect 3286 3659 3292 3660
rect 3494 3664 3500 3665
rect 3494 3660 3495 3664
rect 3499 3660 3500 3664
rect 3494 3659 3500 3660
rect 3678 3664 3684 3665
rect 3678 3660 3679 3664
rect 3683 3660 3684 3664
rect 3798 3661 3799 3665
rect 3803 3661 3804 3665
rect 3798 3660 3804 3661
rect 3678 3659 3684 3660
rect 2202 3649 2208 3650
rect 1974 3648 1980 3649
rect 1974 3644 1975 3648
rect 1979 3644 1980 3648
rect 2202 3645 2203 3649
rect 2207 3645 2208 3649
rect 2202 3644 2208 3645
rect 2418 3649 2424 3650
rect 2418 3645 2419 3649
rect 2423 3645 2424 3649
rect 2418 3644 2424 3645
rect 2634 3649 2640 3650
rect 2634 3645 2635 3649
rect 2639 3645 2640 3649
rect 2634 3644 2640 3645
rect 2842 3649 2848 3650
rect 2842 3645 2843 3649
rect 2847 3645 2848 3649
rect 2842 3644 2848 3645
rect 3050 3649 3056 3650
rect 3050 3645 3051 3649
rect 3055 3645 3056 3649
rect 3050 3644 3056 3645
rect 3258 3649 3264 3650
rect 3258 3645 3259 3649
rect 3263 3645 3264 3649
rect 3258 3644 3264 3645
rect 3466 3649 3472 3650
rect 3466 3645 3467 3649
rect 3471 3645 3472 3649
rect 3466 3644 3472 3645
rect 3650 3649 3656 3650
rect 3838 3649 3844 3650
rect 5662 3649 5668 3650
rect 3650 3645 3651 3649
rect 3655 3645 3656 3649
rect 3650 3644 3656 3645
rect 3798 3648 3804 3649
rect 3798 3644 3799 3648
rect 3803 3644 3804 3648
rect 3838 3645 3839 3649
rect 3843 3645 3844 3649
rect 3838 3644 3844 3645
rect 3886 3648 3892 3649
rect 3886 3644 3887 3648
rect 3891 3644 3892 3648
rect 1974 3643 1980 3644
rect 3798 3643 3804 3644
rect 3886 3643 3892 3644
rect 4046 3648 4052 3649
rect 4046 3644 4047 3648
rect 4051 3644 4052 3648
rect 4046 3643 4052 3644
rect 4246 3648 4252 3649
rect 4246 3644 4247 3648
rect 4251 3644 4252 3648
rect 4246 3643 4252 3644
rect 4478 3648 4484 3649
rect 4478 3644 4479 3648
rect 4483 3644 4484 3648
rect 4478 3643 4484 3644
rect 4726 3648 4732 3649
rect 4726 3644 4727 3648
rect 4731 3644 4732 3648
rect 4726 3643 4732 3644
rect 4998 3648 5004 3649
rect 4998 3644 4999 3648
rect 5003 3644 5004 3648
rect 4998 3643 5004 3644
rect 5278 3648 5284 3649
rect 5278 3644 5279 3648
rect 5283 3644 5284 3648
rect 5278 3643 5284 3644
rect 5542 3648 5548 3649
rect 5542 3644 5543 3648
rect 5547 3644 5548 3648
rect 5662 3645 5663 3649
rect 5667 3645 5668 3649
rect 5662 3644 5668 3645
rect 5542 3643 5548 3644
rect 3858 3633 3864 3634
rect 3838 3632 3844 3633
rect 3838 3628 3839 3632
rect 3843 3628 3844 3632
rect 3858 3629 3859 3633
rect 3863 3629 3864 3633
rect 3858 3628 3864 3629
rect 4018 3633 4024 3634
rect 4018 3629 4019 3633
rect 4023 3629 4024 3633
rect 4018 3628 4024 3629
rect 4218 3633 4224 3634
rect 4218 3629 4219 3633
rect 4223 3629 4224 3633
rect 4218 3628 4224 3629
rect 4450 3633 4456 3634
rect 4450 3629 4451 3633
rect 4455 3629 4456 3633
rect 4450 3628 4456 3629
rect 4698 3633 4704 3634
rect 4698 3629 4699 3633
rect 4703 3629 4704 3633
rect 4698 3628 4704 3629
rect 4970 3633 4976 3634
rect 4970 3629 4971 3633
rect 4975 3629 4976 3633
rect 4970 3628 4976 3629
rect 5250 3633 5256 3634
rect 5250 3629 5251 3633
rect 5255 3629 5256 3633
rect 5250 3628 5256 3629
rect 5514 3633 5520 3634
rect 5514 3629 5515 3633
rect 5519 3629 5520 3633
rect 5514 3628 5520 3629
rect 5662 3632 5668 3633
rect 5662 3628 5663 3632
rect 5667 3628 5668 3632
rect 3838 3627 3844 3628
rect 5662 3627 5668 3628
rect 110 3564 116 3565
rect 1934 3564 1940 3565
rect 110 3560 111 3564
rect 115 3560 116 3564
rect 110 3559 116 3560
rect 130 3563 136 3564
rect 130 3559 131 3563
rect 135 3559 136 3563
rect 130 3558 136 3559
rect 314 3563 320 3564
rect 314 3559 315 3563
rect 319 3559 320 3563
rect 314 3558 320 3559
rect 538 3563 544 3564
rect 538 3559 539 3563
rect 543 3559 544 3563
rect 538 3558 544 3559
rect 786 3563 792 3564
rect 786 3559 787 3563
rect 791 3559 792 3563
rect 786 3558 792 3559
rect 1042 3563 1048 3564
rect 1042 3559 1043 3563
rect 1047 3559 1048 3563
rect 1042 3558 1048 3559
rect 1314 3563 1320 3564
rect 1314 3559 1315 3563
rect 1319 3559 1320 3563
rect 1314 3558 1320 3559
rect 1586 3563 1592 3564
rect 1586 3559 1587 3563
rect 1591 3559 1592 3563
rect 1934 3560 1935 3564
rect 1939 3560 1940 3564
rect 1934 3559 1940 3560
rect 1586 3558 1592 3559
rect 158 3548 164 3549
rect 110 3547 116 3548
rect 110 3543 111 3547
rect 115 3543 116 3547
rect 158 3544 159 3548
rect 163 3544 164 3548
rect 158 3543 164 3544
rect 342 3548 348 3549
rect 342 3544 343 3548
rect 347 3544 348 3548
rect 342 3543 348 3544
rect 566 3548 572 3549
rect 566 3544 567 3548
rect 571 3544 572 3548
rect 566 3543 572 3544
rect 814 3548 820 3549
rect 814 3544 815 3548
rect 819 3544 820 3548
rect 814 3543 820 3544
rect 1070 3548 1076 3549
rect 1070 3544 1071 3548
rect 1075 3544 1076 3548
rect 1070 3543 1076 3544
rect 1342 3548 1348 3549
rect 1342 3544 1343 3548
rect 1347 3544 1348 3548
rect 1342 3543 1348 3544
rect 1614 3548 1620 3549
rect 1614 3544 1615 3548
rect 1619 3544 1620 3548
rect 1614 3543 1620 3544
rect 1934 3547 1940 3548
rect 1934 3543 1935 3547
rect 1939 3543 1940 3547
rect 110 3542 116 3543
rect 1934 3542 1940 3543
rect 1974 3500 1980 3501
rect 3798 3500 3804 3501
rect 1974 3496 1975 3500
rect 1979 3496 1980 3500
rect 1974 3495 1980 3496
rect 2162 3499 2168 3500
rect 2162 3495 2163 3499
rect 2167 3495 2168 3499
rect 2162 3494 2168 3495
rect 2298 3499 2304 3500
rect 2298 3495 2299 3499
rect 2303 3495 2304 3499
rect 2298 3494 2304 3495
rect 2434 3499 2440 3500
rect 2434 3495 2435 3499
rect 2439 3495 2440 3499
rect 2434 3494 2440 3495
rect 2570 3499 2576 3500
rect 2570 3495 2571 3499
rect 2575 3495 2576 3499
rect 3798 3496 3799 3500
rect 3803 3496 3804 3500
rect 3798 3495 3804 3496
rect 2570 3494 2576 3495
rect 3838 3488 3844 3489
rect 5662 3488 5668 3489
rect 2190 3484 2196 3485
rect 1974 3483 1980 3484
rect 1974 3479 1975 3483
rect 1979 3479 1980 3483
rect 2190 3480 2191 3484
rect 2195 3480 2196 3484
rect 2190 3479 2196 3480
rect 2326 3484 2332 3485
rect 2326 3480 2327 3484
rect 2331 3480 2332 3484
rect 2326 3479 2332 3480
rect 2462 3484 2468 3485
rect 2462 3480 2463 3484
rect 2467 3480 2468 3484
rect 2462 3479 2468 3480
rect 2598 3484 2604 3485
rect 3838 3484 3839 3488
rect 3843 3484 3844 3488
rect 2598 3480 2599 3484
rect 2603 3480 2604 3484
rect 2598 3479 2604 3480
rect 3798 3483 3804 3484
rect 3838 3483 3844 3484
rect 3858 3487 3864 3488
rect 3858 3483 3859 3487
rect 3863 3483 3864 3487
rect 3798 3479 3799 3483
rect 3803 3479 3804 3483
rect 3858 3482 3864 3483
rect 3994 3487 4000 3488
rect 3994 3483 3995 3487
rect 3999 3483 4000 3487
rect 3994 3482 4000 3483
rect 4130 3487 4136 3488
rect 4130 3483 4131 3487
rect 4135 3483 4136 3487
rect 4130 3482 4136 3483
rect 4266 3487 4272 3488
rect 4266 3483 4267 3487
rect 4271 3483 4272 3487
rect 4266 3482 4272 3483
rect 4402 3487 4408 3488
rect 4402 3483 4403 3487
rect 4407 3483 4408 3487
rect 4402 3482 4408 3483
rect 4538 3487 4544 3488
rect 4538 3483 4539 3487
rect 4543 3483 4544 3487
rect 4538 3482 4544 3483
rect 4698 3487 4704 3488
rect 4698 3483 4699 3487
rect 4703 3483 4704 3487
rect 4698 3482 4704 3483
rect 4890 3487 4896 3488
rect 4890 3483 4891 3487
rect 4895 3483 4896 3487
rect 4890 3482 4896 3483
rect 5098 3487 5104 3488
rect 5098 3483 5099 3487
rect 5103 3483 5104 3487
rect 5098 3482 5104 3483
rect 5314 3487 5320 3488
rect 5314 3483 5315 3487
rect 5319 3483 5320 3487
rect 5314 3482 5320 3483
rect 5514 3487 5520 3488
rect 5514 3483 5515 3487
rect 5519 3483 5520 3487
rect 5662 3484 5663 3488
rect 5667 3484 5668 3488
rect 5662 3483 5668 3484
rect 5514 3482 5520 3483
rect 1974 3478 1980 3479
rect 3798 3478 3804 3479
rect 110 3477 116 3478
rect 1934 3477 1940 3478
rect 110 3473 111 3477
rect 115 3473 116 3477
rect 110 3472 116 3473
rect 158 3476 164 3477
rect 158 3472 159 3476
rect 163 3472 164 3476
rect 158 3471 164 3472
rect 334 3476 340 3477
rect 334 3472 335 3476
rect 339 3472 340 3476
rect 334 3471 340 3472
rect 550 3476 556 3477
rect 550 3472 551 3476
rect 555 3472 556 3476
rect 550 3471 556 3472
rect 790 3476 796 3477
rect 790 3472 791 3476
rect 795 3472 796 3476
rect 790 3471 796 3472
rect 1038 3476 1044 3477
rect 1038 3472 1039 3476
rect 1043 3472 1044 3476
rect 1038 3471 1044 3472
rect 1294 3476 1300 3477
rect 1294 3472 1295 3476
rect 1299 3472 1300 3476
rect 1294 3471 1300 3472
rect 1558 3476 1564 3477
rect 1558 3472 1559 3476
rect 1563 3472 1564 3476
rect 1934 3473 1935 3477
rect 1939 3473 1940 3477
rect 1934 3472 1940 3473
rect 3886 3472 3892 3473
rect 1558 3471 1564 3472
rect 3838 3471 3844 3472
rect 3838 3467 3839 3471
rect 3843 3467 3844 3471
rect 3886 3468 3887 3472
rect 3891 3468 3892 3472
rect 3886 3467 3892 3468
rect 4022 3472 4028 3473
rect 4022 3468 4023 3472
rect 4027 3468 4028 3472
rect 4022 3467 4028 3468
rect 4158 3472 4164 3473
rect 4158 3468 4159 3472
rect 4163 3468 4164 3472
rect 4158 3467 4164 3468
rect 4294 3472 4300 3473
rect 4294 3468 4295 3472
rect 4299 3468 4300 3472
rect 4294 3467 4300 3468
rect 4430 3472 4436 3473
rect 4430 3468 4431 3472
rect 4435 3468 4436 3472
rect 4430 3467 4436 3468
rect 4566 3472 4572 3473
rect 4566 3468 4567 3472
rect 4571 3468 4572 3472
rect 4566 3467 4572 3468
rect 4726 3472 4732 3473
rect 4726 3468 4727 3472
rect 4731 3468 4732 3472
rect 4726 3467 4732 3468
rect 4918 3472 4924 3473
rect 4918 3468 4919 3472
rect 4923 3468 4924 3472
rect 4918 3467 4924 3468
rect 5126 3472 5132 3473
rect 5126 3468 5127 3472
rect 5131 3468 5132 3472
rect 5126 3467 5132 3468
rect 5342 3472 5348 3473
rect 5342 3468 5343 3472
rect 5347 3468 5348 3472
rect 5342 3467 5348 3468
rect 5542 3472 5548 3473
rect 5542 3468 5543 3472
rect 5547 3468 5548 3472
rect 5542 3467 5548 3468
rect 5662 3471 5668 3472
rect 5662 3467 5663 3471
rect 5667 3467 5668 3471
rect 3838 3466 3844 3467
rect 5662 3466 5668 3467
rect 130 3461 136 3462
rect 110 3460 116 3461
rect 110 3456 111 3460
rect 115 3456 116 3460
rect 130 3457 131 3461
rect 135 3457 136 3461
rect 130 3456 136 3457
rect 306 3461 312 3462
rect 306 3457 307 3461
rect 311 3457 312 3461
rect 306 3456 312 3457
rect 522 3461 528 3462
rect 522 3457 523 3461
rect 527 3457 528 3461
rect 522 3456 528 3457
rect 762 3461 768 3462
rect 762 3457 763 3461
rect 767 3457 768 3461
rect 762 3456 768 3457
rect 1010 3461 1016 3462
rect 1010 3457 1011 3461
rect 1015 3457 1016 3461
rect 1010 3456 1016 3457
rect 1266 3461 1272 3462
rect 1266 3457 1267 3461
rect 1271 3457 1272 3461
rect 1266 3456 1272 3457
rect 1530 3461 1536 3462
rect 1530 3457 1531 3461
rect 1535 3457 1536 3461
rect 1530 3456 1536 3457
rect 1934 3460 1940 3461
rect 1934 3456 1935 3460
rect 1939 3456 1940 3460
rect 110 3455 116 3456
rect 1934 3455 1940 3456
rect 3838 3405 3844 3406
rect 5662 3405 5668 3406
rect 3838 3401 3839 3405
rect 3843 3401 3844 3405
rect 3838 3400 3844 3401
rect 3886 3404 3892 3405
rect 3886 3400 3887 3404
rect 3891 3400 3892 3404
rect 3886 3399 3892 3400
rect 4022 3404 4028 3405
rect 4022 3400 4023 3404
rect 4027 3400 4028 3404
rect 4022 3399 4028 3400
rect 4158 3404 4164 3405
rect 4158 3400 4159 3404
rect 4163 3400 4164 3404
rect 4158 3399 4164 3400
rect 4294 3404 4300 3405
rect 4294 3400 4295 3404
rect 4299 3400 4300 3404
rect 4294 3399 4300 3400
rect 4430 3404 4436 3405
rect 4430 3400 4431 3404
rect 4435 3400 4436 3404
rect 4430 3399 4436 3400
rect 4582 3404 4588 3405
rect 4582 3400 4583 3404
rect 4587 3400 4588 3404
rect 4582 3399 4588 3400
rect 4758 3404 4764 3405
rect 4758 3400 4759 3404
rect 4763 3400 4764 3404
rect 4758 3399 4764 3400
rect 4950 3404 4956 3405
rect 4950 3400 4951 3404
rect 4955 3400 4956 3404
rect 4950 3399 4956 3400
rect 5150 3404 5156 3405
rect 5150 3400 5151 3404
rect 5155 3400 5156 3404
rect 5150 3399 5156 3400
rect 5358 3404 5364 3405
rect 5358 3400 5359 3404
rect 5363 3400 5364 3404
rect 5358 3399 5364 3400
rect 5542 3404 5548 3405
rect 5542 3400 5543 3404
rect 5547 3400 5548 3404
rect 5662 3401 5663 3405
rect 5667 3401 5668 3405
rect 5662 3400 5668 3401
rect 5542 3399 5548 3400
rect 1974 3389 1980 3390
rect 3798 3389 3804 3390
rect 3858 3389 3864 3390
rect 1974 3385 1975 3389
rect 1979 3385 1980 3389
rect 1974 3384 1980 3385
rect 2230 3388 2236 3389
rect 2230 3384 2231 3388
rect 2235 3384 2236 3388
rect 2230 3383 2236 3384
rect 2582 3388 2588 3389
rect 2582 3384 2583 3388
rect 2587 3384 2588 3388
rect 2582 3383 2588 3384
rect 2950 3388 2956 3389
rect 2950 3384 2951 3388
rect 2955 3384 2956 3388
rect 2950 3383 2956 3384
rect 3326 3388 3332 3389
rect 3326 3384 3327 3388
rect 3331 3384 3332 3388
rect 3326 3383 3332 3384
rect 3678 3388 3684 3389
rect 3678 3384 3679 3388
rect 3683 3384 3684 3388
rect 3798 3385 3799 3389
rect 3803 3385 3804 3389
rect 3798 3384 3804 3385
rect 3838 3388 3844 3389
rect 3838 3384 3839 3388
rect 3843 3384 3844 3388
rect 3858 3385 3859 3389
rect 3863 3385 3864 3389
rect 3858 3384 3864 3385
rect 3994 3389 4000 3390
rect 3994 3385 3995 3389
rect 3999 3385 4000 3389
rect 3994 3384 4000 3385
rect 4130 3389 4136 3390
rect 4130 3385 4131 3389
rect 4135 3385 4136 3389
rect 4130 3384 4136 3385
rect 4266 3389 4272 3390
rect 4266 3385 4267 3389
rect 4271 3385 4272 3389
rect 4266 3384 4272 3385
rect 4402 3389 4408 3390
rect 4402 3385 4403 3389
rect 4407 3385 4408 3389
rect 4402 3384 4408 3385
rect 4554 3389 4560 3390
rect 4554 3385 4555 3389
rect 4559 3385 4560 3389
rect 4554 3384 4560 3385
rect 4730 3389 4736 3390
rect 4730 3385 4731 3389
rect 4735 3385 4736 3389
rect 4730 3384 4736 3385
rect 4922 3389 4928 3390
rect 4922 3385 4923 3389
rect 4927 3385 4928 3389
rect 4922 3384 4928 3385
rect 5122 3389 5128 3390
rect 5122 3385 5123 3389
rect 5127 3385 5128 3389
rect 5122 3384 5128 3385
rect 5330 3389 5336 3390
rect 5330 3385 5331 3389
rect 5335 3385 5336 3389
rect 5330 3384 5336 3385
rect 5514 3389 5520 3390
rect 5514 3385 5515 3389
rect 5519 3385 5520 3389
rect 5514 3384 5520 3385
rect 5662 3388 5668 3389
rect 5662 3384 5663 3388
rect 5667 3384 5668 3388
rect 3678 3383 3684 3384
rect 3838 3383 3844 3384
rect 5662 3383 5668 3384
rect 2202 3373 2208 3374
rect 1974 3372 1980 3373
rect 1974 3368 1975 3372
rect 1979 3368 1980 3372
rect 2202 3369 2203 3373
rect 2207 3369 2208 3373
rect 2202 3368 2208 3369
rect 2554 3373 2560 3374
rect 2554 3369 2555 3373
rect 2559 3369 2560 3373
rect 2554 3368 2560 3369
rect 2922 3373 2928 3374
rect 2922 3369 2923 3373
rect 2927 3369 2928 3373
rect 2922 3368 2928 3369
rect 3298 3373 3304 3374
rect 3298 3369 3299 3373
rect 3303 3369 3304 3373
rect 3298 3368 3304 3369
rect 3650 3373 3656 3374
rect 3650 3369 3651 3373
rect 3655 3369 3656 3373
rect 3650 3368 3656 3369
rect 3798 3372 3804 3373
rect 3798 3368 3799 3372
rect 3803 3368 3804 3372
rect 1974 3367 1980 3368
rect 3798 3367 3804 3368
rect 110 3320 116 3321
rect 1934 3320 1940 3321
rect 110 3316 111 3320
rect 115 3316 116 3320
rect 110 3315 116 3316
rect 130 3319 136 3320
rect 130 3315 131 3319
rect 135 3315 136 3319
rect 130 3314 136 3315
rect 298 3319 304 3320
rect 298 3315 299 3319
rect 303 3315 304 3319
rect 298 3314 304 3315
rect 506 3319 512 3320
rect 506 3315 507 3319
rect 511 3315 512 3319
rect 506 3314 512 3315
rect 730 3319 736 3320
rect 730 3315 731 3319
rect 735 3315 736 3319
rect 730 3314 736 3315
rect 970 3319 976 3320
rect 970 3315 971 3319
rect 975 3315 976 3319
rect 970 3314 976 3315
rect 1218 3319 1224 3320
rect 1218 3315 1219 3319
rect 1223 3315 1224 3319
rect 1218 3314 1224 3315
rect 1474 3319 1480 3320
rect 1474 3315 1475 3319
rect 1479 3315 1480 3319
rect 1934 3316 1935 3320
rect 1939 3316 1940 3320
rect 1934 3315 1940 3316
rect 1474 3314 1480 3315
rect 158 3304 164 3305
rect 110 3303 116 3304
rect 110 3299 111 3303
rect 115 3299 116 3303
rect 158 3300 159 3304
rect 163 3300 164 3304
rect 158 3299 164 3300
rect 326 3304 332 3305
rect 326 3300 327 3304
rect 331 3300 332 3304
rect 326 3299 332 3300
rect 534 3304 540 3305
rect 534 3300 535 3304
rect 539 3300 540 3304
rect 534 3299 540 3300
rect 758 3304 764 3305
rect 758 3300 759 3304
rect 763 3300 764 3304
rect 758 3299 764 3300
rect 998 3304 1004 3305
rect 998 3300 999 3304
rect 1003 3300 1004 3304
rect 998 3299 1004 3300
rect 1246 3304 1252 3305
rect 1246 3300 1247 3304
rect 1251 3300 1252 3304
rect 1246 3299 1252 3300
rect 1502 3304 1508 3305
rect 1502 3300 1503 3304
rect 1507 3300 1508 3304
rect 1502 3299 1508 3300
rect 1934 3303 1940 3304
rect 1934 3299 1935 3303
rect 1939 3299 1940 3303
rect 110 3298 116 3299
rect 1934 3298 1940 3299
rect 110 3241 116 3242
rect 1934 3241 1940 3242
rect 110 3237 111 3241
rect 115 3237 116 3241
rect 110 3236 116 3237
rect 238 3240 244 3241
rect 238 3236 239 3240
rect 243 3236 244 3240
rect 238 3235 244 3236
rect 462 3240 468 3241
rect 462 3236 463 3240
rect 467 3236 468 3240
rect 462 3235 468 3236
rect 702 3240 708 3241
rect 702 3236 703 3240
rect 707 3236 708 3240
rect 702 3235 708 3236
rect 950 3240 956 3241
rect 950 3236 951 3240
rect 955 3236 956 3240
rect 950 3235 956 3236
rect 1198 3240 1204 3241
rect 1198 3236 1199 3240
rect 1203 3236 1204 3240
rect 1198 3235 1204 3236
rect 1454 3240 1460 3241
rect 1454 3236 1455 3240
rect 1459 3236 1460 3240
rect 1934 3237 1935 3241
rect 1939 3237 1940 3241
rect 1934 3236 1940 3237
rect 1974 3240 1980 3241
rect 3798 3240 3804 3241
rect 1974 3236 1975 3240
rect 1979 3236 1980 3240
rect 1454 3235 1460 3236
rect 1974 3235 1980 3236
rect 2250 3239 2256 3240
rect 2250 3235 2251 3239
rect 2255 3235 2256 3239
rect 2250 3234 2256 3235
rect 2474 3239 2480 3240
rect 2474 3235 2475 3239
rect 2479 3235 2480 3239
rect 2474 3234 2480 3235
rect 2690 3239 2696 3240
rect 2690 3235 2691 3239
rect 2695 3235 2696 3239
rect 2690 3234 2696 3235
rect 2898 3239 2904 3240
rect 2898 3235 2899 3239
rect 2903 3235 2904 3239
rect 2898 3234 2904 3235
rect 3098 3239 3104 3240
rect 3098 3235 3099 3239
rect 3103 3235 3104 3239
rect 3098 3234 3104 3235
rect 3290 3239 3296 3240
rect 3290 3235 3291 3239
rect 3295 3235 3296 3239
rect 3290 3234 3296 3235
rect 3482 3239 3488 3240
rect 3482 3235 3483 3239
rect 3487 3235 3488 3239
rect 3482 3234 3488 3235
rect 3650 3239 3656 3240
rect 3650 3235 3651 3239
rect 3655 3235 3656 3239
rect 3798 3236 3799 3240
rect 3803 3236 3804 3240
rect 3798 3235 3804 3236
rect 3838 3240 3844 3241
rect 5662 3240 5668 3241
rect 3838 3236 3839 3240
rect 3843 3236 3844 3240
rect 3838 3235 3844 3236
rect 4690 3239 4696 3240
rect 4690 3235 4691 3239
rect 4695 3235 4696 3239
rect 3650 3234 3656 3235
rect 4690 3234 4696 3235
rect 4826 3239 4832 3240
rect 4826 3235 4827 3239
rect 4831 3235 4832 3239
rect 4826 3234 4832 3235
rect 4962 3239 4968 3240
rect 4962 3235 4963 3239
rect 4967 3235 4968 3239
rect 4962 3234 4968 3235
rect 5098 3239 5104 3240
rect 5098 3235 5099 3239
rect 5103 3235 5104 3239
rect 5098 3234 5104 3235
rect 5234 3239 5240 3240
rect 5234 3235 5235 3239
rect 5239 3235 5240 3239
rect 5662 3236 5663 3240
rect 5667 3236 5668 3240
rect 5662 3235 5668 3236
rect 5234 3234 5240 3235
rect 210 3225 216 3226
rect 110 3224 116 3225
rect 110 3220 111 3224
rect 115 3220 116 3224
rect 210 3221 211 3225
rect 215 3221 216 3225
rect 210 3220 216 3221
rect 434 3225 440 3226
rect 434 3221 435 3225
rect 439 3221 440 3225
rect 434 3220 440 3221
rect 674 3225 680 3226
rect 674 3221 675 3225
rect 679 3221 680 3225
rect 674 3220 680 3221
rect 922 3225 928 3226
rect 922 3221 923 3225
rect 927 3221 928 3225
rect 922 3220 928 3221
rect 1170 3225 1176 3226
rect 1170 3221 1171 3225
rect 1175 3221 1176 3225
rect 1170 3220 1176 3221
rect 1426 3225 1432 3226
rect 1426 3221 1427 3225
rect 1431 3221 1432 3225
rect 1426 3220 1432 3221
rect 1934 3224 1940 3225
rect 2278 3224 2284 3225
rect 1934 3220 1935 3224
rect 1939 3220 1940 3224
rect 110 3219 116 3220
rect 1934 3219 1940 3220
rect 1974 3223 1980 3224
rect 1974 3219 1975 3223
rect 1979 3219 1980 3223
rect 2278 3220 2279 3224
rect 2283 3220 2284 3224
rect 2278 3219 2284 3220
rect 2502 3224 2508 3225
rect 2502 3220 2503 3224
rect 2507 3220 2508 3224
rect 2502 3219 2508 3220
rect 2718 3224 2724 3225
rect 2718 3220 2719 3224
rect 2723 3220 2724 3224
rect 2718 3219 2724 3220
rect 2926 3224 2932 3225
rect 2926 3220 2927 3224
rect 2931 3220 2932 3224
rect 2926 3219 2932 3220
rect 3126 3224 3132 3225
rect 3126 3220 3127 3224
rect 3131 3220 3132 3224
rect 3126 3219 3132 3220
rect 3318 3224 3324 3225
rect 3318 3220 3319 3224
rect 3323 3220 3324 3224
rect 3318 3219 3324 3220
rect 3510 3224 3516 3225
rect 3510 3220 3511 3224
rect 3515 3220 3516 3224
rect 3510 3219 3516 3220
rect 3678 3224 3684 3225
rect 4718 3224 4724 3225
rect 3678 3220 3679 3224
rect 3683 3220 3684 3224
rect 3678 3219 3684 3220
rect 3798 3223 3804 3224
rect 3798 3219 3799 3223
rect 3803 3219 3804 3223
rect 1974 3218 1980 3219
rect 3798 3218 3804 3219
rect 3838 3223 3844 3224
rect 3838 3219 3839 3223
rect 3843 3219 3844 3223
rect 4718 3220 4719 3224
rect 4723 3220 4724 3224
rect 4718 3219 4724 3220
rect 4854 3224 4860 3225
rect 4854 3220 4855 3224
rect 4859 3220 4860 3224
rect 4854 3219 4860 3220
rect 4990 3224 4996 3225
rect 4990 3220 4991 3224
rect 4995 3220 4996 3224
rect 4990 3219 4996 3220
rect 5126 3224 5132 3225
rect 5126 3220 5127 3224
rect 5131 3220 5132 3224
rect 5126 3219 5132 3220
rect 5262 3224 5268 3225
rect 5262 3220 5263 3224
rect 5267 3220 5268 3224
rect 5262 3219 5268 3220
rect 5662 3223 5668 3224
rect 5662 3219 5663 3223
rect 5667 3219 5668 3223
rect 3838 3218 3844 3219
rect 5662 3218 5668 3219
rect 1974 3157 1980 3158
rect 3798 3157 3804 3158
rect 1974 3153 1975 3157
rect 1979 3153 1980 3157
rect 1974 3152 1980 3153
rect 2094 3156 2100 3157
rect 2094 3152 2095 3156
rect 2099 3152 2100 3156
rect 2094 3151 2100 3152
rect 2294 3156 2300 3157
rect 2294 3152 2295 3156
rect 2299 3152 2300 3156
rect 2294 3151 2300 3152
rect 2486 3156 2492 3157
rect 2486 3152 2487 3156
rect 2491 3152 2492 3156
rect 2486 3151 2492 3152
rect 2678 3156 2684 3157
rect 2678 3152 2679 3156
rect 2683 3152 2684 3156
rect 2678 3151 2684 3152
rect 2870 3156 2876 3157
rect 2870 3152 2871 3156
rect 2875 3152 2876 3156
rect 2870 3151 2876 3152
rect 3054 3156 3060 3157
rect 3054 3152 3055 3156
rect 3059 3152 3060 3156
rect 3054 3151 3060 3152
rect 3230 3156 3236 3157
rect 3230 3152 3231 3156
rect 3235 3152 3236 3156
rect 3230 3151 3236 3152
rect 3414 3156 3420 3157
rect 3414 3152 3415 3156
rect 3419 3152 3420 3156
rect 3414 3151 3420 3152
rect 3598 3156 3604 3157
rect 3598 3152 3599 3156
rect 3603 3152 3604 3156
rect 3798 3153 3799 3157
rect 3803 3153 3804 3157
rect 3798 3152 3804 3153
rect 3838 3157 3844 3158
rect 5662 3157 5668 3158
rect 3838 3153 3839 3157
rect 3843 3153 3844 3157
rect 3838 3152 3844 3153
rect 4862 3156 4868 3157
rect 4862 3152 4863 3156
rect 4867 3152 4868 3156
rect 3598 3151 3604 3152
rect 4862 3151 4868 3152
rect 4998 3156 5004 3157
rect 4998 3152 4999 3156
rect 5003 3152 5004 3156
rect 4998 3151 5004 3152
rect 5134 3156 5140 3157
rect 5134 3152 5135 3156
rect 5139 3152 5140 3156
rect 5134 3151 5140 3152
rect 5270 3156 5276 3157
rect 5270 3152 5271 3156
rect 5275 3152 5276 3156
rect 5270 3151 5276 3152
rect 5406 3156 5412 3157
rect 5406 3152 5407 3156
rect 5411 3152 5412 3156
rect 5406 3151 5412 3152
rect 5542 3156 5548 3157
rect 5542 3152 5543 3156
rect 5547 3152 5548 3156
rect 5662 3153 5663 3157
rect 5667 3153 5668 3157
rect 5662 3152 5668 3153
rect 5542 3151 5548 3152
rect 2066 3141 2072 3142
rect 1974 3140 1980 3141
rect 1974 3136 1975 3140
rect 1979 3136 1980 3140
rect 2066 3137 2067 3141
rect 2071 3137 2072 3141
rect 2066 3136 2072 3137
rect 2266 3141 2272 3142
rect 2266 3137 2267 3141
rect 2271 3137 2272 3141
rect 2266 3136 2272 3137
rect 2458 3141 2464 3142
rect 2458 3137 2459 3141
rect 2463 3137 2464 3141
rect 2458 3136 2464 3137
rect 2650 3141 2656 3142
rect 2650 3137 2651 3141
rect 2655 3137 2656 3141
rect 2650 3136 2656 3137
rect 2842 3141 2848 3142
rect 2842 3137 2843 3141
rect 2847 3137 2848 3141
rect 2842 3136 2848 3137
rect 3026 3141 3032 3142
rect 3026 3137 3027 3141
rect 3031 3137 3032 3141
rect 3026 3136 3032 3137
rect 3202 3141 3208 3142
rect 3202 3137 3203 3141
rect 3207 3137 3208 3141
rect 3202 3136 3208 3137
rect 3386 3141 3392 3142
rect 3386 3137 3387 3141
rect 3391 3137 3392 3141
rect 3386 3136 3392 3137
rect 3570 3141 3576 3142
rect 4834 3141 4840 3142
rect 3570 3137 3571 3141
rect 3575 3137 3576 3141
rect 3570 3136 3576 3137
rect 3798 3140 3804 3141
rect 3798 3136 3799 3140
rect 3803 3136 3804 3140
rect 1974 3135 1980 3136
rect 3798 3135 3804 3136
rect 3838 3140 3844 3141
rect 3838 3136 3839 3140
rect 3843 3136 3844 3140
rect 4834 3137 4835 3141
rect 4839 3137 4840 3141
rect 4834 3136 4840 3137
rect 4970 3141 4976 3142
rect 4970 3137 4971 3141
rect 4975 3137 4976 3141
rect 4970 3136 4976 3137
rect 5106 3141 5112 3142
rect 5106 3137 5107 3141
rect 5111 3137 5112 3141
rect 5106 3136 5112 3137
rect 5242 3141 5248 3142
rect 5242 3137 5243 3141
rect 5247 3137 5248 3141
rect 5242 3136 5248 3137
rect 5378 3141 5384 3142
rect 5378 3137 5379 3141
rect 5383 3137 5384 3141
rect 5378 3136 5384 3137
rect 5514 3141 5520 3142
rect 5514 3137 5515 3141
rect 5519 3137 5520 3141
rect 5514 3136 5520 3137
rect 5662 3140 5668 3141
rect 5662 3136 5663 3140
rect 5667 3136 5668 3140
rect 3838 3135 3844 3136
rect 5662 3135 5668 3136
rect 110 3088 116 3089
rect 1934 3088 1940 3089
rect 110 3084 111 3088
rect 115 3084 116 3088
rect 110 3083 116 3084
rect 378 3087 384 3088
rect 378 3083 379 3087
rect 383 3083 384 3087
rect 378 3082 384 3083
rect 562 3087 568 3088
rect 562 3083 563 3087
rect 567 3083 568 3087
rect 562 3082 568 3083
rect 754 3087 760 3088
rect 754 3083 755 3087
rect 759 3083 760 3087
rect 754 3082 760 3083
rect 954 3087 960 3088
rect 954 3083 955 3087
rect 959 3083 960 3087
rect 954 3082 960 3083
rect 1162 3087 1168 3088
rect 1162 3083 1163 3087
rect 1167 3083 1168 3087
rect 1162 3082 1168 3083
rect 1370 3087 1376 3088
rect 1370 3083 1371 3087
rect 1375 3083 1376 3087
rect 1934 3084 1935 3088
rect 1939 3084 1940 3088
rect 1934 3083 1940 3084
rect 1370 3082 1376 3083
rect 406 3072 412 3073
rect 110 3071 116 3072
rect 110 3067 111 3071
rect 115 3067 116 3071
rect 406 3068 407 3072
rect 411 3068 412 3072
rect 406 3067 412 3068
rect 590 3072 596 3073
rect 590 3068 591 3072
rect 595 3068 596 3072
rect 590 3067 596 3068
rect 782 3072 788 3073
rect 782 3068 783 3072
rect 787 3068 788 3072
rect 782 3067 788 3068
rect 982 3072 988 3073
rect 982 3068 983 3072
rect 987 3068 988 3072
rect 982 3067 988 3068
rect 1190 3072 1196 3073
rect 1190 3068 1191 3072
rect 1195 3068 1196 3072
rect 1190 3067 1196 3068
rect 1398 3072 1404 3073
rect 1398 3068 1399 3072
rect 1403 3068 1404 3072
rect 1398 3067 1404 3068
rect 1934 3071 1940 3072
rect 1934 3067 1935 3071
rect 1939 3067 1940 3071
rect 110 3066 116 3067
rect 1934 3066 1940 3067
rect 110 2997 116 2998
rect 1934 2997 1940 2998
rect 110 2993 111 2997
rect 115 2993 116 2997
rect 110 2992 116 2993
rect 574 2996 580 2997
rect 574 2992 575 2996
rect 579 2992 580 2996
rect 574 2991 580 2992
rect 798 2996 804 2997
rect 798 2992 799 2996
rect 803 2992 804 2996
rect 798 2991 804 2992
rect 1046 2996 1052 2997
rect 1046 2992 1047 2996
rect 1051 2992 1052 2996
rect 1046 2991 1052 2992
rect 1302 2996 1308 2997
rect 1302 2992 1303 2996
rect 1307 2992 1308 2996
rect 1302 2991 1308 2992
rect 1566 2996 1572 2997
rect 1566 2992 1567 2996
rect 1571 2992 1572 2996
rect 1566 2991 1572 2992
rect 1814 2996 1820 2997
rect 1814 2992 1815 2996
rect 1819 2992 1820 2996
rect 1934 2993 1935 2997
rect 1939 2993 1940 2997
rect 1934 2992 1940 2993
rect 1974 2996 1980 2997
rect 3798 2996 3804 2997
rect 1974 2992 1975 2996
rect 1979 2992 1980 2996
rect 1814 2991 1820 2992
rect 1974 2991 1980 2992
rect 1994 2995 2000 2996
rect 1994 2991 1995 2995
rect 1999 2991 2000 2995
rect 1994 2990 2000 2991
rect 2130 2995 2136 2996
rect 2130 2991 2131 2995
rect 2135 2991 2136 2995
rect 2130 2990 2136 2991
rect 2266 2995 2272 2996
rect 2266 2991 2267 2995
rect 2271 2991 2272 2995
rect 2266 2990 2272 2991
rect 2402 2995 2408 2996
rect 2402 2991 2403 2995
rect 2407 2991 2408 2995
rect 2402 2990 2408 2991
rect 2538 2995 2544 2996
rect 2538 2991 2539 2995
rect 2543 2991 2544 2995
rect 2538 2990 2544 2991
rect 2682 2995 2688 2996
rect 2682 2991 2683 2995
rect 2687 2991 2688 2995
rect 2682 2990 2688 2991
rect 2834 2995 2840 2996
rect 2834 2991 2835 2995
rect 2839 2991 2840 2995
rect 2834 2990 2840 2991
rect 2986 2995 2992 2996
rect 2986 2991 2987 2995
rect 2991 2991 2992 2995
rect 2986 2990 2992 2991
rect 3138 2995 3144 2996
rect 3138 2991 3139 2995
rect 3143 2991 3144 2995
rect 3138 2990 3144 2991
rect 3290 2995 3296 2996
rect 3290 2991 3291 2995
rect 3295 2991 3296 2995
rect 3798 2992 3799 2996
rect 3803 2992 3804 2996
rect 3798 2991 3804 2992
rect 3838 2996 3844 2997
rect 5662 2996 5668 2997
rect 3838 2992 3839 2996
rect 3843 2992 3844 2996
rect 3838 2991 3844 2992
rect 4482 2995 4488 2996
rect 4482 2991 4483 2995
rect 4487 2991 4488 2995
rect 3290 2990 3296 2991
rect 4482 2990 4488 2991
rect 4634 2995 4640 2996
rect 4634 2991 4635 2995
rect 4639 2991 4640 2995
rect 4634 2990 4640 2991
rect 4802 2995 4808 2996
rect 4802 2991 4803 2995
rect 4807 2991 4808 2995
rect 4802 2990 4808 2991
rect 4978 2995 4984 2996
rect 4978 2991 4979 2995
rect 4983 2991 4984 2995
rect 4978 2990 4984 2991
rect 5162 2995 5168 2996
rect 5162 2991 5163 2995
rect 5167 2991 5168 2995
rect 5162 2990 5168 2991
rect 5346 2995 5352 2996
rect 5346 2991 5347 2995
rect 5351 2991 5352 2995
rect 5346 2990 5352 2991
rect 5514 2995 5520 2996
rect 5514 2991 5515 2995
rect 5519 2991 5520 2995
rect 5662 2992 5663 2996
rect 5667 2992 5668 2996
rect 5662 2991 5668 2992
rect 5514 2990 5520 2991
rect 546 2981 552 2982
rect 110 2980 116 2981
rect 110 2976 111 2980
rect 115 2976 116 2980
rect 546 2977 547 2981
rect 551 2977 552 2981
rect 546 2976 552 2977
rect 770 2981 776 2982
rect 770 2977 771 2981
rect 775 2977 776 2981
rect 770 2976 776 2977
rect 1018 2981 1024 2982
rect 1018 2977 1019 2981
rect 1023 2977 1024 2981
rect 1018 2976 1024 2977
rect 1274 2981 1280 2982
rect 1274 2977 1275 2981
rect 1279 2977 1280 2981
rect 1274 2976 1280 2977
rect 1538 2981 1544 2982
rect 1538 2977 1539 2981
rect 1543 2977 1544 2981
rect 1538 2976 1544 2977
rect 1786 2981 1792 2982
rect 1786 2977 1787 2981
rect 1791 2977 1792 2981
rect 1786 2976 1792 2977
rect 1934 2980 1940 2981
rect 2022 2980 2028 2981
rect 1934 2976 1935 2980
rect 1939 2976 1940 2980
rect 110 2975 116 2976
rect 1934 2975 1940 2976
rect 1974 2979 1980 2980
rect 1974 2975 1975 2979
rect 1979 2975 1980 2979
rect 2022 2976 2023 2980
rect 2027 2976 2028 2980
rect 2022 2975 2028 2976
rect 2158 2980 2164 2981
rect 2158 2976 2159 2980
rect 2163 2976 2164 2980
rect 2158 2975 2164 2976
rect 2294 2980 2300 2981
rect 2294 2976 2295 2980
rect 2299 2976 2300 2980
rect 2294 2975 2300 2976
rect 2430 2980 2436 2981
rect 2430 2976 2431 2980
rect 2435 2976 2436 2980
rect 2430 2975 2436 2976
rect 2566 2980 2572 2981
rect 2566 2976 2567 2980
rect 2571 2976 2572 2980
rect 2566 2975 2572 2976
rect 2710 2980 2716 2981
rect 2710 2976 2711 2980
rect 2715 2976 2716 2980
rect 2710 2975 2716 2976
rect 2862 2980 2868 2981
rect 2862 2976 2863 2980
rect 2867 2976 2868 2980
rect 2862 2975 2868 2976
rect 3014 2980 3020 2981
rect 3014 2976 3015 2980
rect 3019 2976 3020 2980
rect 3014 2975 3020 2976
rect 3166 2980 3172 2981
rect 3166 2976 3167 2980
rect 3171 2976 3172 2980
rect 3166 2975 3172 2976
rect 3318 2980 3324 2981
rect 4510 2980 4516 2981
rect 3318 2976 3319 2980
rect 3323 2976 3324 2980
rect 3318 2975 3324 2976
rect 3798 2979 3804 2980
rect 3798 2975 3799 2979
rect 3803 2975 3804 2979
rect 1974 2974 1980 2975
rect 3798 2974 3804 2975
rect 3838 2979 3844 2980
rect 3838 2975 3839 2979
rect 3843 2975 3844 2979
rect 4510 2976 4511 2980
rect 4515 2976 4516 2980
rect 4510 2975 4516 2976
rect 4662 2980 4668 2981
rect 4662 2976 4663 2980
rect 4667 2976 4668 2980
rect 4662 2975 4668 2976
rect 4830 2980 4836 2981
rect 4830 2976 4831 2980
rect 4835 2976 4836 2980
rect 4830 2975 4836 2976
rect 5006 2980 5012 2981
rect 5006 2976 5007 2980
rect 5011 2976 5012 2980
rect 5006 2975 5012 2976
rect 5190 2980 5196 2981
rect 5190 2976 5191 2980
rect 5195 2976 5196 2980
rect 5190 2975 5196 2976
rect 5374 2980 5380 2981
rect 5374 2976 5375 2980
rect 5379 2976 5380 2980
rect 5374 2975 5380 2976
rect 5542 2980 5548 2981
rect 5542 2976 5543 2980
rect 5547 2976 5548 2980
rect 5542 2975 5548 2976
rect 5662 2979 5668 2980
rect 5662 2975 5663 2979
rect 5667 2975 5668 2979
rect 3838 2974 3844 2975
rect 5662 2974 5668 2975
rect 1974 2921 1980 2922
rect 3798 2921 3804 2922
rect 1974 2917 1975 2921
rect 1979 2917 1980 2921
rect 1974 2916 1980 2917
rect 2022 2920 2028 2921
rect 2022 2916 2023 2920
rect 2027 2916 2028 2920
rect 2022 2915 2028 2916
rect 2294 2920 2300 2921
rect 2294 2916 2295 2920
rect 2299 2916 2300 2920
rect 2294 2915 2300 2916
rect 2590 2920 2596 2921
rect 2590 2916 2591 2920
rect 2595 2916 2596 2920
rect 2590 2915 2596 2916
rect 2886 2920 2892 2921
rect 2886 2916 2887 2920
rect 2891 2916 2892 2920
rect 2886 2915 2892 2916
rect 3182 2920 3188 2921
rect 3182 2916 3183 2920
rect 3187 2916 3188 2920
rect 3798 2917 3799 2921
rect 3803 2917 3804 2921
rect 3798 2916 3804 2917
rect 3182 2915 3188 2916
rect 1994 2905 2000 2906
rect 1974 2904 1980 2905
rect 1974 2900 1975 2904
rect 1979 2900 1980 2904
rect 1994 2901 1995 2905
rect 1999 2901 2000 2905
rect 1994 2900 2000 2901
rect 2266 2905 2272 2906
rect 2266 2901 2267 2905
rect 2271 2901 2272 2905
rect 2266 2900 2272 2901
rect 2562 2905 2568 2906
rect 2562 2901 2563 2905
rect 2567 2901 2568 2905
rect 2562 2900 2568 2901
rect 2858 2905 2864 2906
rect 2858 2901 2859 2905
rect 2863 2901 2864 2905
rect 2858 2900 2864 2901
rect 3154 2905 3160 2906
rect 3154 2901 3155 2905
rect 3159 2901 3160 2905
rect 3154 2900 3160 2901
rect 3798 2904 3804 2905
rect 3798 2900 3799 2904
rect 3803 2900 3804 2904
rect 1974 2899 1980 2900
rect 3798 2899 3804 2900
rect 3838 2897 3844 2898
rect 5662 2897 5668 2898
rect 3838 2893 3839 2897
rect 3843 2893 3844 2897
rect 3838 2892 3844 2893
rect 4046 2896 4052 2897
rect 4046 2892 4047 2896
rect 4051 2892 4052 2896
rect 4046 2891 4052 2892
rect 4294 2896 4300 2897
rect 4294 2892 4295 2896
rect 4299 2892 4300 2896
rect 4294 2891 4300 2892
rect 4582 2896 4588 2897
rect 4582 2892 4583 2896
rect 4587 2892 4588 2896
rect 4582 2891 4588 2892
rect 4894 2896 4900 2897
rect 4894 2892 4895 2896
rect 4899 2892 4900 2896
rect 4894 2891 4900 2892
rect 5230 2896 5236 2897
rect 5230 2892 5231 2896
rect 5235 2892 5236 2896
rect 5230 2891 5236 2892
rect 5542 2896 5548 2897
rect 5542 2892 5543 2896
rect 5547 2892 5548 2896
rect 5662 2893 5663 2897
rect 5667 2893 5668 2897
rect 5662 2892 5668 2893
rect 5542 2891 5548 2892
rect 4018 2881 4024 2882
rect 3838 2880 3844 2881
rect 3838 2876 3839 2880
rect 3843 2876 3844 2880
rect 4018 2877 4019 2881
rect 4023 2877 4024 2881
rect 4018 2876 4024 2877
rect 4266 2881 4272 2882
rect 4266 2877 4267 2881
rect 4271 2877 4272 2881
rect 4266 2876 4272 2877
rect 4554 2881 4560 2882
rect 4554 2877 4555 2881
rect 4559 2877 4560 2881
rect 4554 2876 4560 2877
rect 4866 2881 4872 2882
rect 4866 2877 4867 2881
rect 4871 2877 4872 2881
rect 4866 2876 4872 2877
rect 5202 2881 5208 2882
rect 5202 2877 5203 2881
rect 5207 2877 5208 2881
rect 5202 2876 5208 2877
rect 5514 2881 5520 2882
rect 5514 2877 5515 2881
rect 5519 2877 5520 2881
rect 5514 2876 5520 2877
rect 5662 2880 5668 2881
rect 5662 2876 5663 2880
rect 5667 2876 5668 2880
rect 3838 2875 3844 2876
rect 5662 2875 5668 2876
rect 110 2840 116 2841
rect 1934 2840 1940 2841
rect 110 2836 111 2840
rect 115 2836 116 2840
rect 110 2835 116 2836
rect 426 2839 432 2840
rect 426 2835 427 2839
rect 431 2835 432 2839
rect 426 2834 432 2835
rect 562 2839 568 2840
rect 562 2835 563 2839
rect 567 2835 568 2839
rect 562 2834 568 2835
rect 698 2839 704 2840
rect 698 2835 699 2839
rect 703 2835 704 2839
rect 698 2834 704 2835
rect 834 2839 840 2840
rect 834 2835 835 2839
rect 839 2835 840 2839
rect 834 2834 840 2835
rect 970 2839 976 2840
rect 970 2835 971 2839
rect 975 2835 976 2839
rect 970 2834 976 2835
rect 1106 2839 1112 2840
rect 1106 2835 1107 2839
rect 1111 2835 1112 2839
rect 1106 2834 1112 2835
rect 1242 2839 1248 2840
rect 1242 2835 1243 2839
rect 1247 2835 1248 2839
rect 1242 2834 1248 2835
rect 1378 2839 1384 2840
rect 1378 2835 1379 2839
rect 1383 2835 1384 2839
rect 1378 2834 1384 2835
rect 1514 2839 1520 2840
rect 1514 2835 1515 2839
rect 1519 2835 1520 2839
rect 1514 2834 1520 2835
rect 1650 2839 1656 2840
rect 1650 2835 1651 2839
rect 1655 2835 1656 2839
rect 1650 2834 1656 2835
rect 1786 2839 1792 2840
rect 1786 2835 1787 2839
rect 1791 2835 1792 2839
rect 1934 2836 1935 2840
rect 1939 2836 1940 2840
rect 1934 2835 1940 2836
rect 1786 2834 1792 2835
rect 454 2824 460 2825
rect 110 2823 116 2824
rect 110 2819 111 2823
rect 115 2819 116 2823
rect 454 2820 455 2824
rect 459 2820 460 2824
rect 454 2819 460 2820
rect 590 2824 596 2825
rect 590 2820 591 2824
rect 595 2820 596 2824
rect 590 2819 596 2820
rect 726 2824 732 2825
rect 726 2820 727 2824
rect 731 2820 732 2824
rect 726 2819 732 2820
rect 862 2824 868 2825
rect 862 2820 863 2824
rect 867 2820 868 2824
rect 862 2819 868 2820
rect 998 2824 1004 2825
rect 998 2820 999 2824
rect 1003 2820 1004 2824
rect 998 2819 1004 2820
rect 1134 2824 1140 2825
rect 1134 2820 1135 2824
rect 1139 2820 1140 2824
rect 1134 2819 1140 2820
rect 1270 2824 1276 2825
rect 1270 2820 1271 2824
rect 1275 2820 1276 2824
rect 1270 2819 1276 2820
rect 1406 2824 1412 2825
rect 1406 2820 1407 2824
rect 1411 2820 1412 2824
rect 1406 2819 1412 2820
rect 1542 2824 1548 2825
rect 1542 2820 1543 2824
rect 1547 2820 1548 2824
rect 1542 2819 1548 2820
rect 1678 2824 1684 2825
rect 1678 2820 1679 2824
rect 1683 2820 1684 2824
rect 1678 2819 1684 2820
rect 1814 2824 1820 2825
rect 1814 2820 1815 2824
rect 1819 2820 1820 2824
rect 1814 2819 1820 2820
rect 1934 2823 1940 2824
rect 1934 2819 1935 2823
rect 1939 2819 1940 2823
rect 110 2818 116 2819
rect 1934 2818 1940 2819
rect 110 2757 116 2758
rect 1934 2757 1940 2758
rect 110 2753 111 2757
rect 115 2753 116 2757
rect 110 2752 116 2753
rect 462 2756 468 2757
rect 462 2752 463 2756
rect 467 2752 468 2756
rect 462 2751 468 2752
rect 622 2756 628 2757
rect 622 2752 623 2756
rect 627 2752 628 2756
rect 622 2751 628 2752
rect 782 2756 788 2757
rect 782 2752 783 2756
rect 787 2752 788 2756
rect 782 2751 788 2752
rect 934 2756 940 2757
rect 934 2752 935 2756
rect 939 2752 940 2756
rect 934 2751 940 2752
rect 1086 2756 1092 2757
rect 1086 2752 1087 2756
rect 1091 2752 1092 2756
rect 1086 2751 1092 2752
rect 1238 2756 1244 2757
rect 1238 2752 1239 2756
rect 1243 2752 1244 2756
rect 1238 2751 1244 2752
rect 1382 2756 1388 2757
rect 1382 2752 1383 2756
rect 1387 2752 1388 2756
rect 1382 2751 1388 2752
rect 1534 2756 1540 2757
rect 1534 2752 1535 2756
rect 1539 2752 1540 2756
rect 1534 2751 1540 2752
rect 1678 2756 1684 2757
rect 1678 2752 1679 2756
rect 1683 2752 1684 2756
rect 1678 2751 1684 2752
rect 1814 2756 1820 2757
rect 1814 2752 1815 2756
rect 1819 2752 1820 2756
rect 1934 2753 1935 2757
rect 1939 2753 1940 2757
rect 1934 2752 1940 2753
rect 1814 2751 1820 2752
rect 3838 2744 3844 2745
rect 5662 2744 5668 2745
rect 434 2741 440 2742
rect 110 2740 116 2741
rect 110 2736 111 2740
rect 115 2736 116 2740
rect 434 2737 435 2741
rect 439 2737 440 2741
rect 434 2736 440 2737
rect 594 2741 600 2742
rect 594 2737 595 2741
rect 599 2737 600 2741
rect 594 2736 600 2737
rect 754 2741 760 2742
rect 754 2737 755 2741
rect 759 2737 760 2741
rect 754 2736 760 2737
rect 906 2741 912 2742
rect 906 2737 907 2741
rect 911 2737 912 2741
rect 906 2736 912 2737
rect 1058 2741 1064 2742
rect 1058 2737 1059 2741
rect 1063 2737 1064 2741
rect 1058 2736 1064 2737
rect 1210 2741 1216 2742
rect 1210 2737 1211 2741
rect 1215 2737 1216 2741
rect 1210 2736 1216 2737
rect 1354 2741 1360 2742
rect 1354 2737 1355 2741
rect 1359 2737 1360 2741
rect 1354 2736 1360 2737
rect 1506 2741 1512 2742
rect 1506 2737 1507 2741
rect 1511 2737 1512 2741
rect 1506 2736 1512 2737
rect 1650 2741 1656 2742
rect 1650 2737 1651 2741
rect 1655 2737 1656 2741
rect 1650 2736 1656 2737
rect 1786 2741 1792 2742
rect 1786 2737 1787 2741
rect 1791 2737 1792 2741
rect 1786 2736 1792 2737
rect 1934 2740 1940 2741
rect 1934 2736 1935 2740
rect 1939 2736 1940 2740
rect 3838 2740 3839 2744
rect 3843 2740 3844 2744
rect 3838 2739 3844 2740
rect 3858 2743 3864 2744
rect 3858 2739 3859 2743
rect 3863 2739 3864 2743
rect 3858 2738 3864 2739
rect 3994 2743 4000 2744
rect 3994 2739 3995 2743
rect 3999 2739 4000 2743
rect 3994 2738 4000 2739
rect 4130 2743 4136 2744
rect 4130 2739 4131 2743
rect 4135 2739 4136 2743
rect 4130 2738 4136 2739
rect 4266 2743 4272 2744
rect 4266 2739 4267 2743
rect 4271 2739 4272 2743
rect 4266 2738 4272 2739
rect 4402 2743 4408 2744
rect 4402 2739 4403 2743
rect 4407 2739 4408 2743
rect 4402 2738 4408 2739
rect 4538 2743 4544 2744
rect 4538 2739 4539 2743
rect 4543 2739 4544 2743
rect 4538 2738 4544 2739
rect 4674 2743 4680 2744
rect 4674 2739 4675 2743
rect 4679 2739 4680 2743
rect 4674 2738 4680 2739
rect 4810 2743 4816 2744
rect 4810 2739 4811 2743
rect 4815 2739 4816 2743
rect 5662 2740 5663 2744
rect 5667 2740 5668 2744
rect 5662 2739 5668 2740
rect 4810 2738 4816 2739
rect 110 2735 116 2736
rect 1934 2735 1940 2736
rect 3886 2728 3892 2729
rect 3838 2727 3844 2728
rect 3838 2723 3839 2727
rect 3843 2723 3844 2727
rect 3886 2724 3887 2728
rect 3891 2724 3892 2728
rect 3886 2723 3892 2724
rect 4022 2728 4028 2729
rect 4022 2724 4023 2728
rect 4027 2724 4028 2728
rect 4022 2723 4028 2724
rect 4158 2728 4164 2729
rect 4158 2724 4159 2728
rect 4163 2724 4164 2728
rect 4158 2723 4164 2724
rect 4294 2728 4300 2729
rect 4294 2724 4295 2728
rect 4299 2724 4300 2728
rect 4294 2723 4300 2724
rect 4430 2728 4436 2729
rect 4430 2724 4431 2728
rect 4435 2724 4436 2728
rect 4430 2723 4436 2724
rect 4566 2728 4572 2729
rect 4566 2724 4567 2728
rect 4571 2724 4572 2728
rect 4566 2723 4572 2724
rect 4702 2728 4708 2729
rect 4702 2724 4703 2728
rect 4707 2724 4708 2728
rect 4702 2723 4708 2724
rect 4838 2728 4844 2729
rect 4838 2724 4839 2728
rect 4843 2724 4844 2728
rect 4838 2723 4844 2724
rect 5662 2727 5668 2728
rect 5662 2723 5663 2727
rect 5667 2723 5668 2727
rect 3838 2722 3844 2723
rect 5662 2722 5668 2723
rect 1974 2716 1980 2717
rect 3798 2716 3804 2717
rect 1974 2712 1975 2716
rect 1979 2712 1980 2716
rect 1974 2711 1980 2712
rect 3058 2715 3064 2716
rect 3058 2711 3059 2715
rect 3063 2711 3064 2715
rect 3058 2710 3064 2711
rect 3194 2715 3200 2716
rect 3194 2711 3195 2715
rect 3199 2711 3200 2715
rect 3194 2710 3200 2711
rect 3330 2715 3336 2716
rect 3330 2711 3331 2715
rect 3335 2711 3336 2715
rect 3798 2712 3799 2716
rect 3803 2712 3804 2716
rect 3798 2711 3804 2712
rect 3330 2710 3336 2711
rect 3086 2700 3092 2701
rect 1974 2699 1980 2700
rect 1974 2695 1975 2699
rect 1979 2695 1980 2699
rect 3086 2696 3087 2700
rect 3091 2696 3092 2700
rect 3086 2695 3092 2696
rect 3222 2700 3228 2701
rect 3222 2696 3223 2700
rect 3227 2696 3228 2700
rect 3222 2695 3228 2696
rect 3358 2700 3364 2701
rect 3358 2696 3359 2700
rect 3363 2696 3364 2700
rect 3358 2695 3364 2696
rect 3798 2699 3804 2700
rect 3798 2695 3799 2699
rect 3803 2695 3804 2699
rect 1974 2694 1980 2695
rect 3798 2694 3804 2695
rect 3838 2669 3844 2670
rect 5662 2669 5668 2670
rect 3838 2665 3839 2669
rect 3843 2665 3844 2669
rect 3838 2664 3844 2665
rect 4054 2668 4060 2669
rect 4054 2664 4055 2668
rect 4059 2664 4060 2668
rect 4054 2663 4060 2664
rect 4302 2668 4308 2669
rect 4302 2664 4303 2668
rect 4307 2664 4308 2668
rect 4302 2663 4308 2664
rect 4582 2668 4588 2669
rect 4582 2664 4583 2668
rect 4587 2664 4588 2668
rect 4582 2663 4588 2664
rect 4894 2668 4900 2669
rect 4894 2664 4895 2668
rect 4899 2664 4900 2668
rect 4894 2663 4900 2664
rect 5230 2668 5236 2669
rect 5230 2664 5231 2668
rect 5235 2664 5236 2668
rect 5230 2663 5236 2664
rect 5542 2668 5548 2669
rect 5542 2664 5543 2668
rect 5547 2664 5548 2668
rect 5662 2665 5663 2669
rect 5667 2665 5668 2669
rect 5662 2664 5668 2665
rect 5542 2663 5548 2664
rect 4026 2653 4032 2654
rect 3838 2652 3844 2653
rect 3838 2648 3839 2652
rect 3843 2648 3844 2652
rect 4026 2649 4027 2653
rect 4031 2649 4032 2653
rect 4026 2648 4032 2649
rect 4274 2653 4280 2654
rect 4274 2649 4275 2653
rect 4279 2649 4280 2653
rect 4274 2648 4280 2649
rect 4554 2653 4560 2654
rect 4554 2649 4555 2653
rect 4559 2649 4560 2653
rect 4554 2648 4560 2649
rect 4866 2653 4872 2654
rect 4866 2649 4867 2653
rect 4871 2649 4872 2653
rect 4866 2648 4872 2649
rect 5202 2653 5208 2654
rect 5202 2649 5203 2653
rect 5207 2649 5208 2653
rect 5202 2648 5208 2649
rect 5514 2653 5520 2654
rect 5514 2649 5515 2653
rect 5519 2649 5520 2653
rect 5514 2648 5520 2649
rect 5662 2652 5668 2653
rect 5662 2648 5663 2652
rect 5667 2648 5668 2652
rect 3838 2647 3844 2648
rect 5662 2647 5668 2648
rect 1974 2617 1980 2618
rect 3798 2617 3804 2618
rect 1974 2613 1975 2617
rect 1979 2613 1980 2617
rect 1974 2612 1980 2613
rect 3134 2616 3140 2617
rect 3134 2612 3135 2616
rect 3139 2612 3140 2616
rect 3134 2611 3140 2612
rect 3270 2616 3276 2617
rect 3270 2612 3271 2616
rect 3275 2612 3276 2616
rect 3270 2611 3276 2612
rect 3406 2616 3412 2617
rect 3406 2612 3407 2616
rect 3411 2612 3412 2616
rect 3406 2611 3412 2612
rect 3542 2616 3548 2617
rect 3542 2612 3543 2616
rect 3547 2612 3548 2616
rect 3542 2611 3548 2612
rect 3678 2616 3684 2617
rect 3678 2612 3679 2616
rect 3683 2612 3684 2616
rect 3798 2613 3799 2617
rect 3803 2613 3804 2617
rect 3798 2612 3804 2613
rect 3678 2611 3684 2612
rect 110 2604 116 2605
rect 1934 2604 1940 2605
rect 110 2600 111 2604
rect 115 2600 116 2604
rect 110 2599 116 2600
rect 354 2603 360 2604
rect 354 2599 355 2603
rect 359 2599 360 2603
rect 354 2598 360 2599
rect 538 2603 544 2604
rect 538 2599 539 2603
rect 543 2599 544 2603
rect 538 2598 544 2599
rect 714 2603 720 2604
rect 714 2599 715 2603
rect 719 2599 720 2603
rect 714 2598 720 2599
rect 882 2603 888 2604
rect 882 2599 883 2603
rect 887 2599 888 2603
rect 882 2598 888 2599
rect 1042 2603 1048 2604
rect 1042 2599 1043 2603
rect 1047 2599 1048 2603
rect 1042 2598 1048 2599
rect 1202 2603 1208 2604
rect 1202 2599 1203 2603
rect 1207 2599 1208 2603
rect 1202 2598 1208 2599
rect 1354 2603 1360 2604
rect 1354 2599 1355 2603
rect 1359 2599 1360 2603
rect 1354 2598 1360 2599
rect 1506 2603 1512 2604
rect 1506 2599 1507 2603
rect 1511 2599 1512 2603
rect 1506 2598 1512 2599
rect 1650 2603 1656 2604
rect 1650 2599 1651 2603
rect 1655 2599 1656 2603
rect 1650 2598 1656 2599
rect 1786 2603 1792 2604
rect 1786 2599 1787 2603
rect 1791 2599 1792 2603
rect 1934 2600 1935 2604
rect 1939 2600 1940 2604
rect 3106 2601 3112 2602
rect 1934 2599 1940 2600
rect 1974 2600 1980 2601
rect 1786 2598 1792 2599
rect 1974 2596 1975 2600
rect 1979 2596 1980 2600
rect 3106 2597 3107 2601
rect 3111 2597 3112 2601
rect 3106 2596 3112 2597
rect 3242 2601 3248 2602
rect 3242 2597 3243 2601
rect 3247 2597 3248 2601
rect 3242 2596 3248 2597
rect 3378 2601 3384 2602
rect 3378 2597 3379 2601
rect 3383 2597 3384 2601
rect 3378 2596 3384 2597
rect 3514 2601 3520 2602
rect 3514 2597 3515 2601
rect 3519 2597 3520 2601
rect 3514 2596 3520 2597
rect 3650 2601 3656 2602
rect 3650 2597 3651 2601
rect 3655 2597 3656 2601
rect 3650 2596 3656 2597
rect 3798 2600 3804 2601
rect 3798 2596 3799 2600
rect 3803 2596 3804 2600
rect 1974 2595 1980 2596
rect 3798 2595 3804 2596
rect 382 2588 388 2589
rect 110 2587 116 2588
rect 110 2583 111 2587
rect 115 2583 116 2587
rect 382 2584 383 2588
rect 387 2584 388 2588
rect 382 2583 388 2584
rect 566 2588 572 2589
rect 566 2584 567 2588
rect 571 2584 572 2588
rect 566 2583 572 2584
rect 742 2588 748 2589
rect 742 2584 743 2588
rect 747 2584 748 2588
rect 742 2583 748 2584
rect 910 2588 916 2589
rect 910 2584 911 2588
rect 915 2584 916 2588
rect 910 2583 916 2584
rect 1070 2588 1076 2589
rect 1070 2584 1071 2588
rect 1075 2584 1076 2588
rect 1070 2583 1076 2584
rect 1230 2588 1236 2589
rect 1230 2584 1231 2588
rect 1235 2584 1236 2588
rect 1230 2583 1236 2584
rect 1382 2588 1388 2589
rect 1382 2584 1383 2588
rect 1387 2584 1388 2588
rect 1382 2583 1388 2584
rect 1534 2588 1540 2589
rect 1534 2584 1535 2588
rect 1539 2584 1540 2588
rect 1534 2583 1540 2584
rect 1678 2588 1684 2589
rect 1678 2584 1679 2588
rect 1683 2584 1684 2588
rect 1678 2583 1684 2584
rect 1814 2588 1820 2589
rect 1814 2584 1815 2588
rect 1819 2584 1820 2588
rect 1814 2583 1820 2584
rect 1934 2587 1940 2588
rect 1934 2583 1935 2587
rect 1939 2583 1940 2587
rect 110 2582 116 2583
rect 1934 2582 1940 2583
rect 110 2529 116 2530
rect 1934 2529 1940 2530
rect 110 2525 111 2529
rect 115 2525 116 2529
rect 110 2524 116 2525
rect 230 2528 236 2529
rect 230 2524 231 2528
rect 235 2524 236 2528
rect 230 2523 236 2524
rect 422 2528 428 2529
rect 422 2524 423 2528
rect 427 2524 428 2528
rect 422 2523 428 2524
rect 622 2528 628 2529
rect 622 2524 623 2528
rect 627 2524 628 2528
rect 622 2523 628 2524
rect 822 2528 828 2529
rect 822 2524 823 2528
rect 827 2524 828 2528
rect 822 2523 828 2524
rect 1022 2528 1028 2529
rect 1022 2524 1023 2528
rect 1027 2524 1028 2528
rect 1022 2523 1028 2524
rect 1222 2528 1228 2529
rect 1222 2524 1223 2528
rect 1227 2524 1228 2528
rect 1222 2523 1228 2524
rect 1422 2528 1428 2529
rect 1422 2524 1423 2528
rect 1427 2524 1428 2528
rect 1422 2523 1428 2524
rect 1630 2528 1636 2529
rect 1630 2524 1631 2528
rect 1635 2524 1636 2528
rect 1630 2523 1636 2524
rect 1814 2528 1820 2529
rect 1814 2524 1815 2528
rect 1819 2524 1820 2528
rect 1934 2525 1935 2529
rect 1939 2525 1940 2529
rect 1934 2524 1940 2525
rect 1814 2523 1820 2524
rect 3838 2516 3844 2517
rect 5662 2516 5668 2517
rect 202 2513 208 2514
rect 110 2512 116 2513
rect 110 2508 111 2512
rect 115 2508 116 2512
rect 202 2509 203 2513
rect 207 2509 208 2513
rect 202 2508 208 2509
rect 394 2513 400 2514
rect 394 2509 395 2513
rect 399 2509 400 2513
rect 394 2508 400 2509
rect 594 2513 600 2514
rect 594 2509 595 2513
rect 599 2509 600 2513
rect 594 2508 600 2509
rect 794 2513 800 2514
rect 794 2509 795 2513
rect 799 2509 800 2513
rect 794 2508 800 2509
rect 994 2513 1000 2514
rect 994 2509 995 2513
rect 999 2509 1000 2513
rect 994 2508 1000 2509
rect 1194 2513 1200 2514
rect 1194 2509 1195 2513
rect 1199 2509 1200 2513
rect 1194 2508 1200 2509
rect 1394 2513 1400 2514
rect 1394 2509 1395 2513
rect 1399 2509 1400 2513
rect 1394 2508 1400 2509
rect 1602 2513 1608 2514
rect 1602 2509 1603 2513
rect 1607 2509 1608 2513
rect 1602 2508 1608 2509
rect 1786 2513 1792 2514
rect 1786 2509 1787 2513
rect 1791 2509 1792 2513
rect 1786 2508 1792 2509
rect 1934 2512 1940 2513
rect 1934 2508 1935 2512
rect 1939 2508 1940 2512
rect 3838 2512 3839 2516
rect 3843 2512 3844 2516
rect 3838 2511 3844 2512
rect 4258 2515 4264 2516
rect 4258 2511 4259 2515
rect 4263 2511 4264 2515
rect 4258 2510 4264 2511
rect 4474 2515 4480 2516
rect 4474 2511 4475 2515
rect 4479 2511 4480 2515
rect 4474 2510 4480 2511
rect 4714 2515 4720 2516
rect 4714 2511 4715 2515
rect 4719 2511 4720 2515
rect 4714 2510 4720 2511
rect 4978 2515 4984 2516
rect 4978 2511 4979 2515
rect 4983 2511 4984 2515
rect 4978 2510 4984 2511
rect 5258 2515 5264 2516
rect 5258 2511 5259 2515
rect 5263 2511 5264 2515
rect 5258 2510 5264 2511
rect 5514 2515 5520 2516
rect 5514 2511 5515 2515
rect 5519 2511 5520 2515
rect 5662 2512 5663 2516
rect 5667 2512 5668 2516
rect 5662 2511 5668 2512
rect 5514 2510 5520 2511
rect 110 2507 116 2508
rect 1934 2507 1940 2508
rect 4286 2500 4292 2501
rect 3838 2499 3844 2500
rect 3838 2495 3839 2499
rect 3843 2495 3844 2499
rect 4286 2496 4287 2500
rect 4291 2496 4292 2500
rect 4286 2495 4292 2496
rect 4502 2500 4508 2501
rect 4502 2496 4503 2500
rect 4507 2496 4508 2500
rect 4502 2495 4508 2496
rect 4742 2500 4748 2501
rect 4742 2496 4743 2500
rect 4747 2496 4748 2500
rect 4742 2495 4748 2496
rect 5006 2500 5012 2501
rect 5006 2496 5007 2500
rect 5011 2496 5012 2500
rect 5006 2495 5012 2496
rect 5286 2500 5292 2501
rect 5286 2496 5287 2500
rect 5291 2496 5292 2500
rect 5286 2495 5292 2496
rect 5542 2500 5548 2501
rect 5542 2496 5543 2500
rect 5547 2496 5548 2500
rect 5542 2495 5548 2496
rect 5662 2499 5668 2500
rect 5662 2495 5663 2499
rect 5667 2495 5668 2499
rect 3838 2494 3844 2495
rect 5662 2494 5668 2495
rect 1974 2460 1980 2461
rect 3798 2460 3804 2461
rect 1974 2456 1975 2460
rect 1979 2456 1980 2460
rect 1974 2455 1980 2456
rect 1994 2459 2000 2460
rect 1994 2455 1995 2459
rect 1999 2455 2000 2459
rect 1994 2454 2000 2455
rect 2234 2459 2240 2460
rect 2234 2455 2235 2459
rect 2239 2455 2240 2459
rect 2234 2454 2240 2455
rect 2482 2459 2488 2460
rect 2482 2455 2483 2459
rect 2487 2455 2488 2459
rect 2482 2454 2488 2455
rect 2714 2459 2720 2460
rect 2714 2455 2715 2459
rect 2719 2455 2720 2459
rect 2714 2454 2720 2455
rect 2938 2459 2944 2460
rect 2938 2455 2939 2459
rect 2943 2455 2944 2459
rect 2938 2454 2944 2455
rect 3154 2459 3160 2460
rect 3154 2455 3155 2459
rect 3159 2455 3160 2459
rect 3154 2454 3160 2455
rect 3362 2459 3368 2460
rect 3362 2455 3363 2459
rect 3367 2455 3368 2459
rect 3362 2454 3368 2455
rect 3578 2459 3584 2460
rect 3578 2455 3579 2459
rect 3583 2455 3584 2459
rect 3798 2456 3799 2460
rect 3803 2456 3804 2460
rect 3798 2455 3804 2456
rect 3578 2454 3584 2455
rect 2022 2444 2028 2445
rect 1974 2443 1980 2444
rect 1974 2439 1975 2443
rect 1979 2439 1980 2443
rect 2022 2440 2023 2444
rect 2027 2440 2028 2444
rect 2022 2439 2028 2440
rect 2262 2444 2268 2445
rect 2262 2440 2263 2444
rect 2267 2440 2268 2444
rect 2262 2439 2268 2440
rect 2510 2444 2516 2445
rect 2510 2440 2511 2444
rect 2515 2440 2516 2444
rect 2510 2439 2516 2440
rect 2742 2444 2748 2445
rect 2742 2440 2743 2444
rect 2747 2440 2748 2444
rect 2742 2439 2748 2440
rect 2966 2444 2972 2445
rect 2966 2440 2967 2444
rect 2971 2440 2972 2444
rect 2966 2439 2972 2440
rect 3182 2444 3188 2445
rect 3182 2440 3183 2444
rect 3187 2440 3188 2444
rect 3182 2439 3188 2440
rect 3390 2444 3396 2445
rect 3390 2440 3391 2444
rect 3395 2440 3396 2444
rect 3390 2439 3396 2440
rect 3606 2444 3612 2445
rect 3606 2440 3607 2444
rect 3611 2440 3612 2444
rect 3606 2439 3612 2440
rect 3798 2443 3804 2444
rect 3798 2439 3799 2443
rect 3803 2439 3804 2443
rect 1974 2438 1980 2439
rect 3798 2438 3804 2439
rect 3838 2437 3844 2438
rect 5662 2437 5668 2438
rect 3838 2433 3839 2437
rect 3843 2433 3844 2437
rect 3838 2432 3844 2433
rect 4662 2436 4668 2437
rect 4662 2432 4663 2436
rect 4667 2432 4668 2436
rect 4662 2431 4668 2432
rect 4846 2436 4852 2437
rect 4846 2432 4847 2436
rect 4851 2432 4852 2436
rect 4846 2431 4852 2432
rect 5022 2436 5028 2437
rect 5022 2432 5023 2436
rect 5027 2432 5028 2436
rect 5022 2431 5028 2432
rect 5198 2436 5204 2437
rect 5198 2432 5199 2436
rect 5203 2432 5204 2436
rect 5198 2431 5204 2432
rect 5382 2436 5388 2437
rect 5382 2432 5383 2436
rect 5387 2432 5388 2436
rect 5382 2431 5388 2432
rect 5542 2436 5548 2437
rect 5542 2432 5543 2436
rect 5547 2432 5548 2436
rect 5662 2433 5663 2437
rect 5667 2433 5668 2437
rect 5662 2432 5668 2433
rect 5542 2431 5548 2432
rect 4634 2421 4640 2422
rect 3838 2420 3844 2421
rect 3838 2416 3839 2420
rect 3843 2416 3844 2420
rect 4634 2417 4635 2421
rect 4639 2417 4640 2421
rect 4634 2416 4640 2417
rect 4818 2421 4824 2422
rect 4818 2417 4819 2421
rect 4823 2417 4824 2421
rect 4818 2416 4824 2417
rect 4994 2421 5000 2422
rect 4994 2417 4995 2421
rect 4999 2417 5000 2421
rect 4994 2416 5000 2417
rect 5170 2421 5176 2422
rect 5170 2417 5171 2421
rect 5175 2417 5176 2421
rect 5170 2416 5176 2417
rect 5354 2421 5360 2422
rect 5354 2417 5355 2421
rect 5359 2417 5360 2421
rect 5354 2416 5360 2417
rect 5514 2421 5520 2422
rect 5514 2417 5515 2421
rect 5519 2417 5520 2421
rect 5514 2416 5520 2417
rect 5662 2420 5668 2421
rect 5662 2416 5663 2420
rect 5667 2416 5668 2420
rect 3838 2415 3844 2416
rect 5662 2415 5668 2416
rect 1974 2385 1980 2386
rect 3798 2385 3804 2386
rect 1974 2381 1975 2385
rect 1979 2381 1980 2385
rect 1974 2380 1980 2381
rect 2022 2384 2028 2385
rect 2022 2380 2023 2384
rect 2027 2380 2028 2384
rect 2022 2379 2028 2380
rect 2158 2384 2164 2385
rect 2158 2380 2159 2384
rect 2163 2380 2164 2384
rect 2158 2379 2164 2380
rect 2294 2384 2300 2385
rect 2294 2380 2295 2384
rect 2299 2380 2300 2384
rect 2294 2379 2300 2380
rect 2430 2384 2436 2385
rect 2430 2380 2431 2384
rect 2435 2380 2436 2384
rect 2430 2379 2436 2380
rect 2566 2384 2572 2385
rect 2566 2380 2567 2384
rect 2571 2380 2572 2384
rect 2566 2379 2572 2380
rect 2710 2384 2716 2385
rect 2710 2380 2711 2384
rect 2715 2380 2716 2384
rect 2710 2379 2716 2380
rect 2854 2384 2860 2385
rect 2854 2380 2855 2384
rect 2859 2380 2860 2384
rect 2854 2379 2860 2380
rect 3006 2384 3012 2385
rect 3006 2380 3007 2384
rect 3011 2380 3012 2384
rect 3006 2379 3012 2380
rect 3158 2384 3164 2385
rect 3158 2380 3159 2384
rect 3163 2380 3164 2384
rect 3158 2379 3164 2380
rect 3310 2384 3316 2385
rect 3310 2380 3311 2384
rect 3315 2380 3316 2384
rect 3798 2381 3799 2385
rect 3803 2381 3804 2385
rect 3798 2380 3804 2381
rect 3310 2379 3316 2380
rect 1994 2369 2000 2370
rect 1974 2368 1980 2369
rect 1974 2364 1975 2368
rect 1979 2364 1980 2368
rect 1994 2365 1995 2369
rect 1999 2365 2000 2369
rect 1994 2364 2000 2365
rect 2130 2369 2136 2370
rect 2130 2365 2131 2369
rect 2135 2365 2136 2369
rect 2130 2364 2136 2365
rect 2266 2369 2272 2370
rect 2266 2365 2267 2369
rect 2271 2365 2272 2369
rect 2266 2364 2272 2365
rect 2402 2369 2408 2370
rect 2402 2365 2403 2369
rect 2407 2365 2408 2369
rect 2402 2364 2408 2365
rect 2538 2369 2544 2370
rect 2538 2365 2539 2369
rect 2543 2365 2544 2369
rect 2538 2364 2544 2365
rect 2682 2369 2688 2370
rect 2682 2365 2683 2369
rect 2687 2365 2688 2369
rect 2682 2364 2688 2365
rect 2826 2369 2832 2370
rect 2826 2365 2827 2369
rect 2831 2365 2832 2369
rect 2826 2364 2832 2365
rect 2978 2369 2984 2370
rect 2978 2365 2979 2369
rect 2983 2365 2984 2369
rect 2978 2364 2984 2365
rect 3130 2369 3136 2370
rect 3130 2365 3131 2369
rect 3135 2365 3136 2369
rect 3130 2364 3136 2365
rect 3282 2369 3288 2370
rect 3282 2365 3283 2369
rect 3287 2365 3288 2369
rect 3282 2364 3288 2365
rect 3798 2368 3804 2369
rect 3798 2364 3799 2368
rect 3803 2364 3804 2368
rect 1974 2363 1980 2364
rect 3798 2363 3804 2364
rect 110 2360 116 2361
rect 1934 2360 1940 2361
rect 110 2356 111 2360
rect 115 2356 116 2360
rect 110 2355 116 2356
rect 218 2359 224 2360
rect 218 2355 219 2359
rect 223 2355 224 2359
rect 218 2354 224 2355
rect 402 2359 408 2360
rect 402 2355 403 2359
rect 407 2355 408 2359
rect 402 2354 408 2355
rect 594 2359 600 2360
rect 594 2355 595 2359
rect 599 2355 600 2359
rect 594 2354 600 2355
rect 786 2359 792 2360
rect 786 2355 787 2359
rect 791 2355 792 2359
rect 786 2354 792 2355
rect 978 2359 984 2360
rect 978 2355 979 2359
rect 983 2355 984 2359
rect 1934 2356 1935 2360
rect 1939 2356 1940 2360
rect 1934 2355 1940 2356
rect 978 2354 984 2355
rect 246 2344 252 2345
rect 110 2343 116 2344
rect 110 2339 111 2343
rect 115 2339 116 2343
rect 246 2340 247 2344
rect 251 2340 252 2344
rect 246 2339 252 2340
rect 430 2344 436 2345
rect 430 2340 431 2344
rect 435 2340 436 2344
rect 430 2339 436 2340
rect 622 2344 628 2345
rect 622 2340 623 2344
rect 627 2340 628 2344
rect 622 2339 628 2340
rect 814 2344 820 2345
rect 814 2340 815 2344
rect 819 2340 820 2344
rect 814 2339 820 2340
rect 1006 2344 1012 2345
rect 1006 2340 1007 2344
rect 1011 2340 1012 2344
rect 1006 2339 1012 2340
rect 1934 2343 1940 2344
rect 1934 2339 1935 2343
rect 1939 2339 1940 2343
rect 110 2338 116 2339
rect 1934 2338 1940 2339
rect 3838 2284 3844 2285
rect 5662 2284 5668 2285
rect 110 2281 116 2282
rect 1934 2281 1940 2282
rect 110 2277 111 2281
rect 115 2277 116 2281
rect 110 2276 116 2277
rect 398 2280 404 2281
rect 398 2276 399 2280
rect 403 2276 404 2280
rect 398 2275 404 2276
rect 534 2280 540 2281
rect 534 2276 535 2280
rect 539 2276 540 2280
rect 534 2275 540 2276
rect 670 2280 676 2281
rect 670 2276 671 2280
rect 675 2276 676 2280
rect 670 2275 676 2276
rect 806 2280 812 2281
rect 806 2276 807 2280
rect 811 2276 812 2280
rect 806 2275 812 2276
rect 942 2280 948 2281
rect 942 2276 943 2280
rect 947 2276 948 2280
rect 1934 2277 1935 2281
rect 1939 2277 1940 2281
rect 3838 2280 3839 2284
rect 3843 2280 3844 2284
rect 3838 2279 3844 2280
rect 4674 2283 4680 2284
rect 4674 2279 4675 2283
rect 4679 2279 4680 2283
rect 4674 2278 4680 2279
rect 4818 2283 4824 2284
rect 4818 2279 4819 2283
rect 4823 2279 4824 2283
rect 4818 2278 4824 2279
rect 4962 2283 4968 2284
rect 4962 2279 4963 2283
rect 4967 2279 4968 2283
rect 4962 2278 4968 2279
rect 5114 2283 5120 2284
rect 5114 2279 5115 2283
rect 5119 2279 5120 2283
rect 5114 2278 5120 2279
rect 5266 2283 5272 2284
rect 5266 2279 5267 2283
rect 5271 2279 5272 2283
rect 5266 2278 5272 2279
rect 5418 2283 5424 2284
rect 5418 2279 5419 2283
rect 5423 2279 5424 2283
rect 5662 2280 5663 2284
rect 5667 2280 5668 2284
rect 5662 2279 5668 2280
rect 5418 2278 5424 2279
rect 1934 2276 1940 2277
rect 942 2275 948 2276
rect 4702 2268 4708 2269
rect 3838 2267 3844 2268
rect 370 2265 376 2266
rect 110 2264 116 2265
rect 110 2260 111 2264
rect 115 2260 116 2264
rect 370 2261 371 2265
rect 375 2261 376 2265
rect 370 2260 376 2261
rect 506 2265 512 2266
rect 506 2261 507 2265
rect 511 2261 512 2265
rect 506 2260 512 2261
rect 642 2265 648 2266
rect 642 2261 643 2265
rect 647 2261 648 2265
rect 642 2260 648 2261
rect 778 2265 784 2266
rect 778 2261 779 2265
rect 783 2261 784 2265
rect 778 2260 784 2261
rect 914 2265 920 2266
rect 914 2261 915 2265
rect 919 2261 920 2265
rect 914 2260 920 2261
rect 1934 2264 1940 2265
rect 1934 2260 1935 2264
rect 1939 2260 1940 2264
rect 3838 2263 3839 2267
rect 3843 2263 3844 2267
rect 4702 2264 4703 2268
rect 4707 2264 4708 2268
rect 4702 2263 4708 2264
rect 4846 2268 4852 2269
rect 4846 2264 4847 2268
rect 4851 2264 4852 2268
rect 4846 2263 4852 2264
rect 4990 2268 4996 2269
rect 4990 2264 4991 2268
rect 4995 2264 4996 2268
rect 4990 2263 4996 2264
rect 5142 2268 5148 2269
rect 5142 2264 5143 2268
rect 5147 2264 5148 2268
rect 5142 2263 5148 2264
rect 5294 2268 5300 2269
rect 5294 2264 5295 2268
rect 5299 2264 5300 2268
rect 5294 2263 5300 2264
rect 5446 2268 5452 2269
rect 5446 2264 5447 2268
rect 5451 2264 5452 2268
rect 5446 2263 5452 2264
rect 5662 2267 5668 2268
rect 5662 2263 5663 2267
rect 5667 2263 5668 2267
rect 3838 2262 3844 2263
rect 5662 2262 5668 2263
rect 110 2259 116 2260
rect 1934 2259 1940 2260
rect 1974 2232 1980 2233
rect 3798 2232 3804 2233
rect 1974 2228 1975 2232
rect 1979 2228 1980 2232
rect 1974 2227 1980 2228
rect 2042 2231 2048 2232
rect 2042 2227 2043 2231
rect 2047 2227 2048 2231
rect 2042 2226 2048 2227
rect 2178 2231 2184 2232
rect 2178 2227 2179 2231
rect 2183 2227 2184 2231
rect 2178 2226 2184 2227
rect 2314 2231 2320 2232
rect 2314 2227 2315 2231
rect 2319 2227 2320 2231
rect 2314 2226 2320 2227
rect 2450 2231 2456 2232
rect 2450 2227 2451 2231
rect 2455 2227 2456 2231
rect 2450 2226 2456 2227
rect 2586 2231 2592 2232
rect 2586 2227 2587 2231
rect 2591 2227 2592 2231
rect 2586 2226 2592 2227
rect 2722 2231 2728 2232
rect 2722 2227 2723 2231
rect 2727 2227 2728 2231
rect 2722 2226 2728 2227
rect 2858 2231 2864 2232
rect 2858 2227 2859 2231
rect 2863 2227 2864 2231
rect 2858 2226 2864 2227
rect 2994 2231 3000 2232
rect 2994 2227 2995 2231
rect 2999 2227 3000 2231
rect 2994 2226 3000 2227
rect 3130 2231 3136 2232
rect 3130 2227 3131 2231
rect 3135 2227 3136 2231
rect 3798 2228 3799 2232
rect 3803 2228 3804 2232
rect 3798 2227 3804 2228
rect 3130 2226 3136 2227
rect 2070 2216 2076 2217
rect 1974 2215 1980 2216
rect 1974 2211 1975 2215
rect 1979 2211 1980 2215
rect 2070 2212 2071 2216
rect 2075 2212 2076 2216
rect 2070 2211 2076 2212
rect 2206 2216 2212 2217
rect 2206 2212 2207 2216
rect 2211 2212 2212 2216
rect 2206 2211 2212 2212
rect 2342 2216 2348 2217
rect 2342 2212 2343 2216
rect 2347 2212 2348 2216
rect 2342 2211 2348 2212
rect 2478 2216 2484 2217
rect 2478 2212 2479 2216
rect 2483 2212 2484 2216
rect 2478 2211 2484 2212
rect 2614 2216 2620 2217
rect 2614 2212 2615 2216
rect 2619 2212 2620 2216
rect 2614 2211 2620 2212
rect 2750 2216 2756 2217
rect 2750 2212 2751 2216
rect 2755 2212 2756 2216
rect 2750 2211 2756 2212
rect 2886 2216 2892 2217
rect 2886 2212 2887 2216
rect 2891 2212 2892 2216
rect 2886 2211 2892 2212
rect 3022 2216 3028 2217
rect 3022 2212 3023 2216
rect 3027 2212 3028 2216
rect 3022 2211 3028 2212
rect 3158 2216 3164 2217
rect 3158 2212 3159 2216
rect 3163 2212 3164 2216
rect 3158 2211 3164 2212
rect 3798 2215 3804 2216
rect 3798 2211 3799 2215
rect 3803 2211 3804 2215
rect 1974 2210 1980 2211
rect 3798 2210 3804 2211
rect 3838 2197 3844 2198
rect 5662 2197 5668 2198
rect 3838 2193 3839 2197
rect 3843 2193 3844 2197
rect 3838 2192 3844 2193
rect 3886 2196 3892 2197
rect 3886 2192 3887 2196
rect 3891 2192 3892 2196
rect 3886 2191 3892 2192
rect 4166 2196 4172 2197
rect 4166 2192 4167 2196
rect 4171 2192 4172 2196
rect 4166 2191 4172 2192
rect 4454 2196 4460 2197
rect 4454 2192 4455 2196
rect 4459 2192 4460 2196
rect 4454 2191 4460 2192
rect 4718 2196 4724 2197
rect 4718 2192 4719 2196
rect 4723 2192 4724 2196
rect 4718 2191 4724 2192
rect 4974 2196 4980 2197
rect 4974 2192 4975 2196
rect 4979 2192 4980 2196
rect 4974 2191 4980 2192
rect 5230 2196 5236 2197
rect 5230 2192 5231 2196
rect 5235 2192 5236 2196
rect 5230 2191 5236 2192
rect 5486 2196 5492 2197
rect 5486 2192 5487 2196
rect 5491 2192 5492 2196
rect 5662 2193 5663 2197
rect 5667 2193 5668 2197
rect 5662 2192 5668 2193
rect 5486 2191 5492 2192
rect 3858 2181 3864 2182
rect 3838 2180 3844 2181
rect 3838 2176 3839 2180
rect 3843 2176 3844 2180
rect 3858 2177 3859 2181
rect 3863 2177 3864 2181
rect 3858 2176 3864 2177
rect 4138 2181 4144 2182
rect 4138 2177 4139 2181
rect 4143 2177 4144 2181
rect 4138 2176 4144 2177
rect 4426 2181 4432 2182
rect 4426 2177 4427 2181
rect 4431 2177 4432 2181
rect 4426 2176 4432 2177
rect 4690 2181 4696 2182
rect 4690 2177 4691 2181
rect 4695 2177 4696 2181
rect 4690 2176 4696 2177
rect 4946 2181 4952 2182
rect 4946 2177 4947 2181
rect 4951 2177 4952 2181
rect 4946 2176 4952 2177
rect 5202 2181 5208 2182
rect 5202 2177 5203 2181
rect 5207 2177 5208 2181
rect 5202 2176 5208 2177
rect 5458 2181 5464 2182
rect 5458 2177 5459 2181
rect 5463 2177 5464 2181
rect 5458 2176 5464 2177
rect 5662 2180 5668 2181
rect 5662 2176 5663 2180
rect 5667 2176 5668 2180
rect 3838 2175 3844 2176
rect 5662 2175 5668 2176
rect 1974 2157 1980 2158
rect 3798 2157 3804 2158
rect 1974 2153 1975 2157
rect 1979 2153 1980 2157
rect 1974 2152 1980 2153
rect 2022 2156 2028 2157
rect 2022 2152 2023 2156
rect 2027 2152 2028 2156
rect 2022 2151 2028 2152
rect 2238 2156 2244 2157
rect 2238 2152 2239 2156
rect 2243 2152 2244 2156
rect 2238 2151 2244 2152
rect 2486 2156 2492 2157
rect 2486 2152 2487 2156
rect 2491 2152 2492 2156
rect 2486 2151 2492 2152
rect 2726 2156 2732 2157
rect 2726 2152 2727 2156
rect 2731 2152 2732 2156
rect 2726 2151 2732 2152
rect 2966 2156 2972 2157
rect 2966 2152 2967 2156
rect 2971 2152 2972 2156
rect 2966 2151 2972 2152
rect 3206 2156 3212 2157
rect 3206 2152 3207 2156
rect 3211 2152 3212 2156
rect 3206 2151 3212 2152
rect 3454 2156 3460 2157
rect 3454 2152 3455 2156
rect 3459 2152 3460 2156
rect 3454 2151 3460 2152
rect 3678 2156 3684 2157
rect 3678 2152 3679 2156
rect 3683 2152 3684 2156
rect 3798 2153 3799 2157
rect 3803 2153 3804 2157
rect 3798 2152 3804 2153
rect 3678 2151 3684 2152
rect 1994 2141 2000 2142
rect 1974 2140 1980 2141
rect 1974 2136 1975 2140
rect 1979 2136 1980 2140
rect 1994 2137 1995 2141
rect 1999 2137 2000 2141
rect 1994 2136 2000 2137
rect 2210 2141 2216 2142
rect 2210 2137 2211 2141
rect 2215 2137 2216 2141
rect 2210 2136 2216 2137
rect 2458 2141 2464 2142
rect 2458 2137 2459 2141
rect 2463 2137 2464 2141
rect 2458 2136 2464 2137
rect 2698 2141 2704 2142
rect 2698 2137 2699 2141
rect 2703 2137 2704 2141
rect 2698 2136 2704 2137
rect 2938 2141 2944 2142
rect 2938 2137 2939 2141
rect 2943 2137 2944 2141
rect 2938 2136 2944 2137
rect 3178 2141 3184 2142
rect 3178 2137 3179 2141
rect 3183 2137 3184 2141
rect 3178 2136 3184 2137
rect 3426 2141 3432 2142
rect 3426 2137 3427 2141
rect 3431 2137 3432 2141
rect 3426 2136 3432 2137
rect 3650 2141 3656 2142
rect 3650 2137 3651 2141
rect 3655 2137 3656 2141
rect 3650 2136 3656 2137
rect 3798 2140 3804 2141
rect 3798 2136 3799 2140
rect 3803 2136 3804 2140
rect 1974 2135 1980 2136
rect 3798 2135 3804 2136
rect 110 2124 116 2125
rect 1934 2124 1940 2125
rect 110 2120 111 2124
rect 115 2120 116 2124
rect 110 2119 116 2120
rect 322 2123 328 2124
rect 322 2119 323 2123
rect 327 2119 328 2123
rect 322 2118 328 2119
rect 458 2123 464 2124
rect 458 2119 459 2123
rect 463 2119 464 2123
rect 458 2118 464 2119
rect 594 2123 600 2124
rect 594 2119 595 2123
rect 599 2119 600 2123
rect 594 2118 600 2119
rect 730 2123 736 2124
rect 730 2119 731 2123
rect 735 2119 736 2123
rect 730 2118 736 2119
rect 866 2123 872 2124
rect 866 2119 867 2123
rect 871 2119 872 2123
rect 1934 2120 1935 2124
rect 1939 2120 1940 2124
rect 1934 2119 1940 2120
rect 866 2118 872 2119
rect 350 2108 356 2109
rect 110 2107 116 2108
rect 110 2103 111 2107
rect 115 2103 116 2107
rect 350 2104 351 2108
rect 355 2104 356 2108
rect 350 2103 356 2104
rect 486 2108 492 2109
rect 486 2104 487 2108
rect 491 2104 492 2108
rect 486 2103 492 2104
rect 622 2108 628 2109
rect 622 2104 623 2108
rect 627 2104 628 2108
rect 622 2103 628 2104
rect 758 2108 764 2109
rect 758 2104 759 2108
rect 763 2104 764 2108
rect 758 2103 764 2104
rect 894 2108 900 2109
rect 894 2104 895 2108
rect 899 2104 900 2108
rect 894 2103 900 2104
rect 1934 2107 1940 2108
rect 1934 2103 1935 2107
rect 1939 2103 1940 2107
rect 110 2102 116 2103
rect 1934 2102 1940 2103
rect 3838 2048 3844 2049
rect 5662 2048 5668 2049
rect 3838 2044 3839 2048
rect 3843 2044 3844 2048
rect 3838 2043 3844 2044
rect 3858 2047 3864 2048
rect 3858 2043 3859 2047
rect 3863 2043 3864 2047
rect 3858 2042 3864 2043
rect 4082 2047 4088 2048
rect 4082 2043 4083 2047
rect 4087 2043 4088 2047
rect 4082 2042 4088 2043
rect 4322 2047 4328 2048
rect 4322 2043 4323 2047
rect 4327 2043 4328 2047
rect 4322 2042 4328 2043
rect 4546 2047 4552 2048
rect 4546 2043 4547 2047
rect 4551 2043 4552 2047
rect 4546 2042 4552 2043
rect 4754 2047 4760 2048
rect 4754 2043 4755 2047
rect 4759 2043 4760 2047
rect 4754 2042 4760 2043
rect 4946 2047 4952 2048
rect 4946 2043 4947 2047
rect 4951 2043 4952 2047
rect 4946 2042 4952 2043
rect 5138 2047 5144 2048
rect 5138 2043 5139 2047
rect 5143 2043 5144 2047
rect 5138 2042 5144 2043
rect 5322 2047 5328 2048
rect 5322 2043 5323 2047
rect 5327 2043 5328 2047
rect 5322 2042 5328 2043
rect 5514 2047 5520 2048
rect 5514 2043 5515 2047
rect 5519 2043 5520 2047
rect 5662 2044 5663 2048
rect 5667 2044 5668 2048
rect 5662 2043 5668 2044
rect 5514 2042 5520 2043
rect 3886 2032 3892 2033
rect 3838 2031 3844 2032
rect 3838 2027 3839 2031
rect 3843 2027 3844 2031
rect 3886 2028 3887 2032
rect 3891 2028 3892 2032
rect 3886 2027 3892 2028
rect 4110 2032 4116 2033
rect 4110 2028 4111 2032
rect 4115 2028 4116 2032
rect 4110 2027 4116 2028
rect 4350 2032 4356 2033
rect 4350 2028 4351 2032
rect 4355 2028 4356 2032
rect 4350 2027 4356 2028
rect 4574 2032 4580 2033
rect 4574 2028 4575 2032
rect 4579 2028 4580 2032
rect 4574 2027 4580 2028
rect 4782 2032 4788 2033
rect 4782 2028 4783 2032
rect 4787 2028 4788 2032
rect 4782 2027 4788 2028
rect 4974 2032 4980 2033
rect 4974 2028 4975 2032
rect 4979 2028 4980 2032
rect 4974 2027 4980 2028
rect 5166 2032 5172 2033
rect 5166 2028 5167 2032
rect 5171 2028 5172 2032
rect 5166 2027 5172 2028
rect 5350 2032 5356 2033
rect 5350 2028 5351 2032
rect 5355 2028 5356 2032
rect 5350 2027 5356 2028
rect 5542 2032 5548 2033
rect 5542 2028 5543 2032
rect 5547 2028 5548 2032
rect 5542 2027 5548 2028
rect 5662 2031 5668 2032
rect 5662 2027 5663 2031
rect 5667 2027 5668 2031
rect 3838 2026 3844 2027
rect 5662 2026 5668 2027
rect 110 2017 116 2018
rect 1934 2017 1940 2018
rect 110 2013 111 2017
rect 115 2013 116 2017
rect 110 2012 116 2013
rect 318 2016 324 2017
rect 318 2012 319 2016
rect 323 2012 324 2016
rect 318 2011 324 2012
rect 478 2016 484 2017
rect 478 2012 479 2016
rect 483 2012 484 2016
rect 478 2011 484 2012
rect 662 2016 668 2017
rect 662 2012 663 2016
rect 667 2012 668 2016
rect 662 2011 668 2012
rect 870 2016 876 2017
rect 870 2012 871 2016
rect 875 2012 876 2016
rect 870 2011 876 2012
rect 1094 2016 1100 2017
rect 1094 2012 1095 2016
rect 1099 2012 1100 2016
rect 1094 2011 1100 2012
rect 1334 2016 1340 2017
rect 1334 2012 1335 2016
rect 1339 2012 1340 2016
rect 1334 2011 1340 2012
rect 1582 2016 1588 2017
rect 1582 2012 1583 2016
rect 1587 2012 1588 2016
rect 1582 2011 1588 2012
rect 1814 2016 1820 2017
rect 1814 2012 1815 2016
rect 1819 2012 1820 2016
rect 1934 2013 1935 2017
rect 1939 2013 1940 2017
rect 1934 2012 1940 2013
rect 1814 2011 1820 2012
rect 290 2001 296 2002
rect 110 2000 116 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 290 1997 291 2001
rect 295 1997 296 2001
rect 290 1996 296 1997
rect 450 2001 456 2002
rect 450 1997 451 2001
rect 455 1997 456 2001
rect 450 1996 456 1997
rect 634 2001 640 2002
rect 634 1997 635 2001
rect 639 1997 640 2001
rect 634 1996 640 1997
rect 842 2001 848 2002
rect 842 1997 843 2001
rect 847 1997 848 2001
rect 842 1996 848 1997
rect 1066 2001 1072 2002
rect 1066 1997 1067 2001
rect 1071 1997 1072 2001
rect 1066 1996 1072 1997
rect 1306 2001 1312 2002
rect 1306 1997 1307 2001
rect 1311 1997 1312 2001
rect 1306 1996 1312 1997
rect 1554 2001 1560 2002
rect 1554 1997 1555 2001
rect 1559 1997 1560 2001
rect 1554 1996 1560 1997
rect 1786 2001 1792 2002
rect 1786 1997 1787 2001
rect 1791 1997 1792 2001
rect 1786 1996 1792 1997
rect 1934 2000 1940 2001
rect 1934 1996 1935 2000
rect 1939 1996 1940 2000
rect 110 1995 116 1996
rect 1934 1995 1940 1996
rect 1974 1992 1980 1993
rect 3798 1992 3804 1993
rect 1974 1988 1975 1992
rect 1979 1988 1980 1992
rect 1974 1987 1980 1988
rect 1994 1991 2000 1992
rect 1994 1987 1995 1991
rect 1999 1987 2000 1991
rect 1994 1986 2000 1987
rect 2210 1991 2216 1992
rect 2210 1987 2211 1991
rect 2215 1987 2216 1991
rect 2210 1986 2216 1987
rect 2458 1991 2464 1992
rect 2458 1987 2459 1991
rect 2463 1987 2464 1991
rect 2458 1986 2464 1987
rect 2706 1991 2712 1992
rect 2706 1987 2707 1991
rect 2711 1987 2712 1991
rect 2706 1986 2712 1987
rect 2962 1991 2968 1992
rect 2962 1987 2963 1991
rect 2967 1987 2968 1991
rect 2962 1986 2968 1987
rect 3218 1991 3224 1992
rect 3218 1987 3219 1991
rect 3223 1987 3224 1991
rect 3218 1986 3224 1987
rect 3482 1991 3488 1992
rect 3482 1987 3483 1991
rect 3487 1987 3488 1991
rect 3798 1988 3799 1992
rect 3803 1988 3804 1992
rect 3798 1987 3804 1988
rect 3482 1986 3488 1987
rect 2022 1976 2028 1977
rect 1974 1975 1980 1976
rect 1974 1971 1975 1975
rect 1979 1971 1980 1975
rect 2022 1972 2023 1976
rect 2027 1972 2028 1976
rect 2022 1971 2028 1972
rect 2238 1976 2244 1977
rect 2238 1972 2239 1976
rect 2243 1972 2244 1976
rect 2238 1971 2244 1972
rect 2486 1976 2492 1977
rect 2486 1972 2487 1976
rect 2491 1972 2492 1976
rect 2486 1971 2492 1972
rect 2734 1976 2740 1977
rect 2734 1972 2735 1976
rect 2739 1972 2740 1976
rect 2734 1971 2740 1972
rect 2990 1976 2996 1977
rect 2990 1972 2991 1976
rect 2995 1972 2996 1976
rect 2990 1971 2996 1972
rect 3246 1976 3252 1977
rect 3246 1972 3247 1976
rect 3251 1972 3252 1976
rect 3246 1971 3252 1972
rect 3510 1976 3516 1977
rect 3510 1972 3511 1976
rect 3515 1972 3516 1976
rect 3510 1971 3516 1972
rect 3798 1975 3804 1976
rect 3798 1971 3799 1975
rect 3803 1971 3804 1975
rect 1974 1970 1980 1971
rect 3798 1970 3804 1971
rect 3838 1973 3844 1974
rect 5662 1973 5668 1974
rect 3838 1969 3839 1973
rect 3843 1969 3844 1973
rect 3838 1968 3844 1969
rect 3886 1972 3892 1973
rect 3886 1968 3887 1972
rect 3891 1968 3892 1972
rect 3886 1967 3892 1968
rect 4166 1972 4172 1973
rect 4166 1968 4167 1972
rect 4171 1968 4172 1972
rect 4166 1967 4172 1968
rect 4462 1972 4468 1973
rect 4462 1968 4463 1972
rect 4467 1968 4468 1972
rect 4462 1967 4468 1968
rect 4742 1972 4748 1973
rect 4742 1968 4743 1972
rect 4747 1968 4748 1972
rect 4742 1967 4748 1968
rect 5006 1972 5012 1973
rect 5006 1968 5007 1972
rect 5011 1968 5012 1972
rect 5006 1967 5012 1968
rect 5270 1972 5276 1973
rect 5270 1968 5271 1972
rect 5275 1968 5276 1972
rect 5270 1967 5276 1968
rect 5542 1972 5548 1973
rect 5542 1968 5543 1972
rect 5547 1968 5548 1972
rect 5662 1969 5663 1973
rect 5667 1969 5668 1973
rect 5662 1968 5668 1969
rect 5542 1967 5548 1968
rect 3858 1957 3864 1958
rect 3838 1956 3844 1957
rect 3838 1952 3839 1956
rect 3843 1952 3844 1956
rect 3858 1953 3859 1957
rect 3863 1953 3864 1957
rect 3858 1952 3864 1953
rect 4138 1957 4144 1958
rect 4138 1953 4139 1957
rect 4143 1953 4144 1957
rect 4138 1952 4144 1953
rect 4434 1957 4440 1958
rect 4434 1953 4435 1957
rect 4439 1953 4440 1957
rect 4434 1952 4440 1953
rect 4714 1957 4720 1958
rect 4714 1953 4715 1957
rect 4719 1953 4720 1957
rect 4714 1952 4720 1953
rect 4978 1957 4984 1958
rect 4978 1953 4979 1957
rect 4983 1953 4984 1957
rect 4978 1952 4984 1953
rect 5242 1957 5248 1958
rect 5242 1953 5243 1957
rect 5247 1953 5248 1957
rect 5242 1952 5248 1953
rect 5514 1957 5520 1958
rect 5514 1953 5515 1957
rect 5519 1953 5520 1957
rect 5514 1952 5520 1953
rect 5662 1956 5668 1957
rect 5662 1952 5663 1956
rect 5667 1952 5668 1956
rect 3838 1951 3844 1952
rect 5662 1951 5668 1952
rect 1974 1909 1980 1910
rect 3798 1909 3804 1910
rect 1974 1905 1975 1909
rect 1979 1905 1980 1909
rect 1974 1904 1980 1905
rect 2158 1908 2164 1909
rect 2158 1904 2159 1908
rect 2163 1904 2164 1908
rect 2158 1903 2164 1904
rect 2438 1908 2444 1909
rect 2438 1904 2439 1908
rect 2443 1904 2444 1908
rect 2438 1903 2444 1904
rect 2702 1908 2708 1909
rect 2702 1904 2703 1908
rect 2707 1904 2708 1908
rect 2702 1903 2708 1904
rect 2958 1908 2964 1909
rect 2958 1904 2959 1908
rect 2963 1904 2964 1908
rect 2958 1903 2964 1904
rect 3206 1908 3212 1909
rect 3206 1904 3207 1908
rect 3211 1904 3212 1908
rect 3206 1903 3212 1904
rect 3454 1908 3460 1909
rect 3454 1904 3455 1908
rect 3459 1904 3460 1908
rect 3454 1903 3460 1904
rect 3678 1908 3684 1909
rect 3678 1904 3679 1908
rect 3683 1904 3684 1908
rect 3798 1905 3799 1909
rect 3803 1905 3804 1909
rect 3798 1904 3804 1905
rect 3678 1903 3684 1904
rect 2130 1893 2136 1894
rect 1974 1892 1980 1893
rect 1974 1888 1975 1892
rect 1979 1888 1980 1892
rect 2130 1889 2131 1893
rect 2135 1889 2136 1893
rect 2130 1888 2136 1889
rect 2410 1893 2416 1894
rect 2410 1889 2411 1893
rect 2415 1889 2416 1893
rect 2410 1888 2416 1889
rect 2674 1893 2680 1894
rect 2674 1889 2675 1893
rect 2679 1889 2680 1893
rect 2674 1888 2680 1889
rect 2930 1893 2936 1894
rect 2930 1889 2931 1893
rect 2935 1889 2936 1893
rect 2930 1888 2936 1889
rect 3178 1893 3184 1894
rect 3178 1889 3179 1893
rect 3183 1889 3184 1893
rect 3178 1888 3184 1889
rect 3426 1893 3432 1894
rect 3426 1889 3427 1893
rect 3431 1889 3432 1893
rect 3426 1888 3432 1889
rect 3650 1893 3656 1894
rect 3650 1889 3651 1893
rect 3655 1889 3656 1893
rect 3650 1888 3656 1889
rect 3798 1892 3804 1893
rect 3798 1888 3799 1892
rect 3803 1888 3804 1892
rect 1974 1887 1980 1888
rect 3798 1887 3804 1888
rect 110 1860 116 1861
rect 1934 1860 1940 1861
rect 110 1856 111 1860
rect 115 1856 116 1860
rect 110 1855 116 1856
rect 186 1859 192 1860
rect 186 1855 187 1859
rect 191 1855 192 1859
rect 186 1854 192 1855
rect 418 1859 424 1860
rect 418 1855 419 1859
rect 423 1855 424 1859
rect 418 1854 424 1855
rect 650 1859 656 1860
rect 650 1855 651 1859
rect 655 1855 656 1859
rect 650 1854 656 1855
rect 882 1859 888 1860
rect 882 1855 883 1859
rect 887 1855 888 1859
rect 882 1854 888 1855
rect 1114 1859 1120 1860
rect 1114 1855 1115 1859
rect 1119 1855 1120 1859
rect 1114 1854 1120 1855
rect 1346 1859 1352 1860
rect 1346 1855 1347 1859
rect 1351 1855 1352 1859
rect 1346 1854 1352 1855
rect 1578 1859 1584 1860
rect 1578 1855 1579 1859
rect 1583 1855 1584 1859
rect 1578 1854 1584 1855
rect 1786 1859 1792 1860
rect 1786 1855 1787 1859
rect 1791 1855 1792 1859
rect 1934 1856 1935 1860
rect 1939 1856 1940 1860
rect 1934 1855 1940 1856
rect 1786 1854 1792 1855
rect 214 1844 220 1845
rect 110 1843 116 1844
rect 110 1839 111 1843
rect 115 1839 116 1843
rect 214 1840 215 1844
rect 219 1840 220 1844
rect 214 1839 220 1840
rect 446 1844 452 1845
rect 446 1840 447 1844
rect 451 1840 452 1844
rect 446 1839 452 1840
rect 678 1844 684 1845
rect 678 1840 679 1844
rect 683 1840 684 1844
rect 678 1839 684 1840
rect 910 1844 916 1845
rect 910 1840 911 1844
rect 915 1840 916 1844
rect 910 1839 916 1840
rect 1142 1844 1148 1845
rect 1142 1840 1143 1844
rect 1147 1840 1148 1844
rect 1142 1839 1148 1840
rect 1374 1844 1380 1845
rect 1374 1840 1375 1844
rect 1379 1840 1380 1844
rect 1374 1839 1380 1840
rect 1606 1844 1612 1845
rect 1606 1840 1607 1844
rect 1611 1840 1612 1844
rect 1606 1839 1612 1840
rect 1814 1844 1820 1845
rect 1814 1840 1815 1844
rect 1819 1840 1820 1844
rect 1814 1839 1820 1840
rect 1934 1843 1940 1844
rect 1934 1839 1935 1843
rect 1939 1839 1940 1843
rect 110 1838 116 1839
rect 1934 1838 1940 1839
rect 3838 1812 3844 1813
rect 5662 1812 5668 1813
rect 3838 1808 3839 1812
rect 3843 1808 3844 1812
rect 3838 1807 3844 1808
rect 4538 1811 4544 1812
rect 4538 1807 4539 1811
rect 4543 1807 4544 1811
rect 4538 1806 4544 1807
rect 4722 1811 4728 1812
rect 4722 1807 4723 1811
rect 4727 1807 4728 1811
rect 4722 1806 4728 1807
rect 4914 1811 4920 1812
rect 4914 1807 4915 1811
rect 4919 1807 4920 1811
rect 4914 1806 4920 1807
rect 5114 1811 5120 1812
rect 5114 1807 5115 1811
rect 5119 1807 5120 1811
rect 5114 1806 5120 1807
rect 5322 1811 5328 1812
rect 5322 1807 5323 1811
rect 5327 1807 5328 1811
rect 5322 1806 5328 1807
rect 5514 1811 5520 1812
rect 5514 1807 5515 1811
rect 5519 1807 5520 1811
rect 5662 1808 5663 1812
rect 5667 1808 5668 1812
rect 5662 1807 5668 1808
rect 5514 1806 5520 1807
rect 4566 1796 4572 1797
rect 3838 1795 3844 1796
rect 3838 1791 3839 1795
rect 3843 1791 3844 1795
rect 4566 1792 4567 1796
rect 4571 1792 4572 1796
rect 4566 1791 4572 1792
rect 4750 1796 4756 1797
rect 4750 1792 4751 1796
rect 4755 1792 4756 1796
rect 4750 1791 4756 1792
rect 4942 1796 4948 1797
rect 4942 1792 4943 1796
rect 4947 1792 4948 1796
rect 4942 1791 4948 1792
rect 5142 1796 5148 1797
rect 5142 1792 5143 1796
rect 5147 1792 5148 1796
rect 5142 1791 5148 1792
rect 5350 1796 5356 1797
rect 5350 1792 5351 1796
rect 5355 1792 5356 1796
rect 5350 1791 5356 1792
rect 5542 1796 5548 1797
rect 5542 1792 5543 1796
rect 5547 1792 5548 1796
rect 5542 1791 5548 1792
rect 5662 1795 5668 1796
rect 5662 1791 5663 1795
rect 5667 1791 5668 1795
rect 3838 1790 3844 1791
rect 5662 1790 5668 1791
rect 110 1773 116 1774
rect 1934 1773 1940 1774
rect 110 1769 111 1773
rect 115 1769 116 1773
rect 110 1768 116 1769
rect 158 1772 164 1773
rect 158 1768 159 1772
rect 163 1768 164 1772
rect 158 1767 164 1768
rect 366 1772 372 1773
rect 366 1768 367 1772
rect 371 1768 372 1772
rect 366 1767 372 1768
rect 590 1772 596 1773
rect 590 1768 591 1772
rect 595 1768 596 1772
rect 590 1767 596 1768
rect 798 1772 804 1773
rect 798 1768 799 1772
rect 803 1768 804 1772
rect 798 1767 804 1768
rect 998 1772 1004 1773
rect 998 1768 999 1772
rect 1003 1768 1004 1772
rect 998 1767 1004 1768
rect 1190 1772 1196 1773
rect 1190 1768 1191 1772
rect 1195 1768 1196 1772
rect 1190 1767 1196 1768
rect 1374 1772 1380 1773
rect 1374 1768 1375 1772
rect 1379 1768 1380 1772
rect 1374 1767 1380 1768
rect 1558 1772 1564 1773
rect 1558 1768 1559 1772
rect 1563 1768 1564 1772
rect 1558 1767 1564 1768
rect 1750 1772 1756 1773
rect 1750 1768 1751 1772
rect 1755 1768 1756 1772
rect 1934 1769 1935 1773
rect 1939 1769 1940 1773
rect 1934 1768 1940 1769
rect 1750 1767 1756 1768
rect 130 1757 136 1758
rect 110 1756 116 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 130 1753 131 1757
rect 135 1753 136 1757
rect 130 1752 136 1753
rect 338 1757 344 1758
rect 338 1753 339 1757
rect 343 1753 344 1757
rect 338 1752 344 1753
rect 562 1757 568 1758
rect 562 1753 563 1757
rect 567 1753 568 1757
rect 562 1752 568 1753
rect 770 1757 776 1758
rect 770 1753 771 1757
rect 775 1753 776 1757
rect 770 1752 776 1753
rect 970 1757 976 1758
rect 970 1753 971 1757
rect 975 1753 976 1757
rect 970 1752 976 1753
rect 1162 1757 1168 1758
rect 1162 1753 1163 1757
rect 1167 1753 1168 1757
rect 1162 1752 1168 1753
rect 1346 1757 1352 1758
rect 1346 1753 1347 1757
rect 1351 1753 1352 1757
rect 1346 1752 1352 1753
rect 1530 1757 1536 1758
rect 1530 1753 1531 1757
rect 1535 1753 1536 1757
rect 1530 1752 1536 1753
rect 1722 1757 1728 1758
rect 1722 1753 1723 1757
rect 1727 1753 1728 1757
rect 1722 1752 1728 1753
rect 1934 1756 1940 1757
rect 1934 1752 1935 1756
rect 1939 1752 1940 1756
rect 110 1751 116 1752
rect 1934 1751 1940 1752
rect 1974 1752 1980 1753
rect 3798 1752 3804 1753
rect 1974 1748 1975 1752
rect 1979 1748 1980 1752
rect 1974 1747 1980 1748
rect 2306 1751 2312 1752
rect 2306 1747 2307 1751
rect 2311 1747 2312 1751
rect 2306 1746 2312 1747
rect 2498 1751 2504 1752
rect 2498 1747 2499 1751
rect 2503 1747 2504 1751
rect 2498 1746 2504 1747
rect 2690 1751 2696 1752
rect 2690 1747 2691 1751
rect 2695 1747 2696 1751
rect 2690 1746 2696 1747
rect 2882 1751 2888 1752
rect 2882 1747 2883 1751
rect 2887 1747 2888 1751
rect 2882 1746 2888 1747
rect 3066 1751 3072 1752
rect 3066 1747 3067 1751
rect 3071 1747 3072 1751
rect 3066 1746 3072 1747
rect 3250 1751 3256 1752
rect 3250 1747 3251 1751
rect 3255 1747 3256 1751
rect 3250 1746 3256 1747
rect 3442 1751 3448 1752
rect 3442 1747 3443 1751
rect 3447 1747 3448 1751
rect 3442 1746 3448 1747
rect 3634 1751 3640 1752
rect 3634 1747 3635 1751
rect 3639 1747 3640 1751
rect 3798 1748 3799 1752
rect 3803 1748 3804 1752
rect 3798 1747 3804 1748
rect 3634 1746 3640 1747
rect 2334 1736 2340 1737
rect 1974 1735 1980 1736
rect 1974 1731 1975 1735
rect 1979 1731 1980 1735
rect 2334 1732 2335 1736
rect 2339 1732 2340 1736
rect 2334 1731 2340 1732
rect 2526 1736 2532 1737
rect 2526 1732 2527 1736
rect 2531 1732 2532 1736
rect 2526 1731 2532 1732
rect 2718 1736 2724 1737
rect 2718 1732 2719 1736
rect 2723 1732 2724 1736
rect 2718 1731 2724 1732
rect 2910 1736 2916 1737
rect 2910 1732 2911 1736
rect 2915 1732 2916 1736
rect 2910 1731 2916 1732
rect 3094 1736 3100 1737
rect 3094 1732 3095 1736
rect 3099 1732 3100 1736
rect 3094 1731 3100 1732
rect 3278 1736 3284 1737
rect 3278 1732 3279 1736
rect 3283 1732 3284 1736
rect 3278 1731 3284 1732
rect 3470 1736 3476 1737
rect 3470 1732 3471 1736
rect 3475 1732 3476 1736
rect 3470 1731 3476 1732
rect 3662 1736 3668 1737
rect 3662 1732 3663 1736
rect 3667 1732 3668 1736
rect 3662 1731 3668 1732
rect 3798 1735 3804 1736
rect 3798 1731 3799 1735
rect 3803 1731 3804 1735
rect 1974 1730 1980 1731
rect 3798 1730 3804 1731
rect 3838 1729 3844 1730
rect 5662 1729 5668 1730
rect 3838 1725 3839 1729
rect 3843 1725 3844 1729
rect 3838 1724 3844 1725
rect 4382 1728 4388 1729
rect 4382 1724 4383 1728
rect 4387 1724 4388 1728
rect 4382 1723 4388 1724
rect 4598 1728 4604 1729
rect 4598 1724 4599 1728
rect 4603 1724 4604 1728
rect 4598 1723 4604 1724
rect 4830 1728 4836 1729
rect 4830 1724 4831 1728
rect 4835 1724 4836 1728
rect 4830 1723 4836 1724
rect 5070 1728 5076 1729
rect 5070 1724 5071 1728
rect 5075 1724 5076 1728
rect 5070 1723 5076 1724
rect 5318 1728 5324 1729
rect 5318 1724 5319 1728
rect 5323 1724 5324 1728
rect 5318 1723 5324 1724
rect 5542 1728 5548 1729
rect 5542 1724 5543 1728
rect 5547 1724 5548 1728
rect 5662 1725 5663 1729
rect 5667 1725 5668 1729
rect 5662 1724 5668 1725
rect 5542 1723 5548 1724
rect 4354 1713 4360 1714
rect 3838 1712 3844 1713
rect 3838 1708 3839 1712
rect 3843 1708 3844 1712
rect 4354 1709 4355 1713
rect 4359 1709 4360 1713
rect 4354 1708 4360 1709
rect 4570 1713 4576 1714
rect 4570 1709 4571 1713
rect 4575 1709 4576 1713
rect 4570 1708 4576 1709
rect 4802 1713 4808 1714
rect 4802 1709 4803 1713
rect 4807 1709 4808 1713
rect 4802 1708 4808 1709
rect 5042 1713 5048 1714
rect 5042 1709 5043 1713
rect 5047 1709 5048 1713
rect 5042 1708 5048 1709
rect 5290 1713 5296 1714
rect 5290 1709 5291 1713
rect 5295 1709 5296 1713
rect 5290 1708 5296 1709
rect 5514 1713 5520 1714
rect 5514 1709 5515 1713
rect 5519 1709 5520 1713
rect 5514 1708 5520 1709
rect 5662 1712 5668 1713
rect 5662 1708 5663 1712
rect 5667 1708 5668 1712
rect 3838 1707 3844 1708
rect 5662 1707 5668 1708
rect 1974 1677 1980 1678
rect 3798 1677 3804 1678
rect 1974 1673 1975 1677
rect 1979 1673 1980 1677
rect 1974 1672 1980 1673
rect 2470 1676 2476 1677
rect 2470 1672 2471 1676
rect 2475 1672 2476 1676
rect 2470 1671 2476 1672
rect 2606 1676 2612 1677
rect 2606 1672 2607 1676
rect 2611 1672 2612 1676
rect 2606 1671 2612 1672
rect 2742 1676 2748 1677
rect 2742 1672 2743 1676
rect 2747 1672 2748 1676
rect 2742 1671 2748 1672
rect 2878 1676 2884 1677
rect 2878 1672 2879 1676
rect 2883 1672 2884 1676
rect 2878 1671 2884 1672
rect 3022 1676 3028 1677
rect 3022 1672 3023 1676
rect 3027 1672 3028 1676
rect 3022 1671 3028 1672
rect 3174 1676 3180 1677
rect 3174 1672 3175 1676
rect 3179 1672 3180 1676
rect 3174 1671 3180 1672
rect 3326 1676 3332 1677
rect 3326 1672 3327 1676
rect 3331 1672 3332 1676
rect 3798 1673 3799 1677
rect 3803 1673 3804 1677
rect 3798 1672 3804 1673
rect 3326 1671 3332 1672
rect 2442 1661 2448 1662
rect 1974 1660 1980 1661
rect 1974 1656 1975 1660
rect 1979 1656 1980 1660
rect 2442 1657 2443 1661
rect 2447 1657 2448 1661
rect 2442 1656 2448 1657
rect 2578 1661 2584 1662
rect 2578 1657 2579 1661
rect 2583 1657 2584 1661
rect 2578 1656 2584 1657
rect 2714 1661 2720 1662
rect 2714 1657 2715 1661
rect 2719 1657 2720 1661
rect 2714 1656 2720 1657
rect 2850 1661 2856 1662
rect 2850 1657 2851 1661
rect 2855 1657 2856 1661
rect 2850 1656 2856 1657
rect 2994 1661 3000 1662
rect 2994 1657 2995 1661
rect 2999 1657 3000 1661
rect 2994 1656 3000 1657
rect 3146 1661 3152 1662
rect 3146 1657 3147 1661
rect 3151 1657 3152 1661
rect 3146 1656 3152 1657
rect 3298 1661 3304 1662
rect 3298 1657 3299 1661
rect 3303 1657 3304 1661
rect 3298 1656 3304 1657
rect 3798 1660 3804 1661
rect 3798 1656 3799 1660
rect 3803 1656 3804 1660
rect 1974 1655 1980 1656
rect 3798 1655 3804 1656
rect 110 1616 116 1617
rect 1934 1616 1940 1617
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 354 1615 360 1616
rect 354 1611 355 1615
rect 359 1611 360 1615
rect 354 1610 360 1611
rect 594 1615 600 1616
rect 594 1611 595 1615
rect 599 1611 600 1615
rect 594 1610 600 1611
rect 834 1615 840 1616
rect 834 1611 835 1615
rect 839 1611 840 1615
rect 834 1610 840 1611
rect 1066 1615 1072 1616
rect 1066 1611 1067 1615
rect 1071 1611 1072 1615
rect 1066 1610 1072 1611
rect 1306 1615 1312 1616
rect 1306 1611 1307 1615
rect 1311 1611 1312 1615
rect 1306 1610 1312 1611
rect 1546 1615 1552 1616
rect 1546 1611 1547 1615
rect 1551 1611 1552 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 1546 1610 1552 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 382 1600 388 1601
rect 382 1596 383 1600
rect 387 1596 388 1600
rect 382 1595 388 1596
rect 622 1600 628 1601
rect 622 1596 623 1600
rect 627 1596 628 1600
rect 622 1595 628 1596
rect 862 1600 868 1601
rect 862 1596 863 1600
rect 867 1596 868 1600
rect 862 1595 868 1596
rect 1094 1600 1100 1601
rect 1094 1596 1095 1600
rect 1099 1596 1100 1600
rect 1094 1595 1100 1596
rect 1334 1600 1340 1601
rect 1334 1596 1335 1600
rect 1339 1596 1340 1600
rect 1334 1595 1340 1596
rect 1574 1600 1580 1601
rect 1574 1596 1575 1600
rect 1579 1596 1580 1600
rect 1574 1595 1580 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 110 1594 116 1595
rect 1934 1594 1940 1595
rect 3838 1568 3844 1569
rect 5662 1568 5668 1569
rect 3838 1564 3839 1568
rect 3843 1564 3844 1568
rect 3838 1563 3844 1564
rect 3906 1567 3912 1568
rect 3906 1563 3907 1567
rect 3911 1563 3912 1567
rect 3906 1562 3912 1563
rect 4122 1567 4128 1568
rect 4122 1563 4123 1567
rect 4127 1563 4128 1567
rect 4122 1562 4128 1563
rect 4362 1567 4368 1568
rect 4362 1563 4363 1567
rect 4367 1563 4368 1567
rect 4362 1562 4368 1563
rect 4626 1567 4632 1568
rect 4626 1563 4627 1567
rect 4631 1563 4632 1567
rect 4626 1562 4632 1563
rect 4906 1567 4912 1568
rect 4906 1563 4907 1567
rect 4911 1563 4912 1567
rect 4906 1562 4912 1563
rect 5194 1567 5200 1568
rect 5194 1563 5195 1567
rect 5199 1563 5200 1567
rect 5194 1562 5200 1563
rect 5490 1567 5496 1568
rect 5490 1563 5491 1567
rect 5495 1563 5496 1567
rect 5662 1564 5663 1568
rect 5667 1564 5668 1568
rect 5662 1563 5668 1564
rect 5490 1562 5496 1563
rect 3934 1552 3940 1553
rect 3838 1551 3844 1552
rect 3838 1547 3839 1551
rect 3843 1547 3844 1551
rect 3934 1548 3935 1552
rect 3939 1548 3940 1552
rect 3934 1547 3940 1548
rect 4150 1552 4156 1553
rect 4150 1548 4151 1552
rect 4155 1548 4156 1552
rect 4150 1547 4156 1548
rect 4390 1552 4396 1553
rect 4390 1548 4391 1552
rect 4395 1548 4396 1552
rect 4390 1547 4396 1548
rect 4654 1552 4660 1553
rect 4654 1548 4655 1552
rect 4659 1548 4660 1552
rect 4654 1547 4660 1548
rect 4934 1552 4940 1553
rect 4934 1548 4935 1552
rect 4939 1548 4940 1552
rect 4934 1547 4940 1548
rect 5222 1552 5228 1553
rect 5222 1548 5223 1552
rect 5227 1548 5228 1552
rect 5222 1547 5228 1548
rect 5518 1552 5524 1553
rect 5518 1548 5519 1552
rect 5523 1548 5524 1552
rect 5518 1547 5524 1548
rect 5662 1551 5668 1552
rect 5662 1547 5663 1551
rect 5667 1547 5668 1551
rect 3838 1546 3844 1547
rect 5662 1546 5668 1547
rect 110 1537 116 1538
rect 1934 1537 1940 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 110 1532 116 1533
rect 158 1536 164 1537
rect 158 1532 159 1536
rect 163 1532 164 1536
rect 158 1531 164 1532
rect 358 1536 364 1537
rect 358 1532 359 1536
rect 363 1532 364 1536
rect 358 1531 364 1532
rect 574 1536 580 1537
rect 574 1532 575 1536
rect 579 1532 580 1536
rect 574 1531 580 1532
rect 782 1536 788 1537
rect 782 1532 783 1536
rect 787 1532 788 1536
rect 782 1531 788 1532
rect 982 1536 988 1537
rect 982 1532 983 1536
rect 987 1532 988 1536
rect 982 1531 988 1532
rect 1182 1536 1188 1537
rect 1182 1532 1183 1536
rect 1187 1532 1188 1536
rect 1182 1531 1188 1532
rect 1374 1536 1380 1537
rect 1374 1532 1375 1536
rect 1379 1532 1380 1536
rect 1374 1531 1380 1532
rect 1574 1536 1580 1537
rect 1574 1532 1575 1536
rect 1579 1532 1580 1536
rect 1934 1533 1935 1537
rect 1939 1533 1940 1537
rect 1934 1532 1940 1533
rect 1574 1531 1580 1532
rect 1974 1528 1980 1529
rect 3798 1528 3804 1529
rect 1974 1524 1975 1528
rect 1979 1524 1980 1528
rect 1974 1523 1980 1524
rect 2354 1527 2360 1528
rect 2354 1523 2355 1527
rect 2359 1523 2360 1527
rect 2354 1522 2360 1523
rect 2562 1527 2568 1528
rect 2562 1523 2563 1527
rect 2567 1523 2568 1527
rect 2562 1522 2568 1523
rect 2778 1527 2784 1528
rect 2778 1523 2779 1527
rect 2783 1523 2784 1527
rect 2778 1522 2784 1523
rect 3002 1527 3008 1528
rect 3002 1523 3003 1527
rect 3007 1523 3008 1527
rect 3002 1522 3008 1523
rect 3226 1527 3232 1528
rect 3226 1523 3227 1527
rect 3231 1523 3232 1527
rect 3226 1522 3232 1523
rect 3458 1527 3464 1528
rect 3458 1523 3459 1527
rect 3463 1523 3464 1527
rect 3798 1524 3799 1528
rect 3803 1524 3804 1528
rect 3798 1523 3804 1524
rect 3458 1522 3464 1523
rect 130 1521 136 1522
rect 110 1520 116 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 130 1517 131 1521
rect 135 1517 136 1521
rect 130 1516 136 1517
rect 330 1521 336 1522
rect 330 1517 331 1521
rect 335 1517 336 1521
rect 330 1516 336 1517
rect 546 1521 552 1522
rect 546 1517 547 1521
rect 551 1517 552 1521
rect 546 1516 552 1517
rect 754 1521 760 1522
rect 754 1517 755 1521
rect 759 1517 760 1521
rect 754 1516 760 1517
rect 954 1521 960 1522
rect 954 1517 955 1521
rect 959 1517 960 1521
rect 954 1516 960 1517
rect 1154 1521 1160 1522
rect 1154 1517 1155 1521
rect 1159 1517 1160 1521
rect 1154 1516 1160 1517
rect 1346 1521 1352 1522
rect 1346 1517 1347 1521
rect 1351 1517 1352 1521
rect 1346 1516 1352 1517
rect 1546 1521 1552 1522
rect 1546 1517 1547 1521
rect 1551 1517 1552 1521
rect 1546 1516 1552 1517
rect 1934 1520 1940 1521
rect 1934 1516 1935 1520
rect 1939 1516 1940 1520
rect 110 1515 116 1516
rect 1934 1515 1940 1516
rect 2382 1512 2388 1513
rect 1974 1511 1980 1512
rect 1974 1507 1975 1511
rect 1979 1507 1980 1511
rect 2382 1508 2383 1512
rect 2387 1508 2388 1512
rect 2382 1507 2388 1508
rect 2590 1512 2596 1513
rect 2590 1508 2591 1512
rect 2595 1508 2596 1512
rect 2590 1507 2596 1508
rect 2806 1512 2812 1513
rect 2806 1508 2807 1512
rect 2811 1508 2812 1512
rect 2806 1507 2812 1508
rect 3030 1512 3036 1513
rect 3030 1508 3031 1512
rect 3035 1508 3036 1512
rect 3030 1507 3036 1508
rect 3254 1512 3260 1513
rect 3254 1508 3255 1512
rect 3259 1508 3260 1512
rect 3254 1507 3260 1508
rect 3486 1512 3492 1513
rect 3486 1508 3487 1512
rect 3491 1508 3492 1512
rect 3486 1507 3492 1508
rect 3798 1511 3804 1512
rect 3798 1507 3799 1511
rect 3803 1507 3804 1511
rect 1974 1506 1980 1507
rect 3798 1506 3804 1507
rect 3838 1493 3844 1494
rect 5662 1493 5668 1494
rect 3838 1489 3839 1493
rect 3843 1489 3844 1493
rect 3838 1488 3844 1489
rect 3886 1492 3892 1493
rect 3886 1488 3887 1492
rect 3891 1488 3892 1492
rect 3886 1487 3892 1488
rect 4022 1492 4028 1493
rect 4022 1488 4023 1492
rect 4027 1488 4028 1492
rect 4022 1487 4028 1488
rect 4158 1492 4164 1493
rect 4158 1488 4159 1492
rect 4163 1488 4164 1492
rect 4158 1487 4164 1488
rect 4294 1492 4300 1493
rect 4294 1488 4295 1492
rect 4299 1488 4300 1492
rect 4294 1487 4300 1488
rect 4478 1492 4484 1493
rect 4478 1488 4479 1492
rect 4483 1488 4484 1492
rect 4478 1487 4484 1488
rect 4694 1492 4700 1493
rect 4694 1488 4695 1492
rect 4699 1488 4700 1492
rect 4694 1487 4700 1488
rect 4934 1492 4940 1493
rect 4934 1488 4935 1492
rect 4939 1488 4940 1492
rect 4934 1487 4940 1488
rect 5190 1492 5196 1493
rect 5190 1488 5191 1492
rect 5195 1488 5196 1492
rect 5190 1487 5196 1488
rect 5446 1492 5452 1493
rect 5446 1488 5447 1492
rect 5451 1488 5452 1492
rect 5662 1489 5663 1493
rect 5667 1489 5668 1493
rect 5662 1488 5668 1489
rect 5446 1487 5452 1488
rect 3858 1477 3864 1478
rect 3838 1476 3844 1477
rect 3838 1472 3839 1476
rect 3843 1472 3844 1476
rect 3858 1473 3859 1477
rect 3863 1473 3864 1477
rect 3858 1472 3864 1473
rect 3994 1477 4000 1478
rect 3994 1473 3995 1477
rect 3999 1473 4000 1477
rect 3994 1472 4000 1473
rect 4130 1477 4136 1478
rect 4130 1473 4131 1477
rect 4135 1473 4136 1477
rect 4130 1472 4136 1473
rect 4266 1477 4272 1478
rect 4266 1473 4267 1477
rect 4271 1473 4272 1477
rect 4266 1472 4272 1473
rect 4450 1477 4456 1478
rect 4450 1473 4451 1477
rect 4455 1473 4456 1477
rect 4450 1472 4456 1473
rect 4666 1477 4672 1478
rect 4666 1473 4667 1477
rect 4671 1473 4672 1477
rect 4666 1472 4672 1473
rect 4906 1477 4912 1478
rect 4906 1473 4907 1477
rect 4911 1473 4912 1477
rect 4906 1472 4912 1473
rect 5162 1477 5168 1478
rect 5162 1473 5163 1477
rect 5167 1473 5168 1477
rect 5162 1472 5168 1473
rect 5418 1477 5424 1478
rect 5418 1473 5419 1477
rect 5423 1473 5424 1477
rect 5418 1472 5424 1473
rect 5662 1476 5668 1477
rect 5662 1472 5663 1476
rect 5667 1472 5668 1476
rect 3838 1471 3844 1472
rect 5662 1471 5668 1472
rect 1974 1453 1980 1454
rect 3798 1453 3804 1454
rect 1974 1449 1975 1453
rect 1979 1449 1980 1453
rect 1974 1448 1980 1449
rect 2022 1452 2028 1453
rect 2022 1448 2023 1452
rect 2027 1448 2028 1452
rect 2022 1447 2028 1448
rect 2158 1452 2164 1453
rect 2158 1448 2159 1452
rect 2163 1448 2164 1452
rect 2158 1447 2164 1448
rect 2326 1452 2332 1453
rect 2326 1448 2327 1452
rect 2331 1448 2332 1452
rect 2326 1447 2332 1448
rect 2542 1452 2548 1453
rect 2542 1448 2543 1452
rect 2547 1448 2548 1452
rect 2542 1447 2548 1448
rect 2798 1452 2804 1453
rect 2798 1448 2799 1452
rect 2803 1448 2804 1452
rect 2798 1447 2804 1448
rect 3086 1452 3092 1453
rect 3086 1448 3087 1452
rect 3091 1448 3092 1452
rect 3086 1447 3092 1448
rect 3390 1452 3396 1453
rect 3390 1448 3391 1452
rect 3395 1448 3396 1452
rect 3390 1447 3396 1448
rect 3678 1452 3684 1453
rect 3678 1448 3679 1452
rect 3683 1448 3684 1452
rect 3798 1449 3799 1453
rect 3803 1449 3804 1453
rect 3798 1448 3804 1449
rect 3678 1447 3684 1448
rect 1994 1437 2000 1438
rect 1974 1436 1980 1437
rect 1974 1432 1975 1436
rect 1979 1432 1980 1436
rect 1994 1433 1995 1437
rect 1999 1433 2000 1437
rect 1994 1432 2000 1433
rect 2130 1437 2136 1438
rect 2130 1433 2131 1437
rect 2135 1433 2136 1437
rect 2130 1432 2136 1433
rect 2298 1437 2304 1438
rect 2298 1433 2299 1437
rect 2303 1433 2304 1437
rect 2298 1432 2304 1433
rect 2514 1437 2520 1438
rect 2514 1433 2515 1437
rect 2519 1433 2520 1437
rect 2514 1432 2520 1433
rect 2770 1437 2776 1438
rect 2770 1433 2771 1437
rect 2775 1433 2776 1437
rect 2770 1432 2776 1433
rect 3058 1437 3064 1438
rect 3058 1433 3059 1437
rect 3063 1433 3064 1437
rect 3058 1432 3064 1433
rect 3362 1437 3368 1438
rect 3362 1433 3363 1437
rect 3367 1433 3368 1437
rect 3362 1432 3368 1433
rect 3650 1437 3656 1438
rect 3650 1433 3651 1437
rect 3655 1433 3656 1437
rect 3650 1432 3656 1433
rect 3798 1436 3804 1437
rect 3798 1432 3799 1436
rect 3803 1432 3804 1436
rect 1974 1431 1980 1432
rect 3798 1431 3804 1432
rect 110 1368 116 1369
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 234 1367 240 1368
rect 234 1363 235 1367
rect 239 1363 240 1367
rect 234 1362 240 1363
rect 506 1367 512 1368
rect 506 1363 507 1367
rect 511 1363 512 1367
rect 506 1362 512 1363
rect 778 1367 784 1368
rect 778 1363 779 1367
rect 783 1363 784 1367
rect 778 1362 784 1363
rect 1058 1367 1064 1368
rect 1058 1363 1059 1367
rect 1063 1363 1064 1367
rect 1058 1362 1064 1363
rect 1338 1367 1344 1368
rect 1338 1363 1339 1367
rect 1343 1363 1344 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1338 1362 1344 1363
rect 262 1352 268 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 262 1348 263 1352
rect 267 1348 268 1352
rect 262 1347 268 1348
rect 534 1352 540 1353
rect 534 1348 535 1352
rect 539 1348 540 1352
rect 534 1347 540 1348
rect 806 1352 812 1353
rect 806 1348 807 1352
rect 811 1348 812 1352
rect 806 1347 812 1348
rect 1086 1352 1092 1353
rect 1086 1348 1087 1352
rect 1091 1348 1092 1352
rect 1086 1347 1092 1348
rect 1366 1352 1372 1353
rect 1366 1348 1367 1352
rect 1371 1348 1372 1352
rect 1366 1347 1372 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 110 1346 116 1347
rect 1934 1346 1940 1347
rect 3838 1332 3844 1333
rect 5662 1332 5668 1333
rect 3838 1328 3839 1332
rect 3843 1328 3844 1332
rect 3838 1327 3844 1328
rect 3858 1331 3864 1332
rect 3858 1327 3859 1331
rect 3863 1327 3864 1331
rect 3858 1326 3864 1327
rect 3994 1331 4000 1332
rect 3994 1327 3995 1331
rect 3999 1327 4000 1331
rect 3994 1326 4000 1327
rect 4146 1331 4152 1332
rect 4146 1327 4147 1331
rect 4151 1327 4152 1331
rect 4146 1326 4152 1327
rect 4362 1331 4368 1332
rect 4362 1327 4363 1331
rect 4367 1327 4368 1331
rect 4362 1326 4368 1327
rect 4610 1331 4616 1332
rect 4610 1327 4611 1331
rect 4615 1327 4616 1331
rect 4610 1326 4616 1327
rect 4890 1331 4896 1332
rect 4890 1327 4891 1331
rect 4895 1327 4896 1331
rect 4890 1326 4896 1327
rect 5194 1331 5200 1332
rect 5194 1327 5195 1331
rect 5199 1327 5200 1331
rect 5194 1326 5200 1327
rect 5498 1331 5504 1332
rect 5498 1327 5499 1331
rect 5503 1327 5504 1331
rect 5662 1328 5663 1332
rect 5667 1328 5668 1332
rect 5662 1327 5668 1328
rect 5498 1326 5504 1327
rect 3886 1316 3892 1317
rect 3838 1315 3844 1316
rect 3838 1311 3839 1315
rect 3843 1311 3844 1315
rect 3886 1312 3887 1316
rect 3891 1312 3892 1316
rect 3886 1311 3892 1312
rect 4022 1316 4028 1317
rect 4022 1312 4023 1316
rect 4027 1312 4028 1316
rect 4022 1311 4028 1312
rect 4174 1316 4180 1317
rect 4174 1312 4175 1316
rect 4179 1312 4180 1316
rect 4174 1311 4180 1312
rect 4390 1316 4396 1317
rect 4390 1312 4391 1316
rect 4395 1312 4396 1316
rect 4390 1311 4396 1312
rect 4638 1316 4644 1317
rect 4638 1312 4639 1316
rect 4643 1312 4644 1316
rect 4638 1311 4644 1312
rect 4918 1316 4924 1317
rect 4918 1312 4919 1316
rect 4923 1312 4924 1316
rect 4918 1311 4924 1312
rect 5222 1316 5228 1317
rect 5222 1312 5223 1316
rect 5227 1312 5228 1316
rect 5222 1311 5228 1312
rect 5526 1316 5532 1317
rect 5526 1312 5527 1316
rect 5531 1312 5532 1316
rect 5526 1311 5532 1312
rect 5662 1315 5668 1316
rect 5662 1311 5663 1315
rect 5667 1311 5668 1315
rect 3838 1310 3844 1311
rect 5662 1310 5668 1311
rect 1974 1304 1980 1305
rect 3798 1304 3804 1305
rect 1974 1300 1975 1304
rect 1979 1300 1980 1304
rect 1974 1299 1980 1300
rect 1994 1303 2000 1304
rect 1994 1299 1995 1303
rect 1999 1299 2000 1303
rect 1994 1298 2000 1299
rect 2490 1303 2496 1304
rect 2490 1299 2491 1303
rect 2495 1299 2496 1303
rect 2490 1298 2496 1299
rect 3018 1303 3024 1304
rect 3018 1299 3019 1303
rect 3023 1299 3024 1303
rect 3018 1298 3024 1299
rect 3554 1303 3560 1304
rect 3554 1299 3555 1303
rect 3559 1299 3560 1303
rect 3798 1300 3799 1304
rect 3803 1300 3804 1304
rect 3798 1299 3804 1300
rect 3554 1298 3560 1299
rect 110 1289 116 1290
rect 1934 1289 1940 1290
rect 110 1285 111 1289
rect 115 1285 116 1289
rect 110 1284 116 1285
rect 158 1288 164 1289
rect 158 1284 159 1288
rect 163 1284 164 1288
rect 158 1283 164 1284
rect 382 1288 388 1289
rect 382 1284 383 1288
rect 387 1284 388 1288
rect 382 1283 388 1284
rect 598 1288 604 1289
rect 598 1284 599 1288
rect 603 1284 604 1288
rect 598 1283 604 1284
rect 798 1288 804 1289
rect 798 1284 799 1288
rect 803 1284 804 1288
rect 798 1283 804 1284
rect 990 1288 996 1289
rect 990 1284 991 1288
rect 995 1284 996 1288
rect 990 1283 996 1284
rect 1166 1288 1172 1289
rect 1166 1284 1167 1288
rect 1171 1284 1172 1288
rect 1166 1283 1172 1284
rect 1334 1288 1340 1289
rect 1334 1284 1335 1288
rect 1339 1284 1340 1288
rect 1334 1283 1340 1284
rect 1502 1288 1508 1289
rect 1502 1284 1503 1288
rect 1507 1284 1508 1288
rect 1502 1283 1508 1284
rect 1670 1288 1676 1289
rect 1670 1284 1671 1288
rect 1675 1284 1676 1288
rect 1670 1283 1676 1284
rect 1814 1288 1820 1289
rect 1814 1284 1815 1288
rect 1819 1284 1820 1288
rect 1934 1285 1935 1289
rect 1939 1285 1940 1289
rect 2022 1288 2028 1289
rect 1934 1284 1940 1285
rect 1974 1287 1980 1288
rect 1814 1283 1820 1284
rect 1974 1283 1975 1287
rect 1979 1283 1980 1287
rect 2022 1284 2023 1288
rect 2027 1284 2028 1288
rect 2022 1283 2028 1284
rect 2518 1288 2524 1289
rect 2518 1284 2519 1288
rect 2523 1284 2524 1288
rect 2518 1283 2524 1284
rect 3046 1288 3052 1289
rect 3046 1284 3047 1288
rect 3051 1284 3052 1288
rect 3046 1283 3052 1284
rect 3582 1288 3588 1289
rect 3582 1284 3583 1288
rect 3587 1284 3588 1288
rect 3582 1283 3588 1284
rect 3798 1287 3804 1288
rect 3798 1283 3799 1287
rect 3803 1283 3804 1287
rect 1974 1282 1980 1283
rect 3798 1282 3804 1283
rect 130 1273 136 1274
rect 110 1272 116 1273
rect 110 1268 111 1272
rect 115 1268 116 1272
rect 130 1269 131 1273
rect 135 1269 136 1273
rect 130 1268 136 1269
rect 354 1273 360 1274
rect 354 1269 355 1273
rect 359 1269 360 1273
rect 354 1268 360 1269
rect 570 1273 576 1274
rect 570 1269 571 1273
rect 575 1269 576 1273
rect 570 1268 576 1269
rect 770 1273 776 1274
rect 770 1269 771 1273
rect 775 1269 776 1273
rect 770 1268 776 1269
rect 962 1273 968 1274
rect 962 1269 963 1273
rect 967 1269 968 1273
rect 962 1268 968 1269
rect 1138 1273 1144 1274
rect 1138 1269 1139 1273
rect 1143 1269 1144 1273
rect 1138 1268 1144 1269
rect 1306 1273 1312 1274
rect 1306 1269 1307 1273
rect 1311 1269 1312 1273
rect 1306 1268 1312 1269
rect 1474 1273 1480 1274
rect 1474 1269 1475 1273
rect 1479 1269 1480 1273
rect 1474 1268 1480 1269
rect 1642 1273 1648 1274
rect 1642 1269 1643 1273
rect 1647 1269 1648 1273
rect 1642 1268 1648 1269
rect 1786 1273 1792 1274
rect 1786 1269 1787 1273
rect 1791 1269 1792 1273
rect 1786 1268 1792 1269
rect 1934 1272 1940 1273
rect 1934 1268 1935 1272
rect 1939 1268 1940 1272
rect 110 1267 116 1268
rect 1934 1267 1940 1268
rect 3838 1257 3844 1258
rect 5662 1257 5668 1258
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 3886 1256 3892 1257
rect 3886 1252 3887 1256
rect 3891 1252 3892 1256
rect 3886 1251 3892 1252
rect 4022 1256 4028 1257
rect 4022 1252 4023 1256
rect 4027 1252 4028 1256
rect 4022 1251 4028 1252
rect 4166 1256 4172 1257
rect 4166 1252 4167 1256
rect 4171 1252 4172 1256
rect 4166 1251 4172 1252
rect 4334 1256 4340 1257
rect 4334 1252 4335 1256
rect 4339 1252 4340 1256
rect 4334 1251 4340 1252
rect 4510 1256 4516 1257
rect 4510 1252 4511 1256
rect 4515 1252 4516 1256
rect 4510 1251 4516 1252
rect 4702 1256 4708 1257
rect 4702 1252 4703 1256
rect 4707 1252 4708 1256
rect 4702 1251 4708 1252
rect 4902 1256 4908 1257
rect 4902 1252 4903 1256
rect 4907 1252 4908 1256
rect 4902 1251 4908 1252
rect 5118 1256 5124 1257
rect 5118 1252 5119 1256
rect 5123 1252 5124 1256
rect 5118 1251 5124 1252
rect 5342 1256 5348 1257
rect 5342 1252 5343 1256
rect 5347 1252 5348 1256
rect 5342 1251 5348 1252
rect 5542 1256 5548 1257
rect 5542 1252 5543 1256
rect 5547 1252 5548 1256
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5542 1251 5548 1252
rect 3858 1241 3864 1242
rect 3838 1240 3844 1241
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 3858 1237 3859 1241
rect 3863 1237 3864 1241
rect 3858 1236 3864 1237
rect 3994 1241 4000 1242
rect 3994 1237 3995 1241
rect 3999 1237 4000 1241
rect 3994 1236 4000 1237
rect 4138 1241 4144 1242
rect 4138 1237 4139 1241
rect 4143 1237 4144 1241
rect 4138 1236 4144 1237
rect 4306 1241 4312 1242
rect 4306 1237 4307 1241
rect 4311 1237 4312 1241
rect 4306 1236 4312 1237
rect 4482 1241 4488 1242
rect 4482 1237 4483 1241
rect 4487 1237 4488 1241
rect 4482 1236 4488 1237
rect 4674 1241 4680 1242
rect 4674 1237 4675 1241
rect 4679 1237 4680 1241
rect 4674 1236 4680 1237
rect 4874 1241 4880 1242
rect 4874 1237 4875 1241
rect 4879 1237 4880 1241
rect 4874 1236 4880 1237
rect 5090 1241 5096 1242
rect 5090 1237 5091 1241
rect 5095 1237 5096 1241
rect 5090 1236 5096 1237
rect 5314 1241 5320 1242
rect 5314 1237 5315 1241
rect 5319 1237 5320 1241
rect 5314 1236 5320 1237
rect 5514 1241 5520 1242
rect 5514 1237 5515 1241
rect 5519 1237 5520 1241
rect 5514 1236 5520 1237
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 3838 1235 3844 1236
rect 5662 1235 5668 1236
rect 1974 1165 1980 1166
rect 3798 1165 3804 1166
rect 1974 1161 1975 1165
rect 1979 1161 1980 1165
rect 1974 1160 1980 1161
rect 2742 1164 2748 1165
rect 2742 1160 2743 1164
rect 2747 1160 2748 1164
rect 2742 1159 2748 1160
rect 3046 1164 3052 1165
rect 3046 1160 3047 1164
rect 3051 1160 3052 1164
rect 3046 1159 3052 1160
rect 3358 1164 3364 1165
rect 3358 1160 3359 1164
rect 3363 1160 3364 1164
rect 3358 1159 3364 1160
rect 3678 1164 3684 1165
rect 3678 1160 3679 1164
rect 3683 1160 3684 1164
rect 3798 1161 3799 1165
rect 3803 1161 3804 1165
rect 3798 1160 3804 1161
rect 3678 1159 3684 1160
rect 2714 1149 2720 1150
rect 1974 1148 1980 1149
rect 1974 1144 1975 1148
rect 1979 1144 1980 1148
rect 2714 1145 2715 1149
rect 2719 1145 2720 1149
rect 2714 1144 2720 1145
rect 3018 1149 3024 1150
rect 3018 1145 3019 1149
rect 3023 1145 3024 1149
rect 3018 1144 3024 1145
rect 3330 1149 3336 1150
rect 3330 1145 3331 1149
rect 3335 1145 3336 1149
rect 3330 1144 3336 1145
rect 3650 1149 3656 1150
rect 3650 1145 3651 1149
rect 3655 1145 3656 1149
rect 3650 1144 3656 1145
rect 3798 1148 3804 1149
rect 3798 1144 3799 1148
rect 3803 1144 3804 1148
rect 1974 1143 1980 1144
rect 3798 1143 3804 1144
rect 110 1132 116 1133
rect 1934 1132 1940 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 146 1131 152 1132
rect 146 1127 147 1131
rect 151 1127 152 1131
rect 146 1126 152 1127
rect 322 1131 328 1132
rect 322 1127 323 1131
rect 327 1127 328 1131
rect 322 1126 328 1127
rect 498 1131 504 1132
rect 498 1127 499 1131
rect 503 1127 504 1131
rect 498 1126 504 1127
rect 674 1131 680 1132
rect 674 1127 675 1131
rect 679 1127 680 1131
rect 674 1126 680 1127
rect 850 1131 856 1132
rect 850 1127 851 1131
rect 855 1127 856 1131
rect 850 1126 856 1127
rect 1018 1131 1024 1132
rect 1018 1127 1019 1131
rect 1023 1127 1024 1131
rect 1018 1126 1024 1127
rect 1178 1131 1184 1132
rect 1178 1127 1179 1131
rect 1183 1127 1184 1131
rect 1178 1126 1184 1127
rect 1330 1131 1336 1132
rect 1330 1127 1331 1131
rect 1335 1127 1336 1131
rect 1330 1126 1336 1127
rect 1482 1131 1488 1132
rect 1482 1127 1483 1131
rect 1487 1127 1488 1131
rect 1482 1126 1488 1127
rect 1642 1131 1648 1132
rect 1642 1127 1643 1131
rect 1647 1127 1648 1131
rect 1642 1126 1648 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1786 1126 1792 1127
rect 174 1116 180 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 174 1112 175 1116
rect 179 1112 180 1116
rect 174 1111 180 1112
rect 350 1116 356 1117
rect 350 1112 351 1116
rect 355 1112 356 1116
rect 350 1111 356 1112
rect 526 1116 532 1117
rect 526 1112 527 1116
rect 531 1112 532 1116
rect 526 1111 532 1112
rect 702 1116 708 1117
rect 702 1112 703 1116
rect 707 1112 708 1116
rect 702 1111 708 1112
rect 878 1116 884 1117
rect 878 1112 879 1116
rect 883 1112 884 1116
rect 878 1111 884 1112
rect 1046 1116 1052 1117
rect 1046 1112 1047 1116
rect 1051 1112 1052 1116
rect 1046 1111 1052 1112
rect 1206 1116 1212 1117
rect 1206 1112 1207 1116
rect 1211 1112 1212 1116
rect 1206 1111 1212 1112
rect 1358 1116 1364 1117
rect 1358 1112 1359 1116
rect 1363 1112 1364 1116
rect 1358 1111 1364 1112
rect 1510 1116 1516 1117
rect 1510 1112 1511 1116
rect 1515 1112 1516 1116
rect 1510 1111 1516 1112
rect 1670 1116 1676 1117
rect 1670 1112 1671 1116
rect 1675 1112 1676 1116
rect 1670 1111 1676 1112
rect 1814 1116 1820 1117
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 110 1110 116 1111
rect 1934 1110 1940 1111
rect 3838 1104 3844 1105
rect 5662 1104 5668 1105
rect 3838 1100 3839 1104
rect 3843 1100 3844 1104
rect 3838 1099 3844 1100
rect 4810 1103 4816 1104
rect 4810 1099 4811 1103
rect 4815 1099 4816 1103
rect 4810 1098 4816 1099
rect 4946 1103 4952 1104
rect 4946 1099 4947 1103
rect 4951 1099 4952 1103
rect 4946 1098 4952 1099
rect 5082 1103 5088 1104
rect 5082 1099 5083 1103
rect 5087 1099 5088 1103
rect 5082 1098 5088 1099
rect 5226 1103 5232 1104
rect 5226 1099 5227 1103
rect 5231 1099 5232 1103
rect 5226 1098 5232 1099
rect 5378 1103 5384 1104
rect 5378 1099 5379 1103
rect 5383 1099 5384 1103
rect 5378 1098 5384 1099
rect 5514 1103 5520 1104
rect 5514 1099 5515 1103
rect 5519 1099 5520 1103
rect 5662 1100 5663 1104
rect 5667 1100 5668 1104
rect 5662 1099 5668 1100
rect 5514 1098 5520 1099
rect 4838 1088 4844 1089
rect 3838 1087 3844 1088
rect 3838 1083 3839 1087
rect 3843 1083 3844 1087
rect 4838 1084 4839 1088
rect 4843 1084 4844 1088
rect 4838 1083 4844 1084
rect 4974 1088 4980 1089
rect 4974 1084 4975 1088
rect 4979 1084 4980 1088
rect 4974 1083 4980 1084
rect 5110 1088 5116 1089
rect 5110 1084 5111 1088
rect 5115 1084 5116 1088
rect 5110 1083 5116 1084
rect 5254 1088 5260 1089
rect 5254 1084 5255 1088
rect 5259 1084 5260 1088
rect 5254 1083 5260 1084
rect 5406 1088 5412 1089
rect 5406 1084 5407 1088
rect 5411 1084 5412 1088
rect 5406 1083 5412 1084
rect 5542 1088 5548 1089
rect 5542 1084 5543 1088
rect 5547 1084 5548 1088
rect 5542 1083 5548 1084
rect 5662 1087 5668 1088
rect 5662 1083 5663 1087
rect 5667 1083 5668 1087
rect 3838 1082 3844 1083
rect 5662 1082 5668 1083
rect 110 1037 116 1038
rect 1934 1037 1940 1038
rect 110 1033 111 1037
rect 115 1033 116 1037
rect 110 1032 116 1033
rect 158 1036 164 1037
rect 158 1032 159 1036
rect 163 1032 164 1036
rect 158 1031 164 1032
rect 446 1036 452 1037
rect 446 1032 447 1036
rect 451 1032 452 1036
rect 446 1031 452 1032
rect 774 1036 780 1037
rect 774 1032 775 1036
rect 779 1032 780 1036
rect 774 1031 780 1032
rect 1110 1036 1116 1037
rect 1110 1032 1111 1036
rect 1115 1032 1116 1036
rect 1110 1031 1116 1032
rect 1454 1036 1460 1037
rect 1454 1032 1455 1036
rect 1459 1032 1460 1036
rect 1454 1031 1460 1032
rect 1806 1036 1812 1037
rect 1806 1032 1807 1036
rect 1811 1032 1812 1036
rect 1934 1033 1935 1037
rect 1939 1033 1940 1037
rect 1934 1032 1940 1033
rect 1806 1031 1812 1032
rect 3838 1025 3844 1026
rect 5662 1025 5668 1026
rect 130 1021 136 1022
rect 110 1020 116 1021
rect 110 1016 111 1020
rect 115 1016 116 1020
rect 130 1017 131 1021
rect 135 1017 136 1021
rect 130 1016 136 1017
rect 418 1021 424 1022
rect 418 1017 419 1021
rect 423 1017 424 1021
rect 418 1016 424 1017
rect 746 1021 752 1022
rect 746 1017 747 1021
rect 751 1017 752 1021
rect 746 1016 752 1017
rect 1082 1021 1088 1022
rect 1082 1017 1083 1021
rect 1087 1017 1088 1021
rect 1082 1016 1088 1017
rect 1426 1021 1432 1022
rect 1426 1017 1427 1021
rect 1431 1017 1432 1021
rect 1426 1016 1432 1017
rect 1778 1021 1784 1022
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 1778 1017 1779 1021
rect 1783 1017 1784 1021
rect 1778 1016 1784 1017
rect 1934 1020 1940 1021
rect 3838 1020 3844 1021
rect 4806 1024 4812 1025
rect 4806 1020 4807 1024
rect 4811 1020 4812 1024
rect 1934 1016 1935 1020
rect 1939 1016 1940 1020
rect 4806 1019 4812 1020
rect 4942 1024 4948 1025
rect 4942 1020 4943 1024
rect 4947 1020 4948 1024
rect 4942 1019 4948 1020
rect 5078 1024 5084 1025
rect 5078 1020 5079 1024
rect 5083 1020 5084 1024
rect 5078 1019 5084 1020
rect 5214 1024 5220 1025
rect 5214 1020 5215 1024
rect 5219 1020 5220 1024
rect 5214 1019 5220 1020
rect 5350 1024 5356 1025
rect 5350 1020 5351 1024
rect 5355 1020 5356 1024
rect 5350 1019 5356 1020
rect 5486 1024 5492 1025
rect 5486 1020 5487 1024
rect 5491 1020 5492 1024
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5486 1019 5492 1020
rect 110 1015 116 1016
rect 1934 1015 1940 1016
rect 1974 1016 1980 1017
rect 3798 1016 3804 1017
rect 1974 1012 1975 1016
rect 1979 1012 1980 1016
rect 1974 1011 1980 1012
rect 2242 1015 2248 1016
rect 2242 1011 2243 1015
rect 2247 1011 2248 1015
rect 2242 1010 2248 1011
rect 2378 1015 2384 1016
rect 2378 1011 2379 1015
rect 2383 1011 2384 1015
rect 2378 1010 2384 1011
rect 2522 1015 2528 1016
rect 2522 1011 2523 1015
rect 2527 1011 2528 1015
rect 2522 1010 2528 1011
rect 2674 1015 2680 1016
rect 2674 1011 2675 1015
rect 2679 1011 2680 1015
rect 2674 1010 2680 1011
rect 2826 1015 2832 1016
rect 2826 1011 2827 1015
rect 2831 1011 2832 1015
rect 2826 1010 2832 1011
rect 2986 1015 2992 1016
rect 2986 1011 2987 1015
rect 2991 1011 2992 1015
rect 2986 1010 2992 1011
rect 3154 1015 3160 1016
rect 3154 1011 3155 1015
rect 3159 1011 3160 1015
rect 3154 1010 3160 1011
rect 3322 1015 3328 1016
rect 3322 1011 3323 1015
rect 3327 1011 3328 1015
rect 3322 1010 3328 1011
rect 3498 1015 3504 1016
rect 3498 1011 3499 1015
rect 3503 1011 3504 1015
rect 3498 1010 3504 1011
rect 3650 1015 3656 1016
rect 3650 1011 3651 1015
rect 3655 1011 3656 1015
rect 3798 1012 3799 1016
rect 3803 1012 3804 1016
rect 3798 1011 3804 1012
rect 3650 1010 3656 1011
rect 4778 1009 4784 1010
rect 3838 1008 3844 1009
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 4778 1005 4779 1009
rect 4783 1005 4784 1009
rect 4778 1004 4784 1005
rect 4914 1009 4920 1010
rect 4914 1005 4915 1009
rect 4919 1005 4920 1009
rect 4914 1004 4920 1005
rect 5050 1009 5056 1010
rect 5050 1005 5051 1009
rect 5055 1005 5056 1009
rect 5050 1004 5056 1005
rect 5186 1009 5192 1010
rect 5186 1005 5187 1009
rect 5191 1005 5192 1009
rect 5186 1004 5192 1005
rect 5322 1009 5328 1010
rect 5322 1005 5323 1009
rect 5327 1005 5328 1009
rect 5322 1004 5328 1005
rect 5458 1009 5464 1010
rect 5458 1005 5459 1009
rect 5463 1005 5464 1009
rect 5458 1004 5464 1005
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 3838 1003 3844 1004
rect 5662 1003 5668 1004
rect 2270 1000 2276 1001
rect 1974 999 1980 1000
rect 1974 995 1975 999
rect 1979 995 1980 999
rect 2270 996 2271 1000
rect 2275 996 2276 1000
rect 2270 995 2276 996
rect 2406 1000 2412 1001
rect 2406 996 2407 1000
rect 2411 996 2412 1000
rect 2406 995 2412 996
rect 2550 1000 2556 1001
rect 2550 996 2551 1000
rect 2555 996 2556 1000
rect 2550 995 2556 996
rect 2702 1000 2708 1001
rect 2702 996 2703 1000
rect 2707 996 2708 1000
rect 2702 995 2708 996
rect 2854 1000 2860 1001
rect 2854 996 2855 1000
rect 2859 996 2860 1000
rect 2854 995 2860 996
rect 3014 1000 3020 1001
rect 3014 996 3015 1000
rect 3019 996 3020 1000
rect 3014 995 3020 996
rect 3182 1000 3188 1001
rect 3182 996 3183 1000
rect 3187 996 3188 1000
rect 3182 995 3188 996
rect 3350 1000 3356 1001
rect 3350 996 3351 1000
rect 3355 996 3356 1000
rect 3350 995 3356 996
rect 3526 1000 3532 1001
rect 3526 996 3527 1000
rect 3531 996 3532 1000
rect 3526 995 3532 996
rect 3678 1000 3684 1001
rect 3678 996 3679 1000
rect 3683 996 3684 1000
rect 3678 995 3684 996
rect 3798 999 3804 1000
rect 3798 995 3799 999
rect 3803 995 3804 999
rect 1974 994 1980 995
rect 3798 994 3804 995
rect 1974 937 1980 938
rect 3798 937 3804 938
rect 1974 933 1975 937
rect 1979 933 1980 937
rect 1974 932 1980 933
rect 2278 936 2284 937
rect 2278 932 2279 936
rect 2283 932 2284 936
rect 2278 931 2284 932
rect 2494 936 2500 937
rect 2494 932 2495 936
rect 2499 932 2500 936
rect 2494 931 2500 932
rect 2710 936 2716 937
rect 2710 932 2711 936
rect 2715 932 2716 936
rect 2710 931 2716 932
rect 2910 936 2916 937
rect 2910 932 2911 936
rect 2915 932 2916 936
rect 2910 931 2916 932
rect 3102 936 3108 937
rect 3102 932 3103 936
rect 3107 932 3108 936
rect 3102 931 3108 932
rect 3294 936 3300 937
rect 3294 932 3295 936
rect 3299 932 3300 936
rect 3294 931 3300 932
rect 3478 936 3484 937
rect 3478 932 3479 936
rect 3483 932 3484 936
rect 3478 931 3484 932
rect 3670 936 3676 937
rect 3670 932 3671 936
rect 3675 932 3676 936
rect 3798 933 3799 937
rect 3803 933 3804 937
rect 3798 932 3804 933
rect 3670 931 3676 932
rect 2250 921 2256 922
rect 1974 920 1980 921
rect 1974 916 1975 920
rect 1979 916 1980 920
rect 2250 917 2251 921
rect 2255 917 2256 921
rect 2250 916 2256 917
rect 2466 921 2472 922
rect 2466 917 2467 921
rect 2471 917 2472 921
rect 2466 916 2472 917
rect 2682 921 2688 922
rect 2682 917 2683 921
rect 2687 917 2688 921
rect 2682 916 2688 917
rect 2882 921 2888 922
rect 2882 917 2883 921
rect 2887 917 2888 921
rect 2882 916 2888 917
rect 3074 921 3080 922
rect 3074 917 3075 921
rect 3079 917 3080 921
rect 3074 916 3080 917
rect 3266 921 3272 922
rect 3266 917 3267 921
rect 3271 917 3272 921
rect 3266 916 3272 917
rect 3450 921 3456 922
rect 3450 917 3451 921
rect 3455 917 3456 921
rect 3450 916 3456 917
rect 3642 921 3648 922
rect 3642 917 3643 921
rect 3647 917 3648 921
rect 3642 916 3648 917
rect 3798 920 3804 921
rect 3798 916 3799 920
rect 3803 916 3804 920
rect 1974 915 1980 916
rect 3798 915 3804 916
rect 110 884 116 885
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 130 883 136 884
rect 130 879 131 883
rect 135 879 136 883
rect 130 878 136 879
rect 338 883 344 884
rect 338 879 339 883
rect 343 879 344 883
rect 338 878 344 879
rect 594 883 600 884
rect 594 879 595 883
rect 599 879 600 883
rect 594 878 600 879
rect 874 883 880 884
rect 874 879 875 883
rect 879 879 880 883
rect 874 878 880 879
rect 1178 883 1184 884
rect 1178 879 1179 883
rect 1183 879 1184 883
rect 1178 878 1184 879
rect 1490 883 1496 884
rect 1490 879 1491 883
rect 1495 879 1496 883
rect 1490 878 1496 879
rect 1786 883 1792 884
rect 1786 879 1787 883
rect 1791 879 1792 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 1786 878 1792 879
rect 3838 872 3844 873
rect 5662 872 5668 873
rect 158 868 164 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 158 864 159 868
rect 163 864 164 868
rect 158 863 164 864
rect 366 868 372 869
rect 366 864 367 868
rect 371 864 372 868
rect 366 863 372 864
rect 622 868 628 869
rect 622 864 623 868
rect 627 864 628 868
rect 622 863 628 864
rect 902 868 908 869
rect 902 864 903 868
rect 907 864 908 868
rect 902 863 908 864
rect 1206 868 1212 869
rect 1206 864 1207 868
rect 1211 864 1212 868
rect 1206 863 1212 864
rect 1518 868 1524 869
rect 1518 864 1519 868
rect 1523 864 1524 868
rect 1518 863 1524 864
rect 1814 868 1820 869
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 1814 864 1815 868
rect 1819 864 1820 868
rect 1814 863 1820 864
rect 1934 867 1940 868
rect 3838 867 3844 868
rect 4354 871 4360 872
rect 4354 867 4355 871
rect 4359 867 4360 871
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 4354 866 4360 867
rect 4570 871 4576 872
rect 4570 867 4571 871
rect 4575 867 4576 871
rect 4570 866 4576 867
rect 4802 871 4808 872
rect 4802 867 4803 871
rect 4807 867 4808 871
rect 4802 866 4808 867
rect 5042 871 5048 872
rect 5042 867 5043 871
rect 5047 867 5048 871
rect 5042 866 5048 867
rect 5290 871 5296 872
rect 5290 867 5291 871
rect 5295 867 5296 871
rect 5290 866 5296 867
rect 5514 871 5520 872
rect 5514 867 5515 871
rect 5519 867 5520 871
rect 5662 868 5663 872
rect 5667 868 5668 872
rect 5662 867 5668 868
rect 5514 866 5520 867
rect 110 862 116 863
rect 1934 862 1940 863
rect 4382 856 4388 857
rect 3838 855 3844 856
rect 3838 851 3839 855
rect 3843 851 3844 855
rect 4382 852 4383 856
rect 4387 852 4388 856
rect 4382 851 4388 852
rect 4598 856 4604 857
rect 4598 852 4599 856
rect 4603 852 4604 856
rect 4598 851 4604 852
rect 4830 856 4836 857
rect 4830 852 4831 856
rect 4835 852 4836 856
rect 4830 851 4836 852
rect 5070 856 5076 857
rect 5070 852 5071 856
rect 5075 852 5076 856
rect 5070 851 5076 852
rect 5318 856 5324 857
rect 5318 852 5319 856
rect 5323 852 5324 856
rect 5318 851 5324 852
rect 5542 856 5548 857
rect 5542 852 5543 856
rect 5547 852 5548 856
rect 5542 851 5548 852
rect 5662 855 5668 856
rect 5662 851 5663 855
rect 5667 851 5668 855
rect 3838 850 3844 851
rect 5662 850 5668 851
rect 110 797 116 798
rect 1934 797 1940 798
rect 110 793 111 797
rect 115 793 116 797
rect 110 792 116 793
rect 158 796 164 797
rect 158 792 159 796
rect 163 792 164 796
rect 158 791 164 792
rect 382 796 388 797
rect 382 792 383 796
rect 387 792 388 796
rect 382 791 388 792
rect 630 796 636 797
rect 630 792 631 796
rect 635 792 636 796
rect 630 791 636 792
rect 886 796 892 797
rect 886 792 887 796
rect 891 792 892 796
rect 886 791 892 792
rect 1142 796 1148 797
rect 1142 792 1143 796
rect 1147 792 1148 796
rect 1934 793 1935 797
rect 1939 793 1940 797
rect 1934 792 1940 793
rect 3838 793 3844 794
rect 5662 793 5668 794
rect 1142 791 1148 792
rect 3838 789 3839 793
rect 3843 789 3844 793
rect 3838 788 3844 789
rect 3958 792 3964 793
rect 3958 788 3959 792
rect 3963 788 3964 792
rect 3958 787 3964 788
rect 4206 792 4212 793
rect 4206 788 4207 792
rect 4211 788 4212 792
rect 4206 787 4212 788
rect 4494 792 4500 793
rect 4494 788 4495 792
rect 4499 788 4500 792
rect 4494 787 4500 788
rect 4814 792 4820 793
rect 4814 788 4815 792
rect 4819 788 4820 792
rect 4814 787 4820 788
rect 5150 792 5156 793
rect 5150 788 5151 792
rect 5155 788 5156 792
rect 5150 787 5156 788
rect 5486 792 5492 793
rect 5486 788 5487 792
rect 5491 788 5492 792
rect 5662 789 5663 793
rect 5667 789 5668 793
rect 5662 788 5668 789
rect 5486 787 5492 788
rect 1974 784 1980 785
rect 3798 784 3804 785
rect 130 781 136 782
rect 110 780 116 781
rect 110 776 111 780
rect 115 776 116 780
rect 130 777 131 781
rect 135 777 136 781
rect 130 776 136 777
rect 354 781 360 782
rect 354 777 355 781
rect 359 777 360 781
rect 354 776 360 777
rect 602 781 608 782
rect 602 777 603 781
rect 607 777 608 781
rect 602 776 608 777
rect 858 781 864 782
rect 858 777 859 781
rect 863 777 864 781
rect 858 776 864 777
rect 1114 781 1120 782
rect 1114 777 1115 781
rect 1119 777 1120 781
rect 1114 776 1120 777
rect 1934 780 1940 781
rect 1934 776 1935 780
rect 1939 776 1940 780
rect 1974 780 1975 784
rect 1979 780 1980 784
rect 1974 779 1980 780
rect 1994 783 2000 784
rect 1994 779 1995 783
rect 1999 779 2000 783
rect 1994 778 2000 779
rect 2130 783 2136 784
rect 2130 779 2131 783
rect 2135 779 2136 783
rect 2130 778 2136 779
rect 2282 783 2288 784
rect 2282 779 2283 783
rect 2287 779 2288 783
rect 2282 778 2288 779
rect 2442 783 2448 784
rect 2442 779 2443 783
rect 2447 779 2448 783
rect 2442 778 2448 779
rect 2602 783 2608 784
rect 2602 779 2603 783
rect 2607 779 2608 783
rect 2602 778 2608 779
rect 2762 783 2768 784
rect 2762 779 2763 783
rect 2767 779 2768 783
rect 2762 778 2768 779
rect 2922 783 2928 784
rect 2922 779 2923 783
rect 2927 779 2928 783
rect 2922 778 2928 779
rect 3082 783 3088 784
rect 3082 779 3083 783
rect 3087 779 3088 783
rect 3082 778 3088 779
rect 3242 783 3248 784
rect 3242 779 3243 783
rect 3247 779 3248 783
rect 3242 778 3248 779
rect 3402 783 3408 784
rect 3402 779 3403 783
rect 3407 779 3408 783
rect 3798 780 3799 784
rect 3803 780 3804 784
rect 3798 779 3804 780
rect 3402 778 3408 779
rect 3930 777 3936 778
rect 110 775 116 776
rect 1934 775 1940 776
rect 3838 776 3844 777
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3930 773 3931 777
rect 3935 773 3936 777
rect 3930 772 3936 773
rect 4178 777 4184 778
rect 4178 773 4179 777
rect 4183 773 4184 777
rect 4178 772 4184 773
rect 4466 777 4472 778
rect 4466 773 4467 777
rect 4471 773 4472 777
rect 4466 772 4472 773
rect 4786 777 4792 778
rect 4786 773 4787 777
rect 4791 773 4792 777
rect 4786 772 4792 773
rect 5122 777 5128 778
rect 5122 773 5123 777
rect 5127 773 5128 777
rect 5122 772 5128 773
rect 5458 777 5464 778
rect 5458 773 5459 777
rect 5463 773 5464 777
rect 5458 772 5464 773
rect 5662 776 5668 777
rect 5662 772 5663 776
rect 5667 772 5668 776
rect 3838 771 3844 772
rect 5662 771 5668 772
rect 2022 768 2028 769
rect 1974 767 1980 768
rect 1974 763 1975 767
rect 1979 763 1980 767
rect 2022 764 2023 768
rect 2027 764 2028 768
rect 2022 763 2028 764
rect 2158 768 2164 769
rect 2158 764 2159 768
rect 2163 764 2164 768
rect 2158 763 2164 764
rect 2310 768 2316 769
rect 2310 764 2311 768
rect 2315 764 2316 768
rect 2310 763 2316 764
rect 2470 768 2476 769
rect 2470 764 2471 768
rect 2475 764 2476 768
rect 2470 763 2476 764
rect 2630 768 2636 769
rect 2630 764 2631 768
rect 2635 764 2636 768
rect 2630 763 2636 764
rect 2790 768 2796 769
rect 2790 764 2791 768
rect 2795 764 2796 768
rect 2790 763 2796 764
rect 2950 768 2956 769
rect 2950 764 2951 768
rect 2955 764 2956 768
rect 2950 763 2956 764
rect 3110 768 3116 769
rect 3110 764 3111 768
rect 3115 764 3116 768
rect 3110 763 3116 764
rect 3270 768 3276 769
rect 3270 764 3271 768
rect 3275 764 3276 768
rect 3270 763 3276 764
rect 3430 768 3436 769
rect 3430 764 3431 768
rect 3435 764 3436 768
rect 3430 763 3436 764
rect 3798 767 3804 768
rect 3798 763 3799 767
rect 3803 763 3804 767
rect 1974 762 1980 763
rect 3798 762 3804 763
rect 1974 709 1980 710
rect 3798 709 3804 710
rect 1974 705 1975 709
rect 1979 705 1980 709
rect 1974 704 1980 705
rect 2182 708 2188 709
rect 2182 704 2183 708
rect 2187 704 2188 708
rect 2182 703 2188 704
rect 2438 708 2444 709
rect 2438 704 2439 708
rect 2443 704 2444 708
rect 2438 703 2444 704
rect 2678 708 2684 709
rect 2678 704 2679 708
rect 2683 704 2684 708
rect 2678 703 2684 704
rect 2902 708 2908 709
rect 2902 704 2903 708
rect 2907 704 2908 708
rect 2902 703 2908 704
rect 3110 708 3116 709
rect 3110 704 3111 708
rect 3115 704 3116 708
rect 3110 703 3116 704
rect 3310 708 3316 709
rect 3310 704 3311 708
rect 3315 704 3316 708
rect 3310 703 3316 704
rect 3502 708 3508 709
rect 3502 704 3503 708
rect 3507 704 3508 708
rect 3502 703 3508 704
rect 3678 708 3684 709
rect 3678 704 3679 708
rect 3683 704 3684 708
rect 3798 705 3799 709
rect 3803 705 3804 709
rect 3798 704 3804 705
rect 3678 703 3684 704
rect 2154 693 2160 694
rect 1974 692 1980 693
rect 1974 688 1975 692
rect 1979 688 1980 692
rect 2154 689 2155 693
rect 2159 689 2160 693
rect 2154 688 2160 689
rect 2410 693 2416 694
rect 2410 689 2411 693
rect 2415 689 2416 693
rect 2410 688 2416 689
rect 2650 693 2656 694
rect 2650 689 2651 693
rect 2655 689 2656 693
rect 2650 688 2656 689
rect 2874 693 2880 694
rect 2874 689 2875 693
rect 2879 689 2880 693
rect 2874 688 2880 689
rect 3082 693 3088 694
rect 3082 689 3083 693
rect 3087 689 3088 693
rect 3082 688 3088 689
rect 3282 693 3288 694
rect 3282 689 3283 693
rect 3287 689 3288 693
rect 3282 688 3288 689
rect 3474 693 3480 694
rect 3474 689 3475 693
rect 3479 689 3480 693
rect 3474 688 3480 689
rect 3650 693 3656 694
rect 3650 689 3651 693
rect 3655 689 3656 693
rect 3650 688 3656 689
rect 3798 692 3804 693
rect 3798 688 3799 692
rect 3803 688 3804 692
rect 1974 687 1980 688
rect 3798 687 3804 688
rect 110 648 116 649
rect 1934 648 1940 649
rect 110 644 111 648
rect 115 644 116 648
rect 110 643 116 644
rect 698 647 704 648
rect 698 643 699 647
rect 703 643 704 647
rect 698 642 704 643
rect 834 647 840 648
rect 834 643 835 647
rect 839 643 840 647
rect 834 642 840 643
rect 970 647 976 648
rect 970 643 971 647
rect 975 643 976 647
rect 970 642 976 643
rect 1106 647 1112 648
rect 1106 643 1107 647
rect 1111 643 1112 647
rect 1106 642 1112 643
rect 1242 647 1248 648
rect 1242 643 1243 647
rect 1247 643 1248 647
rect 1242 642 1248 643
rect 1378 647 1384 648
rect 1378 643 1379 647
rect 1383 643 1384 647
rect 1378 642 1384 643
rect 1514 647 1520 648
rect 1514 643 1515 647
rect 1519 643 1520 647
rect 1514 642 1520 643
rect 1650 647 1656 648
rect 1650 643 1651 647
rect 1655 643 1656 647
rect 1650 642 1656 643
rect 1786 647 1792 648
rect 1786 643 1787 647
rect 1791 643 1792 647
rect 1934 644 1935 648
rect 1939 644 1940 648
rect 1934 643 1940 644
rect 1786 642 1792 643
rect 726 632 732 633
rect 110 631 116 632
rect 110 627 111 631
rect 115 627 116 631
rect 726 628 727 632
rect 731 628 732 632
rect 726 627 732 628
rect 862 632 868 633
rect 862 628 863 632
rect 867 628 868 632
rect 862 627 868 628
rect 998 632 1004 633
rect 998 628 999 632
rect 1003 628 1004 632
rect 998 627 1004 628
rect 1134 632 1140 633
rect 1134 628 1135 632
rect 1139 628 1140 632
rect 1134 627 1140 628
rect 1270 632 1276 633
rect 1270 628 1271 632
rect 1275 628 1276 632
rect 1270 627 1276 628
rect 1406 632 1412 633
rect 1406 628 1407 632
rect 1411 628 1412 632
rect 1406 627 1412 628
rect 1542 632 1548 633
rect 1542 628 1543 632
rect 1547 628 1548 632
rect 1542 627 1548 628
rect 1678 632 1684 633
rect 1678 628 1679 632
rect 1683 628 1684 632
rect 1678 627 1684 628
rect 1814 632 1820 633
rect 3838 632 3844 633
rect 5662 632 5668 633
rect 1814 628 1815 632
rect 1819 628 1820 632
rect 1814 627 1820 628
rect 1934 631 1940 632
rect 1934 627 1935 631
rect 1939 627 1940 631
rect 3838 628 3839 632
rect 3843 628 3844 632
rect 3838 627 3844 628
rect 3858 631 3864 632
rect 3858 627 3859 631
rect 3863 627 3864 631
rect 110 626 116 627
rect 1934 626 1940 627
rect 3858 626 3864 627
rect 3994 631 4000 632
rect 3994 627 3995 631
rect 3999 627 4000 631
rect 3994 626 4000 627
rect 4146 631 4152 632
rect 4146 627 4147 631
rect 4151 627 4152 631
rect 4146 626 4152 627
rect 4354 631 4360 632
rect 4354 627 4355 631
rect 4359 627 4360 631
rect 4354 626 4360 627
rect 4594 631 4600 632
rect 4594 627 4595 631
rect 4599 627 4600 631
rect 4594 626 4600 627
rect 4866 631 4872 632
rect 4866 627 4867 631
rect 4871 627 4872 631
rect 4866 626 4872 627
rect 5162 631 5168 632
rect 5162 627 5163 631
rect 5167 627 5168 631
rect 5162 626 5168 627
rect 5458 631 5464 632
rect 5458 627 5459 631
rect 5463 627 5464 631
rect 5662 628 5663 632
rect 5667 628 5668 632
rect 5662 627 5668 628
rect 5458 626 5464 627
rect 3886 616 3892 617
rect 3838 615 3844 616
rect 3838 611 3839 615
rect 3843 611 3844 615
rect 3886 612 3887 616
rect 3891 612 3892 616
rect 3886 611 3892 612
rect 4022 616 4028 617
rect 4022 612 4023 616
rect 4027 612 4028 616
rect 4022 611 4028 612
rect 4174 616 4180 617
rect 4174 612 4175 616
rect 4179 612 4180 616
rect 4174 611 4180 612
rect 4382 616 4388 617
rect 4382 612 4383 616
rect 4387 612 4388 616
rect 4382 611 4388 612
rect 4622 616 4628 617
rect 4622 612 4623 616
rect 4627 612 4628 616
rect 4622 611 4628 612
rect 4894 616 4900 617
rect 4894 612 4895 616
rect 4899 612 4900 616
rect 4894 611 4900 612
rect 5190 616 5196 617
rect 5190 612 5191 616
rect 5195 612 5196 616
rect 5190 611 5196 612
rect 5486 616 5492 617
rect 5486 612 5487 616
rect 5491 612 5492 616
rect 5486 611 5492 612
rect 5662 615 5668 616
rect 5662 611 5663 615
rect 5667 611 5668 615
rect 3838 610 3844 611
rect 5662 610 5668 611
rect 110 573 116 574
rect 1934 573 1940 574
rect 110 569 111 573
rect 115 569 116 573
rect 110 568 116 569
rect 158 572 164 573
rect 158 568 159 572
rect 163 568 164 572
rect 158 567 164 568
rect 374 572 380 573
rect 374 568 375 572
rect 379 568 380 572
rect 374 567 380 568
rect 598 572 604 573
rect 598 568 599 572
rect 603 568 604 572
rect 598 567 604 568
rect 806 572 812 573
rect 806 568 807 572
rect 811 568 812 572
rect 806 567 812 568
rect 998 572 1004 573
rect 998 568 999 572
rect 1003 568 1004 572
rect 998 567 1004 568
rect 1174 572 1180 573
rect 1174 568 1175 572
rect 1179 568 1180 572
rect 1174 567 1180 568
rect 1342 572 1348 573
rect 1342 568 1343 572
rect 1347 568 1348 572
rect 1342 567 1348 568
rect 1510 572 1516 573
rect 1510 568 1511 572
rect 1515 568 1516 572
rect 1510 567 1516 568
rect 1670 572 1676 573
rect 1670 568 1671 572
rect 1675 568 1676 572
rect 1670 567 1676 568
rect 1814 572 1820 573
rect 1814 568 1815 572
rect 1819 568 1820 572
rect 1934 569 1935 573
rect 1939 569 1940 573
rect 1934 568 1940 569
rect 1814 567 1820 568
rect 130 557 136 558
rect 110 556 116 557
rect 110 552 111 556
rect 115 552 116 556
rect 130 553 131 557
rect 135 553 136 557
rect 130 552 136 553
rect 346 557 352 558
rect 346 553 347 557
rect 351 553 352 557
rect 346 552 352 553
rect 570 557 576 558
rect 570 553 571 557
rect 575 553 576 557
rect 570 552 576 553
rect 778 557 784 558
rect 778 553 779 557
rect 783 553 784 557
rect 778 552 784 553
rect 970 557 976 558
rect 970 553 971 557
rect 975 553 976 557
rect 970 552 976 553
rect 1146 557 1152 558
rect 1146 553 1147 557
rect 1151 553 1152 557
rect 1146 552 1152 553
rect 1314 557 1320 558
rect 1314 553 1315 557
rect 1319 553 1320 557
rect 1314 552 1320 553
rect 1482 557 1488 558
rect 1482 553 1483 557
rect 1487 553 1488 557
rect 1482 552 1488 553
rect 1642 557 1648 558
rect 1642 553 1643 557
rect 1647 553 1648 557
rect 1642 552 1648 553
rect 1786 557 1792 558
rect 3838 557 3844 558
rect 5662 557 5668 558
rect 1786 553 1787 557
rect 1791 553 1792 557
rect 1786 552 1792 553
rect 1934 556 1940 557
rect 1934 552 1935 556
rect 1939 552 1940 556
rect 3838 553 3839 557
rect 3843 553 3844 557
rect 3838 552 3844 553
rect 3886 556 3892 557
rect 3886 552 3887 556
rect 3891 552 3892 556
rect 110 551 116 552
rect 1934 551 1940 552
rect 3886 551 3892 552
rect 4022 556 4028 557
rect 4022 552 4023 556
rect 4027 552 4028 556
rect 4022 551 4028 552
rect 4158 556 4164 557
rect 4158 552 4159 556
rect 4163 552 4164 556
rect 4158 551 4164 552
rect 4294 556 4300 557
rect 4294 552 4295 556
rect 4299 552 4300 556
rect 4294 551 4300 552
rect 4430 556 4436 557
rect 4430 552 4431 556
rect 4435 552 4436 556
rect 4430 551 4436 552
rect 4566 556 4572 557
rect 4566 552 4567 556
rect 4571 552 4572 556
rect 4566 551 4572 552
rect 4710 556 4716 557
rect 4710 552 4711 556
rect 4715 552 4716 556
rect 4710 551 4716 552
rect 4878 556 4884 557
rect 4878 552 4879 556
rect 4883 552 4884 556
rect 4878 551 4884 552
rect 5062 556 5068 557
rect 5062 552 5063 556
rect 5067 552 5068 556
rect 5062 551 5068 552
rect 5254 556 5260 557
rect 5254 552 5255 556
rect 5259 552 5260 556
rect 5254 551 5260 552
rect 5446 556 5452 557
rect 5446 552 5447 556
rect 5451 552 5452 556
rect 5662 553 5663 557
rect 5667 553 5668 557
rect 5662 552 5668 553
rect 5446 551 5452 552
rect 3858 541 3864 542
rect 3838 540 3844 541
rect 3838 536 3839 540
rect 3843 536 3844 540
rect 3858 537 3859 541
rect 3863 537 3864 541
rect 3858 536 3864 537
rect 3994 541 4000 542
rect 3994 537 3995 541
rect 3999 537 4000 541
rect 3994 536 4000 537
rect 4130 541 4136 542
rect 4130 537 4131 541
rect 4135 537 4136 541
rect 4130 536 4136 537
rect 4266 541 4272 542
rect 4266 537 4267 541
rect 4271 537 4272 541
rect 4266 536 4272 537
rect 4402 541 4408 542
rect 4402 537 4403 541
rect 4407 537 4408 541
rect 4402 536 4408 537
rect 4538 541 4544 542
rect 4538 537 4539 541
rect 4543 537 4544 541
rect 4538 536 4544 537
rect 4682 541 4688 542
rect 4682 537 4683 541
rect 4687 537 4688 541
rect 4682 536 4688 537
rect 4850 541 4856 542
rect 4850 537 4851 541
rect 4855 537 4856 541
rect 4850 536 4856 537
rect 5034 541 5040 542
rect 5034 537 5035 541
rect 5039 537 5040 541
rect 5034 536 5040 537
rect 5226 541 5232 542
rect 5226 537 5227 541
rect 5231 537 5232 541
rect 5226 536 5232 537
rect 5418 541 5424 542
rect 5418 537 5419 541
rect 5423 537 5424 541
rect 5418 536 5424 537
rect 5662 540 5668 541
rect 5662 536 5663 540
rect 5667 536 5668 540
rect 3838 535 3844 536
rect 5662 535 5668 536
rect 110 424 116 425
rect 1934 424 1940 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 130 423 136 424
rect 130 419 131 423
rect 135 419 136 423
rect 130 418 136 419
rect 354 423 360 424
rect 354 419 355 423
rect 359 419 360 423
rect 354 418 360 419
rect 602 423 608 424
rect 602 419 603 423
rect 607 419 608 423
rect 602 418 608 419
rect 842 423 848 424
rect 842 419 843 423
rect 847 419 848 423
rect 842 418 848 419
rect 1082 423 1088 424
rect 1082 419 1083 423
rect 1087 419 1088 423
rect 1082 418 1088 419
rect 1322 423 1328 424
rect 1322 419 1323 423
rect 1327 419 1328 423
rect 1322 418 1328 419
rect 1562 423 1568 424
rect 1562 419 1563 423
rect 1567 419 1568 423
rect 1562 418 1568 419
rect 1786 423 1792 424
rect 1786 419 1787 423
rect 1791 419 1792 423
rect 1934 420 1935 424
rect 1939 420 1940 424
rect 1934 419 1940 420
rect 1786 418 1792 419
rect 158 408 164 409
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 158 404 159 408
rect 163 404 164 408
rect 158 403 164 404
rect 382 408 388 409
rect 382 404 383 408
rect 387 404 388 408
rect 382 403 388 404
rect 630 408 636 409
rect 630 404 631 408
rect 635 404 636 408
rect 630 403 636 404
rect 870 408 876 409
rect 870 404 871 408
rect 875 404 876 408
rect 870 403 876 404
rect 1110 408 1116 409
rect 1110 404 1111 408
rect 1115 404 1116 408
rect 1110 403 1116 404
rect 1350 408 1356 409
rect 1350 404 1351 408
rect 1355 404 1356 408
rect 1350 403 1356 404
rect 1590 408 1596 409
rect 1590 404 1591 408
rect 1595 404 1596 408
rect 1590 403 1596 404
rect 1814 408 1820 409
rect 3838 408 3844 409
rect 5662 408 5668 409
rect 1814 404 1815 408
rect 1819 404 1820 408
rect 1814 403 1820 404
rect 1934 407 1940 408
rect 1934 403 1935 407
rect 1939 403 1940 407
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 3858 407 3864 408
rect 3858 403 3859 407
rect 3863 403 3864 407
rect 110 402 116 403
rect 1934 402 1940 403
rect 3858 402 3864 403
rect 4114 407 4120 408
rect 4114 403 4115 407
rect 4119 403 4120 407
rect 4114 402 4120 403
rect 4394 407 4400 408
rect 4394 403 4395 407
rect 4399 403 4400 407
rect 4394 402 4400 403
rect 4674 407 4680 408
rect 4674 403 4675 407
rect 4679 403 4680 407
rect 4674 402 4680 403
rect 4946 407 4952 408
rect 4946 403 4947 407
rect 4951 403 4952 407
rect 4946 402 4952 403
rect 5226 407 5232 408
rect 5226 403 5227 407
rect 5231 403 5232 407
rect 5226 402 5232 403
rect 5506 407 5512 408
rect 5506 403 5507 407
rect 5511 403 5512 407
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5506 402 5512 403
rect 3886 392 3892 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 3886 388 3887 392
rect 3891 388 3892 392
rect 3886 387 3892 388
rect 4142 392 4148 393
rect 4142 388 4143 392
rect 4147 388 4148 392
rect 4142 387 4148 388
rect 4422 392 4428 393
rect 4422 388 4423 392
rect 4427 388 4428 392
rect 4422 387 4428 388
rect 4702 392 4708 393
rect 4702 388 4703 392
rect 4707 388 4708 392
rect 4702 387 4708 388
rect 4974 392 4980 393
rect 4974 388 4975 392
rect 4979 388 4980 392
rect 4974 387 4980 388
rect 5254 392 5260 393
rect 5254 388 5255 392
rect 5259 388 5260 392
rect 5254 387 5260 388
rect 5534 392 5540 393
rect 5534 388 5535 392
rect 5539 388 5540 392
rect 5534 387 5540 388
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 3838 386 3844 387
rect 5662 386 5668 387
rect 1974 384 1980 385
rect 3798 384 3804 385
rect 1974 380 1975 384
rect 1979 380 1980 384
rect 1974 379 1980 380
rect 1994 383 2000 384
rect 1994 379 1995 383
rect 1999 379 2000 383
rect 1994 378 2000 379
rect 2250 383 2256 384
rect 2250 379 2251 383
rect 2255 379 2256 383
rect 2250 378 2256 379
rect 2522 383 2528 384
rect 2522 379 2523 383
rect 2527 379 2528 383
rect 2522 378 2528 379
rect 2770 383 2776 384
rect 2770 379 2771 383
rect 2775 379 2776 383
rect 2770 378 2776 379
rect 3002 383 3008 384
rect 3002 379 3003 383
rect 3007 379 3008 383
rect 3002 378 3008 379
rect 3226 383 3232 384
rect 3226 379 3227 383
rect 3231 379 3232 383
rect 3226 378 3232 379
rect 3450 383 3456 384
rect 3450 379 3451 383
rect 3455 379 3456 383
rect 3450 378 3456 379
rect 3650 383 3656 384
rect 3650 379 3651 383
rect 3655 379 3656 383
rect 3798 380 3799 384
rect 3803 380 3804 384
rect 3798 379 3804 380
rect 3650 378 3656 379
rect 2022 368 2028 369
rect 1974 367 1980 368
rect 1974 363 1975 367
rect 1979 363 1980 367
rect 2022 364 2023 368
rect 2027 364 2028 368
rect 2022 363 2028 364
rect 2278 368 2284 369
rect 2278 364 2279 368
rect 2283 364 2284 368
rect 2278 363 2284 364
rect 2550 368 2556 369
rect 2550 364 2551 368
rect 2555 364 2556 368
rect 2550 363 2556 364
rect 2798 368 2804 369
rect 2798 364 2799 368
rect 2803 364 2804 368
rect 2798 363 2804 364
rect 3030 368 3036 369
rect 3030 364 3031 368
rect 3035 364 3036 368
rect 3030 363 3036 364
rect 3254 368 3260 369
rect 3254 364 3255 368
rect 3259 364 3260 368
rect 3254 363 3260 364
rect 3478 368 3484 369
rect 3478 364 3479 368
rect 3483 364 3484 368
rect 3478 363 3484 364
rect 3678 368 3684 369
rect 3678 364 3679 368
rect 3683 364 3684 368
rect 3678 363 3684 364
rect 3798 367 3804 368
rect 3798 363 3799 367
rect 3803 363 3804 367
rect 1974 362 1980 363
rect 3798 362 3804 363
rect 110 333 116 334
rect 1934 333 1940 334
rect 110 329 111 333
rect 115 329 116 333
rect 110 328 116 329
rect 158 332 164 333
rect 158 328 159 332
rect 163 328 164 332
rect 158 327 164 328
rect 302 332 308 333
rect 302 328 303 332
rect 307 328 308 332
rect 302 327 308 328
rect 478 332 484 333
rect 478 328 479 332
rect 483 328 484 332
rect 478 327 484 328
rect 654 332 660 333
rect 654 328 655 332
rect 659 328 660 332
rect 654 327 660 328
rect 830 332 836 333
rect 830 328 831 332
rect 835 328 836 332
rect 1934 329 1935 333
rect 1939 329 1940 333
rect 1934 328 1940 329
rect 830 327 836 328
rect 3838 325 3844 326
rect 5662 325 5668 326
rect 3838 321 3839 325
rect 3843 321 3844 325
rect 3838 320 3844 321
rect 4726 324 4732 325
rect 4726 320 4727 324
rect 4731 320 4732 324
rect 4726 319 4732 320
rect 4894 324 4900 325
rect 4894 320 4895 324
rect 4899 320 4900 324
rect 4894 319 4900 320
rect 5062 324 5068 325
rect 5062 320 5063 324
rect 5067 320 5068 324
rect 5062 319 5068 320
rect 5230 324 5236 325
rect 5230 320 5231 324
rect 5235 320 5236 324
rect 5230 319 5236 320
rect 5398 324 5404 325
rect 5398 320 5399 324
rect 5403 320 5404 324
rect 5398 319 5404 320
rect 5542 324 5548 325
rect 5542 320 5543 324
rect 5547 320 5548 324
rect 5662 321 5663 325
rect 5667 321 5668 325
rect 5662 320 5668 321
rect 5542 319 5548 320
rect 130 317 136 318
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 130 313 131 317
rect 135 313 136 317
rect 130 312 136 313
rect 274 317 280 318
rect 274 313 275 317
rect 279 313 280 317
rect 274 312 280 313
rect 450 317 456 318
rect 450 313 451 317
rect 455 313 456 317
rect 450 312 456 313
rect 626 317 632 318
rect 626 313 627 317
rect 631 313 632 317
rect 626 312 632 313
rect 802 317 808 318
rect 802 313 803 317
rect 807 313 808 317
rect 802 312 808 313
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 110 311 116 312
rect 1934 311 1940 312
rect 4698 309 4704 310
rect 3838 308 3844 309
rect 1974 305 1980 306
rect 3798 305 3804 306
rect 1974 301 1975 305
rect 1979 301 1980 305
rect 1974 300 1980 301
rect 2022 304 2028 305
rect 2022 300 2023 304
rect 2027 300 2028 304
rect 2022 299 2028 300
rect 2158 304 2164 305
rect 2158 300 2159 304
rect 2163 300 2164 304
rect 2158 299 2164 300
rect 2294 304 2300 305
rect 2294 300 2295 304
rect 2299 300 2300 304
rect 2294 299 2300 300
rect 2430 304 2436 305
rect 2430 300 2431 304
rect 2435 300 2436 304
rect 2430 299 2436 300
rect 2566 304 2572 305
rect 2566 300 2567 304
rect 2571 300 2572 304
rect 2566 299 2572 300
rect 2702 304 2708 305
rect 2702 300 2703 304
rect 2707 300 2708 304
rect 2702 299 2708 300
rect 2838 304 2844 305
rect 2838 300 2839 304
rect 2843 300 2844 304
rect 2838 299 2844 300
rect 2974 304 2980 305
rect 2974 300 2975 304
rect 2979 300 2980 304
rect 2974 299 2980 300
rect 3110 304 3116 305
rect 3110 300 3111 304
rect 3115 300 3116 304
rect 3110 299 3116 300
rect 3246 304 3252 305
rect 3246 300 3247 304
rect 3251 300 3252 304
rect 3246 299 3252 300
rect 3382 304 3388 305
rect 3382 300 3383 304
rect 3387 300 3388 304
rect 3382 299 3388 300
rect 3518 304 3524 305
rect 3518 300 3519 304
rect 3523 300 3524 304
rect 3518 299 3524 300
rect 3654 304 3660 305
rect 3654 300 3655 304
rect 3659 300 3660 304
rect 3798 301 3799 305
rect 3803 301 3804 305
rect 3838 304 3839 308
rect 3843 304 3844 308
rect 4698 305 4699 309
rect 4703 305 4704 309
rect 4698 304 4704 305
rect 4866 309 4872 310
rect 4866 305 4867 309
rect 4871 305 4872 309
rect 4866 304 4872 305
rect 5034 309 5040 310
rect 5034 305 5035 309
rect 5039 305 5040 309
rect 5034 304 5040 305
rect 5202 309 5208 310
rect 5202 305 5203 309
rect 5207 305 5208 309
rect 5202 304 5208 305
rect 5370 309 5376 310
rect 5370 305 5371 309
rect 5375 305 5376 309
rect 5370 304 5376 305
rect 5514 309 5520 310
rect 5514 305 5515 309
rect 5519 305 5520 309
rect 5514 304 5520 305
rect 5662 308 5668 309
rect 5662 304 5663 308
rect 5667 304 5668 308
rect 3838 303 3844 304
rect 5662 303 5668 304
rect 3798 300 3804 301
rect 3654 299 3660 300
rect 1994 289 2000 290
rect 1974 288 1980 289
rect 1974 284 1975 288
rect 1979 284 1980 288
rect 1994 285 1995 289
rect 1999 285 2000 289
rect 1994 284 2000 285
rect 2130 289 2136 290
rect 2130 285 2131 289
rect 2135 285 2136 289
rect 2130 284 2136 285
rect 2266 289 2272 290
rect 2266 285 2267 289
rect 2271 285 2272 289
rect 2266 284 2272 285
rect 2402 289 2408 290
rect 2402 285 2403 289
rect 2407 285 2408 289
rect 2402 284 2408 285
rect 2538 289 2544 290
rect 2538 285 2539 289
rect 2543 285 2544 289
rect 2538 284 2544 285
rect 2674 289 2680 290
rect 2674 285 2675 289
rect 2679 285 2680 289
rect 2674 284 2680 285
rect 2810 289 2816 290
rect 2810 285 2811 289
rect 2815 285 2816 289
rect 2810 284 2816 285
rect 2946 289 2952 290
rect 2946 285 2947 289
rect 2951 285 2952 289
rect 2946 284 2952 285
rect 3082 289 3088 290
rect 3082 285 3083 289
rect 3087 285 3088 289
rect 3082 284 3088 285
rect 3218 289 3224 290
rect 3218 285 3219 289
rect 3223 285 3224 289
rect 3218 284 3224 285
rect 3354 289 3360 290
rect 3354 285 3355 289
rect 3359 285 3360 289
rect 3354 284 3360 285
rect 3490 289 3496 290
rect 3490 285 3491 289
rect 3495 285 3496 289
rect 3490 284 3496 285
rect 3626 289 3632 290
rect 3626 285 3627 289
rect 3631 285 3632 289
rect 3626 284 3632 285
rect 3798 288 3804 289
rect 3798 284 3799 288
rect 3803 284 3804 288
rect 1974 283 1980 284
rect 3798 283 3804 284
rect 110 144 116 145
rect 1934 144 1940 145
rect 110 140 111 144
rect 115 140 116 144
rect 110 139 116 140
rect 130 143 136 144
rect 130 139 131 143
rect 135 139 136 143
rect 130 138 136 139
rect 266 143 272 144
rect 266 139 267 143
rect 271 139 272 143
rect 266 138 272 139
rect 402 143 408 144
rect 402 139 403 143
rect 407 139 408 143
rect 402 138 408 139
rect 538 143 544 144
rect 538 139 539 143
rect 543 139 544 143
rect 538 138 544 139
rect 674 143 680 144
rect 674 139 675 143
rect 679 139 680 143
rect 674 138 680 139
rect 810 143 816 144
rect 810 139 811 143
rect 815 139 816 143
rect 810 138 816 139
rect 946 143 952 144
rect 946 139 947 143
rect 951 139 952 143
rect 946 138 952 139
rect 1082 143 1088 144
rect 1082 139 1083 143
rect 1087 139 1088 143
rect 1934 140 1935 144
rect 1939 140 1940 144
rect 1934 139 1940 140
rect 1082 138 1088 139
rect 3838 136 3844 137
rect 5662 136 5668 137
rect 3838 132 3839 136
rect 3843 132 3844 136
rect 3838 131 3844 132
rect 4290 135 4296 136
rect 4290 131 4291 135
rect 4295 131 4296 135
rect 4290 130 4296 131
rect 4426 135 4432 136
rect 4426 131 4427 135
rect 4431 131 4432 135
rect 4426 130 4432 131
rect 4562 135 4568 136
rect 4562 131 4563 135
rect 4567 131 4568 135
rect 4562 130 4568 131
rect 4698 135 4704 136
rect 4698 131 4699 135
rect 4703 131 4704 135
rect 4698 130 4704 131
rect 4834 135 4840 136
rect 4834 131 4835 135
rect 4839 131 4840 135
rect 4834 130 4840 131
rect 4970 135 4976 136
rect 4970 131 4971 135
rect 4975 131 4976 135
rect 4970 130 4976 131
rect 5106 135 5112 136
rect 5106 131 5107 135
rect 5111 131 5112 135
rect 5106 130 5112 131
rect 5242 135 5248 136
rect 5242 131 5243 135
rect 5247 131 5248 135
rect 5242 130 5248 131
rect 5378 135 5384 136
rect 5378 131 5379 135
rect 5383 131 5384 135
rect 5378 130 5384 131
rect 5514 135 5520 136
rect 5514 131 5515 135
rect 5519 131 5520 135
rect 5662 132 5663 136
rect 5667 132 5668 136
rect 5662 131 5668 132
rect 5514 130 5520 131
rect 158 128 164 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 158 124 159 128
rect 163 124 164 128
rect 158 123 164 124
rect 294 128 300 129
rect 294 124 295 128
rect 299 124 300 128
rect 294 123 300 124
rect 430 128 436 129
rect 430 124 431 128
rect 435 124 436 128
rect 430 123 436 124
rect 566 128 572 129
rect 566 124 567 128
rect 571 124 572 128
rect 566 123 572 124
rect 702 128 708 129
rect 702 124 703 128
rect 707 124 708 128
rect 702 123 708 124
rect 838 128 844 129
rect 838 124 839 128
rect 843 124 844 128
rect 838 123 844 124
rect 974 128 980 129
rect 974 124 975 128
rect 979 124 980 128
rect 974 123 980 124
rect 1110 128 1116 129
rect 1110 124 1111 128
rect 1115 124 1116 128
rect 1110 123 1116 124
rect 1934 127 1940 128
rect 1934 123 1935 127
rect 1939 123 1940 127
rect 110 122 116 123
rect 1934 122 1940 123
rect 1974 124 1980 125
rect 3798 124 3804 125
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 4318 120 4324 121
rect 3798 119 3804 120
rect 3838 119 3844 120
rect 3626 118 3632 119
rect 3838 115 3839 119
rect 3843 115 3844 119
rect 4318 116 4319 120
rect 4323 116 4324 120
rect 4318 115 4324 116
rect 4454 120 4460 121
rect 4454 116 4455 120
rect 4459 116 4460 120
rect 4454 115 4460 116
rect 4590 120 4596 121
rect 4590 116 4591 120
rect 4595 116 4596 120
rect 4590 115 4596 116
rect 4726 120 4732 121
rect 4726 116 4727 120
rect 4731 116 4732 120
rect 4726 115 4732 116
rect 4862 120 4868 121
rect 4862 116 4863 120
rect 4867 116 4868 120
rect 4862 115 4868 116
rect 4998 120 5004 121
rect 4998 116 4999 120
rect 5003 116 5004 120
rect 4998 115 5004 116
rect 5134 120 5140 121
rect 5134 116 5135 120
rect 5139 116 5140 120
rect 5134 115 5140 116
rect 5270 120 5276 121
rect 5270 116 5271 120
rect 5275 116 5276 120
rect 5270 115 5276 116
rect 5406 120 5412 121
rect 5406 116 5407 120
rect 5411 116 5412 120
rect 5406 115 5412 116
rect 5542 120 5548 121
rect 5542 116 5543 120
rect 5547 116 5548 120
rect 5542 115 5548 116
rect 5662 119 5668 120
rect 5662 115 5663 119
rect 5667 115 5668 119
rect 3838 114 3844 115
rect 5662 114 5668 115
rect 2022 108 2028 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2158 108 2164 109
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2430 108 2436 109
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2566 108 2572 109
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2838 108 2844 109
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2974 108 2980 109
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3110 108 3116 109
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3246 108 3252 109
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3382 108 3388 109
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3518 108 3524 109
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3654 108 3660 109
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 1974 102 1980 103
rect 3798 102 3804 103
<< m3c >>
rect 1975 5725 1979 5729
rect 2375 5724 2379 5728
rect 2511 5724 2515 5728
rect 2655 5724 2659 5728
rect 2807 5724 2811 5728
rect 2959 5724 2963 5728
rect 3119 5724 3123 5728
rect 3799 5725 3803 5729
rect 1975 5708 1979 5712
rect 2347 5709 2351 5713
rect 2483 5709 2487 5713
rect 2627 5709 2631 5713
rect 2779 5709 2783 5713
rect 2931 5709 2935 5713
rect 3091 5709 3095 5713
rect 3799 5708 3803 5712
rect 111 5685 115 5689
rect 159 5684 163 5688
rect 295 5684 299 5688
rect 431 5684 435 5688
rect 567 5684 571 5688
rect 703 5684 707 5688
rect 839 5684 843 5688
rect 975 5684 979 5688
rect 1935 5685 1939 5689
rect 111 5668 115 5672
rect 131 5669 135 5673
rect 267 5669 271 5673
rect 403 5669 407 5673
rect 539 5669 543 5673
rect 675 5669 679 5673
rect 811 5669 815 5673
rect 947 5669 951 5673
rect 1935 5668 1939 5672
rect 3839 5649 3843 5653
rect 4335 5648 4339 5652
rect 4471 5648 4475 5652
rect 4607 5648 4611 5652
rect 4743 5648 4747 5652
rect 4879 5648 4883 5652
rect 5015 5648 5019 5652
rect 5663 5649 5667 5653
rect 3839 5632 3843 5636
rect 4307 5633 4311 5637
rect 4443 5633 4447 5637
rect 4579 5633 4583 5637
rect 4715 5633 4719 5637
rect 4851 5633 4855 5637
rect 4987 5633 4991 5637
rect 5663 5632 5667 5636
rect 1975 5576 1979 5580
rect 1995 5575 1999 5579
rect 2203 5575 2207 5579
rect 2427 5575 2431 5579
rect 2651 5575 2655 5579
rect 2867 5575 2871 5579
rect 3075 5575 3079 5579
rect 3275 5575 3279 5579
rect 3475 5575 3479 5579
rect 3651 5575 3655 5579
rect 3799 5576 3803 5580
rect 1975 5559 1979 5563
rect 2023 5560 2027 5564
rect 2231 5560 2235 5564
rect 2455 5560 2459 5564
rect 2679 5560 2683 5564
rect 2895 5560 2899 5564
rect 3103 5560 3107 5564
rect 3303 5560 3307 5564
rect 3503 5560 3507 5564
rect 3679 5560 3683 5564
rect 3799 5559 3803 5563
rect 111 5508 115 5512
rect 619 5507 623 5511
rect 755 5507 759 5511
rect 899 5507 903 5511
rect 1051 5507 1055 5511
rect 1203 5507 1207 5511
rect 1355 5507 1359 5511
rect 1507 5507 1511 5511
rect 1651 5507 1655 5511
rect 1787 5507 1791 5511
rect 1935 5508 1939 5512
rect 1975 5501 1979 5505
rect 2951 5500 2955 5504
rect 3103 5500 3107 5504
rect 3255 5500 3259 5504
rect 3415 5500 3419 5504
rect 3799 5501 3803 5505
rect 3839 5500 3843 5504
rect 4211 5499 4215 5503
rect 4403 5499 4407 5503
rect 4595 5499 4599 5503
rect 4795 5499 4799 5503
rect 4995 5499 4999 5503
rect 5195 5499 5199 5503
rect 5663 5500 5667 5504
rect 111 5491 115 5495
rect 647 5492 651 5496
rect 783 5492 787 5496
rect 927 5492 931 5496
rect 1079 5492 1083 5496
rect 1231 5492 1235 5496
rect 1383 5492 1387 5496
rect 1535 5492 1539 5496
rect 1679 5492 1683 5496
rect 1815 5492 1819 5496
rect 1935 5491 1939 5495
rect 1975 5484 1979 5488
rect 2923 5485 2927 5489
rect 3075 5485 3079 5489
rect 3227 5485 3231 5489
rect 3387 5485 3391 5489
rect 3799 5484 3803 5488
rect 3839 5483 3843 5487
rect 4239 5484 4243 5488
rect 4431 5484 4435 5488
rect 4623 5484 4627 5488
rect 4823 5484 4827 5488
rect 5023 5484 5027 5488
rect 5223 5484 5227 5488
rect 5663 5483 5667 5487
rect 111 5425 115 5429
rect 591 5424 595 5428
rect 727 5424 731 5428
rect 863 5424 867 5428
rect 999 5424 1003 5428
rect 1135 5424 1139 5428
rect 1271 5424 1275 5428
rect 1407 5424 1411 5428
rect 1543 5424 1547 5428
rect 1679 5424 1683 5428
rect 1815 5424 1819 5428
rect 1935 5425 1939 5429
rect 111 5408 115 5412
rect 563 5409 567 5413
rect 699 5409 703 5413
rect 835 5409 839 5413
rect 971 5409 975 5413
rect 1107 5409 1111 5413
rect 1243 5409 1247 5413
rect 1379 5409 1383 5413
rect 1515 5409 1519 5413
rect 1651 5409 1655 5413
rect 1787 5409 1791 5413
rect 1935 5408 1939 5412
rect 3839 5389 3843 5393
rect 4303 5388 4307 5392
rect 4519 5388 4523 5392
rect 4735 5388 4739 5392
rect 4951 5388 4955 5392
rect 5175 5388 5179 5392
rect 5399 5388 5403 5392
rect 5663 5389 5667 5393
rect 3839 5372 3843 5376
rect 4275 5373 4279 5377
rect 4491 5373 4495 5377
rect 4707 5373 4711 5377
rect 4923 5373 4927 5377
rect 5147 5373 5151 5377
rect 5371 5373 5375 5377
rect 5663 5372 5667 5376
rect 1975 5304 1979 5308
rect 2643 5303 2647 5307
rect 2811 5303 2815 5307
rect 2979 5303 2983 5307
rect 3139 5303 3143 5307
rect 3307 5303 3311 5307
rect 3475 5303 3479 5307
rect 3643 5303 3647 5307
rect 3799 5304 3803 5308
rect 1975 5287 1979 5291
rect 2671 5288 2675 5292
rect 2839 5288 2843 5292
rect 3007 5288 3011 5292
rect 3167 5288 3171 5292
rect 3335 5288 3339 5292
rect 3503 5288 3507 5292
rect 3671 5288 3675 5292
rect 3799 5287 3803 5291
rect 111 5252 115 5256
rect 411 5251 415 5255
rect 587 5251 591 5255
rect 763 5251 767 5255
rect 939 5251 943 5255
rect 1107 5251 1111 5255
rect 1275 5251 1279 5255
rect 1443 5251 1447 5255
rect 1611 5251 1615 5255
rect 1787 5251 1791 5255
rect 1935 5252 1939 5256
rect 111 5235 115 5239
rect 439 5236 443 5240
rect 615 5236 619 5240
rect 791 5236 795 5240
rect 967 5236 971 5240
rect 1135 5236 1139 5240
rect 1303 5236 1307 5240
rect 1471 5236 1475 5240
rect 1639 5236 1643 5240
rect 1815 5236 1819 5240
rect 1935 5235 1939 5239
rect 1975 5229 1979 5233
rect 2511 5228 2515 5232
rect 2687 5228 2691 5232
rect 2863 5228 2867 5232
rect 3039 5228 3043 5232
rect 3207 5228 3211 5232
rect 3367 5228 3371 5232
rect 3535 5228 3539 5232
rect 3679 5228 3683 5232
rect 3799 5229 3803 5233
rect 1975 5212 1979 5216
rect 2483 5213 2487 5217
rect 2659 5213 2663 5217
rect 2835 5213 2839 5217
rect 3011 5213 3015 5217
rect 3179 5213 3183 5217
rect 3339 5213 3343 5217
rect 3507 5213 3511 5217
rect 3651 5213 3655 5217
rect 3799 5212 3803 5216
rect 3839 5208 3843 5212
rect 4371 5207 4375 5211
rect 4563 5207 4567 5211
rect 4771 5207 4775 5211
rect 4979 5207 4983 5211
rect 5195 5207 5199 5211
rect 5419 5207 5423 5211
rect 5663 5208 5667 5212
rect 3839 5191 3843 5195
rect 4399 5192 4403 5196
rect 4591 5192 4595 5196
rect 4799 5192 4803 5196
rect 5007 5192 5011 5196
rect 5223 5192 5227 5196
rect 5447 5192 5451 5196
rect 5663 5191 5667 5195
rect 111 5169 115 5173
rect 207 5168 211 5172
rect 343 5168 347 5172
rect 479 5168 483 5172
rect 615 5168 619 5172
rect 751 5168 755 5172
rect 887 5168 891 5172
rect 1023 5168 1027 5172
rect 1935 5169 1939 5173
rect 111 5152 115 5156
rect 179 5153 183 5157
rect 315 5153 319 5157
rect 451 5153 455 5157
rect 587 5153 591 5157
rect 723 5153 727 5157
rect 859 5153 863 5157
rect 995 5153 999 5157
rect 1935 5152 1939 5156
rect 3839 5109 3843 5113
rect 3887 5108 3891 5112
rect 4087 5108 4091 5112
rect 4311 5108 4315 5112
rect 4535 5108 4539 5112
rect 4759 5108 4763 5112
rect 4983 5108 4987 5112
rect 5207 5108 5211 5112
rect 5439 5108 5443 5112
rect 5663 5109 5667 5113
rect 3839 5092 3843 5096
rect 3859 5093 3863 5097
rect 4059 5093 4063 5097
rect 4283 5093 4287 5097
rect 4507 5093 4511 5097
rect 4731 5093 4735 5097
rect 4955 5093 4959 5097
rect 5179 5093 5183 5097
rect 5411 5093 5415 5097
rect 5663 5092 5667 5096
rect 1975 5072 1979 5076
rect 2139 5071 2143 5075
rect 2307 5071 2311 5075
rect 2491 5071 2495 5075
rect 2691 5071 2695 5075
rect 2915 5071 2919 5075
rect 3163 5071 3167 5075
rect 3419 5071 3423 5075
rect 3651 5071 3655 5075
rect 3799 5072 3803 5076
rect 1975 5055 1979 5059
rect 2167 5056 2171 5060
rect 2335 5056 2339 5060
rect 2519 5056 2523 5060
rect 2719 5056 2723 5060
rect 2943 5056 2947 5060
rect 3191 5056 3195 5060
rect 3447 5056 3451 5060
rect 3679 5056 3683 5060
rect 3799 5055 3803 5059
rect 111 5000 115 5004
rect 147 4999 151 5003
rect 339 4999 343 5003
rect 531 4999 535 5003
rect 731 4999 735 5003
rect 931 4999 935 5003
rect 1131 4999 1135 5003
rect 1935 5000 1939 5004
rect 111 4983 115 4987
rect 175 4984 179 4988
rect 367 4984 371 4988
rect 559 4984 563 4988
rect 759 4984 763 4988
rect 959 4984 963 4988
rect 1159 4984 1163 4988
rect 1935 4983 1939 4987
rect 1975 4973 1979 4977
rect 2023 4972 2027 4976
rect 2167 4972 2171 4976
rect 2351 4972 2355 4976
rect 2543 4972 2547 4976
rect 2751 4972 2755 4976
rect 2967 4972 2971 4976
rect 3183 4972 3187 4976
rect 3799 4973 3803 4977
rect 1975 4956 1979 4960
rect 1995 4957 1999 4961
rect 2139 4957 2143 4961
rect 2323 4957 2327 4961
rect 2515 4957 2519 4961
rect 2723 4957 2727 4961
rect 2939 4957 2943 4961
rect 3155 4957 3159 4961
rect 3799 4956 3803 4960
rect 3839 4944 3843 4948
rect 3859 4943 3863 4947
rect 3995 4943 3999 4947
rect 4131 4943 4135 4947
rect 4283 4943 4287 4947
rect 4443 4943 4447 4947
rect 4611 4943 4615 4947
rect 4787 4943 4791 4947
rect 4971 4943 4975 4947
rect 5155 4943 5159 4947
rect 5339 4943 5343 4947
rect 5515 4943 5519 4947
rect 5663 4944 5667 4948
rect 3839 4927 3843 4931
rect 3887 4928 3891 4932
rect 4023 4928 4027 4932
rect 4159 4928 4163 4932
rect 4311 4928 4315 4932
rect 4471 4928 4475 4932
rect 4639 4928 4643 4932
rect 4815 4928 4819 4932
rect 4999 4928 5003 4932
rect 5183 4928 5187 4932
rect 5367 4928 5371 4932
rect 5543 4928 5547 4932
rect 5663 4927 5667 4931
rect 111 4913 115 4917
rect 159 4912 163 4916
rect 391 4912 395 4916
rect 647 4912 651 4916
rect 895 4912 899 4916
rect 1135 4912 1139 4916
rect 1367 4912 1371 4916
rect 1599 4912 1603 4916
rect 1815 4912 1819 4916
rect 1935 4913 1939 4917
rect 111 4896 115 4900
rect 131 4897 135 4901
rect 363 4897 367 4901
rect 619 4897 623 4901
rect 867 4897 871 4901
rect 1107 4897 1111 4901
rect 1339 4897 1343 4901
rect 1571 4897 1575 4901
rect 1787 4897 1791 4901
rect 1935 4896 1939 4900
rect 3839 4853 3843 4857
rect 3943 4852 3947 4856
rect 4183 4852 4187 4856
rect 4431 4852 4435 4856
rect 4687 4852 4691 4856
rect 4959 4852 4963 4856
rect 5239 4852 5243 4856
rect 5519 4852 5523 4856
rect 5663 4853 5667 4857
rect 3839 4836 3843 4840
rect 3915 4837 3919 4841
rect 4155 4837 4159 4841
rect 4403 4837 4407 4841
rect 4659 4837 4663 4841
rect 4931 4837 4935 4841
rect 5211 4837 5215 4841
rect 5491 4837 5495 4841
rect 5663 4836 5667 4840
rect 1975 4816 1979 4820
rect 1995 4815 1999 4819
rect 2323 4815 2327 4819
rect 2667 4815 2671 4819
rect 3019 4815 3023 4819
rect 3371 4815 3375 4819
rect 3799 4816 3803 4820
rect 1975 4799 1979 4803
rect 2023 4800 2027 4804
rect 2351 4800 2355 4804
rect 2695 4800 2699 4804
rect 3047 4800 3051 4804
rect 3399 4800 3403 4804
rect 3799 4799 3803 4803
rect 111 4764 115 4768
rect 131 4763 135 4767
rect 475 4763 479 4767
rect 859 4763 863 4767
rect 1251 4763 1255 4767
rect 1643 4763 1647 4767
rect 1935 4764 1939 4768
rect 111 4747 115 4751
rect 159 4748 163 4752
rect 503 4748 507 4752
rect 887 4748 891 4752
rect 1279 4748 1283 4752
rect 1671 4748 1675 4752
rect 1935 4747 1939 4751
rect 1975 4693 1979 4697
rect 2079 4692 2083 4696
rect 2231 4692 2235 4696
rect 2391 4692 2395 4696
rect 2559 4692 2563 4696
rect 2727 4692 2731 4696
rect 2903 4692 2907 4696
rect 3079 4692 3083 4696
rect 3255 4692 3259 4696
rect 3439 4692 3443 4696
rect 3623 4692 3627 4696
rect 3799 4693 3803 4697
rect 3839 4696 3843 4700
rect 3939 4695 3943 4699
rect 4179 4695 4183 4699
rect 4435 4695 4439 4699
rect 4691 4695 4695 4699
rect 4955 4695 4959 4699
rect 5227 4695 5231 4699
rect 5507 4695 5511 4699
rect 5663 4696 5667 4700
rect 1975 4676 1979 4680
rect 2051 4677 2055 4681
rect 2203 4677 2207 4681
rect 2363 4677 2367 4681
rect 2531 4677 2535 4681
rect 2699 4677 2703 4681
rect 2875 4677 2879 4681
rect 3051 4677 3055 4681
rect 3227 4677 3231 4681
rect 3411 4677 3415 4681
rect 3595 4677 3599 4681
rect 3799 4676 3803 4680
rect 3839 4679 3843 4683
rect 3967 4680 3971 4684
rect 4207 4680 4211 4684
rect 4463 4680 4467 4684
rect 4719 4680 4723 4684
rect 4983 4680 4987 4684
rect 5255 4680 5259 4684
rect 5535 4680 5539 4684
rect 5663 4679 5667 4683
rect 111 4669 115 4673
rect 159 4668 163 4672
rect 295 4668 299 4672
rect 431 4668 435 4672
rect 567 4668 571 4672
rect 703 4668 707 4672
rect 1935 4669 1939 4673
rect 111 4652 115 4656
rect 131 4653 135 4657
rect 267 4653 271 4657
rect 403 4653 407 4657
rect 539 4653 543 4657
rect 675 4653 679 4657
rect 1935 4652 1939 4656
rect 3839 4617 3843 4621
rect 4175 4616 4179 4620
rect 4455 4616 4459 4620
rect 4735 4616 4739 4620
rect 5015 4616 5019 4620
rect 5303 4616 5307 4620
rect 5663 4617 5667 4621
rect 3839 4600 3843 4604
rect 4147 4601 4151 4605
rect 4427 4601 4431 4605
rect 4707 4601 4711 4605
rect 4987 4601 4991 4605
rect 5275 4601 5279 4605
rect 5663 4600 5667 4604
rect 1975 4540 1979 4544
rect 2123 4539 2127 4543
rect 2275 4539 2279 4543
rect 2443 4539 2447 4543
rect 2611 4539 2615 4543
rect 2787 4539 2791 4543
rect 2963 4539 2967 4543
rect 3139 4539 3143 4543
rect 3315 4539 3319 4543
rect 3491 4539 3495 4543
rect 3651 4539 3655 4543
rect 3799 4540 3803 4544
rect 1975 4523 1979 4527
rect 2151 4524 2155 4528
rect 2303 4524 2307 4528
rect 2471 4524 2475 4528
rect 2639 4524 2643 4528
rect 2815 4524 2819 4528
rect 2991 4524 2995 4528
rect 3167 4524 3171 4528
rect 3343 4524 3347 4528
rect 3519 4524 3523 4528
rect 3679 4524 3683 4528
rect 3799 4523 3803 4527
rect 111 4504 115 4508
rect 291 4503 295 4507
rect 427 4503 431 4507
rect 563 4503 567 4507
rect 699 4503 703 4507
rect 835 4503 839 4507
rect 1935 4504 1939 4508
rect 111 4487 115 4491
rect 319 4488 323 4492
rect 455 4488 459 4492
rect 591 4488 595 4492
rect 727 4488 731 4492
rect 863 4488 867 4492
rect 1935 4487 1939 4491
rect 3839 4464 3843 4468
rect 3859 4463 3863 4467
rect 4155 4463 4159 4467
rect 4483 4463 4487 4467
rect 4819 4463 4823 4467
rect 5163 4463 5167 4467
rect 5515 4463 5519 4467
rect 5663 4464 5667 4468
rect 1975 4457 1979 4461
rect 2023 4456 2027 4460
rect 2159 4456 2163 4460
rect 2295 4456 2299 4460
rect 2431 4456 2435 4460
rect 2567 4456 2571 4460
rect 2703 4456 2707 4460
rect 2839 4456 2843 4460
rect 2975 4456 2979 4460
rect 3799 4457 3803 4461
rect 3839 4447 3843 4451
rect 3887 4448 3891 4452
rect 4183 4448 4187 4452
rect 4511 4448 4515 4452
rect 4847 4448 4851 4452
rect 5191 4448 5195 4452
rect 5543 4448 5547 4452
rect 5663 4447 5667 4451
rect 1975 4440 1979 4444
rect 1995 4441 1999 4445
rect 2131 4441 2135 4445
rect 2267 4441 2271 4445
rect 2403 4441 2407 4445
rect 2539 4441 2543 4445
rect 2675 4441 2679 4445
rect 2811 4441 2815 4445
rect 2947 4441 2951 4445
rect 3799 4440 3803 4444
rect 111 4413 115 4417
rect 519 4412 523 4416
rect 743 4412 747 4416
rect 991 4412 995 4416
rect 1263 4412 1267 4416
rect 1551 4412 1555 4416
rect 1815 4412 1819 4416
rect 1935 4413 1939 4417
rect 111 4396 115 4400
rect 491 4397 495 4401
rect 715 4397 719 4401
rect 963 4397 967 4401
rect 1235 4397 1239 4401
rect 1523 4397 1527 4401
rect 1787 4397 1791 4401
rect 1935 4396 1939 4400
rect 3839 4389 3843 4393
rect 3887 4388 3891 4392
rect 4143 4388 4147 4392
rect 4423 4388 4427 4392
rect 4703 4388 4707 4392
rect 4983 4388 4987 4392
rect 5263 4388 5267 4392
rect 5543 4388 5547 4392
rect 5663 4389 5667 4393
rect 3839 4372 3843 4376
rect 3859 4373 3863 4377
rect 4115 4373 4119 4377
rect 4395 4373 4399 4377
rect 4675 4373 4679 4377
rect 4955 4373 4959 4377
rect 5235 4373 5239 4377
rect 5515 4373 5519 4377
rect 5663 4372 5667 4376
rect 1975 4292 1979 4296
rect 2779 4291 2783 4295
rect 2995 4291 2999 4295
rect 3219 4291 3223 4295
rect 3443 4291 3447 4295
rect 3651 4291 3655 4295
rect 3799 4292 3803 4296
rect 1975 4275 1979 4279
rect 2807 4276 2811 4280
rect 3023 4276 3027 4280
rect 3247 4276 3251 4280
rect 3471 4276 3475 4280
rect 3679 4276 3683 4280
rect 3799 4275 3803 4279
rect 111 4264 115 4268
rect 563 4263 567 4267
rect 699 4263 703 4267
rect 835 4263 839 4267
rect 971 4263 975 4267
rect 1107 4263 1111 4267
rect 1243 4263 1247 4267
rect 1379 4263 1383 4267
rect 1515 4263 1519 4267
rect 1651 4263 1655 4267
rect 1787 4263 1791 4267
rect 1935 4264 1939 4268
rect 111 4247 115 4251
rect 591 4248 595 4252
rect 727 4248 731 4252
rect 863 4248 867 4252
rect 999 4248 1003 4252
rect 1135 4248 1139 4252
rect 1271 4248 1275 4252
rect 1407 4248 1411 4252
rect 1543 4248 1547 4252
rect 1679 4248 1683 4252
rect 1815 4248 1819 4252
rect 1935 4247 1939 4251
rect 3839 4228 3843 4232
rect 4571 4227 4575 4231
rect 4739 4227 4743 4231
rect 4915 4227 4919 4231
rect 5107 4227 5111 4231
rect 5307 4227 5311 4231
rect 5515 4227 5519 4231
rect 5663 4228 5667 4232
rect 3839 4211 3843 4215
rect 4599 4212 4603 4216
rect 4767 4212 4771 4216
rect 4943 4212 4947 4216
rect 5135 4212 5139 4216
rect 5335 4212 5339 4216
rect 5543 4212 5547 4216
rect 5663 4211 5667 4215
rect 1975 4189 1979 4193
rect 2951 4188 2955 4192
rect 3095 4188 3099 4192
rect 3239 4188 3243 4192
rect 3391 4188 3395 4192
rect 3543 4188 3547 4192
rect 3679 4188 3683 4192
rect 3799 4189 3803 4193
rect 111 4177 115 4181
rect 591 4176 595 4180
rect 727 4176 731 4180
rect 863 4176 867 4180
rect 999 4176 1003 4180
rect 1135 4176 1139 4180
rect 1271 4176 1275 4180
rect 1407 4176 1411 4180
rect 1543 4176 1547 4180
rect 1679 4176 1683 4180
rect 1815 4176 1819 4180
rect 1935 4177 1939 4181
rect 1975 4172 1979 4176
rect 2923 4173 2927 4177
rect 3067 4173 3071 4177
rect 3211 4173 3215 4177
rect 3363 4173 3367 4177
rect 3515 4173 3519 4177
rect 3651 4173 3655 4177
rect 3799 4172 3803 4176
rect 111 4160 115 4164
rect 563 4161 567 4165
rect 699 4161 703 4165
rect 835 4161 839 4165
rect 971 4161 975 4165
rect 1107 4161 1111 4165
rect 1243 4161 1247 4165
rect 1379 4161 1383 4165
rect 1515 4161 1519 4165
rect 1651 4161 1655 4165
rect 1787 4161 1791 4165
rect 1935 4160 1939 4164
rect 3839 4153 3843 4157
rect 4655 4152 4659 4156
rect 4815 4152 4819 4156
rect 4983 4152 4987 4156
rect 5167 4152 5171 4156
rect 5359 4152 5363 4156
rect 5543 4152 5547 4156
rect 5663 4153 5667 4157
rect 3839 4136 3843 4140
rect 4627 4137 4631 4141
rect 4787 4137 4791 4141
rect 4955 4137 4959 4141
rect 5139 4137 5143 4141
rect 5331 4137 5335 4141
rect 5515 4137 5519 4141
rect 5663 4136 5667 4140
rect 111 4028 115 4032
rect 699 4027 703 4031
rect 835 4027 839 4031
rect 971 4027 975 4031
rect 1107 4027 1111 4031
rect 1243 4027 1247 4031
rect 1379 4027 1383 4031
rect 1515 4027 1519 4031
rect 1651 4027 1655 4031
rect 1787 4027 1791 4031
rect 1935 4028 1939 4032
rect 111 4011 115 4015
rect 727 4012 731 4016
rect 863 4012 867 4016
rect 999 4012 1003 4016
rect 1135 4012 1139 4016
rect 1271 4012 1275 4016
rect 1407 4012 1411 4016
rect 1543 4012 1547 4016
rect 1679 4012 1683 4016
rect 1815 4012 1819 4016
rect 1935 4011 1939 4015
rect 1975 4004 1979 4008
rect 2899 4003 2903 4007
rect 3043 4003 3047 4007
rect 3187 4003 3191 4007
rect 3339 4003 3343 4007
rect 3491 4003 3495 4007
rect 3643 4003 3647 4007
rect 3799 4004 3803 4008
rect 1975 3987 1979 3991
rect 2927 3988 2931 3992
rect 3071 3988 3075 3992
rect 3215 3988 3219 3992
rect 3367 3988 3371 3992
rect 3519 3988 3523 3992
rect 3671 3988 3675 3992
rect 3799 3987 3803 3991
rect 3839 3968 3843 3972
rect 4939 3967 4943 3971
rect 5075 3967 5079 3971
rect 5211 3967 5215 3971
rect 5347 3967 5351 3971
rect 5663 3968 5667 3972
rect 111 3949 115 3953
rect 695 3948 699 3952
rect 831 3948 835 3952
rect 967 3948 971 3952
rect 1111 3948 1115 3952
rect 1255 3948 1259 3952
rect 1399 3948 1403 3952
rect 1543 3948 1547 3952
rect 1679 3948 1683 3952
rect 1815 3948 1819 3952
rect 1935 3949 1939 3953
rect 3839 3951 3843 3955
rect 4967 3952 4971 3956
rect 5103 3952 5107 3956
rect 5239 3952 5243 3956
rect 5375 3952 5379 3956
rect 5663 3951 5667 3955
rect 111 3932 115 3936
rect 667 3933 671 3937
rect 803 3933 807 3937
rect 939 3933 943 3937
rect 1083 3933 1087 3937
rect 1227 3933 1231 3937
rect 1371 3933 1375 3937
rect 1515 3933 1519 3937
rect 1651 3933 1655 3937
rect 1787 3933 1791 3937
rect 1935 3932 1939 3936
rect 1975 3901 1979 3905
rect 2759 3900 2763 3904
rect 2911 3900 2915 3904
rect 3071 3900 3075 3904
rect 3239 3900 3243 3904
rect 3415 3900 3419 3904
rect 3591 3900 3595 3904
rect 3799 3901 3803 3905
rect 3839 3893 3843 3897
rect 4687 3892 4691 3896
rect 4847 3892 4851 3896
rect 5015 3892 5019 3896
rect 5191 3892 5195 3896
rect 5375 3892 5379 3896
rect 5543 3892 5547 3896
rect 5663 3893 5667 3897
rect 1975 3884 1979 3888
rect 2731 3885 2735 3889
rect 2883 3885 2887 3889
rect 3043 3885 3047 3889
rect 3211 3885 3215 3889
rect 3387 3885 3391 3889
rect 3563 3885 3567 3889
rect 3799 3884 3803 3888
rect 3839 3876 3843 3880
rect 4659 3877 4663 3881
rect 4819 3877 4823 3881
rect 4987 3877 4991 3881
rect 5163 3877 5167 3881
rect 5347 3877 5351 3881
rect 5515 3877 5519 3881
rect 5663 3876 5667 3880
rect 111 3796 115 3800
rect 435 3795 439 3799
rect 619 3795 623 3799
rect 819 3795 823 3799
rect 1027 3795 1031 3799
rect 1251 3795 1255 3799
rect 1483 3795 1487 3799
rect 1723 3795 1727 3799
rect 1935 3796 1939 3800
rect 111 3779 115 3783
rect 463 3780 467 3784
rect 647 3780 651 3784
rect 847 3780 851 3784
rect 1055 3780 1059 3784
rect 1279 3780 1283 3784
rect 1511 3780 1515 3784
rect 1751 3780 1755 3784
rect 1935 3779 1939 3783
rect 1975 3744 1979 3748
rect 2115 3743 2119 3747
rect 2251 3743 2255 3747
rect 2387 3743 2391 3747
rect 2523 3743 2527 3747
rect 2659 3743 2663 3747
rect 2795 3743 2799 3747
rect 2939 3743 2943 3747
rect 3083 3743 3087 3747
rect 3235 3743 3239 3747
rect 3395 3743 3399 3747
rect 3555 3743 3559 3747
rect 3799 3744 3803 3748
rect 3839 3744 3843 3748
rect 4411 3743 4415 3747
rect 4619 3743 4623 3747
rect 4835 3743 4839 3747
rect 5067 3743 5071 3747
rect 5299 3743 5303 3747
rect 5515 3743 5519 3747
rect 5663 3744 5667 3748
rect 1975 3727 1979 3731
rect 2143 3728 2147 3732
rect 2279 3728 2283 3732
rect 2415 3728 2419 3732
rect 2551 3728 2555 3732
rect 2687 3728 2691 3732
rect 2823 3728 2827 3732
rect 2967 3728 2971 3732
rect 3111 3728 3115 3732
rect 3263 3728 3267 3732
rect 3423 3728 3427 3732
rect 3583 3728 3587 3732
rect 3799 3727 3803 3731
rect 3839 3727 3843 3731
rect 4439 3728 4443 3732
rect 4647 3728 4651 3732
rect 4863 3728 4867 3732
rect 5095 3728 5099 3732
rect 5327 3728 5331 3732
rect 5543 3728 5547 3732
rect 5663 3727 5667 3731
rect 111 3717 115 3721
rect 231 3716 235 3720
rect 431 3716 435 3720
rect 655 3716 659 3720
rect 895 3716 899 3720
rect 1151 3716 1155 3720
rect 1415 3716 1419 3720
rect 1679 3716 1683 3720
rect 1935 3717 1939 3721
rect 111 3700 115 3704
rect 203 3701 207 3705
rect 403 3701 407 3705
rect 627 3701 631 3705
rect 867 3701 871 3705
rect 1123 3701 1127 3705
rect 1387 3701 1391 3705
rect 1651 3701 1655 3705
rect 1935 3700 1939 3704
rect 1975 3661 1979 3665
rect 2231 3660 2235 3664
rect 2447 3660 2451 3664
rect 2663 3660 2667 3664
rect 2871 3660 2875 3664
rect 3079 3660 3083 3664
rect 3287 3660 3291 3664
rect 3495 3660 3499 3664
rect 3679 3660 3683 3664
rect 3799 3661 3803 3665
rect 1975 3644 1979 3648
rect 2203 3645 2207 3649
rect 2419 3645 2423 3649
rect 2635 3645 2639 3649
rect 2843 3645 2847 3649
rect 3051 3645 3055 3649
rect 3259 3645 3263 3649
rect 3467 3645 3471 3649
rect 3651 3645 3655 3649
rect 3799 3644 3803 3648
rect 3839 3645 3843 3649
rect 3887 3644 3891 3648
rect 4047 3644 4051 3648
rect 4247 3644 4251 3648
rect 4479 3644 4483 3648
rect 4727 3644 4731 3648
rect 4999 3644 5003 3648
rect 5279 3644 5283 3648
rect 5543 3644 5547 3648
rect 5663 3645 5667 3649
rect 3839 3628 3843 3632
rect 3859 3629 3863 3633
rect 4019 3629 4023 3633
rect 4219 3629 4223 3633
rect 4451 3629 4455 3633
rect 4699 3629 4703 3633
rect 4971 3629 4975 3633
rect 5251 3629 5255 3633
rect 5515 3629 5519 3633
rect 5663 3628 5667 3632
rect 111 3560 115 3564
rect 131 3559 135 3563
rect 315 3559 319 3563
rect 539 3559 543 3563
rect 787 3559 791 3563
rect 1043 3559 1047 3563
rect 1315 3559 1319 3563
rect 1587 3559 1591 3563
rect 1935 3560 1939 3564
rect 111 3543 115 3547
rect 159 3544 163 3548
rect 343 3544 347 3548
rect 567 3544 571 3548
rect 815 3544 819 3548
rect 1071 3544 1075 3548
rect 1343 3544 1347 3548
rect 1615 3544 1619 3548
rect 1935 3543 1939 3547
rect 1975 3496 1979 3500
rect 2163 3495 2167 3499
rect 2299 3495 2303 3499
rect 2435 3495 2439 3499
rect 2571 3495 2575 3499
rect 3799 3496 3803 3500
rect 1975 3479 1979 3483
rect 2191 3480 2195 3484
rect 2327 3480 2331 3484
rect 2463 3480 2467 3484
rect 3839 3484 3843 3488
rect 2599 3480 2603 3484
rect 3859 3483 3863 3487
rect 3799 3479 3803 3483
rect 3995 3483 3999 3487
rect 4131 3483 4135 3487
rect 4267 3483 4271 3487
rect 4403 3483 4407 3487
rect 4539 3483 4543 3487
rect 4699 3483 4703 3487
rect 4891 3483 4895 3487
rect 5099 3483 5103 3487
rect 5315 3483 5319 3487
rect 5515 3483 5519 3487
rect 5663 3484 5667 3488
rect 111 3473 115 3477
rect 159 3472 163 3476
rect 335 3472 339 3476
rect 551 3472 555 3476
rect 791 3472 795 3476
rect 1039 3472 1043 3476
rect 1295 3472 1299 3476
rect 1559 3472 1563 3476
rect 1935 3473 1939 3477
rect 3839 3467 3843 3471
rect 3887 3468 3891 3472
rect 4023 3468 4027 3472
rect 4159 3468 4163 3472
rect 4295 3468 4299 3472
rect 4431 3468 4435 3472
rect 4567 3468 4571 3472
rect 4727 3468 4731 3472
rect 4919 3468 4923 3472
rect 5127 3468 5131 3472
rect 5343 3468 5347 3472
rect 5543 3468 5547 3472
rect 5663 3467 5667 3471
rect 111 3456 115 3460
rect 131 3457 135 3461
rect 307 3457 311 3461
rect 523 3457 527 3461
rect 763 3457 767 3461
rect 1011 3457 1015 3461
rect 1267 3457 1271 3461
rect 1531 3457 1535 3461
rect 1935 3456 1939 3460
rect 3839 3401 3843 3405
rect 3887 3400 3891 3404
rect 4023 3400 4027 3404
rect 4159 3400 4163 3404
rect 4295 3400 4299 3404
rect 4431 3400 4435 3404
rect 4583 3400 4587 3404
rect 4759 3400 4763 3404
rect 4951 3400 4955 3404
rect 5151 3400 5155 3404
rect 5359 3400 5363 3404
rect 5543 3400 5547 3404
rect 5663 3401 5667 3405
rect 1975 3385 1979 3389
rect 2231 3384 2235 3388
rect 2583 3384 2587 3388
rect 2951 3384 2955 3388
rect 3327 3384 3331 3388
rect 3679 3384 3683 3388
rect 3799 3385 3803 3389
rect 3839 3384 3843 3388
rect 3859 3385 3863 3389
rect 3995 3385 3999 3389
rect 4131 3385 4135 3389
rect 4267 3385 4271 3389
rect 4403 3385 4407 3389
rect 4555 3385 4559 3389
rect 4731 3385 4735 3389
rect 4923 3385 4927 3389
rect 5123 3385 5127 3389
rect 5331 3385 5335 3389
rect 5515 3385 5519 3389
rect 5663 3384 5667 3388
rect 1975 3368 1979 3372
rect 2203 3369 2207 3373
rect 2555 3369 2559 3373
rect 2923 3369 2927 3373
rect 3299 3369 3303 3373
rect 3651 3369 3655 3373
rect 3799 3368 3803 3372
rect 111 3316 115 3320
rect 131 3315 135 3319
rect 299 3315 303 3319
rect 507 3315 511 3319
rect 731 3315 735 3319
rect 971 3315 975 3319
rect 1219 3315 1223 3319
rect 1475 3315 1479 3319
rect 1935 3316 1939 3320
rect 111 3299 115 3303
rect 159 3300 163 3304
rect 327 3300 331 3304
rect 535 3300 539 3304
rect 759 3300 763 3304
rect 999 3300 1003 3304
rect 1247 3300 1251 3304
rect 1503 3300 1507 3304
rect 1935 3299 1939 3303
rect 111 3237 115 3241
rect 239 3236 243 3240
rect 463 3236 467 3240
rect 703 3236 707 3240
rect 951 3236 955 3240
rect 1199 3236 1203 3240
rect 1455 3236 1459 3240
rect 1935 3237 1939 3241
rect 1975 3236 1979 3240
rect 2251 3235 2255 3239
rect 2475 3235 2479 3239
rect 2691 3235 2695 3239
rect 2899 3235 2903 3239
rect 3099 3235 3103 3239
rect 3291 3235 3295 3239
rect 3483 3235 3487 3239
rect 3651 3235 3655 3239
rect 3799 3236 3803 3240
rect 3839 3236 3843 3240
rect 4691 3235 4695 3239
rect 4827 3235 4831 3239
rect 4963 3235 4967 3239
rect 5099 3235 5103 3239
rect 5235 3235 5239 3239
rect 5663 3236 5667 3240
rect 111 3220 115 3224
rect 211 3221 215 3225
rect 435 3221 439 3225
rect 675 3221 679 3225
rect 923 3221 927 3225
rect 1171 3221 1175 3225
rect 1427 3221 1431 3225
rect 1935 3220 1939 3224
rect 1975 3219 1979 3223
rect 2279 3220 2283 3224
rect 2503 3220 2507 3224
rect 2719 3220 2723 3224
rect 2927 3220 2931 3224
rect 3127 3220 3131 3224
rect 3319 3220 3323 3224
rect 3511 3220 3515 3224
rect 3679 3220 3683 3224
rect 3799 3219 3803 3223
rect 3839 3219 3843 3223
rect 4719 3220 4723 3224
rect 4855 3220 4859 3224
rect 4991 3220 4995 3224
rect 5127 3220 5131 3224
rect 5263 3220 5267 3224
rect 5663 3219 5667 3223
rect 1975 3153 1979 3157
rect 2095 3152 2099 3156
rect 2295 3152 2299 3156
rect 2487 3152 2491 3156
rect 2679 3152 2683 3156
rect 2871 3152 2875 3156
rect 3055 3152 3059 3156
rect 3231 3152 3235 3156
rect 3415 3152 3419 3156
rect 3599 3152 3603 3156
rect 3799 3153 3803 3157
rect 3839 3153 3843 3157
rect 4863 3152 4867 3156
rect 4999 3152 5003 3156
rect 5135 3152 5139 3156
rect 5271 3152 5275 3156
rect 5407 3152 5411 3156
rect 5543 3152 5547 3156
rect 5663 3153 5667 3157
rect 1975 3136 1979 3140
rect 2067 3137 2071 3141
rect 2267 3137 2271 3141
rect 2459 3137 2463 3141
rect 2651 3137 2655 3141
rect 2843 3137 2847 3141
rect 3027 3137 3031 3141
rect 3203 3137 3207 3141
rect 3387 3137 3391 3141
rect 3571 3137 3575 3141
rect 3799 3136 3803 3140
rect 3839 3136 3843 3140
rect 4835 3137 4839 3141
rect 4971 3137 4975 3141
rect 5107 3137 5111 3141
rect 5243 3137 5247 3141
rect 5379 3137 5383 3141
rect 5515 3137 5519 3141
rect 5663 3136 5667 3140
rect 111 3084 115 3088
rect 379 3083 383 3087
rect 563 3083 567 3087
rect 755 3083 759 3087
rect 955 3083 959 3087
rect 1163 3083 1167 3087
rect 1371 3083 1375 3087
rect 1935 3084 1939 3088
rect 111 3067 115 3071
rect 407 3068 411 3072
rect 591 3068 595 3072
rect 783 3068 787 3072
rect 983 3068 987 3072
rect 1191 3068 1195 3072
rect 1399 3068 1403 3072
rect 1935 3067 1939 3071
rect 111 2993 115 2997
rect 575 2992 579 2996
rect 799 2992 803 2996
rect 1047 2992 1051 2996
rect 1303 2992 1307 2996
rect 1567 2992 1571 2996
rect 1815 2992 1819 2996
rect 1935 2993 1939 2997
rect 1975 2992 1979 2996
rect 1995 2991 1999 2995
rect 2131 2991 2135 2995
rect 2267 2991 2271 2995
rect 2403 2991 2407 2995
rect 2539 2991 2543 2995
rect 2683 2991 2687 2995
rect 2835 2991 2839 2995
rect 2987 2991 2991 2995
rect 3139 2991 3143 2995
rect 3291 2991 3295 2995
rect 3799 2992 3803 2996
rect 3839 2992 3843 2996
rect 4483 2991 4487 2995
rect 4635 2991 4639 2995
rect 4803 2991 4807 2995
rect 4979 2991 4983 2995
rect 5163 2991 5167 2995
rect 5347 2991 5351 2995
rect 5515 2991 5519 2995
rect 5663 2992 5667 2996
rect 111 2976 115 2980
rect 547 2977 551 2981
rect 771 2977 775 2981
rect 1019 2977 1023 2981
rect 1275 2977 1279 2981
rect 1539 2977 1543 2981
rect 1787 2977 1791 2981
rect 1935 2976 1939 2980
rect 1975 2975 1979 2979
rect 2023 2976 2027 2980
rect 2159 2976 2163 2980
rect 2295 2976 2299 2980
rect 2431 2976 2435 2980
rect 2567 2976 2571 2980
rect 2711 2976 2715 2980
rect 2863 2976 2867 2980
rect 3015 2976 3019 2980
rect 3167 2976 3171 2980
rect 3319 2976 3323 2980
rect 3799 2975 3803 2979
rect 3839 2975 3843 2979
rect 4511 2976 4515 2980
rect 4663 2976 4667 2980
rect 4831 2976 4835 2980
rect 5007 2976 5011 2980
rect 5191 2976 5195 2980
rect 5375 2976 5379 2980
rect 5543 2976 5547 2980
rect 5663 2975 5667 2979
rect 1975 2917 1979 2921
rect 2023 2916 2027 2920
rect 2295 2916 2299 2920
rect 2591 2916 2595 2920
rect 2887 2916 2891 2920
rect 3183 2916 3187 2920
rect 3799 2917 3803 2921
rect 1975 2900 1979 2904
rect 1995 2901 1999 2905
rect 2267 2901 2271 2905
rect 2563 2901 2567 2905
rect 2859 2901 2863 2905
rect 3155 2901 3159 2905
rect 3799 2900 3803 2904
rect 3839 2893 3843 2897
rect 4047 2892 4051 2896
rect 4295 2892 4299 2896
rect 4583 2892 4587 2896
rect 4895 2892 4899 2896
rect 5231 2892 5235 2896
rect 5543 2892 5547 2896
rect 5663 2893 5667 2897
rect 3839 2876 3843 2880
rect 4019 2877 4023 2881
rect 4267 2877 4271 2881
rect 4555 2877 4559 2881
rect 4867 2877 4871 2881
rect 5203 2877 5207 2881
rect 5515 2877 5519 2881
rect 5663 2876 5667 2880
rect 111 2836 115 2840
rect 427 2835 431 2839
rect 563 2835 567 2839
rect 699 2835 703 2839
rect 835 2835 839 2839
rect 971 2835 975 2839
rect 1107 2835 1111 2839
rect 1243 2835 1247 2839
rect 1379 2835 1383 2839
rect 1515 2835 1519 2839
rect 1651 2835 1655 2839
rect 1787 2835 1791 2839
rect 1935 2836 1939 2840
rect 111 2819 115 2823
rect 455 2820 459 2824
rect 591 2820 595 2824
rect 727 2820 731 2824
rect 863 2820 867 2824
rect 999 2820 1003 2824
rect 1135 2820 1139 2824
rect 1271 2820 1275 2824
rect 1407 2820 1411 2824
rect 1543 2820 1547 2824
rect 1679 2820 1683 2824
rect 1815 2820 1819 2824
rect 1935 2819 1939 2823
rect 111 2753 115 2757
rect 463 2752 467 2756
rect 623 2752 627 2756
rect 783 2752 787 2756
rect 935 2752 939 2756
rect 1087 2752 1091 2756
rect 1239 2752 1243 2756
rect 1383 2752 1387 2756
rect 1535 2752 1539 2756
rect 1679 2752 1683 2756
rect 1815 2752 1819 2756
rect 1935 2753 1939 2757
rect 111 2736 115 2740
rect 435 2737 439 2741
rect 595 2737 599 2741
rect 755 2737 759 2741
rect 907 2737 911 2741
rect 1059 2737 1063 2741
rect 1211 2737 1215 2741
rect 1355 2737 1359 2741
rect 1507 2737 1511 2741
rect 1651 2737 1655 2741
rect 1787 2737 1791 2741
rect 1935 2736 1939 2740
rect 3839 2740 3843 2744
rect 3859 2739 3863 2743
rect 3995 2739 3999 2743
rect 4131 2739 4135 2743
rect 4267 2739 4271 2743
rect 4403 2739 4407 2743
rect 4539 2739 4543 2743
rect 4675 2739 4679 2743
rect 4811 2739 4815 2743
rect 5663 2740 5667 2744
rect 3839 2723 3843 2727
rect 3887 2724 3891 2728
rect 4023 2724 4027 2728
rect 4159 2724 4163 2728
rect 4295 2724 4299 2728
rect 4431 2724 4435 2728
rect 4567 2724 4571 2728
rect 4703 2724 4707 2728
rect 4839 2724 4843 2728
rect 5663 2723 5667 2727
rect 1975 2712 1979 2716
rect 3059 2711 3063 2715
rect 3195 2711 3199 2715
rect 3331 2711 3335 2715
rect 3799 2712 3803 2716
rect 1975 2695 1979 2699
rect 3087 2696 3091 2700
rect 3223 2696 3227 2700
rect 3359 2696 3363 2700
rect 3799 2695 3803 2699
rect 3839 2665 3843 2669
rect 4055 2664 4059 2668
rect 4303 2664 4307 2668
rect 4583 2664 4587 2668
rect 4895 2664 4899 2668
rect 5231 2664 5235 2668
rect 5543 2664 5547 2668
rect 5663 2665 5667 2669
rect 3839 2648 3843 2652
rect 4027 2649 4031 2653
rect 4275 2649 4279 2653
rect 4555 2649 4559 2653
rect 4867 2649 4871 2653
rect 5203 2649 5207 2653
rect 5515 2649 5519 2653
rect 5663 2648 5667 2652
rect 1975 2613 1979 2617
rect 3135 2612 3139 2616
rect 3271 2612 3275 2616
rect 3407 2612 3411 2616
rect 3543 2612 3547 2616
rect 3679 2612 3683 2616
rect 3799 2613 3803 2617
rect 111 2600 115 2604
rect 355 2599 359 2603
rect 539 2599 543 2603
rect 715 2599 719 2603
rect 883 2599 887 2603
rect 1043 2599 1047 2603
rect 1203 2599 1207 2603
rect 1355 2599 1359 2603
rect 1507 2599 1511 2603
rect 1651 2599 1655 2603
rect 1787 2599 1791 2603
rect 1935 2600 1939 2604
rect 1975 2596 1979 2600
rect 3107 2597 3111 2601
rect 3243 2597 3247 2601
rect 3379 2597 3383 2601
rect 3515 2597 3519 2601
rect 3651 2597 3655 2601
rect 3799 2596 3803 2600
rect 111 2583 115 2587
rect 383 2584 387 2588
rect 567 2584 571 2588
rect 743 2584 747 2588
rect 911 2584 915 2588
rect 1071 2584 1075 2588
rect 1231 2584 1235 2588
rect 1383 2584 1387 2588
rect 1535 2584 1539 2588
rect 1679 2584 1683 2588
rect 1815 2584 1819 2588
rect 1935 2583 1939 2587
rect 111 2525 115 2529
rect 231 2524 235 2528
rect 423 2524 427 2528
rect 623 2524 627 2528
rect 823 2524 827 2528
rect 1023 2524 1027 2528
rect 1223 2524 1227 2528
rect 1423 2524 1427 2528
rect 1631 2524 1635 2528
rect 1815 2524 1819 2528
rect 1935 2525 1939 2529
rect 111 2508 115 2512
rect 203 2509 207 2513
rect 395 2509 399 2513
rect 595 2509 599 2513
rect 795 2509 799 2513
rect 995 2509 999 2513
rect 1195 2509 1199 2513
rect 1395 2509 1399 2513
rect 1603 2509 1607 2513
rect 1787 2509 1791 2513
rect 1935 2508 1939 2512
rect 3839 2512 3843 2516
rect 4259 2511 4263 2515
rect 4475 2511 4479 2515
rect 4715 2511 4719 2515
rect 4979 2511 4983 2515
rect 5259 2511 5263 2515
rect 5515 2511 5519 2515
rect 5663 2512 5667 2516
rect 3839 2495 3843 2499
rect 4287 2496 4291 2500
rect 4503 2496 4507 2500
rect 4743 2496 4747 2500
rect 5007 2496 5011 2500
rect 5287 2496 5291 2500
rect 5543 2496 5547 2500
rect 5663 2495 5667 2499
rect 1975 2456 1979 2460
rect 1995 2455 1999 2459
rect 2235 2455 2239 2459
rect 2483 2455 2487 2459
rect 2715 2455 2719 2459
rect 2939 2455 2943 2459
rect 3155 2455 3159 2459
rect 3363 2455 3367 2459
rect 3579 2455 3583 2459
rect 3799 2456 3803 2460
rect 1975 2439 1979 2443
rect 2023 2440 2027 2444
rect 2263 2440 2267 2444
rect 2511 2440 2515 2444
rect 2743 2440 2747 2444
rect 2967 2440 2971 2444
rect 3183 2440 3187 2444
rect 3391 2440 3395 2444
rect 3607 2440 3611 2444
rect 3799 2439 3803 2443
rect 3839 2433 3843 2437
rect 4663 2432 4667 2436
rect 4847 2432 4851 2436
rect 5023 2432 5027 2436
rect 5199 2432 5203 2436
rect 5383 2432 5387 2436
rect 5543 2432 5547 2436
rect 5663 2433 5667 2437
rect 3839 2416 3843 2420
rect 4635 2417 4639 2421
rect 4819 2417 4823 2421
rect 4995 2417 4999 2421
rect 5171 2417 5175 2421
rect 5355 2417 5359 2421
rect 5515 2417 5519 2421
rect 5663 2416 5667 2420
rect 1975 2381 1979 2385
rect 2023 2380 2027 2384
rect 2159 2380 2163 2384
rect 2295 2380 2299 2384
rect 2431 2380 2435 2384
rect 2567 2380 2571 2384
rect 2711 2380 2715 2384
rect 2855 2380 2859 2384
rect 3007 2380 3011 2384
rect 3159 2380 3163 2384
rect 3311 2380 3315 2384
rect 3799 2381 3803 2385
rect 1975 2364 1979 2368
rect 1995 2365 1999 2369
rect 2131 2365 2135 2369
rect 2267 2365 2271 2369
rect 2403 2365 2407 2369
rect 2539 2365 2543 2369
rect 2683 2365 2687 2369
rect 2827 2365 2831 2369
rect 2979 2365 2983 2369
rect 3131 2365 3135 2369
rect 3283 2365 3287 2369
rect 3799 2364 3803 2368
rect 111 2356 115 2360
rect 219 2355 223 2359
rect 403 2355 407 2359
rect 595 2355 599 2359
rect 787 2355 791 2359
rect 979 2355 983 2359
rect 1935 2356 1939 2360
rect 111 2339 115 2343
rect 247 2340 251 2344
rect 431 2340 435 2344
rect 623 2340 627 2344
rect 815 2340 819 2344
rect 1007 2340 1011 2344
rect 1935 2339 1939 2343
rect 111 2277 115 2281
rect 399 2276 403 2280
rect 535 2276 539 2280
rect 671 2276 675 2280
rect 807 2276 811 2280
rect 943 2276 947 2280
rect 1935 2277 1939 2281
rect 3839 2280 3843 2284
rect 4675 2279 4679 2283
rect 4819 2279 4823 2283
rect 4963 2279 4967 2283
rect 5115 2279 5119 2283
rect 5267 2279 5271 2283
rect 5419 2279 5423 2283
rect 5663 2280 5667 2284
rect 111 2260 115 2264
rect 371 2261 375 2265
rect 507 2261 511 2265
rect 643 2261 647 2265
rect 779 2261 783 2265
rect 915 2261 919 2265
rect 1935 2260 1939 2264
rect 3839 2263 3843 2267
rect 4703 2264 4707 2268
rect 4847 2264 4851 2268
rect 4991 2264 4995 2268
rect 5143 2264 5147 2268
rect 5295 2264 5299 2268
rect 5447 2264 5451 2268
rect 5663 2263 5667 2267
rect 1975 2228 1979 2232
rect 2043 2227 2047 2231
rect 2179 2227 2183 2231
rect 2315 2227 2319 2231
rect 2451 2227 2455 2231
rect 2587 2227 2591 2231
rect 2723 2227 2727 2231
rect 2859 2227 2863 2231
rect 2995 2227 2999 2231
rect 3131 2227 3135 2231
rect 3799 2228 3803 2232
rect 1975 2211 1979 2215
rect 2071 2212 2075 2216
rect 2207 2212 2211 2216
rect 2343 2212 2347 2216
rect 2479 2212 2483 2216
rect 2615 2212 2619 2216
rect 2751 2212 2755 2216
rect 2887 2212 2891 2216
rect 3023 2212 3027 2216
rect 3159 2212 3163 2216
rect 3799 2211 3803 2215
rect 3839 2193 3843 2197
rect 3887 2192 3891 2196
rect 4167 2192 4171 2196
rect 4455 2192 4459 2196
rect 4719 2192 4723 2196
rect 4975 2192 4979 2196
rect 5231 2192 5235 2196
rect 5487 2192 5491 2196
rect 5663 2193 5667 2197
rect 3839 2176 3843 2180
rect 3859 2177 3863 2181
rect 4139 2177 4143 2181
rect 4427 2177 4431 2181
rect 4691 2177 4695 2181
rect 4947 2177 4951 2181
rect 5203 2177 5207 2181
rect 5459 2177 5463 2181
rect 5663 2176 5667 2180
rect 1975 2153 1979 2157
rect 2023 2152 2027 2156
rect 2239 2152 2243 2156
rect 2487 2152 2491 2156
rect 2727 2152 2731 2156
rect 2967 2152 2971 2156
rect 3207 2152 3211 2156
rect 3455 2152 3459 2156
rect 3679 2152 3683 2156
rect 3799 2153 3803 2157
rect 1975 2136 1979 2140
rect 1995 2137 1999 2141
rect 2211 2137 2215 2141
rect 2459 2137 2463 2141
rect 2699 2137 2703 2141
rect 2939 2137 2943 2141
rect 3179 2137 3183 2141
rect 3427 2137 3431 2141
rect 3651 2137 3655 2141
rect 3799 2136 3803 2140
rect 111 2120 115 2124
rect 323 2119 327 2123
rect 459 2119 463 2123
rect 595 2119 599 2123
rect 731 2119 735 2123
rect 867 2119 871 2123
rect 1935 2120 1939 2124
rect 111 2103 115 2107
rect 351 2104 355 2108
rect 487 2104 491 2108
rect 623 2104 627 2108
rect 759 2104 763 2108
rect 895 2104 899 2108
rect 1935 2103 1939 2107
rect 3839 2044 3843 2048
rect 3859 2043 3863 2047
rect 4083 2043 4087 2047
rect 4323 2043 4327 2047
rect 4547 2043 4551 2047
rect 4755 2043 4759 2047
rect 4947 2043 4951 2047
rect 5139 2043 5143 2047
rect 5323 2043 5327 2047
rect 5515 2043 5519 2047
rect 5663 2044 5667 2048
rect 3839 2027 3843 2031
rect 3887 2028 3891 2032
rect 4111 2028 4115 2032
rect 4351 2028 4355 2032
rect 4575 2028 4579 2032
rect 4783 2028 4787 2032
rect 4975 2028 4979 2032
rect 5167 2028 5171 2032
rect 5351 2028 5355 2032
rect 5543 2028 5547 2032
rect 5663 2027 5667 2031
rect 111 2013 115 2017
rect 319 2012 323 2016
rect 479 2012 483 2016
rect 663 2012 667 2016
rect 871 2012 875 2016
rect 1095 2012 1099 2016
rect 1335 2012 1339 2016
rect 1583 2012 1587 2016
rect 1815 2012 1819 2016
rect 1935 2013 1939 2017
rect 111 1996 115 2000
rect 291 1997 295 2001
rect 451 1997 455 2001
rect 635 1997 639 2001
rect 843 1997 847 2001
rect 1067 1997 1071 2001
rect 1307 1997 1311 2001
rect 1555 1997 1559 2001
rect 1787 1997 1791 2001
rect 1935 1996 1939 2000
rect 1975 1988 1979 1992
rect 1995 1987 1999 1991
rect 2211 1987 2215 1991
rect 2459 1987 2463 1991
rect 2707 1987 2711 1991
rect 2963 1987 2967 1991
rect 3219 1987 3223 1991
rect 3483 1987 3487 1991
rect 3799 1988 3803 1992
rect 1975 1971 1979 1975
rect 2023 1972 2027 1976
rect 2239 1972 2243 1976
rect 2487 1972 2491 1976
rect 2735 1972 2739 1976
rect 2991 1972 2995 1976
rect 3247 1972 3251 1976
rect 3511 1972 3515 1976
rect 3799 1971 3803 1975
rect 3839 1969 3843 1973
rect 3887 1968 3891 1972
rect 4167 1968 4171 1972
rect 4463 1968 4467 1972
rect 4743 1968 4747 1972
rect 5007 1968 5011 1972
rect 5271 1968 5275 1972
rect 5543 1968 5547 1972
rect 5663 1969 5667 1973
rect 3839 1952 3843 1956
rect 3859 1953 3863 1957
rect 4139 1953 4143 1957
rect 4435 1953 4439 1957
rect 4715 1953 4719 1957
rect 4979 1953 4983 1957
rect 5243 1953 5247 1957
rect 5515 1953 5519 1957
rect 5663 1952 5667 1956
rect 1975 1905 1979 1909
rect 2159 1904 2163 1908
rect 2439 1904 2443 1908
rect 2703 1904 2707 1908
rect 2959 1904 2963 1908
rect 3207 1904 3211 1908
rect 3455 1904 3459 1908
rect 3679 1904 3683 1908
rect 3799 1905 3803 1909
rect 1975 1888 1979 1892
rect 2131 1889 2135 1893
rect 2411 1889 2415 1893
rect 2675 1889 2679 1893
rect 2931 1889 2935 1893
rect 3179 1889 3183 1893
rect 3427 1889 3431 1893
rect 3651 1889 3655 1893
rect 3799 1888 3803 1892
rect 111 1856 115 1860
rect 187 1855 191 1859
rect 419 1855 423 1859
rect 651 1855 655 1859
rect 883 1855 887 1859
rect 1115 1855 1119 1859
rect 1347 1855 1351 1859
rect 1579 1855 1583 1859
rect 1787 1855 1791 1859
rect 1935 1856 1939 1860
rect 111 1839 115 1843
rect 215 1840 219 1844
rect 447 1840 451 1844
rect 679 1840 683 1844
rect 911 1840 915 1844
rect 1143 1840 1147 1844
rect 1375 1840 1379 1844
rect 1607 1840 1611 1844
rect 1815 1840 1819 1844
rect 1935 1839 1939 1843
rect 3839 1808 3843 1812
rect 4539 1807 4543 1811
rect 4723 1807 4727 1811
rect 4915 1807 4919 1811
rect 5115 1807 5119 1811
rect 5323 1807 5327 1811
rect 5515 1807 5519 1811
rect 5663 1808 5667 1812
rect 3839 1791 3843 1795
rect 4567 1792 4571 1796
rect 4751 1792 4755 1796
rect 4943 1792 4947 1796
rect 5143 1792 5147 1796
rect 5351 1792 5355 1796
rect 5543 1792 5547 1796
rect 5663 1791 5667 1795
rect 111 1769 115 1773
rect 159 1768 163 1772
rect 367 1768 371 1772
rect 591 1768 595 1772
rect 799 1768 803 1772
rect 999 1768 1003 1772
rect 1191 1768 1195 1772
rect 1375 1768 1379 1772
rect 1559 1768 1563 1772
rect 1751 1768 1755 1772
rect 1935 1769 1939 1773
rect 111 1752 115 1756
rect 131 1753 135 1757
rect 339 1753 343 1757
rect 563 1753 567 1757
rect 771 1753 775 1757
rect 971 1753 975 1757
rect 1163 1753 1167 1757
rect 1347 1753 1351 1757
rect 1531 1753 1535 1757
rect 1723 1753 1727 1757
rect 1935 1752 1939 1756
rect 1975 1748 1979 1752
rect 2307 1747 2311 1751
rect 2499 1747 2503 1751
rect 2691 1747 2695 1751
rect 2883 1747 2887 1751
rect 3067 1747 3071 1751
rect 3251 1747 3255 1751
rect 3443 1747 3447 1751
rect 3635 1747 3639 1751
rect 3799 1748 3803 1752
rect 1975 1731 1979 1735
rect 2335 1732 2339 1736
rect 2527 1732 2531 1736
rect 2719 1732 2723 1736
rect 2911 1732 2915 1736
rect 3095 1732 3099 1736
rect 3279 1732 3283 1736
rect 3471 1732 3475 1736
rect 3663 1732 3667 1736
rect 3799 1731 3803 1735
rect 3839 1725 3843 1729
rect 4383 1724 4387 1728
rect 4599 1724 4603 1728
rect 4831 1724 4835 1728
rect 5071 1724 5075 1728
rect 5319 1724 5323 1728
rect 5543 1724 5547 1728
rect 5663 1725 5667 1729
rect 3839 1708 3843 1712
rect 4355 1709 4359 1713
rect 4571 1709 4575 1713
rect 4803 1709 4807 1713
rect 5043 1709 5047 1713
rect 5291 1709 5295 1713
rect 5515 1709 5519 1713
rect 5663 1708 5667 1712
rect 1975 1673 1979 1677
rect 2471 1672 2475 1676
rect 2607 1672 2611 1676
rect 2743 1672 2747 1676
rect 2879 1672 2883 1676
rect 3023 1672 3027 1676
rect 3175 1672 3179 1676
rect 3327 1672 3331 1676
rect 3799 1673 3803 1677
rect 1975 1656 1979 1660
rect 2443 1657 2447 1661
rect 2579 1657 2583 1661
rect 2715 1657 2719 1661
rect 2851 1657 2855 1661
rect 2995 1657 2999 1661
rect 3147 1657 3151 1661
rect 3299 1657 3303 1661
rect 3799 1656 3803 1660
rect 111 1612 115 1616
rect 131 1611 135 1615
rect 355 1611 359 1615
rect 595 1611 599 1615
rect 835 1611 839 1615
rect 1067 1611 1071 1615
rect 1307 1611 1311 1615
rect 1547 1611 1551 1615
rect 1935 1612 1939 1616
rect 111 1595 115 1599
rect 159 1596 163 1600
rect 383 1596 387 1600
rect 623 1596 627 1600
rect 863 1596 867 1600
rect 1095 1596 1099 1600
rect 1335 1596 1339 1600
rect 1575 1596 1579 1600
rect 1935 1595 1939 1599
rect 3839 1564 3843 1568
rect 3907 1563 3911 1567
rect 4123 1563 4127 1567
rect 4363 1563 4367 1567
rect 4627 1563 4631 1567
rect 4907 1563 4911 1567
rect 5195 1563 5199 1567
rect 5491 1563 5495 1567
rect 5663 1564 5667 1568
rect 3839 1547 3843 1551
rect 3935 1548 3939 1552
rect 4151 1548 4155 1552
rect 4391 1548 4395 1552
rect 4655 1548 4659 1552
rect 4935 1548 4939 1552
rect 5223 1548 5227 1552
rect 5519 1548 5523 1552
rect 5663 1547 5667 1551
rect 111 1533 115 1537
rect 159 1532 163 1536
rect 359 1532 363 1536
rect 575 1532 579 1536
rect 783 1532 787 1536
rect 983 1532 987 1536
rect 1183 1532 1187 1536
rect 1375 1532 1379 1536
rect 1575 1532 1579 1536
rect 1935 1533 1939 1537
rect 1975 1524 1979 1528
rect 2355 1523 2359 1527
rect 2563 1523 2567 1527
rect 2779 1523 2783 1527
rect 3003 1523 3007 1527
rect 3227 1523 3231 1527
rect 3459 1523 3463 1527
rect 3799 1524 3803 1528
rect 111 1516 115 1520
rect 131 1517 135 1521
rect 331 1517 335 1521
rect 547 1517 551 1521
rect 755 1517 759 1521
rect 955 1517 959 1521
rect 1155 1517 1159 1521
rect 1347 1517 1351 1521
rect 1547 1517 1551 1521
rect 1935 1516 1939 1520
rect 1975 1507 1979 1511
rect 2383 1508 2387 1512
rect 2591 1508 2595 1512
rect 2807 1508 2811 1512
rect 3031 1508 3035 1512
rect 3255 1508 3259 1512
rect 3487 1508 3491 1512
rect 3799 1507 3803 1511
rect 3839 1489 3843 1493
rect 3887 1488 3891 1492
rect 4023 1488 4027 1492
rect 4159 1488 4163 1492
rect 4295 1488 4299 1492
rect 4479 1488 4483 1492
rect 4695 1488 4699 1492
rect 4935 1488 4939 1492
rect 5191 1488 5195 1492
rect 5447 1488 5451 1492
rect 5663 1489 5667 1493
rect 3839 1472 3843 1476
rect 3859 1473 3863 1477
rect 3995 1473 3999 1477
rect 4131 1473 4135 1477
rect 4267 1473 4271 1477
rect 4451 1473 4455 1477
rect 4667 1473 4671 1477
rect 4907 1473 4911 1477
rect 5163 1473 5167 1477
rect 5419 1473 5423 1477
rect 5663 1472 5667 1476
rect 1975 1449 1979 1453
rect 2023 1448 2027 1452
rect 2159 1448 2163 1452
rect 2327 1448 2331 1452
rect 2543 1448 2547 1452
rect 2799 1448 2803 1452
rect 3087 1448 3091 1452
rect 3391 1448 3395 1452
rect 3679 1448 3683 1452
rect 3799 1449 3803 1453
rect 1975 1432 1979 1436
rect 1995 1433 1999 1437
rect 2131 1433 2135 1437
rect 2299 1433 2303 1437
rect 2515 1433 2519 1437
rect 2771 1433 2775 1437
rect 3059 1433 3063 1437
rect 3363 1433 3367 1437
rect 3651 1433 3655 1437
rect 3799 1432 3803 1436
rect 111 1364 115 1368
rect 235 1363 239 1367
rect 507 1363 511 1367
rect 779 1363 783 1367
rect 1059 1363 1063 1367
rect 1339 1363 1343 1367
rect 1935 1364 1939 1368
rect 111 1347 115 1351
rect 263 1348 267 1352
rect 535 1348 539 1352
rect 807 1348 811 1352
rect 1087 1348 1091 1352
rect 1367 1348 1371 1352
rect 1935 1347 1939 1351
rect 3839 1328 3843 1332
rect 3859 1327 3863 1331
rect 3995 1327 3999 1331
rect 4147 1327 4151 1331
rect 4363 1327 4367 1331
rect 4611 1327 4615 1331
rect 4891 1327 4895 1331
rect 5195 1327 5199 1331
rect 5499 1327 5503 1331
rect 5663 1328 5667 1332
rect 3839 1311 3843 1315
rect 3887 1312 3891 1316
rect 4023 1312 4027 1316
rect 4175 1312 4179 1316
rect 4391 1312 4395 1316
rect 4639 1312 4643 1316
rect 4919 1312 4923 1316
rect 5223 1312 5227 1316
rect 5527 1312 5531 1316
rect 5663 1311 5667 1315
rect 1975 1300 1979 1304
rect 1995 1299 1999 1303
rect 2491 1299 2495 1303
rect 3019 1299 3023 1303
rect 3555 1299 3559 1303
rect 3799 1300 3803 1304
rect 111 1285 115 1289
rect 159 1284 163 1288
rect 383 1284 387 1288
rect 599 1284 603 1288
rect 799 1284 803 1288
rect 991 1284 995 1288
rect 1167 1284 1171 1288
rect 1335 1284 1339 1288
rect 1503 1284 1507 1288
rect 1671 1284 1675 1288
rect 1815 1284 1819 1288
rect 1935 1285 1939 1289
rect 1975 1283 1979 1287
rect 2023 1284 2027 1288
rect 2519 1284 2523 1288
rect 3047 1284 3051 1288
rect 3583 1284 3587 1288
rect 3799 1283 3803 1287
rect 111 1268 115 1272
rect 131 1269 135 1273
rect 355 1269 359 1273
rect 571 1269 575 1273
rect 771 1269 775 1273
rect 963 1269 967 1273
rect 1139 1269 1143 1273
rect 1307 1269 1311 1273
rect 1475 1269 1479 1273
rect 1643 1269 1647 1273
rect 1787 1269 1791 1273
rect 1935 1268 1939 1272
rect 3839 1253 3843 1257
rect 3887 1252 3891 1256
rect 4023 1252 4027 1256
rect 4167 1252 4171 1256
rect 4335 1252 4339 1256
rect 4511 1252 4515 1256
rect 4703 1252 4707 1256
rect 4903 1252 4907 1256
rect 5119 1252 5123 1256
rect 5343 1252 5347 1256
rect 5543 1252 5547 1256
rect 5663 1253 5667 1257
rect 3839 1236 3843 1240
rect 3859 1237 3863 1241
rect 3995 1237 3999 1241
rect 4139 1237 4143 1241
rect 4307 1237 4311 1241
rect 4483 1237 4487 1241
rect 4675 1237 4679 1241
rect 4875 1237 4879 1241
rect 5091 1237 5095 1241
rect 5315 1237 5319 1241
rect 5515 1237 5519 1241
rect 5663 1236 5667 1240
rect 1975 1161 1979 1165
rect 2743 1160 2747 1164
rect 3047 1160 3051 1164
rect 3359 1160 3363 1164
rect 3679 1160 3683 1164
rect 3799 1161 3803 1165
rect 1975 1144 1979 1148
rect 2715 1145 2719 1149
rect 3019 1145 3023 1149
rect 3331 1145 3335 1149
rect 3651 1145 3655 1149
rect 3799 1144 3803 1148
rect 111 1128 115 1132
rect 147 1127 151 1131
rect 323 1127 327 1131
rect 499 1127 503 1131
rect 675 1127 679 1131
rect 851 1127 855 1131
rect 1019 1127 1023 1131
rect 1179 1127 1183 1131
rect 1331 1127 1335 1131
rect 1483 1127 1487 1131
rect 1643 1127 1647 1131
rect 1787 1127 1791 1131
rect 1935 1128 1939 1132
rect 111 1111 115 1115
rect 175 1112 179 1116
rect 351 1112 355 1116
rect 527 1112 531 1116
rect 703 1112 707 1116
rect 879 1112 883 1116
rect 1047 1112 1051 1116
rect 1207 1112 1211 1116
rect 1359 1112 1363 1116
rect 1511 1112 1515 1116
rect 1671 1112 1675 1116
rect 1815 1112 1819 1116
rect 1935 1111 1939 1115
rect 3839 1100 3843 1104
rect 4811 1099 4815 1103
rect 4947 1099 4951 1103
rect 5083 1099 5087 1103
rect 5227 1099 5231 1103
rect 5379 1099 5383 1103
rect 5515 1099 5519 1103
rect 5663 1100 5667 1104
rect 3839 1083 3843 1087
rect 4839 1084 4843 1088
rect 4975 1084 4979 1088
rect 5111 1084 5115 1088
rect 5255 1084 5259 1088
rect 5407 1084 5411 1088
rect 5543 1084 5547 1088
rect 5663 1083 5667 1087
rect 111 1033 115 1037
rect 159 1032 163 1036
rect 447 1032 451 1036
rect 775 1032 779 1036
rect 1111 1032 1115 1036
rect 1455 1032 1459 1036
rect 1807 1032 1811 1036
rect 1935 1033 1939 1037
rect 111 1016 115 1020
rect 131 1017 135 1021
rect 419 1017 423 1021
rect 747 1017 751 1021
rect 1083 1017 1087 1021
rect 1427 1017 1431 1021
rect 3839 1021 3843 1025
rect 1779 1017 1783 1021
rect 4807 1020 4811 1024
rect 1935 1016 1939 1020
rect 4943 1020 4947 1024
rect 5079 1020 5083 1024
rect 5215 1020 5219 1024
rect 5351 1020 5355 1024
rect 5487 1020 5491 1024
rect 5663 1021 5667 1025
rect 1975 1012 1979 1016
rect 2243 1011 2247 1015
rect 2379 1011 2383 1015
rect 2523 1011 2527 1015
rect 2675 1011 2679 1015
rect 2827 1011 2831 1015
rect 2987 1011 2991 1015
rect 3155 1011 3159 1015
rect 3323 1011 3327 1015
rect 3499 1011 3503 1015
rect 3651 1011 3655 1015
rect 3799 1012 3803 1016
rect 3839 1004 3843 1008
rect 4779 1005 4783 1009
rect 4915 1005 4919 1009
rect 5051 1005 5055 1009
rect 5187 1005 5191 1009
rect 5323 1005 5327 1009
rect 5459 1005 5463 1009
rect 5663 1004 5667 1008
rect 1975 995 1979 999
rect 2271 996 2275 1000
rect 2407 996 2411 1000
rect 2551 996 2555 1000
rect 2703 996 2707 1000
rect 2855 996 2859 1000
rect 3015 996 3019 1000
rect 3183 996 3187 1000
rect 3351 996 3355 1000
rect 3527 996 3531 1000
rect 3679 996 3683 1000
rect 3799 995 3803 999
rect 1975 933 1979 937
rect 2279 932 2283 936
rect 2495 932 2499 936
rect 2711 932 2715 936
rect 2911 932 2915 936
rect 3103 932 3107 936
rect 3295 932 3299 936
rect 3479 932 3483 936
rect 3671 932 3675 936
rect 3799 933 3803 937
rect 1975 916 1979 920
rect 2251 917 2255 921
rect 2467 917 2471 921
rect 2683 917 2687 921
rect 2883 917 2887 921
rect 3075 917 3079 921
rect 3267 917 3271 921
rect 3451 917 3455 921
rect 3643 917 3647 921
rect 3799 916 3803 920
rect 111 880 115 884
rect 131 879 135 883
rect 339 879 343 883
rect 595 879 599 883
rect 875 879 879 883
rect 1179 879 1183 883
rect 1491 879 1495 883
rect 1787 879 1791 883
rect 1935 880 1939 884
rect 111 863 115 867
rect 159 864 163 868
rect 367 864 371 868
rect 623 864 627 868
rect 903 864 907 868
rect 1207 864 1211 868
rect 1519 864 1523 868
rect 3839 868 3843 872
rect 1815 864 1819 868
rect 4355 867 4359 871
rect 1935 863 1939 867
rect 4571 867 4575 871
rect 4803 867 4807 871
rect 5043 867 5047 871
rect 5291 867 5295 871
rect 5515 867 5519 871
rect 5663 868 5667 872
rect 3839 851 3843 855
rect 4383 852 4387 856
rect 4599 852 4603 856
rect 4831 852 4835 856
rect 5071 852 5075 856
rect 5319 852 5323 856
rect 5543 852 5547 856
rect 5663 851 5667 855
rect 111 793 115 797
rect 159 792 163 796
rect 383 792 387 796
rect 631 792 635 796
rect 887 792 891 796
rect 1143 792 1147 796
rect 1935 793 1939 797
rect 3839 789 3843 793
rect 3959 788 3963 792
rect 4207 788 4211 792
rect 4495 788 4499 792
rect 4815 788 4819 792
rect 5151 788 5155 792
rect 5487 788 5491 792
rect 5663 789 5667 793
rect 111 776 115 780
rect 131 777 135 781
rect 355 777 359 781
rect 603 777 607 781
rect 859 777 863 781
rect 1115 777 1119 781
rect 1935 776 1939 780
rect 1975 780 1979 784
rect 1995 779 1999 783
rect 2131 779 2135 783
rect 2283 779 2287 783
rect 2443 779 2447 783
rect 2603 779 2607 783
rect 2763 779 2767 783
rect 2923 779 2927 783
rect 3083 779 3087 783
rect 3243 779 3247 783
rect 3403 779 3407 783
rect 3799 780 3803 784
rect 3839 772 3843 776
rect 3931 773 3935 777
rect 4179 773 4183 777
rect 4467 773 4471 777
rect 4787 773 4791 777
rect 5123 773 5127 777
rect 5459 773 5463 777
rect 5663 772 5667 776
rect 1975 763 1979 767
rect 2023 764 2027 768
rect 2159 764 2163 768
rect 2311 764 2315 768
rect 2471 764 2475 768
rect 2631 764 2635 768
rect 2791 764 2795 768
rect 2951 764 2955 768
rect 3111 764 3115 768
rect 3271 764 3275 768
rect 3431 764 3435 768
rect 3799 763 3803 767
rect 1975 705 1979 709
rect 2183 704 2187 708
rect 2439 704 2443 708
rect 2679 704 2683 708
rect 2903 704 2907 708
rect 3111 704 3115 708
rect 3311 704 3315 708
rect 3503 704 3507 708
rect 3679 704 3683 708
rect 3799 705 3803 709
rect 1975 688 1979 692
rect 2155 689 2159 693
rect 2411 689 2415 693
rect 2651 689 2655 693
rect 2875 689 2879 693
rect 3083 689 3087 693
rect 3283 689 3287 693
rect 3475 689 3479 693
rect 3651 689 3655 693
rect 3799 688 3803 692
rect 111 644 115 648
rect 699 643 703 647
rect 835 643 839 647
rect 971 643 975 647
rect 1107 643 1111 647
rect 1243 643 1247 647
rect 1379 643 1383 647
rect 1515 643 1519 647
rect 1651 643 1655 647
rect 1787 643 1791 647
rect 1935 644 1939 648
rect 111 627 115 631
rect 727 628 731 632
rect 863 628 867 632
rect 999 628 1003 632
rect 1135 628 1139 632
rect 1271 628 1275 632
rect 1407 628 1411 632
rect 1543 628 1547 632
rect 1679 628 1683 632
rect 1815 628 1819 632
rect 1935 627 1939 631
rect 3839 628 3843 632
rect 3859 627 3863 631
rect 3995 627 3999 631
rect 4147 627 4151 631
rect 4355 627 4359 631
rect 4595 627 4599 631
rect 4867 627 4871 631
rect 5163 627 5167 631
rect 5459 627 5463 631
rect 5663 628 5667 632
rect 3839 611 3843 615
rect 3887 612 3891 616
rect 4023 612 4027 616
rect 4175 612 4179 616
rect 4383 612 4387 616
rect 4623 612 4627 616
rect 4895 612 4899 616
rect 5191 612 5195 616
rect 5487 612 5491 616
rect 5663 611 5667 615
rect 111 569 115 573
rect 159 568 163 572
rect 375 568 379 572
rect 599 568 603 572
rect 807 568 811 572
rect 999 568 1003 572
rect 1175 568 1179 572
rect 1343 568 1347 572
rect 1511 568 1515 572
rect 1671 568 1675 572
rect 1815 568 1819 572
rect 1935 569 1939 573
rect 111 552 115 556
rect 131 553 135 557
rect 347 553 351 557
rect 571 553 575 557
rect 779 553 783 557
rect 971 553 975 557
rect 1147 553 1151 557
rect 1315 553 1319 557
rect 1483 553 1487 557
rect 1643 553 1647 557
rect 1787 553 1791 557
rect 1935 552 1939 556
rect 3839 553 3843 557
rect 3887 552 3891 556
rect 4023 552 4027 556
rect 4159 552 4163 556
rect 4295 552 4299 556
rect 4431 552 4435 556
rect 4567 552 4571 556
rect 4711 552 4715 556
rect 4879 552 4883 556
rect 5063 552 5067 556
rect 5255 552 5259 556
rect 5447 552 5451 556
rect 5663 553 5667 557
rect 3839 536 3843 540
rect 3859 537 3863 541
rect 3995 537 3999 541
rect 4131 537 4135 541
rect 4267 537 4271 541
rect 4403 537 4407 541
rect 4539 537 4543 541
rect 4683 537 4687 541
rect 4851 537 4855 541
rect 5035 537 5039 541
rect 5227 537 5231 541
rect 5419 537 5423 541
rect 5663 536 5667 540
rect 111 420 115 424
rect 131 419 135 423
rect 355 419 359 423
rect 603 419 607 423
rect 843 419 847 423
rect 1083 419 1087 423
rect 1323 419 1327 423
rect 1563 419 1567 423
rect 1787 419 1791 423
rect 1935 420 1939 424
rect 111 403 115 407
rect 159 404 163 408
rect 383 404 387 408
rect 631 404 635 408
rect 871 404 875 408
rect 1111 404 1115 408
rect 1351 404 1355 408
rect 1591 404 1595 408
rect 1815 404 1819 408
rect 1935 403 1939 407
rect 3839 404 3843 408
rect 3859 403 3863 407
rect 4115 403 4119 407
rect 4395 403 4399 407
rect 4675 403 4679 407
rect 4947 403 4951 407
rect 5227 403 5231 407
rect 5507 403 5511 407
rect 5663 404 5667 408
rect 3839 387 3843 391
rect 3887 388 3891 392
rect 4143 388 4147 392
rect 4423 388 4427 392
rect 4703 388 4707 392
rect 4975 388 4979 392
rect 5255 388 5259 392
rect 5535 388 5539 392
rect 5663 387 5667 391
rect 1975 380 1979 384
rect 1995 379 1999 383
rect 2251 379 2255 383
rect 2523 379 2527 383
rect 2771 379 2775 383
rect 3003 379 3007 383
rect 3227 379 3231 383
rect 3451 379 3455 383
rect 3651 379 3655 383
rect 3799 380 3803 384
rect 1975 363 1979 367
rect 2023 364 2027 368
rect 2279 364 2283 368
rect 2551 364 2555 368
rect 2799 364 2803 368
rect 3031 364 3035 368
rect 3255 364 3259 368
rect 3479 364 3483 368
rect 3679 364 3683 368
rect 3799 363 3803 367
rect 111 329 115 333
rect 159 328 163 332
rect 303 328 307 332
rect 479 328 483 332
rect 655 328 659 332
rect 831 328 835 332
rect 1935 329 1939 333
rect 3839 321 3843 325
rect 4727 320 4731 324
rect 4895 320 4899 324
rect 5063 320 5067 324
rect 5231 320 5235 324
rect 5399 320 5403 324
rect 5543 320 5547 324
rect 5663 321 5667 325
rect 111 312 115 316
rect 131 313 135 317
rect 275 313 279 317
rect 451 313 455 317
rect 627 313 631 317
rect 803 313 807 317
rect 1935 312 1939 316
rect 1975 301 1979 305
rect 2023 300 2027 304
rect 2159 300 2163 304
rect 2295 300 2299 304
rect 2431 300 2435 304
rect 2567 300 2571 304
rect 2703 300 2707 304
rect 2839 300 2843 304
rect 2975 300 2979 304
rect 3111 300 3115 304
rect 3247 300 3251 304
rect 3383 300 3387 304
rect 3519 300 3523 304
rect 3655 300 3659 304
rect 3799 301 3803 305
rect 3839 304 3843 308
rect 4699 305 4703 309
rect 4867 305 4871 309
rect 5035 305 5039 309
rect 5203 305 5207 309
rect 5371 305 5375 309
rect 5515 305 5519 309
rect 5663 304 5667 308
rect 1975 284 1979 288
rect 1995 285 1999 289
rect 2131 285 2135 289
rect 2267 285 2271 289
rect 2403 285 2407 289
rect 2539 285 2543 289
rect 2675 285 2679 289
rect 2811 285 2815 289
rect 2947 285 2951 289
rect 3083 285 3087 289
rect 3219 285 3223 289
rect 3355 285 3359 289
rect 3491 285 3495 289
rect 3627 285 3631 289
rect 3799 284 3803 288
rect 111 140 115 144
rect 131 139 135 143
rect 267 139 271 143
rect 403 139 407 143
rect 539 139 543 143
rect 675 139 679 143
rect 811 139 815 143
rect 947 139 951 143
rect 1083 139 1087 143
rect 1935 140 1939 144
rect 3839 132 3843 136
rect 4291 131 4295 135
rect 4427 131 4431 135
rect 4563 131 4567 135
rect 4699 131 4703 135
rect 4835 131 4839 135
rect 4971 131 4975 135
rect 5107 131 5111 135
rect 5243 131 5247 135
rect 5379 131 5383 135
rect 5515 131 5519 135
rect 5663 132 5667 136
rect 111 123 115 127
rect 159 124 163 128
rect 295 124 299 128
rect 431 124 435 128
rect 567 124 571 128
rect 703 124 707 128
rect 839 124 843 128
rect 975 124 979 128
rect 1111 124 1115 128
rect 1935 123 1939 127
rect 1975 120 1979 124
rect 1995 119 1999 123
rect 2131 119 2135 123
rect 2267 119 2271 123
rect 2403 119 2407 123
rect 2539 119 2543 123
rect 2675 119 2679 123
rect 2811 119 2815 123
rect 2947 119 2951 123
rect 3083 119 3087 123
rect 3219 119 3223 123
rect 3355 119 3359 123
rect 3491 119 3495 123
rect 3627 119 3631 123
rect 3799 120 3803 124
rect 3839 115 3843 119
rect 4319 116 4323 120
rect 4455 116 4459 120
rect 4591 116 4595 120
rect 4727 116 4731 120
rect 4863 116 4867 120
rect 4999 116 5003 120
rect 5135 116 5139 120
rect 5271 116 5275 120
rect 5407 116 5411 120
rect 5543 116 5547 120
rect 5663 115 5667 119
rect 1975 103 1979 107
rect 2023 104 2027 108
rect 2159 104 2163 108
rect 2295 104 2299 108
rect 2431 104 2435 108
rect 2567 104 2571 108
rect 2703 104 2707 108
rect 2839 104 2843 108
rect 2975 104 2979 108
rect 3111 104 3115 108
rect 3247 104 3251 108
rect 3383 104 3387 108
rect 3519 104 3523 108
rect 3655 104 3659 108
rect 3799 103 3803 107
<< m3 >>
rect 1975 5758 1979 5759
rect 1975 5753 1979 5754
rect 2375 5758 2379 5759
rect 2375 5753 2379 5754
rect 2511 5758 2515 5759
rect 2511 5753 2515 5754
rect 2655 5758 2659 5759
rect 2655 5753 2659 5754
rect 2807 5758 2811 5759
rect 2807 5753 2811 5754
rect 2959 5758 2963 5759
rect 2959 5753 2963 5754
rect 3119 5758 3123 5759
rect 3119 5753 3123 5754
rect 3799 5758 3803 5759
rect 3799 5753 3803 5754
rect 1976 5730 1978 5753
rect 1974 5729 1980 5730
rect 2376 5729 2378 5753
rect 2512 5729 2514 5753
rect 2656 5729 2658 5753
rect 2808 5729 2810 5753
rect 2960 5729 2962 5753
rect 3120 5729 3122 5753
rect 3800 5730 3802 5753
rect 3798 5729 3804 5730
rect 1974 5725 1975 5729
rect 1979 5725 1980 5729
rect 1974 5724 1980 5725
rect 2374 5728 2380 5729
rect 2374 5724 2375 5728
rect 2379 5724 2380 5728
rect 2374 5723 2380 5724
rect 2510 5728 2516 5729
rect 2510 5724 2511 5728
rect 2515 5724 2516 5728
rect 2510 5723 2516 5724
rect 2654 5728 2660 5729
rect 2654 5724 2655 5728
rect 2659 5724 2660 5728
rect 2654 5723 2660 5724
rect 2806 5728 2812 5729
rect 2806 5724 2807 5728
rect 2811 5724 2812 5728
rect 2806 5723 2812 5724
rect 2958 5728 2964 5729
rect 2958 5724 2959 5728
rect 2963 5724 2964 5728
rect 2958 5723 2964 5724
rect 3118 5728 3124 5729
rect 3118 5724 3119 5728
rect 3123 5724 3124 5728
rect 3798 5725 3799 5729
rect 3803 5725 3804 5729
rect 3798 5724 3804 5725
rect 3118 5723 3124 5724
rect 111 5718 115 5719
rect 111 5713 115 5714
rect 159 5718 163 5719
rect 159 5713 163 5714
rect 295 5718 299 5719
rect 295 5713 299 5714
rect 431 5718 435 5719
rect 431 5713 435 5714
rect 567 5718 571 5719
rect 567 5713 571 5714
rect 703 5718 707 5719
rect 703 5713 707 5714
rect 839 5718 843 5719
rect 839 5713 843 5714
rect 975 5718 979 5719
rect 975 5713 979 5714
rect 1935 5718 1939 5719
rect 1935 5713 1939 5714
rect 2346 5713 2352 5714
rect 112 5690 114 5713
rect 110 5689 116 5690
rect 160 5689 162 5713
rect 296 5689 298 5713
rect 432 5689 434 5713
rect 568 5689 570 5713
rect 704 5689 706 5713
rect 840 5689 842 5713
rect 976 5689 978 5713
rect 1936 5690 1938 5713
rect 1974 5712 1980 5713
rect 1974 5708 1975 5712
rect 1979 5708 1980 5712
rect 2346 5709 2347 5713
rect 2351 5709 2352 5713
rect 2346 5708 2352 5709
rect 2482 5713 2488 5714
rect 2482 5709 2483 5713
rect 2487 5709 2488 5713
rect 2482 5708 2488 5709
rect 2626 5713 2632 5714
rect 2626 5709 2627 5713
rect 2631 5709 2632 5713
rect 2626 5708 2632 5709
rect 2778 5713 2784 5714
rect 2778 5709 2779 5713
rect 2783 5709 2784 5713
rect 2778 5708 2784 5709
rect 2930 5713 2936 5714
rect 2930 5709 2931 5713
rect 2935 5709 2936 5713
rect 2930 5708 2936 5709
rect 3090 5713 3096 5714
rect 3090 5709 3091 5713
rect 3095 5709 3096 5713
rect 3090 5708 3096 5709
rect 3798 5712 3804 5713
rect 3798 5708 3799 5712
rect 3803 5708 3804 5712
rect 1974 5707 1980 5708
rect 1934 5689 1940 5690
rect 110 5685 111 5689
rect 115 5685 116 5689
rect 110 5684 116 5685
rect 158 5688 164 5689
rect 158 5684 159 5688
rect 163 5684 164 5688
rect 158 5683 164 5684
rect 294 5688 300 5689
rect 294 5684 295 5688
rect 299 5684 300 5688
rect 294 5683 300 5684
rect 430 5688 436 5689
rect 430 5684 431 5688
rect 435 5684 436 5688
rect 430 5683 436 5684
rect 566 5688 572 5689
rect 566 5684 567 5688
rect 571 5684 572 5688
rect 566 5683 572 5684
rect 702 5688 708 5689
rect 702 5684 703 5688
rect 707 5684 708 5688
rect 702 5683 708 5684
rect 838 5688 844 5689
rect 838 5684 839 5688
rect 843 5684 844 5688
rect 838 5683 844 5684
rect 974 5688 980 5689
rect 974 5684 975 5688
rect 979 5684 980 5688
rect 1934 5685 1935 5689
rect 1939 5685 1940 5689
rect 1934 5684 1940 5685
rect 974 5683 980 5684
rect 130 5673 136 5674
rect 110 5672 116 5673
rect 110 5668 111 5672
rect 115 5668 116 5672
rect 130 5669 131 5673
rect 135 5669 136 5673
rect 130 5668 136 5669
rect 266 5673 272 5674
rect 266 5669 267 5673
rect 271 5669 272 5673
rect 266 5668 272 5669
rect 402 5673 408 5674
rect 402 5669 403 5673
rect 407 5669 408 5673
rect 402 5668 408 5669
rect 538 5673 544 5674
rect 538 5669 539 5673
rect 543 5669 544 5673
rect 538 5668 544 5669
rect 674 5673 680 5674
rect 674 5669 675 5673
rect 679 5669 680 5673
rect 674 5668 680 5669
rect 810 5673 816 5674
rect 810 5669 811 5673
rect 815 5669 816 5673
rect 810 5668 816 5669
rect 946 5673 952 5674
rect 946 5669 947 5673
rect 951 5669 952 5673
rect 946 5668 952 5669
rect 1934 5672 1940 5673
rect 1934 5668 1935 5672
rect 1939 5668 1940 5672
rect 110 5667 116 5668
rect 112 5579 114 5667
rect 132 5579 134 5668
rect 268 5579 270 5668
rect 404 5579 406 5668
rect 540 5579 542 5668
rect 676 5579 678 5668
rect 812 5579 814 5668
rect 948 5579 950 5668
rect 1934 5667 1940 5668
rect 1936 5579 1938 5667
rect 1976 5647 1978 5707
rect 2348 5647 2350 5708
rect 2484 5647 2486 5708
rect 2628 5647 2630 5708
rect 2780 5647 2782 5708
rect 2932 5647 2934 5708
rect 3092 5647 3094 5708
rect 3798 5707 3804 5708
rect 3800 5647 3802 5707
rect 3839 5682 3843 5683
rect 3839 5677 3843 5678
rect 4335 5682 4339 5683
rect 4335 5677 4339 5678
rect 4471 5682 4475 5683
rect 4471 5677 4475 5678
rect 4607 5682 4611 5683
rect 4607 5677 4611 5678
rect 4743 5682 4747 5683
rect 4743 5677 4747 5678
rect 4879 5682 4883 5683
rect 4879 5677 4883 5678
rect 5015 5682 5019 5683
rect 5015 5677 5019 5678
rect 5663 5682 5667 5683
rect 5663 5677 5667 5678
rect 3840 5654 3842 5677
rect 3838 5653 3844 5654
rect 4336 5653 4338 5677
rect 4472 5653 4474 5677
rect 4608 5653 4610 5677
rect 4744 5653 4746 5677
rect 4880 5653 4882 5677
rect 5016 5653 5018 5677
rect 5664 5654 5666 5677
rect 5662 5653 5668 5654
rect 3838 5649 3839 5653
rect 3843 5649 3844 5653
rect 3838 5648 3844 5649
rect 4334 5652 4340 5653
rect 4334 5648 4335 5652
rect 4339 5648 4340 5652
rect 4334 5647 4340 5648
rect 4470 5652 4476 5653
rect 4470 5648 4471 5652
rect 4475 5648 4476 5652
rect 4470 5647 4476 5648
rect 4606 5652 4612 5653
rect 4606 5648 4607 5652
rect 4611 5648 4612 5652
rect 4606 5647 4612 5648
rect 4742 5652 4748 5653
rect 4742 5648 4743 5652
rect 4747 5648 4748 5652
rect 4742 5647 4748 5648
rect 4878 5652 4884 5653
rect 4878 5648 4879 5652
rect 4883 5648 4884 5652
rect 4878 5647 4884 5648
rect 5014 5652 5020 5653
rect 5014 5648 5015 5652
rect 5019 5648 5020 5652
rect 5662 5649 5663 5653
rect 5667 5649 5668 5653
rect 5662 5648 5668 5649
rect 5014 5647 5020 5648
rect 1975 5646 1979 5647
rect 1975 5641 1979 5642
rect 1995 5646 1999 5647
rect 1995 5641 1999 5642
rect 2203 5646 2207 5647
rect 2203 5641 2207 5642
rect 2347 5646 2351 5647
rect 2347 5641 2351 5642
rect 2427 5646 2431 5647
rect 2427 5641 2431 5642
rect 2483 5646 2487 5647
rect 2483 5641 2487 5642
rect 2627 5646 2631 5647
rect 2627 5641 2631 5642
rect 2651 5646 2655 5647
rect 2651 5641 2655 5642
rect 2779 5646 2783 5647
rect 2779 5641 2783 5642
rect 2867 5646 2871 5647
rect 2867 5641 2871 5642
rect 2931 5646 2935 5647
rect 2931 5641 2935 5642
rect 3075 5646 3079 5647
rect 3075 5641 3079 5642
rect 3091 5646 3095 5647
rect 3091 5641 3095 5642
rect 3275 5646 3279 5647
rect 3275 5641 3279 5642
rect 3475 5646 3479 5647
rect 3475 5641 3479 5642
rect 3651 5646 3655 5647
rect 3651 5641 3655 5642
rect 3799 5646 3803 5647
rect 3799 5641 3803 5642
rect 1976 5581 1978 5641
rect 1974 5580 1980 5581
rect 1996 5580 1998 5641
rect 2204 5580 2206 5641
rect 2428 5580 2430 5641
rect 2652 5580 2654 5641
rect 2868 5580 2870 5641
rect 3076 5580 3078 5641
rect 3276 5580 3278 5641
rect 3476 5580 3478 5641
rect 3652 5580 3654 5641
rect 3800 5581 3802 5641
rect 4306 5637 4312 5638
rect 3838 5636 3844 5637
rect 3838 5632 3839 5636
rect 3843 5632 3844 5636
rect 4306 5633 4307 5637
rect 4311 5633 4312 5637
rect 4306 5632 4312 5633
rect 4442 5637 4448 5638
rect 4442 5633 4443 5637
rect 4447 5633 4448 5637
rect 4442 5632 4448 5633
rect 4578 5637 4584 5638
rect 4578 5633 4579 5637
rect 4583 5633 4584 5637
rect 4578 5632 4584 5633
rect 4714 5637 4720 5638
rect 4714 5633 4715 5637
rect 4719 5633 4720 5637
rect 4714 5632 4720 5633
rect 4850 5637 4856 5638
rect 4850 5633 4851 5637
rect 4855 5633 4856 5637
rect 4850 5632 4856 5633
rect 4986 5637 4992 5638
rect 4986 5633 4987 5637
rect 4991 5633 4992 5637
rect 4986 5632 4992 5633
rect 5662 5636 5668 5637
rect 5662 5632 5663 5636
rect 5667 5632 5668 5636
rect 3838 5631 3844 5632
rect 3798 5580 3804 5581
rect 111 5578 115 5579
rect 111 5573 115 5574
rect 131 5578 135 5579
rect 131 5573 135 5574
rect 267 5578 271 5579
rect 267 5573 271 5574
rect 403 5578 407 5579
rect 403 5573 407 5574
rect 539 5578 543 5579
rect 539 5573 543 5574
rect 619 5578 623 5579
rect 619 5573 623 5574
rect 675 5578 679 5579
rect 675 5573 679 5574
rect 755 5578 759 5579
rect 755 5573 759 5574
rect 811 5578 815 5579
rect 811 5573 815 5574
rect 899 5578 903 5579
rect 899 5573 903 5574
rect 947 5578 951 5579
rect 947 5573 951 5574
rect 1051 5578 1055 5579
rect 1051 5573 1055 5574
rect 1203 5578 1207 5579
rect 1203 5573 1207 5574
rect 1355 5578 1359 5579
rect 1355 5573 1359 5574
rect 1507 5578 1511 5579
rect 1507 5573 1511 5574
rect 1651 5578 1655 5579
rect 1651 5573 1655 5574
rect 1787 5578 1791 5579
rect 1787 5573 1791 5574
rect 1935 5578 1939 5579
rect 1974 5576 1975 5580
rect 1979 5576 1980 5580
rect 1974 5575 1980 5576
rect 1994 5579 2000 5580
rect 1994 5575 1995 5579
rect 1999 5575 2000 5579
rect 1994 5574 2000 5575
rect 2202 5579 2208 5580
rect 2202 5575 2203 5579
rect 2207 5575 2208 5579
rect 2202 5574 2208 5575
rect 2426 5579 2432 5580
rect 2426 5575 2427 5579
rect 2431 5575 2432 5579
rect 2426 5574 2432 5575
rect 2650 5579 2656 5580
rect 2650 5575 2651 5579
rect 2655 5575 2656 5579
rect 2650 5574 2656 5575
rect 2866 5579 2872 5580
rect 2866 5575 2867 5579
rect 2871 5575 2872 5579
rect 2866 5574 2872 5575
rect 3074 5579 3080 5580
rect 3074 5575 3075 5579
rect 3079 5575 3080 5579
rect 3074 5574 3080 5575
rect 3274 5579 3280 5580
rect 3274 5575 3275 5579
rect 3279 5575 3280 5579
rect 3274 5574 3280 5575
rect 3474 5579 3480 5580
rect 3474 5575 3475 5579
rect 3479 5575 3480 5579
rect 3474 5574 3480 5575
rect 3650 5579 3656 5580
rect 3650 5575 3651 5579
rect 3655 5575 3656 5579
rect 3798 5576 3799 5580
rect 3803 5576 3804 5580
rect 3798 5575 3804 5576
rect 3650 5574 3656 5575
rect 1935 5573 1939 5574
rect 112 5513 114 5573
rect 110 5512 116 5513
rect 620 5512 622 5573
rect 756 5512 758 5573
rect 900 5512 902 5573
rect 1052 5512 1054 5573
rect 1204 5512 1206 5573
rect 1356 5512 1358 5573
rect 1508 5512 1510 5573
rect 1652 5512 1654 5573
rect 1788 5512 1790 5573
rect 1936 5513 1938 5573
rect 3840 5571 3842 5631
rect 4308 5571 4310 5632
rect 4444 5571 4446 5632
rect 4580 5571 4582 5632
rect 4716 5571 4718 5632
rect 4852 5571 4854 5632
rect 4988 5571 4990 5632
rect 5662 5631 5668 5632
rect 5664 5571 5666 5631
rect 3839 5570 3843 5571
rect 3839 5565 3843 5566
rect 4211 5570 4215 5571
rect 4211 5565 4215 5566
rect 4307 5570 4311 5571
rect 4307 5565 4311 5566
rect 4403 5570 4407 5571
rect 4403 5565 4407 5566
rect 4443 5570 4447 5571
rect 4443 5565 4447 5566
rect 4579 5570 4583 5571
rect 4579 5565 4583 5566
rect 4595 5570 4599 5571
rect 4595 5565 4599 5566
rect 4715 5570 4719 5571
rect 4715 5565 4719 5566
rect 4795 5570 4799 5571
rect 4795 5565 4799 5566
rect 4851 5570 4855 5571
rect 4851 5565 4855 5566
rect 4987 5570 4991 5571
rect 4987 5565 4991 5566
rect 4995 5570 4999 5571
rect 4995 5565 4999 5566
rect 5195 5570 5199 5571
rect 5195 5565 5199 5566
rect 5663 5570 5667 5571
rect 5663 5565 5667 5566
rect 2022 5564 2028 5565
rect 1974 5563 1980 5564
rect 1974 5559 1975 5563
rect 1979 5559 1980 5563
rect 2022 5560 2023 5564
rect 2027 5560 2028 5564
rect 2022 5559 2028 5560
rect 2230 5564 2236 5565
rect 2230 5560 2231 5564
rect 2235 5560 2236 5564
rect 2230 5559 2236 5560
rect 2454 5564 2460 5565
rect 2454 5560 2455 5564
rect 2459 5560 2460 5564
rect 2454 5559 2460 5560
rect 2678 5564 2684 5565
rect 2678 5560 2679 5564
rect 2683 5560 2684 5564
rect 2678 5559 2684 5560
rect 2894 5564 2900 5565
rect 2894 5560 2895 5564
rect 2899 5560 2900 5564
rect 2894 5559 2900 5560
rect 3102 5564 3108 5565
rect 3102 5560 3103 5564
rect 3107 5560 3108 5564
rect 3102 5559 3108 5560
rect 3302 5564 3308 5565
rect 3302 5560 3303 5564
rect 3307 5560 3308 5564
rect 3302 5559 3308 5560
rect 3502 5564 3508 5565
rect 3502 5560 3503 5564
rect 3507 5560 3508 5564
rect 3502 5559 3508 5560
rect 3678 5564 3684 5565
rect 3678 5560 3679 5564
rect 3683 5560 3684 5564
rect 3678 5559 3684 5560
rect 3798 5563 3804 5564
rect 3798 5559 3799 5563
rect 3803 5559 3804 5563
rect 1974 5558 1980 5559
rect 1976 5535 1978 5558
rect 2024 5535 2026 5559
rect 2232 5535 2234 5559
rect 2456 5535 2458 5559
rect 2680 5535 2682 5559
rect 2896 5535 2898 5559
rect 3104 5535 3106 5559
rect 3304 5535 3306 5559
rect 3504 5535 3506 5559
rect 3680 5535 3682 5559
rect 3798 5558 3804 5559
rect 3800 5535 3802 5558
rect 1975 5534 1979 5535
rect 1975 5529 1979 5530
rect 2023 5534 2027 5535
rect 2023 5529 2027 5530
rect 2231 5534 2235 5535
rect 2231 5529 2235 5530
rect 2455 5534 2459 5535
rect 2455 5529 2459 5530
rect 2679 5534 2683 5535
rect 2679 5529 2683 5530
rect 2895 5534 2899 5535
rect 2895 5529 2899 5530
rect 2951 5534 2955 5535
rect 2951 5529 2955 5530
rect 3103 5534 3107 5535
rect 3103 5529 3107 5530
rect 3255 5534 3259 5535
rect 3255 5529 3259 5530
rect 3303 5534 3307 5535
rect 3303 5529 3307 5530
rect 3415 5534 3419 5535
rect 3415 5529 3419 5530
rect 3503 5534 3507 5535
rect 3503 5529 3507 5530
rect 3679 5534 3683 5535
rect 3679 5529 3683 5530
rect 3799 5534 3803 5535
rect 3799 5529 3803 5530
rect 1934 5512 1940 5513
rect 110 5508 111 5512
rect 115 5508 116 5512
rect 110 5507 116 5508
rect 618 5511 624 5512
rect 618 5507 619 5511
rect 623 5507 624 5511
rect 618 5506 624 5507
rect 754 5511 760 5512
rect 754 5507 755 5511
rect 759 5507 760 5511
rect 754 5506 760 5507
rect 898 5511 904 5512
rect 898 5507 899 5511
rect 903 5507 904 5511
rect 898 5506 904 5507
rect 1050 5511 1056 5512
rect 1050 5507 1051 5511
rect 1055 5507 1056 5511
rect 1050 5506 1056 5507
rect 1202 5511 1208 5512
rect 1202 5507 1203 5511
rect 1207 5507 1208 5511
rect 1202 5506 1208 5507
rect 1354 5511 1360 5512
rect 1354 5507 1355 5511
rect 1359 5507 1360 5511
rect 1354 5506 1360 5507
rect 1506 5511 1512 5512
rect 1506 5507 1507 5511
rect 1511 5507 1512 5511
rect 1506 5506 1512 5507
rect 1650 5511 1656 5512
rect 1650 5507 1651 5511
rect 1655 5507 1656 5511
rect 1650 5506 1656 5507
rect 1786 5511 1792 5512
rect 1786 5507 1787 5511
rect 1791 5507 1792 5511
rect 1934 5508 1935 5512
rect 1939 5508 1940 5512
rect 1934 5507 1940 5508
rect 1786 5506 1792 5507
rect 1976 5506 1978 5529
rect 1974 5505 1980 5506
rect 2952 5505 2954 5529
rect 3104 5505 3106 5529
rect 3256 5505 3258 5529
rect 3416 5505 3418 5529
rect 3800 5506 3802 5529
rect 3798 5505 3804 5506
rect 3840 5505 3842 5565
rect 1974 5501 1975 5505
rect 1979 5501 1980 5505
rect 1974 5500 1980 5501
rect 2950 5504 2956 5505
rect 2950 5500 2951 5504
rect 2955 5500 2956 5504
rect 2950 5499 2956 5500
rect 3102 5504 3108 5505
rect 3102 5500 3103 5504
rect 3107 5500 3108 5504
rect 3102 5499 3108 5500
rect 3254 5504 3260 5505
rect 3254 5500 3255 5504
rect 3259 5500 3260 5504
rect 3254 5499 3260 5500
rect 3414 5504 3420 5505
rect 3414 5500 3415 5504
rect 3419 5500 3420 5504
rect 3798 5501 3799 5505
rect 3803 5501 3804 5505
rect 3798 5500 3804 5501
rect 3838 5504 3844 5505
rect 4212 5504 4214 5565
rect 4404 5504 4406 5565
rect 4596 5504 4598 5565
rect 4796 5504 4798 5565
rect 4996 5504 4998 5565
rect 5196 5504 5198 5565
rect 5664 5505 5666 5565
rect 5662 5504 5668 5505
rect 3838 5500 3839 5504
rect 3843 5500 3844 5504
rect 3414 5499 3420 5500
rect 3838 5499 3844 5500
rect 4210 5503 4216 5504
rect 4210 5499 4211 5503
rect 4215 5499 4216 5503
rect 4210 5498 4216 5499
rect 4402 5503 4408 5504
rect 4402 5499 4403 5503
rect 4407 5499 4408 5503
rect 4402 5498 4408 5499
rect 4594 5503 4600 5504
rect 4594 5499 4595 5503
rect 4599 5499 4600 5503
rect 4594 5498 4600 5499
rect 4794 5503 4800 5504
rect 4794 5499 4795 5503
rect 4799 5499 4800 5503
rect 4794 5498 4800 5499
rect 4994 5503 5000 5504
rect 4994 5499 4995 5503
rect 4999 5499 5000 5503
rect 4994 5498 5000 5499
rect 5194 5503 5200 5504
rect 5194 5499 5195 5503
rect 5199 5499 5200 5503
rect 5662 5500 5663 5504
rect 5667 5500 5668 5504
rect 5662 5499 5668 5500
rect 5194 5498 5200 5499
rect 646 5496 652 5497
rect 110 5495 116 5496
rect 110 5491 111 5495
rect 115 5491 116 5495
rect 646 5492 647 5496
rect 651 5492 652 5496
rect 646 5491 652 5492
rect 782 5496 788 5497
rect 782 5492 783 5496
rect 787 5492 788 5496
rect 782 5491 788 5492
rect 926 5496 932 5497
rect 926 5492 927 5496
rect 931 5492 932 5496
rect 926 5491 932 5492
rect 1078 5496 1084 5497
rect 1078 5492 1079 5496
rect 1083 5492 1084 5496
rect 1078 5491 1084 5492
rect 1230 5496 1236 5497
rect 1230 5492 1231 5496
rect 1235 5492 1236 5496
rect 1230 5491 1236 5492
rect 1382 5496 1388 5497
rect 1382 5492 1383 5496
rect 1387 5492 1388 5496
rect 1382 5491 1388 5492
rect 1534 5496 1540 5497
rect 1534 5492 1535 5496
rect 1539 5492 1540 5496
rect 1534 5491 1540 5492
rect 1678 5496 1684 5497
rect 1678 5492 1679 5496
rect 1683 5492 1684 5496
rect 1678 5491 1684 5492
rect 1814 5496 1820 5497
rect 1814 5492 1815 5496
rect 1819 5492 1820 5496
rect 1814 5491 1820 5492
rect 1934 5495 1940 5496
rect 1934 5491 1935 5495
rect 1939 5491 1940 5495
rect 110 5490 116 5491
rect 112 5459 114 5490
rect 648 5459 650 5491
rect 784 5459 786 5491
rect 928 5459 930 5491
rect 1080 5459 1082 5491
rect 1232 5459 1234 5491
rect 1384 5459 1386 5491
rect 1536 5459 1538 5491
rect 1680 5459 1682 5491
rect 1816 5459 1818 5491
rect 1934 5490 1940 5491
rect 1936 5459 1938 5490
rect 2922 5489 2928 5490
rect 1974 5488 1980 5489
rect 1974 5484 1975 5488
rect 1979 5484 1980 5488
rect 2922 5485 2923 5489
rect 2927 5485 2928 5489
rect 2922 5484 2928 5485
rect 3074 5489 3080 5490
rect 3074 5485 3075 5489
rect 3079 5485 3080 5489
rect 3074 5484 3080 5485
rect 3226 5489 3232 5490
rect 3226 5485 3227 5489
rect 3231 5485 3232 5489
rect 3226 5484 3232 5485
rect 3386 5489 3392 5490
rect 3386 5485 3387 5489
rect 3391 5485 3392 5489
rect 3386 5484 3392 5485
rect 3798 5488 3804 5489
rect 4238 5488 4244 5489
rect 3798 5484 3799 5488
rect 3803 5484 3804 5488
rect 1974 5483 1980 5484
rect 111 5458 115 5459
rect 111 5453 115 5454
rect 591 5458 595 5459
rect 591 5453 595 5454
rect 647 5458 651 5459
rect 647 5453 651 5454
rect 727 5458 731 5459
rect 727 5453 731 5454
rect 783 5458 787 5459
rect 783 5453 787 5454
rect 863 5458 867 5459
rect 863 5453 867 5454
rect 927 5458 931 5459
rect 927 5453 931 5454
rect 999 5458 1003 5459
rect 999 5453 1003 5454
rect 1079 5458 1083 5459
rect 1079 5453 1083 5454
rect 1135 5458 1139 5459
rect 1135 5453 1139 5454
rect 1231 5458 1235 5459
rect 1231 5453 1235 5454
rect 1271 5458 1275 5459
rect 1271 5453 1275 5454
rect 1383 5458 1387 5459
rect 1383 5453 1387 5454
rect 1407 5458 1411 5459
rect 1407 5453 1411 5454
rect 1535 5458 1539 5459
rect 1535 5453 1539 5454
rect 1543 5458 1547 5459
rect 1543 5453 1547 5454
rect 1679 5458 1683 5459
rect 1679 5453 1683 5454
rect 1815 5458 1819 5459
rect 1815 5453 1819 5454
rect 1935 5458 1939 5459
rect 1935 5453 1939 5454
rect 112 5430 114 5453
rect 110 5429 116 5430
rect 592 5429 594 5453
rect 728 5429 730 5453
rect 864 5429 866 5453
rect 1000 5429 1002 5453
rect 1136 5429 1138 5453
rect 1272 5429 1274 5453
rect 1408 5429 1410 5453
rect 1544 5429 1546 5453
rect 1680 5429 1682 5453
rect 1816 5429 1818 5453
rect 1936 5430 1938 5453
rect 1934 5429 1940 5430
rect 110 5425 111 5429
rect 115 5425 116 5429
rect 110 5424 116 5425
rect 590 5428 596 5429
rect 590 5424 591 5428
rect 595 5424 596 5428
rect 590 5423 596 5424
rect 726 5428 732 5429
rect 726 5424 727 5428
rect 731 5424 732 5428
rect 726 5423 732 5424
rect 862 5428 868 5429
rect 862 5424 863 5428
rect 867 5424 868 5428
rect 862 5423 868 5424
rect 998 5428 1004 5429
rect 998 5424 999 5428
rect 1003 5424 1004 5428
rect 998 5423 1004 5424
rect 1134 5428 1140 5429
rect 1134 5424 1135 5428
rect 1139 5424 1140 5428
rect 1134 5423 1140 5424
rect 1270 5428 1276 5429
rect 1270 5424 1271 5428
rect 1275 5424 1276 5428
rect 1270 5423 1276 5424
rect 1406 5428 1412 5429
rect 1406 5424 1407 5428
rect 1411 5424 1412 5428
rect 1406 5423 1412 5424
rect 1542 5428 1548 5429
rect 1542 5424 1543 5428
rect 1547 5424 1548 5428
rect 1542 5423 1548 5424
rect 1678 5428 1684 5429
rect 1678 5424 1679 5428
rect 1683 5424 1684 5428
rect 1678 5423 1684 5424
rect 1814 5428 1820 5429
rect 1814 5424 1815 5428
rect 1819 5424 1820 5428
rect 1934 5425 1935 5429
rect 1939 5425 1940 5429
rect 1934 5424 1940 5425
rect 1814 5423 1820 5424
rect 562 5413 568 5414
rect 110 5412 116 5413
rect 110 5408 111 5412
rect 115 5408 116 5412
rect 562 5409 563 5413
rect 567 5409 568 5413
rect 562 5408 568 5409
rect 698 5413 704 5414
rect 698 5409 699 5413
rect 703 5409 704 5413
rect 698 5408 704 5409
rect 834 5413 840 5414
rect 834 5409 835 5413
rect 839 5409 840 5413
rect 834 5408 840 5409
rect 970 5413 976 5414
rect 970 5409 971 5413
rect 975 5409 976 5413
rect 970 5408 976 5409
rect 1106 5413 1112 5414
rect 1106 5409 1107 5413
rect 1111 5409 1112 5413
rect 1106 5408 1112 5409
rect 1242 5413 1248 5414
rect 1242 5409 1243 5413
rect 1247 5409 1248 5413
rect 1242 5408 1248 5409
rect 1378 5413 1384 5414
rect 1378 5409 1379 5413
rect 1383 5409 1384 5413
rect 1378 5408 1384 5409
rect 1514 5413 1520 5414
rect 1514 5409 1515 5413
rect 1519 5409 1520 5413
rect 1514 5408 1520 5409
rect 1650 5413 1656 5414
rect 1650 5409 1651 5413
rect 1655 5409 1656 5413
rect 1650 5408 1656 5409
rect 1786 5413 1792 5414
rect 1786 5409 1787 5413
rect 1791 5409 1792 5413
rect 1786 5408 1792 5409
rect 1934 5412 1940 5413
rect 1934 5408 1935 5412
rect 1939 5408 1940 5412
rect 110 5407 116 5408
rect 112 5323 114 5407
rect 564 5323 566 5408
rect 700 5323 702 5408
rect 836 5323 838 5408
rect 972 5323 974 5408
rect 1108 5323 1110 5408
rect 1244 5323 1246 5408
rect 1380 5323 1382 5408
rect 1516 5323 1518 5408
rect 1652 5323 1654 5408
rect 1788 5323 1790 5408
rect 1934 5407 1940 5408
rect 1936 5323 1938 5407
rect 1976 5375 1978 5483
rect 2924 5375 2926 5484
rect 3076 5375 3078 5484
rect 3228 5375 3230 5484
rect 3388 5375 3390 5484
rect 3798 5483 3804 5484
rect 3838 5487 3844 5488
rect 3838 5483 3839 5487
rect 3843 5483 3844 5487
rect 4238 5484 4239 5488
rect 4243 5484 4244 5488
rect 4238 5483 4244 5484
rect 4430 5488 4436 5489
rect 4430 5484 4431 5488
rect 4435 5484 4436 5488
rect 4430 5483 4436 5484
rect 4622 5488 4628 5489
rect 4622 5484 4623 5488
rect 4627 5484 4628 5488
rect 4622 5483 4628 5484
rect 4822 5488 4828 5489
rect 4822 5484 4823 5488
rect 4827 5484 4828 5488
rect 4822 5483 4828 5484
rect 5022 5488 5028 5489
rect 5022 5484 5023 5488
rect 5027 5484 5028 5488
rect 5022 5483 5028 5484
rect 5222 5488 5228 5489
rect 5222 5484 5223 5488
rect 5227 5484 5228 5488
rect 5222 5483 5228 5484
rect 5662 5487 5668 5488
rect 5662 5483 5663 5487
rect 5667 5483 5668 5487
rect 3800 5375 3802 5483
rect 3838 5482 3844 5483
rect 3840 5423 3842 5482
rect 4240 5423 4242 5483
rect 4432 5423 4434 5483
rect 4624 5423 4626 5483
rect 4824 5423 4826 5483
rect 5024 5423 5026 5483
rect 5224 5423 5226 5483
rect 5662 5482 5668 5483
rect 5664 5423 5666 5482
rect 3839 5422 3843 5423
rect 3839 5417 3843 5418
rect 4239 5422 4243 5423
rect 4239 5417 4243 5418
rect 4303 5422 4307 5423
rect 4303 5417 4307 5418
rect 4431 5422 4435 5423
rect 4431 5417 4435 5418
rect 4519 5422 4523 5423
rect 4519 5417 4523 5418
rect 4623 5422 4627 5423
rect 4623 5417 4627 5418
rect 4735 5422 4739 5423
rect 4735 5417 4739 5418
rect 4823 5422 4827 5423
rect 4823 5417 4827 5418
rect 4951 5422 4955 5423
rect 4951 5417 4955 5418
rect 5023 5422 5027 5423
rect 5023 5417 5027 5418
rect 5175 5422 5179 5423
rect 5175 5417 5179 5418
rect 5223 5422 5227 5423
rect 5223 5417 5227 5418
rect 5399 5422 5403 5423
rect 5399 5417 5403 5418
rect 5663 5422 5667 5423
rect 5663 5417 5667 5418
rect 3840 5394 3842 5417
rect 3838 5393 3844 5394
rect 4304 5393 4306 5417
rect 4520 5393 4522 5417
rect 4736 5393 4738 5417
rect 4952 5393 4954 5417
rect 5176 5393 5178 5417
rect 5400 5393 5402 5417
rect 5664 5394 5666 5417
rect 5662 5393 5668 5394
rect 3838 5389 3839 5393
rect 3843 5389 3844 5393
rect 3838 5388 3844 5389
rect 4302 5392 4308 5393
rect 4302 5388 4303 5392
rect 4307 5388 4308 5392
rect 4302 5387 4308 5388
rect 4518 5392 4524 5393
rect 4518 5388 4519 5392
rect 4523 5388 4524 5392
rect 4518 5387 4524 5388
rect 4734 5392 4740 5393
rect 4734 5388 4735 5392
rect 4739 5388 4740 5392
rect 4734 5387 4740 5388
rect 4950 5392 4956 5393
rect 4950 5388 4951 5392
rect 4955 5388 4956 5392
rect 4950 5387 4956 5388
rect 5174 5392 5180 5393
rect 5174 5388 5175 5392
rect 5179 5388 5180 5392
rect 5174 5387 5180 5388
rect 5398 5392 5404 5393
rect 5398 5388 5399 5392
rect 5403 5388 5404 5392
rect 5662 5389 5663 5393
rect 5667 5389 5668 5393
rect 5662 5388 5668 5389
rect 5398 5387 5404 5388
rect 4274 5377 4280 5378
rect 3838 5376 3844 5377
rect 1975 5374 1979 5375
rect 1975 5369 1979 5370
rect 2643 5374 2647 5375
rect 2643 5369 2647 5370
rect 2811 5374 2815 5375
rect 2811 5369 2815 5370
rect 2923 5374 2927 5375
rect 2923 5369 2927 5370
rect 2979 5374 2983 5375
rect 2979 5369 2983 5370
rect 3075 5374 3079 5375
rect 3075 5369 3079 5370
rect 3139 5374 3143 5375
rect 3139 5369 3143 5370
rect 3227 5374 3231 5375
rect 3227 5369 3231 5370
rect 3307 5374 3311 5375
rect 3307 5369 3311 5370
rect 3387 5374 3391 5375
rect 3387 5369 3391 5370
rect 3475 5374 3479 5375
rect 3475 5369 3479 5370
rect 3643 5374 3647 5375
rect 3643 5369 3647 5370
rect 3799 5374 3803 5375
rect 3838 5372 3839 5376
rect 3843 5372 3844 5376
rect 4274 5373 4275 5377
rect 4279 5373 4280 5377
rect 4274 5372 4280 5373
rect 4490 5377 4496 5378
rect 4490 5373 4491 5377
rect 4495 5373 4496 5377
rect 4490 5372 4496 5373
rect 4706 5377 4712 5378
rect 4706 5373 4707 5377
rect 4711 5373 4712 5377
rect 4706 5372 4712 5373
rect 4922 5377 4928 5378
rect 4922 5373 4923 5377
rect 4927 5373 4928 5377
rect 4922 5372 4928 5373
rect 5146 5377 5152 5378
rect 5146 5373 5147 5377
rect 5151 5373 5152 5377
rect 5146 5372 5152 5373
rect 5370 5377 5376 5378
rect 5370 5373 5371 5377
rect 5375 5373 5376 5377
rect 5370 5372 5376 5373
rect 5662 5376 5668 5377
rect 5662 5372 5663 5376
rect 5667 5372 5668 5376
rect 3838 5371 3844 5372
rect 3799 5369 3803 5370
rect 111 5322 115 5323
rect 111 5317 115 5318
rect 411 5322 415 5323
rect 411 5317 415 5318
rect 563 5322 567 5323
rect 563 5317 567 5318
rect 587 5322 591 5323
rect 587 5317 591 5318
rect 699 5322 703 5323
rect 699 5317 703 5318
rect 763 5322 767 5323
rect 763 5317 767 5318
rect 835 5322 839 5323
rect 835 5317 839 5318
rect 939 5322 943 5323
rect 939 5317 943 5318
rect 971 5322 975 5323
rect 971 5317 975 5318
rect 1107 5322 1111 5323
rect 1107 5317 1111 5318
rect 1243 5322 1247 5323
rect 1243 5317 1247 5318
rect 1275 5322 1279 5323
rect 1275 5317 1279 5318
rect 1379 5322 1383 5323
rect 1379 5317 1383 5318
rect 1443 5322 1447 5323
rect 1443 5317 1447 5318
rect 1515 5322 1519 5323
rect 1515 5317 1519 5318
rect 1611 5322 1615 5323
rect 1611 5317 1615 5318
rect 1651 5322 1655 5323
rect 1651 5317 1655 5318
rect 1787 5322 1791 5323
rect 1787 5317 1791 5318
rect 1935 5322 1939 5323
rect 1935 5317 1939 5318
rect 112 5257 114 5317
rect 110 5256 116 5257
rect 412 5256 414 5317
rect 588 5256 590 5317
rect 764 5256 766 5317
rect 940 5256 942 5317
rect 1108 5256 1110 5317
rect 1276 5256 1278 5317
rect 1444 5256 1446 5317
rect 1612 5256 1614 5317
rect 1788 5256 1790 5317
rect 1936 5257 1938 5317
rect 1976 5309 1978 5369
rect 1974 5308 1980 5309
rect 2644 5308 2646 5369
rect 2812 5308 2814 5369
rect 2980 5308 2982 5369
rect 3140 5308 3142 5369
rect 3308 5308 3310 5369
rect 3476 5308 3478 5369
rect 3644 5308 3646 5369
rect 3800 5309 3802 5369
rect 3798 5308 3804 5309
rect 1974 5304 1975 5308
rect 1979 5304 1980 5308
rect 1974 5303 1980 5304
rect 2642 5307 2648 5308
rect 2642 5303 2643 5307
rect 2647 5303 2648 5307
rect 2642 5302 2648 5303
rect 2810 5307 2816 5308
rect 2810 5303 2811 5307
rect 2815 5303 2816 5307
rect 2810 5302 2816 5303
rect 2978 5307 2984 5308
rect 2978 5303 2979 5307
rect 2983 5303 2984 5307
rect 2978 5302 2984 5303
rect 3138 5307 3144 5308
rect 3138 5303 3139 5307
rect 3143 5303 3144 5307
rect 3138 5302 3144 5303
rect 3306 5307 3312 5308
rect 3306 5303 3307 5307
rect 3311 5303 3312 5307
rect 3306 5302 3312 5303
rect 3474 5307 3480 5308
rect 3474 5303 3475 5307
rect 3479 5303 3480 5307
rect 3474 5302 3480 5303
rect 3642 5307 3648 5308
rect 3642 5303 3643 5307
rect 3647 5303 3648 5307
rect 3798 5304 3799 5308
rect 3803 5304 3804 5308
rect 3798 5303 3804 5304
rect 3642 5302 3648 5303
rect 2670 5292 2676 5293
rect 1974 5291 1980 5292
rect 1974 5287 1975 5291
rect 1979 5287 1980 5291
rect 2670 5288 2671 5292
rect 2675 5288 2676 5292
rect 2670 5287 2676 5288
rect 2838 5292 2844 5293
rect 2838 5288 2839 5292
rect 2843 5288 2844 5292
rect 2838 5287 2844 5288
rect 3006 5292 3012 5293
rect 3006 5288 3007 5292
rect 3011 5288 3012 5292
rect 3006 5287 3012 5288
rect 3166 5292 3172 5293
rect 3166 5288 3167 5292
rect 3171 5288 3172 5292
rect 3166 5287 3172 5288
rect 3334 5292 3340 5293
rect 3334 5288 3335 5292
rect 3339 5288 3340 5292
rect 3334 5287 3340 5288
rect 3502 5292 3508 5293
rect 3502 5288 3503 5292
rect 3507 5288 3508 5292
rect 3502 5287 3508 5288
rect 3670 5292 3676 5293
rect 3670 5288 3671 5292
rect 3675 5288 3676 5292
rect 3670 5287 3676 5288
rect 3798 5291 3804 5292
rect 3798 5287 3799 5291
rect 3803 5287 3804 5291
rect 1974 5286 1980 5287
rect 1976 5263 1978 5286
rect 2672 5263 2674 5287
rect 2840 5263 2842 5287
rect 3008 5263 3010 5287
rect 3168 5263 3170 5287
rect 3336 5263 3338 5287
rect 3504 5263 3506 5287
rect 3672 5263 3674 5287
rect 3798 5286 3804 5287
rect 3800 5263 3802 5286
rect 3840 5279 3842 5371
rect 4276 5279 4278 5372
rect 4492 5279 4494 5372
rect 4708 5279 4710 5372
rect 4924 5279 4926 5372
rect 5148 5279 5150 5372
rect 5372 5279 5374 5372
rect 5662 5371 5668 5372
rect 5664 5279 5666 5371
rect 3839 5278 3843 5279
rect 3839 5273 3843 5274
rect 4275 5278 4279 5279
rect 4275 5273 4279 5274
rect 4371 5278 4375 5279
rect 4371 5273 4375 5274
rect 4491 5278 4495 5279
rect 4491 5273 4495 5274
rect 4563 5278 4567 5279
rect 4563 5273 4567 5274
rect 4707 5278 4711 5279
rect 4707 5273 4711 5274
rect 4771 5278 4775 5279
rect 4771 5273 4775 5274
rect 4923 5278 4927 5279
rect 4923 5273 4927 5274
rect 4979 5278 4983 5279
rect 4979 5273 4983 5274
rect 5147 5278 5151 5279
rect 5147 5273 5151 5274
rect 5195 5278 5199 5279
rect 5195 5273 5199 5274
rect 5371 5278 5375 5279
rect 5371 5273 5375 5274
rect 5419 5278 5423 5279
rect 5419 5273 5423 5274
rect 5663 5278 5667 5279
rect 5663 5273 5667 5274
rect 1975 5262 1979 5263
rect 1975 5257 1979 5258
rect 2511 5262 2515 5263
rect 2511 5257 2515 5258
rect 2671 5262 2675 5263
rect 2671 5257 2675 5258
rect 2687 5262 2691 5263
rect 2687 5257 2691 5258
rect 2839 5262 2843 5263
rect 2839 5257 2843 5258
rect 2863 5262 2867 5263
rect 2863 5257 2867 5258
rect 3007 5262 3011 5263
rect 3007 5257 3011 5258
rect 3039 5262 3043 5263
rect 3039 5257 3043 5258
rect 3167 5262 3171 5263
rect 3167 5257 3171 5258
rect 3207 5262 3211 5263
rect 3207 5257 3211 5258
rect 3335 5262 3339 5263
rect 3335 5257 3339 5258
rect 3367 5262 3371 5263
rect 3367 5257 3371 5258
rect 3503 5262 3507 5263
rect 3503 5257 3507 5258
rect 3535 5262 3539 5263
rect 3535 5257 3539 5258
rect 3671 5262 3675 5263
rect 3671 5257 3675 5258
rect 3679 5262 3683 5263
rect 3679 5257 3683 5258
rect 3799 5262 3803 5263
rect 3799 5257 3803 5258
rect 1934 5256 1940 5257
rect 110 5252 111 5256
rect 115 5252 116 5256
rect 110 5251 116 5252
rect 410 5255 416 5256
rect 410 5251 411 5255
rect 415 5251 416 5255
rect 410 5250 416 5251
rect 586 5255 592 5256
rect 586 5251 587 5255
rect 591 5251 592 5255
rect 586 5250 592 5251
rect 762 5255 768 5256
rect 762 5251 763 5255
rect 767 5251 768 5255
rect 762 5250 768 5251
rect 938 5255 944 5256
rect 938 5251 939 5255
rect 943 5251 944 5255
rect 938 5250 944 5251
rect 1106 5255 1112 5256
rect 1106 5251 1107 5255
rect 1111 5251 1112 5255
rect 1106 5250 1112 5251
rect 1274 5255 1280 5256
rect 1274 5251 1275 5255
rect 1279 5251 1280 5255
rect 1274 5250 1280 5251
rect 1442 5255 1448 5256
rect 1442 5251 1443 5255
rect 1447 5251 1448 5255
rect 1442 5250 1448 5251
rect 1610 5255 1616 5256
rect 1610 5251 1611 5255
rect 1615 5251 1616 5255
rect 1610 5250 1616 5251
rect 1786 5255 1792 5256
rect 1786 5251 1787 5255
rect 1791 5251 1792 5255
rect 1934 5252 1935 5256
rect 1939 5252 1940 5256
rect 1934 5251 1940 5252
rect 1786 5250 1792 5251
rect 438 5240 444 5241
rect 110 5239 116 5240
rect 110 5235 111 5239
rect 115 5235 116 5239
rect 438 5236 439 5240
rect 443 5236 444 5240
rect 438 5235 444 5236
rect 614 5240 620 5241
rect 614 5236 615 5240
rect 619 5236 620 5240
rect 614 5235 620 5236
rect 790 5240 796 5241
rect 790 5236 791 5240
rect 795 5236 796 5240
rect 790 5235 796 5236
rect 966 5240 972 5241
rect 966 5236 967 5240
rect 971 5236 972 5240
rect 966 5235 972 5236
rect 1134 5240 1140 5241
rect 1134 5236 1135 5240
rect 1139 5236 1140 5240
rect 1134 5235 1140 5236
rect 1302 5240 1308 5241
rect 1302 5236 1303 5240
rect 1307 5236 1308 5240
rect 1302 5235 1308 5236
rect 1470 5240 1476 5241
rect 1470 5236 1471 5240
rect 1475 5236 1476 5240
rect 1470 5235 1476 5236
rect 1638 5240 1644 5241
rect 1638 5236 1639 5240
rect 1643 5236 1644 5240
rect 1638 5235 1644 5236
rect 1814 5240 1820 5241
rect 1814 5236 1815 5240
rect 1819 5236 1820 5240
rect 1814 5235 1820 5236
rect 1934 5239 1940 5240
rect 1934 5235 1935 5239
rect 1939 5235 1940 5239
rect 110 5234 116 5235
rect 112 5203 114 5234
rect 440 5203 442 5235
rect 616 5203 618 5235
rect 792 5203 794 5235
rect 968 5203 970 5235
rect 1136 5203 1138 5235
rect 1304 5203 1306 5235
rect 1472 5203 1474 5235
rect 1640 5203 1642 5235
rect 1816 5203 1818 5235
rect 1934 5234 1940 5235
rect 1976 5234 1978 5257
rect 1936 5203 1938 5234
rect 1974 5233 1980 5234
rect 2512 5233 2514 5257
rect 2688 5233 2690 5257
rect 2864 5233 2866 5257
rect 3040 5233 3042 5257
rect 3208 5233 3210 5257
rect 3368 5233 3370 5257
rect 3536 5233 3538 5257
rect 3680 5233 3682 5257
rect 3800 5234 3802 5257
rect 3798 5233 3804 5234
rect 1974 5229 1975 5233
rect 1979 5229 1980 5233
rect 1974 5228 1980 5229
rect 2510 5232 2516 5233
rect 2510 5228 2511 5232
rect 2515 5228 2516 5232
rect 2510 5227 2516 5228
rect 2686 5232 2692 5233
rect 2686 5228 2687 5232
rect 2691 5228 2692 5232
rect 2686 5227 2692 5228
rect 2862 5232 2868 5233
rect 2862 5228 2863 5232
rect 2867 5228 2868 5232
rect 2862 5227 2868 5228
rect 3038 5232 3044 5233
rect 3038 5228 3039 5232
rect 3043 5228 3044 5232
rect 3038 5227 3044 5228
rect 3206 5232 3212 5233
rect 3206 5228 3207 5232
rect 3211 5228 3212 5232
rect 3206 5227 3212 5228
rect 3366 5232 3372 5233
rect 3366 5228 3367 5232
rect 3371 5228 3372 5232
rect 3366 5227 3372 5228
rect 3534 5232 3540 5233
rect 3534 5228 3535 5232
rect 3539 5228 3540 5232
rect 3534 5227 3540 5228
rect 3678 5232 3684 5233
rect 3678 5228 3679 5232
rect 3683 5228 3684 5232
rect 3798 5229 3799 5233
rect 3803 5229 3804 5233
rect 3798 5228 3804 5229
rect 3678 5227 3684 5228
rect 2482 5217 2488 5218
rect 1974 5216 1980 5217
rect 1974 5212 1975 5216
rect 1979 5212 1980 5216
rect 2482 5213 2483 5217
rect 2487 5213 2488 5217
rect 2482 5212 2488 5213
rect 2658 5217 2664 5218
rect 2658 5213 2659 5217
rect 2663 5213 2664 5217
rect 2658 5212 2664 5213
rect 2834 5217 2840 5218
rect 2834 5213 2835 5217
rect 2839 5213 2840 5217
rect 2834 5212 2840 5213
rect 3010 5217 3016 5218
rect 3010 5213 3011 5217
rect 3015 5213 3016 5217
rect 3010 5212 3016 5213
rect 3178 5217 3184 5218
rect 3178 5213 3179 5217
rect 3183 5213 3184 5217
rect 3178 5212 3184 5213
rect 3338 5217 3344 5218
rect 3338 5213 3339 5217
rect 3343 5213 3344 5217
rect 3338 5212 3344 5213
rect 3506 5217 3512 5218
rect 3506 5213 3507 5217
rect 3511 5213 3512 5217
rect 3506 5212 3512 5213
rect 3650 5217 3656 5218
rect 3650 5213 3651 5217
rect 3655 5213 3656 5217
rect 3650 5212 3656 5213
rect 3798 5216 3804 5217
rect 3798 5212 3799 5216
rect 3803 5212 3804 5216
rect 3840 5213 3842 5273
rect 1974 5211 1980 5212
rect 111 5202 115 5203
rect 111 5197 115 5198
rect 207 5202 211 5203
rect 207 5197 211 5198
rect 343 5202 347 5203
rect 343 5197 347 5198
rect 439 5202 443 5203
rect 439 5197 443 5198
rect 479 5202 483 5203
rect 479 5197 483 5198
rect 615 5202 619 5203
rect 615 5197 619 5198
rect 751 5202 755 5203
rect 751 5197 755 5198
rect 791 5202 795 5203
rect 791 5197 795 5198
rect 887 5202 891 5203
rect 887 5197 891 5198
rect 967 5202 971 5203
rect 967 5197 971 5198
rect 1023 5202 1027 5203
rect 1023 5197 1027 5198
rect 1135 5202 1139 5203
rect 1135 5197 1139 5198
rect 1303 5202 1307 5203
rect 1303 5197 1307 5198
rect 1471 5202 1475 5203
rect 1471 5197 1475 5198
rect 1639 5202 1643 5203
rect 1639 5197 1643 5198
rect 1815 5202 1819 5203
rect 1815 5197 1819 5198
rect 1935 5202 1939 5203
rect 1935 5197 1939 5198
rect 112 5174 114 5197
rect 110 5173 116 5174
rect 208 5173 210 5197
rect 344 5173 346 5197
rect 480 5173 482 5197
rect 616 5173 618 5197
rect 752 5173 754 5197
rect 888 5173 890 5197
rect 1024 5173 1026 5197
rect 1936 5174 1938 5197
rect 1934 5173 1940 5174
rect 110 5169 111 5173
rect 115 5169 116 5173
rect 110 5168 116 5169
rect 206 5172 212 5173
rect 206 5168 207 5172
rect 211 5168 212 5172
rect 206 5167 212 5168
rect 342 5172 348 5173
rect 342 5168 343 5172
rect 347 5168 348 5172
rect 342 5167 348 5168
rect 478 5172 484 5173
rect 478 5168 479 5172
rect 483 5168 484 5172
rect 478 5167 484 5168
rect 614 5172 620 5173
rect 614 5168 615 5172
rect 619 5168 620 5172
rect 614 5167 620 5168
rect 750 5172 756 5173
rect 750 5168 751 5172
rect 755 5168 756 5172
rect 750 5167 756 5168
rect 886 5172 892 5173
rect 886 5168 887 5172
rect 891 5168 892 5172
rect 886 5167 892 5168
rect 1022 5172 1028 5173
rect 1022 5168 1023 5172
rect 1027 5168 1028 5172
rect 1934 5169 1935 5173
rect 1939 5169 1940 5173
rect 1934 5168 1940 5169
rect 1022 5167 1028 5168
rect 178 5157 184 5158
rect 110 5156 116 5157
rect 110 5152 111 5156
rect 115 5152 116 5156
rect 178 5153 179 5157
rect 183 5153 184 5157
rect 178 5152 184 5153
rect 314 5157 320 5158
rect 314 5153 315 5157
rect 319 5153 320 5157
rect 314 5152 320 5153
rect 450 5157 456 5158
rect 450 5153 451 5157
rect 455 5153 456 5157
rect 450 5152 456 5153
rect 586 5157 592 5158
rect 586 5153 587 5157
rect 591 5153 592 5157
rect 586 5152 592 5153
rect 722 5157 728 5158
rect 722 5153 723 5157
rect 727 5153 728 5157
rect 722 5152 728 5153
rect 858 5157 864 5158
rect 858 5153 859 5157
rect 863 5153 864 5157
rect 858 5152 864 5153
rect 994 5157 1000 5158
rect 994 5153 995 5157
rect 999 5153 1000 5157
rect 994 5152 1000 5153
rect 1934 5156 1940 5157
rect 1934 5152 1935 5156
rect 1939 5152 1940 5156
rect 110 5151 116 5152
rect 112 5071 114 5151
rect 180 5071 182 5152
rect 316 5071 318 5152
rect 452 5071 454 5152
rect 588 5071 590 5152
rect 724 5071 726 5152
rect 860 5071 862 5152
rect 996 5071 998 5152
rect 1934 5151 1940 5152
rect 1936 5071 1938 5151
rect 1976 5143 1978 5211
rect 2484 5143 2486 5212
rect 2660 5143 2662 5212
rect 2836 5143 2838 5212
rect 3012 5143 3014 5212
rect 3180 5143 3182 5212
rect 3340 5143 3342 5212
rect 3508 5143 3510 5212
rect 3652 5143 3654 5212
rect 3798 5211 3804 5212
rect 3838 5212 3844 5213
rect 4372 5212 4374 5273
rect 4564 5212 4566 5273
rect 4772 5212 4774 5273
rect 4980 5212 4982 5273
rect 5196 5212 5198 5273
rect 5420 5212 5422 5273
rect 5664 5213 5666 5273
rect 5662 5212 5668 5213
rect 3800 5143 3802 5211
rect 3838 5208 3839 5212
rect 3843 5208 3844 5212
rect 3838 5207 3844 5208
rect 4370 5211 4376 5212
rect 4370 5207 4371 5211
rect 4375 5207 4376 5211
rect 4370 5206 4376 5207
rect 4562 5211 4568 5212
rect 4562 5207 4563 5211
rect 4567 5207 4568 5211
rect 4562 5206 4568 5207
rect 4770 5211 4776 5212
rect 4770 5207 4771 5211
rect 4775 5207 4776 5211
rect 4770 5206 4776 5207
rect 4978 5211 4984 5212
rect 4978 5207 4979 5211
rect 4983 5207 4984 5211
rect 4978 5206 4984 5207
rect 5194 5211 5200 5212
rect 5194 5207 5195 5211
rect 5199 5207 5200 5211
rect 5194 5206 5200 5207
rect 5418 5211 5424 5212
rect 5418 5207 5419 5211
rect 5423 5207 5424 5211
rect 5662 5208 5663 5212
rect 5667 5208 5668 5212
rect 5662 5207 5668 5208
rect 5418 5206 5424 5207
rect 4398 5196 4404 5197
rect 3838 5195 3844 5196
rect 3838 5191 3839 5195
rect 3843 5191 3844 5195
rect 4398 5192 4399 5196
rect 4403 5192 4404 5196
rect 4398 5191 4404 5192
rect 4590 5196 4596 5197
rect 4590 5192 4591 5196
rect 4595 5192 4596 5196
rect 4590 5191 4596 5192
rect 4798 5196 4804 5197
rect 4798 5192 4799 5196
rect 4803 5192 4804 5196
rect 4798 5191 4804 5192
rect 5006 5196 5012 5197
rect 5006 5192 5007 5196
rect 5011 5192 5012 5196
rect 5006 5191 5012 5192
rect 5222 5196 5228 5197
rect 5222 5192 5223 5196
rect 5227 5192 5228 5196
rect 5222 5191 5228 5192
rect 5446 5196 5452 5197
rect 5446 5192 5447 5196
rect 5451 5192 5452 5196
rect 5446 5191 5452 5192
rect 5662 5195 5668 5196
rect 5662 5191 5663 5195
rect 5667 5191 5668 5195
rect 3838 5190 3844 5191
rect 3840 5143 3842 5190
rect 4400 5143 4402 5191
rect 4592 5143 4594 5191
rect 4800 5143 4802 5191
rect 5008 5143 5010 5191
rect 5224 5143 5226 5191
rect 5448 5143 5450 5191
rect 5662 5190 5668 5191
rect 5664 5143 5666 5190
rect 1975 5142 1979 5143
rect 1975 5137 1979 5138
rect 2139 5142 2143 5143
rect 2139 5137 2143 5138
rect 2307 5142 2311 5143
rect 2307 5137 2311 5138
rect 2483 5142 2487 5143
rect 2483 5137 2487 5138
rect 2491 5142 2495 5143
rect 2491 5137 2495 5138
rect 2659 5142 2663 5143
rect 2659 5137 2663 5138
rect 2691 5142 2695 5143
rect 2691 5137 2695 5138
rect 2835 5142 2839 5143
rect 2835 5137 2839 5138
rect 2915 5142 2919 5143
rect 2915 5137 2919 5138
rect 3011 5142 3015 5143
rect 3011 5137 3015 5138
rect 3163 5142 3167 5143
rect 3163 5137 3167 5138
rect 3179 5142 3183 5143
rect 3179 5137 3183 5138
rect 3339 5142 3343 5143
rect 3339 5137 3343 5138
rect 3419 5142 3423 5143
rect 3419 5137 3423 5138
rect 3507 5142 3511 5143
rect 3507 5137 3511 5138
rect 3651 5142 3655 5143
rect 3651 5137 3655 5138
rect 3799 5142 3803 5143
rect 3799 5137 3803 5138
rect 3839 5142 3843 5143
rect 3839 5137 3843 5138
rect 3887 5142 3891 5143
rect 3887 5137 3891 5138
rect 4087 5142 4091 5143
rect 4087 5137 4091 5138
rect 4311 5142 4315 5143
rect 4311 5137 4315 5138
rect 4399 5142 4403 5143
rect 4399 5137 4403 5138
rect 4535 5142 4539 5143
rect 4535 5137 4539 5138
rect 4591 5142 4595 5143
rect 4591 5137 4595 5138
rect 4759 5142 4763 5143
rect 4759 5137 4763 5138
rect 4799 5142 4803 5143
rect 4799 5137 4803 5138
rect 4983 5142 4987 5143
rect 4983 5137 4987 5138
rect 5007 5142 5011 5143
rect 5007 5137 5011 5138
rect 5207 5142 5211 5143
rect 5207 5137 5211 5138
rect 5223 5142 5227 5143
rect 5223 5137 5227 5138
rect 5439 5142 5443 5143
rect 5439 5137 5443 5138
rect 5447 5142 5451 5143
rect 5447 5137 5451 5138
rect 5663 5142 5667 5143
rect 5663 5137 5667 5138
rect 1976 5077 1978 5137
rect 1974 5076 1980 5077
rect 2140 5076 2142 5137
rect 2308 5076 2310 5137
rect 2492 5076 2494 5137
rect 2692 5076 2694 5137
rect 2916 5076 2918 5137
rect 3164 5076 3166 5137
rect 3420 5076 3422 5137
rect 3652 5076 3654 5137
rect 3800 5077 3802 5137
rect 3840 5114 3842 5137
rect 3838 5113 3844 5114
rect 3888 5113 3890 5137
rect 4088 5113 4090 5137
rect 4312 5113 4314 5137
rect 4536 5113 4538 5137
rect 4760 5113 4762 5137
rect 4984 5113 4986 5137
rect 5208 5113 5210 5137
rect 5440 5113 5442 5137
rect 5664 5114 5666 5137
rect 5662 5113 5668 5114
rect 3838 5109 3839 5113
rect 3843 5109 3844 5113
rect 3838 5108 3844 5109
rect 3886 5112 3892 5113
rect 3886 5108 3887 5112
rect 3891 5108 3892 5112
rect 3886 5107 3892 5108
rect 4086 5112 4092 5113
rect 4086 5108 4087 5112
rect 4091 5108 4092 5112
rect 4086 5107 4092 5108
rect 4310 5112 4316 5113
rect 4310 5108 4311 5112
rect 4315 5108 4316 5112
rect 4310 5107 4316 5108
rect 4534 5112 4540 5113
rect 4534 5108 4535 5112
rect 4539 5108 4540 5112
rect 4534 5107 4540 5108
rect 4758 5112 4764 5113
rect 4758 5108 4759 5112
rect 4763 5108 4764 5112
rect 4758 5107 4764 5108
rect 4982 5112 4988 5113
rect 4982 5108 4983 5112
rect 4987 5108 4988 5112
rect 4982 5107 4988 5108
rect 5206 5112 5212 5113
rect 5206 5108 5207 5112
rect 5211 5108 5212 5112
rect 5206 5107 5212 5108
rect 5438 5112 5444 5113
rect 5438 5108 5439 5112
rect 5443 5108 5444 5112
rect 5662 5109 5663 5113
rect 5667 5109 5668 5113
rect 5662 5108 5668 5109
rect 5438 5107 5444 5108
rect 3858 5097 3864 5098
rect 3838 5096 3844 5097
rect 3838 5092 3839 5096
rect 3843 5092 3844 5096
rect 3858 5093 3859 5097
rect 3863 5093 3864 5097
rect 3858 5092 3864 5093
rect 4058 5097 4064 5098
rect 4058 5093 4059 5097
rect 4063 5093 4064 5097
rect 4058 5092 4064 5093
rect 4282 5097 4288 5098
rect 4282 5093 4283 5097
rect 4287 5093 4288 5097
rect 4282 5092 4288 5093
rect 4506 5097 4512 5098
rect 4506 5093 4507 5097
rect 4511 5093 4512 5097
rect 4506 5092 4512 5093
rect 4730 5097 4736 5098
rect 4730 5093 4731 5097
rect 4735 5093 4736 5097
rect 4730 5092 4736 5093
rect 4954 5097 4960 5098
rect 4954 5093 4955 5097
rect 4959 5093 4960 5097
rect 4954 5092 4960 5093
rect 5178 5097 5184 5098
rect 5178 5093 5179 5097
rect 5183 5093 5184 5097
rect 5178 5092 5184 5093
rect 5410 5097 5416 5098
rect 5410 5093 5411 5097
rect 5415 5093 5416 5097
rect 5410 5092 5416 5093
rect 5662 5096 5668 5097
rect 5662 5092 5663 5096
rect 5667 5092 5668 5096
rect 3838 5091 3844 5092
rect 3798 5076 3804 5077
rect 1974 5072 1975 5076
rect 1979 5072 1980 5076
rect 1974 5071 1980 5072
rect 2138 5075 2144 5076
rect 2138 5071 2139 5075
rect 2143 5071 2144 5075
rect 111 5070 115 5071
rect 111 5065 115 5066
rect 147 5070 151 5071
rect 147 5065 151 5066
rect 179 5070 183 5071
rect 179 5065 183 5066
rect 315 5070 319 5071
rect 315 5065 319 5066
rect 339 5070 343 5071
rect 339 5065 343 5066
rect 451 5070 455 5071
rect 451 5065 455 5066
rect 531 5070 535 5071
rect 531 5065 535 5066
rect 587 5070 591 5071
rect 587 5065 591 5066
rect 723 5070 727 5071
rect 723 5065 727 5066
rect 731 5070 735 5071
rect 731 5065 735 5066
rect 859 5070 863 5071
rect 859 5065 863 5066
rect 931 5070 935 5071
rect 931 5065 935 5066
rect 995 5070 999 5071
rect 995 5065 999 5066
rect 1131 5070 1135 5071
rect 1131 5065 1135 5066
rect 1935 5070 1939 5071
rect 2138 5070 2144 5071
rect 2306 5075 2312 5076
rect 2306 5071 2307 5075
rect 2311 5071 2312 5075
rect 2306 5070 2312 5071
rect 2490 5075 2496 5076
rect 2490 5071 2491 5075
rect 2495 5071 2496 5075
rect 2490 5070 2496 5071
rect 2690 5075 2696 5076
rect 2690 5071 2691 5075
rect 2695 5071 2696 5075
rect 2690 5070 2696 5071
rect 2914 5075 2920 5076
rect 2914 5071 2915 5075
rect 2919 5071 2920 5075
rect 2914 5070 2920 5071
rect 3162 5075 3168 5076
rect 3162 5071 3163 5075
rect 3167 5071 3168 5075
rect 3162 5070 3168 5071
rect 3418 5075 3424 5076
rect 3418 5071 3419 5075
rect 3423 5071 3424 5075
rect 3418 5070 3424 5071
rect 3650 5075 3656 5076
rect 3650 5071 3651 5075
rect 3655 5071 3656 5075
rect 3798 5072 3799 5076
rect 3803 5072 3804 5076
rect 3798 5071 3804 5072
rect 3650 5070 3656 5071
rect 1935 5065 1939 5066
rect 112 5005 114 5065
rect 110 5004 116 5005
rect 148 5004 150 5065
rect 340 5004 342 5065
rect 532 5004 534 5065
rect 732 5004 734 5065
rect 932 5004 934 5065
rect 1132 5004 1134 5065
rect 1936 5005 1938 5065
rect 2166 5060 2172 5061
rect 1974 5059 1980 5060
rect 1974 5055 1975 5059
rect 1979 5055 1980 5059
rect 2166 5056 2167 5060
rect 2171 5056 2172 5060
rect 2166 5055 2172 5056
rect 2334 5060 2340 5061
rect 2334 5056 2335 5060
rect 2339 5056 2340 5060
rect 2334 5055 2340 5056
rect 2518 5060 2524 5061
rect 2518 5056 2519 5060
rect 2523 5056 2524 5060
rect 2518 5055 2524 5056
rect 2718 5060 2724 5061
rect 2718 5056 2719 5060
rect 2723 5056 2724 5060
rect 2718 5055 2724 5056
rect 2942 5060 2948 5061
rect 2942 5056 2943 5060
rect 2947 5056 2948 5060
rect 2942 5055 2948 5056
rect 3190 5060 3196 5061
rect 3190 5056 3191 5060
rect 3195 5056 3196 5060
rect 3190 5055 3196 5056
rect 3446 5060 3452 5061
rect 3446 5056 3447 5060
rect 3451 5056 3452 5060
rect 3446 5055 3452 5056
rect 3678 5060 3684 5061
rect 3678 5056 3679 5060
rect 3683 5056 3684 5060
rect 3678 5055 3684 5056
rect 3798 5059 3804 5060
rect 3798 5055 3799 5059
rect 3803 5055 3804 5059
rect 1974 5054 1980 5055
rect 1976 5007 1978 5054
rect 2168 5007 2170 5055
rect 2336 5007 2338 5055
rect 2520 5007 2522 5055
rect 2720 5007 2722 5055
rect 2944 5007 2946 5055
rect 3192 5007 3194 5055
rect 3448 5007 3450 5055
rect 3680 5007 3682 5055
rect 3798 5054 3804 5055
rect 3800 5007 3802 5054
rect 3840 5015 3842 5091
rect 3860 5015 3862 5092
rect 4060 5015 4062 5092
rect 4284 5015 4286 5092
rect 4508 5015 4510 5092
rect 4732 5015 4734 5092
rect 4956 5015 4958 5092
rect 5180 5015 5182 5092
rect 5412 5015 5414 5092
rect 5662 5091 5668 5092
rect 5664 5015 5666 5091
rect 3839 5014 3843 5015
rect 3839 5009 3843 5010
rect 3859 5014 3863 5015
rect 3859 5009 3863 5010
rect 3995 5014 3999 5015
rect 3995 5009 3999 5010
rect 4059 5014 4063 5015
rect 4059 5009 4063 5010
rect 4131 5014 4135 5015
rect 4131 5009 4135 5010
rect 4283 5014 4287 5015
rect 4283 5009 4287 5010
rect 4443 5014 4447 5015
rect 4443 5009 4447 5010
rect 4507 5014 4511 5015
rect 4507 5009 4511 5010
rect 4611 5014 4615 5015
rect 4611 5009 4615 5010
rect 4731 5014 4735 5015
rect 4731 5009 4735 5010
rect 4787 5014 4791 5015
rect 4787 5009 4791 5010
rect 4955 5014 4959 5015
rect 4955 5009 4959 5010
rect 4971 5014 4975 5015
rect 4971 5009 4975 5010
rect 5155 5014 5159 5015
rect 5155 5009 5159 5010
rect 5179 5014 5183 5015
rect 5179 5009 5183 5010
rect 5339 5014 5343 5015
rect 5339 5009 5343 5010
rect 5411 5014 5415 5015
rect 5411 5009 5415 5010
rect 5515 5014 5519 5015
rect 5515 5009 5519 5010
rect 5663 5014 5667 5015
rect 5663 5009 5667 5010
rect 1975 5006 1979 5007
rect 1934 5004 1940 5005
rect 110 5000 111 5004
rect 115 5000 116 5004
rect 110 4999 116 5000
rect 146 5003 152 5004
rect 146 4999 147 5003
rect 151 4999 152 5003
rect 146 4998 152 4999
rect 338 5003 344 5004
rect 338 4999 339 5003
rect 343 4999 344 5003
rect 338 4998 344 4999
rect 530 5003 536 5004
rect 530 4999 531 5003
rect 535 4999 536 5003
rect 530 4998 536 4999
rect 730 5003 736 5004
rect 730 4999 731 5003
rect 735 4999 736 5003
rect 730 4998 736 4999
rect 930 5003 936 5004
rect 930 4999 931 5003
rect 935 4999 936 5003
rect 930 4998 936 4999
rect 1130 5003 1136 5004
rect 1130 4999 1131 5003
rect 1135 4999 1136 5003
rect 1934 5000 1935 5004
rect 1939 5000 1940 5004
rect 1975 5001 1979 5002
rect 2023 5006 2027 5007
rect 2023 5001 2027 5002
rect 2167 5006 2171 5007
rect 2167 5001 2171 5002
rect 2335 5006 2339 5007
rect 2335 5001 2339 5002
rect 2351 5006 2355 5007
rect 2351 5001 2355 5002
rect 2519 5006 2523 5007
rect 2519 5001 2523 5002
rect 2543 5006 2547 5007
rect 2543 5001 2547 5002
rect 2719 5006 2723 5007
rect 2719 5001 2723 5002
rect 2751 5006 2755 5007
rect 2751 5001 2755 5002
rect 2943 5006 2947 5007
rect 2943 5001 2947 5002
rect 2967 5006 2971 5007
rect 2967 5001 2971 5002
rect 3183 5006 3187 5007
rect 3183 5001 3187 5002
rect 3191 5006 3195 5007
rect 3191 5001 3195 5002
rect 3447 5006 3451 5007
rect 3447 5001 3451 5002
rect 3679 5006 3683 5007
rect 3679 5001 3683 5002
rect 3799 5006 3803 5007
rect 3799 5001 3803 5002
rect 1934 4999 1940 5000
rect 1130 4998 1136 4999
rect 174 4988 180 4989
rect 110 4987 116 4988
rect 110 4983 111 4987
rect 115 4983 116 4987
rect 174 4984 175 4988
rect 179 4984 180 4988
rect 174 4983 180 4984
rect 366 4988 372 4989
rect 366 4984 367 4988
rect 371 4984 372 4988
rect 366 4983 372 4984
rect 558 4988 564 4989
rect 558 4984 559 4988
rect 563 4984 564 4988
rect 558 4983 564 4984
rect 758 4988 764 4989
rect 758 4984 759 4988
rect 763 4984 764 4988
rect 758 4983 764 4984
rect 958 4988 964 4989
rect 958 4984 959 4988
rect 963 4984 964 4988
rect 958 4983 964 4984
rect 1158 4988 1164 4989
rect 1158 4984 1159 4988
rect 1163 4984 1164 4988
rect 1158 4983 1164 4984
rect 1934 4987 1940 4988
rect 1934 4983 1935 4987
rect 1939 4983 1940 4987
rect 110 4982 116 4983
rect 112 4947 114 4982
rect 176 4947 178 4983
rect 368 4947 370 4983
rect 560 4947 562 4983
rect 760 4947 762 4983
rect 960 4947 962 4983
rect 1160 4947 1162 4983
rect 1934 4982 1940 4983
rect 1936 4947 1938 4982
rect 1976 4978 1978 5001
rect 1974 4977 1980 4978
rect 2024 4977 2026 5001
rect 2168 4977 2170 5001
rect 2352 4977 2354 5001
rect 2544 4977 2546 5001
rect 2752 4977 2754 5001
rect 2968 4977 2970 5001
rect 3184 4977 3186 5001
rect 3800 4978 3802 5001
rect 3798 4977 3804 4978
rect 1974 4973 1975 4977
rect 1979 4973 1980 4977
rect 1974 4972 1980 4973
rect 2022 4976 2028 4977
rect 2022 4972 2023 4976
rect 2027 4972 2028 4976
rect 2022 4971 2028 4972
rect 2166 4976 2172 4977
rect 2166 4972 2167 4976
rect 2171 4972 2172 4976
rect 2166 4971 2172 4972
rect 2350 4976 2356 4977
rect 2350 4972 2351 4976
rect 2355 4972 2356 4976
rect 2350 4971 2356 4972
rect 2542 4976 2548 4977
rect 2542 4972 2543 4976
rect 2547 4972 2548 4976
rect 2542 4971 2548 4972
rect 2750 4976 2756 4977
rect 2750 4972 2751 4976
rect 2755 4972 2756 4976
rect 2750 4971 2756 4972
rect 2966 4976 2972 4977
rect 2966 4972 2967 4976
rect 2971 4972 2972 4976
rect 2966 4971 2972 4972
rect 3182 4976 3188 4977
rect 3182 4972 3183 4976
rect 3187 4972 3188 4976
rect 3798 4973 3799 4977
rect 3803 4973 3804 4977
rect 3798 4972 3804 4973
rect 3182 4971 3188 4972
rect 1994 4961 2000 4962
rect 1974 4960 1980 4961
rect 1974 4956 1975 4960
rect 1979 4956 1980 4960
rect 1994 4957 1995 4961
rect 1999 4957 2000 4961
rect 1994 4956 2000 4957
rect 2138 4961 2144 4962
rect 2138 4957 2139 4961
rect 2143 4957 2144 4961
rect 2138 4956 2144 4957
rect 2322 4961 2328 4962
rect 2322 4957 2323 4961
rect 2327 4957 2328 4961
rect 2322 4956 2328 4957
rect 2514 4961 2520 4962
rect 2514 4957 2515 4961
rect 2519 4957 2520 4961
rect 2514 4956 2520 4957
rect 2722 4961 2728 4962
rect 2722 4957 2723 4961
rect 2727 4957 2728 4961
rect 2722 4956 2728 4957
rect 2938 4961 2944 4962
rect 2938 4957 2939 4961
rect 2943 4957 2944 4961
rect 2938 4956 2944 4957
rect 3154 4961 3160 4962
rect 3154 4957 3155 4961
rect 3159 4957 3160 4961
rect 3154 4956 3160 4957
rect 3798 4960 3804 4961
rect 3798 4956 3799 4960
rect 3803 4956 3804 4960
rect 1974 4955 1980 4956
rect 111 4946 115 4947
rect 111 4941 115 4942
rect 159 4946 163 4947
rect 159 4941 163 4942
rect 175 4946 179 4947
rect 175 4941 179 4942
rect 367 4946 371 4947
rect 367 4941 371 4942
rect 391 4946 395 4947
rect 391 4941 395 4942
rect 559 4946 563 4947
rect 559 4941 563 4942
rect 647 4946 651 4947
rect 647 4941 651 4942
rect 759 4946 763 4947
rect 759 4941 763 4942
rect 895 4946 899 4947
rect 895 4941 899 4942
rect 959 4946 963 4947
rect 959 4941 963 4942
rect 1135 4946 1139 4947
rect 1135 4941 1139 4942
rect 1159 4946 1163 4947
rect 1159 4941 1163 4942
rect 1367 4946 1371 4947
rect 1367 4941 1371 4942
rect 1599 4946 1603 4947
rect 1599 4941 1603 4942
rect 1815 4946 1819 4947
rect 1815 4941 1819 4942
rect 1935 4946 1939 4947
rect 1935 4941 1939 4942
rect 112 4918 114 4941
rect 110 4917 116 4918
rect 160 4917 162 4941
rect 392 4917 394 4941
rect 648 4917 650 4941
rect 896 4917 898 4941
rect 1136 4917 1138 4941
rect 1368 4917 1370 4941
rect 1600 4917 1602 4941
rect 1816 4917 1818 4941
rect 1936 4918 1938 4941
rect 1934 4917 1940 4918
rect 110 4913 111 4917
rect 115 4913 116 4917
rect 110 4912 116 4913
rect 158 4916 164 4917
rect 158 4912 159 4916
rect 163 4912 164 4916
rect 158 4911 164 4912
rect 390 4916 396 4917
rect 390 4912 391 4916
rect 395 4912 396 4916
rect 390 4911 396 4912
rect 646 4916 652 4917
rect 646 4912 647 4916
rect 651 4912 652 4916
rect 646 4911 652 4912
rect 894 4916 900 4917
rect 894 4912 895 4916
rect 899 4912 900 4916
rect 894 4911 900 4912
rect 1134 4916 1140 4917
rect 1134 4912 1135 4916
rect 1139 4912 1140 4916
rect 1134 4911 1140 4912
rect 1366 4916 1372 4917
rect 1366 4912 1367 4916
rect 1371 4912 1372 4916
rect 1366 4911 1372 4912
rect 1598 4916 1604 4917
rect 1598 4912 1599 4916
rect 1603 4912 1604 4916
rect 1598 4911 1604 4912
rect 1814 4916 1820 4917
rect 1814 4912 1815 4916
rect 1819 4912 1820 4916
rect 1934 4913 1935 4917
rect 1939 4913 1940 4917
rect 1934 4912 1940 4913
rect 1814 4911 1820 4912
rect 130 4901 136 4902
rect 110 4900 116 4901
rect 110 4896 111 4900
rect 115 4896 116 4900
rect 130 4897 131 4901
rect 135 4897 136 4901
rect 130 4896 136 4897
rect 362 4901 368 4902
rect 362 4897 363 4901
rect 367 4897 368 4901
rect 362 4896 368 4897
rect 618 4901 624 4902
rect 618 4897 619 4901
rect 623 4897 624 4901
rect 618 4896 624 4897
rect 866 4901 872 4902
rect 866 4897 867 4901
rect 871 4897 872 4901
rect 866 4896 872 4897
rect 1106 4901 1112 4902
rect 1106 4897 1107 4901
rect 1111 4897 1112 4901
rect 1106 4896 1112 4897
rect 1338 4901 1344 4902
rect 1338 4897 1339 4901
rect 1343 4897 1344 4901
rect 1338 4896 1344 4897
rect 1570 4901 1576 4902
rect 1570 4897 1571 4901
rect 1575 4897 1576 4901
rect 1570 4896 1576 4897
rect 1786 4901 1792 4902
rect 1786 4897 1787 4901
rect 1791 4897 1792 4901
rect 1786 4896 1792 4897
rect 1934 4900 1940 4901
rect 1934 4896 1935 4900
rect 1939 4896 1940 4900
rect 110 4895 116 4896
rect 112 4835 114 4895
rect 132 4835 134 4896
rect 364 4835 366 4896
rect 620 4835 622 4896
rect 868 4835 870 4896
rect 1108 4835 1110 4896
rect 1340 4835 1342 4896
rect 1572 4835 1574 4896
rect 1788 4835 1790 4896
rect 1934 4895 1940 4896
rect 1936 4835 1938 4895
rect 1976 4887 1978 4955
rect 1996 4887 1998 4956
rect 2140 4887 2142 4956
rect 2324 4887 2326 4956
rect 2516 4887 2518 4956
rect 2724 4887 2726 4956
rect 2940 4887 2942 4956
rect 3156 4887 3158 4956
rect 3798 4955 3804 4956
rect 3800 4887 3802 4955
rect 3840 4949 3842 5009
rect 3838 4948 3844 4949
rect 3860 4948 3862 5009
rect 3996 4948 3998 5009
rect 4132 4948 4134 5009
rect 4284 4948 4286 5009
rect 4444 4948 4446 5009
rect 4612 4948 4614 5009
rect 4788 4948 4790 5009
rect 4972 4948 4974 5009
rect 5156 4948 5158 5009
rect 5340 4948 5342 5009
rect 5516 4948 5518 5009
rect 5664 4949 5666 5009
rect 5662 4948 5668 4949
rect 3838 4944 3839 4948
rect 3843 4944 3844 4948
rect 3838 4943 3844 4944
rect 3858 4947 3864 4948
rect 3858 4943 3859 4947
rect 3863 4943 3864 4947
rect 3858 4942 3864 4943
rect 3994 4947 4000 4948
rect 3994 4943 3995 4947
rect 3999 4943 4000 4947
rect 3994 4942 4000 4943
rect 4130 4947 4136 4948
rect 4130 4943 4131 4947
rect 4135 4943 4136 4947
rect 4130 4942 4136 4943
rect 4282 4947 4288 4948
rect 4282 4943 4283 4947
rect 4287 4943 4288 4947
rect 4282 4942 4288 4943
rect 4442 4947 4448 4948
rect 4442 4943 4443 4947
rect 4447 4943 4448 4947
rect 4442 4942 4448 4943
rect 4610 4947 4616 4948
rect 4610 4943 4611 4947
rect 4615 4943 4616 4947
rect 4610 4942 4616 4943
rect 4786 4947 4792 4948
rect 4786 4943 4787 4947
rect 4791 4943 4792 4947
rect 4786 4942 4792 4943
rect 4970 4947 4976 4948
rect 4970 4943 4971 4947
rect 4975 4943 4976 4947
rect 4970 4942 4976 4943
rect 5154 4947 5160 4948
rect 5154 4943 5155 4947
rect 5159 4943 5160 4947
rect 5154 4942 5160 4943
rect 5338 4947 5344 4948
rect 5338 4943 5339 4947
rect 5343 4943 5344 4947
rect 5338 4942 5344 4943
rect 5514 4947 5520 4948
rect 5514 4943 5515 4947
rect 5519 4943 5520 4947
rect 5662 4944 5663 4948
rect 5667 4944 5668 4948
rect 5662 4943 5668 4944
rect 5514 4942 5520 4943
rect 3886 4932 3892 4933
rect 3838 4931 3844 4932
rect 3838 4927 3839 4931
rect 3843 4927 3844 4931
rect 3886 4928 3887 4932
rect 3891 4928 3892 4932
rect 3886 4927 3892 4928
rect 4022 4932 4028 4933
rect 4022 4928 4023 4932
rect 4027 4928 4028 4932
rect 4022 4927 4028 4928
rect 4158 4932 4164 4933
rect 4158 4928 4159 4932
rect 4163 4928 4164 4932
rect 4158 4927 4164 4928
rect 4310 4932 4316 4933
rect 4310 4928 4311 4932
rect 4315 4928 4316 4932
rect 4310 4927 4316 4928
rect 4470 4932 4476 4933
rect 4470 4928 4471 4932
rect 4475 4928 4476 4932
rect 4470 4927 4476 4928
rect 4638 4932 4644 4933
rect 4638 4928 4639 4932
rect 4643 4928 4644 4932
rect 4638 4927 4644 4928
rect 4814 4932 4820 4933
rect 4814 4928 4815 4932
rect 4819 4928 4820 4932
rect 4814 4927 4820 4928
rect 4998 4932 5004 4933
rect 4998 4928 4999 4932
rect 5003 4928 5004 4932
rect 4998 4927 5004 4928
rect 5182 4932 5188 4933
rect 5182 4928 5183 4932
rect 5187 4928 5188 4932
rect 5182 4927 5188 4928
rect 5366 4932 5372 4933
rect 5366 4928 5367 4932
rect 5371 4928 5372 4932
rect 5366 4927 5372 4928
rect 5542 4932 5548 4933
rect 5542 4928 5543 4932
rect 5547 4928 5548 4932
rect 5542 4927 5548 4928
rect 5662 4931 5668 4932
rect 5662 4927 5663 4931
rect 5667 4927 5668 4931
rect 3838 4926 3844 4927
rect 3840 4887 3842 4926
rect 3888 4887 3890 4927
rect 4024 4887 4026 4927
rect 4160 4887 4162 4927
rect 4312 4887 4314 4927
rect 4472 4887 4474 4927
rect 4640 4887 4642 4927
rect 4816 4887 4818 4927
rect 5000 4887 5002 4927
rect 5184 4887 5186 4927
rect 5368 4887 5370 4927
rect 5544 4887 5546 4927
rect 5662 4926 5668 4927
rect 5664 4887 5666 4926
rect 1975 4886 1979 4887
rect 1975 4881 1979 4882
rect 1995 4886 1999 4887
rect 1995 4881 1999 4882
rect 2139 4886 2143 4887
rect 2139 4881 2143 4882
rect 2323 4886 2327 4887
rect 2323 4881 2327 4882
rect 2515 4886 2519 4887
rect 2515 4881 2519 4882
rect 2667 4886 2671 4887
rect 2667 4881 2671 4882
rect 2723 4886 2727 4887
rect 2723 4881 2727 4882
rect 2939 4886 2943 4887
rect 2939 4881 2943 4882
rect 3019 4886 3023 4887
rect 3019 4881 3023 4882
rect 3155 4886 3159 4887
rect 3155 4881 3159 4882
rect 3371 4886 3375 4887
rect 3371 4881 3375 4882
rect 3799 4886 3803 4887
rect 3799 4881 3803 4882
rect 3839 4886 3843 4887
rect 3839 4881 3843 4882
rect 3887 4886 3891 4887
rect 3887 4881 3891 4882
rect 3943 4886 3947 4887
rect 3943 4881 3947 4882
rect 4023 4886 4027 4887
rect 4023 4881 4027 4882
rect 4159 4886 4163 4887
rect 4159 4881 4163 4882
rect 4183 4886 4187 4887
rect 4183 4881 4187 4882
rect 4311 4886 4315 4887
rect 4311 4881 4315 4882
rect 4431 4886 4435 4887
rect 4431 4881 4435 4882
rect 4471 4886 4475 4887
rect 4471 4881 4475 4882
rect 4639 4886 4643 4887
rect 4639 4881 4643 4882
rect 4687 4886 4691 4887
rect 4687 4881 4691 4882
rect 4815 4886 4819 4887
rect 4815 4881 4819 4882
rect 4959 4886 4963 4887
rect 4959 4881 4963 4882
rect 4999 4886 5003 4887
rect 4999 4881 5003 4882
rect 5183 4886 5187 4887
rect 5183 4881 5187 4882
rect 5239 4886 5243 4887
rect 5239 4881 5243 4882
rect 5367 4886 5371 4887
rect 5367 4881 5371 4882
rect 5519 4886 5523 4887
rect 5519 4881 5523 4882
rect 5543 4886 5547 4887
rect 5543 4881 5547 4882
rect 5663 4886 5667 4887
rect 5663 4881 5667 4882
rect 111 4834 115 4835
rect 111 4829 115 4830
rect 131 4834 135 4835
rect 131 4829 135 4830
rect 363 4834 367 4835
rect 363 4829 367 4830
rect 475 4834 479 4835
rect 475 4829 479 4830
rect 619 4834 623 4835
rect 619 4829 623 4830
rect 859 4834 863 4835
rect 859 4829 863 4830
rect 867 4834 871 4835
rect 867 4829 871 4830
rect 1107 4834 1111 4835
rect 1107 4829 1111 4830
rect 1251 4834 1255 4835
rect 1251 4829 1255 4830
rect 1339 4834 1343 4835
rect 1339 4829 1343 4830
rect 1571 4834 1575 4835
rect 1571 4829 1575 4830
rect 1643 4834 1647 4835
rect 1643 4829 1647 4830
rect 1787 4834 1791 4835
rect 1787 4829 1791 4830
rect 1935 4834 1939 4835
rect 1935 4829 1939 4830
rect 112 4769 114 4829
rect 110 4768 116 4769
rect 132 4768 134 4829
rect 476 4768 478 4829
rect 860 4768 862 4829
rect 1252 4768 1254 4829
rect 1644 4768 1646 4829
rect 1936 4769 1938 4829
rect 1976 4821 1978 4881
rect 1974 4820 1980 4821
rect 1996 4820 1998 4881
rect 2324 4820 2326 4881
rect 2668 4820 2670 4881
rect 3020 4820 3022 4881
rect 3372 4820 3374 4881
rect 3800 4821 3802 4881
rect 3840 4858 3842 4881
rect 3838 4857 3844 4858
rect 3944 4857 3946 4881
rect 4184 4857 4186 4881
rect 4432 4857 4434 4881
rect 4688 4857 4690 4881
rect 4960 4857 4962 4881
rect 5240 4857 5242 4881
rect 5520 4857 5522 4881
rect 5664 4858 5666 4881
rect 5662 4857 5668 4858
rect 3838 4853 3839 4857
rect 3843 4853 3844 4857
rect 3838 4852 3844 4853
rect 3942 4856 3948 4857
rect 3942 4852 3943 4856
rect 3947 4852 3948 4856
rect 3942 4851 3948 4852
rect 4182 4856 4188 4857
rect 4182 4852 4183 4856
rect 4187 4852 4188 4856
rect 4182 4851 4188 4852
rect 4430 4856 4436 4857
rect 4430 4852 4431 4856
rect 4435 4852 4436 4856
rect 4430 4851 4436 4852
rect 4686 4856 4692 4857
rect 4686 4852 4687 4856
rect 4691 4852 4692 4856
rect 4686 4851 4692 4852
rect 4958 4856 4964 4857
rect 4958 4852 4959 4856
rect 4963 4852 4964 4856
rect 4958 4851 4964 4852
rect 5238 4856 5244 4857
rect 5238 4852 5239 4856
rect 5243 4852 5244 4856
rect 5238 4851 5244 4852
rect 5518 4856 5524 4857
rect 5518 4852 5519 4856
rect 5523 4852 5524 4856
rect 5662 4853 5663 4857
rect 5667 4853 5668 4857
rect 5662 4852 5668 4853
rect 5518 4851 5524 4852
rect 3914 4841 3920 4842
rect 3838 4840 3844 4841
rect 3838 4836 3839 4840
rect 3843 4836 3844 4840
rect 3914 4837 3915 4841
rect 3919 4837 3920 4841
rect 3914 4836 3920 4837
rect 4154 4841 4160 4842
rect 4154 4837 4155 4841
rect 4159 4837 4160 4841
rect 4154 4836 4160 4837
rect 4402 4841 4408 4842
rect 4402 4837 4403 4841
rect 4407 4837 4408 4841
rect 4402 4836 4408 4837
rect 4658 4841 4664 4842
rect 4658 4837 4659 4841
rect 4663 4837 4664 4841
rect 4658 4836 4664 4837
rect 4930 4841 4936 4842
rect 4930 4837 4931 4841
rect 4935 4837 4936 4841
rect 4930 4836 4936 4837
rect 5210 4841 5216 4842
rect 5210 4837 5211 4841
rect 5215 4837 5216 4841
rect 5210 4836 5216 4837
rect 5490 4841 5496 4842
rect 5490 4837 5491 4841
rect 5495 4837 5496 4841
rect 5490 4836 5496 4837
rect 5662 4840 5668 4841
rect 5662 4836 5663 4840
rect 5667 4836 5668 4840
rect 3838 4835 3844 4836
rect 3798 4820 3804 4821
rect 1974 4816 1975 4820
rect 1979 4816 1980 4820
rect 1974 4815 1980 4816
rect 1994 4819 2000 4820
rect 1994 4815 1995 4819
rect 1999 4815 2000 4819
rect 1994 4814 2000 4815
rect 2322 4819 2328 4820
rect 2322 4815 2323 4819
rect 2327 4815 2328 4819
rect 2322 4814 2328 4815
rect 2666 4819 2672 4820
rect 2666 4815 2667 4819
rect 2671 4815 2672 4819
rect 2666 4814 2672 4815
rect 3018 4819 3024 4820
rect 3018 4815 3019 4819
rect 3023 4815 3024 4819
rect 3018 4814 3024 4815
rect 3370 4819 3376 4820
rect 3370 4815 3371 4819
rect 3375 4815 3376 4819
rect 3798 4816 3799 4820
rect 3803 4816 3804 4820
rect 3798 4815 3804 4816
rect 3370 4814 3376 4815
rect 2022 4804 2028 4805
rect 1974 4803 1980 4804
rect 1974 4799 1975 4803
rect 1979 4799 1980 4803
rect 2022 4800 2023 4804
rect 2027 4800 2028 4804
rect 2022 4799 2028 4800
rect 2350 4804 2356 4805
rect 2350 4800 2351 4804
rect 2355 4800 2356 4804
rect 2350 4799 2356 4800
rect 2694 4804 2700 4805
rect 2694 4800 2695 4804
rect 2699 4800 2700 4804
rect 2694 4799 2700 4800
rect 3046 4804 3052 4805
rect 3046 4800 3047 4804
rect 3051 4800 3052 4804
rect 3046 4799 3052 4800
rect 3398 4804 3404 4805
rect 3398 4800 3399 4804
rect 3403 4800 3404 4804
rect 3398 4799 3404 4800
rect 3798 4803 3804 4804
rect 3798 4799 3799 4803
rect 3803 4799 3804 4803
rect 1974 4798 1980 4799
rect 1934 4768 1940 4769
rect 110 4764 111 4768
rect 115 4764 116 4768
rect 110 4763 116 4764
rect 130 4767 136 4768
rect 130 4763 131 4767
rect 135 4763 136 4767
rect 130 4762 136 4763
rect 474 4767 480 4768
rect 474 4763 475 4767
rect 479 4763 480 4767
rect 474 4762 480 4763
rect 858 4767 864 4768
rect 858 4763 859 4767
rect 863 4763 864 4767
rect 858 4762 864 4763
rect 1250 4767 1256 4768
rect 1250 4763 1251 4767
rect 1255 4763 1256 4767
rect 1250 4762 1256 4763
rect 1642 4767 1648 4768
rect 1642 4763 1643 4767
rect 1647 4763 1648 4767
rect 1934 4764 1935 4768
rect 1939 4764 1940 4768
rect 1934 4763 1940 4764
rect 1642 4762 1648 4763
rect 158 4752 164 4753
rect 110 4751 116 4752
rect 110 4747 111 4751
rect 115 4747 116 4751
rect 158 4748 159 4752
rect 163 4748 164 4752
rect 158 4747 164 4748
rect 502 4752 508 4753
rect 502 4748 503 4752
rect 507 4748 508 4752
rect 502 4747 508 4748
rect 886 4752 892 4753
rect 886 4748 887 4752
rect 891 4748 892 4752
rect 886 4747 892 4748
rect 1278 4752 1284 4753
rect 1278 4748 1279 4752
rect 1283 4748 1284 4752
rect 1278 4747 1284 4748
rect 1670 4752 1676 4753
rect 1670 4748 1671 4752
rect 1675 4748 1676 4752
rect 1670 4747 1676 4748
rect 1934 4751 1940 4752
rect 1934 4747 1935 4751
rect 1939 4747 1940 4751
rect 110 4746 116 4747
rect 112 4703 114 4746
rect 160 4703 162 4747
rect 504 4703 506 4747
rect 888 4703 890 4747
rect 1280 4703 1282 4747
rect 1672 4703 1674 4747
rect 1934 4746 1940 4747
rect 1936 4703 1938 4746
rect 1976 4727 1978 4798
rect 2024 4727 2026 4799
rect 2352 4727 2354 4799
rect 2696 4727 2698 4799
rect 3048 4727 3050 4799
rect 3400 4727 3402 4799
rect 3798 4798 3804 4799
rect 3800 4727 3802 4798
rect 3840 4767 3842 4835
rect 3916 4767 3918 4836
rect 4156 4767 4158 4836
rect 4404 4767 4406 4836
rect 4660 4767 4662 4836
rect 4932 4767 4934 4836
rect 5212 4767 5214 4836
rect 5492 4767 5494 4836
rect 5662 4835 5668 4836
rect 5664 4767 5666 4835
rect 3839 4766 3843 4767
rect 3839 4761 3843 4762
rect 3915 4766 3919 4767
rect 3915 4761 3919 4762
rect 3939 4766 3943 4767
rect 3939 4761 3943 4762
rect 4155 4766 4159 4767
rect 4155 4761 4159 4762
rect 4179 4766 4183 4767
rect 4179 4761 4183 4762
rect 4403 4766 4407 4767
rect 4403 4761 4407 4762
rect 4435 4766 4439 4767
rect 4435 4761 4439 4762
rect 4659 4766 4663 4767
rect 4659 4761 4663 4762
rect 4691 4766 4695 4767
rect 4691 4761 4695 4762
rect 4931 4766 4935 4767
rect 4931 4761 4935 4762
rect 4955 4766 4959 4767
rect 4955 4761 4959 4762
rect 5211 4766 5215 4767
rect 5211 4761 5215 4762
rect 5227 4766 5231 4767
rect 5227 4761 5231 4762
rect 5491 4766 5495 4767
rect 5491 4761 5495 4762
rect 5507 4766 5511 4767
rect 5507 4761 5511 4762
rect 5663 4766 5667 4767
rect 5663 4761 5667 4762
rect 1975 4726 1979 4727
rect 1975 4721 1979 4722
rect 2023 4726 2027 4727
rect 2023 4721 2027 4722
rect 2079 4726 2083 4727
rect 2079 4721 2083 4722
rect 2231 4726 2235 4727
rect 2231 4721 2235 4722
rect 2351 4726 2355 4727
rect 2351 4721 2355 4722
rect 2391 4726 2395 4727
rect 2391 4721 2395 4722
rect 2559 4726 2563 4727
rect 2559 4721 2563 4722
rect 2695 4726 2699 4727
rect 2695 4721 2699 4722
rect 2727 4726 2731 4727
rect 2727 4721 2731 4722
rect 2903 4726 2907 4727
rect 2903 4721 2907 4722
rect 3047 4726 3051 4727
rect 3047 4721 3051 4722
rect 3079 4726 3083 4727
rect 3079 4721 3083 4722
rect 3255 4726 3259 4727
rect 3255 4721 3259 4722
rect 3399 4726 3403 4727
rect 3399 4721 3403 4722
rect 3439 4726 3443 4727
rect 3439 4721 3443 4722
rect 3623 4726 3627 4727
rect 3623 4721 3627 4722
rect 3799 4726 3803 4727
rect 3799 4721 3803 4722
rect 111 4702 115 4703
rect 111 4697 115 4698
rect 159 4702 163 4703
rect 159 4697 163 4698
rect 295 4702 299 4703
rect 295 4697 299 4698
rect 431 4702 435 4703
rect 431 4697 435 4698
rect 503 4702 507 4703
rect 503 4697 507 4698
rect 567 4702 571 4703
rect 567 4697 571 4698
rect 703 4702 707 4703
rect 703 4697 707 4698
rect 887 4702 891 4703
rect 887 4697 891 4698
rect 1279 4702 1283 4703
rect 1279 4697 1283 4698
rect 1671 4702 1675 4703
rect 1671 4697 1675 4698
rect 1935 4702 1939 4703
rect 1976 4698 1978 4721
rect 1935 4697 1939 4698
rect 1974 4697 1980 4698
rect 2080 4697 2082 4721
rect 2232 4697 2234 4721
rect 2392 4697 2394 4721
rect 2560 4697 2562 4721
rect 2728 4697 2730 4721
rect 2904 4697 2906 4721
rect 3080 4697 3082 4721
rect 3256 4697 3258 4721
rect 3440 4697 3442 4721
rect 3624 4697 3626 4721
rect 3800 4698 3802 4721
rect 3840 4701 3842 4761
rect 3838 4700 3844 4701
rect 3940 4700 3942 4761
rect 4180 4700 4182 4761
rect 4436 4700 4438 4761
rect 4692 4700 4694 4761
rect 4956 4700 4958 4761
rect 5228 4700 5230 4761
rect 5508 4700 5510 4761
rect 5664 4701 5666 4761
rect 5662 4700 5668 4701
rect 3798 4697 3804 4698
rect 112 4674 114 4697
rect 110 4673 116 4674
rect 160 4673 162 4697
rect 296 4673 298 4697
rect 432 4673 434 4697
rect 568 4673 570 4697
rect 704 4673 706 4697
rect 1936 4674 1938 4697
rect 1974 4693 1975 4697
rect 1979 4693 1980 4697
rect 1974 4692 1980 4693
rect 2078 4696 2084 4697
rect 2078 4692 2079 4696
rect 2083 4692 2084 4696
rect 2078 4691 2084 4692
rect 2230 4696 2236 4697
rect 2230 4692 2231 4696
rect 2235 4692 2236 4696
rect 2230 4691 2236 4692
rect 2390 4696 2396 4697
rect 2390 4692 2391 4696
rect 2395 4692 2396 4696
rect 2390 4691 2396 4692
rect 2558 4696 2564 4697
rect 2558 4692 2559 4696
rect 2563 4692 2564 4696
rect 2558 4691 2564 4692
rect 2726 4696 2732 4697
rect 2726 4692 2727 4696
rect 2731 4692 2732 4696
rect 2726 4691 2732 4692
rect 2902 4696 2908 4697
rect 2902 4692 2903 4696
rect 2907 4692 2908 4696
rect 2902 4691 2908 4692
rect 3078 4696 3084 4697
rect 3078 4692 3079 4696
rect 3083 4692 3084 4696
rect 3078 4691 3084 4692
rect 3254 4696 3260 4697
rect 3254 4692 3255 4696
rect 3259 4692 3260 4696
rect 3254 4691 3260 4692
rect 3438 4696 3444 4697
rect 3438 4692 3439 4696
rect 3443 4692 3444 4696
rect 3438 4691 3444 4692
rect 3622 4696 3628 4697
rect 3622 4692 3623 4696
rect 3627 4692 3628 4696
rect 3798 4693 3799 4697
rect 3803 4693 3804 4697
rect 3838 4696 3839 4700
rect 3843 4696 3844 4700
rect 3838 4695 3844 4696
rect 3938 4699 3944 4700
rect 3938 4695 3939 4699
rect 3943 4695 3944 4699
rect 3938 4694 3944 4695
rect 4178 4699 4184 4700
rect 4178 4695 4179 4699
rect 4183 4695 4184 4699
rect 4178 4694 4184 4695
rect 4434 4699 4440 4700
rect 4434 4695 4435 4699
rect 4439 4695 4440 4699
rect 4434 4694 4440 4695
rect 4690 4699 4696 4700
rect 4690 4695 4691 4699
rect 4695 4695 4696 4699
rect 4690 4694 4696 4695
rect 4954 4699 4960 4700
rect 4954 4695 4955 4699
rect 4959 4695 4960 4699
rect 4954 4694 4960 4695
rect 5226 4699 5232 4700
rect 5226 4695 5227 4699
rect 5231 4695 5232 4699
rect 5226 4694 5232 4695
rect 5506 4699 5512 4700
rect 5506 4695 5507 4699
rect 5511 4695 5512 4699
rect 5662 4696 5663 4700
rect 5667 4696 5668 4700
rect 5662 4695 5668 4696
rect 5506 4694 5512 4695
rect 3798 4692 3804 4693
rect 3622 4691 3628 4692
rect 3966 4684 3972 4685
rect 3838 4683 3844 4684
rect 2050 4681 2056 4682
rect 1974 4680 1980 4681
rect 1974 4676 1975 4680
rect 1979 4676 1980 4680
rect 2050 4677 2051 4681
rect 2055 4677 2056 4681
rect 2050 4676 2056 4677
rect 2202 4681 2208 4682
rect 2202 4677 2203 4681
rect 2207 4677 2208 4681
rect 2202 4676 2208 4677
rect 2362 4681 2368 4682
rect 2362 4677 2363 4681
rect 2367 4677 2368 4681
rect 2362 4676 2368 4677
rect 2530 4681 2536 4682
rect 2530 4677 2531 4681
rect 2535 4677 2536 4681
rect 2530 4676 2536 4677
rect 2698 4681 2704 4682
rect 2698 4677 2699 4681
rect 2703 4677 2704 4681
rect 2698 4676 2704 4677
rect 2874 4681 2880 4682
rect 2874 4677 2875 4681
rect 2879 4677 2880 4681
rect 2874 4676 2880 4677
rect 3050 4681 3056 4682
rect 3050 4677 3051 4681
rect 3055 4677 3056 4681
rect 3050 4676 3056 4677
rect 3226 4681 3232 4682
rect 3226 4677 3227 4681
rect 3231 4677 3232 4681
rect 3226 4676 3232 4677
rect 3410 4681 3416 4682
rect 3410 4677 3411 4681
rect 3415 4677 3416 4681
rect 3410 4676 3416 4677
rect 3594 4681 3600 4682
rect 3594 4677 3595 4681
rect 3599 4677 3600 4681
rect 3594 4676 3600 4677
rect 3798 4680 3804 4681
rect 3798 4676 3799 4680
rect 3803 4676 3804 4680
rect 3838 4679 3839 4683
rect 3843 4679 3844 4683
rect 3966 4680 3967 4684
rect 3971 4680 3972 4684
rect 3966 4679 3972 4680
rect 4206 4684 4212 4685
rect 4206 4680 4207 4684
rect 4211 4680 4212 4684
rect 4206 4679 4212 4680
rect 4462 4684 4468 4685
rect 4462 4680 4463 4684
rect 4467 4680 4468 4684
rect 4462 4679 4468 4680
rect 4718 4684 4724 4685
rect 4718 4680 4719 4684
rect 4723 4680 4724 4684
rect 4718 4679 4724 4680
rect 4982 4684 4988 4685
rect 4982 4680 4983 4684
rect 4987 4680 4988 4684
rect 4982 4679 4988 4680
rect 5254 4684 5260 4685
rect 5254 4680 5255 4684
rect 5259 4680 5260 4684
rect 5254 4679 5260 4680
rect 5534 4684 5540 4685
rect 5534 4680 5535 4684
rect 5539 4680 5540 4684
rect 5534 4679 5540 4680
rect 5662 4683 5668 4684
rect 5662 4679 5663 4683
rect 5667 4679 5668 4683
rect 3838 4678 3844 4679
rect 1974 4675 1980 4676
rect 1934 4673 1940 4674
rect 110 4669 111 4673
rect 115 4669 116 4673
rect 110 4668 116 4669
rect 158 4672 164 4673
rect 158 4668 159 4672
rect 163 4668 164 4672
rect 158 4667 164 4668
rect 294 4672 300 4673
rect 294 4668 295 4672
rect 299 4668 300 4672
rect 294 4667 300 4668
rect 430 4672 436 4673
rect 430 4668 431 4672
rect 435 4668 436 4672
rect 430 4667 436 4668
rect 566 4672 572 4673
rect 566 4668 567 4672
rect 571 4668 572 4672
rect 566 4667 572 4668
rect 702 4672 708 4673
rect 702 4668 703 4672
rect 707 4668 708 4672
rect 1934 4669 1935 4673
rect 1939 4669 1940 4673
rect 1934 4668 1940 4669
rect 702 4667 708 4668
rect 130 4657 136 4658
rect 110 4656 116 4657
rect 110 4652 111 4656
rect 115 4652 116 4656
rect 130 4653 131 4657
rect 135 4653 136 4657
rect 130 4652 136 4653
rect 266 4657 272 4658
rect 266 4653 267 4657
rect 271 4653 272 4657
rect 266 4652 272 4653
rect 402 4657 408 4658
rect 402 4653 403 4657
rect 407 4653 408 4657
rect 402 4652 408 4653
rect 538 4657 544 4658
rect 538 4653 539 4657
rect 543 4653 544 4657
rect 538 4652 544 4653
rect 674 4657 680 4658
rect 674 4653 675 4657
rect 679 4653 680 4657
rect 674 4652 680 4653
rect 1934 4656 1940 4657
rect 1934 4652 1935 4656
rect 1939 4652 1940 4656
rect 110 4651 116 4652
rect 112 4575 114 4651
rect 132 4575 134 4652
rect 268 4575 270 4652
rect 404 4575 406 4652
rect 540 4575 542 4652
rect 676 4575 678 4652
rect 1934 4651 1940 4652
rect 1936 4575 1938 4651
rect 1976 4611 1978 4675
rect 2052 4611 2054 4676
rect 2204 4611 2206 4676
rect 2364 4611 2366 4676
rect 2532 4611 2534 4676
rect 2700 4611 2702 4676
rect 2876 4611 2878 4676
rect 3052 4611 3054 4676
rect 3228 4611 3230 4676
rect 3412 4611 3414 4676
rect 3596 4611 3598 4676
rect 3798 4675 3804 4676
rect 3800 4611 3802 4675
rect 3840 4651 3842 4678
rect 3968 4651 3970 4679
rect 4208 4651 4210 4679
rect 4464 4651 4466 4679
rect 4720 4651 4722 4679
rect 4984 4651 4986 4679
rect 5256 4651 5258 4679
rect 5536 4651 5538 4679
rect 5662 4678 5668 4679
rect 5664 4651 5666 4678
rect 3839 4650 3843 4651
rect 3839 4645 3843 4646
rect 3967 4650 3971 4651
rect 3967 4645 3971 4646
rect 4175 4650 4179 4651
rect 4175 4645 4179 4646
rect 4207 4650 4211 4651
rect 4207 4645 4211 4646
rect 4455 4650 4459 4651
rect 4455 4645 4459 4646
rect 4463 4650 4467 4651
rect 4463 4645 4467 4646
rect 4719 4650 4723 4651
rect 4719 4645 4723 4646
rect 4735 4650 4739 4651
rect 4735 4645 4739 4646
rect 4983 4650 4987 4651
rect 4983 4645 4987 4646
rect 5015 4650 5019 4651
rect 5015 4645 5019 4646
rect 5255 4650 5259 4651
rect 5255 4645 5259 4646
rect 5303 4650 5307 4651
rect 5303 4645 5307 4646
rect 5535 4650 5539 4651
rect 5535 4645 5539 4646
rect 5663 4650 5667 4651
rect 5663 4645 5667 4646
rect 3840 4622 3842 4645
rect 3838 4621 3844 4622
rect 4176 4621 4178 4645
rect 4456 4621 4458 4645
rect 4736 4621 4738 4645
rect 5016 4621 5018 4645
rect 5304 4621 5306 4645
rect 5664 4622 5666 4645
rect 5662 4621 5668 4622
rect 3838 4617 3839 4621
rect 3843 4617 3844 4621
rect 3838 4616 3844 4617
rect 4174 4620 4180 4621
rect 4174 4616 4175 4620
rect 4179 4616 4180 4620
rect 4174 4615 4180 4616
rect 4454 4620 4460 4621
rect 4454 4616 4455 4620
rect 4459 4616 4460 4620
rect 4454 4615 4460 4616
rect 4734 4620 4740 4621
rect 4734 4616 4735 4620
rect 4739 4616 4740 4620
rect 4734 4615 4740 4616
rect 5014 4620 5020 4621
rect 5014 4616 5015 4620
rect 5019 4616 5020 4620
rect 5014 4615 5020 4616
rect 5302 4620 5308 4621
rect 5302 4616 5303 4620
rect 5307 4616 5308 4620
rect 5662 4617 5663 4621
rect 5667 4617 5668 4621
rect 5662 4616 5668 4617
rect 5302 4615 5308 4616
rect 1975 4610 1979 4611
rect 1975 4605 1979 4606
rect 2051 4610 2055 4611
rect 2051 4605 2055 4606
rect 2123 4610 2127 4611
rect 2123 4605 2127 4606
rect 2203 4610 2207 4611
rect 2203 4605 2207 4606
rect 2275 4610 2279 4611
rect 2275 4605 2279 4606
rect 2363 4610 2367 4611
rect 2363 4605 2367 4606
rect 2443 4610 2447 4611
rect 2443 4605 2447 4606
rect 2531 4610 2535 4611
rect 2531 4605 2535 4606
rect 2611 4610 2615 4611
rect 2611 4605 2615 4606
rect 2699 4610 2703 4611
rect 2699 4605 2703 4606
rect 2787 4610 2791 4611
rect 2787 4605 2791 4606
rect 2875 4610 2879 4611
rect 2875 4605 2879 4606
rect 2963 4610 2967 4611
rect 2963 4605 2967 4606
rect 3051 4610 3055 4611
rect 3051 4605 3055 4606
rect 3139 4610 3143 4611
rect 3139 4605 3143 4606
rect 3227 4610 3231 4611
rect 3227 4605 3231 4606
rect 3315 4610 3319 4611
rect 3315 4605 3319 4606
rect 3411 4610 3415 4611
rect 3411 4605 3415 4606
rect 3491 4610 3495 4611
rect 3491 4605 3495 4606
rect 3595 4610 3599 4611
rect 3595 4605 3599 4606
rect 3651 4610 3655 4611
rect 3651 4605 3655 4606
rect 3799 4610 3803 4611
rect 3799 4605 3803 4606
rect 4146 4605 4152 4606
rect 111 4574 115 4575
rect 111 4569 115 4570
rect 131 4574 135 4575
rect 131 4569 135 4570
rect 267 4574 271 4575
rect 267 4569 271 4570
rect 291 4574 295 4575
rect 291 4569 295 4570
rect 403 4574 407 4575
rect 403 4569 407 4570
rect 427 4574 431 4575
rect 427 4569 431 4570
rect 539 4574 543 4575
rect 539 4569 543 4570
rect 563 4574 567 4575
rect 563 4569 567 4570
rect 675 4574 679 4575
rect 675 4569 679 4570
rect 699 4574 703 4575
rect 699 4569 703 4570
rect 835 4574 839 4575
rect 835 4569 839 4570
rect 1935 4574 1939 4575
rect 1935 4569 1939 4570
rect 112 4509 114 4569
rect 110 4508 116 4509
rect 292 4508 294 4569
rect 428 4508 430 4569
rect 564 4508 566 4569
rect 700 4508 702 4569
rect 836 4508 838 4569
rect 1936 4509 1938 4569
rect 1976 4545 1978 4605
rect 1974 4544 1980 4545
rect 2124 4544 2126 4605
rect 2276 4544 2278 4605
rect 2444 4544 2446 4605
rect 2612 4544 2614 4605
rect 2788 4544 2790 4605
rect 2964 4544 2966 4605
rect 3140 4544 3142 4605
rect 3316 4544 3318 4605
rect 3492 4544 3494 4605
rect 3652 4544 3654 4605
rect 3800 4545 3802 4605
rect 3838 4604 3844 4605
rect 3838 4600 3839 4604
rect 3843 4600 3844 4604
rect 4146 4601 4147 4605
rect 4151 4601 4152 4605
rect 4146 4600 4152 4601
rect 4426 4605 4432 4606
rect 4426 4601 4427 4605
rect 4431 4601 4432 4605
rect 4426 4600 4432 4601
rect 4706 4605 4712 4606
rect 4706 4601 4707 4605
rect 4711 4601 4712 4605
rect 4706 4600 4712 4601
rect 4986 4605 4992 4606
rect 4986 4601 4987 4605
rect 4991 4601 4992 4605
rect 4986 4600 4992 4601
rect 5274 4605 5280 4606
rect 5274 4601 5275 4605
rect 5279 4601 5280 4605
rect 5274 4600 5280 4601
rect 5662 4604 5668 4605
rect 5662 4600 5663 4604
rect 5667 4600 5668 4604
rect 3838 4599 3844 4600
rect 3798 4544 3804 4545
rect 1974 4540 1975 4544
rect 1979 4540 1980 4544
rect 1974 4539 1980 4540
rect 2122 4543 2128 4544
rect 2122 4539 2123 4543
rect 2127 4539 2128 4543
rect 2122 4538 2128 4539
rect 2274 4543 2280 4544
rect 2274 4539 2275 4543
rect 2279 4539 2280 4543
rect 2274 4538 2280 4539
rect 2442 4543 2448 4544
rect 2442 4539 2443 4543
rect 2447 4539 2448 4543
rect 2442 4538 2448 4539
rect 2610 4543 2616 4544
rect 2610 4539 2611 4543
rect 2615 4539 2616 4543
rect 2610 4538 2616 4539
rect 2786 4543 2792 4544
rect 2786 4539 2787 4543
rect 2791 4539 2792 4543
rect 2786 4538 2792 4539
rect 2962 4543 2968 4544
rect 2962 4539 2963 4543
rect 2967 4539 2968 4543
rect 2962 4538 2968 4539
rect 3138 4543 3144 4544
rect 3138 4539 3139 4543
rect 3143 4539 3144 4543
rect 3138 4538 3144 4539
rect 3314 4543 3320 4544
rect 3314 4539 3315 4543
rect 3319 4539 3320 4543
rect 3314 4538 3320 4539
rect 3490 4543 3496 4544
rect 3490 4539 3491 4543
rect 3495 4539 3496 4543
rect 3490 4538 3496 4539
rect 3650 4543 3656 4544
rect 3650 4539 3651 4543
rect 3655 4539 3656 4543
rect 3798 4540 3799 4544
rect 3803 4540 3804 4544
rect 3798 4539 3804 4540
rect 3650 4538 3656 4539
rect 3840 4535 3842 4599
rect 4148 4535 4150 4600
rect 4428 4535 4430 4600
rect 4708 4535 4710 4600
rect 4988 4535 4990 4600
rect 5276 4535 5278 4600
rect 5662 4599 5668 4600
rect 5664 4535 5666 4599
rect 3839 4534 3843 4535
rect 3839 4529 3843 4530
rect 3859 4534 3863 4535
rect 3859 4529 3863 4530
rect 4147 4534 4151 4535
rect 4147 4529 4151 4530
rect 4155 4534 4159 4535
rect 4155 4529 4159 4530
rect 4427 4534 4431 4535
rect 4427 4529 4431 4530
rect 4483 4534 4487 4535
rect 4483 4529 4487 4530
rect 4707 4534 4711 4535
rect 4707 4529 4711 4530
rect 4819 4534 4823 4535
rect 4819 4529 4823 4530
rect 4987 4534 4991 4535
rect 4987 4529 4991 4530
rect 5163 4534 5167 4535
rect 5163 4529 5167 4530
rect 5275 4534 5279 4535
rect 5275 4529 5279 4530
rect 5515 4534 5519 4535
rect 5515 4529 5519 4530
rect 5663 4534 5667 4535
rect 5663 4529 5667 4530
rect 2150 4528 2156 4529
rect 1974 4527 1980 4528
rect 1974 4523 1975 4527
rect 1979 4523 1980 4527
rect 2150 4524 2151 4528
rect 2155 4524 2156 4528
rect 2150 4523 2156 4524
rect 2302 4528 2308 4529
rect 2302 4524 2303 4528
rect 2307 4524 2308 4528
rect 2302 4523 2308 4524
rect 2470 4528 2476 4529
rect 2470 4524 2471 4528
rect 2475 4524 2476 4528
rect 2470 4523 2476 4524
rect 2638 4528 2644 4529
rect 2638 4524 2639 4528
rect 2643 4524 2644 4528
rect 2638 4523 2644 4524
rect 2814 4528 2820 4529
rect 2814 4524 2815 4528
rect 2819 4524 2820 4528
rect 2814 4523 2820 4524
rect 2990 4528 2996 4529
rect 2990 4524 2991 4528
rect 2995 4524 2996 4528
rect 2990 4523 2996 4524
rect 3166 4528 3172 4529
rect 3166 4524 3167 4528
rect 3171 4524 3172 4528
rect 3166 4523 3172 4524
rect 3342 4528 3348 4529
rect 3342 4524 3343 4528
rect 3347 4524 3348 4528
rect 3342 4523 3348 4524
rect 3518 4528 3524 4529
rect 3518 4524 3519 4528
rect 3523 4524 3524 4528
rect 3518 4523 3524 4524
rect 3678 4528 3684 4529
rect 3678 4524 3679 4528
rect 3683 4524 3684 4528
rect 3678 4523 3684 4524
rect 3798 4527 3804 4528
rect 3798 4523 3799 4527
rect 3803 4523 3804 4527
rect 1974 4522 1980 4523
rect 1934 4508 1940 4509
rect 110 4504 111 4508
rect 115 4504 116 4508
rect 110 4503 116 4504
rect 290 4507 296 4508
rect 290 4503 291 4507
rect 295 4503 296 4507
rect 290 4502 296 4503
rect 426 4507 432 4508
rect 426 4503 427 4507
rect 431 4503 432 4507
rect 426 4502 432 4503
rect 562 4507 568 4508
rect 562 4503 563 4507
rect 567 4503 568 4507
rect 562 4502 568 4503
rect 698 4507 704 4508
rect 698 4503 699 4507
rect 703 4503 704 4507
rect 698 4502 704 4503
rect 834 4507 840 4508
rect 834 4503 835 4507
rect 839 4503 840 4507
rect 1934 4504 1935 4508
rect 1939 4504 1940 4508
rect 1934 4503 1940 4504
rect 834 4502 840 4503
rect 318 4492 324 4493
rect 110 4491 116 4492
rect 110 4487 111 4491
rect 115 4487 116 4491
rect 318 4488 319 4492
rect 323 4488 324 4492
rect 318 4487 324 4488
rect 454 4492 460 4493
rect 454 4488 455 4492
rect 459 4488 460 4492
rect 454 4487 460 4488
rect 590 4492 596 4493
rect 590 4488 591 4492
rect 595 4488 596 4492
rect 590 4487 596 4488
rect 726 4492 732 4493
rect 726 4488 727 4492
rect 731 4488 732 4492
rect 726 4487 732 4488
rect 862 4492 868 4493
rect 862 4488 863 4492
rect 867 4488 868 4492
rect 862 4487 868 4488
rect 1934 4491 1940 4492
rect 1976 4491 1978 4522
rect 2152 4491 2154 4523
rect 2304 4491 2306 4523
rect 2472 4491 2474 4523
rect 2640 4491 2642 4523
rect 2816 4491 2818 4523
rect 2992 4491 2994 4523
rect 3168 4491 3170 4523
rect 3344 4491 3346 4523
rect 3520 4491 3522 4523
rect 3680 4491 3682 4523
rect 3798 4522 3804 4523
rect 3800 4491 3802 4522
rect 1934 4487 1935 4491
rect 1939 4487 1940 4491
rect 110 4486 116 4487
rect 112 4447 114 4486
rect 320 4447 322 4487
rect 456 4447 458 4487
rect 592 4447 594 4487
rect 728 4447 730 4487
rect 864 4447 866 4487
rect 1934 4486 1940 4487
rect 1975 4490 1979 4491
rect 1936 4447 1938 4486
rect 1975 4485 1979 4486
rect 2023 4490 2027 4491
rect 2023 4485 2027 4486
rect 2151 4490 2155 4491
rect 2151 4485 2155 4486
rect 2159 4490 2163 4491
rect 2159 4485 2163 4486
rect 2295 4490 2299 4491
rect 2295 4485 2299 4486
rect 2303 4490 2307 4491
rect 2303 4485 2307 4486
rect 2431 4490 2435 4491
rect 2431 4485 2435 4486
rect 2471 4490 2475 4491
rect 2471 4485 2475 4486
rect 2567 4490 2571 4491
rect 2567 4485 2571 4486
rect 2639 4490 2643 4491
rect 2639 4485 2643 4486
rect 2703 4490 2707 4491
rect 2703 4485 2707 4486
rect 2815 4490 2819 4491
rect 2815 4485 2819 4486
rect 2839 4490 2843 4491
rect 2839 4485 2843 4486
rect 2975 4490 2979 4491
rect 2975 4485 2979 4486
rect 2991 4490 2995 4491
rect 2991 4485 2995 4486
rect 3167 4490 3171 4491
rect 3167 4485 3171 4486
rect 3343 4490 3347 4491
rect 3343 4485 3347 4486
rect 3519 4490 3523 4491
rect 3519 4485 3523 4486
rect 3679 4490 3683 4491
rect 3679 4485 3683 4486
rect 3799 4490 3803 4491
rect 3799 4485 3803 4486
rect 1976 4462 1978 4485
rect 1974 4461 1980 4462
rect 2024 4461 2026 4485
rect 2160 4461 2162 4485
rect 2296 4461 2298 4485
rect 2432 4461 2434 4485
rect 2568 4461 2570 4485
rect 2704 4461 2706 4485
rect 2840 4461 2842 4485
rect 2976 4461 2978 4485
rect 3800 4462 3802 4485
rect 3840 4469 3842 4529
rect 3838 4468 3844 4469
rect 3860 4468 3862 4529
rect 4156 4468 4158 4529
rect 4484 4468 4486 4529
rect 4820 4468 4822 4529
rect 5164 4468 5166 4529
rect 5516 4468 5518 4529
rect 5664 4469 5666 4529
rect 5662 4468 5668 4469
rect 3838 4464 3839 4468
rect 3843 4464 3844 4468
rect 3838 4463 3844 4464
rect 3858 4467 3864 4468
rect 3858 4463 3859 4467
rect 3863 4463 3864 4467
rect 3858 4462 3864 4463
rect 4154 4467 4160 4468
rect 4154 4463 4155 4467
rect 4159 4463 4160 4467
rect 4154 4462 4160 4463
rect 4482 4467 4488 4468
rect 4482 4463 4483 4467
rect 4487 4463 4488 4467
rect 4482 4462 4488 4463
rect 4818 4467 4824 4468
rect 4818 4463 4819 4467
rect 4823 4463 4824 4467
rect 4818 4462 4824 4463
rect 5162 4467 5168 4468
rect 5162 4463 5163 4467
rect 5167 4463 5168 4467
rect 5162 4462 5168 4463
rect 5514 4467 5520 4468
rect 5514 4463 5515 4467
rect 5519 4463 5520 4467
rect 5662 4464 5663 4468
rect 5667 4464 5668 4468
rect 5662 4463 5668 4464
rect 5514 4462 5520 4463
rect 3798 4461 3804 4462
rect 1974 4457 1975 4461
rect 1979 4457 1980 4461
rect 1974 4456 1980 4457
rect 2022 4460 2028 4461
rect 2022 4456 2023 4460
rect 2027 4456 2028 4460
rect 2022 4455 2028 4456
rect 2158 4460 2164 4461
rect 2158 4456 2159 4460
rect 2163 4456 2164 4460
rect 2158 4455 2164 4456
rect 2294 4460 2300 4461
rect 2294 4456 2295 4460
rect 2299 4456 2300 4460
rect 2294 4455 2300 4456
rect 2430 4460 2436 4461
rect 2430 4456 2431 4460
rect 2435 4456 2436 4460
rect 2430 4455 2436 4456
rect 2566 4460 2572 4461
rect 2566 4456 2567 4460
rect 2571 4456 2572 4460
rect 2566 4455 2572 4456
rect 2702 4460 2708 4461
rect 2702 4456 2703 4460
rect 2707 4456 2708 4460
rect 2702 4455 2708 4456
rect 2838 4460 2844 4461
rect 2838 4456 2839 4460
rect 2843 4456 2844 4460
rect 2838 4455 2844 4456
rect 2974 4460 2980 4461
rect 2974 4456 2975 4460
rect 2979 4456 2980 4460
rect 3798 4457 3799 4461
rect 3803 4457 3804 4461
rect 3798 4456 3804 4457
rect 2974 4455 2980 4456
rect 3886 4452 3892 4453
rect 3838 4451 3844 4452
rect 3838 4447 3839 4451
rect 3843 4447 3844 4451
rect 3886 4448 3887 4452
rect 3891 4448 3892 4452
rect 3886 4447 3892 4448
rect 4182 4452 4188 4453
rect 4182 4448 4183 4452
rect 4187 4448 4188 4452
rect 4182 4447 4188 4448
rect 4510 4452 4516 4453
rect 4510 4448 4511 4452
rect 4515 4448 4516 4452
rect 4510 4447 4516 4448
rect 4846 4452 4852 4453
rect 4846 4448 4847 4452
rect 4851 4448 4852 4452
rect 4846 4447 4852 4448
rect 5190 4452 5196 4453
rect 5190 4448 5191 4452
rect 5195 4448 5196 4452
rect 5190 4447 5196 4448
rect 5542 4452 5548 4453
rect 5542 4448 5543 4452
rect 5547 4448 5548 4452
rect 5542 4447 5548 4448
rect 5662 4451 5668 4452
rect 5662 4447 5663 4451
rect 5667 4447 5668 4451
rect 111 4446 115 4447
rect 111 4441 115 4442
rect 319 4446 323 4447
rect 319 4441 323 4442
rect 455 4446 459 4447
rect 455 4441 459 4442
rect 519 4446 523 4447
rect 519 4441 523 4442
rect 591 4446 595 4447
rect 591 4441 595 4442
rect 727 4446 731 4447
rect 727 4441 731 4442
rect 743 4446 747 4447
rect 743 4441 747 4442
rect 863 4446 867 4447
rect 863 4441 867 4442
rect 991 4446 995 4447
rect 991 4441 995 4442
rect 1263 4446 1267 4447
rect 1263 4441 1267 4442
rect 1551 4446 1555 4447
rect 1551 4441 1555 4442
rect 1815 4446 1819 4447
rect 1815 4441 1819 4442
rect 1935 4446 1939 4447
rect 3838 4446 3844 4447
rect 1994 4445 2000 4446
rect 1935 4441 1939 4442
rect 1974 4444 1980 4445
rect 112 4418 114 4441
rect 110 4417 116 4418
rect 520 4417 522 4441
rect 744 4417 746 4441
rect 992 4417 994 4441
rect 1264 4417 1266 4441
rect 1552 4417 1554 4441
rect 1816 4417 1818 4441
rect 1936 4418 1938 4441
rect 1974 4440 1975 4444
rect 1979 4440 1980 4444
rect 1994 4441 1995 4445
rect 1999 4441 2000 4445
rect 1994 4440 2000 4441
rect 2130 4445 2136 4446
rect 2130 4441 2131 4445
rect 2135 4441 2136 4445
rect 2130 4440 2136 4441
rect 2266 4445 2272 4446
rect 2266 4441 2267 4445
rect 2271 4441 2272 4445
rect 2266 4440 2272 4441
rect 2402 4445 2408 4446
rect 2402 4441 2403 4445
rect 2407 4441 2408 4445
rect 2402 4440 2408 4441
rect 2538 4445 2544 4446
rect 2538 4441 2539 4445
rect 2543 4441 2544 4445
rect 2538 4440 2544 4441
rect 2674 4445 2680 4446
rect 2674 4441 2675 4445
rect 2679 4441 2680 4445
rect 2674 4440 2680 4441
rect 2810 4445 2816 4446
rect 2810 4441 2811 4445
rect 2815 4441 2816 4445
rect 2810 4440 2816 4441
rect 2946 4445 2952 4446
rect 2946 4441 2947 4445
rect 2951 4441 2952 4445
rect 2946 4440 2952 4441
rect 3798 4444 3804 4445
rect 3798 4440 3799 4444
rect 3803 4440 3804 4444
rect 1974 4439 1980 4440
rect 1934 4417 1940 4418
rect 110 4413 111 4417
rect 115 4413 116 4417
rect 110 4412 116 4413
rect 518 4416 524 4417
rect 518 4412 519 4416
rect 523 4412 524 4416
rect 518 4411 524 4412
rect 742 4416 748 4417
rect 742 4412 743 4416
rect 747 4412 748 4416
rect 742 4411 748 4412
rect 990 4416 996 4417
rect 990 4412 991 4416
rect 995 4412 996 4416
rect 990 4411 996 4412
rect 1262 4416 1268 4417
rect 1262 4412 1263 4416
rect 1267 4412 1268 4416
rect 1262 4411 1268 4412
rect 1550 4416 1556 4417
rect 1550 4412 1551 4416
rect 1555 4412 1556 4416
rect 1550 4411 1556 4412
rect 1814 4416 1820 4417
rect 1814 4412 1815 4416
rect 1819 4412 1820 4416
rect 1934 4413 1935 4417
rect 1939 4413 1940 4417
rect 1934 4412 1940 4413
rect 1814 4411 1820 4412
rect 490 4401 496 4402
rect 110 4400 116 4401
rect 110 4396 111 4400
rect 115 4396 116 4400
rect 490 4397 491 4401
rect 495 4397 496 4401
rect 490 4396 496 4397
rect 714 4401 720 4402
rect 714 4397 715 4401
rect 719 4397 720 4401
rect 714 4396 720 4397
rect 962 4401 968 4402
rect 962 4397 963 4401
rect 967 4397 968 4401
rect 962 4396 968 4397
rect 1234 4401 1240 4402
rect 1234 4397 1235 4401
rect 1239 4397 1240 4401
rect 1234 4396 1240 4397
rect 1522 4401 1528 4402
rect 1522 4397 1523 4401
rect 1527 4397 1528 4401
rect 1522 4396 1528 4397
rect 1786 4401 1792 4402
rect 1786 4397 1787 4401
rect 1791 4397 1792 4401
rect 1786 4396 1792 4397
rect 1934 4400 1940 4401
rect 1934 4396 1935 4400
rect 1939 4396 1940 4400
rect 110 4395 116 4396
rect 112 4335 114 4395
rect 492 4335 494 4396
rect 716 4335 718 4396
rect 964 4335 966 4396
rect 1236 4335 1238 4396
rect 1524 4335 1526 4396
rect 1788 4335 1790 4396
rect 1934 4395 1940 4396
rect 1936 4335 1938 4395
rect 1976 4363 1978 4439
rect 1996 4363 1998 4440
rect 2132 4363 2134 4440
rect 2268 4363 2270 4440
rect 2404 4363 2406 4440
rect 2540 4363 2542 4440
rect 2676 4363 2678 4440
rect 2812 4363 2814 4440
rect 2948 4363 2950 4440
rect 3798 4439 3804 4440
rect 3800 4363 3802 4439
rect 3840 4423 3842 4446
rect 3888 4423 3890 4447
rect 4184 4423 4186 4447
rect 4512 4423 4514 4447
rect 4848 4423 4850 4447
rect 5192 4423 5194 4447
rect 5544 4423 5546 4447
rect 5662 4446 5668 4447
rect 5664 4423 5666 4446
rect 3839 4422 3843 4423
rect 3839 4417 3843 4418
rect 3887 4422 3891 4423
rect 3887 4417 3891 4418
rect 4143 4422 4147 4423
rect 4143 4417 4147 4418
rect 4183 4422 4187 4423
rect 4183 4417 4187 4418
rect 4423 4422 4427 4423
rect 4423 4417 4427 4418
rect 4511 4422 4515 4423
rect 4511 4417 4515 4418
rect 4703 4422 4707 4423
rect 4703 4417 4707 4418
rect 4847 4422 4851 4423
rect 4847 4417 4851 4418
rect 4983 4422 4987 4423
rect 4983 4417 4987 4418
rect 5191 4422 5195 4423
rect 5191 4417 5195 4418
rect 5263 4422 5267 4423
rect 5263 4417 5267 4418
rect 5543 4422 5547 4423
rect 5543 4417 5547 4418
rect 5663 4422 5667 4423
rect 5663 4417 5667 4418
rect 3840 4394 3842 4417
rect 3838 4393 3844 4394
rect 3888 4393 3890 4417
rect 4144 4393 4146 4417
rect 4424 4393 4426 4417
rect 4704 4393 4706 4417
rect 4984 4393 4986 4417
rect 5264 4393 5266 4417
rect 5544 4393 5546 4417
rect 5664 4394 5666 4417
rect 5662 4393 5668 4394
rect 3838 4389 3839 4393
rect 3843 4389 3844 4393
rect 3838 4388 3844 4389
rect 3886 4392 3892 4393
rect 3886 4388 3887 4392
rect 3891 4388 3892 4392
rect 3886 4387 3892 4388
rect 4142 4392 4148 4393
rect 4142 4388 4143 4392
rect 4147 4388 4148 4392
rect 4142 4387 4148 4388
rect 4422 4392 4428 4393
rect 4422 4388 4423 4392
rect 4427 4388 4428 4392
rect 4422 4387 4428 4388
rect 4702 4392 4708 4393
rect 4702 4388 4703 4392
rect 4707 4388 4708 4392
rect 4702 4387 4708 4388
rect 4982 4392 4988 4393
rect 4982 4388 4983 4392
rect 4987 4388 4988 4392
rect 4982 4387 4988 4388
rect 5262 4392 5268 4393
rect 5262 4388 5263 4392
rect 5267 4388 5268 4392
rect 5262 4387 5268 4388
rect 5542 4392 5548 4393
rect 5542 4388 5543 4392
rect 5547 4388 5548 4392
rect 5662 4389 5663 4393
rect 5667 4389 5668 4393
rect 5662 4388 5668 4389
rect 5542 4387 5548 4388
rect 3858 4377 3864 4378
rect 3838 4376 3844 4377
rect 3838 4372 3839 4376
rect 3843 4372 3844 4376
rect 3858 4373 3859 4377
rect 3863 4373 3864 4377
rect 3858 4372 3864 4373
rect 4114 4377 4120 4378
rect 4114 4373 4115 4377
rect 4119 4373 4120 4377
rect 4114 4372 4120 4373
rect 4394 4377 4400 4378
rect 4394 4373 4395 4377
rect 4399 4373 4400 4377
rect 4394 4372 4400 4373
rect 4674 4377 4680 4378
rect 4674 4373 4675 4377
rect 4679 4373 4680 4377
rect 4674 4372 4680 4373
rect 4954 4377 4960 4378
rect 4954 4373 4955 4377
rect 4959 4373 4960 4377
rect 4954 4372 4960 4373
rect 5234 4377 5240 4378
rect 5234 4373 5235 4377
rect 5239 4373 5240 4377
rect 5234 4372 5240 4373
rect 5514 4377 5520 4378
rect 5514 4373 5515 4377
rect 5519 4373 5520 4377
rect 5514 4372 5520 4373
rect 5662 4376 5668 4377
rect 5662 4372 5663 4376
rect 5667 4372 5668 4376
rect 3838 4371 3844 4372
rect 1975 4362 1979 4363
rect 1975 4357 1979 4358
rect 1995 4362 1999 4363
rect 1995 4357 1999 4358
rect 2131 4362 2135 4363
rect 2131 4357 2135 4358
rect 2267 4362 2271 4363
rect 2267 4357 2271 4358
rect 2403 4362 2407 4363
rect 2403 4357 2407 4358
rect 2539 4362 2543 4363
rect 2539 4357 2543 4358
rect 2675 4362 2679 4363
rect 2675 4357 2679 4358
rect 2779 4362 2783 4363
rect 2779 4357 2783 4358
rect 2811 4362 2815 4363
rect 2811 4357 2815 4358
rect 2947 4362 2951 4363
rect 2947 4357 2951 4358
rect 2995 4362 2999 4363
rect 2995 4357 2999 4358
rect 3219 4362 3223 4363
rect 3219 4357 3223 4358
rect 3443 4362 3447 4363
rect 3443 4357 3447 4358
rect 3651 4362 3655 4363
rect 3651 4357 3655 4358
rect 3799 4362 3803 4363
rect 3799 4357 3803 4358
rect 111 4334 115 4335
rect 111 4329 115 4330
rect 491 4334 495 4335
rect 491 4329 495 4330
rect 563 4334 567 4335
rect 563 4329 567 4330
rect 699 4334 703 4335
rect 699 4329 703 4330
rect 715 4334 719 4335
rect 715 4329 719 4330
rect 835 4334 839 4335
rect 835 4329 839 4330
rect 963 4334 967 4335
rect 963 4329 967 4330
rect 971 4334 975 4335
rect 971 4329 975 4330
rect 1107 4334 1111 4335
rect 1107 4329 1111 4330
rect 1235 4334 1239 4335
rect 1235 4329 1239 4330
rect 1243 4334 1247 4335
rect 1243 4329 1247 4330
rect 1379 4334 1383 4335
rect 1379 4329 1383 4330
rect 1515 4334 1519 4335
rect 1515 4329 1519 4330
rect 1523 4334 1527 4335
rect 1523 4329 1527 4330
rect 1651 4334 1655 4335
rect 1651 4329 1655 4330
rect 1787 4334 1791 4335
rect 1787 4329 1791 4330
rect 1935 4334 1939 4335
rect 1935 4329 1939 4330
rect 112 4269 114 4329
rect 110 4268 116 4269
rect 564 4268 566 4329
rect 700 4268 702 4329
rect 836 4268 838 4329
rect 972 4268 974 4329
rect 1108 4268 1110 4329
rect 1244 4268 1246 4329
rect 1380 4268 1382 4329
rect 1516 4268 1518 4329
rect 1652 4268 1654 4329
rect 1788 4268 1790 4329
rect 1936 4269 1938 4329
rect 1976 4297 1978 4357
rect 1974 4296 1980 4297
rect 2780 4296 2782 4357
rect 2996 4296 2998 4357
rect 3220 4296 3222 4357
rect 3444 4296 3446 4357
rect 3652 4296 3654 4357
rect 3800 4297 3802 4357
rect 3840 4299 3842 4371
rect 3860 4299 3862 4372
rect 4116 4299 4118 4372
rect 4396 4299 4398 4372
rect 4676 4299 4678 4372
rect 4956 4299 4958 4372
rect 5236 4299 5238 4372
rect 5516 4299 5518 4372
rect 5662 4371 5668 4372
rect 5664 4299 5666 4371
rect 3839 4298 3843 4299
rect 3798 4296 3804 4297
rect 1974 4292 1975 4296
rect 1979 4292 1980 4296
rect 1974 4291 1980 4292
rect 2778 4295 2784 4296
rect 2778 4291 2779 4295
rect 2783 4291 2784 4295
rect 2778 4290 2784 4291
rect 2994 4295 3000 4296
rect 2994 4291 2995 4295
rect 2999 4291 3000 4295
rect 2994 4290 3000 4291
rect 3218 4295 3224 4296
rect 3218 4291 3219 4295
rect 3223 4291 3224 4295
rect 3218 4290 3224 4291
rect 3442 4295 3448 4296
rect 3442 4291 3443 4295
rect 3447 4291 3448 4295
rect 3442 4290 3448 4291
rect 3650 4295 3656 4296
rect 3650 4291 3651 4295
rect 3655 4291 3656 4295
rect 3798 4292 3799 4296
rect 3803 4292 3804 4296
rect 3839 4293 3843 4294
rect 3859 4298 3863 4299
rect 3859 4293 3863 4294
rect 4115 4298 4119 4299
rect 4115 4293 4119 4294
rect 4395 4298 4399 4299
rect 4395 4293 4399 4294
rect 4571 4298 4575 4299
rect 4571 4293 4575 4294
rect 4675 4298 4679 4299
rect 4675 4293 4679 4294
rect 4739 4298 4743 4299
rect 4739 4293 4743 4294
rect 4915 4298 4919 4299
rect 4915 4293 4919 4294
rect 4955 4298 4959 4299
rect 4955 4293 4959 4294
rect 5107 4298 5111 4299
rect 5107 4293 5111 4294
rect 5235 4298 5239 4299
rect 5235 4293 5239 4294
rect 5307 4298 5311 4299
rect 5307 4293 5311 4294
rect 5515 4298 5519 4299
rect 5515 4293 5519 4294
rect 5663 4298 5667 4299
rect 5663 4293 5667 4294
rect 3798 4291 3804 4292
rect 3650 4290 3656 4291
rect 2806 4280 2812 4281
rect 1974 4279 1980 4280
rect 1974 4275 1975 4279
rect 1979 4275 1980 4279
rect 2806 4276 2807 4280
rect 2811 4276 2812 4280
rect 2806 4275 2812 4276
rect 3022 4280 3028 4281
rect 3022 4276 3023 4280
rect 3027 4276 3028 4280
rect 3022 4275 3028 4276
rect 3246 4280 3252 4281
rect 3246 4276 3247 4280
rect 3251 4276 3252 4280
rect 3246 4275 3252 4276
rect 3470 4280 3476 4281
rect 3470 4276 3471 4280
rect 3475 4276 3476 4280
rect 3470 4275 3476 4276
rect 3678 4280 3684 4281
rect 3678 4276 3679 4280
rect 3683 4276 3684 4280
rect 3678 4275 3684 4276
rect 3798 4279 3804 4280
rect 3798 4275 3799 4279
rect 3803 4275 3804 4279
rect 1974 4274 1980 4275
rect 1934 4268 1940 4269
rect 110 4264 111 4268
rect 115 4264 116 4268
rect 110 4263 116 4264
rect 562 4267 568 4268
rect 562 4263 563 4267
rect 567 4263 568 4267
rect 562 4262 568 4263
rect 698 4267 704 4268
rect 698 4263 699 4267
rect 703 4263 704 4267
rect 698 4262 704 4263
rect 834 4267 840 4268
rect 834 4263 835 4267
rect 839 4263 840 4267
rect 834 4262 840 4263
rect 970 4267 976 4268
rect 970 4263 971 4267
rect 975 4263 976 4267
rect 970 4262 976 4263
rect 1106 4267 1112 4268
rect 1106 4263 1107 4267
rect 1111 4263 1112 4267
rect 1106 4262 1112 4263
rect 1242 4267 1248 4268
rect 1242 4263 1243 4267
rect 1247 4263 1248 4267
rect 1242 4262 1248 4263
rect 1378 4267 1384 4268
rect 1378 4263 1379 4267
rect 1383 4263 1384 4267
rect 1378 4262 1384 4263
rect 1514 4267 1520 4268
rect 1514 4263 1515 4267
rect 1519 4263 1520 4267
rect 1514 4262 1520 4263
rect 1650 4267 1656 4268
rect 1650 4263 1651 4267
rect 1655 4263 1656 4267
rect 1650 4262 1656 4263
rect 1786 4267 1792 4268
rect 1786 4263 1787 4267
rect 1791 4263 1792 4267
rect 1934 4264 1935 4268
rect 1939 4264 1940 4268
rect 1934 4263 1940 4264
rect 1786 4262 1792 4263
rect 590 4252 596 4253
rect 110 4251 116 4252
rect 110 4247 111 4251
rect 115 4247 116 4251
rect 590 4248 591 4252
rect 595 4248 596 4252
rect 590 4247 596 4248
rect 726 4252 732 4253
rect 726 4248 727 4252
rect 731 4248 732 4252
rect 726 4247 732 4248
rect 862 4252 868 4253
rect 862 4248 863 4252
rect 867 4248 868 4252
rect 862 4247 868 4248
rect 998 4252 1004 4253
rect 998 4248 999 4252
rect 1003 4248 1004 4252
rect 998 4247 1004 4248
rect 1134 4252 1140 4253
rect 1134 4248 1135 4252
rect 1139 4248 1140 4252
rect 1134 4247 1140 4248
rect 1270 4252 1276 4253
rect 1270 4248 1271 4252
rect 1275 4248 1276 4252
rect 1270 4247 1276 4248
rect 1406 4252 1412 4253
rect 1406 4248 1407 4252
rect 1411 4248 1412 4252
rect 1406 4247 1412 4248
rect 1542 4252 1548 4253
rect 1542 4248 1543 4252
rect 1547 4248 1548 4252
rect 1542 4247 1548 4248
rect 1678 4252 1684 4253
rect 1678 4248 1679 4252
rect 1683 4248 1684 4252
rect 1678 4247 1684 4248
rect 1814 4252 1820 4253
rect 1814 4248 1815 4252
rect 1819 4248 1820 4252
rect 1814 4247 1820 4248
rect 1934 4251 1940 4252
rect 1934 4247 1935 4251
rect 1939 4247 1940 4251
rect 110 4246 116 4247
rect 112 4211 114 4246
rect 592 4211 594 4247
rect 728 4211 730 4247
rect 864 4211 866 4247
rect 1000 4211 1002 4247
rect 1136 4211 1138 4247
rect 1272 4211 1274 4247
rect 1408 4211 1410 4247
rect 1544 4211 1546 4247
rect 1680 4211 1682 4247
rect 1816 4211 1818 4247
rect 1934 4246 1940 4247
rect 1936 4211 1938 4246
rect 1976 4223 1978 4274
rect 2808 4223 2810 4275
rect 3024 4223 3026 4275
rect 3248 4223 3250 4275
rect 3472 4223 3474 4275
rect 3680 4223 3682 4275
rect 3798 4274 3804 4275
rect 3800 4223 3802 4274
rect 3840 4233 3842 4293
rect 3838 4232 3844 4233
rect 4572 4232 4574 4293
rect 4740 4232 4742 4293
rect 4916 4232 4918 4293
rect 5108 4232 5110 4293
rect 5308 4232 5310 4293
rect 5516 4232 5518 4293
rect 5664 4233 5666 4293
rect 5662 4232 5668 4233
rect 3838 4228 3839 4232
rect 3843 4228 3844 4232
rect 3838 4227 3844 4228
rect 4570 4231 4576 4232
rect 4570 4227 4571 4231
rect 4575 4227 4576 4231
rect 4570 4226 4576 4227
rect 4738 4231 4744 4232
rect 4738 4227 4739 4231
rect 4743 4227 4744 4231
rect 4738 4226 4744 4227
rect 4914 4231 4920 4232
rect 4914 4227 4915 4231
rect 4919 4227 4920 4231
rect 4914 4226 4920 4227
rect 5106 4231 5112 4232
rect 5106 4227 5107 4231
rect 5111 4227 5112 4231
rect 5106 4226 5112 4227
rect 5306 4231 5312 4232
rect 5306 4227 5307 4231
rect 5311 4227 5312 4231
rect 5306 4226 5312 4227
rect 5514 4231 5520 4232
rect 5514 4227 5515 4231
rect 5519 4227 5520 4231
rect 5662 4228 5663 4232
rect 5667 4228 5668 4232
rect 5662 4227 5668 4228
rect 5514 4226 5520 4227
rect 1975 4222 1979 4223
rect 1975 4217 1979 4218
rect 2807 4222 2811 4223
rect 2807 4217 2811 4218
rect 2951 4222 2955 4223
rect 2951 4217 2955 4218
rect 3023 4222 3027 4223
rect 3023 4217 3027 4218
rect 3095 4222 3099 4223
rect 3095 4217 3099 4218
rect 3239 4222 3243 4223
rect 3239 4217 3243 4218
rect 3247 4222 3251 4223
rect 3247 4217 3251 4218
rect 3391 4222 3395 4223
rect 3391 4217 3395 4218
rect 3471 4222 3475 4223
rect 3471 4217 3475 4218
rect 3543 4222 3547 4223
rect 3543 4217 3547 4218
rect 3679 4222 3683 4223
rect 3679 4217 3683 4218
rect 3799 4222 3803 4223
rect 3799 4217 3803 4218
rect 111 4210 115 4211
rect 111 4205 115 4206
rect 591 4210 595 4211
rect 591 4205 595 4206
rect 727 4210 731 4211
rect 727 4205 731 4206
rect 863 4210 867 4211
rect 863 4205 867 4206
rect 999 4210 1003 4211
rect 999 4205 1003 4206
rect 1135 4210 1139 4211
rect 1135 4205 1139 4206
rect 1271 4210 1275 4211
rect 1271 4205 1275 4206
rect 1407 4210 1411 4211
rect 1407 4205 1411 4206
rect 1543 4210 1547 4211
rect 1543 4205 1547 4206
rect 1679 4210 1683 4211
rect 1679 4205 1683 4206
rect 1815 4210 1819 4211
rect 1815 4205 1819 4206
rect 1935 4210 1939 4211
rect 1935 4205 1939 4206
rect 112 4182 114 4205
rect 110 4181 116 4182
rect 592 4181 594 4205
rect 728 4181 730 4205
rect 864 4181 866 4205
rect 1000 4181 1002 4205
rect 1136 4181 1138 4205
rect 1272 4181 1274 4205
rect 1408 4181 1410 4205
rect 1544 4181 1546 4205
rect 1680 4181 1682 4205
rect 1816 4181 1818 4205
rect 1936 4182 1938 4205
rect 1976 4194 1978 4217
rect 1974 4193 1980 4194
rect 2952 4193 2954 4217
rect 3096 4193 3098 4217
rect 3240 4193 3242 4217
rect 3392 4193 3394 4217
rect 3544 4193 3546 4217
rect 3680 4193 3682 4217
rect 3800 4194 3802 4217
rect 4598 4216 4604 4217
rect 3838 4215 3844 4216
rect 3838 4211 3839 4215
rect 3843 4211 3844 4215
rect 4598 4212 4599 4216
rect 4603 4212 4604 4216
rect 4598 4211 4604 4212
rect 4766 4216 4772 4217
rect 4766 4212 4767 4216
rect 4771 4212 4772 4216
rect 4766 4211 4772 4212
rect 4942 4216 4948 4217
rect 4942 4212 4943 4216
rect 4947 4212 4948 4216
rect 4942 4211 4948 4212
rect 5134 4216 5140 4217
rect 5134 4212 5135 4216
rect 5139 4212 5140 4216
rect 5134 4211 5140 4212
rect 5334 4216 5340 4217
rect 5334 4212 5335 4216
rect 5339 4212 5340 4216
rect 5334 4211 5340 4212
rect 5542 4216 5548 4217
rect 5542 4212 5543 4216
rect 5547 4212 5548 4216
rect 5542 4211 5548 4212
rect 5662 4215 5668 4216
rect 5662 4211 5663 4215
rect 5667 4211 5668 4215
rect 3838 4210 3844 4211
rect 3798 4193 3804 4194
rect 1974 4189 1975 4193
rect 1979 4189 1980 4193
rect 1974 4188 1980 4189
rect 2950 4192 2956 4193
rect 2950 4188 2951 4192
rect 2955 4188 2956 4192
rect 2950 4187 2956 4188
rect 3094 4192 3100 4193
rect 3094 4188 3095 4192
rect 3099 4188 3100 4192
rect 3094 4187 3100 4188
rect 3238 4192 3244 4193
rect 3238 4188 3239 4192
rect 3243 4188 3244 4192
rect 3238 4187 3244 4188
rect 3390 4192 3396 4193
rect 3390 4188 3391 4192
rect 3395 4188 3396 4192
rect 3390 4187 3396 4188
rect 3542 4192 3548 4193
rect 3542 4188 3543 4192
rect 3547 4188 3548 4192
rect 3542 4187 3548 4188
rect 3678 4192 3684 4193
rect 3678 4188 3679 4192
rect 3683 4188 3684 4192
rect 3798 4189 3799 4193
rect 3803 4189 3804 4193
rect 3798 4188 3804 4189
rect 3678 4187 3684 4188
rect 3840 4187 3842 4210
rect 4600 4187 4602 4211
rect 4768 4187 4770 4211
rect 4944 4187 4946 4211
rect 5136 4187 5138 4211
rect 5336 4187 5338 4211
rect 5544 4187 5546 4211
rect 5662 4210 5668 4211
rect 5664 4187 5666 4210
rect 3839 4186 3843 4187
rect 1934 4181 1940 4182
rect 3839 4181 3843 4182
rect 4599 4186 4603 4187
rect 4599 4181 4603 4182
rect 4655 4186 4659 4187
rect 4655 4181 4659 4182
rect 4767 4186 4771 4187
rect 4767 4181 4771 4182
rect 4815 4186 4819 4187
rect 4815 4181 4819 4182
rect 4943 4186 4947 4187
rect 4943 4181 4947 4182
rect 4983 4186 4987 4187
rect 4983 4181 4987 4182
rect 5135 4186 5139 4187
rect 5135 4181 5139 4182
rect 5167 4186 5171 4187
rect 5167 4181 5171 4182
rect 5335 4186 5339 4187
rect 5335 4181 5339 4182
rect 5359 4186 5363 4187
rect 5359 4181 5363 4182
rect 5543 4186 5547 4187
rect 5543 4181 5547 4182
rect 5663 4186 5667 4187
rect 5663 4181 5667 4182
rect 110 4177 111 4181
rect 115 4177 116 4181
rect 110 4176 116 4177
rect 590 4180 596 4181
rect 590 4176 591 4180
rect 595 4176 596 4180
rect 590 4175 596 4176
rect 726 4180 732 4181
rect 726 4176 727 4180
rect 731 4176 732 4180
rect 726 4175 732 4176
rect 862 4180 868 4181
rect 862 4176 863 4180
rect 867 4176 868 4180
rect 862 4175 868 4176
rect 998 4180 1004 4181
rect 998 4176 999 4180
rect 1003 4176 1004 4180
rect 998 4175 1004 4176
rect 1134 4180 1140 4181
rect 1134 4176 1135 4180
rect 1139 4176 1140 4180
rect 1134 4175 1140 4176
rect 1270 4180 1276 4181
rect 1270 4176 1271 4180
rect 1275 4176 1276 4180
rect 1270 4175 1276 4176
rect 1406 4180 1412 4181
rect 1406 4176 1407 4180
rect 1411 4176 1412 4180
rect 1406 4175 1412 4176
rect 1542 4180 1548 4181
rect 1542 4176 1543 4180
rect 1547 4176 1548 4180
rect 1542 4175 1548 4176
rect 1678 4180 1684 4181
rect 1678 4176 1679 4180
rect 1683 4176 1684 4180
rect 1678 4175 1684 4176
rect 1814 4180 1820 4181
rect 1814 4176 1815 4180
rect 1819 4176 1820 4180
rect 1934 4177 1935 4181
rect 1939 4177 1940 4181
rect 2922 4177 2928 4178
rect 1934 4176 1940 4177
rect 1974 4176 1980 4177
rect 1814 4175 1820 4176
rect 1974 4172 1975 4176
rect 1979 4172 1980 4176
rect 2922 4173 2923 4177
rect 2927 4173 2928 4177
rect 2922 4172 2928 4173
rect 3066 4177 3072 4178
rect 3066 4173 3067 4177
rect 3071 4173 3072 4177
rect 3066 4172 3072 4173
rect 3210 4177 3216 4178
rect 3210 4173 3211 4177
rect 3215 4173 3216 4177
rect 3210 4172 3216 4173
rect 3362 4177 3368 4178
rect 3362 4173 3363 4177
rect 3367 4173 3368 4177
rect 3362 4172 3368 4173
rect 3514 4177 3520 4178
rect 3514 4173 3515 4177
rect 3519 4173 3520 4177
rect 3514 4172 3520 4173
rect 3650 4177 3656 4178
rect 3650 4173 3651 4177
rect 3655 4173 3656 4177
rect 3650 4172 3656 4173
rect 3798 4176 3804 4177
rect 3798 4172 3799 4176
rect 3803 4172 3804 4176
rect 1974 4171 1980 4172
rect 562 4165 568 4166
rect 110 4164 116 4165
rect 110 4160 111 4164
rect 115 4160 116 4164
rect 562 4161 563 4165
rect 567 4161 568 4165
rect 562 4160 568 4161
rect 698 4165 704 4166
rect 698 4161 699 4165
rect 703 4161 704 4165
rect 698 4160 704 4161
rect 834 4165 840 4166
rect 834 4161 835 4165
rect 839 4161 840 4165
rect 834 4160 840 4161
rect 970 4165 976 4166
rect 970 4161 971 4165
rect 975 4161 976 4165
rect 970 4160 976 4161
rect 1106 4165 1112 4166
rect 1106 4161 1107 4165
rect 1111 4161 1112 4165
rect 1106 4160 1112 4161
rect 1242 4165 1248 4166
rect 1242 4161 1243 4165
rect 1247 4161 1248 4165
rect 1242 4160 1248 4161
rect 1378 4165 1384 4166
rect 1378 4161 1379 4165
rect 1383 4161 1384 4165
rect 1378 4160 1384 4161
rect 1514 4165 1520 4166
rect 1514 4161 1515 4165
rect 1519 4161 1520 4165
rect 1514 4160 1520 4161
rect 1650 4165 1656 4166
rect 1650 4161 1651 4165
rect 1655 4161 1656 4165
rect 1650 4160 1656 4161
rect 1786 4165 1792 4166
rect 1786 4161 1787 4165
rect 1791 4161 1792 4165
rect 1786 4160 1792 4161
rect 1934 4164 1940 4165
rect 1934 4160 1935 4164
rect 1939 4160 1940 4164
rect 110 4159 116 4160
rect 112 4099 114 4159
rect 564 4099 566 4160
rect 700 4099 702 4160
rect 836 4099 838 4160
rect 972 4099 974 4160
rect 1108 4099 1110 4160
rect 1244 4099 1246 4160
rect 1380 4099 1382 4160
rect 1516 4099 1518 4160
rect 1652 4099 1654 4160
rect 1788 4099 1790 4160
rect 1934 4159 1940 4160
rect 1936 4099 1938 4159
rect 111 4098 115 4099
rect 111 4093 115 4094
rect 563 4098 567 4099
rect 563 4093 567 4094
rect 699 4098 703 4099
rect 699 4093 703 4094
rect 835 4098 839 4099
rect 835 4093 839 4094
rect 971 4098 975 4099
rect 971 4093 975 4094
rect 1107 4098 1111 4099
rect 1107 4093 1111 4094
rect 1243 4098 1247 4099
rect 1243 4093 1247 4094
rect 1379 4098 1383 4099
rect 1379 4093 1383 4094
rect 1515 4098 1519 4099
rect 1515 4093 1519 4094
rect 1651 4098 1655 4099
rect 1651 4093 1655 4094
rect 1787 4098 1791 4099
rect 1787 4093 1791 4094
rect 1935 4098 1939 4099
rect 1935 4093 1939 4094
rect 112 4033 114 4093
rect 110 4032 116 4033
rect 700 4032 702 4093
rect 836 4032 838 4093
rect 972 4032 974 4093
rect 1108 4032 1110 4093
rect 1244 4032 1246 4093
rect 1380 4032 1382 4093
rect 1516 4032 1518 4093
rect 1652 4032 1654 4093
rect 1788 4032 1790 4093
rect 1936 4033 1938 4093
rect 1976 4075 1978 4171
rect 2924 4075 2926 4172
rect 3068 4075 3070 4172
rect 3212 4075 3214 4172
rect 3364 4075 3366 4172
rect 3516 4075 3518 4172
rect 3652 4075 3654 4172
rect 3798 4171 3804 4172
rect 3800 4075 3802 4171
rect 3840 4158 3842 4181
rect 3838 4157 3844 4158
rect 4656 4157 4658 4181
rect 4816 4157 4818 4181
rect 4984 4157 4986 4181
rect 5168 4157 5170 4181
rect 5360 4157 5362 4181
rect 5544 4157 5546 4181
rect 5664 4158 5666 4181
rect 5662 4157 5668 4158
rect 3838 4153 3839 4157
rect 3843 4153 3844 4157
rect 3838 4152 3844 4153
rect 4654 4156 4660 4157
rect 4654 4152 4655 4156
rect 4659 4152 4660 4156
rect 4654 4151 4660 4152
rect 4814 4156 4820 4157
rect 4814 4152 4815 4156
rect 4819 4152 4820 4156
rect 4814 4151 4820 4152
rect 4982 4156 4988 4157
rect 4982 4152 4983 4156
rect 4987 4152 4988 4156
rect 4982 4151 4988 4152
rect 5166 4156 5172 4157
rect 5166 4152 5167 4156
rect 5171 4152 5172 4156
rect 5166 4151 5172 4152
rect 5358 4156 5364 4157
rect 5358 4152 5359 4156
rect 5363 4152 5364 4156
rect 5358 4151 5364 4152
rect 5542 4156 5548 4157
rect 5542 4152 5543 4156
rect 5547 4152 5548 4156
rect 5662 4153 5663 4157
rect 5667 4153 5668 4157
rect 5662 4152 5668 4153
rect 5542 4151 5548 4152
rect 4626 4141 4632 4142
rect 3838 4140 3844 4141
rect 3838 4136 3839 4140
rect 3843 4136 3844 4140
rect 4626 4137 4627 4141
rect 4631 4137 4632 4141
rect 4626 4136 4632 4137
rect 4786 4141 4792 4142
rect 4786 4137 4787 4141
rect 4791 4137 4792 4141
rect 4786 4136 4792 4137
rect 4954 4141 4960 4142
rect 4954 4137 4955 4141
rect 4959 4137 4960 4141
rect 4954 4136 4960 4137
rect 5138 4141 5144 4142
rect 5138 4137 5139 4141
rect 5143 4137 5144 4141
rect 5138 4136 5144 4137
rect 5330 4141 5336 4142
rect 5330 4137 5331 4141
rect 5335 4137 5336 4141
rect 5330 4136 5336 4137
rect 5514 4141 5520 4142
rect 5514 4137 5515 4141
rect 5519 4137 5520 4141
rect 5514 4136 5520 4137
rect 5662 4140 5668 4141
rect 5662 4136 5663 4140
rect 5667 4136 5668 4140
rect 3838 4135 3844 4136
rect 1975 4074 1979 4075
rect 1975 4069 1979 4070
rect 2899 4074 2903 4075
rect 2899 4069 2903 4070
rect 2923 4074 2927 4075
rect 2923 4069 2927 4070
rect 3043 4074 3047 4075
rect 3043 4069 3047 4070
rect 3067 4074 3071 4075
rect 3067 4069 3071 4070
rect 3187 4074 3191 4075
rect 3187 4069 3191 4070
rect 3211 4074 3215 4075
rect 3211 4069 3215 4070
rect 3339 4074 3343 4075
rect 3339 4069 3343 4070
rect 3363 4074 3367 4075
rect 3363 4069 3367 4070
rect 3491 4074 3495 4075
rect 3491 4069 3495 4070
rect 3515 4074 3519 4075
rect 3515 4069 3519 4070
rect 3643 4074 3647 4075
rect 3643 4069 3647 4070
rect 3651 4074 3655 4075
rect 3651 4069 3655 4070
rect 3799 4074 3803 4075
rect 3799 4069 3803 4070
rect 1934 4032 1940 4033
rect 110 4028 111 4032
rect 115 4028 116 4032
rect 110 4027 116 4028
rect 698 4031 704 4032
rect 698 4027 699 4031
rect 703 4027 704 4031
rect 698 4026 704 4027
rect 834 4031 840 4032
rect 834 4027 835 4031
rect 839 4027 840 4031
rect 834 4026 840 4027
rect 970 4031 976 4032
rect 970 4027 971 4031
rect 975 4027 976 4031
rect 970 4026 976 4027
rect 1106 4031 1112 4032
rect 1106 4027 1107 4031
rect 1111 4027 1112 4031
rect 1106 4026 1112 4027
rect 1242 4031 1248 4032
rect 1242 4027 1243 4031
rect 1247 4027 1248 4031
rect 1242 4026 1248 4027
rect 1378 4031 1384 4032
rect 1378 4027 1379 4031
rect 1383 4027 1384 4031
rect 1378 4026 1384 4027
rect 1514 4031 1520 4032
rect 1514 4027 1515 4031
rect 1519 4027 1520 4031
rect 1514 4026 1520 4027
rect 1650 4031 1656 4032
rect 1650 4027 1651 4031
rect 1655 4027 1656 4031
rect 1650 4026 1656 4027
rect 1786 4031 1792 4032
rect 1786 4027 1787 4031
rect 1791 4027 1792 4031
rect 1934 4028 1935 4032
rect 1939 4028 1940 4032
rect 1934 4027 1940 4028
rect 1786 4026 1792 4027
rect 726 4016 732 4017
rect 110 4015 116 4016
rect 110 4011 111 4015
rect 115 4011 116 4015
rect 726 4012 727 4016
rect 731 4012 732 4016
rect 726 4011 732 4012
rect 862 4016 868 4017
rect 862 4012 863 4016
rect 867 4012 868 4016
rect 862 4011 868 4012
rect 998 4016 1004 4017
rect 998 4012 999 4016
rect 1003 4012 1004 4016
rect 998 4011 1004 4012
rect 1134 4016 1140 4017
rect 1134 4012 1135 4016
rect 1139 4012 1140 4016
rect 1134 4011 1140 4012
rect 1270 4016 1276 4017
rect 1270 4012 1271 4016
rect 1275 4012 1276 4016
rect 1270 4011 1276 4012
rect 1406 4016 1412 4017
rect 1406 4012 1407 4016
rect 1411 4012 1412 4016
rect 1406 4011 1412 4012
rect 1542 4016 1548 4017
rect 1542 4012 1543 4016
rect 1547 4012 1548 4016
rect 1542 4011 1548 4012
rect 1678 4016 1684 4017
rect 1678 4012 1679 4016
rect 1683 4012 1684 4016
rect 1678 4011 1684 4012
rect 1814 4016 1820 4017
rect 1814 4012 1815 4016
rect 1819 4012 1820 4016
rect 1814 4011 1820 4012
rect 1934 4015 1940 4016
rect 1934 4011 1935 4015
rect 1939 4011 1940 4015
rect 110 4010 116 4011
rect 112 3983 114 4010
rect 728 3983 730 4011
rect 864 3983 866 4011
rect 1000 3983 1002 4011
rect 1136 3983 1138 4011
rect 1272 3983 1274 4011
rect 1408 3983 1410 4011
rect 1544 3983 1546 4011
rect 1680 3983 1682 4011
rect 1816 3983 1818 4011
rect 1934 4010 1940 4011
rect 1936 3983 1938 4010
rect 1976 4009 1978 4069
rect 1974 4008 1980 4009
rect 2900 4008 2902 4069
rect 3044 4008 3046 4069
rect 3188 4008 3190 4069
rect 3340 4008 3342 4069
rect 3492 4008 3494 4069
rect 3644 4008 3646 4069
rect 3800 4009 3802 4069
rect 3840 4039 3842 4135
rect 4628 4039 4630 4136
rect 4788 4039 4790 4136
rect 4956 4039 4958 4136
rect 5140 4039 5142 4136
rect 5332 4039 5334 4136
rect 5516 4039 5518 4136
rect 5662 4135 5668 4136
rect 5664 4039 5666 4135
rect 3839 4038 3843 4039
rect 3839 4033 3843 4034
rect 4627 4038 4631 4039
rect 4627 4033 4631 4034
rect 4787 4038 4791 4039
rect 4787 4033 4791 4034
rect 4939 4038 4943 4039
rect 4939 4033 4943 4034
rect 4955 4038 4959 4039
rect 4955 4033 4959 4034
rect 5075 4038 5079 4039
rect 5075 4033 5079 4034
rect 5139 4038 5143 4039
rect 5139 4033 5143 4034
rect 5211 4038 5215 4039
rect 5211 4033 5215 4034
rect 5331 4038 5335 4039
rect 5331 4033 5335 4034
rect 5347 4038 5351 4039
rect 5347 4033 5351 4034
rect 5515 4038 5519 4039
rect 5515 4033 5519 4034
rect 5663 4038 5667 4039
rect 5663 4033 5667 4034
rect 3798 4008 3804 4009
rect 1974 4004 1975 4008
rect 1979 4004 1980 4008
rect 1974 4003 1980 4004
rect 2898 4007 2904 4008
rect 2898 4003 2899 4007
rect 2903 4003 2904 4007
rect 2898 4002 2904 4003
rect 3042 4007 3048 4008
rect 3042 4003 3043 4007
rect 3047 4003 3048 4007
rect 3042 4002 3048 4003
rect 3186 4007 3192 4008
rect 3186 4003 3187 4007
rect 3191 4003 3192 4007
rect 3186 4002 3192 4003
rect 3338 4007 3344 4008
rect 3338 4003 3339 4007
rect 3343 4003 3344 4007
rect 3338 4002 3344 4003
rect 3490 4007 3496 4008
rect 3490 4003 3491 4007
rect 3495 4003 3496 4007
rect 3490 4002 3496 4003
rect 3642 4007 3648 4008
rect 3642 4003 3643 4007
rect 3647 4003 3648 4007
rect 3798 4004 3799 4008
rect 3803 4004 3804 4008
rect 3798 4003 3804 4004
rect 3642 4002 3648 4003
rect 2926 3992 2932 3993
rect 1974 3991 1980 3992
rect 1974 3987 1975 3991
rect 1979 3987 1980 3991
rect 2926 3988 2927 3992
rect 2931 3988 2932 3992
rect 2926 3987 2932 3988
rect 3070 3992 3076 3993
rect 3070 3988 3071 3992
rect 3075 3988 3076 3992
rect 3070 3987 3076 3988
rect 3214 3992 3220 3993
rect 3214 3988 3215 3992
rect 3219 3988 3220 3992
rect 3214 3987 3220 3988
rect 3366 3992 3372 3993
rect 3366 3988 3367 3992
rect 3371 3988 3372 3992
rect 3366 3987 3372 3988
rect 3518 3992 3524 3993
rect 3518 3988 3519 3992
rect 3523 3988 3524 3992
rect 3518 3987 3524 3988
rect 3670 3992 3676 3993
rect 3670 3988 3671 3992
rect 3675 3988 3676 3992
rect 3670 3987 3676 3988
rect 3798 3991 3804 3992
rect 3798 3987 3799 3991
rect 3803 3987 3804 3991
rect 1974 3986 1980 3987
rect 111 3982 115 3983
rect 111 3977 115 3978
rect 695 3982 699 3983
rect 695 3977 699 3978
rect 727 3982 731 3983
rect 727 3977 731 3978
rect 831 3982 835 3983
rect 831 3977 835 3978
rect 863 3982 867 3983
rect 863 3977 867 3978
rect 967 3982 971 3983
rect 967 3977 971 3978
rect 999 3982 1003 3983
rect 999 3977 1003 3978
rect 1111 3982 1115 3983
rect 1111 3977 1115 3978
rect 1135 3982 1139 3983
rect 1135 3977 1139 3978
rect 1255 3982 1259 3983
rect 1255 3977 1259 3978
rect 1271 3982 1275 3983
rect 1271 3977 1275 3978
rect 1399 3982 1403 3983
rect 1399 3977 1403 3978
rect 1407 3982 1411 3983
rect 1407 3977 1411 3978
rect 1543 3982 1547 3983
rect 1543 3977 1547 3978
rect 1679 3982 1683 3983
rect 1679 3977 1683 3978
rect 1815 3982 1819 3983
rect 1815 3977 1819 3978
rect 1935 3982 1939 3983
rect 1935 3977 1939 3978
rect 112 3954 114 3977
rect 110 3953 116 3954
rect 696 3953 698 3977
rect 832 3953 834 3977
rect 968 3953 970 3977
rect 1112 3953 1114 3977
rect 1256 3953 1258 3977
rect 1400 3953 1402 3977
rect 1544 3953 1546 3977
rect 1680 3953 1682 3977
rect 1816 3953 1818 3977
rect 1936 3954 1938 3977
rect 1934 3953 1940 3954
rect 110 3949 111 3953
rect 115 3949 116 3953
rect 110 3948 116 3949
rect 694 3952 700 3953
rect 694 3948 695 3952
rect 699 3948 700 3952
rect 694 3947 700 3948
rect 830 3952 836 3953
rect 830 3948 831 3952
rect 835 3948 836 3952
rect 830 3947 836 3948
rect 966 3952 972 3953
rect 966 3948 967 3952
rect 971 3948 972 3952
rect 966 3947 972 3948
rect 1110 3952 1116 3953
rect 1110 3948 1111 3952
rect 1115 3948 1116 3952
rect 1110 3947 1116 3948
rect 1254 3952 1260 3953
rect 1254 3948 1255 3952
rect 1259 3948 1260 3952
rect 1254 3947 1260 3948
rect 1398 3952 1404 3953
rect 1398 3948 1399 3952
rect 1403 3948 1404 3952
rect 1398 3947 1404 3948
rect 1542 3952 1548 3953
rect 1542 3948 1543 3952
rect 1547 3948 1548 3952
rect 1542 3947 1548 3948
rect 1678 3952 1684 3953
rect 1678 3948 1679 3952
rect 1683 3948 1684 3952
rect 1678 3947 1684 3948
rect 1814 3952 1820 3953
rect 1814 3948 1815 3952
rect 1819 3948 1820 3952
rect 1934 3949 1935 3953
rect 1939 3949 1940 3953
rect 1934 3948 1940 3949
rect 1814 3947 1820 3948
rect 666 3937 672 3938
rect 110 3936 116 3937
rect 110 3932 111 3936
rect 115 3932 116 3936
rect 666 3933 667 3937
rect 671 3933 672 3937
rect 666 3932 672 3933
rect 802 3937 808 3938
rect 802 3933 803 3937
rect 807 3933 808 3937
rect 802 3932 808 3933
rect 938 3937 944 3938
rect 938 3933 939 3937
rect 943 3933 944 3937
rect 938 3932 944 3933
rect 1082 3937 1088 3938
rect 1082 3933 1083 3937
rect 1087 3933 1088 3937
rect 1082 3932 1088 3933
rect 1226 3937 1232 3938
rect 1226 3933 1227 3937
rect 1231 3933 1232 3937
rect 1226 3932 1232 3933
rect 1370 3937 1376 3938
rect 1370 3933 1371 3937
rect 1375 3933 1376 3937
rect 1370 3932 1376 3933
rect 1514 3937 1520 3938
rect 1514 3933 1515 3937
rect 1519 3933 1520 3937
rect 1514 3932 1520 3933
rect 1650 3937 1656 3938
rect 1650 3933 1651 3937
rect 1655 3933 1656 3937
rect 1650 3932 1656 3933
rect 1786 3937 1792 3938
rect 1786 3933 1787 3937
rect 1791 3933 1792 3937
rect 1786 3932 1792 3933
rect 1934 3936 1940 3937
rect 1934 3932 1935 3936
rect 1939 3932 1940 3936
rect 1976 3935 1978 3986
rect 2928 3935 2930 3987
rect 3072 3935 3074 3987
rect 3216 3935 3218 3987
rect 3368 3935 3370 3987
rect 3520 3935 3522 3987
rect 3672 3935 3674 3987
rect 3798 3986 3804 3987
rect 3800 3935 3802 3986
rect 3840 3973 3842 4033
rect 3838 3972 3844 3973
rect 4940 3972 4942 4033
rect 5076 3972 5078 4033
rect 5212 3972 5214 4033
rect 5348 3972 5350 4033
rect 5664 3973 5666 4033
rect 5662 3972 5668 3973
rect 3838 3968 3839 3972
rect 3843 3968 3844 3972
rect 3838 3967 3844 3968
rect 4938 3971 4944 3972
rect 4938 3967 4939 3971
rect 4943 3967 4944 3971
rect 4938 3966 4944 3967
rect 5074 3971 5080 3972
rect 5074 3967 5075 3971
rect 5079 3967 5080 3971
rect 5074 3966 5080 3967
rect 5210 3971 5216 3972
rect 5210 3967 5211 3971
rect 5215 3967 5216 3971
rect 5210 3966 5216 3967
rect 5346 3971 5352 3972
rect 5346 3967 5347 3971
rect 5351 3967 5352 3971
rect 5662 3968 5663 3972
rect 5667 3968 5668 3972
rect 5662 3967 5668 3968
rect 5346 3966 5352 3967
rect 4966 3956 4972 3957
rect 3838 3955 3844 3956
rect 3838 3951 3839 3955
rect 3843 3951 3844 3955
rect 4966 3952 4967 3956
rect 4971 3952 4972 3956
rect 4966 3951 4972 3952
rect 5102 3956 5108 3957
rect 5102 3952 5103 3956
rect 5107 3952 5108 3956
rect 5102 3951 5108 3952
rect 5238 3956 5244 3957
rect 5238 3952 5239 3956
rect 5243 3952 5244 3956
rect 5238 3951 5244 3952
rect 5374 3956 5380 3957
rect 5374 3952 5375 3956
rect 5379 3952 5380 3956
rect 5374 3951 5380 3952
rect 5662 3955 5668 3956
rect 5662 3951 5663 3955
rect 5667 3951 5668 3955
rect 3838 3950 3844 3951
rect 110 3931 116 3932
rect 112 3867 114 3931
rect 668 3867 670 3932
rect 804 3867 806 3932
rect 940 3867 942 3932
rect 1084 3867 1086 3932
rect 1228 3867 1230 3932
rect 1372 3867 1374 3932
rect 1516 3867 1518 3932
rect 1652 3867 1654 3932
rect 1788 3867 1790 3932
rect 1934 3931 1940 3932
rect 1975 3934 1979 3935
rect 1936 3867 1938 3931
rect 1975 3929 1979 3930
rect 2759 3934 2763 3935
rect 2759 3929 2763 3930
rect 2911 3934 2915 3935
rect 2911 3929 2915 3930
rect 2927 3934 2931 3935
rect 2927 3929 2931 3930
rect 3071 3934 3075 3935
rect 3071 3929 3075 3930
rect 3215 3934 3219 3935
rect 3215 3929 3219 3930
rect 3239 3934 3243 3935
rect 3239 3929 3243 3930
rect 3367 3934 3371 3935
rect 3367 3929 3371 3930
rect 3415 3934 3419 3935
rect 3415 3929 3419 3930
rect 3519 3934 3523 3935
rect 3519 3929 3523 3930
rect 3591 3934 3595 3935
rect 3591 3929 3595 3930
rect 3671 3934 3675 3935
rect 3671 3929 3675 3930
rect 3799 3934 3803 3935
rect 3799 3929 3803 3930
rect 1976 3906 1978 3929
rect 1974 3905 1980 3906
rect 2760 3905 2762 3929
rect 2912 3905 2914 3929
rect 3072 3905 3074 3929
rect 3240 3905 3242 3929
rect 3416 3905 3418 3929
rect 3592 3905 3594 3929
rect 3800 3906 3802 3929
rect 3840 3927 3842 3950
rect 4968 3927 4970 3951
rect 5104 3927 5106 3951
rect 5240 3927 5242 3951
rect 5376 3927 5378 3951
rect 5662 3950 5668 3951
rect 5664 3927 5666 3950
rect 3839 3926 3843 3927
rect 3839 3921 3843 3922
rect 4687 3926 4691 3927
rect 4687 3921 4691 3922
rect 4847 3926 4851 3927
rect 4847 3921 4851 3922
rect 4967 3926 4971 3927
rect 4967 3921 4971 3922
rect 5015 3926 5019 3927
rect 5015 3921 5019 3922
rect 5103 3926 5107 3927
rect 5103 3921 5107 3922
rect 5191 3926 5195 3927
rect 5191 3921 5195 3922
rect 5239 3926 5243 3927
rect 5239 3921 5243 3922
rect 5375 3926 5379 3927
rect 5375 3921 5379 3922
rect 5543 3926 5547 3927
rect 5543 3921 5547 3922
rect 5663 3926 5667 3927
rect 5663 3921 5667 3922
rect 3798 3905 3804 3906
rect 1974 3901 1975 3905
rect 1979 3901 1980 3905
rect 1974 3900 1980 3901
rect 2758 3904 2764 3905
rect 2758 3900 2759 3904
rect 2763 3900 2764 3904
rect 2758 3899 2764 3900
rect 2910 3904 2916 3905
rect 2910 3900 2911 3904
rect 2915 3900 2916 3904
rect 2910 3899 2916 3900
rect 3070 3904 3076 3905
rect 3070 3900 3071 3904
rect 3075 3900 3076 3904
rect 3070 3899 3076 3900
rect 3238 3904 3244 3905
rect 3238 3900 3239 3904
rect 3243 3900 3244 3904
rect 3238 3899 3244 3900
rect 3414 3904 3420 3905
rect 3414 3900 3415 3904
rect 3419 3900 3420 3904
rect 3414 3899 3420 3900
rect 3590 3904 3596 3905
rect 3590 3900 3591 3904
rect 3595 3900 3596 3904
rect 3798 3901 3799 3905
rect 3803 3901 3804 3905
rect 3798 3900 3804 3901
rect 3590 3899 3596 3900
rect 3840 3898 3842 3921
rect 3838 3897 3844 3898
rect 4688 3897 4690 3921
rect 4848 3897 4850 3921
rect 5016 3897 5018 3921
rect 5192 3897 5194 3921
rect 5376 3897 5378 3921
rect 5544 3897 5546 3921
rect 5664 3898 5666 3921
rect 5662 3897 5668 3898
rect 3838 3893 3839 3897
rect 3843 3893 3844 3897
rect 3838 3892 3844 3893
rect 4686 3896 4692 3897
rect 4686 3892 4687 3896
rect 4691 3892 4692 3896
rect 4686 3891 4692 3892
rect 4846 3896 4852 3897
rect 4846 3892 4847 3896
rect 4851 3892 4852 3896
rect 4846 3891 4852 3892
rect 5014 3896 5020 3897
rect 5014 3892 5015 3896
rect 5019 3892 5020 3896
rect 5014 3891 5020 3892
rect 5190 3896 5196 3897
rect 5190 3892 5191 3896
rect 5195 3892 5196 3896
rect 5190 3891 5196 3892
rect 5374 3896 5380 3897
rect 5374 3892 5375 3896
rect 5379 3892 5380 3896
rect 5374 3891 5380 3892
rect 5542 3896 5548 3897
rect 5542 3892 5543 3896
rect 5547 3892 5548 3896
rect 5662 3893 5663 3897
rect 5667 3893 5668 3897
rect 5662 3892 5668 3893
rect 5542 3891 5548 3892
rect 2730 3889 2736 3890
rect 1974 3888 1980 3889
rect 1974 3884 1975 3888
rect 1979 3884 1980 3888
rect 2730 3885 2731 3889
rect 2735 3885 2736 3889
rect 2730 3884 2736 3885
rect 2882 3889 2888 3890
rect 2882 3885 2883 3889
rect 2887 3885 2888 3889
rect 2882 3884 2888 3885
rect 3042 3889 3048 3890
rect 3042 3885 3043 3889
rect 3047 3885 3048 3889
rect 3042 3884 3048 3885
rect 3210 3889 3216 3890
rect 3210 3885 3211 3889
rect 3215 3885 3216 3889
rect 3210 3884 3216 3885
rect 3386 3889 3392 3890
rect 3386 3885 3387 3889
rect 3391 3885 3392 3889
rect 3386 3884 3392 3885
rect 3562 3889 3568 3890
rect 3562 3885 3563 3889
rect 3567 3885 3568 3889
rect 3562 3884 3568 3885
rect 3798 3888 3804 3889
rect 3798 3884 3799 3888
rect 3803 3884 3804 3888
rect 1974 3883 1980 3884
rect 111 3866 115 3867
rect 111 3861 115 3862
rect 435 3866 439 3867
rect 435 3861 439 3862
rect 619 3866 623 3867
rect 619 3861 623 3862
rect 667 3866 671 3867
rect 667 3861 671 3862
rect 803 3866 807 3867
rect 803 3861 807 3862
rect 819 3866 823 3867
rect 819 3861 823 3862
rect 939 3866 943 3867
rect 939 3861 943 3862
rect 1027 3866 1031 3867
rect 1027 3861 1031 3862
rect 1083 3866 1087 3867
rect 1083 3861 1087 3862
rect 1227 3866 1231 3867
rect 1227 3861 1231 3862
rect 1251 3866 1255 3867
rect 1251 3861 1255 3862
rect 1371 3866 1375 3867
rect 1371 3861 1375 3862
rect 1483 3866 1487 3867
rect 1483 3861 1487 3862
rect 1515 3866 1519 3867
rect 1515 3861 1519 3862
rect 1651 3866 1655 3867
rect 1651 3861 1655 3862
rect 1723 3866 1727 3867
rect 1723 3861 1727 3862
rect 1787 3866 1791 3867
rect 1787 3861 1791 3862
rect 1935 3866 1939 3867
rect 1935 3861 1939 3862
rect 112 3801 114 3861
rect 110 3800 116 3801
rect 436 3800 438 3861
rect 620 3800 622 3861
rect 820 3800 822 3861
rect 1028 3800 1030 3861
rect 1252 3800 1254 3861
rect 1484 3800 1486 3861
rect 1724 3800 1726 3861
rect 1936 3801 1938 3861
rect 1976 3815 1978 3883
rect 2732 3815 2734 3884
rect 2884 3815 2886 3884
rect 3044 3815 3046 3884
rect 3212 3815 3214 3884
rect 3388 3815 3390 3884
rect 3564 3815 3566 3884
rect 3798 3883 3804 3884
rect 3800 3815 3802 3883
rect 4658 3881 4664 3882
rect 3838 3880 3844 3881
rect 3838 3876 3839 3880
rect 3843 3876 3844 3880
rect 4658 3877 4659 3881
rect 4663 3877 4664 3881
rect 4658 3876 4664 3877
rect 4818 3881 4824 3882
rect 4818 3877 4819 3881
rect 4823 3877 4824 3881
rect 4818 3876 4824 3877
rect 4986 3881 4992 3882
rect 4986 3877 4987 3881
rect 4991 3877 4992 3881
rect 4986 3876 4992 3877
rect 5162 3881 5168 3882
rect 5162 3877 5163 3881
rect 5167 3877 5168 3881
rect 5162 3876 5168 3877
rect 5346 3881 5352 3882
rect 5346 3877 5347 3881
rect 5351 3877 5352 3881
rect 5346 3876 5352 3877
rect 5514 3881 5520 3882
rect 5514 3877 5515 3881
rect 5519 3877 5520 3881
rect 5514 3876 5520 3877
rect 5662 3880 5668 3881
rect 5662 3876 5663 3880
rect 5667 3876 5668 3880
rect 3838 3875 3844 3876
rect 3840 3815 3842 3875
rect 4660 3815 4662 3876
rect 4820 3815 4822 3876
rect 4988 3815 4990 3876
rect 5164 3815 5166 3876
rect 5348 3815 5350 3876
rect 5516 3815 5518 3876
rect 5662 3875 5668 3876
rect 5664 3815 5666 3875
rect 1975 3814 1979 3815
rect 1975 3809 1979 3810
rect 2115 3814 2119 3815
rect 2115 3809 2119 3810
rect 2251 3814 2255 3815
rect 2251 3809 2255 3810
rect 2387 3814 2391 3815
rect 2387 3809 2391 3810
rect 2523 3814 2527 3815
rect 2523 3809 2527 3810
rect 2659 3814 2663 3815
rect 2659 3809 2663 3810
rect 2731 3814 2735 3815
rect 2731 3809 2735 3810
rect 2795 3814 2799 3815
rect 2795 3809 2799 3810
rect 2883 3814 2887 3815
rect 2883 3809 2887 3810
rect 2939 3814 2943 3815
rect 2939 3809 2943 3810
rect 3043 3814 3047 3815
rect 3043 3809 3047 3810
rect 3083 3814 3087 3815
rect 3083 3809 3087 3810
rect 3211 3814 3215 3815
rect 3211 3809 3215 3810
rect 3235 3814 3239 3815
rect 3235 3809 3239 3810
rect 3387 3814 3391 3815
rect 3387 3809 3391 3810
rect 3395 3814 3399 3815
rect 3395 3809 3399 3810
rect 3555 3814 3559 3815
rect 3555 3809 3559 3810
rect 3563 3814 3567 3815
rect 3563 3809 3567 3810
rect 3799 3814 3803 3815
rect 3799 3809 3803 3810
rect 3839 3814 3843 3815
rect 3839 3809 3843 3810
rect 4411 3814 4415 3815
rect 4411 3809 4415 3810
rect 4619 3814 4623 3815
rect 4619 3809 4623 3810
rect 4659 3814 4663 3815
rect 4659 3809 4663 3810
rect 4819 3814 4823 3815
rect 4819 3809 4823 3810
rect 4835 3814 4839 3815
rect 4835 3809 4839 3810
rect 4987 3814 4991 3815
rect 4987 3809 4991 3810
rect 5067 3814 5071 3815
rect 5067 3809 5071 3810
rect 5163 3814 5167 3815
rect 5163 3809 5167 3810
rect 5299 3814 5303 3815
rect 5299 3809 5303 3810
rect 5347 3814 5351 3815
rect 5347 3809 5351 3810
rect 5515 3814 5519 3815
rect 5515 3809 5519 3810
rect 5663 3814 5667 3815
rect 5663 3809 5667 3810
rect 1934 3800 1940 3801
rect 110 3796 111 3800
rect 115 3796 116 3800
rect 110 3795 116 3796
rect 434 3799 440 3800
rect 434 3795 435 3799
rect 439 3795 440 3799
rect 434 3794 440 3795
rect 618 3799 624 3800
rect 618 3795 619 3799
rect 623 3795 624 3799
rect 618 3794 624 3795
rect 818 3799 824 3800
rect 818 3795 819 3799
rect 823 3795 824 3799
rect 818 3794 824 3795
rect 1026 3799 1032 3800
rect 1026 3795 1027 3799
rect 1031 3795 1032 3799
rect 1026 3794 1032 3795
rect 1250 3799 1256 3800
rect 1250 3795 1251 3799
rect 1255 3795 1256 3799
rect 1250 3794 1256 3795
rect 1482 3799 1488 3800
rect 1482 3795 1483 3799
rect 1487 3795 1488 3799
rect 1482 3794 1488 3795
rect 1722 3799 1728 3800
rect 1722 3795 1723 3799
rect 1727 3795 1728 3799
rect 1934 3796 1935 3800
rect 1939 3796 1940 3800
rect 1934 3795 1940 3796
rect 1722 3794 1728 3795
rect 462 3784 468 3785
rect 110 3783 116 3784
rect 110 3779 111 3783
rect 115 3779 116 3783
rect 462 3780 463 3784
rect 467 3780 468 3784
rect 462 3779 468 3780
rect 646 3784 652 3785
rect 646 3780 647 3784
rect 651 3780 652 3784
rect 646 3779 652 3780
rect 846 3784 852 3785
rect 846 3780 847 3784
rect 851 3780 852 3784
rect 846 3779 852 3780
rect 1054 3784 1060 3785
rect 1054 3780 1055 3784
rect 1059 3780 1060 3784
rect 1054 3779 1060 3780
rect 1278 3784 1284 3785
rect 1278 3780 1279 3784
rect 1283 3780 1284 3784
rect 1278 3779 1284 3780
rect 1510 3784 1516 3785
rect 1510 3780 1511 3784
rect 1515 3780 1516 3784
rect 1510 3779 1516 3780
rect 1750 3784 1756 3785
rect 1750 3780 1751 3784
rect 1755 3780 1756 3784
rect 1750 3779 1756 3780
rect 1934 3783 1940 3784
rect 1934 3779 1935 3783
rect 1939 3779 1940 3783
rect 110 3778 116 3779
rect 112 3751 114 3778
rect 464 3751 466 3779
rect 648 3751 650 3779
rect 848 3751 850 3779
rect 1056 3751 1058 3779
rect 1280 3751 1282 3779
rect 1512 3751 1514 3779
rect 1752 3751 1754 3779
rect 1934 3778 1940 3779
rect 1936 3751 1938 3778
rect 111 3750 115 3751
rect 111 3745 115 3746
rect 231 3750 235 3751
rect 231 3745 235 3746
rect 431 3750 435 3751
rect 431 3745 435 3746
rect 463 3750 467 3751
rect 463 3745 467 3746
rect 647 3750 651 3751
rect 647 3745 651 3746
rect 655 3750 659 3751
rect 655 3745 659 3746
rect 847 3750 851 3751
rect 847 3745 851 3746
rect 895 3750 899 3751
rect 895 3745 899 3746
rect 1055 3750 1059 3751
rect 1055 3745 1059 3746
rect 1151 3750 1155 3751
rect 1151 3745 1155 3746
rect 1279 3750 1283 3751
rect 1279 3745 1283 3746
rect 1415 3750 1419 3751
rect 1415 3745 1419 3746
rect 1511 3750 1515 3751
rect 1511 3745 1515 3746
rect 1679 3750 1683 3751
rect 1679 3745 1683 3746
rect 1751 3750 1755 3751
rect 1751 3745 1755 3746
rect 1935 3750 1939 3751
rect 1976 3749 1978 3809
rect 1935 3745 1939 3746
rect 1974 3748 1980 3749
rect 2116 3748 2118 3809
rect 2252 3748 2254 3809
rect 2388 3748 2390 3809
rect 2524 3748 2526 3809
rect 2660 3748 2662 3809
rect 2796 3748 2798 3809
rect 2940 3748 2942 3809
rect 3084 3748 3086 3809
rect 3236 3748 3238 3809
rect 3396 3748 3398 3809
rect 3556 3748 3558 3809
rect 3800 3749 3802 3809
rect 3840 3749 3842 3809
rect 3798 3748 3804 3749
rect 112 3722 114 3745
rect 110 3721 116 3722
rect 232 3721 234 3745
rect 432 3721 434 3745
rect 656 3721 658 3745
rect 896 3721 898 3745
rect 1152 3721 1154 3745
rect 1416 3721 1418 3745
rect 1680 3721 1682 3745
rect 1936 3722 1938 3745
rect 1974 3744 1975 3748
rect 1979 3744 1980 3748
rect 1974 3743 1980 3744
rect 2114 3747 2120 3748
rect 2114 3743 2115 3747
rect 2119 3743 2120 3747
rect 2114 3742 2120 3743
rect 2250 3747 2256 3748
rect 2250 3743 2251 3747
rect 2255 3743 2256 3747
rect 2250 3742 2256 3743
rect 2386 3747 2392 3748
rect 2386 3743 2387 3747
rect 2391 3743 2392 3747
rect 2386 3742 2392 3743
rect 2522 3747 2528 3748
rect 2522 3743 2523 3747
rect 2527 3743 2528 3747
rect 2522 3742 2528 3743
rect 2658 3747 2664 3748
rect 2658 3743 2659 3747
rect 2663 3743 2664 3747
rect 2658 3742 2664 3743
rect 2794 3747 2800 3748
rect 2794 3743 2795 3747
rect 2799 3743 2800 3747
rect 2794 3742 2800 3743
rect 2938 3747 2944 3748
rect 2938 3743 2939 3747
rect 2943 3743 2944 3747
rect 2938 3742 2944 3743
rect 3082 3747 3088 3748
rect 3082 3743 3083 3747
rect 3087 3743 3088 3747
rect 3082 3742 3088 3743
rect 3234 3747 3240 3748
rect 3234 3743 3235 3747
rect 3239 3743 3240 3747
rect 3234 3742 3240 3743
rect 3394 3747 3400 3748
rect 3394 3743 3395 3747
rect 3399 3743 3400 3747
rect 3394 3742 3400 3743
rect 3554 3747 3560 3748
rect 3554 3743 3555 3747
rect 3559 3743 3560 3747
rect 3798 3744 3799 3748
rect 3803 3744 3804 3748
rect 3798 3743 3804 3744
rect 3838 3748 3844 3749
rect 4412 3748 4414 3809
rect 4620 3748 4622 3809
rect 4836 3748 4838 3809
rect 5068 3748 5070 3809
rect 5300 3748 5302 3809
rect 5516 3748 5518 3809
rect 5664 3749 5666 3809
rect 5662 3748 5668 3749
rect 3838 3744 3839 3748
rect 3843 3744 3844 3748
rect 3838 3743 3844 3744
rect 4410 3747 4416 3748
rect 4410 3743 4411 3747
rect 4415 3743 4416 3747
rect 3554 3742 3560 3743
rect 4410 3742 4416 3743
rect 4618 3747 4624 3748
rect 4618 3743 4619 3747
rect 4623 3743 4624 3747
rect 4618 3742 4624 3743
rect 4834 3747 4840 3748
rect 4834 3743 4835 3747
rect 4839 3743 4840 3747
rect 4834 3742 4840 3743
rect 5066 3747 5072 3748
rect 5066 3743 5067 3747
rect 5071 3743 5072 3747
rect 5066 3742 5072 3743
rect 5298 3747 5304 3748
rect 5298 3743 5299 3747
rect 5303 3743 5304 3747
rect 5298 3742 5304 3743
rect 5514 3747 5520 3748
rect 5514 3743 5515 3747
rect 5519 3743 5520 3747
rect 5662 3744 5663 3748
rect 5667 3744 5668 3748
rect 5662 3743 5668 3744
rect 5514 3742 5520 3743
rect 2142 3732 2148 3733
rect 1974 3731 1980 3732
rect 1974 3727 1975 3731
rect 1979 3727 1980 3731
rect 2142 3728 2143 3732
rect 2147 3728 2148 3732
rect 2142 3727 2148 3728
rect 2278 3732 2284 3733
rect 2278 3728 2279 3732
rect 2283 3728 2284 3732
rect 2278 3727 2284 3728
rect 2414 3732 2420 3733
rect 2414 3728 2415 3732
rect 2419 3728 2420 3732
rect 2414 3727 2420 3728
rect 2550 3732 2556 3733
rect 2550 3728 2551 3732
rect 2555 3728 2556 3732
rect 2550 3727 2556 3728
rect 2686 3732 2692 3733
rect 2686 3728 2687 3732
rect 2691 3728 2692 3732
rect 2686 3727 2692 3728
rect 2822 3732 2828 3733
rect 2822 3728 2823 3732
rect 2827 3728 2828 3732
rect 2822 3727 2828 3728
rect 2966 3732 2972 3733
rect 2966 3728 2967 3732
rect 2971 3728 2972 3732
rect 2966 3727 2972 3728
rect 3110 3732 3116 3733
rect 3110 3728 3111 3732
rect 3115 3728 3116 3732
rect 3110 3727 3116 3728
rect 3262 3732 3268 3733
rect 3262 3728 3263 3732
rect 3267 3728 3268 3732
rect 3262 3727 3268 3728
rect 3422 3732 3428 3733
rect 3422 3728 3423 3732
rect 3427 3728 3428 3732
rect 3422 3727 3428 3728
rect 3582 3732 3588 3733
rect 4438 3732 4444 3733
rect 3582 3728 3583 3732
rect 3587 3728 3588 3732
rect 3582 3727 3588 3728
rect 3798 3731 3804 3732
rect 3798 3727 3799 3731
rect 3803 3727 3804 3731
rect 1974 3726 1980 3727
rect 1934 3721 1940 3722
rect 110 3717 111 3721
rect 115 3717 116 3721
rect 110 3716 116 3717
rect 230 3720 236 3721
rect 230 3716 231 3720
rect 235 3716 236 3720
rect 230 3715 236 3716
rect 430 3720 436 3721
rect 430 3716 431 3720
rect 435 3716 436 3720
rect 430 3715 436 3716
rect 654 3720 660 3721
rect 654 3716 655 3720
rect 659 3716 660 3720
rect 654 3715 660 3716
rect 894 3720 900 3721
rect 894 3716 895 3720
rect 899 3716 900 3720
rect 894 3715 900 3716
rect 1150 3720 1156 3721
rect 1150 3716 1151 3720
rect 1155 3716 1156 3720
rect 1150 3715 1156 3716
rect 1414 3720 1420 3721
rect 1414 3716 1415 3720
rect 1419 3716 1420 3720
rect 1414 3715 1420 3716
rect 1678 3720 1684 3721
rect 1678 3716 1679 3720
rect 1683 3716 1684 3720
rect 1934 3717 1935 3721
rect 1939 3717 1940 3721
rect 1934 3716 1940 3717
rect 1678 3715 1684 3716
rect 202 3705 208 3706
rect 110 3704 116 3705
rect 110 3700 111 3704
rect 115 3700 116 3704
rect 202 3701 203 3705
rect 207 3701 208 3705
rect 202 3700 208 3701
rect 402 3705 408 3706
rect 402 3701 403 3705
rect 407 3701 408 3705
rect 402 3700 408 3701
rect 626 3705 632 3706
rect 626 3701 627 3705
rect 631 3701 632 3705
rect 626 3700 632 3701
rect 866 3705 872 3706
rect 866 3701 867 3705
rect 871 3701 872 3705
rect 866 3700 872 3701
rect 1122 3705 1128 3706
rect 1122 3701 1123 3705
rect 1127 3701 1128 3705
rect 1122 3700 1128 3701
rect 1386 3705 1392 3706
rect 1386 3701 1387 3705
rect 1391 3701 1392 3705
rect 1386 3700 1392 3701
rect 1650 3705 1656 3706
rect 1650 3701 1651 3705
rect 1655 3701 1656 3705
rect 1650 3700 1656 3701
rect 1934 3704 1940 3705
rect 1934 3700 1935 3704
rect 1939 3700 1940 3704
rect 110 3699 116 3700
rect 112 3631 114 3699
rect 204 3631 206 3700
rect 404 3631 406 3700
rect 628 3631 630 3700
rect 868 3631 870 3700
rect 1124 3631 1126 3700
rect 1388 3631 1390 3700
rect 1652 3631 1654 3700
rect 1934 3699 1940 3700
rect 1936 3631 1938 3699
rect 1976 3695 1978 3726
rect 2144 3695 2146 3727
rect 2280 3695 2282 3727
rect 2416 3695 2418 3727
rect 2552 3695 2554 3727
rect 2688 3695 2690 3727
rect 2824 3695 2826 3727
rect 2968 3695 2970 3727
rect 3112 3695 3114 3727
rect 3264 3695 3266 3727
rect 3424 3695 3426 3727
rect 3584 3695 3586 3727
rect 3798 3726 3804 3727
rect 3838 3731 3844 3732
rect 3838 3727 3839 3731
rect 3843 3727 3844 3731
rect 4438 3728 4439 3732
rect 4443 3728 4444 3732
rect 4438 3727 4444 3728
rect 4646 3732 4652 3733
rect 4646 3728 4647 3732
rect 4651 3728 4652 3732
rect 4646 3727 4652 3728
rect 4862 3732 4868 3733
rect 4862 3728 4863 3732
rect 4867 3728 4868 3732
rect 4862 3727 4868 3728
rect 5094 3732 5100 3733
rect 5094 3728 5095 3732
rect 5099 3728 5100 3732
rect 5094 3727 5100 3728
rect 5326 3732 5332 3733
rect 5326 3728 5327 3732
rect 5331 3728 5332 3732
rect 5326 3727 5332 3728
rect 5542 3732 5548 3733
rect 5542 3728 5543 3732
rect 5547 3728 5548 3732
rect 5542 3727 5548 3728
rect 5662 3731 5668 3732
rect 5662 3727 5663 3731
rect 5667 3727 5668 3731
rect 3838 3726 3844 3727
rect 3800 3695 3802 3726
rect 1975 3694 1979 3695
rect 1975 3689 1979 3690
rect 2143 3694 2147 3695
rect 2143 3689 2147 3690
rect 2231 3694 2235 3695
rect 2231 3689 2235 3690
rect 2279 3694 2283 3695
rect 2279 3689 2283 3690
rect 2415 3694 2419 3695
rect 2415 3689 2419 3690
rect 2447 3694 2451 3695
rect 2447 3689 2451 3690
rect 2551 3694 2555 3695
rect 2551 3689 2555 3690
rect 2663 3694 2667 3695
rect 2663 3689 2667 3690
rect 2687 3694 2691 3695
rect 2687 3689 2691 3690
rect 2823 3694 2827 3695
rect 2823 3689 2827 3690
rect 2871 3694 2875 3695
rect 2871 3689 2875 3690
rect 2967 3694 2971 3695
rect 2967 3689 2971 3690
rect 3079 3694 3083 3695
rect 3079 3689 3083 3690
rect 3111 3694 3115 3695
rect 3111 3689 3115 3690
rect 3263 3694 3267 3695
rect 3263 3689 3267 3690
rect 3287 3694 3291 3695
rect 3287 3689 3291 3690
rect 3423 3694 3427 3695
rect 3423 3689 3427 3690
rect 3495 3694 3499 3695
rect 3495 3689 3499 3690
rect 3583 3694 3587 3695
rect 3583 3689 3587 3690
rect 3679 3694 3683 3695
rect 3679 3689 3683 3690
rect 3799 3694 3803 3695
rect 3799 3689 3803 3690
rect 1976 3666 1978 3689
rect 1974 3665 1980 3666
rect 2232 3665 2234 3689
rect 2448 3665 2450 3689
rect 2664 3665 2666 3689
rect 2872 3665 2874 3689
rect 3080 3665 3082 3689
rect 3288 3665 3290 3689
rect 3496 3665 3498 3689
rect 3680 3665 3682 3689
rect 3800 3666 3802 3689
rect 3840 3679 3842 3726
rect 4440 3679 4442 3727
rect 4648 3679 4650 3727
rect 4864 3679 4866 3727
rect 5096 3679 5098 3727
rect 5328 3679 5330 3727
rect 5544 3679 5546 3727
rect 5662 3726 5668 3727
rect 5664 3679 5666 3726
rect 3839 3678 3843 3679
rect 3839 3673 3843 3674
rect 3887 3678 3891 3679
rect 3887 3673 3891 3674
rect 4047 3678 4051 3679
rect 4047 3673 4051 3674
rect 4247 3678 4251 3679
rect 4247 3673 4251 3674
rect 4439 3678 4443 3679
rect 4439 3673 4443 3674
rect 4479 3678 4483 3679
rect 4479 3673 4483 3674
rect 4647 3678 4651 3679
rect 4647 3673 4651 3674
rect 4727 3678 4731 3679
rect 4727 3673 4731 3674
rect 4863 3678 4867 3679
rect 4863 3673 4867 3674
rect 4999 3678 5003 3679
rect 4999 3673 5003 3674
rect 5095 3678 5099 3679
rect 5095 3673 5099 3674
rect 5279 3678 5283 3679
rect 5279 3673 5283 3674
rect 5327 3678 5331 3679
rect 5327 3673 5331 3674
rect 5543 3678 5547 3679
rect 5543 3673 5547 3674
rect 5663 3678 5667 3679
rect 5663 3673 5667 3674
rect 3798 3665 3804 3666
rect 1974 3661 1975 3665
rect 1979 3661 1980 3665
rect 1974 3660 1980 3661
rect 2230 3664 2236 3665
rect 2230 3660 2231 3664
rect 2235 3660 2236 3664
rect 2230 3659 2236 3660
rect 2446 3664 2452 3665
rect 2446 3660 2447 3664
rect 2451 3660 2452 3664
rect 2446 3659 2452 3660
rect 2662 3664 2668 3665
rect 2662 3660 2663 3664
rect 2667 3660 2668 3664
rect 2662 3659 2668 3660
rect 2870 3664 2876 3665
rect 2870 3660 2871 3664
rect 2875 3660 2876 3664
rect 2870 3659 2876 3660
rect 3078 3664 3084 3665
rect 3078 3660 3079 3664
rect 3083 3660 3084 3664
rect 3078 3659 3084 3660
rect 3286 3664 3292 3665
rect 3286 3660 3287 3664
rect 3291 3660 3292 3664
rect 3286 3659 3292 3660
rect 3494 3664 3500 3665
rect 3494 3660 3495 3664
rect 3499 3660 3500 3664
rect 3494 3659 3500 3660
rect 3678 3664 3684 3665
rect 3678 3660 3679 3664
rect 3683 3660 3684 3664
rect 3798 3661 3799 3665
rect 3803 3661 3804 3665
rect 3798 3660 3804 3661
rect 3678 3659 3684 3660
rect 3840 3650 3842 3673
rect 2202 3649 2208 3650
rect 1974 3648 1980 3649
rect 1974 3644 1975 3648
rect 1979 3644 1980 3648
rect 2202 3645 2203 3649
rect 2207 3645 2208 3649
rect 2202 3644 2208 3645
rect 2418 3649 2424 3650
rect 2418 3645 2419 3649
rect 2423 3645 2424 3649
rect 2418 3644 2424 3645
rect 2634 3649 2640 3650
rect 2634 3645 2635 3649
rect 2639 3645 2640 3649
rect 2634 3644 2640 3645
rect 2842 3649 2848 3650
rect 2842 3645 2843 3649
rect 2847 3645 2848 3649
rect 2842 3644 2848 3645
rect 3050 3649 3056 3650
rect 3050 3645 3051 3649
rect 3055 3645 3056 3649
rect 3050 3644 3056 3645
rect 3258 3649 3264 3650
rect 3258 3645 3259 3649
rect 3263 3645 3264 3649
rect 3258 3644 3264 3645
rect 3466 3649 3472 3650
rect 3466 3645 3467 3649
rect 3471 3645 3472 3649
rect 3466 3644 3472 3645
rect 3650 3649 3656 3650
rect 3838 3649 3844 3650
rect 3888 3649 3890 3673
rect 4048 3649 4050 3673
rect 4248 3649 4250 3673
rect 4480 3649 4482 3673
rect 4728 3649 4730 3673
rect 5000 3649 5002 3673
rect 5280 3649 5282 3673
rect 5544 3649 5546 3673
rect 5664 3650 5666 3673
rect 5662 3649 5668 3650
rect 3650 3645 3651 3649
rect 3655 3645 3656 3649
rect 3650 3644 3656 3645
rect 3798 3648 3804 3649
rect 3798 3644 3799 3648
rect 3803 3644 3804 3648
rect 3838 3645 3839 3649
rect 3843 3645 3844 3649
rect 3838 3644 3844 3645
rect 3886 3648 3892 3649
rect 3886 3644 3887 3648
rect 3891 3644 3892 3648
rect 1974 3643 1980 3644
rect 111 3630 115 3631
rect 111 3625 115 3626
rect 131 3630 135 3631
rect 131 3625 135 3626
rect 203 3630 207 3631
rect 203 3625 207 3626
rect 315 3630 319 3631
rect 315 3625 319 3626
rect 403 3630 407 3631
rect 403 3625 407 3626
rect 539 3630 543 3631
rect 539 3625 543 3626
rect 627 3630 631 3631
rect 627 3625 631 3626
rect 787 3630 791 3631
rect 787 3625 791 3626
rect 867 3630 871 3631
rect 867 3625 871 3626
rect 1043 3630 1047 3631
rect 1043 3625 1047 3626
rect 1123 3630 1127 3631
rect 1123 3625 1127 3626
rect 1315 3630 1319 3631
rect 1315 3625 1319 3626
rect 1387 3630 1391 3631
rect 1387 3625 1391 3626
rect 1587 3630 1591 3631
rect 1587 3625 1591 3626
rect 1651 3630 1655 3631
rect 1651 3625 1655 3626
rect 1935 3630 1939 3631
rect 1935 3625 1939 3626
rect 112 3565 114 3625
rect 110 3564 116 3565
rect 132 3564 134 3625
rect 316 3564 318 3625
rect 540 3564 542 3625
rect 788 3564 790 3625
rect 1044 3564 1046 3625
rect 1316 3564 1318 3625
rect 1588 3564 1590 3625
rect 1936 3565 1938 3625
rect 1976 3567 1978 3643
rect 2204 3567 2206 3644
rect 2420 3567 2422 3644
rect 2636 3567 2638 3644
rect 2844 3567 2846 3644
rect 3052 3567 3054 3644
rect 3260 3567 3262 3644
rect 3468 3567 3470 3644
rect 3652 3567 3654 3644
rect 3798 3643 3804 3644
rect 3886 3643 3892 3644
rect 4046 3648 4052 3649
rect 4046 3644 4047 3648
rect 4051 3644 4052 3648
rect 4046 3643 4052 3644
rect 4246 3648 4252 3649
rect 4246 3644 4247 3648
rect 4251 3644 4252 3648
rect 4246 3643 4252 3644
rect 4478 3648 4484 3649
rect 4478 3644 4479 3648
rect 4483 3644 4484 3648
rect 4478 3643 4484 3644
rect 4726 3648 4732 3649
rect 4726 3644 4727 3648
rect 4731 3644 4732 3648
rect 4726 3643 4732 3644
rect 4998 3648 5004 3649
rect 4998 3644 4999 3648
rect 5003 3644 5004 3648
rect 4998 3643 5004 3644
rect 5278 3648 5284 3649
rect 5278 3644 5279 3648
rect 5283 3644 5284 3648
rect 5278 3643 5284 3644
rect 5542 3648 5548 3649
rect 5542 3644 5543 3648
rect 5547 3644 5548 3648
rect 5662 3645 5663 3649
rect 5667 3645 5668 3649
rect 5662 3644 5668 3645
rect 5542 3643 5548 3644
rect 3800 3567 3802 3643
rect 3858 3633 3864 3634
rect 3838 3632 3844 3633
rect 3838 3628 3839 3632
rect 3843 3628 3844 3632
rect 3858 3629 3859 3633
rect 3863 3629 3864 3633
rect 3858 3628 3864 3629
rect 4018 3633 4024 3634
rect 4018 3629 4019 3633
rect 4023 3629 4024 3633
rect 4018 3628 4024 3629
rect 4218 3633 4224 3634
rect 4218 3629 4219 3633
rect 4223 3629 4224 3633
rect 4218 3628 4224 3629
rect 4450 3633 4456 3634
rect 4450 3629 4451 3633
rect 4455 3629 4456 3633
rect 4450 3628 4456 3629
rect 4698 3633 4704 3634
rect 4698 3629 4699 3633
rect 4703 3629 4704 3633
rect 4698 3628 4704 3629
rect 4970 3633 4976 3634
rect 4970 3629 4971 3633
rect 4975 3629 4976 3633
rect 4970 3628 4976 3629
rect 5250 3633 5256 3634
rect 5250 3629 5251 3633
rect 5255 3629 5256 3633
rect 5250 3628 5256 3629
rect 5514 3633 5520 3634
rect 5514 3629 5515 3633
rect 5519 3629 5520 3633
rect 5514 3628 5520 3629
rect 5662 3632 5668 3633
rect 5662 3628 5663 3632
rect 5667 3628 5668 3632
rect 3838 3627 3844 3628
rect 1975 3566 1979 3567
rect 1934 3564 1940 3565
rect 110 3560 111 3564
rect 115 3560 116 3564
rect 110 3559 116 3560
rect 130 3563 136 3564
rect 130 3559 131 3563
rect 135 3559 136 3563
rect 130 3558 136 3559
rect 314 3563 320 3564
rect 314 3559 315 3563
rect 319 3559 320 3563
rect 314 3558 320 3559
rect 538 3563 544 3564
rect 538 3559 539 3563
rect 543 3559 544 3563
rect 538 3558 544 3559
rect 786 3563 792 3564
rect 786 3559 787 3563
rect 791 3559 792 3563
rect 786 3558 792 3559
rect 1042 3563 1048 3564
rect 1042 3559 1043 3563
rect 1047 3559 1048 3563
rect 1042 3558 1048 3559
rect 1314 3563 1320 3564
rect 1314 3559 1315 3563
rect 1319 3559 1320 3563
rect 1314 3558 1320 3559
rect 1586 3563 1592 3564
rect 1586 3559 1587 3563
rect 1591 3559 1592 3563
rect 1934 3560 1935 3564
rect 1939 3560 1940 3564
rect 1975 3561 1979 3562
rect 2163 3566 2167 3567
rect 2163 3561 2167 3562
rect 2203 3566 2207 3567
rect 2203 3561 2207 3562
rect 2299 3566 2303 3567
rect 2299 3561 2303 3562
rect 2419 3566 2423 3567
rect 2419 3561 2423 3562
rect 2435 3566 2439 3567
rect 2435 3561 2439 3562
rect 2571 3566 2575 3567
rect 2571 3561 2575 3562
rect 2635 3566 2639 3567
rect 2635 3561 2639 3562
rect 2843 3566 2847 3567
rect 2843 3561 2847 3562
rect 3051 3566 3055 3567
rect 3051 3561 3055 3562
rect 3259 3566 3263 3567
rect 3259 3561 3263 3562
rect 3467 3566 3471 3567
rect 3467 3561 3471 3562
rect 3651 3566 3655 3567
rect 3651 3561 3655 3562
rect 3799 3566 3803 3567
rect 3799 3561 3803 3562
rect 1934 3559 1940 3560
rect 1586 3558 1592 3559
rect 158 3548 164 3549
rect 110 3547 116 3548
rect 110 3543 111 3547
rect 115 3543 116 3547
rect 158 3544 159 3548
rect 163 3544 164 3548
rect 158 3543 164 3544
rect 342 3548 348 3549
rect 342 3544 343 3548
rect 347 3544 348 3548
rect 342 3543 348 3544
rect 566 3548 572 3549
rect 566 3544 567 3548
rect 571 3544 572 3548
rect 566 3543 572 3544
rect 814 3548 820 3549
rect 814 3544 815 3548
rect 819 3544 820 3548
rect 814 3543 820 3544
rect 1070 3548 1076 3549
rect 1070 3544 1071 3548
rect 1075 3544 1076 3548
rect 1070 3543 1076 3544
rect 1342 3548 1348 3549
rect 1342 3544 1343 3548
rect 1347 3544 1348 3548
rect 1342 3543 1348 3544
rect 1614 3548 1620 3549
rect 1614 3544 1615 3548
rect 1619 3544 1620 3548
rect 1614 3543 1620 3544
rect 1934 3547 1940 3548
rect 1934 3543 1935 3547
rect 1939 3543 1940 3547
rect 110 3542 116 3543
rect 112 3507 114 3542
rect 160 3507 162 3543
rect 344 3507 346 3543
rect 568 3507 570 3543
rect 816 3507 818 3543
rect 1072 3507 1074 3543
rect 1344 3507 1346 3543
rect 1616 3507 1618 3543
rect 1934 3542 1940 3543
rect 1936 3507 1938 3542
rect 111 3506 115 3507
rect 111 3501 115 3502
rect 159 3506 163 3507
rect 159 3501 163 3502
rect 335 3506 339 3507
rect 335 3501 339 3502
rect 343 3506 347 3507
rect 343 3501 347 3502
rect 551 3506 555 3507
rect 551 3501 555 3502
rect 567 3506 571 3507
rect 567 3501 571 3502
rect 791 3506 795 3507
rect 791 3501 795 3502
rect 815 3506 819 3507
rect 815 3501 819 3502
rect 1039 3506 1043 3507
rect 1039 3501 1043 3502
rect 1071 3506 1075 3507
rect 1071 3501 1075 3502
rect 1295 3506 1299 3507
rect 1295 3501 1299 3502
rect 1343 3506 1347 3507
rect 1343 3501 1347 3502
rect 1559 3506 1563 3507
rect 1559 3501 1563 3502
rect 1615 3506 1619 3507
rect 1615 3501 1619 3502
rect 1935 3506 1939 3507
rect 1935 3501 1939 3502
rect 1976 3501 1978 3561
rect 112 3478 114 3501
rect 110 3477 116 3478
rect 160 3477 162 3501
rect 336 3477 338 3501
rect 552 3477 554 3501
rect 792 3477 794 3501
rect 1040 3477 1042 3501
rect 1296 3477 1298 3501
rect 1560 3477 1562 3501
rect 1936 3478 1938 3501
rect 1974 3500 1980 3501
rect 2164 3500 2166 3561
rect 2300 3500 2302 3561
rect 2436 3500 2438 3561
rect 2572 3500 2574 3561
rect 3800 3501 3802 3561
rect 3840 3555 3842 3627
rect 3860 3555 3862 3628
rect 4020 3555 4022 3628
rect 4220 3555 4222 3628
rect 4452 3555 4454 3628
rect 4700 3555 4702 3628
rect 4972 3555 4974 3628
rect 5252 3555 5254 3628
rect 5516 3555 5518 3628
rect 5662 3627 5668 3628
rect 5664 3555 5666 3627
rect 3839 3554 3843 3555
rect 3839 3549 3843 3550
rect 3859 3554 3863 3555
rect 3859 3549 3863 3550
rect 3995 3554 3999 3555
rect 3995 3549 3999 3550
rect 4019 3554 4023 3555
rect 4019 3549 4023 3550
rect 4131 3554 4135 3555
rect 4131 3549 4135 3550
rect 4219 3554 4223 3555
rect 4219 3549 4223 3550
rect 4267 3554 4271 3555
rect 4267 3549 4271 3550
rect 4403 3554 4407 3555
rect 4403 3549 4407 3550
rect 4451 3554 4455 3555
rect 4451 3549 4455 3550
rect 4539 3554 4543 3555
rect 4539 3549 4543 3550
rect 4699 3554 4703 3555
rect 4699 3549 4703 3550
rect 4891 3554 4895 3555
rect 4891 3549 4895 3550
rect 4971 3554 4975 3555
rect 4971 3549 4975 3550
rect 5099 3554 5103 3555
rect 5099 3549 5103 3550
rect 5251 3554 5255 3555
rect 5251 3549 5255 3550
rect 5315 3554 5319 3555
rect 5315 3549 5319 3550
rect 5515 3554 5519 3555
rect 5515 3549 5519 3550
rect 5663 3554 5667 3555
rect 5663 3549 5667 3550
rect 3798 3500 3804 3501
rect 1974 3496 1975 3500
rect 1979 3496 1980 3500
rect 1974 3495 1980 3496
rect 2162 3499 2168 3500
rect 2162 3495 2163 3499
rect 2167 3495 2168 3499
rect 2162 3494 2168 3495
rect 2298 3499 2304 3500
rect 2298 3495 2299 3499
rect 2303 3495 2304 3499
rect 2298 3494 2304 3495
rect 2434 3499 2440 3500
rect 2434 3495 2435 3499
rect 2439 3495 2440 3499
rect 2434 3494 2440 3495
rect 2570 3499 2576 3500
rect 2570 3495 2571 3499
rect 2575 3495 2576 3499
rect 3798 3496 3799 3500
rect 3803 3496 3804 3500
rect 3798 3495 3804 3496
rect 2570 3494 2576 3495
rect 3840 3489 3842 3549
rect 3838 3488 3844 3489
rect 3860 3488 3862 3549
rect 3996 3488 3998 3549
rect 4132 3488 4134 3549
rect 4268 3488 4270 3549
rect 4404 3488 4406 3549
rect 4540 3488 4542 3549
rect 4700 3488 4702 3549
rect 4892 3488 4894 3549
rect 5100 3488 5102 3549
rect 5316 3488 5318 3549
rect 5516 3488 5518 3549
rect 5664 3489 5666 3549
rect 5662 3488 5668 3489
rect 2190 3484 2196 3485
rect 1974 3483 1980 3484
rect 1974 3479 1975 3483
rect 1979 3479 1980 3483
rect 2190 3480 2191 3484
rect 2195 3480 2196 3484
rect 2190 3479 2196 3480
rect 2326 3484 2332 3485
rect 2326 3480 2327 3484
rect 2331 3480 2332 3484
rect 2326 3479 2332 3480
rect 2462 3484 2468 3485
rect 2462 3480 2463 3484
rect 2467 3480 2468 3484
rect 2462 3479 2468 3480
rect 2598 3484 2604 3485
rect 3838 3484 3839 3488
rect 3843 3484 3844 3488
rect 2598 3480 2599 3484
rect 2603 3480 2604 3484
rect 2598 3479 2604 3480
rect 3798 3483 3804 3484
rect 3838 3483 3844 3484
rect 3858 3487 3864 3488
rect 3858 3483 3859 3487
rect 3863 3483 3864 3487
rect 3798 3479 3799 3483
rect 3803 3479 3804 3483
rect 3858 3482 3864 3483
rect 3994 3487 4000 3488
rect 3994 3483 3995 3487
rect 3999 3483 4000 3487
rect 3994 3482 4000 3483
rect 4130 3487 4136 3488
rect 4130 3483 4131 3487
rect 4135 3483 4136 3487
rect 4130 3482 4136 3483
rect 4266 3487 4272 3488
rect 4266 3483 4267 3487
rect 4271 3483 4272 3487
rect 4266 3482 4272 3483
rect 4402 3487 4408 3488
rect 4402 3483 4403 3487
rect 4407 3483 4408 3487
rect 4402 3482 4408 3483
rect 4538 3487 4544 3488
rect 4538 3483 4539 3487
rect 4543 3483 4544 3487
rect 4538 3482 4544 3483
rect 4698 3487 4704 3488
rect 4698 3483 4699 3487
rect 4703 3483 4704 3487
rect 4698 3482 4704 3483
rect 4890 3487 4896 3488
rect 4890 3483 4891 3487
rect 4895 3483 4896 3487
rect 4890 3482 4896 3483
rect 5098 3487 5104 3488
rect 5098 3483 5099 3487
rect 5103 3483 5104 3487
rect 5098 3482 5104 3483
rect 5314 3487 5320 3488
rect 5314 3483 5315 3487
rect 5319 3483 5320 3487
rect 5314 3482 5320 3483
rect 5514 3487 5520 3488
rect 5514 3483 5515 3487
rect 5519 3483 5520 3487
rect 5662 3484 5663 3488
rect 5667 3484 5668 3488
rect 5662 3483 5668 3484
rect 5514 3482 5520 3483
rect 1974 3478 1980 3479
rect 1934 3477 1940 3478
rect 110 3473 111 3477
rect 115 3473 116 3477
rect 110 3472 116 3473
rect 158 3476 164 3477
rect 158 3472 159 3476
rect 163 3472 164 3476
rect 158 3471 164 3472
rect 334 3476 340 3477
rect 334 3472 335 3476
rect 339 3472 340 3476
rect 334 3471 340 3472
rect 550 3476 556 3477
rect 550 3472 551 3476
rect 555 3472 556 3476
rect 550 3471 556 3472
rect 790 3476 796 3477
rect 790 3472 791 3476
rect 795 3472 796 3476
rect 790 3471 796 3472
rect 1038 3476 1044 3477
rect 1038 3472 1039 3476
rect 1043 3472 1044 3476
rect 1038 3471 1044 3472
rect 1294 3476 1300 3477
rect 1294 3472 1295 3476
rect 1299 3472 1300 3476
rect 1294 3471 1300 3472
rect 1558 3476 1564 3477
rect 1558 3472 1559 3476
rect 1563 3472 1564 3476
rect 1934 3473 1935 3477
rect 1939 3473 1940 3477
rect 1934 3472 1940 3473
rect 1558 3471 1564 3472
rect 130 3461 136 3462
rect 110 3460 116 3461
rect 110 3456 111 3460
rect 115 3456 116 3460
rect 130 3457 131 3461
rect 135 3457 136 3461
rect 130 3456 136 3457
rect 306 3461 312 3462
rect 306 3457 307 3461
rect 311 3457 312 3461
rect 306 3456 312 3457
rect 522 3461 528 3462
rect 522 3457 523 3461
rect 527 3457 528 3461
rect 522 3456 528 3457
rect 762 3461 768 3462
rect 762 3457 763 3461
rect 767 3457 768 3461
rect 762 3456 768 3457
rect 1010 3461 1016 3462
rect 1010 3457 1011 3461
rect 1015 3457 1016 3461
rect 1010 3456 1016 3457
rect 1266 3461 1272 3462
rect 1266 3457 1267 3461
rect 1271 3457 1272 3461
rect 1266 3456 1272 3457
rect 1530 3461 1536 3462
rect 1530 3457 1531 3461
rect 1535 3457 1536 3461
rect 1530 3456 1536 3457
rect 1934 3460 1940 3461
rect 1934 3456 1935 3460
rect 1939 3456 1940 3460
rect 110 3455 116 3456
rect 112 3387 114 3455
rect 132 3387 134 3456
rect 308 3387 310 3456
rect 524 3387 526 3456
rect 764 3387 766 3456
rect 1012 3387 1014 3456
rect 1268 3387 1270 3456
rect 1532 3387 1534 3456
rect 1934 3455 1940 3456
rect 1936 3387 1938 3455
rect 1976 3419 1978 3478
rect 2192 3419 2194 3479
rect 2328 3419 2330 3479
rect 2464 3419 2466 3479
rect 2600 3419 2602 3479
rect 3798 3478 3804 3479
rect 3800 3419 3802 3478
rect 3886 3472 3892 3473
rect 3838 3471 3844 3472
rect 3838 3467 3839 3471
rect 3843 3467 3844 3471
rect 3886 3468 3887 3472
rect 3891 3468 3892 3472
rect 3886 3467 3892 3468
rect 4022 3472 4028 3473
rect 4022 3468 4023 3472
rect 4027 3468 4028 3472
rect 4022 3467 4028 3468
rect 4158 3472 4164 3473
rect 4158 3468 4159 3472
rect 4163 3468 4164 3472
rect 4158 3467 4164 3468
rect 4294 3472 4300 3473
rect 4294 3468 4295 3472
rect 4299 3468 4300 3472
rect 4294 3467 4300 3468
rect 4430 3472 4436 3473
rect 4430 3468 4431 3472
rect 4435 3468 4436 3472
rect 4430 3467 4436 3468
rect 4566 3472 4572 3473
rect 4566 3468 4567 3472
rect 4571 3468 4572 3472
rect 4566 3467 4572 3468
rect 4726 3472 4732 3473
rect 4726 3468 4727 3472
rect 4731 3468 4732 3472
rect 4726 3467 4732 3468
rect 4918 3472 4924 3473
rect 4918 3468 4919 3472
rect 4923 3468 4924 3472
rect 4918 3467 4924 3468
rect 5126 3472 5132 3473
rect 5126 3468 5127 3472
rect 5131 3468 5132 3472
rect 5126 3467 5132 3468
rect 5342 3472 5348 3473
rect 5342 3468 5343 3472
rect 5347 3468 5348 3472
rect 5342 3467 5348 3468
rect 5542 3472 5548 3473
rect 5542 3468 5543 3472
rect 5547 3468 5548 3472
rect 5542 3467 5548 3468
rect 5662 3471 5668 3472
rect 5662 3467 5663 3471
rect 5667 3467 5668 3471
rect 3838 3466 3844 3467
rect 3840 3435 3842 3466
rect 3888 3435 3890 3467
rect 4024 3435 4026 3467
rect 4160 3435 4162 3467
rect 4296 3435 4298 3467
rect 4432 3435 4434 3467
rect 4568 3435 4570 3467
rect 4728 3435 4730 3467
rect 4920 3435 4922 3467
rect 5128 3435 5130 3467
rect 5344 3435 5346 3467
rect 5544 3435 5546 3467
rect 5662 3466 5668 3467
rect 5664 3435 5666 3466
rect 3839 3434 3843 3435
rect 3839 3429 3843 3430
rect 3887 3434 3891 3435
rect 3887 3429 3891 3430
rect 4023 3434 4027 3435
rect 4023 3429 4027 3430
rect 4159 3434 4163 3435
rect 4159 3429 4163 3430
rect 4295 3434 4299 3435
rect 4295 3429 4299 3430
rect 4431 3434 4435 3435
rect 4431 3429 4435 3430
rect 4567 3434 4571 3435
rect 4567 3429 4571 3430
rect 4583 3434 4587 3435
rect 4583 3429 4587 3430
rect 4727 3434 4731 3435
rect 4727 3429 4731 3430
rect 4759 3434 4763 3435
rect 4759 3429 4763 3430
rect 4919 3434 4923 3435
rect 4919 3429 4923 3430
rect 4951 3434 4955 3435
rect 4951 3429 4955 3430
rect 5127 3434 5131 3435
rect 5127 3429 5131 3430
rect 5151 3434 5155 3435
rect 5151 3429 5155 3430
rect 5343 3434 5347 3435
rect 5343 3429 5347 3430
rect 5359 3434 5363 3435
rect 5359 3429 5363 3430
rect 5543 3434 5547 3435
rect 5543 3429 5547 3430
rect 5663 3434 5667 3435
rect 5663 3429 5667 3430
rect 1975 3418 1979 3419
rect 1975 3413 1979 3414
rect 2191 3418 2195 3419
rect 2191 3413 2195 3414
rect 2231 3418 2235 3419
rect 2231 3413 2235 3414
rect 2327 3418 2331 3419
rect 2327 3413 2331 3414
rect 2463 3418 2467 3419
rect 2463 3413 2467 3414
rect 2583 3418 2587 3419
rect 2583 3413 2587 3414
rect 2599 3418 2603 3419
rect 2599 3413 2603 3414
rect 2951 3418 2955 3419
rect 2951 3413 2955 3414
rect 3327 3418 3331 3419
rect 3327 3413 3331 3414
rect 3679 3418 3683 3419
rect 3679 3413 3683 3414
rect 3799 3418 3803 3419
rect 3799 3413 3803 3414
rect 1976 3390 1978 3413
rect 1974 3389 1980 3390
rect 2232 3389 2234 3413
rect 2584 3389 2586 3413
rect 2952 3389 2954 3413
rect 3328 3389 3330 3413
rect 3680 3389 3682 3413
rect 3800 3390 3802 3413
rect 3840 3406 3842 3429
rect 3838 3405 3844 3406
rect 3888 3405 3890 3429
rect 4024 3405 4026 3429
rect 4160 3405 4162 3429
rect 4296 3405 4298 3429
rect 4432 3405 4434 3429
rect 4584 3405 4586 3429
rect 4760 3405 4762 3429
rect 4952 3405 4954 3429
rect 5152 3405 5154 3429
rect 5360 3405 5362 3429
rect 5544 3405 5546 3429
rect 5664 3406 5666 3429
rect 5662 3405 5668 3406
rect 3838 3401 3839 3405
rect 3843 3401 3844 3405
rect 3838 3400 3844 3401
rect 3886 3404 3892 3405
rect 3886 3400 3887 3404
rect 3891 3400 3892 3404
rect 3886 3399 3892 3400
rect 4022 3404 4028 3405
rect 4022 3400 4023 3404
rect 4027 3400 4028 3404
rect 4022 3399 4028 3400
rect 4158 3404 4164 3405
rect 4158 3400 4159 3404
rect 4163 3400 4164 3404
rect 4158 3399 4164 3400
rect 4294 3404 4300 3405
rect 4294 3400 4295 3404
rect 4299 3400 4300 3404
rect 4294 3399 4300 3400
rect 4430 3404 4436 3405
rect 4430 3400 4431 3404
rect 4435 3400 4436 3404
rect 4430 3399 4436 3400
rect 4582 3404 4588 3405
rect 4582 3400 4583 3404
rect 4587 3400 4588 3404
rect 4582 3399 4588 3400
rect 4758 3404 4764 3405
rect 4758 3400 4759 3404
rect 4763 3400 4764 3404
rect 4758 3399 4764 3400
rect 4950 3404 4956 3405
rect 4950 3400 4951 3404
rect 4955 3400 4956 3404
rect 4950 3399 4956 3400
rect 5150 3404 5156 3405
rect 5150 3400 5151 3404
rect 5155 3400 5156 3404
rect 5150 3399 5156 3400
rect 5358 3404 5364 3405
rect 5358 3400 5359 3404
rect 5363 3400 5364 3404
rect 5358 3399 5364 3400
rect 5542 3404 5548 3405
rect 5542 3400 5543 3404
rect 5547 3400 5548 3404
rect 5662 3401 5663 3405
rect 5667 3401 5668 3405
rect 5662 3400 5668 3401
rect 5542 3399 5548 3400
rect 3798 3389 3804 3390
rect 3858 3389 3864 3390
rect 111 3386 115 3387
rect 111 3381 115 3382
rect 131 3386 135 3387
rect 131 3381 135 3382
rect 299 3386 303 3387
rect 299 3381 303 3382
rect 307 3386 311 3387
rect 307 3381 311 3382
rect 507 3386 511 3387
rect 507 3381 511 3382
rect 523 3386 527 3387
rect 523 3381 527 3382
rect 731 3386 735 3387
rect 731 3381 735 3382
rect 763 3386 767 3387
rect 763 3381 767 3382
rect 971 3386 975 3387
rect 971 3381 975 3382
rect 1011 3386 1015 3387
rect 1011 3381 1015 3382
rect 1219 3386 1223 3387
rect 1219 3381 1223 3382
rect 1267 3386 1271 3387
rect 1267 3381 1271 3382
rect 1475 3386 1479 3387
rect 1475 3381 1479 3382
rect 1531 3386 1535 3387
rect 1531 3381 1535 3382
rect 1935 3386 1939 3387
rect 1974 3385 1975 3389
rect 1979 3385 1980 3389
rect 1974 3384 1980 3385
rect 2230 3388 2236 3389
rect 2230 3384 2231 3388
rect 2235 3384 2236 3388
rect 2230 3383 2236 3384
rect 2582 3388 2588 3389
rect 2582 3384 2583 3388
rect 2587 3384 2588 3388
rect 2582 3383 2588 3384
rect 2950 3388 2956 3389
rect 2950 3384 2951 3388
rect 2955 3384 2956 3388
rect 2950 3383 2956 3384
rect 3326 3388 3332 3389
rect 3326 3384 3327 3388
rect 3331 3384 3332 3388
rect 3326 3383 3332 3384
rect 3678 3388 3684 3389
rect 3678 3384 3679 3388
rect 3683 3384 3684 3388
rect 3798 3385 3799 3389
rect 3803 3385 3804 3389
rect 3798 3384 3804 3385
rect 3838 3388 3844 3389
rect 3838 3384 3839 3388
rect 3843 3384 3844 3388
rect 3858 3385 3859 3389
rect 3863 3385 3864 3389
rect 3858 3384 3864 3385
rect 3994 3389 4000 3390
rect 3994 3385 3995 3389
rect 3999 3385 4000 3389
rect 3994 3384 4000 3385
rect 4130 3389 4136 3390
rect 4130 3385 4131 3389
rect 4135 3385 4136 3389
rect 4130 3384 4136 3385
rect 4266 3389 4272 3390
rect 4266 3385 4267 3389
rect 4271 3385 4272 3389
rect 4266 3384 4272 3385
rect 4402 3389 4408 3390
rect 4402 3385 4403 3389
rect 4407 3385 4408 3389
rect 4402 3384 4408 3385
rect 4554 3389 4560 3390
rect 4554 3385 4555 3389
rect 4559 3385 4560 3389
rect 4554 3384 4560 3385
rect 4730 3389 4736 3390
rect 4730 3385 4731 3389
rect 4735 3385 4736 3389
rect 4730 3384 4736 3385
rect 4922 3389 4928 3390
rect 4922 3385 4923 3389
rect 4927 3385 4928 3389
rect 4922 3384 4928 3385
rect 5122 3389 5128 3390
rect 5122 3385 5123 3389
rect 5127 3385 5128 3389
rect 5122 3384 5128 3385
rect 5330 3389 5336 3390
rect 5330 3385 5331 3389
rect 5335 3385 5336 3389
rect 5330 3384 5336 3385
rect 5514 3389 5520 3390
rect 5514 3385 5515 3389
rect 5519 3385 5520 3389
rect 5514 3384 5520 3385
rect 5662 3388 5668 3389
rect 5662 3384 5663 3388
rect 5667 3384 5668 3388
rect 3678 3383 3684 3384
rect 3838 3383 3844 3384
rect 1935 3381 1939 3382
rect 112 3321 114 3381
rect 110 3320 116 3321
rect 132 3320 134 3381
rect 300 3320 302 3381
rect 508 3320 510 3381
rect 732 3320 734 3381
rect 972 3320 974 3381
rect 1220 3320 1222 3381
rect 1476 3320 1478 3381
rect 1936 3321 1938 3381
rect 2202 3373 2208 3374
rect 1974 3372 1980 3373
rect 1974 3368 1975 3372
rect 1979 3368 1980 3372
rect 2202 3369 2203 3373
rect 2207 3369 2208 3373
rect 2202 3368 2208 3369
rect 2554 3373 2560 3374
rect 2554 3369 2555 3373
rect 2559 3369 2560 3373
rect 2554 3368 2560 3369
rect 2922 3373 2928 3374
rect 2922 3369 2923 3373
rect 2927 3369 2928 3373
rect 2922 3368 2928 3369
rect 3298 3373 3304 3374
rect 3298 3369 3299 3373
rect 3303 3369 3304 3373
rect 3298 3368 3304 3369
rect 3650 3373 3656 3374
rect 3650 3369 3651 3373
rect 3655 3369 3656 3373
rect 3650 3368 3656 3369
rect 3798 3372 3804 3373
rect 3798 3368 3799 3372
rect 3803 3368 3804 3372
rect 1974 3367 1980 3368
rect 1934 3320 1940 3321
rect 110 3316 111 3320
rect 115 3316 116 3320
rect 110 3315 116 3316
rect 130 3319 136 3320
rect 130 3315 131 3319
rect 135 3315 136 3319
rect 130 3314 136 3315
rect 298 3319 304 3320
rect 298 3315 299 3319
rect 303 3315 304 3319
rect 298 3314 304 3315
rect 506 3319 512 3320
rect 506 3315 507 3319
rect 511 3315 512 3319
rect 506 3314 512 3315
rect 730 3319 736 3320
rect 730 3315 731 3319
rect 735 3315 736 3319
rect 730 3314 736 3315
rect 970 3319 976 3320
rect 970 3315 971 3319
rect 975 3315 976 3319
rect 970 3314 976 3315
rect 1218 3319 1224 3320
rect 1218 3315 1219 3319
rect 1223 3315 1224 3319
rect 1218 3314 1224 3315
rect 1474 3319 1480 3320
rect 1474 3315 1475 3319
rect 1479 3315 1480 3319
rect 1934 3316 1935 3320
rect 1939 3316 1940 3320
rect 1934 3315 1940 3316
rect 1474 3314 1480 3315
rect 1976 3307 1978 3367
rect 2204 3307 2206 3368
rect 2556 3307 2558 3368
rect 2924 3307 2926 3368
rect 3300 3307 3302 3368
rect 3652 3307 3654 3368
rect 3798 3367 3804 3368
rect 3800 3307 3802 3367
rect 3840 3307 3842 3383
rect 3860 3307 3862 3384
rect 3996 3307 3998 3384
rect 4132 3307 4134 3384
rect 4268 3307 4270 3384
rect 4404 3307 4406 3384
rect 4556 3307 4558 3384
rect 4732 3307 4734 3384
rect 4924 3307 4926 3384
rect 5124 3307 5126 3384
rect 5332 3307 5334 3384
rect 5516 3307 5518 3384
rect 5662 3383 5668 3384
rect 5664 3307 5666 3383
rect 1975 3306 1979 3307
rect 158 3304 164 3305
rect 110 3303 116 3304
rect 110 3299 111 3303
rect 115 3299 116 3303
rect 158 3300 159 3304
rect 163 3300 164 3304
rect 158 3299 164 3300
rect 326 3304 332 3305
rect 326 3300 327 3304
rect 331 3300 332 3304
rect 326 3299 332 3300
rect 534 3304 540 3305
rect 534 3300 535 3304
rect 539 3300 540 3304
rect 534 3299 540 3300
rect 758 3304 764 3305
rect 758 3300 759 3304
rect 763 3300 764 3304
rect 758 3299 764 3300
rect 998 3304 1004 3305
rect 998 3300 999 3304
rect 1003 3300 1004 3304
rect 998 3299 1004 3300
rect 1246 3304 1252 3305
rect 1246 3300 1247 3304
rect 1251 3300 1252 3304
rect 1246 3299 1252 3300
rect 1502 3304 1508 3305
rect 1502 3300 1503 3304
rect 1507 3300 1508 3304
rect 1502 3299 1508 3300
rect 1934 3303 1940 3304
rect 1934 3299 1935 3303
rect 1939 3299 1940 3303
rect 1975 3301 1979 3302
rect 2203 3306 2207 3307
rect 2203 3301 2207 3302
rect 2251 3306 2255 3307
rect 2251 3301 2255 3302
rect 2475 3306 2479 3307
rect 2475 3301 2479 3302
rect 2555 3306 2559 3307
rect 2555 3301 2559 3302
rect 2691 3306 2695 3307
rect 2691 3301 2695 3302
rect 2899 3306 2903 3307
rect 2899 3301 2903 3302
rect 2923 3306 2927 3307
rect 2923 3301 2927 3302
rect 3099 3306 3103 3307
rect 3099 3301 3103 3302
rect 3291 3306 3295 3307
rect 3291 3301 3295 3302
rect 3299 3306 3303 3307
rect 3299 3301 3303 3302
rect 3483 3306 3487 3307
rect 3483 3301 3487 3302
rect 3651 3306 3655 3307
rect 3651 3301 3655 3302
rect 3799 3306 3803 3307
rect 3799 3301 3803 3302
rect 3839 3306 3843 3307
rect 3839 3301 3843 3302
rect 3859 3306 3863 3307
rect 3859 3301 3863 3302
rect 3995 3306 3999 3307
rect 3995 3301 3999 3302
rect 4131 3306 4135 3307
rect 4131 3301 4135 3302
rect 4267 3306 4271 3307
rect 4267 3301 4271 3302
rect 4403 3306 4407 3307
rect 4403 3301 4407 3302
rect 4555 3306 4559 3307
rect 4555 3301 4559 3302
rect 4691 3306 4695 3307
rect 4691 3301 4695 3302
rect 4731 3306 4735 3307
rect 4731 3301 4735 3302
rect 4827 3306 4831 3307
rect 4827 3301 4831 3302
rect 4923 3306 4927 3307
rect 4923 3301 4927 3302
rect 4963 3306 4967 3307
rect 4963 3301 4967 3302
rect 5099 3306 5103 3307
rect 5099 3301 5103 3302
rect 5123 3306 5127 3307
rect 5123 3301 5127 3302
rect 5235 3306 5239 3307
rect 5235 3301 5239 3302
rect 5331 3306 5335 3307
rect 5331 3301 5335 3302
rect 5515 3306 5519 3307
rect 5515 3301 5519 3302
rect 5663 3306 5667 3307
rect 5663 3301 5667 3302
rect 110 3298 116 3299
rect 112 3271 114 3298
rect 160 3271 162 3299
rect 328 3271 330 3299
rect 536 3271 538 3299
rect 760 3271 762 3299
rect 1000 3271 1002 3299
rect 1248 3271 1250 3299
rect 1504 3271 1506 3299
rect 1934 3298 1940 3299
rect 1936 3271 1938 3298
rect 111 3270 115 3271
rect 111 3265 115 3266
rect 159 3270 163 3271
rect 159 3265 163 3266
rect 239 3270 243 3271
rect 239 3265 243 3266
rect 327 3270 331 3271
rect 327 3265 331 3266
rect 463 3270 467 3271
rect 463 3265 467 3266
rect 535 3270 539 3271
rect 535 3265 539 3266
rect 703 3270 707 3271
rect 703 3265 707 3266
rect 759 3270 763 3271
rect 759 3265 763 3266
rect 951 3270 955 3271
rect 951 3265 955 3266
rect 999 3270 1003 3271
rect 999 3265 1003 3266
rect 1199 3270 1203 3271
rect 1199 3265 1203 3266
rect 1247 3270 1251 3271
rect 1247 3265 1251 3266
rect 1455 3270 1459 3271
rect 1455 3265 1459 3266
rect 1503 3270 1507 3271
rect 1503 3265 1507 3266
rect 1935 3270 1939 3271
rect 1935 3265 1939 3266
rect 112 3242 114 3265
rect 110 3241 116 3242
rect 240 3241 242 3265
rect 464 3241 466 3265
rect 704 3241 706 3265
rect 952 3241 954 3265
rect 1200 3241 1202 3265
rect 1456 3241 1458 3265
rect 1936 3242 1938 3265
rect 1934 3241 1940 3242
rect 1976 3241 1978 3301
rect 110 3237 111 3241
rect 115 3237 116 3241
rect 110 3236 116 3237
rect 238 3240 244 3241
rect 238 3236 239 3240
rect 243 3236 244 3240
rect 238 3235 244 3236
rect 462 3240 468 3241
rect 462 3236 463 3240
rect 467 3236 468 3240
rect 462 3235 468 3236
rect 702 3240 708 3241
rect 702 3236 703 3240
rect 707 3236 708 3240
rect 702 3235 708 3236
rect 950 3240 956 3241
rect 950 3236 951 3240
rect 955 3236 956 3240
rect 950 3235 956 3236
rect 1198 3240 1204 3241
rect 1198 3236 1199 3240
rect 1203 3236 1204 3240
rect 1198 3235 1204 3236
rect 1454 3240 1460 3241
rect 1454 3236 1455 3240
rect 1459 3236 1460 3240
rect 1934 3237 1935 3241
rect 1939 3237 1940 3241
rect 1934 3236 1940 3237
rect 1974 3240 1980 3241
rect 2252 3240 2254 3301
rect 2476 3240 2478 3301
rect 2692 3240 2694 3301
rect 2900 3240 2902 3301
rect 3100 3240 3102 3301
rect 3292 3240 3294 3301
rect 3484 3240 3486 3301
rect 3652 3240 3654 3301
rect 3800 3241 3802 3301
rect 3840 3241 3842 3301
rect 3798 3240 3804 3241
rect 1974 3236 1975 3240
rect 1979 3236 1980 3240
rect 1454 3235 1460 3236
rect 1974 3235 1980 3236
rect 2250 3239 2256 3240
rect 2250 3235 2251 3239
rect 2255 3235 2256 3239
rect 2250 3234 2256 3235
rect 2474 3239 2480 3240
rect 2474 3235 2475 3239
rect 2479 3235 2480 3239
rect 2474 3234 2480 3235
rect 2690 3239 2696 3240
rect 2690 3235 2691 3239
rect 2695 3235 2696 3239
rect 2690 3234 2696 3235
rect 2898 3239 2904 3240
rect 2898 3235 2899 3239
rect 2903 3235 2904 3239
rect 2898 3234 2904 3235
rect 3098 3239 3104 3240
rect 3098 3235 3099 3239
rect 3103 3235 3104 3239
rect 3098 3234 3104 3235
rect 3290 3239 3296 3240
rect 3290 3235 3291 3239
rect 3295 3235 3296 3239
rect 3290 3234 3296 3235
rect 3482 3239 3488 3240
rect 3482 3235 3483 3239
rect 3487 3235 3488 3239
rect 3482 3234 3488 3235
rect 3650 3239 3656 3240
rect 3650 3235 3651 3239
rect 3655 3235 3656 3239
rect 3798 3236 3799 3240
rect 3803 3236 3804 3240
rect 3798 3235 3804 3236
rect 3838 3240 3844 3241
rect 4692 3240 4694 3301
rect 4828 3240 4830 3301
rect 4964 3240 4966 3301
rect 5100 3240 5102 3301
rect 5236 3240 5238 3301
rect 5664 3241 5666 3301
rect 5662 3240 5668 3241
rect 3838 3236 3839 3240
rect 3843 3236 3844 3240
rect 3838 3235 3844 3236
rect 4690 3239 4696 3240
rect 4690 3235 4691 3239
rect 4695 3235 4696 3239
rect 3650 3234 3656 3235
rect 4690 3234 4696 3235
rect 4826 3239 4832 3240
rect 4826 3235 4827 3239
rect 4831 3235 4832 3239
rect 4826 3234 4832 3235
rect 4962 3239 4968 3240
rect 4962 3235 4963 3239
rect 4967 3235 4968 3239
rect 4962 3234 4968 3235
rect 5098 3239 5104 3240
rect 5098 3235 5099 3239
rect 5103 3235 5104 3239
rect 5098 3234 5104 3235
rect 5234 3239 5240 3240
rect 5234 3235 5235 3239
rect 5239 3235 5240 3239
rect 5662 3236 5663 3240
rect 5667 3236 5668 3240
rect 5662 3235 5668 3236
rect 5234 3234 5240 3235
rect 210 3225 216 3226
rect 110 3224 116 3225
rect 110 3220 111 3224
rect 115 3220 116 3224
rect 210 3221 211 3225
rect 215 3221 216 3225
rect 210 3220 216 3221
rect 434 3225 440 3226
rect 434 3221 435 3225
rect 439 3221 440 3225
rect 434 3220 440 3221
rect 674 3225 680 3226
rect 674 3221 675 3225
rect 679 3221 680 3225
rect 674 3220 680 3221
rect 922 3225 928 3226
rect 922 3221 923 3225
rect 927 3221 928 3225
rect 922 3220 928 3221
rect 1170 3225 1176 3226
rect 1170 3221 1171 3225
rect 1175 3221 1176 3225
rect 1170 3220 1176 3221
rect 1426 3225 1432 3226
rect 1426 3221 1427 3225
rect 1431 3221 1432 3225
rect 1426 3220 1432 3221
rect 1934 3224 1940 3225
rect 2278 3224 2284 3225
rect 1934 3220 1935 3224
rect 1939 3220 1940 3224
rect 110 3219 116 3220
rect 112 3155 114 3219
rect 212 3155 214 3220
rect 436 3155 438 3220
rect 676 3155 678 3220
rect 924 3155 926 3220
rect 1172 3155 1174 3220
rect 1428 3155 1430 3220
rect 1934 3219 1940 3220
rect 1974 3223 1980 3224
rect 1974 3219 1975 3223
rect 1979 3219 1980 3223
rect 2278 3220 2279 3224
rect 2283 3220 2284 3224
rect 2278 3219 2284 3220
rect 2502 3224 2508 3225
rect 2502 3220 2503 3224
rect 2507 3220 2508 3224
rect 2502 3219 2508 3220
rect 2718 3224 2724 3225
rect 2718 3220 2719 3224
rect 2723 3220 2724 3224
rect 2718 3219 2724 3220
rect 2926 3224 2932 3225
rect 2926 3220 2927 3224
rect 2931 3220 2932 3224
rect 2926 3219 2932 3220
rect 3126 3224 3132 3225
rect 3126 3220 3127 3224
rect 3131 3220 3132 3224
rect 3126 3219 3132 3220
rect 3318 3224 3324 3225
rect 3318 3220 3319 3224
rect 3323 3220 3324 3224
rect 3318 3219 3324 3220
rect 3510 3224 3516 3225
rect 3510 3220 3511 3224
rect 3515 3220 3516 3224
rect 3510 3219 3516 3220
rect 3678 3224 3684 3225
rect 4718 3224 4724 3225
rect 3678 3220 3679 3224
rect 3683 3220 3684 3224
rect 3678 3219 3684 3220
rect 3798 3223 3804 3224
rect 3798 3219 3799 3223
rect 3803 3219 3804 3223
rect 1936 3155 1938 3219
rect 1974 3218 1980 3219
rect 1976 3187 1978 3218
rect 2280 3187 2282 3219
rect 2504 3187 2506 3219
rect 2720 3187 2722 3219
rect 2928 3187 2930 3219
rect 3128 3187 3130 3219
rect 3320 3187 3322 3219
rect 3512 3187 3514 3219
rect 3680 3187 3682 3219
rect 3798 3218 3804 3219
rect 3838 3223 3844 3224
rect 3838 3219 3839 3223
rect 3843 3219 3844 3223
rect 4718 3220 4719 3224
rect 4723 3220 4724 3224
rect 4718 3219 4724 3220
rect 4854 3224 4860 3225
rect 4854 3220 4855 3224
rect 4859 3220 4860 3224
rect 4854 3219 4860 3220
rect 4990 3224 4996 3225
rect 4990 3220 4991 3224
rect 4995 3220 4996 3224
rect 4990 3219 4996 3220
rect 5126 3224 5132 3225
rect 5126 3220 5127 3224
rect 5131 3220 5132 3224
rect 5126 3219 5132 3220
rect 5262 3224 5268 3225
rect 5262 3220 5263 3224
rect 5267 3220 5268 3224
rect 5262 3219 5268 3220
rect 5662 3223 5668 3224
rect 5662 3219 5663 3223
rect 5667 3219 5668 3223
rect 3838 3218 3844 3219
rect 3800 3187 3802 3218
rect 3840 3187 3842 3218
rect 4720 3187 4722 3219
rect 4856 3187 4858 3219
rect 4992 3187 4994 3219
rect 5128 3187 5130 3219
rect 5264 3187 5266 3219
rect 5662 3218 5668 3219
rect 5664 3187 5666 3218
rect 1975 3186 1979 3187
rect 1975 3181 1979 3182
rect 2095 3186 2099 3187
rect 2095 3181 2099 3182
rect 2279 3186 2283 3187
rect 2279 3181 2283 3182
rect 2295 3186 2299 3187
rect 2295 3181 2299 3182
rect 2487 3186 2491 3187
rect 2487 3181 2491 3182
rect 2503 3186 2507 3187
rect 2503 3181 2507 3182
rect 2679 3186 2683 3187
rect 2679 3181 2683 3182
rect 2719 3186 2723 3187
rect 2719 3181 2723 3182
rect 2871 3186 2875 3187
rect 2871 3181 2875 3182
rect 2927 3186 2931 3187
rect 2927 3181 2931 3182
rect 3055 3186 3059 3187
rect 3055 3181 3059 3182
rect 3127 3186 3131 3187
rect 3127 3181 3131 3182
rect 3231 3186 3235 3187
rect 3231 3181 3235 3182
rect 3319 3186 3323 3187
rect 3319 3181 3323 3182
rect 3415 3186 3419 3187
rect 3415 3181 3419 3182
rect 3511 3186 3515 3187
rect 3511 3181 3515 3182
rect 3599 3186 3603 3187
rect 3599 3181 3603 3182
rect 3679 3186 3683 3187
rect 3679 3181 3683 3182
rect 3799 3186 3803 3187
rect 3799 3181 3803 3182
rect 3839 3186 3843 3187
rect 3839 3181 3843 3182
rect 4719 3186 4723 3187
rect 4719 3181 4723 3182
rect 4855 3186 4859 3187
rect 4855 3181 4859 3182
rect 4863 3186 4867 3187
rect 4863 3181 4867 3182
rect 4991 3186 4995 3187
rect 4991 3181 4995 3182
rect 4999 3186 5003 3187
rect 4999 3181 5003 3182
rect 5127 3186 5131 3187
rect 5127 3181 5131 3182
rect 5135 3186 5139 3187
rect 5135 3181 5139 3182
rect 5263 3186 5267 3187
rect 5263 3181 5267 3182
rect 5271 3186 5275 3187
rect 5271 3181 5275 3182
rect 5407 3186 5411 3187
rect 5407 3181 5411 3182
rect 5543 3186 5547 3187
rect 5543 3181 5547 3182
rect 5663 3186 5667 3187
rect 5663 3181 5667 3182
rect 1976 3158 1978 3181
rect 1974 3157 1980 3158
rect 2096 3157 2098 3181
rect 2296 3157 2298 3181
rect 2488 3157 2490 3181
rect 2680 3157 2682 3181
rect 2872 3157 2874 3181
rect 3056 3157 3058 3181
rect 3232 3157 3234 3181
rect 3416 3157 3418 3181
rect 3600 3157 3602 3181
rect 3800 3158 3802 3181
rect 3840 3158 3842 3181
rect 3798 3157 3804 3158
rect 111 3154 115 3155
rect 111 3149 115 3150
rect 211 3154 215 3155
rect 211 3149 215 3150
rect 379 3154 383 3155
rect 379 3149 383 3150
rect 435 3154 439 3155
rect 435 3149 439 3150
rect 563 3154 567 3155
rect 563 3149 567 3150
rect 675 3154 679 3155
rect 675 3149 679 3150
rect 755 3154 759 3155
rect 755 3149 759 3150
rect 923 3154 927 3155
rect 923 3149 927 3150
rect 955 3154 959 3155
rect 955 3149 959 3150
rect 1163 3154 1167 3155
rect 1163 3149 1167 3150
rect 1171 3154 1175 3155
rect 1171 3149 1175 3150
rect 1371 3154 1375 3155
rect 1371 3149 1375 3150
rect 1427 3154 1431 3155
rect 1427 3149 1431 3150
rect 1935 3154 1939 3155
rect 1974 3153 1975 3157
rect 1979 3153 1980 3157
rect 1974 3152 1980 3153
rect 2094 3156 2100 3157
rect 2094 3152 2095 3156
rect 2099 3152 2100 3156
rect 2094 3151 2100 3152
rect 2294 3156 2300 3157
rect 2294 3152 2295 3156
rect 2299 3152 2300 3156
rect 2294 3151 2300 3152
rect 2486 3156 2492 3157
rect 2486 3152 2487 3156
rect 2491 3152 2492 3156
rect 2486 3151 2492 3152
rect 2678 3156 2684 3157
rect 2678 3152 2679 3156
rect 2683 3152 2684 3156
rect 2678 3151 2684 3152
rect 2870 3156 2876 3157
rect 2870 3152 2871 3156
rect 2875 3152 2876 3156
rect 2870 3151 2876 3152
rect 3054 3156 3060 3157
rect 3054 3152 3055 3156
rect 3059 3152 3060 3156
rect 3054 3151 3060 3152
rect 3230 3156 3236 3157
rect 3230 3152 3231 3156
rect 3235 3152 3236 3156
rect 3230 3151 3236 3152
rect 3414 3156 3420 3157
rect 3414 3152 3415 3156
rect 3419 3152 3420 3156
rect 3414 3151 3420 3152
rect 3598 3156 3604 3157
rect 3598 3152 3599 3156
rect 3603 3152 3604 3156
rect 3798 3153 3799 3157
rect 3803 3153 3804 3157
rect 3798 3152 3804 3153
rect 3838 3157 3844 3158
rect 4864 3157 4866 3181
rect 5000 3157 5002 3181
rect 5136 3157 5138 3181
rect 5272 3157 5274 3181
rect 5408 3157 5410 3181
rect 5544 3157 5546 3181
rect 5664 3158 5666 3181
rect 5662 3157 5668 3158
rect 3838 3153 3839 3157
rect 3843 3153 3844 3157
rect 3838 3152 3844 3153
rect 4862 3156 4868 3157
rect 4862 3152 4863 3156
rect 4867 3152 4868 3156
rect 3598 3151 3604 3152
rect 4862 3151 4868 3152
rect 4998 3156 5004 3157
rect 4998 3152 4999 3156
rect 5003 3152 5004 3156
rect 4998 3151 5004 3152
rect 5134 3156 5140 3157
rect 5134 3152 5135 3156
rect 5139 3152 5140 3156
rect 5134 3151 5140 3152
rect 5270 3156 5276 3157
rect 5270 3152 5271 3156
rect 5275 3152 5276 3156
rect 5270 3151 5276 3152
rect 5406 3156 5412 3157
rect 5406 3152 5407 3156
rect 5411 3152 5412 3156
rect 5406 3151 5412 3152
rect 5542 3156 5548 3157
rect 5542 3152 5543 3156
rect 5547 3152 5548 3156
rect 5662 3153 5663 3157
rect 5667 3153 5668 3157
rect 5662 3152 5668 3153
rect 5542 3151 5548 3152
rect 1935 3149 1939 3150
rect 112 3089 114 3149
rect 110 3088 116 3089
rect 380 3088 382 3149
rect 564 3088 566 3149
rect 756 3088 758 3149
rect 956 3088 958 3149
rect 1164 3088 1166 3149
rect 1372 3088 1374 3149
rect 1936 3089 1938 3149
rect 2066 3141 2072 3142
rect 1974 3140 1980 3141
rect 1974 3136 1975 3140
rect 1979 3136 1980 3140
rect 2066 3137 2067 3141
rect 2071 3137 2072 3141
rect 2066 3136 2072 3137
rect 2266 3141 2272 3142
rect 2266 3137 2267 3141
rect 2271 3137 2272 3141
rect 2266 3136 2272 3137
rect 2458 3141 2464 3142
rect 2458 3137 2459 3141
rect 2463 3137 2464 3141
rect 2458 3136 2464 3137
rect 2650 3141 2656 3142
rect 2650 3137 2651 3141
rect 2655 3137 2656 3141
rect 2650 3136 2656 3137
rect 2842 3141 2848 3142
rect 2842 3137 2843 3141
rect 2847 3137 2848 3141
rect 2842 3136 2848 3137
rect 3026 3141 3032 3142
rect 3026 3137 3027 3141
rect 3031 3137 3032 3141
rect 3026 3136 3032 3137
rect 3202 3141 3208 3142
rect 3202 3137 3203 3141
rect 3207 3137 3208 3141
rect 3202 3136 3208 3137
rect 3386 3141 3392 3142
rect 3386 3137 3387 3141
rect 3391 3137 3392 3141
rect 3386 3136 3392 3137
rect 3570 3141 3576 3142
rect 4834 3141 4840 3142
rect 3570 3137 3571 3141
rect 3575 3137 3576 3141
rect 3570 3136 3576 3137
rect 3798 3140 3804 3141
rect 3798 3136 3799 3140
rect 3803 3136 3804 3140
rect 1974 3135 1980 3136
rect 1934 3088 1940 3089
rect 110 3084 111 3088
rect 115 3084 116 3088
rect 110 3083 116 3084
rect 378 3087 384 3088
rect 378 3083 379 3087
rect 383 3083 384 3087
rect 378 3082 384 3083
rect 562 3087 568 3088
rect 562 3083 563 3087
rect 567 3083 568 3087
rect 562 3082 568 3083
rect 754 3087 760 3088
rect 754 3083 755 3087
rect 759 3083 760 3087
rect 754 3082 760 3083
rect 954 3087 960 3088
rect 954 3083 955 3087
rect 959 3083 960 3087
rect 954 3082 960 3083
rect 1162 3087 1168 3088
rect 1162 3083 1163 3087
rect 1167 3083 1168 3087
rect 1162 3082 1168 3083
rect 1370 3087 1376 3088
rect 1370 3083 1371 3087
rect 1375 3083 1376 3087
rect 1934 3084 1935 3088
rect 1939 3084 1940 3088
rect 1934 3083 1940 3084
rect 1370 3082 1376 3083
rect 406 3072 412 3073
rect 110 3071 116 3072
rect 110 3067 111 3071
rect 115 3067 116 3071
rect 406 3068 407 3072
rect 411 3068 412 3072
rect 406 3067 412 3068
rect 590 3072 596 3073
rect 590 3068 591 3072
rect 595 3068 596 3072
rect 590 3067 596 3068
rect 782 3072 788 3073
rect 782 3068 783 3072
rect 787 3068 788 3072
rect 782 3067 788 3068
rect 982 3072 988 3073
rect 982 3068 983 3072
rect 987 3068 988 3072
rect 982 3067 988 3068
rect 1190 3072 1196 3073
rect 1190 3068 1191 3072
rect 1195 3068 1196 3072
rect 1190 3067 1196 3068
rect 1398 3072 1404 3073
rect 1398 3068 1399 3072
rect 1403 3068 1404 3072
rect 1398 3067 1404 3068
rect 1934 3071 1940 3072
rect 1934 3067 1935 3071
rect 1939 3067 1940 3071
rect 110 3066 116 3067
rect 112 3027 114 3066
rect 408 3027 410 3067
rect 592 3027 594 3067
rect 784 3027 786 3067
rect 984 3027 986 3067
rect 1192 3027 1194 3067
rect 1400 3027 1402 3067
rect 1934 3066 1940 3067
rect 1936 3027 1938 3066
rect 1976 3063 1978 3135
rect 2068 3063 2070 3136
rect 2268 3063 2270 3136
rect 2460 3063 2462 3136
rect 2652 3063 2654 3136
rect 2844 3063 2846 3136
rect 3028 3063 3030 3136
rect 3204 3063 3206 3136
rect 3388 3063 3390 3136
rect 3572 3063 3574 3136
rect 3798 3135 3804 3136
rect 3838 3140 3844 3141
rect 3838 3136 3839 3140
rect 3843 3136 3844 3140
rect 4834 3137 4835 3141
rect 4839 3137 4840 3141
rect 4834 3136 4840 3137
rect 4970 3141 4976 3142
rect 4970 3137 4971 3141
rect 4975 3137 4976 3141
rect 4970 3136 4976 3137
rect 5106 3141 5112 3142
rect 5106 3137 5107 3141
rect 5111 3137 5112 3141
rect 5106 3136 5112 3137
rect 5242 3141 5248 3142
rect 5242 3137 5243 3141
rect 5247 3137 5248 3141
rect 5242 3136 5248 3137
rect 5378 3141 5384 3142
rect 5378 3137 5379 3141
rect 5383 3137 5384 3141
rect 5378 3136 5384 3137
rect 5514 3141 5520 3142
rect 5514 3137 5515 3141
rect 5519 3137 5520 3141
rect 5514 3136 5520 3137
rect 5662 3140 5668 3141
rect 5662 3136 5663 3140
rect 5667 3136 5668 3140
rect 3838 3135 3844 3136
rect 3800 3063 3802 3135
rect 3840 3063 3842 3135
rect 4836 3063 4838 3136
rect 4972 3063 4974 3136
rect 5108 3063 5110 3136
rect 5244 3063 5246 3136
rect 5380 3063 5382 3136
rect 5516 3063 5518 3136
rect 5662 3135 5668 3136
rect 5664 3063 5666 3135
rect 1975 3062 1979 3063
rect 1975 3057 1979 3058
rect 1995 3062 1999 3063
rect 1995 3057 1999 3058
rect 2067 3062 2071 3063
rect 2067 3057 2071 3058
rect 2131 3062 2135 3063
rect 2131 3057 2135 3058
rect 2267 3062 2271 3063
rect 2267 3057 2271 3058
rect 2403 3062 2407 3063
rect 2403 3057 2407 3058
rect 2459 3062 2463 3063
rect 2459 3057 2463 3058
rect 2539 3062 2543 3063
rect 2539 3057 2543 3058
rect 2651 3062 2655 3063
rect 2651 3057 2655 3058
rect 2683 3062 2687 3063
rect 2683 3057 2687 3058
rect 2835 3062 2839 3063
rect 2835 3057 2839 3058
rect 2843 3062 2847 3063
rect 2843 3057 2847 3058
rect 2987 3062 2991 3063
rect 2987 3057 2991 3058
rect 3027 3062 3031 3063
rect 3027 3057 3031 3058
rect 3139 3062 3143 3063
rect 3139 3057 3143 3058
rect 3203 3062 3207 3063
rect 3203 3057 3207 3058
rect 3291 3062 3295 3063
rect 3291 3057 3295 3058
rect 3387 3062 3391 3063
rect 3387 3057 3391 3058
rect 3571 3062 3575 3063
rect 3571 3057 3575 3058
rect 3799 3062 3803 3063
rect 3799 3057 3803 3058
rect 3839 3062 3843 3063
rect 3839 3057 3843 3058
rect 4483 3062 4487 3063
rect 4483 3057 4487 3058
rect 4635 3062 4639 3063
rect 4635 3057 4639 3058
rect 4803 3062 4807 3063
rect 4803 3057 4807 3058
rect 4835 3062 4839 3063
rect 4835 3057 4839 3058
rect 4971 3062 4975 3063
rect 4971 3057 4975 3058
rect 4979 3062 4983 3063
rect 4979 3057 4983 3058
rect 5107 3062 5111 3063
rect 5107 3057 5111 3058
rect 5163 3062 5167 3063
rect 5163 3057 5167 3058
rect 5243 3062 5247 3063
rect 5243 3057 5247 3058
rect 5347 3062 5351 3063
rect 5347 3057 5351 3058
rect 5379 3062 5383 3063
rect 5379 3057 5383 3058
rect 5515 3062 5519 3063
rect 5515 3057 5519 3058
rect 5663 3062 5667 3063
rect 5663 3057 5667 3058
rect 111 3026 115 3027
rect 111 3021 115 3022
rect 407 3026 411 3027
rect 407 3021 411 3022
rect 575 3026 579 3027
rect 575 3021 579 3022
rect 591 3026 595 3027
rect 591 3021 595 3022
rect 783 3026 787 3027
rect 783 3021 787 3022
rect 799 3026 803 3027
rect 799 3021 803 3022
rect 983 3026 987 3027
rect 983 3021 987 3022
rect 1047 3026 1051 3027
rect 1047 3021 1051 3022
rect 1191 3026 1195 3027
rect 1191 3021 1195 3022
rect 1303 3026 1307 3027
rect 1303 3021 1307 3022
rect 1399 3026 1403 3027
rect 1399 3021 1403 3022
rect 1567 3026 1571 3027
rect 1567 3021 1571 3022
rect 1815 3026 1819 3027
rect 1815 3021 1819 3022
rect 1935 3026 1939 3027
rect 1935 3021 1939 3022
rect 112 2998 114 3021
rect 110 2997 116 2998
rect 576 2997 578 3021
rect 800 2997 802 3021
rect 1048 2997 1050 3021
rect 1304 2997 1306 3021
rect 1568 2997 1570 3021
rect 1816 2997 1818 3021
rect 1936 2998 1938 3021
rect 1934 2997 1940 2998
rect 1976 2997 1978 3057
rect 110 2993 111 2997
rect 115 2993 116 2997
rect 110 2992 116 2993
rect 574 2996 580 2997
rect 574 2992 575 2996
rect 579 2992 580 2996
rect 574 2991 580 2992
rect 798 2996 804 2997
rect 798 2992 799 2996
rect 803 2992 804 2996
rect 798 2991 804 2992
rect 1046 2996 1052 2997
rect 1046 2992 1047 2996
rect 1051 2992 1052 2996
rect 1046 2991 1052 2992
rect 1302 2996 1308 2997
rect 1302 2992 1303 2996
rect 1307 2992 1308 2996
rect 1302 2991 1308 2992
rect 1566 2996 1572 2997
rect 1566 2992 1567 2996
rect 1571 2992 1572 2996
rect 1566 2991 1572 2992
rect 1814 2996 1820 2997
rect 1814 2992 1815 2996
rect 1819 2992 1820 2996
rect 1934 2993 1935 2997
rect 1939 2993 1940 2997
rect 1934 2992 1940 2993
rect 1974 2996 1980 2997
rect 1996 2996 1998 3057
rect 2132 2996 2134 3057
rect 2268 2996 2270 3057
rect 2404 2996 2406 3057
rect 2540 2996 2542 3057
rect 2684 2996 2686 3057
rect 2836 2996 2838 3057
rect 2988 2996 2990 3057
rect 3140 2996 3142 3057
rect 3292 2996 3294 3057
rect 3800 2997 3802 3057
rect 3840 2997 3842 3057
rect 3798 2996 3804 2997
rect 1974 2992 1975 2996
rect 1979 2992 1980 2996
rect 1814 2991 1820 2992
rect 1974 2991 1980 2992
rect 1994 2995 2000 2996
rect 1994 2991 1995 2995
rect 1999 2991 2000 2995
rect 1994 2990 2000 2991
rect 2130 2995 2136 2996
rect 2130 2991 2131 2995
rect 2135 2991 2136 2995
rect 2130 2990 2136 2991
rect 2266 2995 2272 2996
rect 2266 2991 2267 2995
rect 2271 2991 2272 2995
rect 2266 2990 2272 2991
rect 2402 2995 2408 2996
rect 2402 2991 2403 2995
rect 2407 2991 2408 2995
rect 2402 2990 2408 2991
rect 2538 2995 2544 2996
rect 2538 2991 2539 2995
rect 2543 2991 2544 2995
rect 2538 2990 2544 2991
rect 2682 2995 2688 2996
rect 2682 2991 2683 2995
rect 2687 2991 2688 2995
rect 2682 2990 2688 2991
rect 2834 2995 2840 2996
rect 2834 2991 2835 2995
rect 2839 2991 2840 2995
rect 2834 2990 2840 2991
rect 2986 2995 2992 2996
rect 2986 2991 2987 2995
rect 2991 2991 2992 2995
rect 2986 2990 2992 2991
rect 3138 2995 3144 2996
rect 3138 2991 3139 2995
rect 3143 2991 3144 2995
rect 3138 2990 3144 2991
rect 3290 2995 3296 2996
rect 3290 2991 3291 2995
rect 3295 2991 3296 2995
rect 3798 2992 3799 2996
rect 3803 2992 3804 2996
rect 3798 2991 3804 2992
rect 3838 2996 3844 2997
rect 4484 2996 4486 3057
rect 4636 2996 4638 3057
rect 4804 2996 4806 3057
rect 4980 2996 4982 3057
rect 5164 2996 5166 3057
rect 5348 2996 5350 3057
rect 5516 2996 5518 3057
rect 5664 2997 5666 3057
rect 5662 2996 5668 2997
rect 3838 2992 3839 2996
rect 3843 2992 3844 2996
rect 3838 2991 3844 2992
rect 4482 2995 4488 2996
rect 4482 2991 4483 2995
rect 4487 2991 4488 2995
rect 3290 2990 3296 2991
rect 4482 2990 4488 2991
rect 4634 2995 4640 2996
rect 4634 2991 4635 2995
rect 4639 2991 4640 2995
rect 4634 2990 4640 2991
rect 4802 2995 4808 2996
rect 4802 2991 4803 2995
rect 4807 2991 4808 2995
rect 4802 2990 4808 2991
rect 4978 2995 4984 2996
rect 4978 2991 4979 2995
rect 4983 2991 4984 2995
rect 4978 2990 4984 2991
rect 5162 2995 5168 2996
rect 5162 2991 5163 2995
rect 5167 2991 5168 2995
rect 5162 2990 5168 2991
rect 5346 2995 5352 2996
rect 5346 2991 5347 2995
rect 5351 2991 5352 2995
rect 5346 2990 5352 2991
rect 5514 2995 5520 2996
rect 5514 2991 5515 2995
rect 5519 2991 5520 2995
rect 5662 2992 5663 2996
rect 5667 2992 5668 2996
rect 5662 2991 5668 2992
rect 5514 2990 5520 2991
rect 546 2981 552 2982
rect 110 2980 116 2981
rect 110 2976 111 2980
rect 115 2976 116 2980
rect 546 2977 547 2981
rect 551 2977 552 2981
rect 546 2976 552 2977
rect 770 2981 776 2982
rect 770 2977 771 2981
rect 775 2977 776 2981
rect 770 2976 776 2977
rect 1018 2981 1024 2982
rect 1018 2977 1019 2981
rect 1023 2977 1024 2981
rect 1018 2976 1024 2977
rect 1274 2981 1280 2982
rect 1274 2977 1275 2981
rect 1279 2977 1280 2981
rect 1274 2976 1280 2977
rect 1538 2981 1544 2982
rect 1538 2977 1539 2981
rect 1543 2977 1544 2981
rect 1538 2976 1544 2977
rect 1786 2981 1792 2982
rect 1786 2977 1787 2981
rect 1791 2977 1792 2981
rect 1786 2976 1792 2977
rect 1934 2980 1940 2981
rect 2022 2980 2028 2981
rect 1934 2976 1935 2980
rect 1939 2976 1940 2980
rect 110 2975 116 2976
rect 112 2907 114 2975
rect 548 2907 550 2976
rect 772 2907 774 2976
rect 1020 2907 1022 2976
rect 1276 2907 1278 2976
rect 1540 2907 1542 2976
rect 1788 2907 1790 2976
rect 1934 2975 1940 2976
rect 1974 2979 1980 2980
rect 1974 2975 1975 2979
rect 1979 2975 1980 2979
rect 2022 2976 2023 2980
rect 2027 2976 2028 2980
rect 2022 2975 2028 2976
rect 2158 2980 2164 2981
rect 2158 2976 2159 2980
rect 2163 2976 2164 2980
rect 2158 2975 2164 2976
rect 2294 2980 2300 2981
rect 2294 2976 2295 2980
rect 2299 2976 2300 2980
rect 2294 2975 2300 2976
rect 2430 2980 2436 2981
rect 2430 2976 2431 2980
rect 2435 2976 2436 2980
rect 2430 2975 2436 2976
rect 2566 2980 2572 2981
rect 2566 2976 2567 2980
rect 2571 2976 2572 2980
rect 2566 2975 2572 2976
rect 2710 2980 2716 2981
rect 2710 2976 2711 2980
rect 2715 2976 2716 2980
rect 2710 2975 2716 2976
rect 2862 2980 2868 2981
rect 2862 2976 2863 2980
rect 2867 2976 2868 2980
rect 2862 2975 2868 2976
rect 3014 2980 3020 2981
rect 3014 2976 3015 2980
rect 3019 2976 3020 2980
rect 3014 2975 3020 2976
rect 3166 2980 3172 2981
rect 3166 2976 3167 2980
rect 3171 2976 3172 2980
rect 3166 2975 3172 2976
rect 3318 2980 3324 2981
rect 4510 2980 4516 2981
rect 3318 2976 3319 2980
rect 3323 2976 3324 2980
rect 3318 2975 3324 2976
rect 3798 2979 3804 2980
rect 3798 2975 3799 2979
rect 3803 2975 3804 2979
rect 1936 2907 1938 2975
rect 1974 2974 1980 2975
rect 1976 2951 1978 2974
rect 2024 2951 2026 2975
rect 2160 2951 2162 2975
rect 2296 2951 2298 2975
rect 2432 2951 2434 2975
rect 2568 2951 2570 2975
rect 2712 2951 2714 2975
rect 2864 2951 2866 2975
rect 3016 2951 3018 2975
rect 3168 2951 3170 2975
rect 3320 2951 3322 2975
rect 3798 2974 3804 2975
rect 3838 2979 3844 2980
rect 3838 2975 3839 2979
rect 3843 2975 3844 2979
rect 4510 2976 4511 2980
rect 4515 2976 4516 2980
rect 4510 2975 4516 2976
rect 4662 2980 4668 2981
rect 4662 2976 4663 2980
rect 4667 2976 4668 2980
rect 4662 2975 4668 2976
rect 4830 2980 4836 2981
rect 4830 2976 4831 2980
rect 4835 2976 4836 2980
rect 4830 2975 4836 2976
rect 5006 2980 5012 2981
rect 5006 2976 5007 2980
rect 5011 2976 5012 2980
rect 5006 2975 5012 2976
rect 5190 2980 5196 2981
rect 5190 2976 5191 2980
rect 5195 2976 5196 2980
rect 5190 2975 5196 2976
rect 5374 2980 5380 2981
rect 5374 2976 5375 2980
rect 5379 2976 5380 2980
rect 5374 2975 5380 2976
rect 5542 2980 5548 2981
rect 5542 2976 5543 2980
rect 5547 2976 5548 2980
rect 5542 2975 5548 2976
rect 5662 2979 5668 2980
rect 5662 2975 5663 2979
rect 5667 2975 5668 2979
rect 3838 2974 3844 2975
rect 3800 2951 3802 2974
rect 1975 2950 1979 2951
rect 1975 2945 1979 2946
rect 2023 2950 2027 2951
rect 2023 2945 2027 2946
rect 2159 2950 2163 2951
rect 2159 2945 2163 2946
rect 2295 2950 2299 2951
rect 2295 2945 2299 2946
rect 2431 2950 2435 2951
rect 2431 2945 2435 2946
rect 2567 2950 2571 2951
rect 2567 2945 2571 2946
rect 2591 2950 2595 2951
rect 2591 2945 2595 2946
rect 2711 2950 2715 2951
rect 2711 2945 2715 2946
rect 2863 2950 2867 2951
rect 2863 2945 2867 2946
rect 2887 2950 2891 2951
rect 2887 2945 2891 2946
rect 3015 2950 3019 2951
rect 3015 2945 3019 2946
rect 3167 2950 3171 2951
rect 3167 2945 3171 2946
rect 3183 2950 3187 2951
rect 3183 2945 3187 2946
rect 3319 2950 3323 2951
rect 3319 2945 3323 2946
rect 3799 2950 3803 2951
rect 3799 2945 3803 2946
rect 1976 2922 1978 2945
rect 1974 2921 1980 2922
rect 2024 2921 2026 2945
rect 2296 2921 2298 2945
rect 2592 2921 2594 2945
rect 2888 2921 2890 2945
rect 3184 2921 3186 2945
rect 3800 2922 3802 2945
rect 3840 2927 3842 2974
rect 4512 2927 4514 2975
rect 4664 2927 4666 2975
rect 4832 2927 4834 2975
rect 5008 2927 5010 2975
rect 5192 2927 5194 2975
rect 5376 2927 5378 2975
rect 5544 2927 5546 2975
rect 5662 2974 5668 2975
rect 5664 2927 5666 2974
rect 3839 2926 3843 2927
rect 3798 2921 3804 2922
rect 3839 2921 3843 2922
rect 4047 2926 4051 2927
rect 4047 2921 4051 2922
rect 4295 2926 4299 2927
rect 4295 2921 4299 2922
rect 4511 2926 4515 2927
rect 4511 2921 4515 2922
rect 4583 2926 4587 2927
rect 4583 2921 4587 2922
rect 4663 2926 4667 2927
rect 4663 2921 4667 2922
rect 4831 2926 4835 2927
rect 4831 2921 4835 2922
rect 4895 2926 4899 2927
rect 4895 2921 4899 2922
rect 5007 2926 5011 2927
rect 5007 2921 5011 2922
rect 5191 2926 5195 2927
rect 5191 2921 5195 2922
rect 5231 2926 5235 2927
rect 5231 2921 5235 2922
rect 5375 2926 5379 2927
rect 5375 2921 5379 2922
rect 5543 2926 5547 2927
rect 5543 2921 5547 2922
rect 5663 2926 5667 2927
rect 5663 2921 5667 2922
rect 1974 2917 1975 2921
rect 1979 2917 1980 2921
rect 1974 2916 1980 2917
rect 2022 2920 2028 2921
rect 2022 2916 2023 2920
rect 2027 2916 2028 2920
rect 2022 2915 2028 2916
rect 2294 2920 2300 2921
rect 2294 2916 2295 2920
rect 2299 2916 2300 2920
rect 2294 2915 2300 2916
rect 2590 2920 2596 2921
rect 2590 2916 2591 2920
rect 2595 2916 2596 2920
rect 2590 2915 2596 2916
rect 2886 2920 2892 2921
rect 2886 2916 2887 2920
rect 2891 2916 2892 2920
rect 2886 2915 2892 2916
rect 3182 2920 3188 2921
rect 3182 2916 3183 2920
rect 3187 2916 3188 2920
rect 3798 2917 3799 2921
rect 3803 2917 3804 2921
rect 3798 2916 3804 2917
rect 3182 2915 3188 2916
rect 111 2906 115 2907
rect 111 2901 115 2902
rect 427 2906 431 2907
rect 427 2901 431 2902
rect 547 2906 551 2907
rect 547 2901 551 2902
rect 563 2906 567 2907
rect 563 2901 567 2902
rect 699 2906 703 2907
rect 699 2901 703 2902
rect 771 2906 775 2907
rect 771 2901 775 2902
rect 835 2906 839 2907
rect 835 2901 839 2902
rect 971 2906 975 2907
rect 971 2901 975 2902
rect 1019 2906 1023 2907
rect 1019 2901 1023 2902
rect 1107 2906 1111 2907
rect 1107 2901 1111 2902
rect 1243 2906 1247 2907
rect 1243 2901 1247 2902
rect 1275 2906 1279 2907
rect 1275 2901 1279 2902
rect 1379 2906 1383 2907
rect 1379 2901 1383 2902
rect 1515 2906 1519 2907
rect 1515 2901 1519 2902
rect 1539 2906 1543 2907
rect 1539 2901 1543 2902
rect 1651 2906 1655 2907
rect 1651 2901 1655 2902
rect 1787 2906 1791 2907
rect 1787 2901 1791 2902
rect 1935 2906 1939 2907
rect 1994 2905 2000 2906
rect 1935 2901 1939 2902
rect 1974 2904 1980 2905
rect 112 2841 114 2901
rect 110 2840 116 2841
rect 428 2840 430 2901
rect 564 2840 566 2901
rect 700 2840 702 2901
rect 836 2840 838 2901
rect 972 2840 974 2901
rect 1108 2840 1110 2901
rect 1244 2840 1246 2901
rect 1380 2840 1382 2901
rect 1516 2840 1518 2901
rect 1652 2840 1654 2901
rect 1788 2840 1790 2901
rect 1936 2841 1938 2901
rect 1974 2900 1975 2904
rect 1979 2900 1980 2904
rect 1994 2901 1995 2905
rect 1999 2901 2000 2905
rect 1994 2900 2000 2901
rect 2266 2905 2272 2906
rect 2266 2901 2267 2905
rect 2271 2901 2272 2905
rect 2266 2900 2272 2901
rect 2562 2905 2568 2906
rect 2562 2901 2563 2905
rect 2567 2901 2568 2905
rect 2562 2900 2568 2901
rect 2858 2905 2864 2906
rect 2858 2901 2859 2905
rect 2863 2901 2864 2905
rect 2858 2900 2864 2901
rect 3154 2905 3160 2906
rect 3154 2901 3155 2905
rect 3159 2901 3160 2905
rect 3154 2900 3160 2901
rect 3798 2904 3804 2905
rect 3798 2900 3799 2904
rect 3803 2900 3804 2904
rect 1974 2899 1980 2900
rect 1934 2840 1940 2841
rect 110 2836 111 2840
rect 115 2836 116 2840
rect 110 2835 116 2836
rect 426 2839 432 2840
rect 426 2835 427 2839
rect 431 2835 432 2839
rect 426 2834 432 2835
rect 562 2839 568 2840
rect 562 2835 563 2839
rect 567 2835 568 2839
rect 562 2834 568 2835
rect 698 2839 704 2840
rect 698 2835 699 2839
rect 703 2835 704 2839
rect 698 2834 704 2835
rect 834 2839 840 2840
rect 834 2835 835 2839
rect 839 2835 840 2839
rect 834 2834 840 2835
rect 970 2839 976 2840
rect 970 2835 971 2839
rect 975 2835 976 2839
rect 970 2834 976 2835
rect 1106 2839 1112 2840
rect 1106 2835 1107 2839
rect 1111 2835 1112 2839
rect 1106 2834 1112 2835
rect 1242 2839 1248 2840
rect 1242 2835 1243 2839
rect 1247 2835 1248 2839
rect 1242 2834 1248 2835
rect 1378 2839 1384 2840
rect 1378 2835 1379 2839
rect 1383 2835 1384 2839
rect 1378 2834 1384 2835
rect 1514 2839 1520 2840
rect 1514 2835 1515 2839
rect 1519 2835 1520 2839
rect 1514 2834 1520 2835
rect 1650 2839 1656 2840
rect 1650 2835 1651 2839
rect 1655 2835 1656 2839
rect 1650 2834 1656 2835
rect 1786 2839 1792 2840
rect 1786 2835 1787 2839
rect 1791 2835 1792 2839
rect 1934 2836 1935 2840
rect 1939 2836 1940 2840
rect 1934 2835 1940 2836
rect 1786 2834 1792 2835
rect 454 2824 460 2825
rect 110 2823 116 2824
rect 110 2819 111 2823
rect 115 2819 116 2823
rect 454 2820 455 2824
rect 459 2820 460 2824
rect 454 2819 460 2820
rect 590 2824 596 2825
rect 590 2820 591 2824
rect 595 2820 596 2824
rect 590 2819 596 2820
rect 726 2824 732 2825
rect 726 2820 727 2824
rect 731 2820 732 2824
rect 726 2819 732 2820
rect 862 2824 868 2825
rect 862 2820 863 2824
rect 867 2820 868 2824
rect 862 2819 868 2820
rect 998 2824 1004 2825
rect 998 2820 999 2824
rect 1003 2820 1004 2824
rect 998 2819 1004 2820
rect 1134 2824 1140 2825
rect 1134 2820 1135 2824
rect 1139 2820 1140 2824
rect 1134 2819 1140 2820
rect 1270 2824 1276 2825
rect 1270 2820 1271 2824
rect 1275 2820 1276 2824
rect 1270 2819 1276 2820
rect 1406 2824 1412 2825
rect 1406 2820 1407 2824
rect 1411 2820 1412 2824
rect 1406 2819 1412 2820
rect 1542 2824 1548 2825
rect 1542 2820 1543 2824
rect 1547 2820 1548 2824
rect 1542 2819 1548 2820
rect 1678 2824 1684 2825
rect 1678 2820 1679 2824
rect 1683 2820 1684 2824
rect 1678 2819 1684 2820
rect 1814 2824 1820 2825
rect 1814 2820 1815 2824
rect 1819 2820 1820 2824
rect 1814 2819 1820 2820
rect 1934 2823 1940 2824
rect 1934 2819 1935 2823
rect 1939 2819 1940 2823
rect 110 2818 116 2819
rect 112 2787 114 2818
rect 456 2787 458 2819
rect 592 2787 594 2819
rect 728 2787 730 2819
rect 864 2787 866 2819
rect 1000 2787 1002 2819
rect 1136 2787 1138 2819
rect 1272 2787 1274 2819
rect 1408 2787 1410 2819
rect 1544 2787 1546 2819
rect 1680 2787 1682 2819
rect 1816 2787 1818 2819
rect 1934 2818 1940 2819
rect 1936 2787 1938 2818
rect 111 2786 115 2787
rect 111 2781 115 2782
rect 455 2786 459 2787
rect 455 2781 459 2782
rect 463 2786 467 2787
rect 463 2781 467 2782
rect 591 2786 595 2787
rect 591 2781 595 2782
rect 623 2786 627 2787
rect 623 2781 627 2782
rect 727 2786 731 2787
rect 727 2781 731 2782
rect 783 2786 787 2787
rect 783 2781 787 2782
rect 863 2786 867 2787
rect 863 2781 867 2782
rect 935 2786 939 2787
rect 935 2781 939 2782
rect 999 2786 1003 2787
rect 999 2781 1003 2782
rect 1087 2786 1091 2787
rect 1087 2781 1091 2782
rect 1135 2786 1139 2787
rect 1135 2781 1139 2782
rect 1239 2786 1243 2787
rect 1239 2781 1243 2782
rect 1271 2786 1275 2787
rect 1271 2781 1275 2782
rect 1383 2786 1387 2787
rect 1383 2781 1387 2782
rect 1407 2786 1411 2787
rect 1407 2781 1411 2782
rect 1535 2786 1539 2787
rect 1535 2781 1539 2782
rect 1543 2786 1547 2787
rect 1543 2781 1547 2782
rect 1679 2786 1683 2787
rect 1679 2781 1683 2782
rect 1815 2786 1819 2787
rect 1815 2781 1819 2782
rect 1935 2786 1939 2787
rect 1976 2783 1978 2899
rect 1996 2783 1998 2900
rect 2268 2783 2270 2900
rect 2564 2783 2566 2900
rect 2860 2783 2862 2900
rect 3156 2783 3158 2900
rect 3798 2899 3804 2900
rect 3800 2783 3802 2899
rect 3840 2898 3842 2921
rect 3838 2897 3844 2898
rect 4048 2897 4050 2921
rect 4296 2897 4298 2921
rect 4584 2897 4586 2921
rect 4896 2897 4898 2921
rect 5232 2897 5234 2921
rect 5544 2897 5546 2921
rect 5664 2898 5666 2921
rect 5662 2897 5668 2898
rect 3838 2893 3839 2897
rect 3843 2893 3844 2897
rect 3838 2892 3844 2893
rect 4046 2896 4052 2897
rect 4046 2892 4047 2896
rect 4051 2892 4052 2896
rect 4046 2891 4052 2892
rect 4294 2896 4300 2897
rect 4294 2892 4295 2896
rect 4299 2892 4300 2896
rect 4294 2891 4300 2892
rect 4582 2896 4588 2897
rect 4582 2892 4583 2896
rect 4587 2892 4588 2896
rect 4582 2891 4588 2892
rect 4894 2896 4900 2897
rect 4894 2892 4895 2896
rect 4899 2892 4900 2896
rect 4894 2891 4900 2892
rect 5230 2896 5236 2897
rect 5230 2892 5231 2896
rect 5235 2892 5236 2896
rect 5230 2891 5236 2892
rect 5542 2896 5548 2897
rect 5542 2892 5543 2896
rect 5547 2892 5548 2896
rect 5662 2893 5663 2897
rect 5667 2893 5668 2897
rect 5662 2892 5668 2893
rect 5542 2891 5548 2892
rect 4018 2881 4024 2882
rect 3838 2880 3844 2881
rect 3838 2876 3839 2880
rect 3843 2876 3844 2880
rect 4018 2877 4019 2881
rect 4023 2877 4024 2881
rect 4018 2876 4024 2877
rect 4266 2881 4272 2882
rect 4266 2877 4267 2881
rect 4271 2877 4272 2881
rect 4266 2876 4272 2877
rect 4554 2881 4560 2882
rect 4554 2877 4555 2881
rect 4559 2877 4560 2881
rect 4554 2876 4560 2877
rect 4866 2881 4872 2882
rect 4866 2877 4867 2881
rect 4871 2877 4872 2881
rect 4866 2876 4872 2877
rect 5202 2881 5208 2882
rect 5202 2877 5203 2881
rect 5207 2877 5208 2881
rect 5202 2876 5208 2877
rect 5514 2881 5520 2882
rect 5514 2877 5515 2881
rect 5519 2877 5520 2881
rect 5514 2876 5520 2877
rect 5662 2880 5668 2881
rect 5662 2876 5663 2880
rect 5667 2876 5668 2880
rect 3838 2875 3844 2876
rect 3840 2811 3842 2875
rect 4020 2811 4022 2876
rect 4268 2811 4270 2876
rect 4556 2811 4558 2876
rect 4868 2811 4870 2876
rect 5204 2811 5206 2876
rect 5516 2811 5518 2876
rect 5662 2875 5668 2876
rect 5664 2811 5666 2875
rect 3839 2810 3843 2811
rect 3839 2805 3843 2806
rect 3859 2810 3863 2811
rect 3859 2805 3863 2806
rect 3995 2810 3999 2811
rect 3995 2805 3999 2806
rect 4019 2810 4023 2811
rect 4019 2805 4023 2806
rect 4131 2810 4135 2811
rect 4131 2805 4135 2806
rect 4267 2810 4271 2811
rect 4267 2805 4271 2806
rect 4403 2810 4407 2811
rect 4403 2805 4407 2806
rect 4539 2810 4543 2811
rect 4539 2805 4543 2806
rect 4555 2810 4559 2811
rect 4555 2805 4559 2806
rect 4675 2810 4679 2811
rect 4675 2805 4679 2806
rect 4811 2810 4815 2811
rect 4811 2805 4815 2806
rect 4867 2810 4871 2811
rect 4867 2805 4871 2806
rect 5203 2810 5207 2811
rect 5203 2805 5207 2806
rect 5515 2810 5519 2811
rect 5515 2805 5519 2806
rect 5663 2810 5667 2811
rect 5663 2805 5667 2806
rect 1935 2781 1939 2782
rect 1975 2782 1979 2783
rect 112 2758 114 2781
rect 110 2757 116 2758
rect 464 2757 466 2781
rect 624 2757 626 2781
rect 784 2757 786 2781
rect 936 2757 938 2781
rect 1088 2757 1090 2781
rect 1240 2757 1242 2781
rect 1384 2757 1386 2781
rect 1536 2757 1538 2781
rect 1680 2757 1682 2781
rect 1816 2757 1818 2781
rect 1936 2758 1938 2781
rect 1975 2777 1979 2778
rect 1995 2782 1999 2783
rect 1995 2777 1999 2778
rect 2267 2782 2271 2783
rect 2267 2777 2271 2778
rect 2563 2782 2567 2783
rect 2563 2777 2567 2778
rect 2859 2782 2863 2783
rect 2859 2777 2863 2778
rect 3059 2782 3063 2783
rect 3059 2777 3063 2778
rect 3155 2782 3159 2783
rect 3155 2777 3159 2778
rect 3195 2782 3199 2783
rect 3195 2777 3199 2778
rect 3331 2782 3335 2783
rect 3331 2777 3335 2778
rect 3799 2782 3803 2783
rect 3799 2777 3803 2778
rect 1934 2757 1940 2758
rect 110 2753 111 2757
rect 115 2753 116 2757
rect 110 2752 116 2753
rect 462 2756 468 2757
rect 462 2752 463 2756
rect 467 2752 468 2756
rect 462 2751 468 2752
rect 622 2756 628 2757
rect 622 2752 623 2756
rect 627 2752 628 2756
rect 622 2751 628 2752
rect 782 2756 788 2757
rect 782 2752 783 2756
rect 787 2752 788 2756
rect 782 2751 788 2752
rect 934 2756 940 2757
rect 934 2752 935 2756
rect 939 2752 940 2756
rect 934 2751 940 2752
rect 1086 2756 1092 2757
rect 1086 2752 1087 2756
rect 1091 2752 1092 2756
rect 1086 2751 1092 2752
rect 1238 2756 1244 2757
rect 1238 2752 1239 2756
rect 1243 2752 1244 2756
rect 1238 2751 1244 2752
rect 1382 2756 1388 2757
rect 1382 2752 1383 2756
rect 1387 2752 1388 2756
rect 1382 2751 1388 2752
rect 1534 2756 1540 2757
rect 1534 2752 1535 2756
rect 1539 2752 1540 2756
rect 1534 2751 1540 2752
rect 1678 2756 1684 2757
rect 1678 2752 1679 2756
rect 1683 2752 1684 2756
rect 1678 2751 1684 2752
rect 1814 2756 1820 2757
rect 1814 2752 1815 2756
rect 1819 2752 1820 2756
rect 1934 2753 1935 2757
rect 1939 2753 1940 2757
rect 1934 2752 1940 2753
rect 1814 2751 1820 2752
rect 434 2741 440 2742
rect 110 2740 116 2741
rect 110 2736 111 2740
rect 115 2736 116 2740
rect 434 2737 435 2741
rect 439 2737 440 2741
rect 434 2736 440 2737
rect 594 2741 600 2742
rect 594 2737 595 2741
rect 599 2737 600 2741
rect 594 2736 600 2737
rect 754 2741 760 2742
rect 754 2737 755 2741
rect 759 2737 760 2741
rect 754 2736 760 2737
rect 906 2741 912 2742
rect 906 2737 907 2741
rect 911 2737 912 2741
rect 906 2736 912 2737
rect 1058 2741 1064 2742
rect 1058 2737 1059 2741
rect 1063 2737 1064 2741
rect 1058 2736 1064 2737
rect 1210 2741 1216 2742
rect 1210 2737 1211 2741
rect 1215 2737 1216 2741
rect 1210 2736 1216 2737
rect 1354 2741 1360 2742
rect 1354 2737 1355 2741
rect 1359 2737 1360 2741
rect 1354 2736 1360 2737
rect 1506 2741 1512 2742
rect 1506 2737 1507 2741
rect 1511 2737 1512 2741
rect 1506 2736 1512 2737
rect 1650 2741 1656 2742
rect 1650 2737 1651 2741
rect 1655 2737 1656 2741
rect 1650 2736 1656 2737
rect 1786 2741 1792 2742
rect 1786 2737 1787 2741
rect 1791 2737 1792 2741
rect 1786 2736 1792 2737
rect 1934 2740 1940 2741
rect 1934 2736 1935 2740
rect 1939 2736 1940 2740
rect 110 2735 116 2736
rect 112 2671 114 2735
rect 436 2671 438 2736
rect 596 2671 598 2736
rect 756 2671 758 2736
rect 908 2671 910 2736
rect 1060 2671 1062 2736
rect 1212 2671 1214 2736
rect 1356 2671 1358 2736
rect 1508 2671 1510 2736
rect 1652 2671 1654 2736
rect 1788 2671 1790 2736
rect 1934 2735 1940 2736
rect 1936 2671 1938 2735
rect 1976 2717 1978 2777
rect 1974 2716 1980 2717
rect 3060 2716 3062 2777
rect 3196 2716 3198 2777
rect 3332 2716 3334 2777
rect 3800 2717 3802 2777
rect 3840 2745 3842 2805
rect 3838 2744 3844 2745
rect 3860 2744 3862 2805
rect 3996 2744 3998 2805
rect 4132 2744 4134 2805
rect 4268 2744 4270 2805
rect 4404 2744 4406 2805
rect 4540 2744 4542 2805
rect 4676 2744 4678 2805
rect 4812 2744 4814 2805
rect 5664 2745 5666 2805
rect 5662 2744 5668 2745
rect 3838 2740 3839 2744
rect 3843 2740 3844 2744
rect 3838 2739 3844 2740
rect 3858 2743 3864 2744
rect 3858 2739 3859 2743
rect 3863 2739 3864 2743
rect 3858 2738 3864 2739
rect 3994 2743 4000 2744
rect 3994 2739 3995 2743
rect 3999 2739 4000 2743
rect 3994 2738 4000 2739
rect 4130 2743 4136 2744
rect 4130 2739 4131 2743
rect 4135 2739 4136 2743
rect 4130 2738 4136 2739
rect 4266 2743 4272 2744
rect 4266 2739 4267 2743
rect 4271 2739 4272 2743
rect 4266 2738 4272 2739
rect 4402 2743 4408 2744
rect 4402 2739 4403 2743
rect 4407 2739 4408 2743
rect 4402 2738 4408 2739
rect 4538 2743 4544 2744
rect 4538 2739 4539 2743
rect 4543 2739 4544 2743
rect 4538 2738 4544 2739
rect 4674 2743 4680 2744
rect 4674 2739 4675 2743
rect 4679 2739 4680 2743
rect 4674 2738 4680 2739
rect 4810 2743 4816 2744
rect 4810 2739 4811 2743
rect 4815 2739 4816 2743
rect 5662 2740 5663 2744
rect 5667 2740 5668 2744
rect 5662 2739 5668 2740
rect 4810 2738 4816 2739
rect 3886 2728 3892 2729
rect 3838 2727 3844 2728
rect 3838 2723 3839 2727
rect 3843 2723 3844 2727
rect 3886 2724 3887 2728
rect 3891 2724 3892 2728
rect 3886 2723 3892 2724
rect 4022 2728 4028 2729
rect 4022 2724 4023 2728
rect 4027 2724 4028 2728
rect 4022 2723 4028 2724
rect 4158 2728 4164 2729
rect 4158 2724 4159 2728
rect 4163 2724 4164 2728
rect 4158 2723 4164 2724
rect 4294 2728 4300 2729
rect 4294 2724 4295 2728
rect 4299 2724 4300 2728
rect 4294 2723 4300 2724
rect 4430 2728 4436 2729
rect 4430 2724 4431 2728
rect 4435 2724 4436 2728
rect 4430 2723 4436 2724
rect 4566 2728 4572 2729
rect 4566 2724 4567 2728
rect 4571 2724 4572 2728
rect 4566 2723 4572 2724
rect 4702 2728 4708 2729
rect 4702 2724 4703 2728
rect 4707 2724 4708 2728
rect 4702 2723 4708 2724
rect 4838 2728 4844 2729
rect 4838 2724 4839 2728
rect 4843 2724 4844 2728
rect 4838 2723 4844 2724
rect 5662 2727 5668 2728
rect 5662 2723 5663 2727
rect 5667 2723 5668 2727
rect 3838 2722 3844 2723
rect 3798 2716 3804 2717
rect 1974 2712 1975 2716
rect 1979 2712 1980 2716
rect 1974 2711 1980 2712
rect 3058 2715 3064 2716
rect 3058 2711 3059 2715
rect 3063 2711 3064 2715
rect 3058 2710 3064 2711
rect 3194 2715 3200 2716
rect 3194 2711 3195 2715
rect 3199 2711 3200 2715
rect 3194 2710 3200 2711
rect 3330 2715 3336 2716
rect 3330 2711 3331 2715
rect 3335 2711 3336 2715
rect 3798 2712 3799 2716
rect 3803 2712 3804 2716
rect 3798 2711 3804 2712
rect 3330 2710 3336 2711
rect 3086 2700 3092 2701
rect 1974 2699 1980 2700
rect 1974 2695 1975 2699
rect 1979 2695 1980 2699
rect 3086 2696 3087 2700
rect 3091 2696 3092 2700
rect 3086 2695 3092 2696
rect 3222 2700 3228 2701
rect 3222 2696 3223 2700
rect 3227 2696 3228 2700
rect 3222 2695 3228 2696
rect 3358 2700 3364 2701
rect 3358 2696 3359 2700
rect 3363 2696 3364 2700
rect 3358 2695 3364 2696
rect 3798 2699 3804 2700
rect 3840 2699 3842 2722
rect 3888 2699 3890 2723
rect 4024 2699 4026 2723
rect 4160 2699 4162 2723
rect 4296 2699 4298 2723
rect 4432 2699 4434 2723
rect 4568 2699 4570 2723
rect 4704 2699 4706 2723
rect 4840 2699 4842 2723
rect 5662 2722 5668 2723
rect 5664 2699 5666 2722
rect 3798 2695 3799 2699
rect 3803 2695 3804 2699
rect 1974 2694 1980 2695
rect 111 2670 115 2671
rect 111 2665 115 2666
rect 355 2670 359 2671
rect 355 2665 359 2666
rect 435 2670 439 2671
rect 435 2665 439 2666
rect 539 2670 543 2671
rect 539 2665 543 2666
rect 595 2670 599 2671
rect 595 2665 599 2666
rect 715 2670 719 2671
rect 715 2665 719 2666
rect 755 2670 759 2671
rect 755 2665 759 2666
rect 883 2670 887 2671
rect 883 2665 887 2666
rect 907 2670 911 2671
rect 907 2665 911 2666
rect 1043 2670 1047 2671
rect 1043 2665 1047 2666
rect 1059 2670 1063 2671
rect 1059 2665 1063 2666
rect 1203 2670 1207 2671
rect 1203 2665 1207 2666
rect 1211 2670 1215 2671
rect 1211 2665 1215 2666
rect 1355 2670 1359 2671
rect 1355 2665 1359 2666
rect 1507 2670 1511 2671
rect 1507 2665 1511 2666
rect 1651 2670 1655 2671
rect 1651 2665 1655 2666
rect 1787 2670 1791 2671
rect 1787 2665 1791 2666
rect 1935 2670 1939 2671
rect 1935 2665 1939 2666
rect 112 2605 114 2665
rect 110 2604 116 2605
rect 356 2604 358 2665
rect 540 2604 542 2665
rect 716 2604 718 2665
rect 884 2604 886 2665
rect 1044 2604 1046 2665
rect 1204 2604 1206 2665
rect 1356 2604 1358 2665
rect 1508 2604 1510 2665
rect 1652 2604 1654 2665
rect 1788 2604 1790 2665
rect 1936 2605 1938 2665
rect 1976 2647 1978 2694
rect 3088 2647 3090 2695
rect 3224 2647 3226 2695
rect 3360 2647 3362 2695
rect 3798 2694 3804 2695
rect 3839 2698 3843 2699
rect 3800 2647 3802 2694
rect 3839 2693 3843 2694
rect 3887 2698 3891 2699
rect 3887 2693 3891 2694
rect 4023 2698 4027 2699
rect 4023 2693 4027 2694
rect 4055 2698 4059 2699
rect 4055 2693 4059 2694
rect 4159 2698 4163 2699
rect 4159 2693 4163 2694
rect 4295 2698 4299 2699
rect 4295 2693 4299 2694
rect 4303 2698 4307 2699
rect 4303 2693 4307 2694
rect 4431 2698 4435 2699
rect 4431 2693 4435 2694
rect 4567 2698 4571 2699
rect 4567 2693 4571 2694
rect 4583 2698 4587 2699
rect 4583 2693 4587 2694
rect 4703 2698 4707 2699
rect 4703 2693 4707 2694
rect 4839 2698 4843 2699
rect 4839 2693 4843 2694
rect 4895 2698 4899 2699
rect 4895 2693 4899 2694
rect 5231 2698 5235 2699
rect 5231 2693 5235 2694
rect 5543 2698 5547 2699
rect 5543 2693 5547 2694
rect 5663 2698 5667 2699
rect 5663 2693 5667 2694
rect 3840 2670 3842 2693
rect 3838 2669 3844 2670
rect 4056 2669 4058 2693
rect 4304 2669 4306 2693
rect 4584 2669 4586 2693
rect 4896 2669 4898 2693
rect 5232 2669 5234 2693
rect 5544 2669 5546 2693
rect 5664 2670 5666 2693
rect 5662 2669 5668 2670
rect 3838 2665 3839 2669
rect 3843 2665 3844 2669
rect 3838 2664 3844 2665
rect 4054 2668 4060 2669
rect 4054 2664 4055 2668
rect 4059 2664 4060 2668
rect 4054 2663 4060 2664
rect 4302 2668 4308 2669
rect 4302 2664 4303 2668
rect 4307 2664 4308 2668
rect 4302 2663 4308 2664
rect 4582 2668 4588 2669
rect 4582 2664 4583 2668
rect 4587 2664 4588 2668
rect 4582 2663 4588 2664
rect 4894 2668 4900 2669
rect 4894 2664 4895 2668
rect 4899 2664 4900 2668
rect 4894 2663 4900 2664
rect 5230 2668 5236 2669
rect 5230 2664 5231 2668
rect 5235 2664 5236 2668
rect 5230 2663 5236 2664
rect 5542 2668 5548 2669
rect 5542 2664 5543 2668
rect 5547 2664 5548 2668
rect 5662 2665 5663 2669
rect 5667 2665 5668 2669
rect 5662 2664 5668 2665
rect 5542 2663 5548 2664
rect 4026 2653 4032 2654
rect 3838 2652 3844 2653
rect 3838 2648 3839 2652
rect 3843 2648 3844 2652
rect 4026 2649 4027 2653
rect 4031 2649 4032 2653
rect 4026 2648 4032 2649
rect 4274 2653 4280 2654
rect 4274 2649 4275 2653
rect 4279 2649 4280 2653
rect 4274 2648 4280 2649
rect 4554 2653 4560 2654
rect 4554 2649 4555 2653
rect 4559 2649 4560 2653
rect 4554 2648 4560 2649
rect 4866 2653 4872 2654
rect 4866 2649 4867 2653
rect 4871 2649 4872 2653
rect 4866 2648 4872 2649
rect 5202 2653 5208 2654
rect 5202 2649 5203 2653
rect 5207 2649 5208 2653
rect 5202 2648 5208 2649
rect 5514 2653 5520 2654
rect 5514 2649 5515 2653
rect 5519 2649 5520 2653
rect 5514 2648 5520 2649
rect 5662 2652 5668 2653
rect 5662 2648 5663 2652
rect 5667 2648 5668 2652
rect 3838 2647 3844 2648
rect 1975 2646 1979 2647
rect 1975 2641 1979 2642
rect 3087 2646 3091 2647
rect 3087 2641 3091 2642
rect 3135 2646 3139 2647
rect 3135 2641 3139 2642
rect 3223 2646 3227 2647
rect 3223 2641 3227 2642
rect 3271 2646 3275 2647
rect 3271 2641 3275 2642
rect 3359 2646 3363 2647
rect 3359 2641 3363 2642
rect 3407 2646 3411 2647
rect 3407 2641 3411 2642
rect 3543 2646 3547 2647
rect 3543 2641 3547 2642
rect 3679 2646 3683 2647
rect 3679 2641 3683 2642
rect 3799 2646 3803 2647
rect 3799 2641 3803 2642
rect 1976 2618 1978 2641
rect 1974 2617 1980 2618
rect 3136 2617 3138 2641
rect 3272 2617 3274 2641
rect 3408 2617 3410 2641
rect 3544 2617 3546 2641
rect 3680 2617 3682 2641
rect 3800 2618 3802 2641
rect 3798 2617 3804 2618
rect 1974 2613 1975 2617
rect 1979 2613 1980 2617
rect 1974 2612 1980 2613
rect 3134 2616 3140 2617
rect 3134 2612 3135 2616
rect 3139 2612 3140 2616
rect 3134 2611 3140 2612
rect 3270 2616 3276 2617
rect 3270 2612 3271 2616
rect 3275 2612 3276 2616
rect 3270 2611 3276 2612
rect 3406 2616 3412 2617
rect 3406 2612 3407 2616
rect 3411 2612 3412 2616
rect 3406 2611 3412 2612
rect 3542 2616 3548 2617
rect 3542 2612 3543 2616
rect 3547 2612 3548 2616
rect 3542 2611 3548 2612
rect 3678 2616 3684 2617
rect 3678 2612 3679 2616
rect 3683 2612 3684 2616
rect 3798 2613 3799 2617
rect 3803 2613 3804 2617
rect 3798 2612 3804 2613
rect 3678 2611 3684 2612
rect 1934 2604 1940 2605
rect 110 2600 111 2604
rect 115 2600 116 2604
rect 110 2599 116 2600
rect 354 2603 360 2604
rect 354 2599 355 2603
rect 359 2599 360 2603
rect 354 2598 360 2599
rect 538 2603 544 2604
rect 538 2599 539 2603
rect 543 2599 544 2603
rect 538 2598 544 2599
rect 714 2603 720 2604
rect 714 2599 715 2603
rect 719 2599 720 2603
rect 714 2598 720 2599
rect 882 2603 888 2604
rect 882 2599 883 2603
rect 887 2599 888 2603
rect 882 2598 888 2599
rect 1042 2603 1048 2604
rect 1042 2599 1043 2603
rect 1047 2599 1048 2603
rect 1042 2598 1048 2599
rect 1202 2603 1208 2604
rect 1202 2599 1203 2603
rect 1207 2599 1208 2603
rect 1202 2598 1208 2599
rect 1354 2603 1360 2604
rect 1354 2599 1355 2603
rect 1359 2599 1360 2603
rect 1354 2598 1360 2599
rect 1506 2603 1512 2604
rect 1506 2599 1507 2603
rect 1511 2599 1512 2603
rect 1506 2598 1512 2599
rect 1650 2603 1656 2604
rect 1650 2599 1651 2603
rect 1655 2599 1656 2603
rect 1650 2598 1656 2599
rect 1786 2603 1792 2604
rect 1786 2599 1787 2603
rect 1791 2599 1792 2603
rect 1934 2600 1935 2604
rect 1939 2600 1940 2604
rect 3106 2601 3112 2602
rect 1934 2599 1940 2600
rect 1974 2600 1980 2601
rect 1786 2598 1792 2599
rect 1974 2596 1975 2600
rect 1979 2596 1980 2600
rect 3106 2597 3107 2601
rect 3111 2597 3112 2601
rect 3106 2596 3112 2597
rect 3242 2601 3248 2602
rect 3242 2597 3243 2601
rect 3247 2597 3248 2601
rect 3242 2596 3248 2597
rect 3378 2601 3384 2602
rect 3378 2597 3379 2601
rect 3383 2597 3384 2601
rect 3378 2596 3384 2597
rect 3514 2601 3520 2602
rect 3514 2597 3515 2601
rect 3519 2597 3520 2601
rect 3514 2596 3520 2597
rect 3650 2601 3656 2602
rect 3650 2597 3651 2601
rect 3655 2597 3656 2601
rect 3650 2596 3656 2597
rect 3798 2600 3804 2601
rect 3798 2596 3799 2600
rect 3803 2596 3804 2600
rect 1974 2595 1980 2596
rect 382 2588 388 2589
rect 110 2587 116 2588
rect 110 2583 111 2587
rect 115 2583 116 2587
rect 382 2584 383 2588
rect 387 2584 388 2588
rect 382 2583 388 2584
rect 566 2588 572 2589
rect 566 2584 567 2588
rect 571 2584 572 2588
rect 566 2583 572 2584
rect 742 2588 748 2589
rect 742 2584 743 2588
rect 747 2584 748 2588
rect 742 2583 748 2584
rect 910 2588 916 2589
rect 910 2584 911 2588
rect 915 2584 916 2588
rect 910 2583 916 2584
rect 1070 2588 1076 2589
rect 1070 2584 1071 2588
rect 1075 2584 1076 2588
rect 1070 2583 1076 2584
rect 1230 2588 1236 2589
rect 1230 2584 1231 2588
rect 1235 2584 1236 2588
rect 1230 2583 1236 2584
rect 1382 2588 1388 2589
rect 1382 2584 1383 2588
rect 1387 2584 1388 2588
rect 1382 2583 1388 2584
rect 1534 2588 1540 2589
rect 1534 2584 1535 2588
rect 1539 2584 1540 2588
rect 1534 2583 1540 2584
rect 1678 2588 1684 2589
rect 1678 2584 1679 2588
rect 1683 2584 1684 2588
rect 1678 2583 1684 2584
rect 1814 2588 1820 2589
rect 1814 2584 1815 2588
rect 1819 2584 1820 2588
rect 1814 2583 1820 2584
rect 1934 2587 1940 2588
rect 1934 2583 1935 2587
rect 1939 2583 1940 2587
rect 110 2582 116 2583
rect 112 2559 114 2582
rect 384 2559 386 2583
rect 568 2559 570 2583
rect 744 2559 746 2583
rect 912 2559 914 2583
rect 1072 2559 1074 2583
rect 1232 2559 1234 2583
rect 1384 2559 1386 2583
rect 1536 2559 1538 2583
rect 1680 2559 1682 2583
rect 1816 2559 1818 2583
rect 1934 2582 1940 2583
rect 1936 2559 1938 2582
rect 111 2558 115 2559
rect 111 2553 115 2554
rect 231 2558 235 2559
rect 231 2553 235 2554
rect 383 2558 387 2559
rect 383 2553 387 2554
rect 423 2558 427 2559
rect 423 2553 427 2554
rect 567 2558 571 2559
rect 567 2553 571 2554
rect 623 2558 627 2559
rect 623 2553 627 2554
rect 743 2558 747 2559
rect 743 2553 747 2554
rect 823 2558 827 2559
rect 823 2553 827 2554
rect 911 2558 915 2559
rect 911 2553 915 2554
rect 1023 2558 1027 2559
rect 1023 2553 1027 2554
rect 1071 2558 1075 2559
rect 1071 2553 1075 2554
rect 1223 2558 1227 2559
rect 1223 2553 1227 2554
rect 1231 2558 1235 2559
rect 1231 2553 1235 2554
rect 1383 2558 1387 2559
rect 1383 2553 1387 2554
rect 1423 2558 1427 2559
rect 1423 2553 1427 2554
rect 1535 2558 1539 2559
rect 1535 2553 1539 2554
rect 1631 2558 1635 2559
rect 1631 2553 1635 2554
rect 1679 2558 1683 2559
rect 1679 2553 1683 2554
rect 1815 2558 1819 2559
rect 1815 2553 1819 2554
rect 1935 2558 1939 2559
rect 1935 2553 1939 2554
rect 112 2530 114 2553
rect 110 2529 116 2530
rect 232 2529 234 2553
rect 424 2529 426 2553
rect 624 2529 626 2553
rect 824 2529 826 2553
rect 1024 2529 1026 2553
rect 1224 2529 1226 2553
rect 1424 2529 1426 2553
rect 1632 2529 1634 2553
rect 1816 2529 1818 2553
rect 1936 2530 1938 2553
rect 1934 2529 1940 2530
rect 110 2525 111 2529
rect 115 2525 116 2529
rect 110 2524 116 2525
rect 230 2528 236 2529
rect 230 2524 231 2528
rect 235 2524 236 2528
rect 230 2523 236 2524
rect 422 2528 428 2529
rect 422 2524 423 2528
rect 427 2524 428 2528
rect 422 2523 428 2524
rect 622 2528 628 2529
rect 622 2524 623 2528
rect 627 2524 628 2528
rect 622 2523 628 2524
rect 822 2528 828 2529
rect 822 2524 823 2528
rect 827 2524 828 2528
rect 822 2523 828 2524
rect 1022 2528 1028 2529
rect 1022 2524 1023 2528
rect 1027 2524 1028 2528
rect 1022 2523 1028 2524
rect 1222 2528 1228 2529
rect 1222 2524 1223 2528
rect 1227 2524 1228 2528
rect 1222 2523 1228 2524
rect 1422 2528 1428 2529
rect 1422 2524 1423 2528
rect 1427 2524 1428 2528
rect 1422 2523 1428 2524
rect 1630 2528 1636 2529
rect 1630 2524 1631 2528
rect 1635 2524 1636 2528
rect 1630 2523 1636 2524
rect 1814 2528 1820 2529
rect 1814 2524 1815 2528
rect 1819 2524 1820 2528
rect 1934 2525 1935 2529
rect 1939 2525 1940 2529
rect 1976 2527 1978 2595
rect 3108 2527 3110 2596
rect 3244 2527 3246 2596
rect 3380 2527 3382 2596
rect 3516 2527 3518 2596
rect 3652 2527 3654 2596
rect 3798 2595 3804 2596
rect 3800 2527 3802 2595
rect 3840 2583 3842 2647
rect 4028 2583 4030 2648
rect 4276 2583 4278 2648
rect 4556 2583 4558 2648
rect 4868 2583 4870 2648
rect 5204 2583 5206 2648
rect 5516 2583 5518 2648
rect 5662 2647 5668 2648
rect 5664 2583 5666 2647
rect 3839 2582 3843 2583
rect 3839 2577 3843 2578
rect 4027 2582 4031 2583
rect 4027 2577 4031 2578
rect 4259 2582 4263 2583
rect 4259 2577 4263 2578
rect 4275 2582 4279 2583
rect 4275 2577 4279 2578
rect 4475 2582 4479 2583
rect 4475 2577 4479 2578
rect 4555 2582 4559 2583
rect 4555 2577 4559 2578
rect 4715 2582 4719 2583
rect 4715 2577 4719 2578
rect 4867 2582 4871 2583
rect 4867 2577 4871 2578
rect 4979 2582 4983 2583
rect 4979 2577 4983 2578
rect 5203 2582 5207 2583
rect 5203 2577 5207 2578
rect 5259 2582 5263 2583
rect 5259 2577 5263 2578
rect 5515 2582 5519 2583
rect 5515 2577 5519 2578
rect 5663 2582 5667 2583
rect 5663 2577 5667 2578
rect 1934 2524 1940 2525
rect 1975 2526 1979 2527
rect 1814 2523 1820 2524
rect 1975 2521 1979 2522
rect 1995 2526 1999 2527
rect 1995 2521 1999 2522
rect 2235 2526 2239 2527
rect 2235 2521 2239 2522
rect 2483 2526 2487 2527
rect 2483 2521 2487 2522
rect 2715 2526 2719 2527
rect 2715 2521 2719 2522
rect 2939 2526 2943 2527
rect 2939 2521 2943 2522
rect 3107 2526 3111 2527
rect 3107 2521 3111 2522
rect 3155 2526 3159 2527
rect 3155 2521 3159 2522
rect 3243 2526 3247 2527
rect 3243 2521 3247 2522
rect 3363 2526 3367 2527
rect 3363 2521 3367 2522
rect 3379 2526 3383 2527
rect 3379 2521 3383 2522
rect 3515 2526 3519 2527
rect 3515 2521 3519 2522
rect 3579 2526 3583 2527
rect 3579 2521 3583 2522
rect 3651 2526 3655 2527
rect 3651 2521 3655 2522
rect 3799 2526 3803 2527
rect 3799 2521 3803 2522
rect 202 2513 208 2514
rect 110 2512 116 2513
rect 110 2508 111 2512
rect 115 2508 116 2512
rect 202 2509 203 2513
rect 207 2509 208 2513
rect 202 2508 208 2509
rect 394 2513 400 2514
rect 394 2509 395 2513
rect 399 2509 400 2513
rect 394 2508 400 2509
rect 594 2513 600 2514
rect 594 2509 595 2513
rect 599 2509 600 2513
rect 594 2508 600 2509
rect 794 2513 800 2514
rect 794 2509 795 2513
rect 799 2509 800 2513
rect 794 2508 800 2509
rect 994 2513 1000 2514
rect 994 2509 995 2513
rect 999 2509 1000 2513
rect 994 2508 1000 2509
rect 1194 2513 1200 2514
rect 1194 2509 1195 2513
rect 1199 2509 1200 2513
rect 1194 2508 1200 2509
rect 1394 2513 1400 2514
rect 1394 2509 1395 2513
rect 1399 2509 1400 2513
rect 1394 2508 1400 2509
rect 1602 2513 1608 2514
rect 1602 2509 1603 2513
rect 1607 2509 1608 2513
rect 1602 2508 1608 2509
rect 1786 2513 1792 2514
rect 1786 2509 1787 2513
rect 1791 2509 1792 2513
rect 1786 2508 1792 2509
rect 1934 2512 1940 2513
rect 1934 2508 1935 2512
rect 1939 2508 1940 2512
rect 110 2507 116 2508
rect 112 2427 114 2507
rect 204 2427 206 2508
rect 396 2427 398 2508
rect 596 2427 598 2508
rect 796 2427 798 2508
rect 996 2427 998 2508
rect 1196 2427 1198 2508
rect 1396 2427 1398 2508
rect 1604 2427 1606 2508
rect 1788 2427 1790 2508
rect 1934 2507 1940 2508
rect 1936 2427 1938 2507
rect 1976 2461 1978 2521
rect 1974 2460 1980 2461
rect 1996 2460 1998 2521
rect 2236 2460 2238 2521
rect 2484 2460 2486 2521
rect 2716 2460 2718 2521
rect 2940 2460 2942 2521
rect 3156 2460 3158 2521
rect 3364 2460 3366 2521
rect 3580 2460 3582 2521
rect 3800 2461 3802 2521
rect 3840 2517 3842 2577
rect 3838 2516 3844 2517
rect 4260 2516 4262 2577
rect 4476 2516 4478 2577
rect 4716 2516 4718 2577
rect 4980 2516 4982 2577
rect 5260 2516 5262 2577
rect 5516 2516 5518 2577
rect 5664 2517 5666 2577
rect 5662 2516 5668 2517
rect 3838 2512 3839 2516
rect 3843 2512 3844 2516
rect 3838 2511 3844 2512
rect 4258 2515 4264 2516
rect 4258 2511 4259 2515
rect 4263 2511 4264 2515
rect 4258 2510 4264 2511
rect 4474 2515 4480 2516
rect 4474 2511 4475 2515
rect 4479 2511 4480 2515
rect 4474 2510 4480 2511
rect 4714 2515 4720 2516
rect 4714 2511 4715 2515
rect 4719 2511 4720 2515
rect 4714 2510 4720 2511
rect 4978 2515 4984 2516
rect 4978 2511 4979 2515
rect 4983 2511 4984 2515
rect 4978 2510 4984 2511
rect 5258 2515 5264 2516
rect 5258 2511 5259 2515
rect 5263 2511 5264 2515
rect 5258 2510 5264 2511
rect 5514 2515 5520 2516
rect 5514 2511 5515 2515
rect 5519 2511 5520 2515
rect 5662 2512 5663 2516
rect 5667 2512 5668 2516
rect 5662 2511 5668 2512
rect 5514 2510 5520 2511
rect 4286 2500 4292 2501
rect 3838 2499 3844 2500
rect 3838 2495 3839 2499
rect 3843 2495 3844 2499
rect 4286 2496 4287 2500
rect 4291 2496 4292 2500
rect 4286 2495 4292 2496
rect 4502 2500 4508 2501
rect 4502 2496 4503 2500
rect 4507 2496 4508 2500
rect 4502 2495 4508 2496
rect 4742 2500 4748 2501
rect 4742 2496 4743 2500
rect 4747 2496 4748 2500
rect 4742 2495 4748 2496
rect 5006 2500 5012 2501
rect 5006 2496 5007 2500
rect 5011 2496 5012 2500
rect 5006 2495 5012 2496
rect 5286 2500 5292 2501
rect 5286 2496 5287 2500
rect 5291 2496 5292 2500
rect 5286 2495 5292 2496
rect 5542 2500 5548 2501
rect 5542 2496 5543 2500
rect 5547 2496 5548 2500
rect 5542 2495 5548 2496
rect 5662 2499 5668 2500
rect 5662 2495 5663 2499
rect 5667 2495 5668 2499
rect 3838 2494 3844 2495
rect 3840 2467 3842 2494
rect 4288 2467 4290 2495
rect 4504 2467 4506 2495
rect 4744 2467 4746 2495
rect 5008 2467 5010 2495
rect 5288 2467 5290 2495
rect 5544 2467 5546 2495
rect 5662 2494 5668 2495
rect 5664 2467 5666 2494
rect 3839 2466 3843 2467
rect 3839 2461 3843 2462
rect 4287 2466 4291 2467
rect 4287 2461 4291 2462
rect 4503 2466 4507 2467
rect 4503 2461 4507 2462
rect 4663 2466 4667 2467
rect 4663 2461 4667 2462
rect 4743 2466 4747 2467
rect 4743 2461 4747 2462
rect 4847 2466 4851 2467
rect 4847 2461 4851 2462
rect 5007 2466 5011 2467
rect 5007 2461 5011 2462
rect 5023 2466 5027 2467
rect 5023 2461 5027 2462
rect 5199 2466 5203 2467
rect 5199 2461 5203 2462
rect 5287 2466 5291 2467
rect 5287 2461 5291 2462
rect 5383 2466 5387 2467
rect 5383 2461 5387 2462
rect 5543 2466 5547 2467
rect 5543 2461 5547 2462
rect 5663 2466 5667 2467
rect 5663 2461 5667 2462
rect 3798 2460 3804 2461
rect 1974 2456 1975 2460
rect 1979 2456 1980 2460
rect 1974 2455 1980 2456
rect 1994 2459 2000 2460
rect 1994 2455 1995 2459
rect 1999 2455 2000 2459
rect 1994 2454 2000 2455
rect 2234 2459 2240 2460
rect 2234 2455 2235 2459
rect 2239 2455 2240 2459
rect 2234 2454 2240 2455
rect 2482 2459 2488 2460
rect 2482 2455 2483 2459
rect 2487 2455 2488 2459
rect 2482 2454 2488 2455
rect 2714 2459 2720 2460
rect 2714 2455 2715 2459
rect 2719 2455 2720 2459
rect 2714 2454 2720 2455
rect 2938 2459 2944 2460
rect 2938 2455 2939 2459
rect 2943 2455 2944 2459
rect 2938 2454 2944 2455
rect 3154 2459 3160 2460
rect 3154 2455 3155 2459
rect 3159 2455 3160 2459
rect 3154 2454 3160 2455
rect 3362 2459 3368 2460
rect 3362 2455 3363 2459
rect 3367 2455 3368 2459
rect 3362 2454 3368 2455
rect 3578 2459 3584 2460
rect 3578 2455 3579 2459
rect 3583 2455 3584 2459
rect 3798 2456 3799 2460
rect 3803 2456 3804 2460
rect 3798 2455 3804 2456
rect 3578 2454 3584 2455
rect 2022 2444 2028 2445
rect 1974 2443 1980 2444
rect 1974 2439 1975 2443
rect 1979 2439 1980 2443
rect 2022 2440 2023 2444
rect 2027 2440 2028 2444
rect 2022 2439 2028 2440
rect 2262 2444 2268 2445
rect 2262 2440 2263 2444
rect 2267 2440 2268 2444
rect 2262 2439 2268 2440
rect 2510 2444 2516 2445
rect 2510 2440 2511 2444
rect 2515 2440 2516 2444
rect 2510 2439 2516 2440
rect 2742 2444 2748 2445
rect 2742 2440 2743 2444
rect 2747 2440 2748 2444
rect 2742 2439 2748 2440
rect 2966 2444 2972 2445
rect 2966 2440 2967 2444
rect 2971 2440 2972 2444
rect 2966 2439 2972 2440
rect 3182 2444 3188 2445
rect 3182 2440 3183 2444
rect 3187 2440 3188 2444
rect 3182 2439 3188 2440
rect 3390 2444 3396 2445
rect 3390 2440 3391 2444
rect 3395 2440 3396 2444
rect 3390 2439 3396 2440
rect 3606 2444 3612 2445
rect 3606 2440 3607 2444
rect 3611 2440 3612 2444
rect 3606 2439 3612 2440
rect 3798 2443 3804 2444
rect 3798 2439 3799 2443
rect 3803 2439 3804 2443
rect 1974 2438 1980 2439
rect 111 2426 115 2427
rect 111 2421 115 2422
rect 203 2426 207 2427
rect 203 2421 207 2422
rect 219 2426 223 2427
rect 219 2421 223 2422
rect 395 2426 399 2427
rect 395 2421 399 2422
rect 403 2426 407 2427
rect 403 2421 407 2422
rect 595 2426 599 2427
rect 595 2421 599 2422
rect 787 2426 791 2427
rect 787 2421 791 2422
rect 795 2426 799 2427
rect 795 2421 799 2422
rect 979 2426 983 2427
rect 979 2421 983 2422
rect 995 2426 999 2427
rect 995 2421 999 2422
rect 1195 2426 1199 2427
rect 1195 2421 1199 2422
rect 1395 2426 1399 2427
rect 1395 2421 1399 2422
rect 1603 2426 1607 2427
rect 1603 2421 1607 2422
rect 1787 2426 1791 2427
rect 1787 2421 1791 2422
rect 1935 2426 1939 2427
rect 1935 2421 1939 2422
rect 112 2361 114 2421
rect 110 2360 116 2361
rect 220 2360 222 2421
rect 404 2360 406 2421
rect 596 2360 598 2421
rect 788 2360 790 2421
rect 980 2360 982 2421
rect 1936 2361 1938 2421
rect 1976 2415 1978 2438
rect 2024 2415 2026 2439
rect 2264 2415 2266 2439
rect 2512 2415 2514 2439
rect 2744 2415 2746 2439
rect 2968 2415 2970 2439
rect 3184 2415 3186 2439
rect 3392 2415 3394 2439
rect 3608 2415 3610 2439
rect 3798 2438 3804 2439
rect 3840 2438 3842 2461
rect 3800 2415 3802 2438
rect 3838 2437 3844 2438
rect 4664 2437 4666 2461
rect 4848 2437 4850 2461
rect 5024 2437 5026 2461
rect 5200 2437 5202 2461
rect 5384 2437 5386 2461
rect 5544 2437 5546 2461
rect 5664 2438 5666 2461
rect 5662 2437 5668 2438
rect 3838 2433 3839 2437
rect 3843 2433 3844 2437
rect 3838 2432 3844 2433
rect 4662 2436 4668 2437
rect 4662 2432 4663 2436
rect 4667 2432 4668 2436
rect 4662 2431 4668 2432
rect 4846 2436 4852 2437
rect 4846 2432 4847 2436
rect 4851 2432 4852 2436
rect 4846 2431 4852 2432
rect 5022 2436 5028 2437
rect 5022 2432 5023 2436
rect 5027 2432 5028 2436
rect 5022 2431 5028 2432
rect 5198 2436 5204 2437
rect 5198 2432 5199 2436
rect 5203 2432 5204 2436
rect 5198 2431 5204 2432
rect 5382 2436 5388 2437
rect 5382 2432 5383 2436
rect 5387 2432 5388 2436
rect 5382 2431 5388 2432
rect 5542 2436 5548 2437
rect 5542 2432 5543 2436
rect 5547 2432 5548 2436
rect 5662 2433 5663 2437
rect 5667 2433 5668 2437
rect 5662 2432 5668 2433
rect 5542 2431 5548 2432
rect 4634 2421 4640 2422
rect 3838 2420 3844 2421
rect 3838 2416 3839 2420
rect 3843 2416 3844 2420
rect 4634 2417 4635 2421
rect 4639 2417 4640 2421
rect 4634 2416 4640 2417
rect 4818 2421 4824 2422
rect 4818 2417 4819 2421
rect 4823 2417 4824 2421
rect 4818 2416 4824 2417
rect 4994 2421 5000 2422
rect 4994 2417 4995 2421
rect 4999 2417 5000 2421
rect 4994 2416 5000 2417
rect 5170 2421 5176 2422
rect 5170 2417 5171 2421
rect 5175 2417 5176 2421
rect 5170 2416 5176 2417
rect 5354 2421 5360 2422
rect 5354 2417 5355 2421
rect 5359 2417 5360 2421
rect 5354 2416 5360 2417
rect 5514 2421 5520 2422
rect 5514 2417 5515 2421
rect 5519 2417 5520 2421
rect 5514 2416 5520 2417
rect 5662 2420 5668 2421
rect 5662 2416 5663 2420
rect 5667 2416 5668 2420
rect 3838 2415 3844 2416
rect 1975 2414 1979 2415
rect 1975 2409 1979 2410
rect 2023 2414 2027 2415
rect 2023 2409 2027 2410
rect 2159 2414 2163 2415
rect 2159 2409 2163 2410
rect 2263 2414 2267 2415
rect 2263 2409 2267 2410
rect 2295 2414 2299 2415
rect 2295 2409 2299 2410
rect 2431 2414 2435 2415
rect 2431 2409 2435 2410
rect 2511 2414 2515 2415
rect 2511 2409 2515 2410
rect 2567 2414 2571 2415
rect 2567 2409 2571 2410
rect 2711 2414 2715 2415
rect 2711 2409 2715 2410
rect 2743 2414 2747 2415
rect 2743 2409 2747 2410
rect 2855 2414 2859 2415
rect 2855 2409 2859 2410
rect 2967 2414 2971 2415
rect 2967 2409 2971 2410
rect 3007 2414 3011 2415
rect 3007 2409 3011 2410
rect 3159 2414 3163 2415
rect 3159 2409 3163 2410
rect 3183 2414 3187 2415
rect 3183 2409 3187 2410
rect 3311 2414 3315 2415
rect 3311 2409 3315 2410
rect 3391 2414 3395 2415
rect 3391 2409 3395 2410
rect 3607 2414 3611 2415
rect 3607 2409 3611 2410
rect 3799 2414 3803 2415
rect 3799 2409 3803 2410
rect 1976 2386 1978 2409
rect 1974 2385 1980 2386
rect 2024 2385 2026 2409
rect 2160 2385 2162 2409
rect 2296 2385 2298 2409
rect 2432 2385 2434 2409
rect 2568 2385 2570 2409
rect 2712 2385 2714 2409
rect 2856 2385 2858 2409
rect 3008 2385 3010 2409
rect 3160 2385 3162 2409
rect 3312 2385 3314 2409
rect 3800 2386 3802 2409
rect 3798 2385 3804 2386
rect 1974 2381 1975 2385
rect 1979 2381 1980 2385
rect 1974 2380 1980 2381
rect 2022 2384 2028 2385
rect 2022 2380 2023 2384
rect 2027 2380 2028 2384
rect 2022 2379 2028 2380
rect 2158 2384 2164 2385
rect 2158 2380 2159 2384
rect 2163 2380 2164 2384
rect 2158 2379 2164 2380
rect 2294 2384 2300 2385
rect 2294 2380 2295 2384
rect 2299 2380 2300 2384
rect 2294 2379 2300 2380
rect 2430 2384 2436 2385
rect 2430 2380 2431 2384
rect 2435 2380 2436 2384
rect 2430 2379 2436 2380
rect 2566 2384 2572 2385
rect 2566 2380 2567 2384
rect 2571 2380 2572 2384
rect 2566 2379 2572 2380
rect 2710 2384 2716 2385
rect 2710 2380 2711 2384
rect 2715 2380 2716 2384
rect 2710 2379 2716 2380
rect 2854 2384 2860 2385
rect 2854 2380 2855 2384
rect 2859 2380 2860 2384
rect 2854 2379 2860 2380
rect 3006 2384 3012 2385
rect 3006 2380 3007 2384
rect 3011 2380 3012 2384
rect 3006 2379 3012 2380
rect 3158 2384 3164 2385
rect 3158 2380 3159 2384
rect 3163 2380 3164 2384
rect 3158 2379 3164 2380
rect 3310 2384 3316 2385
rect 3310 2380 3311 2384
rect 3315 2380 3316 2384
rect 3798 2381 3799 2385
rect 3803 2381 3804 2385
rect 3798 2380 3804 2381
rect 3310 2379 3316 2380
rect 1994 2369 2000 2370
rect 1974 2368 1980 2369
rect 1974 2364 1975 2368
rect 1979 2364 1980 2368
rect 1994 2365 1995 2369
rect 1999 2365 2000 2369
rect 1994 2364 2000 2365
rect 2130 2369 2136 2370
rect 2130 2365 2131 2369
rect 2135 2365 2136 2369
rect 2130 2364 2136 2365
rect 2266 2369 2272 2370
rect 2266 2365 2267 2369
rect 2271 2365 2272 2369
rect 2266 2364 2272 2365
rect 2402 2369 2408 2370
rect 2402 2365 2403 2369
rect 2407 2365 2408 2369
rect 2402 2364 2408 2365
rect 2538 2369 2544 2370
rect 2538 2365 2539 2369
rect 2543 2365 2544 2369
rect 2538 2364 2544 2365
rect 2682 2369 2688 2370
rect 2682 2365 2683 2369
rect 2687 2365 2688 2369
rect 2682 2364 2688 2365
rect 2826 2369 2832 2370
rect 2826 2365 2827 2369
rect 2831 2365 2832 2369
rect 2826 2364 2832 2365
rect 2978 2369 2984 2370
rect 2978 2365 2979 2369
rect 2983 2365 2984 2369
rect 2978 2364 2984 2365
rect 3130 2369 3136 2370
rect 3130 2365 3131 2369
rect 3135 2365 3136 2369
rect 3130 2364 3136 2365
rect 3282 2369 3288 2370
rect 3282 2365 3283 2369
rect 3287 2365 3288 2369
rect 3282 2364 3288 2365
rect 3798 2368 3804 2369
rect 3798 2364 3799 2368
rect 3803 2364 3804 2368
rect 1974 2363 1980 2364
rect 1934 2360 1940 2361
rect 110 2356 111 2360
rect 115 2356 116 2360
rect 110 2355 116 2356
rect 218 2359 224 2360
rect 218 2355 219 2359
rect 223 2355 224 2359
rect 218 2354 224 2355
rect 402 2359 408 2360
rect 402 2355 403 2359
rect 407 2355 408 2359
rect 402 2354 408 2355
rect 594 2359 600 2360
rect 594 2355 595 2359
rect 599 2355 600 2359
rect 594 2354 600 2355
rect 786 2359 792 2360
rect 786 2355 787 2359
rect 791 2355 792 2359
rect 786 2354 792 2355
rect 978 2359 984 2360
rect 978 2355 979 2359
rect 983 2355 984 2359
rect 1934 2356 1935 2360
rect 1939 2356 1940 2360
rect 1934 2355 1940 2356
rect 978 2354 984 2355
rect 246 2344 252 2345
rect 110 2343 116 2344
rect 110 2339 111 2343
rect 115 2339 116 2343
rect 246 2340 247 2344
rect 251 2340 252 2344
rect 246 2339 252 2340
rect 430 2344 436 2345
rect 430 2340 431 2344
rect 435 2340 436 2344
rect 430 2339 436 2340
rect 622 2344 628 2345
rect 622 2340 623 2344
rect 627 2340 628 2344
rect 622 2339 628 2340
rect 814 2344 820 2345
rect 814 2340 815 2344
rect 819 2340 820 2344
rect 814 2339 820 2340
rect 1006 2344 1012 2345
rect 1006 2340 1007 2344
rect 1011 2340 1012 2344
rect 1006 2339 1012 2340
rect 1934 2343 1940 2344
rect 1934 2339 1935 2343
rect 1939 2339 1940 2343
rect 110 2338 116 2339
rect 112 2311 114 2338
rect 248 2311 250 2339
rect 432 2311 434 2339
rect 624 2311 626 2339
rect 816 2311 818 2339
rect 1008 2311 1010 2339
rect 1934 2338 1940 2339
rect 1936 2311 1938 2338
rect 111 2310 115 2311
rect 111 2305 115 2306
rect 247 2310 251 2311
rect 247 2305 251 2306
rect 399 2310 403 2311
rect 399 2305 403 2306
rect 431 2310 435 2311
rect 431 2305 435 2306
rect 535 2310 539 2311
rect 535 2305 539 2306
rect 623 2310 627 2311
rect 623 2305 627 2306
rect 671 2310 675 2311
rect 671 2305 675 2306
rect 807 2310 811 2311
rect 807 2305 811 2306
rect 815 2310 819 2311
rect 815 2305 819 2306
rect 943 2310 947 2311
rect 943 2305 947 2306
rect 1007 2310 1011 2311
rect 1007 2305 1011 2306
rect 1935 2310 1939 2311
rect 1935 2305 1939 2306
rect 112 2282 114 2305
rect 110 2281 116 2282
rect 400 2281 402 2305
rect 536 2281 538 2305
rect 672 2281 674 2305
rect 808 2281 810 2305
rect 944 2281 946 2305
rect 1936 2282 1938 2305
rect 1976 2299 1978 2363
rect 1996 2299 1998 2364
rect 2132 2299 2134 2364
rect 2268 2299 2270 2364
rect 2404 2299 2406 2364
rect 2540 2299 2542 2364
rect 2684 2299 2686 2364
rect 2828 2299 2830 2364
rect 2980 2299 2982 2364
rect 3132 2299 3134 2364
rect 3284 2299 3286 2364
rect 3798 2363 3804 2364
rect 3800 2299 3802 2363
rect 3840 2351 3842 2415
rect 4636 2351 4638 2416
rect 4820 2351 4822 2416
rect 4996 2351 4998 2416
rect 5172 2351 5174 2416
rect 5356 2351 5358 2416
rect 5516 2351 5518 2416
rect 5662 2415 5668 2416
rect 5664 2351 5666 2415
rect 3839 2350 3843 2351
rect 3839 2345 3843 2346
rect 4635 2350 4639 2351
rect 4635 2345 4639 2346
rect 4675 2350 4679 2351
rect 4675 2345 4679 2346
rect 4819 2350 4823 2351
rect 4819 2345 4823 2346
rect 4963 2350 4967 2351
rect 4963 2345 4967 2346
rect 4995 2350 4999 2351
rect 4995 2345 4999 2346
rect 5115 2350 5119 2351
rect 5115 2345 5119 2346
rect 5171 2350 5175 2351
rect 5171 2345 5175 2346
rect 5267 2350 5271 2351
rect 5267 2345 5271 2346
rect 5355 2350 5359 2351
rect 5355 2345 5359 2346
rect 5419 2350 5423 2351
rect 5419 2345 5423 2346
rect 5515 2350 5519 2351
rect 5515 2345 5519 2346
rect 5663 2350 5667 2351
rect 5663 2345 5667 2346
rect 1975 2298 1979 2299
rect 1975 2293 1979 2294
rect 1995 2298 1999 2299
rect 1995 2293 1999 2294
rect 2043 2298 2047 2299
rect 2043 2293 2047 2294
rect 2131 2298 2135 2299
rect 2131 2293 2135 2294
rect 2179 2298 2183 2299
rect 2179 2293 2183 2294
rect 2267 2298 2271 2299
rect 2267 2293 2271 2294
rect 2315 2298 2319 2299
rect 2315 2293 2319 2294
rect 2403 2298 2407 2299
rect 2403 2293 2407 2294
rect 2451 2298 2455 2299
rect 2451 2293 2455 2294
rect 2539 2298 2543 2299
rect 2539 2293 2543 2294
rect 2587 2298 2591 2299
rect 2587 2293 2591 2294
rect 2683 2298 2687 2299
rect 2683 2293 2687 2294
rect 2723 2298 2727 2299
rect 2723 2293 2727 2294
rect 2827 2298 2831 2299
rect 2827 2293 2831 2294
rect 2859 2298 2863 2299
rect 2859 2293 2863 2294
rect 2979 2298 2983 2299
rect 2979 2293 2983 2294
rect 2995 2298 2999 2299
rect 2995 2293 2999 2294
rect 3131 2298 3135 2299
rect 3131 2293 3135 2294
rect 3283 2298 3287 2299
rect 3283 2293 3287 2294
rect 3799 2298 3803 2299
rect 3799 2293 3803 2294
rect 1934 2281 1940 2282
rect 110 2277 111 2281
rect 115 2277 116 2281
rect 110 2276 116 2277
rect 398 2280 404 2281
rect 398 2276 399 2280
rect 403 2276 404 2280
rect 398 2275 404 2276
rect 534 2280 540 2281
rect 534 2276 535 2280
rect 539 2276 540 2280
rect 534 2275 540 2276
rect 670 2280 676 2281
rect 670 2276 671 2280
rect 675 2276 676 2280
rect 670 2275 676 2276
rect 806 2280 812 2281
rect 806 2276 807 2280
rect 811 2276 812 2280
rect 806 2275 812 2276
rect 942 2280 948 2281
rect 942 2276 943 2280
rect 947 2276 948 2280
rect 1934 2277 1935 2281
rect 1939 2277 1940 2281
rect 1934 2276 1940 2277
rect 942 2275 948 2276
rect 370 2265 376 2266
rect 110 2264 116 2265
rect 110 2260 111 2264
rect 115 2260 116 2264
rect 370 2261 371 2265
rect 375 2261 376 2265
rect 370 2260 376 2261
rect 506 2265 512 2266
rect 506 2261 507 2265
rect 511 2261 512 2265
rect 506 2260 512 2261
rect 642 2265 648 2266
rect 642 2261 643 2265
rect 647 2261 648 2265
rect 642 2260 648 2261
rect 778 2265 784 2266
rect 778 2261 779 2265
rect 783 2261 784 2265
rect 778 2260 784 2261
rect 914 2265 920 2266
rect 914 2261 915 2265
rect 919 2261 920 2265
rect 914 2260 920 2261
rect 1934 2264 1940 2265
rect 1934 2260 1935 2264
rect 1939 2260 1940 2264
rect 110 2259 116 2260
rect 112 2191 114 2259
rect 372 2191 374 2260
rect 508 2191 510 2260
rect 644 2191 646 2260
rect 780 2191 782 2260
rect 916 2191 918 2260
rect 1934 2259 1940 2260
rect 1936 2191 1938 2259
rect 1976 2233 1978 2293
rect 1974 2232 1980 2233
rect 2044 2232 2046 2293
rect 2180 2232 2182 2293
rect 2316 2232 2318 2293
rect 2452 2232 2454 2293
rect 2588 2232 2590 2293
rect 2724 2232 2726 2293
rect 2860 2232 2862 2293
rect 2996 2232 2998 2293
rect 3132 2232 3134 2293
rect 3800 2233 3802 2293
rect 3840 2285 3842 2345
rect 3838 2284 3844 2285
rect 4676 2284 4678 2345
rect 4820 2284 4822 2345
rect 4964 2284 4966 2345
rect 5116 2284 5118 2345
rect 5268 2284 5270 2345
rect 5420 2284 5422 2345
rect 5664 2285 5666 2345
rect 5662 2284 5668 2285
rect 3838 2280 3839 2284
rect 3843 2280 3844 2284
rect 3838 2279 3844 2280
rect 4674 2283 4680 2284
rect 4674 2279 4675 2283
rect 4679 2279 4680 2283
rect 4674 2278 4680 2279
rect 4818 2283 4824 2284
rect 4818 2279 4819 2283
rect 4823 2279 4824 2283
rect 4818 2278 4824 2279
rect 4962 2283 4968 2284
rect 4962 2279 4963 2283
rect 4967 2279 4968 2283
rect 4962 2278 4968 2279
rect 5114 2283 5120 2284
rect 5114 2279 5115 2283
rect 5119 2279 5120 2283
rect 5114 2278 5120 2279
rect 5266 2283 5272 2284
rect 5266 2279 5267 2283
rect 5271 2279 5272 2283
rect 5266 2278 5272 2279
rect 5418 2283 5424 2284
rect 5418 2279 5419 2283
rect 5423 2279 5424 2283
rect 5662 2280 5663 2284
rect 5667 2280 5668 2284
rect 5662 2279 5668 2280
rect 5418 2278 5424 2279
rect 4702 2268 4708 2269
rect 3838 2267 3844 2268
rect 3838 2263 3839 2267
rect 3843 2263 3844 2267
rect 4702 2264 4703 2268
rect 4707 2264 4708 2268
rect 4702 2263 4708 2264
rect 4846 2268 4852 2269
rect 4846 2264 4847 2268
rect 4851 2264 4852 2268
rect 4846 2263 4852 2264
rect 4990 2268 4996 2269
rect 4990 2264 4991 2268
rect 4995 2264 4996 2268
rect 4990 2263 4996 2264
rect 5142 2268 5148 2269
rect 5142 2264 5143 2268
rect 5147 2264 5148 2268
rect 5142 2263 5148 2264
rect 5294 2268 5300 2269
rect 5294 2264 5295 2268
rect 5299 2264 5300 2268
rect 5294 2263 5300 2264
rect 5446 2268 5452 2269
rect 5446 2264 5447 2268
rect 5451 2264 5452 2268
rect 5446 2263 5452 2264
rect 5662 2267 5668 2268
rect 5662 2263 5663 2267
rect 5667 2263 5668 2267
rect 3838 2262 3844 2263
rect 3798 2232 3804 2233
rect 1974 2228 1975 2232
rect 1979 2228 1980 2232
rect 1974 2227 1980 2228
rect 2042 2231 2048 2232
rect 2042 2227 2043 2231
rect 2047 2227 2048 2231
rect 2042 2226 2048 2227
rect 2178 2231 2184 2232
rect 2178 2227 2179 2231
rect 2183 2227 2184 2231
rect 2178 2226 2184 2227
rect 2314 2231 2320 2232
rect 2314 2227 2315 2231
rect 2319 2227 2320 2231
rect 2314 2226 2320 2227
rect 2450 2231 2456 2232
rect 2450 2227 2451 2231
rect 2455 2227 2456 2231
rect 2450 2226 2456 2227
rect 2586 2231 2592 2232
rect 2586 2227 2587 2231
rect 2591 2227 2592 2231
rect 2586 2226 2592 2227
rect 2722 2231 2728 2232
rect 2722 2227 2723 2231
rect 2727 2227 2728 2231
rect 2722 2226 2728 2227
rect 2858 2231 2864 2232
rect 2858 2227 2859 2231
rect 2863 2227 2864 2231
rect 2858 2226 2864 2227
rect 2994 2231 3000 2232
rect 2994 2227 2995 2231
rect 2999 2227 3000 2231
rect 2994 2226 3000 2227
rect 3130 2231 3136 2232
rect 3130 2227 3131 2231
rect 3135 2227 3136 2231
rect 3798 2228 3799 2232
rect 3803 2228 3804 2232
rect 3798 2227 3804 2228
rect 3840 2227 3842 2262
rect 4704 2227 4706 2263
rect 4848 2227 4850 2263
rect 4992 2227 4994 2263
rect 5144 2227 5146 2263
rect 5296 2227 5298 2263
rect 5448 2227 5450 2263
rect 5662 2262 5668 2263
rect 5664 2227 5666 2262
rect 3130 2226 3136 2227
rect 3839 2226 3843 2227
rect 3839 2221 3843 2222
rect 3887 2226 3891 2227
rect 3887 2221 3891 2222
rect 4167 2226 4171 2227
rect 4167 2221 4171 2222
rect 4455 2226 4459 2227
rect 4455 2221 4459 2222
rect 4703 2226 4707 2227
rect 4703 2221 4707 2222
rect 4719 2226 4723 2227
rect 4719 2221 4723 2222
rect 4847 2226 4851 2227
rect 4847 2221 4851 2222
rect 4975 2226 4979 2227
rect 4975 2221 4979 2222
rect 4991 2226 4995 2227
rect 4991 2221 4995 2222
rect 5143 2226 5147 2227
rect 5143 2221 5147 2222
rect 5231 2226 5235 2227
rect 5231 2221 5235 2222
rect 5295 2226 5299 2227
rect 5295 2221 5299 2222
rect 5447 2226 5451 2227
rect 5447 2221 5451 2222
rect 5487 2226 5491 2227
rect 5487 2221 5491 2222
rect 5663 2226 5667 2227
rect 5663 2221 5667 2222
rect 2070 2216 2076 2217
rect 1974 2215 1980 2216
rect 1974 2211 1975 2215
rect 1979 2211 1980 2215
rect 2070 2212 2071 2216
rect 2075 2212 2076 2216
rect 2070 2211 2076 2212
rect 2206 2216 2212 2217
rect 2206 2212 2207 2216
rect 2211 2212 2212 2216
rect 2206 2211 2212 2212
rect 2342 2216 2348 2217
rect 2342 2212 2343 2216
rect 2347 2212 2348 2216
rect 2342 2211 2348 2212
rect 2478 2216 2484 2217
rect 2478 2212 2479 2216
rect 2483 2212 2484 2216
rect 2478 2211 2484 2212
rect 2614 2216 2620 2217
rect 2614 2212 2615 2216
rect 2619 2212 2620 2216
rect 2614 2211 2620 2212
rect 2750 2216 2756 2217
rect 2750 2212 2751 2216
rect 2755 2212 2756 2216
rect 2750 2211 2756 2212
rect 2886 2216 2892 2217
rect 2886 2212 2887 2216
rect 2891 2212 2892 2216
rect 2886 2211 2892 2212
rect 3022 2216 3028 2217
rect 3022 2212 3023 2216
rect 3027 2212 3028 2216
rect 3022 2211 3028 2212
rect 3158 2216 3164 2217
rect 3158 2212 3159 2216
rect 3163 2212 3164 2216
rect 3158 2211 3164 2212
rect 3798 2215 3804 2216
rect 3798 2211 3799 2215
rect 3803 2211 3804 2215
rect 1974 2210 1980 2211
rect 111 2190 115 2191
rect 111 2185 115 2186
rect 323 2190 327 2191
rect 323 2185 327 2186
rect 371 2190 375 2191
rect 371 2185 375 2186
rect 459 2190 463 2191
rect 459 2185 463 2186
rect 507 2190 511 2191
rect 507 2185 511 2186
rect 595 2190 599 2191
rect 595 2185 599 2186
rect 643 2190 647 2191
rect 643 2185 647 2186
rect 731 2190 735 2191
rect 731 2185 735 2186
rect 779 2190 783 2191
rect 779 2185 783 2186
rect 867 2190 871 2191
rect 867 2185 871 2186
rect 915 2190 919 2191
rect 915 2185 919 2186
rect 1935 2190 1939 2191
rect 1976 2187 1978 2210
rect 2072 2187 2074 2211
rect 2208 2187 2210 2211
rect 2344 2187 2346 2211
rect 2480 2187 2482 2211
rect 2616 2187 2618 2211
rect 2752 2187 2754 2211
rect 2888 2187 2890 2211
rect 3024 2187 3026 2211
rect 3160 2187 3162 2211
rect 3798 2210 3804 2211
rect 3800 2187 3802 2210
rect 3840 2198 3842 2221
rect 3838 2197 3844 2198
rect 3888 2197 3890 2221
rect 4168 2197 4170 2221
rect 4456 2197 4458 2221
rect 4720 2197 4722 2221
rect 4976 2197 4978 2221
rect 5232 2197 5234 2221
rect 5488 2197 5490 2221
rect 5664 2198 5666 2221
rect 5662 2197 5668 2198
rect 3838 2193 3839 2197
rect 3843 2193 3844 2197
rect 3838 2192 3844 2193
rect 3886 2196 3892 2197
rect 3886 2192 3887 2196
rect 3891 2192 3892 2196
rect 3886 2191 3892 2192
rect 4166 2196 4172 2197
rect 4166 2192 4167 2196
rect 4171 2192 4172 2196
rect 4166 2191 4172 2192
rect 4454 2196 4460 2197
rect 4454 2192 4455 2196
rect 4459 2192 4460 2196
rect 4454 2191 4460 2192
rect 4718 2196 4724 2197
rect 4718 2192 4719 2196
rect 4723 2192 4724 2196
rect 4718 2191 4724 2192
rect 4974 2196 4980 2197
rect 4974 2192 4975 2196
rect 4979 2192 4980 2196
rect 4974 2191 4980 2192
rect 5230 2196 5236 2197
rect 5230 2192 5231 2196
rect 5235 2192 5236 2196
rect 5230 2191 5236 2192
rect 5486 2196 5492 2197
rect 5486 2192 5487 2196
rect 5491 2192 5492 2196
rect 5662 2193 5663 2197
rect 5667 2193 5668 2197
rect 5662 2192 5668 2193
rect 5486 2191 5492 2192
rect 1935 2185 1939 2186
rect 1975 2186 1979 2187
rect 112 2125 114 2185
rect 110 2124 116 2125
rect 324 2124 326 2185
rect 460 2124 462 2185
rect 596 2124 598 2185
rect 732 2124 734 2185
rect 868 2124 870 2185
rect 1936 2125 1938 2185
rect 1975 2181 1979 2182
rect 2023 2186 2027 2187
rect 2023 2181 2027 2182
rect 2071 2186 2075 2187
rect 2071 2181 2075 2182
rect 2207 2186 2211 2187
rect 2207 2181 2211 2182
rect 2239 2186 2243 2187
rect 2239 2181 2243 2182
rect 2343 2186 2347 2187
rect 2343 2181 2347 2182
rect 2479 2186 2483 2187
rect 2479 2181 2483 2182
rect 2487 2186 2491 2187
rect 2487 2181 2491 2182
rect 2615 2186 2619 2187
rect 2615 2181 2619 2182
rect 2727 2186 2731 2187
rect 2727 2181 2731 2182
rect 2751 2186 2755 2187
rect 2751 2181 2755 2182
rect 2887 2186 2891 2187
rect 2887 2181 2891 2182
rect 2967 2186 2971 2187
rect 2967 2181 2971 2182
rect 3023 2186 3027 2187
rect 3023 2181 3027 2182
rect 3159 2186 3163 2187
rect 3159 2181 3163 2182
rect 3207 2186 3211 2187
rect 3207 2181 3211 2182
rect 3455 2186 3459 2187
rect 3455 2181 3459 2182
rect 3679 2186 3683 2187
rect 3679 2181 3683 2182
rect 3799 2186 3803 2187
rect 3799 2181 3803 2182
rect 3858 2181 3864 2182
rect 1976 2158 1978 2181
rect 1974 2157 1980 2158
rect 2024 2157 2026 2181
rect 2240 2157 2242 2181
rect 2488 2157 2490 2181
rect 2728 2157 2730 2181
rect 2968 2157 2970 2181
rect 3208 2157 3210 2181
rect 3456 2157 3458 2181
rect 3680 2157 3682 2181
rect 3800 2158 3802 2181
rect 3838 2180 3844 2181
rect 3838 2176 3839 2180
rect 3843 2176 3844 2180
rect 3858 2177 3859 2181
rect 3863 2177 3864 2181
rect 3858 2176 3864 2177
rect 4138 2181 4144 2182
rect 4138 2177 4139 2181
rect 4143 2177 4144 2181
rect 4138 2176 4144 2177
rect 4426 2181 4432 2182
rect 4426 2177 4427 2181
rect 4431 2177 4432 2181
rect 4426 2176 4432 2177
rect 4690 2181 4696 2182
rect 4690 2177 4691 2181
rect 4695 2177 4696 2181
rect 4690 2176 4696 2177
rect 4946 2181 4952 2182
rect 4946 2177 4947 2181
rect 4951 2177 4952 2181
rect 4946 2176 4952 2177
rect 5202 2181 5208 2182
rect 5202 2177 5203 2181
rect 5207 2177 5208 2181
rect 5202 2176 5208 2177
rect 5458 2181 5464 2182
rect 5458 2177 5459 2181
rect 5463 2177 5464 2181
rect 5458 2176 5464 2177
rect 5662 2180 5668 2181
rect 5662 2176 5663 2180
rect 5667 2176 5668 2180
rect 3838 2175 3844 2176
rect 3798 2157 3804 2158
rect 1974 2153 1975 2157
rect 1979 2153 1980 2157
rect 1974 2152 1980 2153
rect 2022 2156 2028 2157
rect 2022 2152 2023 2156
rect 2027 2152 2028 2156
rect 2022 2151 2028 2152
rect 2238 2156 2244 2157
rect 2238 2152 2239 2156
rect 2243 2152 2244 2156
rect 2238 2151 2244 2152
rect 2486 2156 2492 2157
rect 2486 2152 2487 2156
rect 2491 2152 2492 2156
rect 2486 2151 2492 2152
rect 2726 2156 2732 2157
rect 2726 2152 2727 2156
rect 2731 2152 2732 2156
rect 2726 2151 2732 2152
rect 2966 2156 2972 2157
rect 2966 2152 2967 2156
rect 2971 2152 2972 2156
rect 2966 2151 2972 2152
rect 3206 2156 3212 2157
rect 3206 2152 3207 2156
rect 3211 2152 3212 2156
rect 3206 2151 3212 2152
rect 3454 2156 3460 2157
rect 3454 2152 3455 2156
rect 3459 2152 3460 2156
rect 3454 2151 3460 2152
rect 3678 2156 3684 2157
rect 3678 2152 3679 2156
rect 3683 2152 3684 2156
rect 3798 2153 3799 2157
rect 3803 2153 3804 2157
rect 3798 2152 3804 2153
rect 3678 2151 3684 2152
rect 1994 2141 2000 2142
rect 1974 2140 1980 2141
rect 1974 2136 1975 2140
rect 1979 2136 1980 2140
rect 1994 2137 1995 2141
rect 1999 2137 2000 2141
rect 1994 2136 2000 2137
rect 2210 2141 2216 2142
rect 2210 2137 2211 2141
rect 2215 2137 2216 2141
rect 2210 2136 2216 2137
rect 2458 2141 2464 2142
rect 2458 2137 2459 2141
rect 2463 2137 2464 2141
rect 2458 2136 2464 2137
rect 2698 2141 2704 2142
rect 2698 2137 2699 2141
rect 2703 2137 2704 2141
rect 2698 2136 2704 2137
rect 2938 2141 2944 2142
rect 2938 2137 2939 2141
rect 2943 2137 2944 2141
rect 2938 2136 2944 2137
rect 3178 2141 3184 2142
rect 3178 2137 3179 2141
rect 3183 2137 3184 2141
rect 3178 2136 3184 2137
rect 3426 2141 3432 2142
rect 3426 2137 3427 2141
rect 3431 2137 3432 2141
rect 3426 2136 3432 2137
rect 3650 2141 3656 2142
rect 3650 2137 3651 2141
rect 3655 2137 3656 2141
rect 3650 2136 3656 2137
rect 3798 2140 3804 2141
rect 3798 2136 3799 2140
rect 3803 2136 3804 2140
rect 1974 2135 1980 2136
rect 1934 2124 1940 2125
rect 110 2120 111 2124
rect 115 2120 116 2124
rect 110 2119 116 2120
rect 322 2123 328 2124
rect 322 2119 323 2123
rect 327 2119 328 2123
rect 322 2118 328 2119
rect 458 2123 464 2124
rect 458 2119 459 2123
rect 463 2119 464 2123
rect 458 2118 464 2119
rect 594 2123 600 2124
rect 594 2119 595 2123
rect 599 2119 600 2123
rect 594 2118 600 2119
rect 730 2123 736 2124
rect 730 2119 731 2123
rect 735 2119 736 2123
rect 730 2118 736 2119
rect 866 2123 872 2124
rect 866 2119 867 2123
rect 871 2119 872 2123
rect 1934 2120 1935 2124
rect 1939 2120 1940 2124
rect 1934 2119 1940 2120
rect 866 2118 872 2119
rect 350 2108 356 2109
rect 110 2107 116 2108
rect 110 2103 111 2107
rect 115 2103 116 2107
rect 350 2104 351 2108
rect 355 2104 356 2108
rect 350 2103 356 2104
rect 486 2108 492 2109
rect 486 2104 487 2108
rect 491 2104 492 2108
rect 486 2103 492 2104
rect 622 2108 628 2109
rect 622 2104 623 2108
rect 627 2104 628 2108
rect 622 2103 628 2104
rect 758 2108 764 2109
rect 758 2104 759 2108
rect 763 2104 764 2108
rect 758 2103 764 2104
rect 894 2108 900 2109
rect 894 2104 895 2108
rect 899 2104 900 2108
rect 894 2103 900 2104
rect 1934 2107 1940 2108
rect 1934 2103 1935 2107
rect 1939 2103 1940 2107
rect 110 2102 116 2103
rect 112 2047 114 2102
rect 352 2047 354 2103
rect 488 2047 490 2103
rect 624 2047 626 2103
rect 760 2047 762 2103
rect 896 2047 898 2103
rect 1934 2102 1940 2103
rect 1936 2047 1938 2102
rect 1976 2059 1978 2135
rect 1996 2059 1998 2136
rect 2212 2059 2214 2136
rect 2460 2059 2462 2136
rect 2700 2059 2702 2136
rect 2940 2059 2942 2136
rect 3180 2059 3182 2136
rect 3428 2059 3430 2136
rect 3652 2059 3654 2136
rect 3798 2135 3804 2136
rect 3800 2059 3802 2135
rect 3840 2115 3842 2175
rect 3860 2115 3862 2176
rect 4140 2115 4142 2176
rect 4428 2115 4430 2176
rect 4692 2115 4694 2176
rect 4948 2115 4950 2176
rect 5204 2115 5206 2176
rect 5460 2115 5462 2176
rect 5662 2175 5668 2176
rect 5664 2115 5666 2175
rect 3839 2114 3843 2115
rect 3839 2109 3843 2110
rect 3859 2114 3863 2115
rect 3859 2109 3863 2110
rect 4083 2114 4087 2115
rect 4083 2109 4087 2110
rect 4139 2114 4143 2115
rect 4139 2109 4143 2110
rect 4323 2114 4327 2115
rect 4323 2109 4327 2110
rect 4427 2114 4431 2115
rect 4427 2109 4431 2110
rect 4547 2114 4551 2115
rect 4547 2109 4551 2110
rect 4691 2114 4695 2115
rect 4691 2109 4695 2110
rect 4755 2114 4759 2115
rect 4755 2109 4759 2110
rect 4947 2114 4951 2115
rect 4947 2109 4951 2110
rect 5139 2114 5143 2115
rect 5139 2109 5143 2110
rect 5203 2114 5207 2115
rect 5203 2109 5207 2110
rect 5323 2114 5327 2115
rect 5323 2109 5327 2110
rect 5459 2114 5463 2115
rect 5459 2109 5463 2110
rect 5515 2114 5519 2115
rect 5515 2109 5519 2110
rect 5663 2114 5667 2115
rect 5663 2109 5667 2110
rect 1975 2058 1979 2059
rect 1975 2053 1979 2054
rect 1995 2058 1999 2059
rect 1995 2053 1999 2054
rect 2211 2058 2215 2059
rect 2211 2053 2215 2054
rect 2459 2058 2463 2059
rect 2459 2053 2463 2054
rect 2699 2058 2703 2059
rect 2699 2053 2703 2054
rect 2707 2058 2711 2059
rect 2707 2053 2711 2054
rect 2939 2058 2943 2059
rect 2939 2053 2943 2054
rect 2963 2058 2967 2059
rect 2963 2053 2967 2054
rect 3179 2058 3183 2059
rect 3179 2053 3183 2054
rect 3219 2058 3223 2059
rect 3219 2053 3223 2054
rect 3427 2058 3431 2059
rect 3427 2053 3431 2054
rect 3483 2058 3487 2059
rect 3483 2053 3487 2054
rect 3651 2058 3655 2059
rect 3651 2053 3655 2054
rect 3799 2058 3803 2059
rect 3799 2053 3803 2054
rect 111 2046 115 2047
rect 111 2041 115 2042
rect 319 2046 323 2047
rect 319 2041 323 2042
rect 351 2046 355 2047
rect 351 2041 355 2042
rect 479 2046 483 2047
rect 479 2041 483 2042
rect 487 2046 491 2047
rect 487 2041 491 2042
rect 623 2046 627 2047
rect 623 2041 627 2042
rect 663 2046 667 2047
rect 663 2041 667 2042
rect 759 2046 763 2047
rect 759 2041 763 2042
rect 871 2046 875 2047
rect 871 2041 875 2042
rect 895 2046 899 2047
rect 895 2041 899 2042
rect 1095 2046 1099 2047
rect 1095 2041 1099 2042
rect 1335 2046 1339 2047
rect 1335 2041 1339 2042
rect 1583 2046 1587 2047
rect 1583 2041 1587 2042
rect 1815 2046 1819 2047
rect 1815 2041 1819 2042
rect 1935 2046 1939 2047
rect 1935 2041 1939 2042
rect 112 2018 114 2041
rect 110 2017 116 2018
rect 320 2017 322 2041
rect 480 2017 482 2041
rect 664 2017 666 2041
rect 872 2017 874 2041
rect 1096 2017 1098 2041
rect 1336 2017 1338 2041
rect 1584 2017 1586 2041
rect 1816 2017 1818 2041
rect 1936 2018 1938 2041
rect 1934 2017 1940 2018
rect 110 2013 111 2017
rect 115 2013 116 2017
rect 110 2012 116 2013
rect 318 2016 324 2017
rect 318 2012 319 2016
rect 323 2012 324 2016
rect 318 2011 324 2012
rect 478 2016 484 2017
rect 478 2012 479 2016
rect 483 2012 484 2016
rect 478 2011 484 2012
rect 662 2016 668 2017
rect 662 2012 663 2016
rect 667 2012 668 2016
rect 662 2011 668 2012
rect 870 2016 876 2017
rect 870 2012 871 2016
rect 875 2012 876 2016
rect 870 2011 876 2012
rect 1094 2016 1100 2017
rect 1094 2012 1095 2016
rect 1099 2012 1100 2016
rect 1094 2011 1100 2012
rect 1334 2016 1340 2017
rect 1334 2012 1335 2016
rect 1339 2012 1340 2016
rect 1334 2011 1340 2012
rect 1582 2016 1588 2017
rect 1582 2012 1583 2016
rect 1587 2012 1588 2016
rect 1582 2011 1588 2012
rect 1814 2016 1820 2017
rect 1814 2012 1815 2016
rect 1819 2012 1820 2016
rect 1934 2013 1935 2017
rect 1939 2013 1940 2017
rect 1934 2012 1940 2013
rect 1814 2011 1820 2012
rect 290 2001 296 2002
rect 110 2000 116 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 290 1997 291 2001
rect 295 1997 296 2001
rect 290 1996 296 1997
rect 450 2001 456 2002
rect 450 1997 451 2001
rect 455 1997 456 2001
rect 450 1996 456 1997
rect 634 2001 640 2002
rect 634 1997 635 2001
rect 639 1997 640 2001
rect 634 1996 640 1997
rect 842 2001 848 2002
rect 842 1997 843 2001
rect 847 1997 848 2001
rect 842 1996 848 1997
rect 1066 2001 1072 2002
rect 1066 1997 1067 2001
rect 1071 1997 1072 2001
rect 1066 1996 1072 1997
rect 1306 2001 1312 2002
rect 1306 1997 1307 2001
rect 1311 1997 1312 2001
rect 1306 1996 1312 1997
rect 1554 2001 1560 2002
rect 1554 1997 1555 2001
rect 1559 1997 1560 2001
rect 1554 1996 1560 1997
rect 1786 2001 1792 2002
rect 1786 1997 1787 2001
rect 1791 1997 1792 2001
rect 1786 1996 1792 1997
rect 1934 2000 1940 2001
rect 1934 1996 1935 2000
rect 1939 1996 1940 2000
rect 110 1995 116 1996
rect 112 1927 114 1995
rect 292 1927 294 1996
rect 452 1927 454 1996
rect 636 1927 638 1996
rect 844 1927 846 1996
rect 1068 1927 1070 1996
rect 1308 1927 1310 1996
rect 1556 1927 1558 1996
rect 1788 1927 1790 1996
rect 1934 1995 1940 1996
rect 1936 1927 1938 1995
rect 1976 1993 1978 2053
rect 1974 1992 1980 1993
rect 1996 1992 1998 2053
rect 2212 1992 2214 2053
rect 2460 1992 2462 2053
rect 2708 1992 2710 2053
rect 2964 1992 2966 2053
rect 3220 1992 3222 2053
rect 3484 1992 3486 2053
rect 3800 1993 3802 2053
rect 3840 2049 3842 2109
rect 3838 2048 3844 2049
rect 3860 2048 3862 2109
rect 4084 2048 4086 2109
rect 4324 2048 4326 2109
rect 4548 2048 4550 2109
rect 4756 2048 4758 2109
rect 4948 2048 4950 2109
rect 5140 2048 5142 2109
rect 5324 2048 5326 2109
rect 5516 2048 5518 2109
rect 5664 2049 5666 2109
rect 5662 2048 5668 2049
rect 3838 2044 3839 2048
rect 3843 2044 3844 2048
rect 3838 2043 3844 2044
rect 3858 2047 3864 2048
rect 3858 2043 3859 2047
rect 3863 2043 3864 2047
rect 3858 2042 3864 2043
rect 4082 2047 4088 2048
rect 4082 2043 4083 2047
rect 4087 2043 4088 2047
rect 4082 2042 4088 2043
rect 4322 2047 4328 2048
rect 4322 2043 4323 2047
rect 4327 2043 4328 2047
rect 4322 2042 4328 2043
rect 4546 2047 4552 2048
rect 4546 2043 4547 2047
rect 4551 2043 4552 2047
rect 4546 2042 4552 2043
rect 4754 2047 4760 2048
rect 4754 2043 4755 2047
rect 4759 2043 4760 2047
rect 4754 2042 4760 2043
rect 4946 2047 4952 2048
rect 4946 2043 4947 2047
rect 4951 2043 4952 2047
rect 4946 2042 4952 2043
rect 5138 2047 5144 2048
rect 5138 2043 5139 2047
rect 5143 2043 5144 2047
rect 5138 2042 5144 2043
rect 5322 2047 5328 2048
rect 5322 2043 5323 2047
rect 5327 2043 5328 2047
rect 5322 2042 5328 2043
rect 5514 2047 5520 2048
rect 5514 2043 5515 2047
rect 5519 2043 5520 2047
rect 5662 2044 5663 2048
rect 5667 2044 5668 2048
rect 5662 2043 5668 2044
rect 5514 2042 5520 2043
rect 3886 2032 3892 2033
rect 3838 2031 3844 2032
rect 3838 2027 3839 2031
rect 3843 2027 3844 2031
rect 3886 2028 3887 2032
rect 3891 2028 3892 2032
rect 3886 2027 3892 2028
rect 4110 2032 4116 2033
rect 4110 2028 4111 2032
rect 4115 2028 4116 2032
rect 4110 2027 4116 2028
rect 4350 2032 4356 2033
rect 4350 2028 4351 2032
rect 4355 2028 4356 2032
rect 4350 2027 4356 2028
rect 4574 2032 4580 2033
rect 4574 2028 4575 2032
rect 4579 2028 4580 2032
rect 4574 2027 4580 2028
rect 4782 2032 4788 2033
rect 4782 2028 4783 2032
rect 4787 2028 4788 2032
rect 4782 2027 4788 2028
rect 4974 2032 4980 2033
rect 4974 2028 4975 2032
rect 4979 2028 4980 2032
rect 4974 2027 4980 2028
rect 5166 2032 5172 2033
rect 5166 2028 5167 2032
rect 5171 2028 5172 2032
rect 5166 2027 5172 2028
rect 5350 2032 5356 2033
rect 5350 2028 5351 2032
rect 5355 2028 5356 2032
rect 5350 2027 5356 2028
rect 5542 2032 5548 2033
rect 5542 2028 5543 2032
rect 5547 2028 5548 2032
rect 5542 2027 5548 2028
rect 5662 2031 5668 2032
rect 5662 2027 5663 2031
rect 5667 2027 5668 2031
rect 3838 2026 3844 2027
rect 3840 2003 3842 2026
rect 3888 2003 3890 2027
rect 4112 2003 4114 2027
rect 4352 2003 4354 2027
rect 4576 2003 4578 2027
rect 4784 2003 4786 2027
rect 4976 2003 4978 2027
rect 5168 2003 5170 2027
rect 5352 2003 5354 2027
rect 5544 2003 5546 2027
rect 5662 2026 5668 2027
rect 5664 2003 5666 2026
rect 3839 2002 3843 2003
rect 3839 1997 3843 1998
rect 3887 2002 3891 2003
rect 3887 1997 3891 1998
rect 4111 2002 4115 2003
rect 4111 1997 4115 1998
rect 4167 2002 4171 2003
rect 4167 1997 4171 1998
rect 4351 2002 4355 2003
rect 4351 1997 4355 1998
rect 4463 2002 4467 2003
rect 4463 1997 4467 1998
rect 4575 2002 4579 2003
rect 4575 1997 4579 1998
rect 4743 2002 4747 2003
rect 4743 1997 4747 1998
rect 4783 2002 4787 2003
rect 4783 1997 4787 1998
rect 4975 2002 4979 2003
rect 4975 1997 4979 1998
rect 5007 2002 5011 2003
rect 5007 1997 5011 1998
rect 5167 2002 5171 2003
rect 5167 1997 5171 1998
rect 5271 2002 5275 2003
rect 5271 1997 5275 1998
rect 5351 2002 5355 2003
rect 5351 1997 5355 1998
rect 5543 2002 5547 2003
rect 5543 1997 5547 1998
rect 5663 2002 5667 2003
rect 5663 1997 5667 1998
rect 3798 1992 3804 1993
rect 1974 1988 1975 1992
rect 1979 1988 1980 1992
rect 1974 1987 1980 1988
rect 1994 1991 2000 1992
rect 1994 1987 1995 1991
rect 1999 1987 2000 1991
rect 1994 1986 2000 1987
rect 2210 1991 2216 1992
rect 2210 1987 2211 1991
rect 2215 1987 2216 1991
rect 2210 1986 2216 1987
rect 2458 1991 2464 1992
rect 2458 1987 2459 1991
rect 2463 1987 2464 1991
rect 2458 1986 2464 1987
rect 2706 1991 2712 1992
rect 2706 1987 2707 1991
rect 2711 1987 2712 1991
rect 2706 1986 2712 1987
rect 2962 1991 2968 1992
rect 2962 1987 2963 1991
rect 2967 1987 2968 1991
rect 2962 1986 2968 1987
rect 3218 1991 3224 1992
rect 3218 1987 3219 1991
rect 3223 1987 3224 1991
rect 3218 1986 3224 1987
rect 3482 1991 3488 1992
rect 3482 1987 3483 1991
rect 3487 1987 3488 1991
rect 3798 1988 3799 1992
rect 3803 1988 3804 1992
rect 3798 1987 3804 1988
rect 3482 1986 3488 1987
rect 2022 1976 2028 1977
rect 1974 1975 1980 1976
rect 1974 1971 1975 1975
rect 1979 1971 1980 1975
rect 2022 1972 2023 1976
rect 2027 1972 2028 1976
rect 2022 1971 2028 1972
rect 2238 1976 2244 1977
rect 2238 1972 2239 1976
rect 2243 1972 2244 1976
rect 2238 1971 2244 1972
rect 2486 1976 2492 1977
rect 2486 1972 2487 1976
rect 2491 1972 2492 1976
rect 2486 1971 2492 1972
rect 2734 1976 2740 1977
rect 2734 1972 2735 1976
rect 2739 1972 2740 1976
rect 2734 1971 2740 1972
rect 2990 1976 2996 1977
rect 2990 1972 2991 1976
rect 2995 1972 2996 1976
rect 2990 1971 2996 1972
rect 3246 1976 3252 1977
rect 3246 1972 3247 1976
rect 3251 1972 3252 1976
rect 3246 1971 3252 1972
rect 3510 1976 3516 1977
rect 3510 1972 3511 1976
rect 3515 1972 3516 1976
rect 3510 1971 3516 1972
rect 3798 1975 3804 1976
rect 3798 1971 3799 1975
rect 3803 1971 3804 1975
rect 3840 1974 3842 1997
rect 1974 1970 1980 1971
rect 1976 1939 1978 1970
rect 2024 1939 2026 1971
rect 2240 1939 2242 1971
rect 2488 1939 2490 1971
rect 2736 1939 2738 1971
rect 2992 1939 2994 1971
rect 3248 1939 3250 1971
rect 3512 1939 3514 1971
rect 3798 1970 3804 1971
rect 3838 1973 3844 1974
rect 3888 1973 3890 1997
rect 4168 1973 4170 1997
rect 4464 1973 4466 1997
rect 4744 1973 4746 1997
rect 5008 1973 5010 1997
rect 5272 1973 5274 1997
rect 5544 1973 5546 1997
rect 5664 1974 5666 1997
rect 5662 1973 5668 1974
rect 3800 1939 3802 1970
rect 3838 1969 3839 1973
rect 3843 1969 3844 1973
rect 3838 1968 3844 1969
rect 3886 1972 3892 1973
rect 3886 1968 3887 1972
rect 3891 1968 3892 1972
rect 3886 1967 3892 1968
rect 4166 1972 4172 1973
rect 4166 1968 4167 1972
rect 4171 1968 4172 1972
rect 4166 1967 4172 1968
rect 4462 1972 4468 1973
rect 4462 1968 4463 1972
rect 4467 1968 4468 1972
rect 4462 1967 4468 1968
rect 4742 1972 4748 1973
rect 4742 1968 4743 1972
rect 4747 1968 4748 1972
rect 4742 1967 4748 1968
rect 5006 1972 5012 1973
rect 5006 1968 5007 1972
rect 5011 1968 5012 1972
rect 5006 1967 5012 1968
rect 5270 1972 5276 1973
rect 5270 1968 5271 1972
rect 5275 1968 5276 1972
rect 5270 1967 5276 1968
rect 5542 1972 5548 1973
rect 5542 1968 5543 1972
rect 5547 1968 5548 1972
rect 5662 1969 5663 1973
rect 5667 1969 5668 1973
rect 5662 1968 5668 1969
rect 5542 1967 5548 1968
rect 3858 1957 3864 1958
rect 3838 1956 3844 1957
rect 3838 1952 3839 1956
rect 3843 1952 3844 1956
rect 3858 1953 3859 1957
rect 3863 1953 3864 1957
rect 3858 1952 3864 1953
rect 4138 1957 4144 1958
rect 4138 1953 4139 1957
rect 4143 1953 4144 1957
rect 4138 1952 4144 1953
rect 4434 1957 4440 1958
rect 4434 1953 4435 1957
rect 4439 1953 4440 1957
rect 4434 1952 4440 1953
rect 4714 1957 4720 1958
rect 4714 1953 4715 1957
rect 4719 1953 4720 1957
rect 4714 1952 4720 1953
rect 4978 1957 4984 1958
rect 4978 1953 4979 1957
rect 4983 1953 4984 1957
rect 4978 1952 4984 1953
rect 5242 1957 5248 1958
rect 5242 1953 5243 1957
rect 5247 1953 5248 1957
rect 5242 1952 5248 1953
rect 5514 1957 5520 1958
rect 5514 1953 5515 1957
rect 5519 1953 5520 1957
rect 5514 1952 5520 1953
rect 5662 1956 5668 1957
rect 5662 1952 5663 1956
rect 5667 1952 5668 1956
rect 3838 1951 3844 1952
rect 1975 1938 1979 1939
rect 1975 1933 1979 1934
rect 2023 1938 2027 1939
rect 2023 1933 2027 1934
rect 2159 1938 2163 1939
rect 2159 1933 2163 1934
rect 2239 1938 2243 1939
rect 2239 1933 2243 1934
rect 2439 1938 2443 1939
rect 2439 1933 2443 1934
rect 2487 1938 2491 1939
rect 2487 1933 2491 1934
rect 2703 1938 2707 1939
rect 2703 1933 2707 1934
rect 2735 1938 2739 1939
rect 2735 1933 2739 1934
rect 2959 1938 2963 1939
rect 2959 1933 2963 1934
rect 2991 1938 2995 1939
rect 2991 1933 2995 1934
rect 3207 1938 3211 1939
rect 3207 1933 3211 1934
rect 3247 1938 3251 1939
rect 3247 1933 3251 1934
rect 3455 1938 3459 1939
rect 3455 1933 3459 1934
rect 3511 1938 3515 1939
rect 3511 1933 3515 1934
rect 3679 1938 3683 1939
rect 3679 1933 3683 1934
rect 3799 1938 3803 1939
rect 3799 1933 3803 1934
rect 111 1926 115 1927
rect 111 1921 115 1922
rect 187 1926 191 1927
rect 187 1921 191 1922
rect 291 1926 295 1927
rect 291 1921 295 1922
rect 419 1926 423 1927
rect 419 1921 423 1922
rect 451 1926 455 1927
rect 451 1921 455 1922
rect 635 1926 639 1927
rect 635 1921 639 1922
rect 651 1926 655 1927
rect 651 1921 655 1922
rect 843 1926 847 1927
rect 843 1921 847 1922
rect 883 1926 887 1927
rect 883 1921 887 1922
rect 1067 1926 1071 1927
rect 1067 1921 1071 1922
rect 1115 1926 1119 1927
rect 1115 1921 1119 1922
rect 1307 1926 1311 1927
rect 1307 1921 1311 1922
rect 1347 1926 1351 1927
rect 1347 1921 1351 1922
rect 1555 1926 1559 1927
rect 1555 1921 1559 1922
rect 1579 1926 1583 1927
rect 1579 1921 1583 1922
rect 1787 1926 1791 1927
rect 1787 1921 1791 1922
rect 1935 1926 1939 1927
rect 1935 1921 1939 1922
rect 112 1861 114 1921
rect 110 1860 116 1861
rect 188 1860 190 1921
rect 420 1860 422 1921
rect 652 1860 654 1921
rect 884 1860 886 1921
rect 1116 1860 1118 1921
rect 1348 1860 1350 1921
rect 1580 1860 1582 1921
rect 1788 1860 1790 1921
rect 1936 1861 1938 1921
rect 1976 1910 1978 1933
rect 1974 1909 1980 1910
rect 2160 1909 2162 1933
rect 2440 1909 2442 1933
rect 2704 1909 2706 1933
rect 2960 1909 2962 1933
rect 3208 1909 3210 1933
rect 3456 1909 3458 1933
rect 3680 1909 3682 1933
rect 3800 1910 3802 1933
rect 3798 1909 3804 1910
rect 1974 1905 1975 1909
rect 1979 1905 1980 1909
rect 1974 1904 1980 1905
rect 2158 1908 2164 1909
rect 2158 1904 2159 1908
rect 2163 1904 2164 1908
rect 2158 1903 2164 1904
rect 2438 1908 2444 1909
rect 2438 1904 2439 1908
rect 2443 1904 2444 1908
rect 2438 1903 2444 1904
rect 2702 1908 2708 1909
rect 2702 1904 2703 1908
rect 2707 1904 2708 1908
rect 2702 1903 2708 1904
rect 2958 1908 2964 1909
rect 2958 1904 2959 1908
rect 2963 1904 2964 1908
rect 2958 1903 2964 1904
rect 3206 1908 3212 1909
rect 3206 1904 3207 1908
rect 3211 1904 3212 1908
rect 3206 1903 3212 1904
rect 3454 1908 3460 1909
rect 3454 1904 3455 1908
rect 3459 1904 3460 1908
rect 3454 1903 3460 1904
rect 3678 1908 3684 1909
rect 3678 1904 3679 1908
rect 3683 1904 3684 1908
rect 3798 1905 3799 1909
rect 3803 1905 3804 1909
rect 3798 1904 3804 1905
rect 3678 1903 3684 1904
rect 2130 1893 2136 1894
rect 1974 1892 1980 1893
rect 1974 1888 1975 1892
rect 1979 1888 1980 1892
rect 2130 1889 2131 1893
rect 2135 1889 2136 1893
rect 2130 1888 2136 1889
rect 2410 1893 2416 1894
rect 2410 1889 2411 1893
rect 2415 1889 2416 1893
rect 2410 1888 2416 1889
rect 2674 1893 2680 1894
rect 2674 1889 2675 1893
rect 2679 1889 2680 1893
rect 2674 1888 2680 1889
rect 2930 1893 2936 1894
rect 2930 1889 2931 1893
rect 2935 1889 2936 1893
rect 2930 1888 2936 1889
rect 3178 1893 3184 1894
rect 3178 1889 3179 1893
rect 3183 1889 3184 1893
rect 3178 1888 3184 1889
rect 3426 1893 3432 1894
rect 3426 1889 3427 1893
rect 3431 1889 3432 1893
rect 3426 1888 3432 1889
rect 3650 1893 3656 1894
rect 3650 1889 3651 1893
rect 3655 1889 3656 1893
rect 3650 1888 3656 1889
rect 3798 1892 3804 1893
rect 3798 1888 3799 1892
rect 3803 1888 3804 1892
rect 1974 1887 1980 1888
rect 1934 1860 1940 1861
rect 110 1856 111 1860
rect 115 1856 116 1860
rect 110 1855 116 1856
rect 186 1859 192 1860
rect 186 1855 187 1859
rect 191 1855 192 1859
rect 186 1854 192 1855
rect 418 1859 424 1860
rect 418 1855 419 1859
rect 423 1855 424 1859
rect 418 1854 424 1855
rect 650 1859 656 1860
rect 650 1855 651 1859
rect 655 1855 656 1859
rect 650 1854 656 1855
rect 882 1859 888 1860
rect 882 1855 883 1859
rect 887 1855 888 1859
rect 882 1854 888 1855
rect 1114 1859 1120 1860
rect 1114 1855 1115 1859
rect 1119 1855 1120 1859
rect 1114 1854 1120 1855
rect 1346 1859 1352 1860
rect 1346 1855 1347 1859
rect 1351 1855 1352 1859
rect 1346 1854 1352 1855
rect 1578 1859 1584 1860
rect 1578 1855 1579 1859
rect 1583 1855 1584 1859
rect 1578 1854 1584 1855
rect 1786 1859 1792 1860
rect 1786 1855 1787 1859
rect 1791 1855 1792 1859
rect 1934 1856 1935 1860
rect 1939 1856 1940 1860
rect 1934 1855 1940 1856
rect 1786 1854 1792 1855
rect 214 1844 220 1845
rect 110 1843 116 1844
rect 110 1839 111 1843
rect 115 1839 116 1843
rect 214 1840 215 1844
rect 219 1840 220 1844
rect 214 1839 220 1840
rect 446 1844 452 1845
rect 446 1840 447 1844
rect 451 1840 452 1844
rect 446 1839 452 1840
rect 678 1844 684 1845
rect 678 1840 679 1844
rect 683 1840 684 1844
rect 678 1839 684 1840
rect 910 1844 916 1845
rect 910 1840 911 1844
rect 915 1840 916 1844
rect 910 1839 916 1840
rect 1142 1844 1148 1845
rect 1142 1840 1143 1844
rect 1147 1840 1148 1844
rect 1142 1839 1148 1840
rect 1374 1844 1380 1845
rect 1374 1840 1375 1844
rect 1379 1840 1380 1844
rect 1374 1839 1380 1840
rect 1606 1844 1612 1845
rect 1606 1840 1607 1844
rect 1611 1840 1612 1844
rect 1606 1839 1612 1840
rect 1814 1844 1820 1845
rect 1814 1840 1815 1844
rect 1819 1840 1820 1844
rect 1814 1839 1820 1840
rect 1934 1843 1940 1844
rect 1934 1839 1935 1843
rect 1939 1839 1940 1843
rect 110 1838 116 1839
rect 112 1803 114 1838
rect 216 1803 218 1839
rect 448 1803 450 1839
rect 680 1803 682 1839
rect 912 1803 914 1839
rect 1144 1803 1146 1839
rect 1376 1803 1378 1839
rect 1608 1803 1610 1839
rect 1816 1803 1818 1839
rect 1934 1838 1940 1839
rect 1936 1803 1938 1838
rect 1976 1819 1978 1887
rect 2132 1819 2134 1888
rect 2412 1819 2414 1888
rect 2676 1819 2678 1888
rect 2932 1819 2934 1888
rect 3180 1819 3182 1888
rect 3428 1819 3430 1888
rect 3652 1819 3654 1888
rect 3798 1887 3804 1888
rect 3800 1819 3802 1887
rect 3840 1879 3842 1951
rect 3860 1879 3862 1952
rect 4140 1879 4142 1952
rect 4436 1879 4438 1952
rect 4716 1879 4718 1952
rect 4980 1879 4982 1952
rect 5244 1879 5246 1952
rect 5516 1879 5518 1952
rect 5662 1951 5668 1952
rect 5664 1879 5666 1951
rect 3839 1878 3843 1879
rect 3839 1873 3843 1874
rect 3859 1878 3863 1879
rect 3859 1873 3863 1874
rect 4139 1878 4143 1879
rect 4139 1873 4143 1874
rect 4435 1878 4439 1879
rect 4435 1873 4439 1874
rect 4539 1878 4543 1879
rect 4539 1873 4543 1874
rect 4715 1878 4719 1879
rect 4715 1873 4719 1874
rect 4723 1878 4727 1879
rect 4723 1873 4727 1874
rect 4915 1878 4919 1879
rect 4915 1873 4919 1874
rect 4979 1878 4983 1879
rect 4979 1873 4983 1874
rect 5115 1878 5119 1879
rect 5115 1873 5119 1874
rect 5243 1878 5247 1879
rect 5243 1873 5247 1874
rect 5323 1878 5327 1879
rect 5323 1873 5327 1874
rect 5515 1878 5519 1879
rect 5515 1873 5519 1874
rect 5663 1878 5667 1879
rect 5663 1873 5667 1874
rect 1975 1818 1979 1819
rect 1975 1813 1979 1814
rect 2131 1818 2135 1819
rect 2131 1813 2135 1814
rect 2307 1818 2311 1819
rect 2307 1813 2311 1814
rect 2411 1818 2415 1819
rect 2411 1813 2415 1814
rect 2499 1818 2503 1819
rect 2499 1813 2503 1814
rect 2675 1818 2679 1819
rect 2675 1813 2679 1814
rect 2691 1818 2695 1819
rect 2691 1813 2695 1814
rect 2883 1818 2887 1819
rect 2883 1813 2887 1814
rect 2931 1818 2935 1819
rect 2931 1813 2935 1814
rect 3067 1818 3071 1819
rect 3067 1813 3071 1814
rect 3179 1818 3183 1819
rect 3179 1813 3183 1814
rect 3251 1818 3255 1819
rect 3251 1813 3255 1814
rect 3427 1818 3431 1819
rect 3427 1813 3431 1814
rect 3443 1818 3447 1819
rect 3443 1813 3447 1814
rect 3635 1818 3639 1819
rect 3635 1813 3639 1814
rect 3651 1818 3655 1819
rect 3651 1813 3655 1814
rect 3799 1818 3803 1819
rect 3799 1813 3803 1814
rect 3840 1813 3842 1873
rect 111 1802 115 1803
rect 111 1797 115 1798
rect 159 1802 163 1803
rect 159 1797 163 1798
rect 215 1802 219 1803
rect 215 1797 219 1798
rect 367 1802 371 1803
rect 367 1797 371 1798
rect 447 1802 451 1803
rect 447 1797 451 1798
rect 591 1802 595 1803
rect 591 1797 595 1798
rect 679 1802 683 1803
rect 679 1797 683 1798
rect 799 1802 803 1803
rect 799 1797 803 1798
rect 911 1802 915 1803
rect 911 1797 915 1798
rect 999 1802 1003 1803
rect 999 1797 1003 1798
rect 1143 1802 1147 1803
rect 1143 1797 1147 1798
rect 1191 1802 1195 1803
rect 1191 1797 1195 1798
rect 1375 1802 1379 1803
rect 1375 1797 1379 1798
rect 1559 1802 1563 1803
rect 1559 1797 1563 1798
rect 1607 1802 1611 1803
rect 1607 1797 1611 1798
rect 1751 1802 1755 1803
rect 1751 1797 1755 1798
rect 1815 1802 1819 1803
rect 1815 1797 1819 1798
rect 1935 1802 1939 1803
rect 1935 1797 1939 1798
rect 112 1774 114 1797
rect 110 1773 116 1774
rect 160 1773 162 1797
rect 368 1773 370 1797
rect 592 1773 594 1797
rect 800 1773 802 1797
rect 1000 1773 1002 1797
rect 1192 1773 1194 1797
rect 1376 1773 1378 1797
rect 1560 1773 1562 1797
rect 1752 1773 1754 1797
rect 1936 1774 1938 1797
rect 1934 1773 1940 1774
rect 110 1769 111 1773
rect 115 1769 116 1773
rect 110 1768 116 1769
rect 158 1772 164 1773
rect 158 1768 159 1772
rect 163 1768 164 1772
rect 158 1767 164 1768
rect 366 1772 372 1773
rect 366 1768 367 1772
rect 371 1768 372 1772
rect 366 1767 372 1768
rect 590 1772 596 1773
rect 590 1768 591 1772
rect 595 1768 596 1772
rect 590 1767 596 1768
rect 798 1772 804 1773
rect 798 1768 799 1772
rect 803 1768 804 1772
rect 798 1767 804 1768
rect 998 1772 1004 1773
rect 998 1768 999 1772
rect 1003 1768 1004 1772
rect 998 1767 1004 1768
rect 1190 1772 1196 1773
rect 1190 1768 1191 1772
rect 1195 1768 1196 1772
rect 1190 1767 1196 1768
rect 1374 1772 1380 1773
rect 1374 1768 1375 1772
rect 1379 1768 1380 1772
rect 1374 1767 1380 1768
rect 1558 1772 1564 1773
rect 1558 1768 1559 1772
rect 1563 1768 1564 1772
rect 1558 1767 1564 1768
rect 1750 1772 1756 1773
rect 1750 1768 1751 1772
rect 1755 1768 1756 1772
rect 1934 1769 1935 1773
rect 1939 1769 1940 1773
rect 1934 1768 1940 1769
rect 1750 1767 1756 1768
rect 130 1757 136 1758
rect 110 1756 116 1757
rect 110 1752 111 1756
rect 115 1752 116 1756
rect 130 1753 131 1757
rect 135 1753 136 1757
rect 130 1752 136 1753
rect 338 1757 344 1758
rect 338 1753 339 1757
rect 343 1753 344 1757
rect 338 1752 344 1753
rect 562 1757 568 1758
rect 562 1753 563 1757
rect 567 1753 568 1757
rect 562 1752 568 1753
rect 770 1757 776 1758
rect 770 1753 771 1757
rect 775 1753 776 1757
rect 770 1752 776 1753
rect 970 1757 976 1758
rect 970 1753 971 1757
rect 975 1753 976 1757
rect 970 1752 976 1753
rect 1162 1757 1168 1758
rect 1162 1753 1163 1757
rect 1167 1753 1168 1757
rect 1162 1752 1168 1753
rect 1346 1757 1352 1758
rect 1346 1753 1347 1757
rect 1351 1753 1352 1757
rect 1346 1752 1352 1753
rect 1530 1757 1536 1758
rect 1530 1753 1531 1757
rect 1535 1753 1536 1757
rect 1530 1752 1536 1753
rect 1722 1757 1728 1758
rect 1722 1753 1723 1757
rect 1727 1753 1728 1757
rect 1722 1752 1728 1753
rect 1934 1756 1940 1757
rect 1934 1752 1935 1756
rect 1939 1752 1940 1756
rect 1976 1753 1978 1813
rect 110 1751 116 1752
rect 112 1683 114 1751
rect 132 1683 134 1752
rect 340 1683 342 1752
rect 564 1683 566 1752
rect 772 1683 774 1752
rect 972 1683 974 1752
rect 1164 1683 1166 1752
rect 1348 1683 1350 1752
rect 1532 1683 1534 1752
rect 1724 1683 1726 1752
rect 1934 1751 1940 1752
rect 1974 1752 1980 1753
rect 2308 1752 2310 1813
rect 2500 1752 2502 1813
rect 2692 1752 2694 1813
rect 2884 1752 2886 1813
rect 3068 1752 3070 1813
rect 3252 1752 3254 1813
rect 3444 1752 3446 1813
rect 3636 1752 3638 1813
rect 3800 1753 3802 1813
rect 3838 1812 3844 1813
rect 4540 1812 4542 1873
rect 4724 1812 4726 1873
rect 4916 1812 4918 1873
rect 5116 1812 5118 1873
rect 5324 1812 5326 1873
rect 5516 1812 5518 1873
rect 5664 1813 5666 1873
rect 5662 1812 5668 1813
rect 3838 1808 3839 1812
rect 3843 1808 3844 1812
rect 3838 1807 3844 1808
rect 4538 1811 4544 1812
rect 4538 1807 4539 1811
rect 4543 1807 4544 1811
rect 4538 1806 4544 1807
rect 4722 1811 4728 1812
rect 4722 1807 4723 1811
rect 4727 1807 4728 1811
rect 4722 1806 4728 1807
rect 4914 1811 4920 1812
rect 4914 1807 4915 1811
rect 4919 1807 4920 1811
rect 4914 1806 4920 1807
rect 5114 1811 5120 1812
rect 5114 1807 5115 1811
rect 5119 1807 5120 1811
rect 5114 1806 5120 1807
rect 5322 1811 5328 1812
rect 5322 1807 5323 1811
rect 5327 1807 5328 1811
rect 5322 1806 5328 1807
rect 5514 1811 5520 1812
rect 5514 1807 5515 1811
rect 5519 1807 5520 1811
rect 5662 1808 5663 1812
rect 5667 1808 5668 1812
rect 5662 1807 5668 1808
rect 5514 1806 5520 1807
rect 4566 1796 4572 1797
rect 3838 1795 3844 1796
rect 3838 1791 3839 1795
rect 3843 1791 3844 1795
rect 4566 1792 4567 1796
rect 4571 1792 4572 1796
rect 4566 1791 4572 1792
rect 4750 1796 4756 1797
rect 4750 1792 4751 1796
rect 4755 1792 4756 1796
rect 4750 1791 4756 1792
rect 4942 1796 4948 1797
rect 4942 1792 4943 1796
rect 4947 1792 4948 1796
rect 4942 1791 4948 1792
rect 5142 1796 5148 1797
rect 5142 1792 5143 1796
rect 5147 1792 5148 1796
rect 5142 1791 5148 1792
rect 5350 1796 5356 1797
rect 5350 1792 5351 1796
rect 5355 1792 5356 1796
rect 5350 1791 5356 1792
rect 5542 1796 5548 1797
rect 5542 1792 5543 1796
rect 5547 1792 5548 1796
rect 5542 1791 5548 1792
rect 5662 1795 5668 1796
rect 5662 1791 5663 1795
rect 5667 1791 5668 1795
rect 3838 1790 3844 1791
rect 3840 1759 3842 1790
rect 4568 1759 4570 1791
rect 4752 1759 4754 1791
rect 4944 1759 4946 1791
rect 5144 1759 5146 1791
rect 5352 1759 5354 1791
rect 5544 1759 5546 1791
rect 5662 1790 5668 1791
rect 5664 1759 5666 1790
rect 3839 1758 3843 1759
rect 3839 1753 3843 1754
rect 4383 1758 4387 1759
rect 4383 1753 4387 1754
rect 4567 1758 4571 1759
rect 4567 1753 4571 1754
rect 4599 1758 4603 1759
rect 4599 1753 4603 1754
rect 4751 1758 4755 1759
rect 4751 1753 4755 1754
rect 4831 1758 4835 1759
rect 4831 1753 4835 1754
rect 4943 1758 4947 1759
rect 4943 1753 4947 1754
rect 5071 1758 5075 1759
rect 5071 1753 5075 1754
rect 5143 1758 5147 1759
rect 5143 1753 5147 1754
rect 5319 1758 5323 1759
rect 5319 1753 5323 1754
rect 5351 1758 5355 1759
rect 5351 1753 5355 1754
rect 5543 1758 5547 1759
rect 5543 1753 5547 1754
rect 5663 1758 5667 1759
rect 5663 1753 5667 1754
rect 3798 1752 3804 1753
rect 1936 1683 1938 1751
rect 1974 1748 1975 1752
rect 1979 1748 1980 1752
rect 1974 1747 1980 1748
rect 2306 1751 2312 1752
rect 2306 1747 2307 1751
rect 2311 1747 2312 1751
rect 2306 1746 2312 1747
rect 2498 1751 2504 1752
rect 2498 1747 2499 1751
rect 2503 1747 2504 1751
rect 2498 1746 2504 1747
rect 2690 1751 2696 1752
rect 2690 1747 2691 1751
rect 2695 1747 2696 1751
rect 2690 1746 2696 1747
rect 2882 1751 2888 1752
rect 2882 1747 2883 1751
rect 2887 1747 2888 1751
rect 2882 1746 2888 1747
rect 3066 1751 3072 1752
rect 3066 1747 3067 1751
rect 3071 1747 3072 1751
rect 3066 1746 3072 1747
rect 3250 1751 3256 1752
rect 3250 1747 3251 1751
rect 3255 1747 3256 1751
rect 3250 1746 3256 1747
rect 3442 1751 3448 1752
rect 3442 1747 3443 1751
rect 3447 1747 3448 1751
rect 3442 1746 3448 1747
rect 3634 1751 3640 1752
rect 3634 1747 3635 1751
rect 3639 1747 3640 1751
rect 3798 1748 3799 1752
rect 3803 1748 3804 1752
rect 3798 1747 3804 1748
rect 3634 1746 3640 1747
rect 2334 1736 2340 1737
rect 1974 1735 1980 1736
rect 1974 1731 1975 1735
rect 1979 1731 1980 1735
rect 2334 1732 2335 1736
rect 2339 1732 2340 1736
rect 2334 1731 2340 1732
rect 2526 1736 2532 1737
rect 2526 1732 2527 1736
rect 2531 1732 2532 1736
rect 2526 1731 2532 1732
rect 2718 1736 2724 1737
rect 2718 1732 2719 1736
rect 2723 1732 2724 1736
rect 2718 1731 2724 1732
rect 2910 1736 2916 1737
rect 2910 1732 2911 1736
rect 2915 1732 2916 1736
rect 2910 1731 2916 1732
rect 3094 1736 3100 1737
rect 3094 1732 3095 1736
rect 3099 1732 3100 1736
rect 3094 1731 3100 1732
rect 3278 1736 3284 1737
rect 3278 1732 3279 1736
rect 3283 1732 3284 1736
rect 3278 1731 3284 1732
rect 3470 1736 3476 1737
rect 3470 1732 3471 1736
rect 3475 1732 3476 1736
rect 3470 1731 3476 1732
rect 3662 1736 3668 1737
rect 3662 1732 3663 1736
rect 3667 1732 3668 1736
rect 3662 1731 3668 1732
rect 3798 1735 3804 1736
rect 3798 1731 3799 1735
rect 3803 1731 3804 1735
rect 1974 1730 1980 1731
rect 1976 1707 1978 1730
rect 2336 1707 2338 1731
rect 2528 1707 2530 1731
rect 2720 1707 2722 1731
rect 2912 1707 2914 1731
rect 3096 1707 3098 1731
rect 3280 1707 3282 1731
rect 3472 1707 3474 1731
rect 3664 1707 3666 1731
rect 3798 1730 3804 1731
rect 3840 1730 3842 1753
rect 3800 1707 3802 1730
rect 3838 1729 3844 1730
rect 4384 1729 4386 1753
rect 4600 1729 4602 1753
rect 4832 1729 4834 1753
rect 5072 1729 5074 1753
rect 5320 1729 5322 1753
rect 5544 1729 5546 1753
rect 5664 1730 5666 1753
rect 5662 1729 5668 1730
rect 3838 1725 3839 1729
rect 3843 1725 3844 1729
rect 3838 1724 3844 1725
rect 4382 1728 4388 1729
rect 4382 1724 4383 1728
rect 4387 1724 4388 1728
rect 4382 1723 4388 1724
rect 4598 1728 4604 1729
rect 4598 1724 4599 1728
rect 4603 1724 4604 1728
rect 4598 1723 4604 1724
rect 4830 1728 4836 1729
rect 4830 1724 4831 1728
rect 4835 1724 4836 1728
rect 4830 1723 4836 1724
rect 5070 1728 5076 1729
rect 5070 1724 5071 1728
rect 5075 1724 5076 1728
rect 5070 1723 5076 1724
rect 5318 1728 5324 1729
rect 5318 1724 5319 1728
rect 5323 1724 5324 1728
rect 5318 1723 5324 1724
rect 5542 1728 5548 1729
rect 5542 1724 5543 1728
rect 5547 1724 5548 1728
rect 5662 1725 5663 1729
rect 5667 1725 5668 1729
rect 5662 1724 5668 1725
rect 5542 1723 5548 1724
rect 4354 1713 4360 1714
rect 3838 1712 3844 1713
rect 3838 1708 3839 1712
rect 3843 1708 3844 1712
rect 4354 1709 4355 1713
rect 4359 1709 4360 1713
rect 4354 1708 4360 1709
rect 4570 1713 4576 1714
rect 4570 1709 4571 1713
rect 4575 1709 4576 1713
rect 4570 1708 4576 1709
rect 4802 1713 4808 1714
rect 4802 1709 4803 1713
rect 4807 1709 4808 1713
rect 4802 1708 4808 1709
rect 5042 1713 5048 1714
rect 5042 1709 5043 1713
rect 5047 1709 5048 1713
rect 5042 1708 5048 1709
rect 5290 1713 5296 1714
rect 5290 1709 5291 1713
rect 5295 1709 5296 1713
rect 5290 1708 5296 1709
rect 5514 1713 5520 1714
rect 5514 1709 5515 1713
rect 5519 1709 5520 1713
rect 5514 1708 5520 1709
rect 5662 1712 5668 1713
rect 5662 1708 5663 1712
rect 5667 1708 5668 1712
rect 3838 1707 3844 1708
rect 1975 1706 1979 1707
rect 1975 1701 1979 1702
rect 2335 1706 2339 1707
rect 2335 1701 2339 1702
rect 2471 1706 2475 1707
rect 2471 1701 2475 1702
rect 2527 1706 2531 1707
rect 2527 1701 2531 1702
rect 2607 1706 2611 1707
rect 2607 1701 2611 1702
rect 2719 1706 2723 1707
rect 2719 1701 2723 1702
rect 2743 1706 2747 1707
rect 2743 1701 2747 1702
rect 2879 1706 2883 1707
rect 2879 1701 2883 1702
rect 2911 1706 2915 1707
rect 2911 1701 2915 1702
rect 3023 1706 3027 1707
rect 3023 1701 3027 1702
rect 3095 1706 3099 1707
rect 3095 1701 3099 1702
rect 3175 1706 3179 1707
rect 3175 1701 3179 1702
rect 3279 1706 3283 1707
rect 3279 1701 3283 1702
rect 3327 1706 3331 1707
rect 3327 1701 3331 1702
rect 3471 1706 3475 1707
rect 3471 1701 3475 1702
rect 3663 1706 3667 1707
rect 3663 1701 3667 1702
rect 3799 1706 3803 1707
rect 3799 1701 3803 1702
rect 111 1682 115 1683
rect 111 1677 115 1678
rect 131 1682 135 1683
rect 131 1677 135 1678
rect 339 1682 343 1683
rect 339 1677 343 1678
rect 355 1682 359 1683
rect 355 1677 359 1678
rect 563 1682 567 1683
rect 563 1677 567 1678
rect 595 1682 599 1683
rect 595 1677 599 1678
rect 771 1682 775 1683
rect 771 1677 775 1678
rect 835 1682 839 1683
rect 835 1677 839 1678
rect 971 1682 975 1683
rect 971 1677 975 1678
rect 1067 1682 1071 1683
rect 1067 1677 1071 1678
rect 1163 1682 1167 1683
rect 1163 1677 1167 1678
rect 1307 1682 1311 1683
rect 1307 1677 1311 1678
rect 1347 1682 1351 1683
rect 1347 1677 1351 1678
rect 1531 1682 1535 1683
rect 1531 1677 1535 1678
rect 1547 1682 1551 1683
rect 1547 1677 1551 1678
rect 1723 1682 1727 1683
rect 1723 1677 1727 1678
rect 1935 1682 1939 1683
rect 1976 1678 1978 1701
rect 1935 1677 1939 1678
rect 1974 1677 1980 1678
rect 2472 1677 2474 1701
rect 2608 1677 2610 1701
rect 2744 1677 2746 1701
rect 2880 1677 2882 1701
rect 3024 1677 3026 1701
rect 3176 1677 3178 1701
rect 3328 1677 3330 1701
rect 3800 1678 3802 1701
rect 3798 1677 3804 1678
rect 112 1617 114 1677
rect 110 1616 116 1617
rect 132 1616 134 1677
rect 356 1616 358 1677
rect 596 1616 598 1677
rect 836 1616 838 1677
rect 1068 1616 1070 1677
rect 1308 1616 1310 1677
rect 1548 1616 1550 1677
rect 1936 1617 1938 1677
rect 1974 1673 1975 1677
rect 1979 1673 1980 1677
rect 1974 1672 1980 1673
rect 2470 1676 2476 1677
rect 2470 1672 2471 1676
rect 2475 1672 2476 1676
rect 2470 1671 2476 1672
rect 2606 1676 2612 1677
rect 2606 1672 2607 1676
rect 2611 1672 2612 1676
rect 2606 1671 2612 1672
rect 2742 1676 2748 1677
rect 2742 1672 2743 1676
rect 2747 1672 2748 1676
rect 2742 1671 2748 1672
rect 2878 1676 2884 1677
rect 2878 1672 2879 1676
rect 2883 1672 2884 1676
rect 2878 1671 2884 1672
rect 3022 1676 3028 1677
rect 3022 1672 3023 1676
rect 3027 1672 3028 1676
rect 3022 1671 3028 1672
rect 3174 1676 3180 1677
rect 3174 1672 3175 1676
rect 3179 1672 3180 1676
rect 3174 1671 3180 1672
rect 3326 1676 3332 1677
rect 3326 1672 3327 1676
rect 3331 1672 3332 1676
rect 3798 1673 3799 1677
rect 3803 1673 3804 1677
rect 3798 1672 3804 1673
rect 3326 1671 3332 1672
rect 2442 1661 2448 1662
rect 1974 1660 1980 1661
rect 1974 1656 1975 1660
rect 1979 1656 1980 1660
rect 2442 1657 2443 1661
rect 2447 1657 2448 1661
rect 2442 1656 2448 1657
rect 2578 1661 2584 1662
rect 2578 1657 2579 1661
rect 2583 1657 2584 1661
rect 2578 1656 2584 1657
rect 2714 1661 2720 1662
rect 2714 1657 2715 1661
rect 2719 1657 2720 1661
rect 2714 1656 2720 1657
rect 2850 1661 2856 1662
rect 2850 1657 2851 1661
rect 2855 1657 2856 1661
rect 2850 1656 2856 1657
rect 2994 1661 3000 1662
rect 2994 1657 2995 1661
rect 2999 1657 3000 1661
rect 2994 1656 3000 1657
rect 3146 1661 3152 1662
rect 3146 1657 3147 1661
rect 3151 1657 3152 1661
rect 3146 1656 3152 1657
rect 3298 1661 3304 1662
rect 3298 1657 3299 1661
rect 3303 1657 3304 1661
rect 3298 1656 3304 1657
rect 3798 1660 3804 1661
rect 3798 1656 3799 1660
rect 3803 1656 3804 1660
rect 1974 1655 1980 1656
rect 1934 1616 1940 1617
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 354 1615 360 1616
rect 354 1611 355 1615
rect 359 1611 360 1615
rect 354 1610 360 1611
rect 594 1615 600 1616
rect 594 1611 595 1615
rect 599 1611 600 1615
rect 594 1610 600 1611
rect 834 1615 840 1616
rect 834 1611 835 1615
rect 839 1611 840 1615
rect 834 1610 840 1611
rect 1066 1615 1072 1616
rect 1066 1611 1067 1615
rect 1071 1611 1072 1615
rect 1066 1610 1072 1611
rect 1306 1615 1312 1616
rect 1306 1611 1307 1615
rect 1311 1611 1312 1615
rect 1306 1610 1312 1611
rect 1546 1615 1552 1616
rect 1546 1611 1547 1615
rect 1551 1611 1552 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 1546 1610 1552 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 382 1600 388 1601
rect 382 1596 383 1600
rect 387 1596 388 1600
rect 382 1595 388 1596
rect 622 1600 628 1601
rect 622 1596 623 1600
rect 627 1596 628 1600
rect 622 1595 628 1596
rect 862 1600 868 1601
rect 862 1596 863 1600
rect 867 1596 868 1600
rect 862 1595 868 1596
rect 1094 1600 1100 1601
rect 1094 1596 1095 1600
rect 1099 1596 1100 1600
rect 1094 1595 1100 1596
rect 1334 1600 1340 1601
rect 1334 1596 1335 1600
rect 1339 1596 1340 1600
rect 1334 1595 1340 1596
rect 1574 1600 1580 1601
rect 1574 1596 1575 1600
rect 1579 1596 1580 1600
rect 1574 1595 1580 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 1976 1595 1978 1655
rect 2444 1595 2446 1656
rect 2580 1595 2582 1656
rect 2716 1595 2718 1656
rect 2852 1595 2854 1656
rect 2996 1595 2998 1656
rect 3148 1595 3150 1656
rect 3300 1595 3302 1656
rect 3798 1655 3804 1656
rect 3800 1595 3802 1655
rect 3840 1635 3842 1707
rect 4356 1635 4358 1708
rect 4572 1635 4574 1708
rect 4804 1635 4806 1708
rect 5044 1635 5046 1708
rect 5292 1635 5294 1708
rect 5516 1635 5518 1708
rect 5662 1707 5668 1708
rect 5664 1635 5666 1707
rect 3839 1634 3843 1635
rect 3839 1629 3843 1630
rect 3907 1634 3911 1635
rect 3907 1629 3911 1630
rect 4123 1634 4127 1635
rect 4123 1629 4127 1630
rect 4355 1634 4359 1635
rect 4355 1629 4359 1630
rect 4363 1634 4367 1635
rect 4363 1629 4367 1630
rect 4571 1634 4575 1635
rect 4571 1629 4575 1630
rect 4627 1634 4631 1635
rect 4627 1629 4631 1630
rect 4803 1634 4807 1635
rect 4803 1629 4807 1630
rect 4907 1634 4911 1635
rect 4907 1629 4911 1630
rect 5043 1634 5047 1635
rect 5043 1629 5047 1630
rect 5195 1634 5199 1635
rect 5195 1629 5199 1630
rect 5291 1634 5295 1635
rect 5291 1629 5295 1630
rect 5491 1634 5495 1635
rect 5491 1629 5495 1630
rect 5515 1634 5519 1635
rect 5515 1629 5519 1630
rect 5663 1634 5667 1635
rect 5663 1629 5667 1630
rect 110 1594 116 1595
rect 112 1567 114 1594
rect 160 1567 162 1595
rect 384 1567 386 1595
rect 624 1567 626 1595
rect 864 1567 866 1595
rect 1096 1567 1098 1595
rect 1336 1567 1338 1595
rect 1576 1567 1578 1595
rect 1934 1594 1940 1595
rect 1975 1594 1979 1595
rect 1936 1567 1938 1594
rect 1975 1589 1979 1590
rect 2355 1594 2359 1595
rect 2355 1589 2359 1590
rect 2443 1594 2447 1595
rect 2443 1589 2447 1590
rect 2563 1594 2567 1595
rect 2563 1589 2567 1590
rect 2579 1594 2583 1595
rect 2579 1589 2583 1590
rect 2715 1594 2719 1595
rect 2715 1589 2719 1590
rect 2779 1594 2783 1595
rect 2779 1589 2783 1590
rect 2851 1594 2855 1595
rect 2851 1589 2855 1590
rect 2995 1594 2999 1595
rect 2995 1589 2999 1590
rect 3003 1594 3007 1595
rect 3003 1589 3007 1590
rect 3147 1594 3151 1595
rect 3147 1589 3151 1590
rect 3227 1594 3231 1595
rect 3227 1589 3231 1590
rect 3299 1594 3303 1595
rect 3299 1589 3303 1590
rect 3459 1594 3463 1595
rect 3459 1589 3463 1590
rect 3799 1594 3803 1595
rect 3799 1589 3803 1590
rect 111 1566 115 1567
rect 111 1561 115 1562
rect 159 1566 163 1567
rect 159 1561 163 1562
rect 359 1566 363 1567
rect 359 1561 363 1562
rect 383 1566 387 1567
rect 383 1561 387 1562
rect 575 1566 579 1567
rect 575 1561 579 1562
rect 623 1566 627 1567
rect 623 1561 627 1562
rect 783 1566 787 1567
rect 783 1561 787 1562
rect 863 1566 867 1567
rect 863 1561 867 1562
rect 983 1566 987 1567
rect 983 1561 987 1562
rect 1095 1566 1099 1567
rect 1095 1561 1099 1562
rect 1183 1566 1187 1567
rect 1183 1561 1187 1562
rect 1335 1566 1339 1567
rect 1335 1561 1339 1562
rect 1375 1566 1379 1567
rect 1375 1561 1379 1562
rect 1575 1566 1579 1567
rect 1575 1561 1579 1562
rect 1935 1566 1939 1567
rect 1935 1561 1939 1562
rect 112 1538 114 1561
rect 110 1537 116 1538
rect 160 1537 162 1561
rect 360 1537 362 1561
rect 576 1537 578 1561
rect 784 1537 786 1561
rect 984 1537 986 1561
rect 1184 1537 1186 1561
rect 1376 1537 1378 1561
rect 1576 1537 1578 1561
rect 1936 1538 1938 1561
rect 1934 1537 1940 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 110 1532 116 1533
rect 158 1536 164 1537
rect 158 1532 159 1536
rect 163 1532 164 1536
rect 158 1531 164 1532
rect 358 1536 364 1537
rect 358 1532 359 1536
rect 363 1532 364 1536
rect 358 1531 364 1532
rect 574 1536 580 1537
rect 574 1532 575 1536
rect 579 1532 580 1536
rect 574 1531 580 1532
rect 782 1536 788 1537
rect 782 1532 783 1536
rect 787 1532 788 1536
rect 782 1531 788 1532
rect 982 1536 988 1537
rect 982 1532 983 1536
rect 987 1532 988 1536
rect 982 1531 988 1532
rect 1182 1536 1188 1537
rect 1182 1532 1183 1536
rect 1187 1532 1188 1536
rect 1182 1531 1188 1532
rect 1374 1536 1380 1537
rect 1374 1532 1375 1536
rect 1379 1532 1380 1536
rect 1374 1531 1380 1532
rect 1574 1536 1580 1537
rect 1574 1532 1575 1536
rect 1579 1532 1580 1536
rect 1934 1533 1935 1537
rect 1939 1533 1940 1537
rect 1934 1532 1940 1533
rect 1574 1531 1580 1532
rect 1976 1529 1978 1589
rect 1974 1528 1980 1529
rect 2356 1528 2358 1589
rect 2564 1528 2566 1589
rect 2780 1528 2782 1589
rect 3004 1528 3006 1589
rect 3228 1528 3230 1589
rect 3460 1528 3462 1589
rect 3800 1529 3802 1589
rect 3840 1569 3842 1629
rect 3838 1568 3844 1569
rect 3908 1568 3910 1629
rect 4124 1568 4126 1629
rect 4364 1568 4366 1629
rect 4628 1568 4630 1629
rect 4908 1568 4910 1629
rect 5196 1568 5198 1629
rect 5492 1568 5494 1629
rect 5664 1569 5666 1629
rect 5662 1568 5668 1569
rect 3838 1564 3839 1568
rect 3843 1564 3844 1568
rect 3838 1563 3844 1564
rect 3906 1567 3912 1568
rect 3906 1563 3907 1567
rect 3911 1563 3912 1567
rect 3906 1562 3912 1563
rect 4122 1567 4128 1568
rect 4122 1563 4123 1567
rect 4127 1563 4128 1567
rect 4122 1562 4128 1563
rect 4362 1567 4368 1568
rect 4362 1563 4363 1567
rect 4367 1563 4368 1567
rect 4362 1562 4368 1563
rect 4626 1567 4632 1568
rect 4626 1563 4627 1567
rect 4631 1563 4632 1567
rect 4626 1562 4632 1563
rect 4906 1567 4912 1568
rect 4906 1563 4907 1567
rect 4911 1563 4912 1567
rect 4906 1562 4912 1563
rect 5194 1567 5200 1568
rect 5194 1563 5195 1567
rect 5199 1563 5200 1567
rect 5194 1562 5200 1563
rect 5490 1567 5496 1568
rect 5490 1563 5491 1567
rect 5495 1563 5496 1567
rect 5662 1564 5663 1568
rect 5667 1564 5668 1568
rect 5662 1563 5668 1564
rect 5490 1562 5496 1563
rect 3934 1552 3940 1553
rect 3838 1551 3844 1552
rect 3838 1547 3839 1551
rect 3843 1547 3844 1551
rect 3934 1548 3935 1552
rect 3939 1548 3940 1552
rect 3934 1547 3940 1548
rect 4150 1552 4156 1553
rect 4150 1548 4151 1552
rect 4155 1548 4156 1552
rect 4150 1547 4156 1548
rect 4390 1552 4396 1553
rect 4390 1548 4391 1552
rect 4395 1548 4396 1552
rect 4390 1547 4396 1548
rect 4654 1552 4660 1553
rect 4654 1548 4655 1552
rect 4659 1548 4660 1552
rect 4654 1547 4660 1548
rect 4934 1552 4940 1553
rect 4934 1548 4935 1552
rect 4939 1548 4940 1552
rect 4934 1547 4940 1548
rect 5222 1552 5228 1553
rect 5222 1548 5223 1552
rect 5227 1548 5228 1552
rect 5222 1547 5228 1548
rect 5518 1552 5524 1553
rect 5518 1548 5519 1552
rect 5523 1548 5524 1552
rect 5518 1547 5524 1548
rect 5662 1551 5668 1552
rect 5662 1547 5663 1551
rect 5667 1547 5668 1551
rect 3838 1546 3844 1547
rect 3798 1528 3804 1529
rect 1974 1524 1975 1528
rect 1979 1524 1980 1528
rect 1974 1523 1980 1524
rect 2354 1527 2360 1528
rect 2354 1523 2355 1527
rect 2359 1523 2360 1527
rect 2354 1522 2360 1523
rect 2562 1527 2568 1528
rect 2562 1523 2563 1527
rect 2567 1523 2568 1527
rect 2562 1522 2568 1523
rect 2778 1527 2784 1528
rect 2778 1523 2779 1527
rect 2783 1523 2784 1527
rect 2778 1522 2784 1523
rect 3002 1527 3008 1528
rect 3002 1523 3003 1527
rect 3007 1523 3008 1527
rect 3002 1522 3008 1523
rect 3226 1527 3232 1528
rect 3226 1523 3227 1527
rect 3231 1523 3232 1527
rect 3226 1522 3232 1523
rect 3458 1527 3464 1528
rect 3458 1523 3459 1527
rect 3463 1523 3464 1527
rect 3798 1524 3799 1528
rect 3803 1524 3804 1528
rect 3798 1523 3804 1524
rect 3840 1523 3842 1546
rect 3936 1523 3938 1547
rect 4152 1523 4154 1547
rect 4392 1523 4394 1547
rect 4656 1523 4658 1547
rect 4936 1523 4938 1547
rect 5224 1523 5226 1547
rect 5520 1523 5522 1547
rect 5662 1546 5668 1547
rect 5664 1523 5666 1546
rect 3458 1522 3464 1523
rect 3839 1522 3843 1523
rect 130 1521 136 1522
rect 110 1520 116 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 130 1517 131 1521
rect 135 1517 136 1521
rect 130 1516 136 1517
rect 330 1521 336 1522
rect 330 1517 331 1521
rect 335 1517 336 1521
rect 330 1516 336 1517
rect 546 1521 552 1522
rect 546 1517 547 1521
rect 551 1517 552 1521
rect 546 1516 552 1517
rect 754 1521 760 1522
rect 754 1517 755 1521
rect 759 1517 760 1521
rect 754 1516 760 1517
rect 954 1521 960 1522
rect 954 1517 955 1521
rect 959 1517 960 1521
rect 954 1516 960 1517
rect 1154 1521 1160 1522
rect 1154 1517 1155 1521
rect 1159 1517 1160 1521
rect 1154 1516 1160 1517
rect 1346 1521 1352 1522
rect 1346 1517 1347 1521
rect 1351 1517 1352 1521
rect 1346 1516 1352 1517
rect 1546 1521 1552 1522
rect 1546 1517 1547 1521
rect 1551 1517 1552 1521
rect 1546 1516 1552 1517
rect 1934 1520 1940 1521
rect 1934 1516 1935 1520
rect 1939 1516 1940 1520
rect 3839 1517 3843 1518
rect 3887 1522 3891 1523
rect 3887 1517 3891 1518
rect 3935 1522 3939 1523
rect 3935 1517 3939 1518
rect 4023 1522 4027 1523
rect 4023 1517 4027 1518
rect 4151 1522 4155 1523
rect 4151 1517 4155 1518
rect 4159 1522 4163 1523
rect 4159 1517 4163 1518
rect 4295 1522 4299 1523
rect 4295 1517 4299 1518
rect 4391 1522 4395 1523
rect 4391 1517 4395 1518
rect 4479 1522 4483 1523
rect 4479 1517 4483 1518
rect 4655 1522 4659 1523
rect 4655 1517 4659 1518
rect 4695 1522 4699 1523
rect 4695 1517 4699 1518
rect 4935 1522 4939 1523
rect 4935 1517 4939 1518
rect 5191 1522 5195 1523
rect 5191 1517 5195 1518
rect 5223 1522 5227 1523
rect 5223 1517 5227 1518
rect 5447 1522 5451 1523
rect 5447 1517 5451 1518
rect 5519 1522 5523 1523
rect 5519 1517 5523 1518
rect 5663 1522 5667 1523
rect 5663 1517 5667 1518
rect 110 1515 116 1516
rect 112 1435 114 1515
rect 132 1435 134 1516
rect 332 1435 334 1516
rect 548 1435 550 1516
rect 756 1435 758 1516
rect 956 1435 958 1516
rect 1156 1435 1158 1516
rect 1348 1435 1350 1516
rect 1548 1435 1550 1516
rect 1934 1515 1940 1516
rect 1936 1435 1938 1515
rect 2382 1512 2388 1513
rect 1974 1511 1980 1512
rect 1974 1507 1975 1511
rect 1979 1507 1980 1511
rect 2382 1508 2383 1512
rect 2387 1508 2388 1512
rect 2382 1507 2388 1508
rect 2590 1512 2596 1513
rect 2590 1508 2591 1512
rect 2595 1508 2596 1512
rect 2590 1507 2596 1508
rect 2806 1512 2812 1513
rect 2806 1508 2807 1512
rect 2811 1508 2812 1512
rect 2806 1507 2812 1508
rect 3030 1512 3036 1513
rect 3030 1508 3031 1512
rect 3035 1508 3036 1512
rect 3030 1507 3036 1508
rect 3254 1512 3260 1513
rect 3254 1508 3255 1512
rect 3259 1508 3260 1512
rect 3254 1507 3260 1508
rect 3486 1512 3492 1513
rect 3486 1508 3487 1512
rect 3491 1508 3492 1512
rect 3486 1507 3492 1508
rect 3798 1511 3804 1512
rect 3798 1507 3799 1511
rect 3803 1507 3804 1511
rect 1974 1506 1980 1507
rect 1976 1483 1978 1506
rect 2384 1483 2386 1507
rect 2592 1483 2594 1507
rect 2808 1483 2810 1507
rect 3032 1483 3034 1507
rect 3256 1483 3258 1507
rect 3488 1483 3490 1507
rect 3798 1506 3804 1507
rect 3800 1483 3802 1506
rect 3840 1494 3842 1517
rect 3838 1493 3844 1494
rect 3888 1493 3890 1517
rect 4024 1493 4026 1517
rect 4160 1493 4162 1517
rect 4296 1493 4298 1517
rect 4480 1493 4482 1517
rect 4696 1493 4698 1517
rect 4936 1493 4938 1517
rect 5192 1493 5194 1517
rect 5448 1493 5450 1517
rect 5664 1494 5666 1517
rect 5662 1493 5668 1494
rect 3838 1489 3839 1493
rect 3843 1489 3844 1493
rect 3838 1488 3844 1489
rect 3886 1492 3892 1493
rect 3886 1488 3887 1492
rect 3891 1488 3892 1492
rect 3886 1487 3892 1488
rect 4022 1492 4028 1493
rect 4022 1488 4023 1492
rect 4027 1488 4028 1492
rect 4022 1487 4028 1488
rect 4158 1492 4164 1493
rect 4158 1488 4159 1492
rect 4163 1488 4164 1492
rect 4158 1487 4164 1488
rect 4294 1492 4300 1493
rect 4294 1488 4295 1492
rect 4299 1488 4300 1492
rect 4294 1487 4300 1488
rect 4478 1492 4484 1493
rect 4478 1488 4479 1492
rect 4483 1488 4484 1492
rect 4478 1487 4484 1488
rect 4694 1492 4700 1493
rect 4694 1488 4695 1492
rect 4699 1488 4700 1492
rect 4694 1487 4700 1488
rect 4934 1492 4940 1493
rect 4934 1488 4935 1492
rect 4939 1488 4940 1492
rect 4934 1487 4940 1488
rect 5190 1492 5196 1493
rect 5190 1488 5191 1492
rect 5195 1488 5196 1492
rect 5190 1487 5196 1488
rect 5446 1492 5452 1493
rect 5446 1488 5447 1492
rect 5451 1488 5452 1492
rect 5662 1489 5663 1493
rect 5667 1489 5668 1493
rect 5662 1488 5668 1489
rect 5446 1487 5452 1488
rect 1975 1482 1979 1483
rect 1975 1477 1979 1478
rect 2023 1482 2027 1483
rect 2023 1477 2027 1478
rect 2159 1482 2163 1483
rect 2159 1477 2163 1478
rect 2327 1482 2331 1483
rect 2327 1477 2331 1478
rect 2383 1482 2387 1483
rect 2383 1477 2387 1478
rect 2543 1482 2547 1483
rect 2543 1477 2547 1478
rect 2591 1482 2595 1483
rect 2591 1477 2595 1478
rect 2799 1482 2803 1483
rect 2799 1477 2803 1478
rect 2807 1482 2811 1483
rect 2807 1477 2811 1478
rect 3031 1482 3035 1483
rect 3031 1477 3035 1478
rect 3087 1482 3091 1483
rect 3087 1477 3091 1478
rect 3255 1482 3259 1483
rect 3255 1477 3259 1478
rect 3391 1482 3395 1483
rect 3391 1477 3395 1478
rect 3487 1482 3491 1483
rect 3487 1477 3491 1478
rect 3679 1482 3683 1483
rect 3679 1477 3683 1478
rect 3799 1482 3803 1483
rect 3799 1477 3803 1478
rect 3858 1477 3864 1478
rect 1976 1454 1978 1477
rect 1974 1453 1980 1454
rect 2024 1453 2026 1477
rect 2160 1453 2162 1477
rect 2328 1453 2330 1477
rect 2544 1453 2546 1477
rect 2800 1453 2802 1477
rect 3088 1453 3090 1477
rect 3392 1453 3394 1477
rect 3680 1453 3682 1477
rect 3800 1454 3802 1477
rect 3838 1476 3844 1477
rect 3838 1472 3839 1476
rect 3843 1472 3844 1476
rect 3858 1473 3859 1477
rect 3863 1473 3864 1477
rect 3858 1472 3864 1473
rect 3994 1477 4000 1478
rect 3994 1473 3995 1477
rect 3999 1473 4000 1477
rect 3994 1472 4000 1473
rect 4130 1477 4136 1478
rect 4130 1473 4131 1477
rect 4135 1473 4136 1477
rect 4130 1472 4136 1473
rect 4266 1477 4272 1478
rect 4266 1473 4267 1477
rect 4271 1473 4272 1477
rect 4266 1472 4272 1473
rect 4450 1477 4456 1478
rect 4450 1473 4451 1477
rect 4455 1473 4456 1477
rect 4450 1472 4456 1473
rect 4666 1477 4672 1478
rect 4666 1473 4667 1477
rect 4671 1473 4672 1477
rect 4666 1472 4672 1473
rect 4906 1477 4912 1478
rect 4906 1473 4907 1477
rect 4911 1473 4912 1477
rect 4906 1472 4912 1473
rect 5162 1477 5168 1478
rect 5162 1473 5163 1477
rect 5167 1473 5168 1477
rect 5162 1472 5168 1473
rect 5418 1477 5424 1478
rect 5418 1473 5419 1477
rect 5423 1473 5424 1477
rect 5418 1472 5424 1473
rect 5662 1476 5668 1477
rect 5662 1472 5663 1476
rect 5667 1472 5668 1476
rect 3838 1471 3844 1472
rect 3798 1453 3804 1454
rect 1974 1449 1975 1453
rect 1979 1449 1980 1453
rect 1974 1448 1980 1449
rect 2022 1452 2028 1453
rect 2022 1448 2023 1452
rect 2027 1448 2028 1452
rect 2022 1447 2028 1448
rect 2158 1452 2164 1453
rect 2158 1448 2159 1452
rect 2163 1448 2164 1452
rect 2158 1447 2164 1448
rect 2326 1452 2332 1453
rect 2326 1448 2327 1452
rect 2331 1448 2332 1452
rect 2326 1447 2332 1448
rect 2542 1452 2548 1453
rect 2542 1448 2543 1452
rect 2547 1448 2548 1452
rect 2542 1447 2548 1448
rect 2798 1452 2804 1453
rect 2798 1448 2799 1452
rect 2803 1448 2804 1452
rect 2798 1447 2804 1448
rect 3086 1452 3092 1453
rect 3086 1448 3087 1452
rect 3091 1448 3092 1452
rect 3086 1447 3092 1448
rect 3390 1452 3396 1453
rect 3390 1448 3391 1452
rect 3395 1448 3396 1452
rect 3390 1447 3396 1448
rect 3678 1452 3684 1453
rect 3678 1448 3679 1452
rect 3683 1448 3684 1452
rect 3798 1449 3799 1453
rect 3803 1449 3804 1453
rect 3798 1448 3804 1449
rect 3678 1447 3684 1448
rect 1994 1437 2000 1438
rect 1974 1436 1980 1437
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 131 1434 135 1435
rect 131 1429 135 1430
rect 235 1434 239 1435
rect 235 1429 239 1430
rect 331 1434 335 1435
rect 331 1429 335 1430
rect 507 1434 511 1435
rect 507 1429 511 1430
rect 547 1434 551 1435
rect 547 1429 551 1430
rect 755 1434 759 1435
rect 755 1429 759 1430
rect 779 1434 783 1435
rect 779 1429 783 1430
rect 955 1434 959 1435
rect 955 1429 959 1430
rect 1059 1434 1063 1435
rect 1059 1429 1063 1430
rect 1155 1434 1159 1435
rect 1155 1429 1159 1430
rect 1339 1434 1343 1435
rect 1339 1429 1343 1430
rect 1347 1434 1351 1435
rect 1347 1429 1351 1430
rect 1547 1434 1551 1435
rect 1547 1429 1551 1430
rect 1935 1434 1939 1435
rect 1974 1432 1975 1436
rect 1979 1432 1980 1436
rect 1994 1433 1995 1437
rect 1999 1433 2000 1437
rect 1994 1432 2000 1433
rect 2130 1437 2136 1438
rect 2130 1433 2131 1437
rect 2135 1433 2136 1437
rect 2130 1432 2136 1433
rect 2298 1437 2304 1438
rect 2298 1433 2299 1437
rect 2303 1433 2304 1437
rect 2298 1432 2304 1433
rect 2514 1437 2520 1438
rect 2514 1433 2515 1437
rect 2519 1433 2520 1437
rect 2514 1432 2520 1433
rect 2770 1437 2776 1438
rect 2770 1433 2771 1437
rect 2775 1433 2776 1437
rect 2770 1432 2776 1433
rect 3058 1437 3064 1438
rect 3058 1433 3059 1437
rect 3063 1433 3064 1437
rect 3058 1432 3064 1433
rect 3362 1437 3368 1438
rect 3362 1433 3363 1437
rect 3367 1433 3368 1437
rect 3362 1432 3368 1433
rect 3650 1437 3656 1438
rect 3650 1433 3651 1437
rect 3655 1433 3656 1437
rect 3650 1432 3656 1433
rect 3798 1436 3804 1437
rect 3798 1432 3799 1436
rect 3803 1432 3804 1436
rect 1974 1431 1980 1432
rect 1935 1429 1939 1430
rect 112 1369 114 1429
rect 110 1368 116 1369
rect 236 1368 238 1429
rect 508 1368 510 1429
rect 780 1368 782 1429
rect 1060 1368 1062 1429
rect 1340 1368 1342 1429
rect 1936 1369 1938 1429
rect 1976 1371 1978 1431
rect 1996 1371 1998 1432
rect 2132 1371 2134 1432
rect 2300 1371 2302 1432
rect 2516 1371 2518 1432
rect 2772 1371 2774 1432
rect 3060 1371 3062 1432
rect 3364 1371 3366 1432
rect 3652 1371 3654 1432
rect 3798 1431 3804 1432
rect 3800 1371 3802 1431
rect 3840 1399 3842 1471
rect 3860 1399 3862 1472
rect 3996 1399 3998 1472
rect 4132 1399 4134 1472
rect 4268 1399 4270 1472
rect 4452 1399 4454 1472
rect 4668 1399 4670 1472
rect 4908 1399 4910 1472
rect 5164 1399 5166 1472
rect 5420 1399 5422 1472
rect 5662 1471 5668 1472
rect 5664 1399 5666 1471
rect 3839 1398 3843 1399
rect 3839 1393 3843 1394
rect 3859 1398 3863 1399
rect 3859 1393 3863 1394
rect 3995 1398 3999 1399
rect 3995 1393 3999 1394
rect 4131 1398 4135 1399
rect 4131 1393 4135 1394
rect 4147 1398 4151 1399
rect 4147 1393 4151 1394
rect 4267 1398 4271 1399
rect 4267 1393 4271 1394
rect 4363 1398 4367 1399
rect 4363 1393 4367 1394
rect 4451 1398 4455 1399
rect 4451 1393 4455 1394
rect 4611 1398 4615 1399
rect 4611 1393 4615 1394
rect 4667 1398 4671 1399
rect 4667 1393 4671 1394
rect 4891 1398 4895 1399
rect 4891 1393 4895 1394
rect 4907 1398 4911 1399
rect 4907 1393 4911 1394
rect 5163 1398 5167 1399
rect 5163 1393 5167 1394
rect 5195 1398 5199 1399
rect 5195 1393 5199 1394
rect 5419 1398 5423 1399
rect 5419 1393 5423 1394
rect 5499 1398 5503 1399
rect 5499 1393 5503 1394
rect 5663 1398 5667 1399
rect 5663 1393 5667 1394
rect 1975 1370 1979 1371
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 234 1367 240 1368
rect 234 1363 235 1367
rect 239 1363 240 1367
rect 234 1362 240 1363
rect 506 1367 512 1368
rect 506 1363 507 1367
rect 511 1363 512 1367
rect 506 1362 512 1363
rect 778 1367 784 1368
rect 778 1363 779 1367
rect 783 1363 784 1367
rect 778 1362 784 1363
rect 1058 1367 1064 1368
rect 1058 1363 1059 1367
rect 1063 1363 1064 1367
rect 1058 1362 1064 1363
rect 1338 1367 1344 1368
rect 1338 1363 1339 1367
rect 1343 1363 1344 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1975 1365 1979 1366
rect 1995 1370 1999 1371
rect 1995 1365 1999 1366
rect 2131 1370 2135 1371
rect 2131 1365 2135 1366
rect 2299 1370 2303 1371
rect 2299 1365 2303 1366
rect 2491 1370 2495 1371
rect 2491 1365 2495 1366
rect 2515 1370 2519 1371
rect 2515 1365 2519 1366
rect 2771 1370 2775 1371
rect 2771 1365 2775 1366
rect 3019 1370 3023 1371
rect 3019 1365 3023 1366
rect 3059 1370 3063 1371
rect 3059 1365 3063 1366
rect 3363 1370 3367 1371
rect 3363 1365 3367 1366
rect 3555 1370 3559 1371
rect 3555 1365 3559 1366
rect 3651 1370 3655 1371
rect 3651 1365 3655 1366
rect 3799 1370 3803 1371
rect 3799 1365 3803 1366
rect 1934 1363 1940 1364
rect 1338 1362 1344 1363
rect 262 1352 268 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 262 1348 263 1352
rect 267 1348 268 1352
rect 262 1347 268 1348
rect 534 1352 540 1353
rect 534 1348 535 1352
rect 539 1348 540 1352
rect 534 1347 540 1348
rect 806 1352 812 1353
rect 806 1348 807 1352
rect 811 1348 812 1352
rect 806 1347 812 1348
rect 1086 1352 1092 1353
rect 1086 1348 1087 1352
rect 1091 1348 1092 1352
rect 1086 1347 1092 1348
rect 1366 1352 1372 1353
rect 1366 1348 1367 1352
rect 1371 1348 1372 1352
rect 1366 1347 1372 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 110 1346 116 1347
rect 112 1319 114 1346
rect 264 1319 266 1347
rect 536 1319 538 1347
rect 808 1319 810 1347
rect 1088 1319 1090 1347
rect 1368 1319 1370 1347
rect 1934 1346 1940 1347
rect 1936 1319 1938 1346
rect 111 1318 115 1319
rect 111 1313 115 1314
rect 159 1318 163 1319
rect 159 1313 163 1314
rect 263 1318 267 1319
rect 263 1313 267 1314
rect 383 1318 387 1319
rect 383 1313 387 1314
rect 535 1318 539 1319
rect 535 1313 539 1314
rect 599 1318 603 1319
rect 599 1313 603 1314
rect 799 1318 803 1319
rect 799 1313 803 1314
rect 807 1318 811 1319
rect 807 1313 811 1314
rect 991 1318 995 1319
rect 991 1313 995 1314
rect 1087 1318 1091 1319
rect 1087 1313 1091 1314
rect 1167 1318 1171 1319
rect 1167 1313 1171 1314
rect 1335 1318 1339 1319
rect 1335 1313 1339 1314
rect 1367 1318 1371 1319
rect 1367 1313 1371 1314
rect 1503 1318 1507 1319
rect 1503 1313 1507 1314
rect 1671 1318 1675 1319
rect 1671 1313 1675 1314
rect 1815 1318 1819 1319
rect 1815 1313 1819 1314
rect 1935 1318 1939 1319
rect 1935 1313 1939 1314
rect 112 1290 114 1313
rect 110 1289 116 1290
rect 160 1289 162 1313
rect 384 1289 386 1313
rect 600 1289 602 1313
rect 800 1289 802 1313
rect 992 1289 994 1313
rect 1168 1289 1170 1313
rect 1336 1289 1338 1313
rect 1504 1289 1506 1313
rect 1672 1289 1674 1313
rect 1816 1289 1818 1313
rect 1936 1290 1938 1313
rect 1976 1305 1978 1365
rect 1974 1304 1980 1305
rect 1996 1304 1998 1365
rect 2492 1304 2494 1365
rect 3020 1304 3022 1365
rect 3556 1304 3558 1365
rect 3800 1305 3802 1365
rect 3840 1333 3842 1393
rect 3838 1332 3844 1333
rect 3860 1332 3862 1393
rect 3996 1332 3998 1393
rect 4148 1332 4150 1393
rect 4364 1332 4366 1393
rect 4612 1332 4614 1393
rect 4892 1332 4894 1393
rect 5196 1332 5198 1393
rect 5500 1332 5502 1393
rect 5664 1333 5666 1393
rect 5662 1332 5668 1333
rect 3838 1328 3839 1332
rect 3843 1328 3844 1332
rect 3838 1327 3844 1328
rect 3858 1331 3864 1332
rect 3858 1327 3859 1331
rect 3863 1327 3864 1331
rect 3858 1326 3864 1327
rect 3994 1331 4000 1332
rect 3994 1327 3995 1331
rect 3999 1327 4000 1331
rect 3994 1326 4000 1327
rect 4146 1331 4152 1332
rect 4146 1327 4147 1331
rect 4151 1327 4152 1331
rect 4146 1326 4152 1327
rect 4362 1331 4368 1332
rect 4362 1327 4363 1331
rect 4367 1327 4368 1331
rect 4362 1326 4368 1327
rect 4610 1331 4616 1332
rect 4610 1327 4611 1331
rect 4615 1327 4616 1331
rect 4610 1326 4616 1327
rect 4890 1331 4896 1332
rect 4890 1327 4891 1331
rect 4895 1327 4896 1331
rect 4890 1326 4896 1327
rect 5194 1331 5200 1332
rect 5194 1327 5195 1331
rect 5199 1327 5200 1331
rect 5194 1326 5200 1327
rect 5498 1331 5504 1332
rect 5498 1327 5499 1331
rect 5503 1327 5504 1331
rect 5662 1328 5663 1332
rect 5667 1328 5668 1332
rect 5662 1327 5668 1328
rect 5498 1326 5504 1327
rect 3886 1316 3892 1317
rect 3838 1315 3844 1316
rect 3838 1311 3839 1315
rect 3843 1311 3844 1315
rect 3886 1312 3887 1316
rect 3891 1312 3892 1316
rect 3886 1311 3892 1312
rect 4022 1316 4028 1317
rect 4022 1312 4023 1316
rect 4027 1312 4028 1316
rect 4022 1311 4028 1312
rect 4174 1316 4180 1317
rect 4174 1312 4175 1316
rect 4179 1312 4180 1316
rect 4174 1311 4180 1312
rect 4390 1316 4396 1317
rect 4390 1312 4391 1316
rect 4395 1312 4396 1316
rect 4390 1311 4396 1312
rect 4638 1316 4644 1317
rect 4638 1312 4639 1316
rect 4643 1312 4644 1316
rect 4638 1311 4644 1312
rect 4918 1316 4924 1317
rect 4918 1312 4919 1316
rect 4923 1312 4924 1316
rect 4918 1311 4924 1312
rect 5222 1316 5228 1317
rect 5222 1312 5223 1316
rect 5227 1312 5228 1316
rect 5222 1311 5228 1312
rect 5526 1316 5532 1317
rect 5526 1312 5527 1316
rect 5531 1312 5532 1316
rect 5526 1311 5532 1312
rect 5662 1315 5668 1316
rect 5662 1311 5663 1315
rect 5667 1311 5668 1315
rect 3838 1310 3844 1311
rect 3798 1304 3804 1305
rect 1974 1300 1975 1304
rect 1979 1300 1980 1304
rect 1974 1299 1980 1300
rect 1994 1303 2000 1304
rect 1994 1299 1995 1303
rect 1999 1299 2000 1303
rect 1994 1298 2000 1299
rect 2490 1303 2496 1304
rect 2490 1299 2491 1303
rect 2495 1299 2496 1303
rect 2490 1298 2496 1299
rect 3018 1303 3024 1304
rect 3018 1299 3019 1303
rect 3023 1299 3024 1303
rect 3018 1298 3024 1299
rect 3554 1303 3560 1304
rect 3554 1299 3555 1303
rect 3559 1299 3560 1303
rect 3798 1300 3799 1304
rect 3803 1300 3804 1304
rect 3798 1299 3804 1300
rect 3554 1298 3560 1299
rect 1934 1289 1940 1290
rect 110 1285 111 1289
rect 115 1285 116 1289
rect 110 1284 116 1285
rect 158 1288 164 1289
rect 158 1284 159 1288
rect 163 1284 164 1288
rect 158 1283 164 1284
rect 382 1288 388 1289
rect 382 1284 383 1288
rect 387 1284 388 1288
rect 382 1283 388 1284
rect 598 1288 604 1289
rect 598 1284 599 1288
rect 603 1284 604 1288
rect 598 1283 604 1284
rect 798 1288 804 1289
rect 798 1284 799 1288
rect 803 1284 804 1288
rect 798 1283 804 1284
rect 990 1288 996 1289
rect 990 1284 991 1288
rect 995 1284 996 1288
rect 990 1283 996 1284
rect 1166 1288 1172 1289
rect 1166 1284 1167 1288
rect 1171 1284 1172 1288
rect 1166 1283 1172 1284
rect 1334 1288 1340 1289
rect 1334 1284 1335 1288
rect 1339 1284 1340 1288
rect 1334 1283 1340 1284
rect 1502 1288 1508 1289
rect 1502 1284 1503 1288
rect 1507 1284 1508 1288
rect 1502 1283 1508 1284
rect 1670 1288 1676 1289
rect 1670 1284 1671 1288
rect 1675 1284 1676 1288
rect 1670 1283 1676 1284
rect 1814 1288 1820 1289
rect 1814 1284 1815 1288
rect 1819 1284 1820 1288
rect 1934 1285 1935 1289
rect 1939 1285 1940 1289
rect 2022 1288 2028 1289
rect 1934 1284 1940 1285
rect 1974 1287 1980 1288
rect 1814 1283 1820 1284
rect 1974 1283 1975 1287
rect 1979 1283 1980 1287
rect 2022 1284 2023 1288
rect 2027 1284 2028 1288
rect 2022 1283 2028 1284
rect 2518 1288 2524 1289
rect 2518 1284 2519 1288
rect 2523 1284 2524 1288
rect 2518 1283 2524 1284
rect 3046 1288 3052 1289
rect 3046 1284 3047 1288
rect 3051 1284 3052 1288
rect 3046 1283 3052 1284
rect 3582 1288 3588 1289
rect 3582 1284 3583 1288
rect 3587 1284 3588 1288
rect 3582 1283 3588 1284
rect 3798 1287 3804 1288
rect 3840 1287 3842 1310
rect 3888 1287 3890 1311
rect 4024 1287 4026 1311
rect 4176 1287 4178 1311
rect 4392 1287 4394 1311
rect 4640 1287 4642 1311
rect 4920 1287 4922 1311
rect 5224 1287 5226 1311
rect 5528 1287 5530 1311
rect 5662 1310 5668 1311
rect 5664 1287 5666 1310
rect 3798 1283 3799 1287
rect 3803 1283 3804 1287
rect 1974 1282 1980 1283
rect 130 1273 136 1274
rect 110 1272 116 1273
rect 110 1268 111 1272
rect 115 1268 116 1272
rect 130 1269 131 1273
rect 135 1269 136 1273
rect 130 1268 136 1269
rect 354 1273 360 1274
rect 354 1269 355 1273
rect 359 1269 360 1273
rect 354 1268 360 1269
rect 570 1273 576 1274
rect 570 1269 571 1273
rect 575 1269 576 1273
rect 570 1268 576 1269
rect 770 1273 776 1274
rect 770 1269 771 1273
rect 775 1269 776 1273
rect 770 1268 776 1269
rect 962 1273 968 1274
rect 962 1269 963 1273
rect 967 1269 968 1273
rect 962 1268 968 1269
rect 1138 1273 1144 1274
rect 1138 1269 1139 1273
rect 1143 1269 1144 1273
rect 1138 1268 1144 1269
rect 1306 1273 1312 1274
rect 1306 1269 1307 1273
rect 1311 1269 1312 1273
rect 1306 1268 1312 1269
rect 1474 1273 1480 1274
rect 1474 1269 1475 1273
rect 1479 1269 1480 1273
rect 1474 1268 1480 1269
rect 1642 1273 1648 1274
rect 1642 1269 1643 1273
rect 1647 1269 1648 1273
rect 1642 1268 1648 1269
rect 1786 1273 1792 1274
rect 1786 1269 1787 1273
rect 1791 1269 1792 1273
rect 1786 1268 1792 1269
rect 1934 1272 1940 1273
rect 1934 1268 1935 1272
rect 1939 1268 1940 1272
rect 110 1267 116 1268
rect 112 1199 114 1267
rect 132 1199 134 1268
rect 356 1199 358 1268
rect 572 1199 574 1268
rect 772 1199 774 1268
rect 964 1199 966 1268
rect 1140 1199 1142 1268
rect 1308 1199 1310 1268
rect 1476 1199 1478 1268
rect 1644 1199 1646 1268
rect 1788 1199 1790 1268
rect 1934 1267 1940 1268
rect 1936 1199 1938 1267
rect 111 1198 115 1199
rect 111 1193 115 1194
rect 131 1198 135 1199
rect 131 1193 135 1194
rect 147 1198 151 1199
rect 147 1193 151 1194
rect 323 1198 327 1199
rect 323 1193 327 1194
rect 355 1198 359 1199
rect 355 1193 359 1194
rect 499 1198 503 1199
rect 499 1193 503 1194
rect 571 1198 575 1199
rect 571 1193 575 1194
rect 675 1198 679 1199
rect 675 1193 679 1194
rect 771 1198 775 1199
rect 771 1193 775 1194
rect 851 1198 855 1199
rect 851 1193 855 1194
rect 963 1198 967 1199
rect 963 1193 967 1194
rect 1019 1198 1023 1199
rect 1019 1193 1023 1194
rect 1139 1198 1143 1199
rect 1139 1193 1143 1194
rect 1179 1198 1183 1199
rect 1179 1193 1183 1194
rect 1307 1198 1311 1199
rect 1307 1193 1311 1194
rect 1331 1198 1335 1199
rect 1331 1193 1335 1194
rect 1475 1198 1479 1199
rect 1475 1193 1479 1194
rect 1483 1198 1487 1199
rect 1483 1193 1487 1194
rect 1643 1198 1647 1199
rect 1643 1193 1647 1194
rect 1787 1198 1791 1199
rect 1787 1193 1791 1194
rect 1935 1198 1939 1199
rect 1976 1195 1978 1282
rect 2024 1195 2026 1283
rect 2520 1195 2522 1283
rect 3048 1195 3050 1283
rect 3584 1195 3586 1283
rect 3798 1282 3804 1283
rect 3839 1286 3843 1287
rect 3800 1195 3802 1282
rect 3839 1281 3843 1282
rect 3887 1286 3891 1287
rect 3887 1281 3891 1282
rect 4023 1286 4027 1287
rect 4023 1281 4027 1282
rect 4167 1286 4171 1287
rect 4167 1281 4171 1282
rect 4175 1286 4179 1287
rect 4175 1281 4179 1282
rect 4335 1286 4339 1287
rect 4335 1281 4339 1282
rect 4391 1286 4395 1287
rect 4391 1281 4395 1282
rect 4511 1286 4515 1287
rect 4511 1281 4515 1282
rect 4639 1286 4643 1287
rect 4639 1281 4643 1282
rect 4703 1286 4707 1287
rect 4703 1281 4707 1282
rect 4903 1286 4907 1287
rect 4903 1281 4907 1282
rect 4919 1286 4923 1287
rect 4919 1281 4923 1282
rect 5119 1286 5123 1287
rect 5119 1281 5123 1282
rect 5223 1286 5227 1287
rect 5223 1281 5227 1282
rect 5343 1286 5347 1287
rect 5343 1281 5347 1282
rect 5527 1286 5531 1287
rect 5527 1281 5531 1282
rect 5543 1286 5547 1287
rect 5543 1281 5547 1282
rect 5663 1286 5667 1287
rect 5663 1281 5667 1282
rect 3840 1258 3842 1281
rect 3838 1257 3844 1258
rect 3888 1257 3890 1281
rect 4024 1257 4026 1281
rect 4168 1257 4170 1281
rect 4336 1257 4338 1281
rect 4512 1257 4514 1281
rect 4704 1257 4706 1281
rect 4904 1257 4906 1281
rect 5120 1257 5122 1281
rect 5344 1257 5346 1281
rect 5544 1257 5546 1281
rect 5664 1258 5666 1281
rect 5662 1257 5668 1258
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 3886 1256 3892 1257
rect 3886 1252 3887 1256
rect 3891 1252 3892 1256
rect 3886 1251 3892 1252
rect 4022 1256 4028 1257
rect 4022 1252 4023 1256
rect 4027 1252 4028 1256
rect 4022 1251 4028 1252
rect 4166 1256 4172 1257
rect 4166 1252 4167 1256
rect 4171 1252 4172 1256
rect 4166 1251 4172 1252
rect 4334 1256 4340 1257
rect 4334 1252 4335 1256
rect 4339 1252 4340 1256
rect 4334 1251 4340 1252
rect 4510 1256 4516 1257
rect 4510 1252 4511 1256
rect 4515 1252 4516 1256
rect 4510 1251 4516 1252
rect 4702 1256 4708 1257
rect 4702 1252 4703 1256
rect 4707 1252 4708 1256
rect 4702 1251 4708 1252
rect 4902 1256 4908 1257
rect 4902 1252 4903 1256
rect 4907 1252 4908 1256
rect 4902 1251 4908 1252
rect 5118 1256 5124 1257
rect 5118 1252 5119 1256
rect 5123 1252 5124 1256
rect 5118 1251 5124 1252
rect 5342 1256 5348 1257
rect 5342 1252 5343 1256
rect 5347 1252 5348 1256
rect 5342 1251 5348 1252
rect 5542 1256 5548 1257
rect 5542 1252 5543 1256
rect 5547 1252 5548 1256
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5542 1251 5548 1252
rect 3858 1241 3864 1242
rect 3838 1240 3844 1241
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 3858 1237 3859 1241
rect 3863 1237 3864 1241
rect 3858 1236 3864 1237
rect 3994 1241 4000 1242
rect 3994 1237 3995 1241
rect 3999 1237 4000 1241
rect 3994 1236 4000 1237
rect 4138 1241 4144 1242
rect 4138 1237 4139 1241
rect 4143 1237 4144 1241
rect 4138 1236 4144 1237
rect 4306 1241 4312 1242
rect 4306 1237 4307 1241
rect 4311 1237 4312 1241
rect 4306 1236 4312 1237
rect 4482 1241 4488 1242
rect 4482 1237 4483 1241
rect 4487 1237 4488 1241
rect 4482 1236 4488 1237
rect 4674 1241 4680 1242
rect 4674 1237 4675 1241
rect 4679 1237 4680 1241
rect 4674 1236 4680 1237
rect 4874 1241 4880 1242
rect 4874 1237 4875 1241
rect 4879 1237 4880 1241
rect 4874 1236 4880 1237
rect 5090 1241 5096 1242
rect 5090 1237 5091 1241
rect 5095 1237 5096 1241
rect 5090 1236 5096 1237
rect 5314 1241 5320 1242
rect 5314 1237 5315 1241
rect 5319 1237 5320 1241
rect 5314 1236 5320 1237
rect 5514 1241 5520 1242
rect 5514 1237 5515 1241
rect 5519 1237 5520 1241
rect 5514 1236 5520 1237
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 3838 1235 3844 1236
rect 1935 1193 1939 1194
rect 1975 1194 1979 1195
rect 112 1133 114 1193
rect 110 1132 116 1133
rect 148 1132 150 1193
rect 324 1132 326 1193
rect 500 1132 502 1193
rect 676 1132 678 1193
rect 852 1132 854 1193
rect 1020 1132 1022 1193
rect 1180 1132 1182 1193
rect 1332 1132 1334 1193
rect 1484 1132 1486 1193
rect 1644 1132 1646 1193
rect 1788 1132 1790 1193
rect 1936 1133 1938 1193
rect 1975 1189 1979 1190
rect 2023 1194 2027 1195
rect 2023 1189 2027 1190
rect 2519 1194 2523 1195
rect 2519 1189 2523 1190
rect 2743 1194 2747 1195
rect 2743 1189 2747 1190
rect 3047 1194 3051 1195
rect 3047 1189 3051 1190
rect 3359 1194 3363 1195
rect 3359 1189 3363 1190
rect 3583 1194 3587 1195
rect 3583 1189 3587 1190
rect 3679 1194 3683 1195
rect 3679 1189 3683 1190
rect 3799 1194 3803 1195
rect 3799 1189 3803 1190
rect 1976 1166 1978 1189
rect 1974 1165 1980 1166
rect 2744 1165 2746 1189
rect 3048 1165 3050 1189
rect 3360 1165 3362 1189
rect 3680 1165 3682 1189
rect 3800 1166 3802 1189
rect 3840 1171 3842 1235
rect 3860 1171 3862 1236
rect 3996 1171 3998 1236
rect 4140 1171 4142 1236
rect 4308 1171 4310 1236
rect 4484 1171 4486 1236
rect 4676 1171 4678 1236
rect 4876 1171 4878 1236
rect 5092 1171 5094 1236
rect 5316 1171 5318 1236
rect 5516 1171 5518 1236
rect 5662 1235 5668 1236
rect 5664 1171 5666 1235
rect 3839 1170 3843 1171
rect 3798 1165 3804 1166
rect 3839 1165 3843 1166
rect 3859 1170 3863 1171
rect 3859 1165 3863 1166
rect 3995 1170 3999 1171
rect 3995 1165 3999 1166
rect 4139 1170 4143 1171
rect 4139 1165 4143 1166
rect 4307 1170 4311 1171
rect 4307 1165 4311 1166
rect 4483 1170 4487 1171
rect 4483 1165 4487 1166
rect 4675 1170 4679 1171
rect 4675 1165 4679 1166
rect 4811 1170 4815 1171
rect 4811 1165 4815 1166
rect 4875 1170 4879 1171
rect 4875 1165 4879 1166
rect 4947 1170 4951 1171
rect 4947 1165 4951 1166
rect 5083 1170 5087 1171
rect 5083 1165 5087 1166
rect 5091 1170 5095 1171
rect 5091 1165 5095 1166
rect 5227 1170 5231 1171
rect 5227 1165 5231 1166
rect 5315 1170 5319 1171
rect 5315 1165 5319 1166
rect 5379 1170 5383 1171
rect 5379 1165 5383 1166
rect 5515 1170 5519 1171
rect 5515 1165 5519 1166
rect 5663 1170 5667 1171
rect 5663 1165 5667 1166
rect 1974 1161 1975 1165
rect 1979 1161 1980 1165
rect 1974 1160 1980 1161
rect 2742 1164 2748 1165
rect 2742 1160 2743 1164
rect 2747 1160 2748 1164
rect 2742 1159 2748 1160
rect 3046 1164 3052 1165
rect 3046 1160 3047 1164
rect 3051 1160 3052 1164
rect 3046 1159 3052 1160
rect 3358 1164 3364 1165
rect 3358 1160 3359 1164
rect 3363 1160 3364 1164
rect 3358 1159 3364 1160
rect 3678 1164 3684 1165
rect 3678 1160 3679 1164
rect 3683 1160 3684 1164
rect 3798 1161 3799 1165
rect 3803 1161 3804 1165
rect 3798 1160 3804 1161
rect 3678 1159 3684 1160
rect 2714 1149 2720 1150
rect 1974 1148 1980 1149
rect 1974 1144 1975 1148
rect 1979 1144 1980 1148
rect 2714 1145 2715 1149
rect 2719 1145 2720 1149
rect 2714 1144 2720 1145
rect 3018 1149 3024 1150
rect 3018 1145 3019 1149
rect 3023 1145 3024 1149
rect 3018 1144 3024 1145
rect 3330 1149 3336 1150
rect 3330 1145 3331 1149
rect 3335 1145 3336 1149
rect 3330 1144 3336 1145
rect 3650 1149 3656 1150
rect 3650 1145 3651 1149
rect 3655 1145 3656 1149
rect 3650 1144 3656 1145
rect 3798 1148 3804 1149
rect 3798 1144 3799 1148
rect 3803 1144 3804 1148
rect 1974 1143 1980 1144
rect 1934 1132 1940 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 146 1131 152 1132
rect 146 1127 147 1131
rect 151 1127 152 1131
rect 146 1126 152 1127
rect 322 1131 328 1132
rect 322 1127 323 1131
rect 327 1127 328 1131
rect 322 1126 328 1127
rect 498 1131 504 1132
rect 498 1127 499 1131
rect 503 1127 504 1131
rect 498 1126 504 1127
rect 674 1131 680 1132
rect 674 1127 675 1131
rect 679 1127 680 1131
rect 674 1126 680 1127
rect 850 1131 856 1132
rect 850 1127 851 1131
rect 855 1127 856 1131
rect 850 1126 856 1127
rect 1018 1131 1024 1132
rect 1018 1127 1019 1131
rect 1023 1127 1024 1131
rect 1018 1126 1024 1127
rect 1178 1131 1184 1132
rect 1178 1127 1179 1131
rect 1183 1127 1184 1131
rect 1178 1126 1184 1127
rect 1330 1131 1336 1132
rect 1330 1127 1331 1131
rect 1335 1127 1336 1131
rect 1330 1126 1336 1127
rect 1482 1131 1488 1132
rect 1482 1127 1483 1131
rect 1487 1127 1488 1131
rect 1482 1126 1488 1127
rect 1642 1131 1648 1132
rect 1642 1127 1643 1131
rect 1647 1127 1648 1131
rect 1642 1126 1648 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1786 1126 1792 1127
rect 174 1116 180 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 174 1112 175 1116
rect 179 1112 180 1116
rect 174 1111 180 1112
rect 350 1116 356 1117
rect 350 1112 351 1116
rect 355 1112 356 1116
rect 350 1111 356 1112
rect 526 1116 532 1117
rect 526 1112 527 1116
rect 531 1112 532 1116
rect 526 1111 532 1112
rect 702 1116 708 1117
rect 702 1112 703 1116
rect 707 1112 708 1116
rect 702 1111 708 1112
rect 878 1116 884 1117
rect 878 1112 879 1116
rect 883 1112 884 1116
rect 878 1111 884 1112
rect 1046 1116 1052 1117
rect 1046 1112 1047 1116
rect 1051 1112 1052 1116
rect 1046 1111 1052 1112
rect 1206 1116 1212 1117
rect 1206 1112 1207 1116
rect 1211 1112 1212 1116
rect 1206 1111 1212 1112
rect 1358 1116 1364 1117
rect 1358 1112 1359 1116
rect 1363 1112 1364 1116
rect 1358 1111 1364 1112
rect 1510 1116 1516 1117
rect 1510 1112 1511 1116
rect 1515 1112 1516 1116
rect 1510 1111 1516 1112
rect 1670 1116 1676 1117
rect 1670 1112 1671 1116
rect 1675 1112 1676 1116
rect 1670 1111 1676 1112
rect 1814 1116 1820 1117
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 110 1110 116 1111
rect 112 1067 114 1110
rect 176 1067 178 1111
rect 352 1067 354 1111
rect 528 1067 530 1111
rect 704 1067 706 1111
rect 880 1067 882 1111
rect 1048 1067 1050 1111
rect 1208 1067 1210 1111
rect 1360 1067 1362 1111
rect 1512 1067 1514 1111
rect 1672 1067 1674 1111
rect 1816 1067 1818 1111
rect 1934 1110 1940 1111
rect 1936 1067 1938 1110
rect 1976 1083 1978 1143
rect 2716 1083 2718 1144
rect 3020 1083 3022 1144
rect 3332 1083 3334 1144
rect 3652 1083 3654 1144
rect 3798 1143 3804 1144
rect 3800 1083 3802 1143
rect 3840 1105 3842 1165
rect 3838 1104 3844 1105
rect 4812 1104 4814 1165
rect 4948 1104 4950 1165
rect 5084 1104 5086 1165
rect 5228 1104 5230 1165
rect 5380 1104 5382 1165
rect 5516 1104 5518 1165
rect 5664 1105 5666 1165
rect 5662 1104 5668 1105
rect 3838 1100 3839 1104
rect 3843 1100 3844 1104
rect 3838 1099 3844 1100
rect 4810 1103 4816 1104
rect 4810 1099 4811 1103
rect 4815 1099 4816 1103
rect 4810 1098 4816 1099
rect 4946 1103 4952 1104
rect 4946 1099 4947 1103
rect 4951 1099 4952 1103
rect 4946 1098 4952 1099
rect 5082 1103 5088 1104
rect 5082 1099 5083 1103
rect 5087 1099 5088 1103
rect 5082 1098 5088 1099
rect 5226 1103 5232 1104
rect 5226 1099 5227 1103
rect 5231 1099 5232 1103
rect 5226 1098 5232 1099
rect 5378 1103 5384 1104
rect 5378 1099 5379 1103
rect 5383 1099 5384 1103
rect 5378 1098 5384 1099
rect 5514 1103 5520 1104
rect 5514 1099 5515 1103
rect 5519 1099 5520 1103
rect 5662 1100 5663 1104
rect 5667 1100 5668 1104
rect 5662 1099 5668 1100
rect 5514 1098 5520 1099
rect 4838 1088 4844 1089
rect 3838 1087 3844 1088
rect 3838 1083 3839 1087
rect 3843 1083 3844 1087
rect 4838 1084 4839 1088
rect 4843 1084 4844 1088
rect 4838 1083 4844 1084
rect 4974 1088 4980 1089
rect 4974 1084 4975 1088
rect 4979 1084 4980 1088
rect 4974 1083 4980 1084
rect 5110 1088 5116 1089
rect 5110 1084 5111 1088
rect 5115 1084 5116 1088
rect 5110 1083 5116 1084
rect 5254 1088 5260 1089
rect 5254 1084 5255 1088
rect 5259 1084 5260 1088
rect 5254 1083 5260 1084
rect 5406 1088 5412 1089
rect 5406 1084 5407 1088
rect 5411 1084 5412 1088
rect 5406 1083 5412 1084
rect 5542 1088 5548 1089
rect 5542 1084 5543 1088
rect 5547 1084 5548 1088
rect 5542 1083 5548 1084
rect 5662 1087 5668 1088
rect 5662 1083 5663 1087
rect 5667 1083 5668 1087
rect 1975 1082 1979 1083
rect 1975 1077 1979 1078
rect 2243 1082 2247 1083
rect 2243 1077 2247 1078
rect 2379 1082 2383 1083
rect 2379 1077 2383 1078
rect 2523 1082 2527 1083
rect 2523 1077 2527 1078
rect 2675 1082 2679 1083
rect 2675 1077 2679 1078
rect 2715 1082 2719 1083
rect 2715 1077 2719 1078
rect 2827 1082 2831 1083
rect 2827 1077 2831 1078
rect 2987 1082 2991 1083
rect 2987 1077 2991 1078
rect 3019 1082 3023 1083
rect 3019 1077 3023 1078
rect 3155 1082 3159 1083
rect 3155 1077 3159 1078
rect 3323 1082 3327 1083
rect 3323 1077 3327 1078
rect 3331 1082 3335 1083
rect 3331 1077 3335 1078
rect 3499 1082 3503 1083
rect 3499 1077 3503 1078
rect 3651 1082 3655 1083
rect 3651 1077 3655 1078
rect 3799 1082 3803 1083
rect 3838 1082 3844 1083
rect 3799 1077 3803 1078
rect 111 1066 115 1067
rect 111 1061 115 1062
rect 159 1066 163 1067
rect 159 1061 163 1062
rect 175 1066 179 1067
rect 175 1061 179 1062
rect 351 1066 355 1067
rect 351 1061 355 1062
rect 447 1066 451 1067
rect 447 1061 451 1062
rect 527 1066 531 1067
rect 527 1061 531 1062
rect 703 1066 707 1067
rect 703 1061 707 1062
rect 775 1066 779 1067
rect 775 1061 779 1062
rect 879 1066 883 1067
rect 879 1061 883 1062
rect 1047 1066 1051 1067
rect 1047 1061 1051 1062
rect 1111 1066 1115 1067
rect 1111 1061 1115 1062
rect 1207 1066 1211 1067
rect 1207 1061 1211 1062
rect 1359 1066 1363 1067
rect 1359 1061 1363 1062
rect 1455 1066 1459 1067
rect 1455 1061 1459 1062
rect 1511 1066 1515 1067
rect 1511 1061 1515 1062
rect 1671 1066 1675 1067
rect 1671 1061 1675 1062
rect 1807 1066 1811 1067
rect 1807 1061 1811 1062
rect 1815 1066 1819 1067
rect 1815 1061 1819 1062
rect 1935 1066 1939 1067
rect 1935 1061 1939 1062
rect 112 1038 114 1061
rect 110 1037 116 1038
rect 160 1037 162 1061
rect 448 1037 450 1061
rect 776 1037 778 1061
rect 1112 1037 1114 1061
rect 1456 1037 1458 1061
rect 1808 1037 1810 1061
rect 1936 1038 1938 1061
rect 1934 1037 1940 1038
rect 110 1033 111 1037
rect 115 1033 116 1037
rect 110 1032 116 1033
rect 158 1036 164 1037
rect 158 1032 159 1036
rect 163 1032 164 1036
rect 158 1031 164 1032
rect 446 1036 452 1037
rect 446 1032 447 1036
rect 451 1032 452 1036
rect 446 1031 452 1032
rect 774 1036 780 1037
rect 774 1032 775 1036
rect 779 1032 780 1036
rect 774 1031 780 1032
rect 1110 1036 1116 1037
rect 1110 1032 1111 1036
rect 1115 1032 1116 1036
rect 1110 1031 1116 1032
rect 1454 1036 1460 1037
rect 1454 1032 1455 1036
rect 1459 1032 1460 1036
rect 1454 1031 1460 1032
rect 1806 1036 1812 1037
rect 1806 1032 1807 1036
rect 1811 1032 1812 1036
rect 1934 1033 1935 1037
rect 1939 1033 1940 1037
rect 1934 1032 1940 1033
rect 1806 1031 1812 1032
rect 130 1021 136 1022
rect 110 1020 116 1021
rect 110 1016 111 1020
rect 115 1016 116 1020
rect 130 1017 131 1021
rect 135 1017 136 1021
rect 130 1016 136 1017
rect 418 1021 424 1022
rect 418 1017 419 1021
rect 423 1017 424 1021
rect 418 1016 424 1017
rect 746 1021 752 1022
rect 746 1017 747 1021
rect 751 1017 752 1021
rect 746 1016 752 1017
rect 1082 1021 1088 1022
rect 1082 1017 1083 1021
rect 1087 1017 1088 1021
rect 1082 1016 1088 1017
rect 1426 1021 1432 1022
rect 1426 1017 1427 1021
rect 1431 1017 1432 1021
rect 1426 1016 1432 1017
rect 1778 1021 1784 1022
rect 1778 1017 1779 1021
rect 1783 1017 1784 1021
rect 1778 1016 1784 1017
rect 1934 1020 1940 1021
rect 1934 1016 1935 1020
rect 1939 1016 1940 1020
rect 1976 1017 1978 1077
rect 110 1015 116 1016
rect 112 951 114 1015
rect 132 951 134 1016
rect 420 951 422 1016
rect 748 951 750 1016
rect 1084 951 1086 1016
rect 1428 951 1430 1016
rect 1780 951 1782 1016
rect 1934 1015 1940 1016
rect 1974 1016 1980 1017
rect 2244 1016 2246 1077
rect 2380 1016 2382 1077
rect 2524 1016 2526 1077
rect 2676 1016 2678 1077
rect 2828 1016 2830 1077
rect 2988 1016 2990 1077
rect 3156 1016 3158 1077
rect 3324 1016 3326 1077
rect 3500 1016 3502 1077
rect 3652 1016 3654 1077
rect 3800 1017 3802 1077
rect 3840 1055 3842 1082
rect 4840 1055 4842 1083
rect 4976 1055 4978 1083
rect 5112 1055 5114 1083
rect 5256 1055 5258 1083
rect 5408 1055 5410 1083
rect 5544 1055 5546 1083
rect 5662 1082 5668 1083
rect 5664 1055 5666 1082
rect 3839 1054 3843 1055
rect 3839 1049 3843 1050
rect 4807 1054 4811 1055
rect 4807 1049 4811 1050
rect 4839 1054 4843 1055
rect 4839 1049 4843 1050
rect 4943 1054 4947 1055
rect 4943 1049 4947 1050
rect 4975 1054 4979 1055
rect 4975 1049 4979 1050
rect 5079 1054 5083 1055
rect 5079 1049 5083 1050
rect 5111 1054 5115 1055
rect 5111 1049 5115 1050
rect 5215 1054 5219 1055
rect 5215 1049 5219 1050
rect 5255 1054 5259 1055
rect 5255 1049 5259 1050
rect 5351 1054 5355 1055
rect 5351 1049 5355 1050
rect 5407 1054 5411 1055
rect 5407 1049 5411 1050
rect 5487 1054 5491 1055
rect 5487 1049 5491 1050
rect 5543 1054 5547 1055
rect 5543 1049 5547 1050
rect 5663 1054 5667 1055
rect 5663 1049 5667 1050
rect 3840 1026 3842 1049
rect 3838 1025 3844 1026
rect 4808 1025 4810 1049
rect 4944 1025 4946 1049
rect 5080 1025 5082 1049
rect 5216 1025 5218 1049
rect 5352 1025 5354 1049
rect 5488 1025 5490 1049
rect 5664 1026 5666 1049
rect 5662 1025 5668 1026
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 4806 1024 4812 1025
rect 4806 1020 4807 1024
rect 4811 1020 4812 1024
rect 4806 1019 4812 1020
rect 4942 1024 4948 1025
rect 4942 1020 4943 1024
rect 4947 1020 4948 1024
rect 4942 1019 4948 1020
rect 5078 1024 5084 1025
rect 5078 1020 5079 1024
rect 5083 1020 5084 1024
rect 5078 1019 5084 1020
rect 5214 1024 5220 1025
rect 5214 1020 5215 1024
rect 5219 1020 5220 1024
rect 5214 1019 5220 1020
rect 5350 1024 5356 1025
rect 5350 1020 5351 1024
rect 5355 1020 5356 1024
rect 5350 1019 5356 1020
rect 5486 1024 5492 1025
rect 5486 1020 5487 1024
rect 5491 1020 5492 1024
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5486 1019 5492 1020
rect 3798 1016 3804 1017
rect 1936 951 1938 1015
rect 1974 1012 1975 1016
rect 1979 1012 1980 1016
rect 1974 1011 1980 1012
rect 2242 1015 2248 1016
rect 2242 1011 2243 1015
rect 2247 1011 2248 1015
rect 2242 1010 2248 1011
rect 2378 1015 2384 1016
rect 2378 1011 2379 1015
rect 2383 1011 2384 1015
rect 2378 1010 2384 1011
rect 2522 1015 2528 1016
rect 2522 1011 2523 1015
rect 2527 1011 2528 1015
rect 2522 1010 2528 1011
rect 2674 1015 2680 1016
rect 2674 1011 2675 1015
rect 2679 1011 2680 1015
rect 2674 1010 2680 1011
rect 2826 1015 2832 1016
rect 2826 1011 2827 1015
rect 2831 1011 2832 1015
rect 2826 1010 2832 1011
rect 2986 1015 2992 1016
rect 2986 1011 2987 1015
rect 2991 1011 2992 1015
rect 2986 1010 2992 1011
rect 3154 1015 3160 1016
rect 3154 1011 3155 1015
rect 3159 1011 3160 1015
rect 3154 1010 3160 1011
rect 3322 1015 3328 1016
rect 3322 1011 3323 1015
rect 3327 1011 3328 1015
rect 3322 1010 3328 1011
rect 3498 1015 3504 1016
rect 3498 1011 3499 1015
rect 3503 1011 3504 1015
rect 3498 1010 3504 1011
rect 3650 1015 3656 1016
rect 3650 1011 3651 1015
rect 3655 1011 3656 1015
rect 3798 1012 3799 1016
rect 3803 1012 3804 1016
rect 3798 1011 3804 1012
rect 3650 1010 3656 1011
rect 4778 1009 4784 1010
rect 3838 1008 3844 1009
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 4778 1005 4779 1009
rect 4783 1005 4784 1009
rect 4778 1004 4784 1005
rect 4914 1009 4920 1010
rect 4914 1005 4915 1009
rect 4919 1005 4920 1009
rect 4914 1004 4920 1005
rect 5050 1009 5056 1010
rect 5050 1005 5051 1009
rect 5055 1005 5056 1009
rect 5050 1004 5056 1005
rect 5186 1009 5192 1010
rect 5186 1005 5187 1009
rect 5191 1005 5192 1009
rect 5186 1004 5192 1005
rect 5322 1009 5328 1010
rect 5322 1005 5323 1009
rect 5327 1005 5328 1009
rect 5322 1004 5328 1005
rect 5458 1009 5464 1010
rect 5458 1005 5459 1009
rect 5463 1005 5464 1009
rect 5458 1004 5464 1005
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 3838 1003 3844 1004
rect 2270 1000 2276 1001
rect 1974 999 1980 1000
rect 1974 995 1975 999
rect 1979 995 1980 999
rect 2270 996 2271 1000
rect 2275 996 2276 1000
rect 2270 995 2276 996
rect 2406 1000 2412 1001
rect 2406 996 2407 1000
rect 2411 996 2412 1000
rect 2406 995 2412 996
rect 2550 1000 2556 1001
rect 2550 996 2551 1000
rect 2555 996 2556 1000
rect 2550 995 2556 996
rect 2702 1000 2708 1001
rect 2702 996 2703 1000
rect 2707 996 2708 1000
rect 2702 995 2708 996
rect 2854 1000 2860 1001
rect 2854 996 2855 1000
rect 2859 996 2860 1000
rect 2854 995 2860 996
rect 3014 1000 3020 1001
rect 3014 996 3015 1000
rect 3019 996 3020 1000
rect 3014 995 3020 996
rect 3182 1000 3188 1001
rect 3182 996 3183 1000
rect 3187 996 3188 1000
rect 3182 995 3188 996
rect 3350 1000 3356 1001
rect 3350 996 3351 1000
rect 3355 996 3356 1000
rect 3350 995 3356 996
rect 3526 1000 3532 1001
rect 3526 996 3527 1000
rect 3531 996 3532 1000
rect 3526 995 3532 996
rect 3678 1000 3684 1001
rect 3678 996 3679 1000
rect 3683 996 3684 1000
rect 3678 995 3684 996
rect 3798 999 3804 1000
rect 3798 995 3799 999
rect 3803 995 3804 999
rect 1974 994 1980 995
rect 1976 967 1978 994
rect 2272 967 2274 995
rect 2408 967 2410 995
rect 2552 967 2554 995
rect 2704 967 2706 995
rect 2856 967 2858 995
rect 3016 967 3018 995
rect 3184 967 3186 995
rect 3352 967 3354 995
rect 3528 967 3530 995
rect 3680 967 3682 995
rect 3798 994 3804 995
rect 3800 967 3802 994
rect 1975 966 1979 967
rect 1975 961 1979 962
rect 2271 966 2275 967
rect 2271 961 2275 962
rect 2279 966 2283 967
rect 2279 961 2283 962
rect 2407 966 2411 967
rect 2407 961 2411 962
rect 2495 966 2499 967
rect 2495 961 2499 962
rect 2551 966 2555 967
rect 2551 961 2555 962
rect 2703 966 2707 967
rect 2703 961 2707 962
rect 2711 966 2715 967
rect 2711 961 2715 962
rect 2855 966 2859 967
rect 2855 961 2859 962
rect 2911 966 2915 967
rect 2911 961 2915 962
rect 3015 966 3019 967
rect 3015 961 3019 962
rect 3103 966 3107 967
rect 3103 961 3107 962
rect 3183 966 3187 967
rect 3183 961 3187 962
rect 3295 966 3299 967
rect 3295 961 3299 962
rect 3351 966 3355 967
rect 3351 961 3355 962
rect 3479 966 3483 967
rect 3479 961 3483 962
rect 3527 966 3531 967
rect 3527 961 3531 962
rect 3671 966 3675 967
rect 3671 961 3675 962
rect 3679 966 3683 967
rect 3679 961 3683 962
rect 3799 966 3803 967
rect 3799 961 3803 962
rect 111 950 115 951
rect 111 945 115 946
rect 131 950 135 951
rect 131 945 135 946
rect 339 950 343 951
rect 339 945 343 946
rect 419 950 423 951
rect 419 945 423 946
rect 595 950 599 951
rect 595 945 599 946
rect 747 950 751 951
rect 747 945 751 946
rect 875 950 879 951
rect 875 945 879 946
rect 1083 950 1087 951
rect 1083 945 1087 946
rect 1179 950 1183 951
rect 1179 945 1183 946
rect 1427 950 1431 951
rect 1427 945 1431 946
rect 1491 950 1495 951
rect 1491 945 1495 946
rect 1779 950 1783 951
rect 1779 945 1783 946
rect 1787 950 1791 951
rect 1787 945 1791 946
rect 1935 950 1939 951
rect 1935 945 1939 946
rect 112 885 114 945
rect 110 884 116 885
rect 132 884 134 945
rect 340 884 342 945
rect 596 884 598 945
rect 876 884 878 945
rect 1180 884 1182 945
rect 1492 884 1494 945
rect 1788 884 1790 945
rect 1936 885 1938 945
rect 1976 938 1978 961
rect 1974 937 1980 938
rect 2280 937 2282 961
rect 2496 937 2498 961
rect 2712 937 2714 961
rect 2912 937 2914 961
rect 3104 937 3106 961
rect 3296 937 3298 961
rect 3480 937 3482 961
rect 3672 937 3674 961
rect 3800 938 3802 961
rect 3840 939 3842 1003
rect 4780 939 4782 1004
rect 4916 939 4918 1004
rect 5052 939 5054 1004
rect 5188 939 5190 1004
rect 5324 939 5326 1004
rect 5460 939 5462 1004
rect 5662 1003 5668 1004
rect 5664 939 5666 1003
rect 3839 938 3843 939
rect 3798 937 3804 938
rect 1974 933 1975 937
rect 1979 933 1980 937
rect 1974 932 1980 933
rect 2278 936 2284 937
rect 2278 932 2279 936
rect 2283 932 2284 936
rect 2278 931 2284 932
rect 2494 936 2500 937
rect 2494 932 2495 936
rect 2499 932 2500 936
rect 2494 931 2500 932
rect 2710 936 2716 937
rect 2710 932 2711 936
rect 2715 932 2716 936
rect 2710 931 2716 932
rect 2910 936 2916 937
rect 2910 932 2911 936
rect 2915 932 2916 936
rect 2910 931 2916 932
rect 3102 936 3108 937
rect 3102 932 3103 936
rect 3107 932 3108 936
rect 3102 931 3108 932
rect 3294 936 3300 937
rect 3294 932 3295 936
rect 3299 932 3300 936
rect 3294 931 3300 932
rect 3478 936 3484 937
rect 3478 932 3479 936
rect 3483 932 3484 936
rect 3478 931 3484 932
rect 3670 936 3676 937
rect 3670 932 3671 936
rect 3675 932 3676 936
rect 3798 933 3799 937
rect 3803 933 3804 937
rect 3839 933 3843 934
rect 4355 938 4359 939
rect 4355 933 4359 934
rect 4571 938 4575 939
rect 4571 933 4575 934
rect 4779 938 4783 939
rect 4779 933 4783 934
rect 4803 938 4807 939
rect 4803 933 4807 934
rect 4915 938 4919 939
rect 4915 933 4919 934
rect 5043 938 5047 939
rect 5043 933 5047 934
rect 5051 938 5055 939
rect 5051 933 5055 934
rect 5187 938 5191 939
rect 5187 933 5191 934
rect 5291 938 5295 939
rect 5291 933 5295 934
rect 5323 938 5327 939
rect 5323 933 5327 934
rect 5459 938 5463 939
rect 5459 933 5463 934
rect 5515 938 5519 939
rect 5515 933 5519 934
rect 5663 938 5667 939
rect 5663 933 5667 934
rect 3798 932 3804 933
rect 3670 931 3676 932
rect 2250 921 2256 922
rect 1974 920 1980 921
rect 1974 916 1975 920
rect 1979 916 1980 920
rect 2250 917 2251 921
rect 2255 917 2256 921
rect 2250 916 2256 917
rect 2466 921 2472 922
rect 2466 917 2467 921
rect 2471 917 2472 921
rect 2466 916 2472 917
rect 2682 921 2688 922
rect 2682 917 2683 921
rect 2687 917 2688 921
rect 2682 916 2688 917
rect 2882 921 2888 922
rect 2882 917 2883 921
rect 2887 917 2888 921
rect 2882 916 2888 917
rect 3074 921 3080 922
rect 3074 917 3075 921
rect 3079 917 3080 921
rect 3074 916 3080 917
rect 3266 921 3272 922
rect 3266 917 3267 921
rect 3271 917 3272 921
rect 3266 916 3272 917
rect 3450 921 3456 922
rect 3450 917 3451 921
rect 3455 917 3456 921
rect 3450 916 3456 917
rect 3642 921 3648 922
rect 3642 917 3643 921
rect 3647 917 3648 921
rect 3642 916 3648 917
rect 3798 920 3804 921
rect 3798 916 3799 920
rect 3803 916 3804 920
rect 1974 915 1980 916
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 130 883 136 884
rect 130 879 131 883
rect 135 879 136 883
rect 130 878 136 879
rect 338 883 344 884
rect 338 879 339 883
rect 343 879 344 883
rect 338 878 344 879
rect 594 883 600 884
rect 594 879 595 883
rect 599 879 600 883
rect 594 878 600 879
rect 874 883 880 884
rect 874 879 875 883
rect 879 879 880 883
rect 874 878 880 879
rect 1178 883 1184 884
rect 1178 879 1179 883
rect 1183 879 1184 883
rect 1178 878 1184 879
rect 1490 883 1496 884
rect 1490 879 1491 883
rect 1495 879 1496 883
rect 1490 878 1496 879
rect 1786 883 1792 884
rect 1786 879 1787 883
rect 1791 879 1792 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 1786 878 1792 879
rect 158 868 164 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 158 864 159 868
rect 163 864 164 868
rect 158 863 164 864
rect 366 868 372 869
rect 366 864 367 868
rect 371 864 372 868
rect 366 863 372 864
rect 622 868 628 869
rect 622 864 623 868
rect 627 864 628 868
rect 622 863 628 864
rect 902 868 908 869
rect 902 864 903 868
rect 907 864 908 868
rect 902 863 908 864
rect 1206 868 1212 869
rect 1206 864 1207 868
rect 1211 864 1212 868
rect 1206 863 1212 864
rect 1518 868 1524 869
rect 1518 864 1519 868
rect 1523 864 1524 868
rect 1518 863 1524 864
rect 1814 868 1820 869
rect 1814 864 1815 868
rect 1819 864 1820 868
rect 1814 863 1820 864
rect 1934 867 1940 868
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 110 862 116 863
rect 112 827 114 862
rect 160 827 162 863
rect 368 827 370 863
rect 624 827 626 863
rect 904 827 906 863
rect 1208 827 1210 863
rect 1520 827 1522 863
rect 1816 827 1818 863
rect 1934 862 1940 863
rect 1936 827 1938 862
rect 1976 851 1978 915
rect 2252 851 2254 916
rect 2468 851 2470 916
rect 2684 851 2686 916
rect 2884 851 2886 916
rect 3076 851 3078 916
rect 3268 851 3270 916
rect 3452 851 3454 916
rect 3644 851 3646 916
rect 3798 915 3804 916
rect 3800 851 3802 915
rect 3840 873 3842 933
rect 3838 872 3844 873
rect 4356 872 4358 933
rect 4572 872 4574 933
rect 4804 872 4806 933
rect 5044 872 5046 933
rect 5292 872 5294 933
rect 5516 872 5518 933
rect 5664 873 5666 933
rect 5662 872 5668 873
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 3838 867 3844 868
rect 4354 871 4360 872
rect 4354 867 4355 871
rect 4359 867 4360 871
rect 4354 866 4360 867
rect 4570 871 4576 872
rect 4570 867 4571 871
rect 4575 867 4576 871
rect 4570 866 4576 867
rect 4802 871 4808 872
rect 4802 867 4803 871
rect 4807 867 4808 871
rect 4802 866 4808 867
rect 5042 871 5048 872
rect 5042 867 5043 871
rect 5047 867 5048 871
rect 5042 866 5048 867
rect 5290 871 5296 872
rect 5290 867 5291 871
rect 5295 867 5296 871
rect 5290 866 5296 867
rect 5514 871 5520 872
rect 5514 867 5515 871
rect 5519 867 5520 871
rect 5662 868 5663 872
rect 5667 868 5668 872
rect 5662 867 5668 868
rect 5514 866 5520 867
rect 4382 856 4388 857
rect 3838 855 3844 856
rect 3838 851 3839 855
rect 3843 851 3844 855
rect 4382 852 4383 856
rect 4387 852 4388 856
rect 4382 851 4388 852
rect 4598 856 4604 857
rect 4598 852 4599 856
rect 4603 852 4604 856
rect 4598 851 4604 852
rect 4830 856 4836 857
rect 4830 852 4831 856
rect 4835 852 4836 856
rect 4830 851 4836 852
rect 5070 856 5076 857
rect 5070 852 5071 856
rect 5075 852 5076 856
rect 5070 851 5076 852
rect 5318 856 5324 857
rect 5318 852 5319 856
rect 5323 852 5324 856
rect 5318 851 5324 852
rect 5542 856 5548 857
rect 5542 852 5543 856
rect 5547 852 5548 856
rect 5542 851 5548 852
rect 5662 855 5668 856
rect 5662 851 5663 855
rect 5667 851 5668 855
rect 1975 850 1979 851
rect 1975 845 1979 846
rect 1995 850 1999 851
rect 1995 845 1999 846
rect 2131 850 2135 851
rect 2131 845 2135 846
rect 2251 850 2255 851
rect 2251 845 2255 846
rect 2283 850 2287 851
rect 2283 845 2287 846
rect 2443 850 2447 851
rect 2443 845 2447 846
rect 2467 850 2471 851
rect 2467 845 2471 846
rect 2603 850 2607 851
rect 2603 845 2607 846
rect 2683 850 2687 851
rect 2683 845 2687 846
rect 2763 850 2767 851
rect 2763 845 2767 846
rect 2883 850 2887 851
rect 2883 845 2887 846
rect 2923 850 2927 851
rect 2923 845 2927 846
rect 3075 850 3079 851
rect 3075 845 3079 846
rect 3083 850 3087 851
rect 3083 845 3087 846
rect 3243 850 3247 851
rect 3243 845 3247 846
rect 3267 850 3271 851
rect 3267 845 3271 846
rect 3403 850 3407 851
rect 3403 845 3407 846
rect 3451 850 3455 851
rect 3451 845 3455 846
rect 3643 850 3647 851
rect 3643 845 3647 846
rect 3799 850 3803 851
rect 3838 850 3844 851
rect 3799 845 3803 846
rect 111 826 115 827
rect 111 821 115 822
rect 159 826 163 827
rect 159 821 163 822
rect 367 826 371 827
rect 367 821 371 822
rect 383 826 387 827
rect 383 821 387 822
rect 623 826 627 827
rect 623 821 627 822
rect 631 826 635 827
rect 631 821 635 822
rect 887 826 891 827
rect 887 821 891 822
rect 903 826 907 827
rect 903 821 907 822
rect 1143 826 1147 827
rect 1143 821 1147 822
rect 1207 826 1211 827
rect 1207 821 1211 822
rect 1519 826 1523 827
rect 1519 821 1523 822
rect 1815 826 1819 827
rect 1815 821 1819 822
rect 1935 826 1939 827
rect 1935 821 1939 822
rect 112 798 114 821
rect 110 797 116 798
rect 160 797 162 821
rect 384 797 386 821
rect 632 797 634 821
rect 888 797 890 821
rect 1144 797 1146 821
rect 1936 798 1938 821
rect 1934 797 1940 798
rect 110 793 111 797
rect 115 793 116 797
rect 110 792 116 793
rect 158 796 164 797
rect 158 792 159 796
rect 163 792 164 796
rect 158 791 164 792
rect 382 796 388 797
rect 382 792 383 796
rect 387 792 388 796
rect 382 791 388 792
rect 630 796 636 797
rect 630 792 631 796
rect 635 792 636 796
rect 630 791 636 792
rect 886 796 892 797
rect 886 792 887 796
rect 891 792 892 796
rect 886 791 892 792
rect 1142 796 1148 797
rect 1142 792 1143 796
rect 1147 792 1148 796
rect 1934 793 1935 797
rect 1939 793 1940 797
rect 1934 792 1940 793
rect 1142 791 1148 792
rect 1976 785 1978 845
rect 1974 784 1980 785
rect 1996 784 1998 845
rect 2132 784 2134 845
rect 2284 784 2286 845
rect 2444 784 2446 845
rect 2604 784 2606 845
rect 2764 784 2766 845
rect 2924 784 2926 845
rect 3084 784 3086 845
rect 3244 784 3246 845
rect 3404 784 3406 845
rect 3800 785 3802 845
rect 3840 823 3842 850
rect 4384 823 4386 851
rect 4600 823 4602 851
rect 4832 823 4834 851
rect 5072 823 5074 851
rect 5320 823 5322 851
rect 5544 823 5546 851
rect 5662 850 5668 851
rect 5664 823 5666 850
rect 3839 822 3843 823
rect 3839 817 3843 818
rect 3959 822 3963 823
rect 3959 817 3963 818
rect 4207 822 4211 823
rect 4207 817 4211 818
rect 4383 822 4387 823
rect 4383 817 4387 818
rect 4495 822 4499 823
rect 4495 817 4499 818
rect 4599 822 4603 823
rect 4599 817 4603 818
rect 4815 822 4819 823
rect 4815 817 4819 818
rect 4831 822 4835 823
rect 4831 817 4835 818
rect 5071 822 5075 823
rect 5071 817 5075 818
rect 5151 822 5155 823
rect 5151 817 5155 818
rect 5319 822 5323 823
rect 5319 817 5323 818
rect 5487 822 5491 823
rect 5487 817 5491 818
rect 5543 822 5547 823
rect 5543 817 5547 818
rect 5663 822 5667 823
rect 5663 817 5667 818
rect 3840 794 3842 817
rect 3838 793 3844 794
rect 3960 793 3962 817
rect 4208 793 4210 817
rect 4496 793 4498 817
rect 4816 793 4818 817
rect 5152 793 5154 817
rect 5488 793 5490 817
rect 5664 794 5666 817
rect 5662 793 5668 794
rect 3838 789 3839 793
rect 3843 789 3844 793
rect 3838 788 3844 789
rect 3958 792 3964 793
rect 3958 788 3959 792
rect 3963 788 3964 792
rect 3958 787 3964 788
rect 4206 792 4212 793
rect 4206 788 4207 792
rect 4211 788 4212 792
rect 4206 787 4212 788
rect 4494 792 4500 793
rect 4494 788 4495 792
rect 4499 788 4500 792
rect 4494 787 4500 788
rect 4814 792 4820 793
rect 4814 788 4815 792
rect 4819 788 4820 792
rect 4814 787 4820 788
rect 5150 792 5156 793
rect 5150 788 5151 792
rect 5155 788 5156 792
rect 5150 787 5156 788
rect 5486 792 5492 793
rect 5486 788 5487 792
rect 5491 788 5492 792
rect 5662 789 5663 793
rect 5667 789 5668 793
rect 5662 788 5668 789
rect 5486 787 5492 788
rect 3798 784 3804 785
rect 130 781 136 782
rect 110 780 116 781
rect 110 776 111 780
rect 115 776 116 780
rect 130 777 131 781
rect 135 777 136 781
rect 130 776 136 777
rect 354 781 360 782
rect 354 777 355 781
rect 359 777 360 781
rect 354 776 360 777
rect 602 781 608 782
rect 602 777 603 781
rect 607 777 608 781
rect 602 776 608 777
rect 858 781 864 782
rect 858 777 859 781
rect 863 777 864 781
rect 858 776 864 777
rect 1114 781 1120 782
rect 1114 777 1115 781
rect 1119 777 1120 781
rect 1114 776 1120 777
rect 1934 780 1940 781
rect 1934 776 1935 780
rect 1939 776 1940 780
rect 1974 780 1975 784
rect 1979 780 1980 784
rect 1974 779 1980 780
rect 1994 783 2000 784
rect 1994 779 1995 783
rect 1999 779 2000 783
rect 1994 778 2000 779
rect 2130 783 2136 784
rect 2130 779 2131 783
rect 2135 779 2136 783
rect 2130 778 2136 779
rect 2282 783 2288 784
rect 2282 779 2283 783
rect 2287 779 2288 783
rect 2282 778 2288 779
rect 2442 783 2448 784
rect 2442 779 2443 783
rect 2447 779 2448 783
rect 2442 778 2448 779
rect 2602 783 2608 784
rect 2602 779 2603 783
rect 2607 779 2608 783
rect 2602 778 2608 779
rect 2762 783 2768 784
rect 2762 779 2763 783
rect 2767 779 2768 783
rect 2762 778 2768 779
rect 2922 783 2928 784
rect 2922 779 2923 783
rect 2927 779 2928 783
rect 2922 778 2928 779
rect 3082 783 3088 784
rect 3082 779 3083 783
rect 3087 779 3088 783
rect 3082 778 3088 779
rect 3242 783 3248 784
rect 3242 779 3243 783
rect 3247 779 3248 783
rect 3242 778 3248 779
rect 3402 783 3408 784
rect 3402 779 3403 783
rect 3407 779 3408 783
rect 3798 780 3799 784
rect 3803 780 3804 784
rect 3798 779 3804 780
rect 3402 778 3408 779
rect 3930 777 3936 778
rect 110 775 116 776
rect 112 715 114 775
rect 132 715 134 776
rect 356 715 358 776
rect 604 715 606 776
rect 860 715 862 776
rect 1116 715 1118 776
rect 1934 775 1940 776
rect 3838 776 3844 777
rect 1936 715 1938 775
rect 3838 772 3839 776
rect 3843 772 3844 776
rect 3930 773 3931 777
rect 3935 773 3936 777
rect 3930 772 3936 773
rect 4178 777 4184 778
rect 4178 773 4179 777
rect 4183 773 4184 777
rect 4178 772 4184 773
rect 4466 777 4472 778
rect 4466 773 4467 777
rect 4471 773 4472 777
rect 4466 772 4472 773
rect 4786 777 4792 778
rect 4786 773 4787 777
rect 4791 773 4792 777
rect 4786 772 4792 773
rect 5122 777 5128 778
rect 5122 773 5123 777
rect 5127 773 5128 777
rect 5122 772 5128 773
rect 5458 777 5464 778
rect 5458 773 5459 777
rect 5463 773 5464 777
rect 5458 772 5464 773
rect 5662 776 5668 777
rect 5662 772 5663 776
rect 5667 772 5668 776
rect 3838 771 3844 772
rect 2022 768 2028 769
rect 1974 767 1980 768
rect 1974 763 1975 767
rect 1979 763 1980 767
rect 2022 764 2023 768
rect 2027 764 2028 768
rect 2022 763 2028 764
rect 2158 768 2164 769
rect 2158 764 2159 768
rect 2163 764 2164 768
rect 2158 763 2164 764
rect 2310 768 2316 769
rect 2310 764 2311 768
rect 2315 764 2316 768
rect 2310 763 2316 764
rect 2470 768 2476 769
rect 2470 764 2471 768
rect 2475 764 2476 768
rect 2470 763 2476 764
rect 2630 768 2636 769
rect 2630 764 2631 768
rect 2635 764 2636 768
rect 2630 763 2636 764
rect 2790 768 2796 769
rect 2790 764 2791 768
rect 2795 764 2796 768
rect 2790 763 2796 764
rect 2950 768 2956 769
rect 2950 764 2951 768
rect 2955 764 2956 768
rect 2950 763 2956 764
rect 3110 768 3116 769
rect 3110 764 3111 768
rect 3115 764 3116 768
rect 3110 763 3116 764
rect 3270 768 3276 769
rect 3270 764 3271 768
rect 3275 764 3276 768
rect 3270 763 3276 764
rect 3430 768 3436 769
rect 3430 764 3431 768
rect 3435 764 3436 768
rect 3430 763 3436 764
rect 3798 767 3804 768
rect 3798 763 3799 767
rect 3803 763 3804 767
rect 1974 762 1980 763
rect 1976 739 1978 762
rect 2024 739 2026 763
rect 2160 739 2162 763
rect 2312 739 2314 763
rect 2472 739 2474 763
rect 2632 739 2634 763
rect 2792 739 2794 763
rect 2952 739 2954 763
rect 3112 739 3114 763
rect 3272 739 3274 763
rect 3432 739 3434 763
rect 3798 762 3804 763
rect 3800 739 3802 762
rect 1975 738 1979 739
rect 1975 733 1979 734
rect 2023 738 2027 739
rect 2023 733 2027 734
rect 2159 738 2163 739
rect 2159 733 2163 734
rect 2183 738 2187 739
rect 2183 733 2187 734
rect 2311 738 2315 739
rect 2311 733 2315 734
rect 2439 738 2443 739
rect 2439 733 2443 734
rect 2471 738 2475 739
rect 2471 733 2475 734
rect 2631 738 2635 739
rect 2631 733 2635 734
rect 2679 738 2683 739
rect 2679 733 2683 734
rect 2791 738 2795 739
rect 2791 733 2795 734
rect 2903 738 2907 739
rect 2903 733 2907 734
rect 2951 738 2955 739
rect 2951 733 2955 734
rect 3111 738 3115 739
rect 3111 733 3115 734
rect 3271 738 3275 739
rect 3271 733 3275 734
rect 3311 738 3315 739
rect 3311 733 3315 734
rect 3431 738 3435 739
rect 3431 733 3435 734
rect 3503 738 3507 739
rect 3503 733 3507 734
rect 3679 738 3683 739
rect 3679 733 3683 734
rect 3799 738 3803 739
rect 3799 733 3803 734
rect 111 714 115 715
rect 111 709 115 710
rect 131 714 135 715
rect 131 709 135 710
rect 355 714 359 715
rect 355 709 359 710
rect 603 714 607 715
rect 603 709 607 710
rect 699 714 703 715
rect 699 709 703 710
rect 835 714 839 715
rect 835 709 839 710
rect 859 714 863 715
rect 859 709 863 710
rect 971 714 975 715
rect 971 709 975 710
rect 1107 714 1111 715
rect 1107 709 1111 710
rect 1115 714 1119 715
rect 1115 709 1119 710
rect 1243 714 1247 715
rect 1243 709 1247 710
rect 1379 714 1383 715
rect 1379 709 1383 710
rect 1515 714 1519 715
rect 1515 709 1519 710
rect 1651 714 1655 715
rect 1651 709 1655 710
rect 1787 714 1791 715
rect 1787 709 1791 710
rect 1935 714 1939 715
rect 1976 710 1978 733
rect 1935 709 1939 710
rect 1974 709 1980 710
rect 2184 709 2186 733
rect 2440 709 2442 733
rect 2680 709 2682 733
rect 2904 709 2906 733
rect 3112 709 3114 733
rect 3312 709 3314 733
rect 3504 709 3506 733
rect 3680 709 3682 733
rect 3800 710 3802 733
rect 3798 709 3804 710
rect 112 649 114 709
rect 110 648 116 649
rect 700 648 702 709
rect 836 648 838 709
rect 972 648 974 709
rect 1108 648 1110 709
rect 1244 648 1246 709
rect 1380 648 1382 709
rect 1516 648 1518 709
rect 1652 648 1654 709
rect 1788 648 1790 709
rect 1936 649 1938 709
rect 1974 705 1975 709
rect 1979 705 1980 709
rect 1974 704 1980 705
rect 2182 708 2188 709
rect 2182 704 2183 708
rect 2187 704 2188 708
rect 2182 703 2188 704
rect 2438 708 2444 709
rect 2438 704 2439 708
rect 2443 704 2444 708
rect 2438 703 2444 704
rect 2678 708 2684 709
rect 2678 704 2679 708
rect 2683 704 2684 708
rect 2678 703 2684 704
rect 2902 708 2908 709
rect 2902 704 2903 708
rect 2907 704 2908 708
rect 2902 703 2908 704
rect 3110 708 3116 709
rect 3110 704 3111 708
rect 3115 704 3116 708
rect 3110 703 3116 704
rect 3310 708 3316 709
rect 3310 704 3311 708
rect 3315 704 3316 708
rect 3310 703 3316 704
rect 3502 708 3508 709
rect 3502 704 3503 708
rect 3507 704 3508 708
rect 3502 703 3508 704
rect 3678 708 3684 709
rect 3678 704 3679 708
rect 3683 704 3684 708
rect 3798 705 3799 709
rect 3803 705 3804 709
rect 3798 704 3804 705
rect 3678 703 3684 704
rect 3840 699 3842 771
rect 3932 699 3934 772
rect 4180 699 4182 772
rect 4468 699 4470 772
rect 4788 699 4790 772
rect 5124 699 5126 772
rect 5460 699 5462 772
rect 5662 771 5668 772
rect 5664 699 5666 771
rect 3839 698 3843 699
rect 2154 693 2160 694
rect 1974 692 1980 693
rect 1974 688 1975 692
rect 1979 688 1980 692
rect 2154 689 2155 693
rect 2159 689 2160 693
rect 2154 688 2160 689
rect 2410 693 2416 694
rect 2410 689 2411 693
rect 2415 689 2416 693
rect 2410 688 2416 689
rect 2650 693 2656 694
rect 2650 689 2651 693
rect 2655 689 2656 693
rect 2650 688 2656 689
rect 2874 693 2880 694
rect 2874 689 2875 693
rect 2879 689 2880 693
rect 2874 688 2880 689
rect 3082 693 3088 694
rect 3082 689 3083 693
rect 3087 689 3088 693
rect 3082 688 3088 689
rect 3282 693 3288 694
rect 3282 689 3283 693
rect 3287 689 3288 693
rect 3282 688 3288 689
rect 3474 693 3480 694
rect 3474 689 3475 693
rect 3479 689 3480 693
rect 3474 688 3480 689
rect 3650 693 3656 694
rect 3839 693 3843 694
rect 3859 698 3863 699
rect 3859 693 3863 694
rect 3931 698 3935 699
rect 3931 693 3935 694
rect 3995 698 3999 699
rect 3995 693 3999 694
rect 4147 698 4151 699
rect 4147 693 4151 694
rect 4179 698 4183 699
rect 4179 693 4183 694
rect 4355 698 4359 699
rect 4355 693 4359 694
rect 4467 698 4471 699
rect 4467 693 4471 694
rect 4595 698 4599 699
rect 4595 693 4599 694
rect 4787 698 4791 699
rect 4787 693 4791 694
rect 4867 698 4871 699
rect 4867 693 4871 694
rect 5123 698 5127 699
rect 5123 693 5127 694
rect 5163 698 5167 699
rect 5163 693 5167 694
rect 5459 698 5463 699
rect 5459 693 5463 694
rect 5663 698 5667 699
rect 5663 693 5667 694
rect 3650 689 3651 693
rect 3655 689 3656 693
rect 3650 688 3656 689
rect 3798 692 3804 693
rect 3798 688 3799 692
rect 3803 688 3804 692
rect 1974 687 1980 688
rect 1934 648 1940 649
rect 110 644 111 648
rect 115 644 116 648
rect 110 643 116 644
rect 698 647 704 648
rect 698 643 699 647
rect 703 643 704 647
rect 698 642 704 643
rect 834 647 840 648
rect 834 643 835 647
rect 839 643 840 647
rect 834 642 840 643
rect 970 647 976 648
rect 970 643 971 647
rect 975 643 976 647
rect 970 642 976 643
rect 1106 647 1112 648
rect 1106 643 1107 647
rect 1111 643 1112 647
rect 1106 642 1112 643
rect 1242 647 1248 648
rect 1242 643 1243 647
rect 1247 643 1248 647
rect 1242 642 1248 643
rect 1378 647 1384 648
rect 1378 643 1379 647
rect 1383 643 1384 647
rect 1378 642 1384 643
rect 1514 647 1520 648
rect 1514 643 1515 647
rect 1519 643 1520 647
rect 1514 642 1520 643
rect 1650 647 1656 648
rect 1650 643 1651 647
rect 1655 643 1656 647
rect 1650 642 1656 643
rect 1786 647 1792 648
rect 1786 643 1787 647
rect 1791 643 1792 647
rect 1934 644 1935 648
rect 1939 644 1940 648
rect 1934 643 1940 644
rect 1786 642 1792 643
rect 726 632 732 633
rect 110 631 116 632
rect 110 627 111 631
rect 115 627 116 631
rect 726 628 727 632
rect 731 628 732 632
rect 726 627 732 628
rect 862 632 868 633
rect 862 628 863 632
rect 867 628 868 632
rect 862 627 868 628
rect 998 632 1004 633
rect 998 628 999 632
rect 1003 628 1004 632
rect 998 627 1004 628
rect 1134 632 1140 633
rect 1134 628 1135 632
rect 1139 628 1140 632
rect 1134 627 1140 628
rect 1270 632 1276 633
rect 1270 628 1271 632
rect 1275 628 1276 632
rect 1270 627 1276 628
rect 1406 632 1412 633
rect 1406 628 1407 632
rect 1411 628 1412 632
rect 1406 627 1412 628
rect 1542 632 1548 633
rect 1542 628 1543 632
rect 1547 628 1548 632
rect 1542 627 1548 628
rect 1678 632 1684 633
rect 1678 628 1679 632
rect 1683 628 1684 632
rect 1678 627 1684 628
rect 1814 632 1820 633
rect 1814 628 1815 632
rect 1819 628 1820 632
rect 1814 627 1820 628
rect 1934 631 1940 632
rect 1934 627 1935 631
rect 1939 627 1940 631
rect 110 626 116 627
rect 112 603 114 626
rect 728 603 730 627
rect 864 603 866 627
rect 1000 603 1002 627
rect 1136 603 1138 627
rect 1272 603 1274 627
rect 1408 603 1410 627
rect 1544 603 1546 627
rect 1680 603 1682 627
rect 1816 603 1818 627
rect 1934 626 1940 627
rect 1936 603 1938 626
rect 111 602 115 603
rect 111 597 115 598
rect 159 602 163 603
rect 159 597 163 598
rect 375 602 379 603
rect 375 597 379 598
rect 599 602 603 603
rect 599 597 603 598
rect 727 602 731 603
rect 727 597 731 598
rect 807 602 811 603
rect 807 597 811 598
rect 863 602 867 603
rect 863 597 867 598
rect 999 602 1003 603
rect 999 597 1003 598
rect 1135 602 1139 603
rect 1135 597 1139 598
rect 1175 602 1179 603
rect 1175 597 1179 598
rect 1271 602 1275 603
rect 1271 597 1275 598
rect 1343 602 1347 603
rect 1343 597 1347 598
rect 1407 602 1411 603
rect 1407 597 1411 598
rect 1511 602 1515 603
rect 1511 597 1515 598
rect 1543 602 1547 603
rect 1543 597 1547 598
rect 1671 602 1675 603
rect 1671 597 1675 598
rect 1679 602 1683 603
rect 1679 597 1683 598
rect 1815 602 1819 603
rect 1815 597 1819 598
rect 1935 602 1939 603
rect 1935 597 1939 598
rect 112 574 114 597
rect 110 573 116 574
rect 160 573 162 597
rect 376 573 378 597
rect 600 573 602 597
rect 808 573 810 597
rect 1000 573 1002 597
rect 1176 573 1178 597
rect 1344 573 1346 597
rect 1512 573 1514 597
rect 1672 573 1674 597
rect 1816 573 1818 597
rect 1936 574 1938 597
rect 1934 573 1940 574
rect 110 569 111 573
rect 115 569 116 573
rect 110 568 116 569
rect 158 572 164 573
rect 158 568 159 572
rect 163 568 164 572
rect 158 567 164 568
rect 374 572 380 573
rect 374 568 375 572
rect 379 568 380 572
rect 374 567 380 568
rect 598 572 604 573
rect 598 568 599 572
rect 603 568 604 572
rect 598 567 604 568
rect 806 572 812 573
rect 806 568 807 572
rect 811 568 812 572
rect 806 567 812 568
rect 998 572 1004 573
rect 998 568 999 572
rect 1003 568 1004 572
rect 998 567 1004 568
rect 1174 572 1180 573
rect 1174 568 1175 572
rect 1179 568 1180 572
rect 1174 567 1180 568
rect 1342 572 1348 573
rect 1342 568 1343 572
rect 1347 568 1348 572
rect 1342 567 1348 568
rect 1510 572 1516 573
rect 1510 568 1511 572
rect 1515 568 1516 572
rect 1510 567 1516 568
rect 1670 572 1676 573
rect 1670 568 1671 572
rect 1675 568 1676 572
rect 1670 567 1676 568
rect 1814 572 1820 573
rect 1814 568 1815 572
rect 1819 568 1820 572
rect 1934 569 1935 573
rect 1939 569 1940 573
rect 1934 568 1940 569
rect 1814 567 1820 568
rect 130 557 136 558
rect 110 556 116 557
rect 110 552 111 556
rect 115 552 116 556
rect 130 553 131 557
rect 135 553 136 557
rect 130 552 136 553
rect 346 557 352 558
rect 346 553 347 557
rect 351 553 352 557
rect 346 552 352 553
rect 570 557 576 558
rect 570 553 571 557
rect 575 553 576 557
rect 570 552 576 553
rect 778 557 784 558
rect 778 553 779 557
rect 783 553 784 557
rect 778 552 784 553
rect 970 557 976 558
rect 970 553 971 557
rect 975 553 976 557
rect 970 552 976 553
rect 1146 557 1152 558
rect 1146 553 1147 557
rect 1151 553 1152 557
rect 1146 552 1152 553
rect 1314 557 1320 558
rect 1314 553 1315 557
rect 1319 553 1320 557
rect 1314 552 1320 553
rect 1482 557 1488 558
rect 1482 553 1483 557
rect 1487 553 1488 557
rect 1482 552 1488 553
rect 1642 557 1648 558
rect 1642 553 1643 557
rect 1647 553 1648 557
rect 1642 552 1648 553
rect 1786 557 1792 558
rect 1786 553 1787 557
rect 1791 553 1792 557
rect 1786 552 1792 553
rect 1934 556 1940 557
rect 1934 552 1935 556
rect 1939 552 1940 556
rect 110 551 116 552
rect 112 491 114 551
rect 132 491 134 552
rect 348 491 350 552
rect 572 491 574 552
rect 780 491 782 552
rect 972 491 974 552
rect 1148 491 1150 552
rect 1316 491 1318 552
rect 1484 491 1486 552
rect 1644 491 1646 552
rect 1788 491 1790 552
rect 1934 551 1940 552
rect 1936 491 1938 551
rect 111 490 115 491
rect 111 485 115 486
rect 131 490 135 491
rect 131 485 135 486
rect 347 490 351 491
rect 347 485 351 486
rect 355 490 359 491
rect 355 485 359 486
rect 571 490 575 491
rect 571 485 575 486
rect 603 490 607 491
rect 603 485 607 486
rect 779 490 783 491
rect 779 485 783 486
rect 843 490 847 491
rect 843 485 847 486
rect 971 490 975 491
rect 971 485 975 486
rect 1083 490 1087 491
rect 1083 485 1087 486
rect 1147 490 1151 491
rect 1147 485 1151 486
rect 1315 490 1319 491
rect 1315 485 1319 486
rect 1323 490 1327 491
rect 1323 485 1327 486
rect 1483 490 1487 491
rect 1483 485 1487 486
rect 1563 490 1567 491
rect 1563 485 1567 486
rect 1643 490 1647 491
rect 1643 485 1647 486
rect 1787 490 1791 491
rect 1787 485 1791 486
rect 1935 490 1939 491
rect 1935 485 1939 486
rect 112 425 114 485
rect 110 424 116 425
rect 132 424 134 485
rect 356 424 358 485
rect 604 424 606 485
rect 844 424 846 485
rect 1084 424 1086 485
rect 1324 424 1326 485
rect 1564 424 1566 485
rect 1788 424 1790 485
rect 1936 425 1938 485
rect 1976 451 1978 687
rect 2156 451 2158 688
rect 2412 451 2414 688
rect 2652 451 2654 688
rect 2876 451 2878 688
rect 3084 451 3086 688
rect 3284 451 3286 688
rect 3476 451 3478 688
rect 3652 451 3654 688
rect 3798 687 3804 688
rect 3800 451 3802 687
rect 3840 633 3842 693
rect 3838 632 3844 633
rect 3860 632 3862 693
rect 3996 632 3998 693
rect 4148 632 4150 693
rect 4356 632 4358 693
rect 4596 632 4598 693
rect 4868 632 4870 693
rect 5164 632 5166 693
rect 5460 632 5462 693
rect 5664 633 5666 693
rect 5662 632 5668 633
rect 3838 628 3839 632
rect 3843 628 3844 632
rect 3838 627 3844 628
rect 3858 631 3864 632
rect 3858 627 3859 631
rect 3863 627 3864 631
rect 3858 626 3864 627
rect 3994 631 4000 632
rect 3994 627 3995 631
rect 3999 627 4000 631
rect 3994 626 4000 627
rect 4146 631 4152 632
rect 4146 627 4147 631
rect 4151 627 4152 631
rect 4146 626 4152 627
rect 4354 631 4360 632
rect 4354 627 4355 631
rect 4359 627 4360 631
rect 4354 626 4360 627
rect 4594 631 4600 632
rect 4594 627 4595 631
rect 4599 627 4600 631
rect 4594 626 4600 627
rect 4866 631 4872 632
rect 4866 627 4867 631
rect 4871 627 4872 631
rect 4866 626 4872 627
rect 5162 631 5168 632
rect 5162 627 5163 631
rect 5167 627 5168 631
rect 5162 626 5168 627
rect 5458 631 5464 632
rect 5458 627 5459 631
rect 5463 627 5464 631
rect 5662 628 5663 632
rect 5667 628 5668 632
rect 5662 627 5668 628
rect 5458 626 5464 627
rect 3886 616 3892 617
rect 3838 615 3844 616
rect 3838 611 3839 615
rect 3843 611 3844 615
rect 3886 612 3887 616
rect 3891 612 3892 616
rect 3886 611 3892 612
rect 4022 616 4028 617
rect 4022 612 4023 616
rect 4027 612 4028 616
rect 4022 611 4028 612
rect 4174 616 4180 617
rect 4174 612 4175 616
rect 4179 612 4180 616
rect 4174 611 4180 612
rect 4382 616 4388 617
rect 4382 612 4383 616
rect 4387 612 4388 616
rect 4382 611 4388 612
rect 4622 616 4628 617
rect 4622 612 4623 616
rect 4627 612 4628 616
rect 4622 611 4628 612
rect 4894 616 4900 617
rect 4894 612 4895 616
rect 4899 612 4900 616
rect 4894 611 4900 612
rect 5190 616 5196 617
rect 5190 612 5191 616
rect 5195 612 5196 616
rect 5190 611 5196 612
rect 5486 616 5492 617
rect 5486 612 5487 616
rect 5491 612 5492 616
rect 5486 611 5492 612
rect 5662 615 5668 616
rect 5662 611 5663 615
rect 5667 611 5668 615
rect 3838 610 3844 611
rect 3840 587 3842 610
rect 3888 587 3890 611
rect 4024 587 4026 611
rect 4176 587 4178 611
rect 4384 587 4386 611
rect 4624 587 4626 611
rect 4896 587 4898 611
rect 5192 587 5194 611
rect 5488 587 5490 611
rect 5662 610 5668 611
rect 5664 587 5666 610
rect 3839 586 3843 587
rect 3839 581 3843 582
rect 3887 586 3891 587
rect 3887 581 3891 582
rect 4023 586 4027 587
rect 4023 581 4027 582
rect 4159 586 4163 587
rect 4159 581 4163 582
rect 4175 586 4179 587
rect 4175 581 4179 582
rect 4295 586 4299 587
rect 4295 581 4299 582
rect 4383 586 4387 587
rect 4383 581 4387 582
rect 4431 586 4435 587
rect 4431 581 4435 582
rect 4567 586 4571 587
rect 4567 581 4571 582
rect 4623 586 4627 587
rect 4623 581 4627 582
rect 4711 586 4715 587
rect 4711 581 4715 582
rect 4879 586 4883 587
rect 4879 581 4883 582
rect 4895 586 4899 587
rect 4895 581 4899 582
rect 5063 586 5067 587
rect 5063 581 5067 582
rect 5191 586 5195 587
rect 5191 581 5195 582
rect 5255 586 5259 587
rect 5255 581 5259 582
rect 5447 586 5451 587
rect 5447 581 5451 582
rect 5487 586 5491 587
rect 5487 581 5491 582
rect 5663 586 5667 587
rect 5663 581 5667 582
rect 3840 558 3842 581
rect 3838 557 3844 558
rect 3888 557 3890 581
rect 4024 557 4026 581
rect 4160 557 4162 581
rect 4296 557 4298 581
rect 4432 557 4434 581
rect 4568 557 4570 581
rect 4712 557 4714 581
rect 4880 557 4882 581
rect 5064 557 5066 581
rect 5256 557 5258 581
rect 5448 557 5450 581
rect 5664 558 5666 581
rect 5662 557 5668 558
rect 3838 553 3839 557
rect 3843 553 3844 557
rect 3838 552 3844 553
rect 3886 556 3892 557
rect 3886 552 3887 556
rect 3891 552 3892 556
rect 3886 551 3892 552
rect 4022 556 4028 557
rect 4022 552 4023 556
rect 4027 552 4028 556
rect 4022 551 4028 552
rect 4158 556 4164 557
rect 4158 552 4159 556
rect 4163 552 4164 556
rect 4158 551 4164 552
rect 4294 556 4300 557
rect 4294 552 4295 556
rect 4299 552 4300 556
rect 4294 551 4300 552
rect 4430 556 4436 557
rect 4430 552 4431 556
rect 4435 552 4436 556
rect 4430 551 4436 552
rect 4566 556 4572 557
rect 4566 552 4567 556
rect 4571 552 4572 556
rect 4566 551 4572 552
rect 4710 556 4716 557
rect 4710 552 4711 556
rect 4715 552 4716 556
rect 4710 551 4716 552
rect 4878 556 4884 557
rect 4878 552 4879 556
rect 4883 552 4884 556
rect 4878 551 4884 552
rect 5062 556 5068 557
rect 5062 552 5063 556
rect 5067 552 5068 556
rect 5062 551 5068 552
rect 5254 556 5260 557
rect 5254 552 5255 556
rect 5259 552 5260 556
rect 5254 551 5260 552
rect 5446 556 5452 557
rect 5446 552 5447 556
rect 5451 552 5452 556
rect 5662 553 5663 557
rect 5667 553 5668 557
rect 5662 552 5668 553
rect 5446 551 5452 552
rect 3858 541 3864 542
rect 3838 540 3844 541
rect 3838 536 3839 540
rect 3843 536 3844 540
rect 3858 537 3859 541
rect 3863 537 3864 541
rect 3858 536 3864 537
rect 3994 541 4000 542
rect 3994 537 3995 541
rect 3999 537 4000 541
rect 3994 536 4000 537
rect 4130 541 4136 542
rect 4130 537 4131 541
rect 4135 537 4136 541
rect 4130 536 4136 537
rect 4266 541 4272 542
rect 4266 537 4267 541
rect 4271 537 4272 541
rect 4266 536 4272 537
rect 4402 541 4408 542
rect 4402 537 4403 541
rect 4407 537 4408 541
rect 4402 536 4408 537
rect 4538 541 4544 542
rect 4538 537 4539 541
rect 4543 537 4544 541
rect 4538 536 4544 537
rect 4682 541 4688 542
rect 4682 537 4683 541
rect 4687 537 4688 541
rect 4682 536 4688 537
rect 4850 541 4856 542
rect 4850 537 4851 541
rect 4855 537 4856 541
rect 4850 536 4856 537
rect 5034 541 5040 542
rect 5034 537 5035 541
rect 5039 537 5040 541
rect 5034 536 5040 537
rect 5226 541 5232 542
rect 5226 537 5227 541
rect 5231 537 5232 541
rect 5226 536 5232 537
rect 5418 541 5424 542
rect 5418 537 5419 541
rect 5423 537 5424 541
rect 5418 536 5424 537
rect 5662 540 5668 541
rect 5662 536 5663 540
rect 5667 536 5668 540
rect 3838 535 3844 536
rect 3840 475 3842 535
rect 3860 475 3862 536
rect 3996 475 3998 536
rect 4132 475 4134 536
rect 4268 475 4270 536
rect 4404 475 4406 536
rect 4540 475 4542 536
rect 4684 475 4686 536
rect 4852 475 4854 536
rect 5036 475 5038 536
rect 5228 475 5230 536
rect 5420 475 5422 536
rect 5662 535 5668 536
rect 5664 475 5666 535
rect 3839 474 3843 475
rect 3839 469 3843 470
rect 3859 474 3863 475
rect 3859 469 3863 470
rect 3995 474 3999 475
rect 3995 469 3999 470
rect 4115 474 4119 475
rect 4115 469 4119 470
rect 4131 474 4135 475
rect 4131 469 4135 470
rect 4267 474 4271 475
rect 4267 469 4271 470
rect 4395 474 4399 475
rect 4395 469 4399 470
rect 4403 474 4407 475
rect 4403 469 4407 470
rect 4539 474 4543 475
rect 4539 469 4543 470
rect 4675 474 4679 475
rect 4675 469 4679 470
rect 4683 474 4687 475
rect 4683 469 4687 470
rect 4851 474 4855 475
rect 4851 469 4855 470
rect 4947 474 4951 475
rect 4947 469 4951 470
rect 5035 474 5039 475
rect 5035 469 5039 470
rect 5227 474 5231 475
rect 5227 469 5231 470
rect 5419 474 5423 475
rect 5419 469 5423 470
rect 5507 474 5511 475
rect 5507 469 5511 470
rect 5663 474 5667 475
rect 5663 469 5667 470
rect 1975 450 1979 451
rect 1975 445 1979 446
rect 1995 450 1999 451
rect 1995 445 1999 446
rect 2155 450 2159 451
rect 2155 445 2159 446
rect 2251 450 2255 451
rect 2251 445 2255 446
rect 2411 450 2415 451
rect 2411 445 2415 446
rect 2523 450 2527 451
rect 2523 445 2527 446
rect 2651 450 2655 451
rect 2651 445 2655 446
rect 2771 450 2775 451
rect 2771 445 2775 446
rect 2875 450 2879 451
rect 2875 445 2879 446
rect 3003 450 3007 451
rect 3003 445 3007 446
rect 3083 450 3087 451
rect 3083 445 3087 446
rect 3227 450 3231 451
rect 3227 445 3231 446
rect 3283 450 3287 451
rect 3283 445 3287 446
rect 3451 450 3455 451
rect 3451 445 3455 446
rect 3475 450 3479 451
rect 3475 445 3479 446
rect 3651 450 3655 451
rect 3651 445 3655 446
rect 3799 450 3803 451
rect 3799 445 3803 446
rect 1934 424 1940 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 130 423 136 424
rect 130 419 131 423
rect 135 419 136 423
rect 130 418 136 419
rect 354 423 360 424
rect 354 419 355 423
rect 359 419 360 423
rect 354 418 360 419
rect 602 423 608 424
rect 602 419 603 423
rect 607 419 608 423
rect 602 418 608 419
rect 842 423 848 424
rect 842 419 843 423
rect 847 419 848 423
rect 842 418 848 419
rect 1082 423 1088 424
rect 1082 419 1083 423
rect 1087 419 1088 423
rect 1082 418 1088 419
rect 1322 423 1328 424
rect 1322 419 1323 423
rect 1327 419 1328 423
rect 1322 418 1328 419
rect 1562 423 1568 424
rect 1562 419 1563 423
rect 1567 419 1568 423
rect 1562 418 1568 419
rect 1786 423 1792 424
rect 1786 419 1787 423
rect 1791 419 1792 423
rect 1934 420 1935 424
rect 1939 420 1940 424
rect 1934 419 1940 420
rect 1786 418 1792 419
rect 158 408 164 409
rect 110 407 116 408
rect 110 403 111 407
rect 115 403 116 407
rect 158 404 159 408
rect 163 404 164 408
rect 158 403 164 404
rect 382 408 388 409
rect 382 404 383 408
rect 387 404 388 408
rect 382 403 388 404
rect 630 408 636 409
rect 630 404 631 408
rect 635 404 636 408
rect 630 403 636 404
rect 870 408 876 409
rect 870 404 871 408
rect 875 404 876 408
rect 870 403 876 404
rect 1110 408 1116 409
rect 1110 404 1111 408
rect 1115 404 1116 408
rect 1110 403 1116 404
rect 1350 408 1356 409
rect 1350 404 1351 408
rect 1355 404 1356 408
rect 1350 403 1356 404
rect 1590 408 1596 409
rect 1590 404 1591 408
rect 1595 404 1596 408
rect 1590 403 1596 404
rect 1814 408 1820 409
rect 1814 404 1815 408
rect 1819 404 1820 408
rect 1814 403 1820 404
rect 1934 407 1940 408
rect 1934 403 1935 407
rect 1939 403 1940 407
rect 110 402 116 403
rect 112 363 114 402
rect 160 363 162 403
rect 384 363 386 403
rect 632 363 634 403
rect 872 363 874 403
rect 1112 363 1114 403
rect 1352 363 1354 403
rect 1592 363 1594 403
rect 1816 363 1818 403
rect 1934 402 1940 403
rect 1936 363 1938 402
rect 1976 385 1978 445
rect 1974 384 1980 385
rect 1996 384 1998 445
rect 2252 384 2254 445
rect 2524 384 2526 445
rect 2772 384 2774 445
rect 3004 384 3006 445
rect 3228 384 3230 445
rect 3452 384 3454 445
rect 3652 384 3654 445
rect 3800 385 3802 445
rect 3840 409 3842 469
rect 3838 408 3844 409
rect 3860 408 3862 469
rect 4116 408 4118 469
rect 4396 408 4398 469
rect 4676 408 4678 469
rect 4948 408 4950 469
rect 5228 408 5230 469
rect 5508 408 5510 469
rect 5664 409 5666 469
rect 5662 408 5668 409
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 3858 407 3864 408
rect 3858 403 3859 407
rect 3863 403 3864 407
rect 3858 402 3864 403
rect 4114 407 4120 408
rect 4114 403 4115 407
rect 4119 403 4120 407
rect 4114 402 4120 403
rect 4394 407 4400 408
rect 4394 403 4395 407
rect 4399 403 4400 407
rect 4394 402 4400 403
rect 4674 407 4680 408
rect 4674 403 4675 407
rect 4679 403 4680 407
rect 4674 402 4680 403
rect 4946 407 4952 408
rect 4946 403 4947 407
rect 4951 403 4952 407
rect 4946 402 4952 403
rect 5226 407 5232 408
rect 5226 403 5227 407
rect 5231 403 5232 407
rect 5226 402 5232 403
rect 5506 407 5512 408
rect 5506 403 5507 407
rect 5511 403 5512 407
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5506 402 5512 403
rect 3886 392 3892 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 3886 388 3887 392
rect 3891 388 3892 392
rect 3886 387 3892 388
rect 4142 392 4148 393
rect 4142 388 4143 392
rect 4147 388 4148 392
rect 4142 387 4148 388
rect 4422 392 4428 393
rect 4422 388 4423 392
rect 4427 388 4428 392
rect 4422 387 4428 388
rect 4702 392 4708 393
rect 4702 388 4703 392
rect 4707 388 4708 392
rect 4702 387 4708 388
rect 4974 392 4980 393
rect 4974 388 4975 392
rect 4979 388 4980 392
rect 4974 387 4980 388
rect 5254 392 5260 393
rect 5254 388 5255 392
rect 5259 388 5260 392
rect 5254 387 5260 388
rect 5534 392 5540 393
rect 5534 388 5535 392
rect 5539 388 5540 392
rect 5534 387 5540 388
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 3838 386 3844 387
rect 3798 384 3804 385
rect 1974 380 1975 384
rect 1979 380 1980 384
rect 1974 379 1980 380
rect 1994 383 2000 384
rect 1994 379 1995 383
rect 1999 379 2000 383
rect 1994 378 2000 379
rect 2250 383 2256 384
rect 2250 379 2251 383
rect 2255 379 2256 383
rect 2250 378 2256 379
rect 2522 383 2528 384
rect 2522 379 2523 383
rect 2527 379 2528 383
rect 2522 378 2528 379
rect 2770 383 2776 384
rect 2770 379 2771 383
rect 2775 379 2776 383
rect 2770 378 2776 379
rect 3002 383 3008 384
rect 3002 379 3003 383
rect 3007 379 3008 383
rect 3002 378 3008 379
rect 3226 383 3232 384
rect 3226 379 3227 383
rect 3231 379 3232 383
rect 3226 378 3232 379
rect 3450 383 3456 384
rect 3450 379 3451 383
rect 3455 379 3456 383
rect 3450 378 3456 379
rect 3650 383 3656 384
rect 3650 379 3651 383
rect 3655 379 3656 383
rect 3798 380 3799 384
rect 3803 380 3804 384
rect 3798 379 3804 380
rect 3650 378 3656 379
rect 2022 368 2028 369
rect 1974 367 1980 368
rect 1974 363 1975 367
rect 1979 363 1980 367
rect 2022 364 2023 368
rect 2027 364 2028 368
rect 2022 363 2028 364
rect 2278 368 2284 369
rect 2278 364 2279 368
rect 2283 364 2284 368
rect 2278 363 2284 364
rect 2550 368 2556 369
rect 2550 364 2551 368
rect 2555 364 2556 368
rect 2550 363 2556 364
rect 2798 368 2804 369
rect 2798 364 2799 368
rect 2803 364 2804 368
rect 2798 363 2804 364
rect 3030 368 3036 369
rect 3030 364 3031 368
rect 3035 364 3036 368
rect 3030 363 3036 364
rect 3254 368 3260 369
rect 3254 364 3255 368
rect 3259 364 3260 368
rect 3254 363 3260 364
rect 3478 368 3484 369
rect 3478 364 3479 368
rect 3483 364 3484 368
rect 3478 363 3484 364
rect 3678 368 3684 369
rect 3678 364 3679 368
rect 3683 364 3684 368
rect 3678 363 3684 364
rect 3798 367 3804 368
rect 3798 363 3799 367
rect 3803 363 3804 367
rect 111 362 115 363
rect 111 357 115 358
rect 159 362 163 363
rect 159 357 163 358
rect 303 362 307 363
rect 303 357 307 358
rect 383 362 387 363
rect 383 357 387 358
rect 479 362 483 363
rect 479 357 483 358
rect 631 362 635 363
rect 631 357 635 358
rect 655 362 659 363
rect 655 357 659 358
rect 831 362 835 363
rect 831 357 835 358
rect 871 362 875 363
rect 871 357 875 358
rect 1111 362 1115 363
rect 1111 357 1115 358
rect 1351 362 1355 363
rect 1351 357 1355 358
rect 1591 362 1595 363
rect 1591 357 1595 358
rect 1815 362 1819 363
rect 1815 357 1819 358
rect 1935 362 1939 363
rect 1974 362 1980 363
rect 1935 357 1939 358
rect 112 334 114 357
rect 110 333 116 334
rect 160 333 162 357
rect 304 333 306 357
rect 480 333 482 357
rect 656 333 658 357
rect 832 333 834 357
rect 1936 334 1938 357
rect 1976 335 1978 362
rect 2024 335 2026 363
rect 2280 335 2282 363
rect 2552 335 2554 363
rect 2800 335 2802 363
rect 3032 335 3034 363
rect 3256 335 3258 363
rect 3480 335 3482 363
rect 3680 335 3682 363
rect 3798 362 3804 363
rect 3800 335 3802 362
rect 3840 355 3842 386
rect 3888 355 3890 387
rect 4144 355 4146 387
rect 4424 355 4426 387
rect 4704 355 4706 387
rect 4976 355 4978 387
rect 5256 355 5258 387
rect 5536 355 5538 387
rect 5662 386 5668 387
rect 5664 355 5666 386
rect 3839 354 3843 355
rect 3839 349 3843 350
rect 3887 354 3891 355
rect 3887 349 3891 350
rect 4143 354 4147 355
rect 4143 349 4147 350
rect 4423 354 4427 355
rect 4423 349 4427 350
rect 4703 354 4707 355
rect 4703 349 4707 350
rect 4727 354 4731 355
rect 4727 349 4731 350
rect 4895 354 4899 355
rect 4895 349 4899 350
rect 4975 354 4979 355
rect 4975 349 4979 350
rect 5063 354 5067 355
rect 5063 349 5067 350
rect 5231 354 5235 355
rect 5231 349 5235 350
rect 5255 354 5259 355
rect 5255 349 5259 350
rect 5399 354 5403 355
rect 5399 349 5403 350
rect 5535 354 5539 355
rect 5535 349 5539 350
rect 5543 354 5547 355
rect 5543 349 5547 350
rect 5663 354 5667 355
rect 5663 349 5667 350
rect 1975 334 1979 335
rect 1934 333 1940 334
rect 110 329 111 333
rect 115 329 116 333
rect 110 328 116 329
rect 158 332 164 333
rect 158 328 159 332
rect 163 328 164 332
rect 158 327 164 328
rect 302 332 308 333
rect 302 328 303 332
rect 307 328 308 332
rect 302 327 308 328
rect 478 332 484 333
rect 478 328 479 332
rect 483 328 484 332
rect 478 327 484 328
rect 654 332 660 333
rect 654 328 655 332
rect 659 328 660 332
rect 654 327 660 328
rect 830 332 836 333
rect 830 328 831 332
rect 835 328 836 332
rect 1934 329 1935 333
rect 1939 329 1940 333
rect 1975 329 1979 330
rect 2023 334 2027 335
rect 2023 329 2027 330
rect 2159 334 2163 335
rect 2159 329 2163 330
rect 2279 334 2283 335
rect 2279 329 2283 330
rect 2295 334 2299 335
rect 2295 329 2299 330
rect 2431 334 2435 335
rect 2431 329 2435 330
rect 2551 334 2555 335
rect 2551 329 2555 330
rect 2567 334 2571 335
rect 2567 329 2571 330
rect 2703 334 2707 335
rect 2703 329 2707 330
rect 2799 334 2803 335
rect 2799 329 2803 330
rect 2839 334 2843 335
rect 2839 329 2843 330
rect 2975 334 2979 335
rect 2975 329 2979 330
rect 3031 334 3035 335
rect 3031 329 3035 330
rect 3111 334 3115 335
rect 3111 329 3115 330
rect 3247 334 3251 335
rect 3247 329 3251 330
rect 3255 334 3259 335
rect 3255 329 3259 330
rect 3383 334 3387 335
rect 3383 329 3387 330
rect 3479 334 3483 335
rect 3479 329 3483 330
rect 3519 334 3523 335
rect 3519 329 3523 330
rect 3655 334 3659 335
rect 3655 329 3659 330
rect 3679 334 3683 335
rect 3679 329 3683 330
rect 3799 334 3803 335
rect 3799 329 3803 330
rect 1934 328 1940 329
rect 830 327 836 328
rect 130 317 136 318
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 130 313 131 317
rect 135 313 136 317
rect 130 312 136 313
rect 274 317 280 318
rect 274 313 275 317
rect 279 313 280 317
rect 274 312 280 313
rect 450 317 456 318
rect 450 313 451 317
rect 455 313 456 317
rect 450 312 456 313
rect 626 317 632 318
rect 626 313 627 317
rect 631 313 632 317
rect 626 312 632 313
rect 802 317 808 318
rect 802 313 803 317
rect 807 313 808 317
rect 802 312 808 313
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 110 311 116 312
rect 112 211 114 311
rect 132 211 134 312
rect 276 211 278 312
rect 452 211 454 312
rect 628 211 630 312
rect 804 211 806 312
rect 1934 311 1940 312
rect 1936 211 1938 311
rect 1976 306 1978 329
rect 1974 305 1980 306
rect 2024 305 2026 329
rect 2160 305 2162 329
rect 2296 305 2298 329
rect 2432 305 2434 329
rect 2568 305 2570 329
rect 2704 305 2706 329
rect 2840 305 2842 329
rect 2976 305 2978 329
rect 3112 305 3114 329
rect 3248 305 3250 329
rect 3384 305 3386 329
rect 3520 305 3522 329
rect 3656 305 3658 329
rect 3800 306 3802 329
rect 3840 326 3842 349
rect 3838 325 3844 326
rect 4728 325 4730 349
rect 4896 325 4898 349
rect 5064 325 5066 349
rect 5232 325 5234 349
rect 5400 325 5402 349
rect 5544 325 5546 349
rect 5664 326 5666 349
rect 5662 325 5668 326
rect 3838 321 3839 325
rect 3843 321 3844 325
rect 3838 320 3844 321
rect 4726 324 4732 325
rect 4726 320 4727 324
rect 4731 320 4732 324
rect 4726 319 4732 320
rect 4894 324 4900 325
rect 4894 320 4895 324
rect 4899 320 4900 324
rect 4894 319 4900 320
rect 5062 324 5068 325
rect 5062 320 5063 324
rect 5067 320 5068 324
rect 5062 319 5068 320
rect 5230 324 5236 325
rect 5230 320 5231 324
rect 5235 320 5236 324
rect 5230 319 5236 320
rect 5398 324 5404 325
rect 5398 320 5399 324
rect 5403 320 5404 324
rect 5398 319 5404 320
rect 5542 324 5548 325
rect 5542 320 5543 324
rect 5547 320 5548 324
rect 5662 321 5663 325
rect 5667 321 5668 325
rect 5662 320 5668 321
rect 5542 319 5548 320
rect 4698 309 4704 310
rect 3838 308 3844 309
rect 3798 305 3804 306
rect 1974 301 1975 305
rect 1979 301 1980 305
rect 1974 300 1980 301
rect 2022 304 2028 305
rect 2022 300 2023 304
rect 2027 300 2028 304
rect 2022 299 2028 300
rect 2158 304 2164 305
rect 2158 300 2159 304
rect 2163 300 2164 304
rect 2158 299 2164 300
rect 2294 304 2300 305
rect 2294 300 2295 304
rect 2299 300 2300 304
rect 2294 299 2300 300
rect 2430 304 2436 305
rect 2430 300 2431 304
rect 2435 300 2436 304
rect 2430 299 2436 300
rect 2566 304 2572 305
rect 2566 300 2567 304
rect 2571 300 2572 304
rect 2566 299 2572 300
rect 2702 304 2708 305
rect 2702 300 2703 304
rect 2707 300 2708 304
rect 2702 299 2708 300
rect 2838 304 2844 305
rect 2838 300 2839 304
rect 2843 300 2844 304
rect 2838 299 2844 300
rect 2974 304 2980 305
rect 2974 300 2975 304
rect 2979 300 2980 304
rect 2974 299 2980 300
rect 3110 304 3116 305
rect 3110 300 3111 304
rect 3115 300 3116 304
rect 3110 299 3116 300
rect 3246 304 3252 305
rect 3246 300 3247 304
rect 3251 300 3252 304
rect 3246 299 3252 300
rect 3382 304 3388 305
rect 3382 300 3383 304
rect 3387 300 3388 304
rect 3382 299 3388 300
rect 3518 304 3524 305
rect 3518 300 3519 304
rect 3523 300 3524 304
rect 3518 299 3524 300
rect 3654 304 3660 305
rect 3654 300 3655 304
rect 3659 300 3660 304
rect 3798 301 3799 305
rect 3803 301 3804 305
rect 3838 304 3839 308
rect 3843 304 3844 308
rect 4698 305 4699 309
rect 4703 305 4704 309
rect 4698 304 4704 305
rect 4866 309 4872 310
rect 4866 305 4867 309
rect 4871 305 4872 309
rect 4866 304 4872 305
rect 5034 309 5040 310
rect 5034 305 5035 309
rect 5039 305 5040 309
rect 5034 304 5040 305
rect 5202 309 5208 310
rect 5202 305 5203 309
rect 5207 305 5208 309
rect 5202 304 5208 305
rect 5370 309 5376 310
rect 5370 305 5371 309
rect 5375 305 5376 309
rect 5370 304 5376 305
rect 5514 309 5520 310
rect 5514 305 5515 309
rect 5519 305 5520 309
rect 5514 304 5520 305
rect 5662 308 5668 309
rect 5662 304 5663 308
rect 5667 304 5668 308
rect 3838 303 3844 304
rect 3798 300 3804 301
rect 3654 299 3660 300
rect 1994 289 2000 290
rect 1974 288 1980 289
rect 1974 284 1975 288
rect 1979 284 1980 288
rect 1994 285 1995 289
rect 1999 285 2000 289
rect 1994 284 2000 285
rect 2130 289 2136 290
rect 2130 285 2131 289
rect 2135 285 2136 289
rect 2130 284 2136 285
rect 2266 289 2272 290
rect 2266 285 2267 289
rect 2271 285 2272 289
rect 2266 284 2272 285
rect 2402 289 2408 290
rect 2402 285 2403 289
rect 2407 285 2408 289
rect 2402 284 2408 285
rect 2538 289 2544 290
rect 2538 285 2539 289
rect 2543 285 2544 289
rect 2538 284 2544 285
rect 2674 289 2680 290
rect 2674 285 2675 289
rect 2679 285 2680 289
rect 2674 284 2680 285
rect 2810 289 2816 290
rect 2810 285 2811 289
rect 2815 285 2816 289
rect 2810 284 2816 285
rect 2946 289 2952 290
rect 2946 285 2947 289
rect 2951 285 2952 289
rect 2946 284 2952 285
rect 3082 289 3088 290
rect 3082 285 3083 289
rect 3087 285 3088 289
rect 3082 284 3088 285
rect 3218 289 3224 290
rect 3218 285 3219 289
rect 3223 285 3224 289
rect 3218 284 3224 285
rect 3354 289 3360 290
rect 3354 285 3355 289
rect 3359 285 3360 289
rect 3354 284 3360 285
rect 3490 289 3496 290
rect 3490 285 3491 289
rect 3495 285 3496 289
rect 3490 284 3496 285
rect 3626 289 3632 290
rect 3626 285 3627 289
rect 3631 285 3632 289
rect 3626 284 3632 285
rect 3798 288 3804 289
rect 3798 284 3799 288
rect 3803 284 3804 288
rect 1974 283 1980 284
rect 111 210 115 211
rect 111 205 115 206
rect 131 210 135 211
rect 131 205 135 206
rect 267 210 271 211
rect 267 205 271 206
rect 275 210 279 211
rect 275 205 279 206
rect 403 210 407 211
rect 403 205 407 206
rect 451 210 455 211
rect 451 205 455 206
rect 539 210 543 211
rect 539 205 543 206
rect 627 210 631 211
rect 627 205 631 206
rect 675 210 679 211
rect 675 205 679 206
rect 803 210 807 211
rect 803 205 807 206
rect 811 210 815 211
rect 811 205 815 206
rect 947 210 951 211
rect 947 205 951 206
rect 1083 210 1087 211
rect 1083 205 1087 206
rect 1935 210 1939 211
rect 1935 205 1939 206
rect 112 145 114 205
rect 110 144 116 145
rect 132 144 134 205
rect 268 144 270 205
rect 404 144 406 205
rect 540 144 542 205
rect 676 144 678 205
rect 812 144 814 205
rect 948 144 950 205
rect 1084 144 1086 205
rect 1936 145 1938 205
rect 1976 191 1978 283
rect 1996 191 1998 284
rect 2132 191 2134 284
rect 2268 191 2270 284
rect 2404 191 2406 284
rect 2540 191 2542 284
rect 2676 191 2678 284
rect 2812 191 2814 284
rect 2948 191 2950 284
rect 3084 191 3086 284
rect 3220 191 3222 284
rect 3356 191 3358 284
rect 3492 191 3494 284
rect 3628 191 3630 284
rect 3798 283 3804 284
rect 3800 191 3802 283
rect 3840 203 3842 303
rect 4700 203 4702 304
rect 4868 203 4870 304
rect 5036 203 5038 304
rect 5204 203 5206 304
rect 5372 203 5374 304
rect 5516 203 5518 304
rect 5662 303 5668 304
rect 5664 203 5666 303
rect 3839 202 3843 203
rect 3839 197 3843 198
rect 4291 202 4295 203
rect 4291 197 4295 198
rect 4427 202 4431 203
rect 4427 197 4431 198
rect 4563 202 4567 203
rect 4563 197 4567 198
rect 4699 202 4703 203
rect 4699 197 4703 198
rect 4835 202 4839 203
rect 4835 197 4839 198
rect 4867 202 4871 203
rect 4867 197 4871 198
rect 4971 202 4975 203
rect 4971 197 4975 198
rect 5035 202 5039 203
rect 5035 197 5039 198
rect 5107 202 5111 203
rect 5107 197 5111 198
rect 5203 202 5207 203
rect 5203 197 5207 198
rect 5243 202 5247 203
rect 5243 197 5247 198
rect 5371 202 5375 203
rect 5371 197 5375 198
rect 5379 202 5383 203
rect 5379 197 5383 198
rect 5515 202 5519 203
rect 5515 197 5519 198
rect 5663 202 5667 203
rect 5663 197 5667 198
rect 1975 190 1979 191
rect 1975 185 1979 186
rect 1995 190 1999 191
rect 1995 185 1999 186
rect 2131 190 2135 191
rect 2131 185 2135 186
rect 2267 190 2271 191
rect 2267 185 2271 186
rect 2403 190 2407 191
rect 2403 185 2407 186
rect 2539 190 2543 191
rect 2539 185 2543 186
rect 2675 190 2679 191
rect 2675 185 2679 186
rect 2811 190 2815 191
rect 2811 185 2815 186
rect 2947 190 2951 191
rect 2947 185 2951 186
rect 3083 190 3087 191
rect 3083 185 3087 186
rect 3219 190 3223 191
rect 3219 185 3223 186
rect 3355 190 3359 191
rect 3355 185 3359 186
rect 3491 190 3495 191
rect 3491 185 3495 186
rect 3627 190 3631 191
rect 3627 185 3631 186
rect 3799 190 3803 191
rect 3799 185 3803 186
rect 1934 144 1940 145
rect 110 140 111 144
rect 115 140 116 144
rect 110 139 116 140
rect 130 143 136 144
rect 130 139 131 143
rect 135 139 136 143
rect 130 138 136 139
rect 266 143 272 144
rect 266 139 267 143
rect 271 139 272 143
rect 266 138 272 139
rect 402 143 408 144
rect 402 139 403 143
rect 407 139 408 143
rect 402 138 408 139
rect 538 143 544 144
rect 538 139 539 143
rect 543 139 544 143
rect 538 138 544 139
rect 674 143 680 144
rect 674 139 675 143
rect 679 139 680 143
rect 674 138 680 139
rect 810 143 816 144
rect 810 139 811 143
rect 815 139 816 143
rect 810 138 816 139
rect 946 143 952 144
rect 946 139 947 143
rect 951 139 952 143
rect 946 138 952 139
rect 1082 143 1088 144
rect 1082 139 1083 143
rect 1087 139 1088 143
rect 1934 140 1935 144
rect 1939 140 1940 144
rect 1934 139 1940 140
rect 1082 138 1088 139
rect 158 128 164 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 158 124 159 128
rect 163 124 164 128
rect 158 123 164 124
rect 294 128 300 129
rect 294 124 295 128
rect 299 124 300 128
rect 294 123 300 124
rect 430 128 436 129
rect 430 124 431 128
rect 435 124 436 128
rect 430 123 436 124
rect 566 128 572 129
rect 566 124 567 128
rect 571 124 572 128
rect 566 123 572 124
rect 702 128 708 129
rect 702 124 703 128
rect 707 124 708 128
rect 702 123 708 124
rect 838 128 844 129
rect 838 124 839 128
rect 843 124 844 128
rect 838 123 844 124
rect 974 128 980 129
rect 974 124 975 128
rect 979 124 980 128
rect 974 123 980 124
rect 1110 128 1116 129
rect 1110 124 1111 128
rect 1115 124 1116 128
rect 1110 123 1116 124
rect 1934 127 1940 128
rect 1934 123 1935 127
rect 1939 123 1940 127
rect 1976 125 1978 185
rect 110 122 116 123
rect 112 99 114 122
rect 160 99 162 123
rect 296 99 298 123
rect 432 99 434 123
rect 568 99 570 123
rect 704 99 706 123
rect 840 99 842 123
rect 976 99 978 123
rect 1112 99 1114 123
rect 1934 122 1940 123
rect 1974 124 1980 125
rect 1996 124 1998 185
rect 2132 124 2134 185
rect 2268 124 2270 185
rect 2404 124 2406 185
rect 2540 124 2542 185
rect 2676 124 2678 185
rect 2812 124 2814 185
rect 2948 124 2950 185
rect 3084 124 3086 185
rect 3220 124 3222 185
rect 3356 124 3358 185
rect 3492 124 3494 185
rect 3628 124 3630 185
rect 3800 125 3802 185
rect 3840 137 3842 197
rect 3838 136 3844 137
rect 4292 136 4294 197
rect 4428 136 4430 197
rect 4564 136 4566 197
rect 4700 136 4702 197
rect 4836 136 4838 197
rect 4972 136 4974 197
rect 5108 136 5110 197
rect 5244 136 5246 197
rect 5380 136 5382 197
rect 5516 136 5518 197
rect 5664 137 5666 197
rect 5662 136 5668 137
rect 3838 132 3839 136
rect 3843 132 3844 136
rect 3838 131 3844 132
rect 4290 135 4296 136
rect 4290 131 4291 135
rect 4295 131 4296 135
rect 4290 130 4296 131
rect 4426 135 4432 136
rect 4426 131 4427 135
rect 4431 131 4432 135
rect 4426 130 4432 131
rect 4562 135 4568 136
rect 4562 131 4563 135
rect 4567 131 4568 135
rect 4562 130 4568 131
rect 4698 135 4704 136
rect 4698 131 4699 135
rect 4703 131 4704 135
rect 4698 130 4704 131
rect 4834 135 4840 136
rect 4834 131 4835 135
rect 4839 131 4840 135
rect 4834 130 4840 131
rect 4970 135 4976 136
rect 4970 131 4971 135
rect 4975 131 4976 135
rect 4970 130 4976 131
rect 5106 135 5112 136
rect 5106 131 5107 135
rect 5111 131 5112 135
rect 5106 130 5112 131
rect 5242 135 5248 136
rect 5242 131 5243 135
rect 5247 131 5248 135
rect 5242 130 5248 131
rect 5378 135 5384 136
rect 5378 131 5379 135
rect 5383 131 5384 135
rect 5378 130 5384 131
rect 5514 135 5520 136
rect 5514 131 5515 135
rect 5519 131 5520 135
rect 5662 132 5663 136
rect 5667 132 5668 136
rect 5662 131 5668 132
rect 5514 130 5520 131
rect 3798 124 3804 125
rect 1936 99 1938 122
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 4318 120 4324 121
rect 3798 119 3804 120
rect 3838 119 3844 120
rect 3626 118 3632 119
rect 3838 115 3839 119
rect 3843 115 3844 119
rect 4318 116 4319 120
rect 4323 116 4324 120
rect 4318 115 4324 116
rect 4454 120 4460 121
rect 4454 116 4455 120
rect 4459 116 4460 120
rect 4454 115 4460 116
rect 4590 120 4596 121
rect 4590 116 4591 120
rect 4595 116 4596 120
rect 4590 115 4596 116
rect 4726 120 4732 121
rect 4726 116 4727 120
rect 4731 116 4732 120
rect 4726 115 4732 116
rect 4862 120 4868 121
rect 4862 116 4863 120
rect 4867 116 4868 120
rect 4862 115 4868 116
rect 4998 120 5004 121
rect 4998 116 4999 120
rect 5003 116 5004 120
rect 4998 115 5004 116
rect 5134 120 5140 121
rect 5134 116 5135 120
rect 5139 116 5140 120
rect 5134 115 5140 116
rect 5270 120 5276 121
rect 5270 116 5271 120
rect 5275 116 5276 120
rect 5270 115 5276 116
rect 5406 120 5412 121
rect 5406 116 5407 120
rect 5411 116 5412 120
rect 5406 115 5412 116
rect 5542 120 5548 121
rect 5542 116 5543 120
rect 5547 116 5548 120
rect 5542 115 5548 116
rect 5662 119 5668 120
rect 5662 115 5663 119
rect 5667 115 5668 119
rect 3838 114 3844 115
rect 2022 108 2028 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2158 108 2164 109
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2430 108 2436 109
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2566 108 2572 109
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2838 108 2844 109
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2974 108 2980 109
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3110 108 3116 109
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3246 108 3252 109
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3382 108 3388 109
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3518 108 3524 109
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3654 108 3660 109
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 1974 102 1980 103
rect 111 98 115 99
rect 111 93 115 94
rect 159 98 163 99
rect 159 93 163 94
rect 295 98 299 99
rect 295 93 299 94
rect 431 98 435 99
rect 431 93 435 94
rect 567 98 571 99
rect 567 93 571 94
rect 703 98 707 99
rect 703 93 707 94
rect 839 98 843 99
rect 839 93 843 94
rect 975 98 979 99
rect 975 93 979 94
rect 1111 98 1115 99
rect 1111 93 1115 94
rect 1935 98 1939 99
rect 1935 93 1939 94
rect 1976 79 1978 102
rect 2024 79 2026 103
rect 2160 79 2162 103
rect 2296 79 2298 103
rect 2432 79 2434 103
rect 2568 79 2570 103
rect 2704 79 2706 103
rect 2840 79 2842 103
rect 2976 79 2978 103
rect 3112 79 3114 103
rect 3248 79 3250 103
rect 3384 79 3386 103
rect 3520 79 3522 103
rect 3656 79 3658 103
rect 3798 102 3804 103
rect 3800 79 3802 102
rect 3840 91 3842 114
rect 4320 91 4322 115
rect 4456 91 4458 115
rect 4592 91 4594 115
rect 4728 91 4730 115
rect 4864 91 4866 115
rect 5000 91 5002 115
rect 5136 91 5138 115
rect 5272 91 5274 115
rect 5408 91 5410 115
rect 5544 91 5546 115
rect 5662 114 5668 115
rect 5664 91 5666 114
rect 3839 90 3843 91
rect 3839 85 3843 86
rect 4319 90 4323 91
rect 4319 85 4323 86
rect 4455 90 4459 91
rect 4455 85 4459 86
rect 4591 90 4595 91
rect 4591 85 4595 86
rect 4727 90 4731 91
rect 4727 85 4731 86
rect 4863 90 4867 91
rect 4863 85 4867 86
rect 4999 90 5003 91
rect 4999 85 5003 86
rect 5135 90 5139 91
rect 5135 85 5139 86
rect 5271 90 5275 91
rect 5271 85 5275 86
rect 5407 90 5411 91
rect 5407 85 5411 86
rect 5543 90 5547 91
rect 5543 85 5547 86
rect 5663 90 5667 91
rect 5663 85 5667 86
rect 1975 78 1979 79
rect 1975 73 1979 74
rect 2023 78 2027 79
rect 2023 73 2027 74
rect 2159 78 2163 79
rect 2159 73 2163 74
rect 2295 78 2299 79
rect 2295 73 2299 74
rect 2431 78 2435 79
rect 2431 73 2435 74
rect 2567 78 2571 79
rect 2567 73 2571 74
rect 2703 78 2707 79
rect 2703 73 2707 74
rect 2839 78 2843 79
rect 2839 73 2843 74
rect 2975 78 2979 79
rect 2975 73 2979 74
rect 3111 78 3115 79
rect 3111 73 3115 74
rect 3247 78 3251 79
rect 3247 73 3251 74
rect 3383 78 3387 79
rect 3383 73 3387 74
rect 3519 78 3523 79
rect 3519 73 3523 74
rect 3655 78 3659 79
rect 3655 73 3659 74
rect 3799 78 3803 79
rect 3799 73 3803 74
<< m4c >>
rect 1975 5754 1979 5758
rect 2375 5754 2379 5758
rect 2511 5754 2515 5758
rect 2655 5754 2659 5758
rect 2807 5754 2811 5758
rect 2959 5754 2963 5758
rect 3119 5754 3123 5758
rect 3799 5754 3803 5758
rect 111 5714 115 5718
rect 159 5714 163 5718
rect 295 5714 299 5718
rect 431 5714 435 5718
rect 567 5714 571 5718
rect 703 5714 707 5718
rect 839 5714 843 5718
rect 975 5714 979 5718
rect 1935 5714 1939 5718
rect 3839 5678 3843 5682
rect 4335 5678 4339 5682
rect 4471 5678 4475 5682
rect 4607 5678 4611 5682
rect 4743 5678 4747 5682
rect 4879 5678 4883 5682
rect 5015 5678 5019 5682
rect 5663 5678 5667 5682
rect 1975 5642 1979 5646
rect 1995 5642 1999 5646
rect 2203 5642 2207 5646
rect 2347 5642 2351 5646
rect 2427 5642 2431 5646
rect 2483 5642 2487 5646
rect 2627 5642 2631 5646
rect 2651 5642 2655 5646
rect 2779 5642 2783 5646
rect 2867 5642 2871 5646
rect 2931 5642 2935 5646
rect 3075 5642 3079 5646
rect 3091 5642 3095 5646
rect 3275 5642 3279 5646
rect 3475 5642 3479 5646
rect 3651 5642 3655 5646
rect 3799 5642 3803 5646
rect 111 5574 115 5578
rect 131 5574 135 5578
rect 267 5574 271 5578
rect 403 5574 407 5578
rect 539 5574 543 5578
rect 619 5574 623 5578
rect 675 5574 679 5578
rect 755 5574 759 5578
rect 811 5574 815 5578
rect 899 5574 903 5578
rect 947 5574 951 5578
rect 1051 5574 1055 5578
rect 1203 5574 1207 5578
rect 1355 5574 1359 5578
rect 1507 5574 1511 5578
rect 1651 5574 1655 5578
rect 1787 5574 1791 5578
rect 1935 5574 1939 5578
rect 3839 5566 3843 5570
rect 4211 5566 4215 5570
rect 4307 5566 4311 5570
rect 4403 5566 4407 5570
rect 4443 5566 4447 5570
rect 4579 5566 4583 5570
rect 4595 5566 4599 5570
rect 4715 5566 4719 5570
rect 4795 5566 4799 5570
rect 4851 5566 4855 5570
rect 4987 5566 4991 5570
rect 4995 5566 4999 5570
rect 5195 5566 5199 5570
rect 5663 5566 5667 5570
rect 1975 5530 1979 5534
rect 2023 5530 2027 5534
rect 2231 5530 2235 5534
rect 2455 5530 2459 5534
rect 2679 5530 2683 5534
rect 2895 5530 2899 5534
rect 2951 5530 2955 5534
rect 3103 5530 3107 5534
rect 3255 5530 3259 5534
rect 3303 5530 3307 5534
rect 3415 5530 3419 5534
rect 3503 5530 3507 5534
rect 3679 5530 3683 5534
rect 3799 5530 3803 5534
rect 111 5454 115 5458
rect 591 5454 595 5458
rect 647 5454 651 5458
rect 727 5454 731 5458
rect 783 5454 787 5458
rect 863 5454 867 5458
rect 927 5454 931 5458
rect 999 5454 1003 5458
rect 1079 5454 1083 5458
rect 1135 5454 1139 5458
rect 1231 5454 1235 5458
rect 1271 5454 1275 5458
rect 1383 5454 1387 5458
rect 1407 5454 1411 5458
rect 1535 5454 1539 5458
rect 1543 5454 1547 5458
rect 1679 5454 1683 5458
rect 1815 5454 1819 5458
rect 1935 5454 1939 5458
rect 3839 5418 3843 5422
rect 4239 5418 4243 5422
rect 4303 5418 4307 5422
rect 4431 5418 4435 5422
rect 4519 5418 4523 5422
rect 4623 5418 4627 5422
rect 4735 5418 4739 5422
rect 4823 5418 4827 5422
rect 4951 5418 4955 5422
rect 5023 5418 5027 5422
rect 5175 5418 5179 5422
rect 5223 5418 5227 5422
rect 5399 5418 5403 5422
rect 5663 5418 5667 5422
rect 1975 5370 1979 5374
rect 2643 5370 2647 5374
rect 2811 5370 2815 5374
rect 2923 5370 2927 5374
rect 2979 5370 2983 5374
rect 3075 5370 3079 5374
rect 3139 5370 3143 5374
rect 3227 5370 3231 5374
rect 3307 5370 3311 5374
rect 3387 5370 3391 5374
rect 3475 5370 3479 5374
rect 3643 5370 3647 5374
rect 3799 5370 3803 5374
rect 111 5318 115 5322
rect 411 5318 415 5322
rect 563 5318 567 5322
rect 587 5318 591 5322
rect 699 5318 703 5322
rect 763 5318 767 5322
rect 835 5318 839 5322
rect 939 5318 943 5322
rect 971 5318 975 5322
rect 1107 5318 1111 5322
rect 1243 5318 1247 5322
rect 1275 5318 1279 5322
rect 1379 5318 1383 5322
rect 1443 5318 1447 5322
rect 1515 5318 1519 5322
rect 1611 5318 1615 5322
rect 1651 5318 1655 5322
rect 1787 5318 1791 5322
rect 1935 5318 1939 5322
rect 3839 5274 3843 5278
rect 4275 5274 4279 5278
rect 4371 5274 4375 5278
rect 4491 5274 4495 5278
rect 4563 5274 4567 5278
rect 4707 5274 4711 5278
rect 4771 5274 4775 5278
rect 4923 5274 4927 5278
rect 4979 5274 4983 5278
rect 5147 5274 5151 5278
rect 5195 5274 5199 5278
rect 5371 5274 5375 5278
rect 5419 5274 5423 5278
rect 5663 5274 5667 5278
rect 1975 5258 1979 5262
rect 2511 5258 2515 5262
rect 2671 5258 2675 5262
rect 2687 5258 2691 5262
rect 2839 5258 2843 5262
rect 2863 5258 2867 5262
rect 3007 5258 3011 5262
rect 3039 5258 3043 5262
rect 3167 5258 3171 5262
rect 3207 5258 3211 5262
rect 3335 5258 3339 5262
rect 3367 5258 3371 5262
rect 3503 5258 3507 5262
rect 3535 5258 3539 5262
rect 3671 5258 3675 5262
rect 3679 5258 3683 5262
rect 3799 5258 3803 5262
rect 111 5198 115 5202
rect 207 5198 211 5202
rect 343 5198 347 5202
rect 439 5198 443 5202
rect 479 5198 483 5202
rect 615 5198 619 5202
rect 751 5198 755 5202
rect 791 5198 795 5202
rect 887 5198 891 5202
rect 967 5198 971 5202
rect 1023 5198 1027 5202
rect 1135 5198 1139 5202
rect 1303 5198 1307 5202
rect 1471 5198 1475 5202
rect 1639 5198 1643 5202
rect 1815 5198 1819 5202
rect 1935 5198 1939 5202
rect 1975 5138 1979 5142
rect 2139 5138 2143 5142
rect 2307 5138 2311 5142
rect 2483 5138 2487 5142
rect 2491 5138 2495 5142
rect 2659 5138 2663 5142
rect 2691 5138 2695 5142
rect 2835 5138 2839 5142
rect 2915 5138 2919 5142
rect 3011 5138 3015 5142
rect 3163 5138 3167 5142
rect 3179 5138 3183 5142
rect 3339 5138 3343 5142
rect 3419 5138 3423 5142
rect 3507 5138 3511 5142
rect 3651 5138 3655 5142
rect 3799 5138 3803 5142
rect 3839 5138 3843 5142
rect 3887 5138 3891 5142
rect 4087 5138 4091 5142
rect 4311 5138 4315 5142
rect 4399 5138 4403 5142
rect 4535 5138 4539 5142
rect 4591 5138 4595 5142
rect 4759 5138 4763 5142
rect 4799 5138 4803 5142
rect 4983 5138 4987 5142
rect 5007 5138 5011 5142
rect 5207 5138 5211 5142
rect 5223 5138 5227 5142
rect 5439 5138 5443 5142
rect 5447 5138 5451 5142
rect 5663 5138 5667 5142
rect 111 5066 115 5070
rect 147 5066 151 5070
rect 179 5066 183 5070
rect 315 5066 319 5070
rect 339 5066 343 5070
rect 451 5066 455 5070
rect 531 5066 535 5070
rect 587 5066 591 5070
rect 723 5066 727 5070
rect 731 5066 735 5070
rect 859 5066 863 5070
rect 931 5066 935 5070
rect 995 5066 999 5070
rect 1131 5066 1135 5070
rect 1935 5066 1939 5070
rect 3839 5010 3843 5014
rect 3859 5010 3863 5014
rect 3995 5010 3999 5014
rect 4059 5010 4063 5014
rect 4131 5010 4135 5014
rect 4283 5010 4287 5014
rect 4443 5010 4447 5014
rect 4507 5010 4511 5014
rect 4611 5010 4615 5014
rect 4731 5010 4735 5014
rect 4787 5010 4791 5014
rect 4955 5010 4959 5014
rect 4971 5010 4975 5014
rect 5155 5010 5159 5014
rect 5179 5010 5183 5014
rect 5339 5010 5343 5014
rect 5411 5010 5415 5014
rect 5515 5010 5519 5014
rect 5663 5010 5667 5014
rect 1975 5002 1979 5006
rect 2023 5002 2027 5006
rect 2167 5002 2171 5006
rect 2335 5002 2339 5006
rect 2351 5002 2355 5006
rect 2519 5002 2523 5006
rect 2543 5002 2547 5006
rect 2719 5002 2723 5006
rect 2751 5002 2755 5006
rect 2943 5002 2947 5006
rect 2967 5002 2971 5006
rect 3183 5002 3187 5006
rect 3191 5002 3195 5006
rect 3447 5002 3451 5006
rect 3679 5002 3683 5006
rect 3799 5002 3803 5006
rect 111 4942 115 4946
rect 159 4942 163 4946
rect 175 4942 179 4946
rect 367 4942 371 4946
rect 391 4942 395 4946
rect 559 4942 563 4946
rect 647 4942 651 4946
rect 759 4942 763 4946
rect 895 4942 899 4946
rect 959 4942 963 4946
rect 1135 4942 1139 4946
rect 1159 4942 1163 4946
rect 1367 4942 1371 4946
rect 1599 4942 1603 4946
rect 1815 4942 1819 4946
rect 1935 4942 1939 4946
rect 1975 4882 1979 4886
rect 1995 4882 1999 4886
rect 2139 4882 2143 4886
rect 2323 4882 2327 4886
rect 2515 4882 2519 4886
rect 2667 4882 2671 4886
rect 2723 4882 2727 4886
rect 2939 4882 2943 4886
rect 3019 4882 3023 4886
rect 3155 4882 3159 4886
rect 3371 4882 3375 4886
rect 3799 4882 3803 4886
rect 3839 4882 3843 4886
rect 3887 4882 3891 4886
rect 3943 4882 3947 4886
rect 4023 4882 4027 4886
rect 4159 4882 4163 4886
rect 4183 4882 4187 4886
rect 4311 4882 4315 4886
rect 4431 4882 4435 4886
rect 4471 4882 4475 4886
rect 4639 4882 4643 4886
rect 4687 4882 4691 4886
rect 4815 4882 4819 4886
rect 4959 4882 4963 4886
rect 4999 4882 5003 4886
rect 5183 4882 5187 4886
rect 5239 4882 5243 4886
rect 5367 4882 5371 4886
rect 5519 4882 5523 4886
rect 5543 4882 5547 4886
rect 5663 4882 5667 4886
rect 111 4830 115 4834
rect 131 4830 135 4834
rect 363 4830 367 4834
rect 475 4830 479 4834
rect 619 4830 623 4834
rect 859 4830 863 4834
rect 867 4830 871 4834
rect 1107 4830 1111 4834
rect 1251 4830 1255 4834
rect 1339 4830 1343 4834
rect 1571 4830 1575 4834
rect 1643 4830 1647 4834
rect 1787 4830 1791 4834
rect 1935 4830 1939 4834
rect 3839 4762 3843 4766
rect 3915 4762 3919 4766
rect 3939 4762 3943 4766
rect 4155 4762 4159 4766
rect 4179 4762 4183 4766
rect 4403 4762 4407 4766
rect 4435 4762 4439 4766
rect 4659 4762 4663 4766
rect 4691 4762 4695 4766
rect 4931 4762 4935 4766
rect 4955 4762 4959 4766
rect 5211 4762 5215 4766
rect 5227 4762 5231 4766
rect 5491 4762 5495 4766
rect 5507 4762 5511 4766
rect 5663 4762 5667 4766
rect 1975 4722 1979 4726
rect 2023 4722 2027 4726
rect 2079 4722 2083 4726
rect 2231 4722 2235 4726
rect 2351 4722 2355 4726
rect 2391 4722 2395 4726
rect 2559 4722 2563 4726
rect 2695 4722 2699 4726
rect 2727 4722 2731 4726
rect 2903 4722 2907 4726
rect 3047 4722 3051 4726
rect 3079 4722 3083 4726
rect 3255 4722 3259 4726
rect 3399 4722 3403 4726
rect 3439 4722 3443 4726
rect 3623 4722 3627 4726
rect 3799 4722 3803 4726
rect 111 4698 115 4702
rect 159 4698 163 4702
rect 295 4698 299 4702
rect 431 4698 435 4702
rect 503 4698 507 4702
rect 567 4698 571 4702
rect 703 4698 707 4702
rect 887 4698 891 4702
rect 1279 4698 1283 4702
rect 1671 4698 1675 4702
rect 1935 4698 1939 4702
rect 3839 4646 3843 4650
rect 3967 4646 3971 4650
rect 4175 4646 4179 4650
rect 4207 4646 4211 4650
rect 4455 4646 4459 4650
rect 4463 4646 4467 4650
rect 4719 4646 4723 4650
rect 4735 4646 4739 4650
rect 4983 4646 4987 4650
rect 5015 4646 5019 4650
rect 5255 4646 5259 4650
rect 5303 4646 5307 4650
rect 5535 4646 5539 4650
rect 5663 4646 5667 4650
rect 1975 4606 1979 4610
rect 2051 4606 2055 4610
rect 2123 4606 2127 4610
rect 2203 4606 2207 4610
rect 2275 4606 2279 4610
rect 2363 4606 2367 4610
rect 2443 4606 2447 4610
rect 2531 4606 2535 4610
rect 2611 4606 2615 4610
rect 2699 4606 2703 4610
rect 2787 4606 2791 4610
rect 2875 4606 2879 4610
rect 2963 4606 2967 4610
rect 3051 4606 3055 4610
rect 3139 4606 3143 4610
rect 3227 4606 3231 4610
rect 3315 4606 3319 4610
rect 3411 4606 3415 4610
rect 3491 4606 3495 4610
rect 3595 4606 3599 4610
rect 3651 4606 3655 4610
rect 3799 4606 3803 4610
rect 111 4570 115 4574
rect 131 4570 135 4574
rect 267 4570 271 4574
rect 291 4570 295 4574
rect 403 4570 407 4574
rect 427 4570 431 4574
rect 539 4570 543 4574
rect 563 4570 567 4574
rect 675 4570 679 4574
rect 699 4570 703 4574
rect 835 4570 839 4574
rect 1935 4570 1939 4574
rect 3839 4530 3843 4534
rect 3859 4530 3863 4534
rect 4147 4530 4151 4534
rect 4155 4530 4159 4534
rect 4427 4530 4431 4534
rect 4483 4530 4487 4534
rect 4707 4530 4711 4534
rect 4819 4530 4823 4534
rect 4987 4530 4991 4534
rect 5163 4530 5167 4534
rect 5275 4530 5279 4534
rect 5515 4530 5519 4534
rect 5663 4530 5667 4534
rect 1975 4486 1979 4490
rect 2023 4486 2027 4490
rect 2151 4486 2155 4490
rect 2159 4486 2163 4490
rect 2295 4486 2299 4490
rect 2303 4486 2307 4490
rect 2431 4486 2435 4490
rect 2471 4486 2475 4490
rect 2567 4486 2571 4490
rect 2639 4486 2643 4490
rect 2703 4486 2707 4490
rect 2815 4486 2819 4490
rect 2839 4486 2843 4490
rect 2975 4486 2979 4490
rect 2991 4486 2995 4490
rect 3167 4486 3171 4490
rect 3343 4486 3347 4490
rect 3519 4486 3523 4490
rect 3679 4486 3683 4490
rect 3799 4486 3803 4490
rect 111 4442 115 4446
rect 319 4442 323 4446
rect 455 4442 459 4446
rect 519 4442 523 4446
rect 591 4442 595 4446
rect 727 4442 731 4446
rect 743 4442 747 4446
rect 863 4442 867 4446
rect 991 4442 995 4446
rect 1263 4442 1267 4446
rect 1551 4442 1555 4446
rect 1815 4442 1819 4446
rect 1935 4442 1939 4446
rect 3839 4418 3843 4422
rect 3887 4418 3891 4422
rect 4143 4418 4147 4422
rect 4183 4418 4187 4422
rect 4423 4418 4427 4422
rect 4511 4418 4515 4422
rect 4703 4418 4707 4422
rect 4847 4418 4851 4422
rect 4983 4418 4987 4422
rect 5191 4418 5195 4422
rect 5263 4418 5267 4422
rect 5543 4418 5547 4422
rect 5663 4418 5667 4422
rect 1975 4358 1979 4362
rect 1995 4358 1999 4362
rect 2131 4358 2135 4362
rect 2267 4358 2271 4362
rect 2403 4358 2407 4362
rect 2539 4358 2543 4362
rect 2675 4358 2679 4362
rect 2779 4358 2783 4362
rect 2811 4358 2815 4362
rect 2947 4358 2951 4362
rect 2995 4358 2999 4362
rect 3219 4358 3223 4362
rect 3443 4358 3447 4362
rect 3651 4358 3655 4362
rect 3799 4358 3803 4362
rect 111 4330 115 4334
rect 491 4330 495 4334
rect 563 4330 567 4334
rect 699 4330 703 4334
rect 715 4330 719 4334
rect 835 4330 839 4334
rect 963 4330 967 4334
rect 971 4330 975 4334
rect 1107 4330 1111 4334
rect 1235 4330 1239 4334
rect 1243 4330 1247 4334
rect 1379 4330 1383 4334
rect 1515 4330 1519 4334
rect 1523 4330 1527 4334
rect 1651 4330 1655 4334
rect 1787 4330 1791 4334
rect 1935 4330 1939 4334
rect 3839 4294 3843 4298
rect 3859 4294 3863 4298
rect 4115 4294 4119 4298
rect 4395 4294 4399 4298
rect 4571 4294 4575 4298
rect 4675 4294 4679 4298
rect 4739 4294 4743 4298
rect 4915 4294 4919 4298
rect 4955 4294 4959 4298
rect 5107 4294 5111 4298
rect 5235 4294 5239 4298
rect 5307 4294 5311 4298
rect 5515 4294 5519 4298
rect 5663 4294 5667 4298
rect 1975 4218 1979 4222
rect 2807 4218 2811 4222
rect 2951 4218 2955 4222
rect 3023 4218 3027 4222
rect 3095 4218 3099 4222
rect 3239 4218 3243 4222
rect 3247 4218 3251 4222
rect 3391 4218 3395 4222
rect 3471 4218 3475 4222
rect 3543 4218 3547 4222
rect 3679 4218 3683 4222
rect 3799 4218 3803 4222
rect 111 4206 115 4210
rect 591 4206 595 4210
rect 727 4206 731 4210
rect 863 4206 867 4210
rect 999 4206 1003 4210
rect 1135 4206 1139 4210
rect 1271 4206 1275 4210
rect 1407 4206 1411 4210
rect 1543 4206 1547 4210
rect 1679 4206 1683 4210
rect 1815 4206 1819 4210
rect 1935 4206 1939 4210
rect 3839 4182 3843 4186
rect 4599 4182 4603 4186
rect 4655 4182 4659 4186
rect 4767 4182 4771 4186
rect 4815 4182 4819 4186
rect 4943 4182 4947 4186
rect 4983 4182 4987 4186
rect 5135 4182 5139 4186
rect 5167 4182 5171 4186
rect 5335 4182 5339 4186
rect 5359 4182 5363 4186
rect 5543 4182 5547 4186
rect 5663 4182 5667 4186
rect 111 4094 115 4098
rect 563 4094 567 4098
rect 699 4094 703 4098
rect 835 4094 839 4098
rect 971 4094 975 4098
rect 1107 4094 1111 4098
rect 1243 4094 1247 4098
rect 1379 4094 1383 4098
rect 1515 4094 1519 4098
rect 1651 4094 1655 4098
rect 1787 4094 1791 4098
rect 1935 4094 1939 4098
rect 1975 4070 1979 4074
rect 2899 4070 2903 4074
rect 2923 4070 2927 4074
rect 3043 4070 3047 4074
rect 3067 4070 3071 4074
rect 3187 4070 3191 4074
rect 3211 4070 3215 4074
rect 3339 4070 3343 4074
rect 3363 4070 3367 4074
rect 3491 4070 3495 4074
rect 3515 4070 3519 4074
rect 3643 4070 3647 4074
rect 3651 4070 3655 4074
rect 3799 4070 3803 4074
rect 3839 4034 3843 4038
rect 4627 4034 4631 4038
rect 4787 4034 4791 4038
rect 4939 4034 4943 4038
rect 4955 4034 4959 4038
rect 5075 4034 5079 4038
rect 5139 4034 5143 4038
rect 5211 4034 5215 4038
rect 5331 4034 5335 4038
rect 5347 4034 5351 4038
rect 5515 4034 5519 4038
rect 5663 4034 5667 4038
rect 111 3978 115 3982
rect 695 3978 699 3982
rect 727 3978 731 3982
rect 831 3978 835 3982
rect 863 3978 867 3982
rect 967 3978 971 3982
rect 999 3978 1003 3982
rect 1111 3978 1115 3982
rect 1135 3978 1139 3982
rect 1255 3978 1259 3982
rect 1271 3978 1275 3982
rect 1399 3978 1403 3982
rect 1407 3978 1411 3982
rect 1543 3978 1547 3982
rect 1679 3978 1683 3982
rect 1815 3978 1819 3982
rect 1935 3978 1939 3982
rect 1975 3930 1979 3934
rect 2759 3930 2763 3934
rect 2911 3930 2915 3934
rect 2927 3930 2931 3934
rect 3071 3930 3075 3934
rect 3215 3930 3219 3934
rect 3239 3930 3243 3934
rect 3367 3930 3371 3934
rect 3415 3930 3419 3934
rect 3519 3930 3523 3934
rect 3591 3930 3595 3934
rect 3671 3930 3675 3934
rect 3799 3930 3803 3934
rect 3839 3922 3843 3926
rect 4687 3922 4691 3926
rect 4847 3922 4851 3926
rect 4967 3922 4971 3926
rect 5015 3922 5019 3926
rect 5103 3922 5107 3926
rect 5191 3922 5195 3926
rect 5239 3922 5243 3926
rect 5375 3922 5379 3926
rect 5543 3922 5547 3926
rect 5663 3922 5667 3926
rect 111 3862 115 3866
rect 435 3862 439 3866
rect 619 3862 623 3866
rect 667 3862 671 3866
rect 803 3862 807 3866
rect 819 3862 823 3866
rect 939 3862 943 3866
rect 1027 3862 1031 3866
rect 1083 3862 1087 3866
rect 1227 3862 1231 3866
rect 1251 3862 1255 3866
rect 1371 3862 1375 3866
rect 1483 3862 1487 3866
rect 1515 3862 1519 3866
rect 1651 3862 1655 3866
rect 1723 3862 1727 3866
rect 1787 3862 1791 3866
rect 1935 3862 1939 3866
rect 1975 3810 1979 3814
rect 2115 3810 2119 3814
rect 2251 3810 2255 3814
rect 2387 3810 2391 3814
rect 2523 3810 2527 3814
rect 2659 3810 2663 3814
rect 2731 3810 2735 3814
rect 2795 3810 2799 3814
rect 2883 3810 2887 3814
rect 2939 3810 2943 3814
rect 3043 3810 3047 3814
rect 3083 3810 3087 3814
rect 3211 3810 3215 3814
rect 3235 3810 3239 3814
rect 3387 3810 3391 3814
rect 3395 3810 3399 3814
rect 3555 3810 3559 3814
rect 3563 3810 3567 3814
rect 3799 3810 3803 3814
rect 3839 3810 3843 3814
rect 4411 3810 4415 3814
rect 4619 3810 4623 3814
rect 4659 3810 4663 3814
rect 4819 3810 4823 3814
rect 4835 3810 4839 3814
rect 4987 3810 4991 3814
rect 5067 3810 5071 3814
rect 5163 3810 5167 3814
rect 5299 3810 5303 3814
rect 5347 3810 5351 3814
rect 5515 3810 5519 3814
rect 5663 3810 5667 3814
rect 111 3746 115 3750
rect 231 3746 235 3750
rect 431 3746 435 3750
rect 463 3746 467 3750
rect 647 3746 651 3750
rect 655 3746 659 3750
rect 847 3746 851 3750
rect 895 3746 899 3750
rect 1055 3746 1059 3750
rect 1151 3746 1155 3750
rect 1279 3746 1283 3750
rect 1415 3746 1419 3750
rect 1511 3746 1515 3750
rect 1679 3746 1683 3750
rect 1751 3746 1755 3750
rect 1935 3746 1939 3750
rect 1975 3690 1979 3694
rect 2143 3690 2147 3694
rect 2231 3690 2235 3694
rect 2279 3690 2283 3694
rect 2415 3690 2419 3694
rect 2447 3690 2451 3694
rect 2551 3690 2555 3694
rect 2663 3690 2667 3694
rect 2687 3690 2691 3694
rect 2823 3690 2827 3694
rect 2871 3690 2875 3694
rect 2967 3690 2971 3694
rect 3079 3690 3083 3694
rect 3111 3690 3115 3694
rect 3263 3690 3267 3694
rect 3287 3690 3291 3694
rect 3423 3690 3427 3694
rect 3495 3690 3499 3694
rect 3583 3690 3587 3694
rect 3679 3690 3683 3694
rect 3799 3690 3803 3694
rect 3839 3674 3843 3678
rect 3887 3674 3891 3678
rect 4047 3674 4051 3678
rect 4247 3674 4251 3678
rect 4439 3674 4443 3678
rect 4479 3674 4483 3678
rect 4647 3674 4651 3678
rect 4727 3674 4731 3678
rect 4863 3674 4867 3678
rect 4999 3674 5003 3678
rect 5095 3674 5099 3678
rect 5279 3674 5283 3678
rect 5327 3674 5331 3678
rect 5543 3674 5547 3678
rect 5663 3674 5667 3678
rect 111 3626 115 3630
rect 131 3626 135 3630
rect 203 3626 207 3630
rect 315 3626 319 3630
rect 403 3626 407 3630
rect 539 3626 543 3630
rect 627 3626 631 3630
rect 787 3626 791 3630
rect 867 3626 871 3630
rect 1043 3626 1047 3630
rect 1123 3626 1127 3630
rect 1315 3626 1319 3630
rect 1387 3626 1391 3630
rect 1587 3626 1591 3630
rect 1651 3626 1655 3630
rect 1935 3626 1939 3630
rect 1975 3562 1979 3566
rect 2163 3562 2167 3566
rect 2203 3562 2207 3566
rect 2299 3562 2303 3566
rect 2419 3562 2423 3566
rect 2435 3562 2439 3566
rect 2571 3562 2575 3566
rect 2635 3562 2639 3566
rect 2843 3562 2847 3566
rect 3051 3562 3055 3566
rect 3259 3562 3263 3566
rect 3467 3562 3471 3566
rect 3651 3562 3655 3566
rect 3799 3562 3803 3566
rect 111 3502 115 3506
rect 159 3502 163 3506
rect 335 3502 339 3506
rect 343 3502 347 3506
rect 551 3502 555 3506
rect 567 3502 571 3506
rect 791 3502 795 3506
rect 815 3502 819 3506
rect 1039 3502 1043 3506
rect 1071 3502 1075 3506
rect 1295 3502 1299 3506
rect 1343 3502 1347 3506
rect 1559 3502 1563 3506
rect 1615 3502 1619 3506
rect 1935 3502 1939 3506
rect 3839 3550 3843 3554
rect 3859 3550 3863 3554
rect 3995 3550 3999 3554
rect 4019 3550 4023 3554
rect 4131 3550 4135 3554
rect 4219 3550 4223 3554
rect 4267 3550 4271 3554
rect 4403 3550 4407 3554
rect 4451 3550 4455 3554
rect 4539 3550 4543 3554
rect 4699 3550 4703 3554
rect 4891 3550 4895 3554
rect 4971 3550 4975 3554
rect 5099 3550 5103 3554
rect 5251 3550 5255 3554
rect 5315 3550 5319 3554
rect 5515 3550 5519 3554
rect 5663 3550 5667 3554
rect 3839 3430 3843 3434
rect 3887 3430 3891 3434
rect 4023 3430 4027 3434
rect 4159 3430 4163 3434
rect 4295 3430 4299 3434
rect 4431 3430 4435 3434
rect 4567 3430 4571 3434
rect 4583 3430 4587 3434
rect 4727 3430 4731 3434
rect 4759 3430 4763 3434
rect 4919 3430 4923 3434
rect 4951 3430 4955 3434
rect 5127 3430 5131 3434
rect 5151 3430 5155 3434
rect 5343 3430 5347 3434
rect 5359 3430 5363 3434
rect 5543 3430 5547 3434
rect 5663 3430 5667 3434
rect 1975 3414 1979 3418
rect 2191 3414 2195 3418
rect 2231 3414 2235 3418
rect 2327 3414 2331 3418
rect 2463 3414 2467 3418
rect 2583 3414 2587 3418
rect 2599 3414 2603 3418
rect 2951 3414 2955 3418
rect 3327 3414 3331 3418
rect 3679 3414 3683 3418
rect 3799 3414 3803 3418
rect 111 3382 115 3386
rect 131 3382 135 3386
rect 299 3382 303 3386
rect 307 3382 311 3386
rect 507 3382 511 3386
rect 523 3382 527 3386
rect 731 3382 735 3386
rect 763 3382 767 3386
rect 971 3382 975 3386
rect 1011 3382 1015 3386
rect 1219 3382 1223 3386
rect 1267 3382 1271 3386
rect 1475 3382 1479 3386
rect 1531 3382 1535 3386
rect 1935 3382 1939 3386
rect 1975 3302 1979 3306
rect 2203 3302 2207 3306
rect 2251 3302 2255 3306
rect 2475 3302 2479 3306
rect 2555 3302 2559 3306
rect 2691 3302 2695 3306
rect 2899 3302 2903 3306
rect 2923 3302 2927 3306
rect 3099 3302 3103 3306
rect 3291 3302 3295 3306
rect 3299 3302 3303 3306
rect 3483 3302 3487 3306
rect 3651 3302 3655 3306
rect 3799 3302 3803 3306
rect 3839 3302 3843 3306
rect 3859 3302 3863 3306
rect 3995 3302 3999 3306
rect 4131 3302 4135 3306
rect 4267 3302 4271 3306
rect 4403 3302 4407 3306
rect 4555 3302 4559 3306
rect 4691 3302 4695 3306
rect 4731 3302 4735 3306
rect 4827 3302 4831 3306
rect 4923 3302 4927 3306
rect 4963 3302 4967 3306
rect 5099 3302 5103 3306
rect 5123 3302 5127 3306
rect 5235 3302 5239 3306
rect 5331 3302 5335 3306
rect 5515 3302 5519 3306
rect 5663 3302 5667 3306
rect 111 3266 115 3270
rect 159 3266 163 3270
rect 239 3266 243 3270
rect 327 3266 331 3270
rect 463 3266 467 3270
rect 535 3266 539 3270
rect 703 3266 707 3270
rect 759 3266 763 3270
rect 951 3266 955 3270
rect 999 3266 1003 3270
rect 1199 3266 1203 3270
rect 1247 3266 1251 3270
rect 1455 3266 1459 3270
rect 1503 3266 1507 3270
rect 1935 3266 1939 3270
rect 1975 3182 1979 3186
rect 2095 3182 2099 3186
rect 2279 3182 2283 3186
rect 2295 3182 2299 3186
rect 2487 3182 2491 3186
rect 2503 3182 2507 3186
rect 2679 3182 2683 3186
rect 2719 3182 2723 3186
rect 2871 3182 2875 3186
rect 2927 3182 2931 3186
rect 3055 3182 3059 3186
rect 3127 3182 3131 3186
rect 3231 3182 3235 3186
rect 3319 3182 3323 3186
rect 3415 3182 3419 3186
rect 3511 3182 3515 3186
rect 3599 3182 3603 3186
rect 3679 3182 3683 3186
rect 3799 3182 3803 3186
rect 3839 3182 3843 3186
rect 4719 3182 4723 3186
rect 4855 3182 4859 3186
rect 4863 3182 4867 3186
rect 4991 3182 4995 3186
rect 4999 3182 5003 3186
rect 5127 3182 5131 3186
rect 5135 3182 5139 3186
rect 5263 3182 5267 3186
rect 5271 3182 5275 3186
rect 5407 3182 5411 3186
rect 5543 3182 5547 3186
rect 5663 3182 5667 3186
rect 111 3150 115 3154
rect 211 3150 215 3154
rect 379 3150 383 3154
rect 435 3150 439 3154
rect 563 3150 567 3154
rect 675 3150 679 3154
rect 755 3150 759 3154
rect 923 3150 927 3154
rect 955 3150 959 3154
rect 1163 3150 1167 3154
rect 1171 3150 1175 3154
rect 1371 3150 1375 3154
rect 1427 3150 1431 3154
rect 1935 3150 1939 3154
rect 1975 3058 1979 3062
rect 1995 3058 1999 3062
rect 2067 3058 2071 3062
rect 2131 3058 2135 3062
rect 2267 3058 2271 3062
rect 2403 3058 2407 3062
rect 2459 3058 2463 3062
rect 2539 3058 2543 3062
rect 2651 3058 2655 3062
rect 2683 3058 2687 3062
rect 2835 3058 2839 3062
rect 2843 3058 2847 3062
rect 2987 3058 2991 3062
rect 3027 3058 3031 3062
rect 3139 3058 3143 3062
rect 3203 3058 3207 3062
rect 3291 3058 3295 3062
rect 3387 3058 3391 3062
rect 3571 3058 3575 3062
rect 3799 3058 3803 3062
rect 3839 3058 3843 3062
rect 4483 3058 4487 3062
rect 4635 3058 4639 3062
rect 4803 3058 4807 3062
rect 4835 3058 4839 3062
rect 4971 3058 4975 3062
rect 4979 3058 4983 3062
rect 5107 3058 5111 3062
rect 5163 3058 5167 3062
rect 5243 3058 5247 3062
rect 5347 3058 5351 3062
rect 5379 3058 5383 3062
rect 5515 3058 5519 3062
rect 5663 3058 5667 3062
rect 111 3022 115 3026
rect 407 3022 411 3026
rect 575 3022 579 3026
rect 591 3022 595 3026
rect 783 3022 787 3026
rect 799 3022 803 3026
rect 983 3022 987 3026
rect 1047 3022 1051 3026
rect 1191 3022 1195 3026
rect 1303 3022 1307 3026
rect 1399 3022 1403 3026
rect 1567 3022 1571 3026
rect 1815 3022 1819 3026
rect 1935 3022 1939 3026
rect 1975 2946 1979 2950
rect 2023 2946 2027 2950
rect 2159 2946 2163 2950
rect 2295 2946 2299 2950
rect 2431 2946 2435 2950
rect 2567 2946 2571 2950
rect 2591 2946 2595 2950
rect 2711 2946 2715 2950
rect 2863 2946 2867 2950
rect 2887 2946 2891 2950
rect 3015 2946 3019 2950
rect 3167 2946 3171 2950
rect 3183 2946 3187 2950
rect 3319 2946 3323 2950
rect 3799 2946 3803 2950
rect 3839 2922 3843 2926
rect 4047 2922 4051 2926
rect 4295 2922 4299 2926
rect 4511 2922 4515 2926
rect 4583 2922 4587 2926
rect 4663 2922 4667 2926
rect 4831 2922 4835 2926
rect 4895 2922 4899 2926
rect 5007 2922 5011 2926
rect 5191 2922 5195 2926
rect 5231 2922 5235 2926
rect 5375 2922 5379 2926
rect 5543 2922 5547 2926
rect 5663 2922 5667 2926
rect 111 2902 115 2906
rect 427 2902 431 2906
rect 547 2902 551 2906
rect 563 2902 567 2906
rect 699 2902 703 2906
rect 771 2902 775 2906
rect 835 2902 839 2906
rect 971 2902 975 2906
rect 1019 2902 1023 2906
rect 1107 2902 1111 2906
rect 1243 2902 1247 2906
rect 1275 2902 1279 2906
rect 1379 2902 1383 2906
rect 1515 2902 1519 2906
rect 1539 2902 1543 2906
rect 1651 2902 1655 2906
rect 1787 2902 1791 2906
rect 1935 2902 1939 2906
rect 111 2782 115 2786
rect 455 2782 459 2786
rect 463 2782 467 2786
rect 591 2782 595 2786
rect 623 2782 627 2786
rect 727 2782 731 2786
rect 783 2782 787 2786
rect 863 2782 867 2786
rect 935 2782 939 2786
rect 999 2782 1003 2786
rect 1087 2782 1091 2786
rect 1135 2782 1139 2786
rect 1239 2782 1243 2786
rect 1271 2782 1275 2786
rect 1383 2782 1387 2786
rect 1407 2782 1411 2786
rect 1535 2782 1539 2786
rect 1543 2782 1547 2786
rect 1679 2782 1683 2786
rect 1815 2782 1819 2786
rect 1935 2782 1939 2786
rect 3839 2806 3843 2810
rect 3859 2806 3863 2810
rect 3995 2806 3999 2810
rect 4019 2806 4023 2810
rect 4131 2806 4135 2810
rect 4267 2806 4271 2810
rect 4403 2806 4407 2810
rect 4539 2806 4543 2810
rect 4555 2806 4559 2810
rect 4675 2806 4679 2810
rect 4811 2806 4815 2810
rect 4867 2806 4871 2810
rect 5203 2806 5207 2810
rect 5515 2806 5519 2810
rect 5663 2806 5667 2810
rect 1975 2778 1979 2782
rect 1995 2778 1999 2782
rect 2267 2778 2271 2782
rect 2563 2778 2567 2782
rect 2859 2778 2863 2782
rect 3059 2778 3063 2782
rect 3155 2778 3159 2782
rect 3195 2778 3199 2782
rect 3331 2778 3335 2782
rect 3799 2778 3803 2782
rect 111 2666 115 2670
rect 355 2666 359 2670
rect 435 2666 439 2670
rect 539 2666 543 2670
rect 595 2666 599 2670
rect 715 2666 719 2670
rect 755 2666 759 2670
rect 883 2666 887 2670
rect 907 2666 911 2670
rect 1043 2666 1047 2670
rect 1059 2666 1063 2670
rect 1203 2666 1207 2670
rect 1211 2666 1215 2670
rect 1355 2666 1359 2670
rect 1507 2666 1511 2670
rect 1651 2666 1655 2670
rect 1787 2666 1791 2670
rect 1935 2666 1939 2670
rect 3839 2694 3843 2698
rect 3887 2694 3891 2698
rect 4023 2694 4027 2698
rect 4055 2694 4059 2698
rect 4159 2694 4163 2698
rect 4295 2694 4299 2698
rect 4303 2694 4307 2698
rect 4431 2694 4435 2698
rect 4567 2694 4571 2698
rect 4583 2694 4587 2698
rect 4703 2694 4707 2698
rect 4839 2694 4843 2698
rect 4895 2694 4899 2698
rect 5231 2694 5235 2698
rect 5543 2694 5547 2698
rect 5663 2694 5667 2698
rect 1975 2642 1979 2646
rect 3087 2642 3091 2646
rect 3135 2642 3139 2646
rect 3223 2642 3227 2646
rect 3271 2642 3275 2646
rect 3359 2642 3363 2646
rect 3407 2642 3411 2646
rect 3543 2642 3547 2646
rect 3679 2642 3683 2646
rect 3799 2642 3803 2646
rect 111 2554 115 2558
rect 231 2554 235 2558
rect 383 2554 387 2558
rect 423 2554 427 2558
rect 567 2554 571 2558
rect 623 2554 627 2558
rect 743 2554 747 2558
rect 823 2554 827 2558
rect 911 2554 915 2558
rect 1023 2554 1027 2558
rect 1071 2554 1075 2558
rect 1223 2554 1227 2558
rect 1231 2554 1235 2558
rect 1383 2554 1387 2558
rect 1423 2554 1427 2558
rect 1535 2554 1539 2558
rect 1631 2554 1635 2558
rect 1679 2554 1683 2558
rect 1815 2554 1819 2558
rect 1935 2554 1939 2558
rect 3839 2578 3843 2582
rect 4027 2578 4031 2582
rect 4259 2578 4263 2582
rect 4275 2578 4279 2582
rect 4475 2578 4479 2582
rect 4555 2578 4559 2582
rect 4715 2578 4719 2582
rect 4867 2578 4871 2582
rect 4979 2578 4983 2582
rect 5203 2578 5207 2582
rect 5259 2578 5263 2582
rect 5515 2578 5519 2582
rect 5663 2578 5667 2582
rect 1975 2522 1979 2526
rect 1995 2522 1999 2526
rect 2235 2522 2239 2526
rect 2483 2522 2487 2526
rect 2715 2522 2719 2526
rect 2939 2522 2943 2526
rect 3107 2522 3111 2526
rect 3155 2522 3159 2526
rect 3243 2522 3247 2526
rect 3363 2522 3367 2526
rect 3379 2522 3383 2526
rect 3515 2522 3519 2526
rect 3579 2522 3583 2526
rect 3651 2522 3655 2526
rect 3799 2522 3803 2526
rect 3839 2462 3843 2466
rect 4287 2462 4291 2466
rect 4503 2462 4507 2466
rect 4663 2462 4667 2466
rect 4743 2462 4747 2466
rect 4847 2462 4851 2466
rect 5007 2462 5011 2466
rect 5023 2462 5027 2466
rect 5199 2462 5203 2466
rect 5287 2462 5291 2466
rect 5383 2462 5387 2466
rect 5543 2462 5547 2466
rect 5663 2462 5667 2466
rect 111 2422 115 2426
rect 203 2422 207 2426
rect 219 2422 223 2426
rect 395 2422 399 2426
rect 403 2422 407 2426
rect 595 2422 599 2426
rect 787 2422 791 2426
rect 795 2422 799 2426
rect 979 2422 983 2426
rect 995 2422 999 2426
rect 1195 2422 1199 2426
rect 1395 2422 1399 2426
rect 1603 2422 1607 2426
rect 1787 2422 1791 2426
rect 1935 2422 1939 2426
rect 1975 2410 1979 2414
rect 2023 2410 2027 2414
rect 2159 2410 2163 2414
rect 2263 2410 2267 2414
rect 2295 2410 2299 2414
rect 2431 2410 2435 2414
rect 2511 2410 2515 2414
rect 2567 2410 2571 2414
rect 2711 2410 2715 2414
rect 2743 2410 2747 2414
rect 2855 2410 2859 2414
rect 2967 2410 2971 2414
rect 3007 2410 3011 2414
rect 3159 2410 3163 2414
rect 3183 2410 3187 2414
rect 3311 2410 3315 2414
rect 3391 2410 3395 2414
rect 3607 2410 3611 2414
rect 3799 2410 3803 2414
rect 111 2306 115 2310
rect 247 2306 251 2310
rect 399 2306 403 2310
rect 431 2306 435 2310
rect 535 2306 539 2310
rect 623 2306 627 2310
rect 671 2306 675 2310
rect 807 2306 811 2310
rect 815 2306 819 2310
rect 943 2306 947 2310
rect 1007 2306 1011 2310
rect 1935 2306 1939 2310
rect 3839 2346 3843 2350
rect 4635 2346 4639 2350
rect 4675 2346 4679 2350
rect 4819 2346 4823 2350
rect 4963 2346 4967 2350
rect 4995 2346 4999 2350
rect 5115 2346 5119 2350
rect 5171 2346 5175 2350
rect 5267 2346 5271 2350
rect 5355 2346 5359 2350
rect 5419 2346 5423 2350
rect 5515 2346 5519 2350
rect 5663 2346 5667 2350
rect 1975 2294 1979 2298
rect 1995 2294 1999 2298
rect 2043 2294 2047 2298
rect 2131 2294 2135 2298
rect 2179 2294 2183 2298
rect 2267 2294 2271 2298
rect 2315 2294 2319 2298
rect 2403 2294 2407 2298
rect 2451 2294 2455 2298
rect 2539 2294 2543 2298
rect 2587 2294 2591 2298
rect 2683 2294 2687 2298
rect 2723 2294 2727 2298
rect 2827 2294 2831 2298
rect 2859 2294 2863 2298
rect 2979 2294 2983 2298
rect 2995 2294 2999 2298
rect 3131 2294 3135 2298
rect 3283 2294 3287 2298
rect 3799 2294 3803 2298
rect 3839 2222 3843 2226
rect 3887 2222 3891 2226
rect 4167 2222 4171 2226
rect 4455 2222 4459 2226
rect 4703 2222 4707 2226
rect 4719 2222 4723 2226
rect 4847 2222 4851 2226
rect 4975 2222 4979 2226
rect 4991 2222 4995 2226
rect 5143 2222 5147 2226
rect 5231 2222 5235 2226
rect 5295 2222 5299 2226
rect 5447 2222 5451 2226
rect 5487 2222 5491 2226
rect 5663 2222 5667 2226
rect 111 2186 115 2190
rect 323 2186 327 2190
rect 371 2186 375 2190
rect 459 2186 463 2190
rect 507 2186 511 2190
rect 595 2186 599 2190
rect 643 2186 647 2190
rect 731 2186 735 2190
rect 779 2186 783 2190
rect 867 2186 871 2190
rect 915 2186 919 2190
rect 1935 2186 1939 2190
rect 1975 2182 1979 2186
rect 2023 2182 2027 2186
rect 2071 2182 2075 2186
rect 2207 2182 2211 2186
rect 2239 2182 2243 2186
rect 2343 2182 2347 2186
rect 2479 2182 2483 2186
rect 2487 2182 2491 2186
rect 2615 2182 2619 2186
rect 2727 2182 2731 2186
rect 2751 2182 2755 2186
rect 2887 2182 2891 2186
rect 2967 2182 2971 2186
rect 3023 2182 3027 2186
rect 3159 2182 3163 2186
rect 3207 2182 3211 2186
rect 3455 2182 3459 2186
rect 3679 2182 3683 2186
rect 3799 2182 3803 2186
rect 3839 2110 3843 2114
rect 3859 2110 3863 2114
rect 4083 2110 4087 2114
rect 4139 2110 4143 2114
rect 4323 2110 4327 2114
rect 4427 2110 4431 2114
rect 4547 2110 4551 2114
rect 4691 2110 4695 2114
rect 4755 2110 4759 2114
rect 4947 2110 4951 2114
rect 5139 2110 5143 2114
rect 5203 2110 5207 2114
rect 5323 2110 5327 2114
rect 5459 2110 5463 2114
rect 5515 2110 5519 2114
rect 5663 2110 5667 2114
rect 1975 2054 1979 2058
rect 1995 2054 1999 2058
rect 2211 2054 2215 2058
rect 2459 2054 2463 2058
rect 2699 2054 2703 2058
rect 2707 2054 2711 2058
rect 2939 2054 2943 2058
rect 2963 2054 2967 2058
rect 3179 2054 3183 2058
rect 3219 2054 3223 2058
rect 3427 2054 3431 2058
rect 3483 2054 3487 2058
rect 3651 2054 3655 2058
rect 3799 2054 3803 2058
rect 111 2042 115 2046
rect 319 2042 323 2046
rect 351 2042 355 2046
rect 479 2042 483 2046
rect 487 2042 491 2046
rect 623 2042 627 2046
rect 663 2042 667 2046
rect 759 2042 763 2046
rect 871 2042 875 2046
rect 895 2042 899 2046
rect 1095 2042 1099 2046
rect 1335 2042 1339 2046
rect 1583 2042 1587 2046
rect 1815 2042 1819 2046
rect 1935 2042 1939 2046
rect 3839 1998 3843 2002
rect 3887 1998 3891 2002
rect 4111 1998 4115 2002
rect 4167 1998 4171 2002
rect 4351 1998 4355 2002
rect 4463 1998 4467 2002
rect 4575 1998 4579 2002
rect 4743 1998 4747 2002
rect 4783 1998 4787 2002
rect 4975 1998 4979 2002
rect 5007 1998 5011 2002
rect 5167 1998 5171 2002
rect 5271 1998 5275 2002
rect 5351 1998 5355 2002
rect 5543 1998 5547 2002
rect 5663 1998 5667 2002
rect 1975 1934 1979 1938
rect 2023 1934 2027 1938
rect 2159 1934 2163 1938
rect 2239 1934 2243 1938
rect 2439 1934 2443 1938
rect 2487 1934 2491 1938
rect 2703 1934 2707 1938
rect 2735 1934 2739 1938
rect 2959 1934 2963 1938
rect 2991 1934 2995 1938
rect 3207 1934 3211 1938
rect 3247 1934 3251 1938
rect 3455 1934 3459 1938
rect 3511 1934 3515 1938
rect 3679 1934 3683 1938
rect 3799 1934 3803 1938
rect 111 1922 115 1926
rect 187 1922 191 1926
rect 291 1922 295 1926
rect 419 1922 423 1926
rect 451 1922 455 1926
rect 635 1922 639 1926
rect 651 1922 655 1926
rect 843 1922 847 1926
rect 883 1922 887 1926
rect 1067 1922 1071 1926
rect 1115 1922 1119 1926
rect 1307 1922 1311 1926
rect 1347 1922 1351 1926
rect 1555 1922 1559 1926
rect 1579 1922 1583 1926
rect 1787 1922 1791 1926
rect 1935 1922 1939 1926
rect 3839 1874 3843 1878
rect 3859 1874 3863 1878
rect 4139 1874 4143 1878
rect 4435 1874 4439 1878
rect 4539 1874 4543 1878
rect 4715 1874 4719 1878
rect 4723 1874 4727 1878
rect 4915 1874 4919 1878
rect 4979 1874 4983 1878
rect 5115 1874 5119 1878
rect 5243 1874 5247 1878
rect 5323 1874 5327 1878
rect 5515 1874 5519 1878
rect 5663 1874 5667 1878
rect 1975 1814 1979 1818
rect 2131 1814 2135 1818
rect 2307 1814 2311 1818
rect 2411 1814 2415 1818
rect 2499 1814 2503 1818
rect 2675 1814 2679 1818
rect 2691 1814 2695 1818
rect 2883 1814 2887 1818
rect 2931 1814 2935 1818
rect 3067 1814 3071 1818
rect 3179 1814 3183 1818
rect 3251 1814 3255 1818
rect 3427 1814 3431 1818
rect 3443 1814 3447 1818
rect 3635 1814 3639 1818
rect 3651 1814 3655 1818
rect 3799 1814 3803 1818
rect 111 1798 115 1802
rect 159 1798 163 1802
rect 215 1798 219 1802
rect 367 1798 371 1802
rect 447 1798 451 1802
rect 591 1798 595 1802
rect 679 1798 683 1802
rect 799 1798 803 1802
rect 911 1798 915 1802
rect 999 1798 1003 1802
rect 1143 1798 1147 1802
rect 1191 1798 1195 1802
rect 1375 1798 1379 1802
rect 1559 1798 1563 1802
rect 1607 1798 1611 1802
rect 1751 1798 1755 1802
rect 1815 1798 1819 1802
rect 1935 1798 1939 1802
rect 3839 1754 3843 1758
rect 4383 1754 4387 1758
rect 4567 1754 4571 1758
rect 4599 1754 4603 1758
rect 4751 1754 4755 1758
rect 4831 1754 4835 1758
rect 4943 1754 4947 1758
rect 5071 1754 5075 1758
rect 5143 1754 5147 1758
rect 5319 1754 5323 1758
rect 5351 1754 5355 1758
rect 5543 1754 5547 1758
rect 5663 1754 5667 1758
rect 1975 1702 1979 1706
rect 2335 1702 2339 1706
rect 2471 1702 2475 1706
rect 2527 1702 2531 1706
rect 2607 1702 2611 1706
rect 2719 1702 2723 1706
rect 2743 1702 2747 1706
rect 2879 1702 2883 1706
rect 2911 1702 2915 1706
rect 3023 1702 3027 1706
rect 3095 1702 3099 1706
rect 3175 1702 3179 1706
rect 3279 1702 3283 1706
rect 3327 1702 3331 1706
rect 3471 1702 3475 1706
rect 3663 1702 3667 1706
rect 3799 1702 3803 1706
rect 111 1678 115 1682
rect 131 1678 135 1682
rect 339 1678 343 1682
rect 355 1678 359 1682
rect 563 1678 567 1682
rect 595 1678 599 1682
rect 771 1678 775 1682
rect 835 1678 839 1682
rect 971 1678 975 1682
rect 1067 1678 1071 1682
rect 1163 1678 1167 1682
rect 1307 1678 1311 1682
rect 1347 1678 1351 1682
rect 1531 1678 1535 1682
rect 1547 1678 1551 1682
rect 1723 1678 1727 1682
rect 1935 1678 1939 1682
rect 3839 1630 3843 1634
rect 3907 1630 3911 1634
rect 4123 1630 4127 1634
rect 4355 1630 4359 1634
rect 4363 1630 4367 1634
rect 4571 1630 4575 1634
rect 4627 1630 4631 1634
rect 4803 1630 4807 1634
rect 4907 1630 4911 1634
rect 5043 1630 5047 1634
rect 5195 1630 5199 1634
rect 5291 1630 5295 1634
rect 5491 1630 5495 1634
rect 5515 1630 5519 1634
rect 5663 1630 5667 1634
rect 1975 1590 1979 1594
rect 2355 1590 2359 1594
rect 2443 1590 2447 1594
rect 2563 1590 2567 1594
rect 2579 1590 2583 1594
rect 2715 1590 2719 1594
rect 2779 1590 2783 1594
rect 2851 1590 2855 1594
rect 2995 1590 2999 1594
rect 3003 1590 3007 1594
rect 3147 1590 3151 1594
rect 3227 1590 3231 1594
rect 3299 1590 3303 1594
rect 3459 1590 3463 1594
rect 3799 1590 3803 1594
rect 111 1562 115 1566
rect 159 1562 163 1566
rect 359 1562 363 1566
rect 383 1562 387 1566
rect 575 1562 579 1566
rect 623 1562 627 1566
rect 783 1562 787 1566
rect 863 1562 867 1566
rect 983 1562 987 1566
rect 1095 1562 1099 1566
rect 1183 1562 1187 1566
rect 1335 1562 1339 1566
rect 1375 1562 1379 1566
rect 1575 1562 1579 1566
rect 1935 1562 1939 1566
rect 3839 1518 3843 1522
rect 3887 1518 3891 1522
rect 3935 1518 3939 1522
rect 4023 1518 4027 1522
rect 4151 1518 4155 1522
rect 4159 1518 4163 1522
rect 4295 1518 4299 1522
rect 4391 1518 4395 1522
rect 4479 1518 4483 1522
rect 4655 1518 4659 1522
rect 4695 1518 4699 1522
rect 4935 1518 4939 1522
rect 5191 1518 5195 1522
rect 5223 1518 5227 1522
rect 5447 1518 5451 1522
rect 5519 1518 5523 1522
rect 5663 1518 5667 1522
rect 1975 1478 1979 1482
rect 2023 1478 2027 1482
rect 2159 1478 2163 1482
rect 2327 1478 2331 1482
rect 2383 1478 2387 1482
rect 2543 1478 2547 1482
rect 2591 1478 2595 1482
rect 2799 1478 2803 1482
rect 2807 1478 2811 1482
rect 3031 1478 3035 1482
rect 3087 1478 3091 1482
rect 3255 1478 3259 1482
rect 3391 1478 3395 1482
rect 3487 1478 3491 1482
rect 3679 1478 3683 1482
rect 3799 1478 3803 1482
rect 111 1430 115 1434
rect 131 1430 135 1434
rect 235 1430 239 1434
rect 331 1430 335 1434
rect 507 1430 511 1434
rect 547 1430 551 1434
rect 755 1430 759 1434
rect 779 1430 783 1434
rect 955 1430 959 1434
rect 1059 1430 1063 1434
rect 1155 1430 1159 1434
rect 1339 1430 1343 1434
rect 1347 1430 1351 1434
rect 1547 1430 1551 1434
rect 1935 1430 1939 1434
rect 3839 1394 3843 1398
rect 3859 1394 3863 1398
rect 3995 1394 3999 1398
rect 4131 1394 4135 1398
rect 4147 1394 4151 1398
rect 4267 1394 4271 1398
rect 4363 1394 4367 1398
rect 4451 1394 4455 1398
rect 4611 1394 4615 1398
rect 4667 1394 4671 1398
rect 4891 1394 4895 1398
rect 4907 1394 4911 1398
rect 5163 1394 5167 1398
rect 5195 1394 5199 1398
rect 5419 1394 5423 1398
rect 5499 1394 5503 1398
rect 5663 1394 5667 1398
rect 1975 1366 1979 1370
rect 1995 1366 1999 1370
rect 2131 1366 2135 1370
rect 2299 1366 2303 1370
rect 2491 1366 2495 1370
rect 2515 1366 2519 1370
rect 2771 1366 2775 1370
rect 3019 1366 3023 1370
rect 3059 1366 3063 1370
rect 3363 1366 3367 1370
rect 3555 1366 3559 1370
rect 3651 1366 3655 1370
rect 3799 1366 3803 1370
rect 111 1314 115 1318
rect 159 1314 163 1318
rect 263 1314 267 1318
rect 383 1314 387 1318
rect 535 1314 539 1318
rect 599 1314 603 1318
rect 799 1314 803 1318
rect 807 1314 811 1318
rect 991 1314 995 1318
rect 1087 1314 1091 1318
rect 1167 1314 1171 1318
rect 1335 1314 1339 1318
rect 1367 1314 1371 1318
rect 1503 1314 1507 1318
rect 1671 1314 1675 1318
rect 1815 1314 1819 1318
rect 1935 1314 1939 1318
rect 111 1194 115 1198
rect 131 1194 135 1198
rect 147 1194 151 1198
rect 323 1194 327 1198
rect 355 1194 359 1198
rect 499 1194 503 1198
rect 571 1194 575 1198
rect 675 1194 679 1198
rect 771 1194 775 1198
rect 851 1194 855 1198
rect 963 1194 967 1198
rect 1019 1194 1023 1198
rect 1139 1194 1143 1198
rect 1179 1194 1183 1198
rect 1307 1194 1311 1198
rect 1331 1194 1335 1198
rect 1475 1194 1479 1198
rect 1483 1194 1487 1198
rect 1643 1194 1647 1198
rect 1787 1194 1791 1198
rect 1935 1194 1939 1198
rect 3839 1282 3843 1286
rect 3887 1282 3891 1286
rect 4023 1282 4027 1286
rect 4167 1282 4171 1286
rect 4175 1282 4179 1286
rect 4335 1282 4339 1286
rect 4391 1282 4395 1286
rect 4511 1282 4515 1286
rect 4639 1282 4643 1286
rect 4703 1282 4707 1286
rect 4903 1282 4907 1286
rect 4919 1282 4923 1286
rect 5119 1282 5123 1286
rect 5223 1282 5227 1286
rect 5343 1282 5347 1286
rect 5527 1282 5531 1286
rect 5543 1282 5547 1286
rect 5663 1282 5667 1286
rect 1975 1190 1979 1194
rect 2023 1190 2027 1194
rect 2519 1190 2523 1194
rect 2743 1190 2747 1194
rect 3047 1190 3051 1194
rect 3359 1190 3363 1194
rect 3583 1190 3587 1194
rect 3679 1190 3683 1194
rect 3799 1190 3803 1194
rect 3839 1166 3843 1170
rect 3859 1166 3863 1170
rect 3995 1166 3999 1170
rect 4139 1166 4143 1170
rect 4307 1166 4311 1170
rect 4483 1166 4487 1170
rect 4675 1166 4679 1170
rect 4811 1166 4815 1170
rect 4875 1166 4879 1170
rect 4947 1166 4951 1170
rect 5083 1166 5087 1170
rect 5091 1166 5095 1170
rect 5227 1166 5231 1170
rect 5315 1166 5319 1170
rect 5379 1166 5383 1170
rect 5515 1166 5519 1170
rect 5663 1166 5667 1170
rect 1975 1078 1979 1082
rect 2243 1078 2247 1082
rect 2379 1078 2383 1082
rect 2523 1078 2527 1082
rect 2675 1078 2679 1082
rect 2715 1078 2719 1082
rect 2827 1078 2831 1082
rect 2987 1078 2991 1082
rect 3019 1078 3023 1082
rect 3155 1078 3159 1082
rect 3323 1078 3327 1082
rect 3331 1078 3335 1082
rect 3499 1078 3503 1082
rect 3651 1078 3655 1082
rect 3799 1078 3803 1082
rect 111 1062 115 1066
rect 159 1062 163 1066
rect 175 1062 179 1066
rect 351 1062 355 1066
rect 447 1062 451 1066
rect 527 1062 531 1066
rect 703 1062 707 1066
rect 775 1062 779 1066
rect 879 1062 883 1066
rect 1047 1062 1051 1066
rect 1111 1062 1115 1066
rect 1207 1062 1211 1066
rect 1359 1062 1363 1066
rect 1455 1062 1459 1066
rect 1511 1062 1515 1066
rect 1671 1062 1675 1066
rect 1807 1062 1811 1066
rect 1815 1062 1819 1066
rect 1935 1062 1939 1066
rect 3839 1050 3843 1054
rect 4807 1050 4811 1054
rect 4839 1050 4843 1054
rect 4943 1050 4947 1054
rect 4975 1050 4979 1054
rect 5079 1050 5083 1054
rect 5111 1050 5115 1054
rect 5215 1050 5219 1054
rect 5255 1050 5259 1054
rect 5351 1050 5355 1054
rect 5407 1050 5411 1054
rect 5487 1050 5491 1054
rect 5543 1050 5547 1054
rect 5663 1050 5667 1054
rect 1975 962 1979 966
rect 2271 962 2275 966
rect 2279 962 2283 966
rect 2407 962 2411 966
rect 2495 962 2499 966
rect 2551 962 2555 966
rect 2703 962 2707 966
rect 2711 962 2715 966
rect 2855 962 2859 966
rect 2911 962 2915 966
rect 3015 962 3019 966
rect 3103 962 3107 966
rect 3183 962 3187 966
rect 3295 962 3299 966
rect 3351 962 3355 966
rect 3479 962 3483 966
rect 3527 962 3531 966
rect 3671 962 3675 966
rect 3679 962 3683 966
rect 3799 962 3803 966
rect 111 946 115 950
rect 131 946 135 950
rect 339 946 343 950
rect 419 946 423 950
rect 595 946 599 950
rect 747 946 751 950
rect 875 946 879 950
rect 1083 946 1087 950
rect 1179 946 1183 950
rect 1427 946 1431 950
rect 1491 946 1495 950
rect 1779 946 1783 950
rect 1787 946 1791 950
rect 1935 946 1939 950
rect 3839 934 3843 938
rect 4355 934 4359 938
rect 4571 934 4575 938
rect 4779 934 4783 938
rect 4803 934 4807 938
rect 4915 934 4919 938
rect 5043 934 5047 938
rect 5051 934 5055 938
rect 5187 934 5191 938
rect 5291 934 5295 938
rect 5323 934 5327 938
rect 5459 934 5463 938
rect 5515 934 5519 938
rect 5663 934 5667 938
rect 1975 846 1979 850
rect 1995 846 1999 850
rect 2131 846 2135 850
rect 2251 846 2255 850
rect 2283 846 2287 850
rect 2443 846 2447 850
rect 2467 846 2471 850
rect 2603 846 2607 850
rect 2683 846 2687 850
rect 2763 846 2767 850
rect 2883 846 2887 850
rect 2923 846 2927 850
rect 3075 846 3079 850
rect 3083 846 3087 850
rect 3243 846 3247 850
rect 3267 846 3271 850
rect 3403 846 3407 850
rect 3451 846 3455 850
rect 3643 846 3647 850
rect 3799 846 3803 850
rect 111 822 115 826
rect 159 822 163 826
rect 367 822 371 826
rect 383 822 387 826
rect 623 822 627 826
rect 631 822 635 826
rect 887 822 891 826
rect 903 822 907 826
rect 1143 822 1147 826
rect 1207 822 1211 826
rect 1519 822 1523 826
rect 1815 822 1819 826
rect 1935 822 1939 826
rect 3839 818 3843 822
rect 3959 818 3963 822
rect 4207 818 4211 822
rect 4383 818 4387 822
rect 4495 818 4499 822
rect 4599 818 4603 822
rect 4815 818 4819 822
rect 4831 818 4835 822
rect 5071 818 5075 822
rect 5151 818 5155 822
rect 5319 818 5323 822
rect 5487 818 5491 822
rect 5543 818 5547 822
rect 5663 818 5667 822
rect 1975 734 1979 738
rect 2023 734 2027 738
rect 2159 734 2163 738
rect 2183 734 2187 738
rect 2311 734 2315 738
rect 2439 734 2443 738
rect 2471 734 2475 738
rect 2631 734 2635 738
rect 2679 734 2683 738
rect 2791 734 2795 738
rect 2903 734 2907 738
rect 2951 734 2955 738
rect 3111 734 3115 738
rect 3271 734 3275 738
rect 3311 734 3315 738
rect 3431 734 3435 738
rect 3503 734 3507 738
rect 3679 734 3683 738
rect 3799 734 3803 738
rect 111 710 115 714
rect 131 710 135 714
rect 355 710 359 714
rect 603 710 607 714
rect 699 710 703 714
rect 835 710 839 714
rect 859 710 863 714
rect 971 710 975 714
rect 1107 710 1111 714
rect 1115 710 1119 714
rect 1243 710 1247 714
rect 1379 710 1383 714
rect 1515 710 1519 714
rect 1651 710 1655 714
rect 1787 710 1791 714
rect 1935 710 1939 714
rect 3839 694 3843 698
rect 3859 694 3863 698
rect 3931 694 3935 698
rect 3995 694 3999 698
rect 4147 694 4151 698
rect 4179 694 4183 698
rect 4355 694 4359 698
rect 4467 694 4471 698
rect 4595 694 4599 698
rect 4787 694 4791 698
rect 4867 694 4871 698
rect 5123 694 5127 698
rect 5163 694 5167 698
rect 5459 694 5463 698
rect 5663 694 5667 698
rect 111 598 115 602
rect 159 598 163 602
rect 375 598 379 602
rect 599 598 603 602
rect 727 598 731 602
rect 807 598 811 602
rect 863 598 867 602
rect 999 598 1003 602
rect 1135 598 1139 602
rect 1175 598 1179 602
rect 1271 598 1275 602
rect 1343 598 1347 602
rect 1407 598 1411 602
rect 1511 598 1515 602
rect 1543 598 1547 602
rect 1671 598 1675 602
rect 1679 598 1683 602
rect 1815 598 1819 602
rect 1935 598 1939 602
rect 111 486 115 490
rect 131 486 135 490
rect 347 486 351 490
rect 355 486 359 490
rect 571 486 575 490
rect 603 486 607 490
rect 779 486 783 490
rect 843 486 847 490
rect 971 486 975 490
rect 1083 486 1087 490
rect 1147 486 1151 490
rect 1315 486 1319 490
rect 1323 486 1327 490
rect 1483 486 1487 490
rect 1563 486 1567 490
rect 1643 486 1647 490
rect 1787 486 1791 490
rect 1935 486 1939 490
rect 3839 582 3843 586
rect 3887 582 3891 586
rect 4023 582 4027 586
rect 4159 582 4163 586
rect 4175 582 4179 586
rect 4295 582 4299 586
rect 4383 582 4387 586
rect 4431 582 4435 586
rect 4567 582 4571 586
rect 4623 582 4627 586
rect 4711 582 4715 586
rect 4879 582 4883 586
rect 4895 582 4899 586
rect 5063 582 5067 586
rect 5191 582 5195 586
rect 5255 582 5259 586
rect 5447 582 5451 586
rect 5487 582 5491 586
rect 5663 582 5667 586
rect 3839 470 3843 474
rect 3859 470 3863 474
rect 3995 470 3999 474
rect 4115 470 4119 474
rect 4131 470 4135 474
rect 4267 470 4271 474
rect 4395 470 4399 474
rect 4403 470 4407 474
rect 4539 470 4543 474
rect 4675 470 4679 474
rect 4683 470 4687 474
rect 4851 470 4855 474
rect 4947 470 4951 474
rect 5035 470 5039 474
rect 5227 470 5231 474
rect 5419 470 5423 474
rect 5507 470 5511 474
rect 5663 470 5667 474
rect 1975 446 1979 450
rect 1995 446 1999 450
rect 2155 446 2159 450
rect 2251 446 2255 450
rect 2411 446 2415 450
rect 2523 446 2527 450
rect 2651 446 2655 450
rect 2771 446 2775 450
rect 2875 446 2879 450
rect 3003 446 3007 450
rect 3083 446 3087 450
rect 3227 446 3231 450
rect 3283 446 3287 450
rect 3451 446 3455 450
rect 3475 446 3479 450
rect 3651 446 3655 450
rect 3799 446 3803 450
rect 111 358 115 362
rect 159 358 163 362
rect 303 358 307 362
rect 383 358 387 362
rect 479 358 483 362
rect 631 358 635 362
rect 655 358 659 362
rect 831 358 835 362
rect 871 358 875 362
rect 1111 358 1115 362
rect 1351 358 1355 362
rect 1591 358 1595 362
rect 1815 358 1819 362
rect 1935 358 1939 362
rect 3839 350 3843 354
rect 3887 350 3891 354
rect 4143 350 4147 354
rect 4423 350 4427 354
rect 4703 350 4707 354
rect 4727 350 4731 354
rect 4895 350 4899 354
rect 4975 350 4979 354
rect 5063 350 5067 354
rect 5231 350 5235 354
rect 5255 350 5259 354
rect 5399 350 5403 354
rect 5535 350 5539 354
rect 5543 350 5547 354
rect 5663 350 5667 354
rect 1975 330 1979 334
rect 2023 330 2027 334
rect 2159 330 2163 334
rect 2279 330 2283 334
rect 2295 330 2299 334
rect 2431 330 2435 334
rect 2551 330 2555 334
rect 2567 330 2571 334
rect 2703 330 2707 334
rect 2799 330 2803 334
rect 2839 330 2843 334
rect 2975 330 2979 334
rect 3031 330 3035 334
rect 3111 330 3115 334
rect 3247 330 3251 334
rect 3255 330 3259 334
rect 3383 330 3387 334
rect 3479 330 3483 334
rect 3519 330 3523 334
rect 3655 330 3659 334
rect 3679 330 3683 334
rect 3799 330 3803 334
rect 111 206 115 210
rect 131 206 135 210
rect 267 206 271 210
rect 275 206 279 210
rect 403 206 407 210
rect 451 206 455 210
rect 539 206 543 210
rect 627 206 631 210
rect 675 206 679 210
rect 803 206 807 210
rect 811 206 815 210
rect 947 206 951 210
rect 1083 206 1087 210
rect 1935 206 1939 210
rect 3839 198 3843 202
rect 4291 198 4295 202
rect 4427 198 4431 202
rect 4563 198 4567 202
rect 4699 198 4703 202
rect 4835 198 4839 202
rect 4867 198 4871 202
rect 4971 198 4975 202
rect 5035 198 5039 202
rect 5107 198 5111 202
rect 5203 198 5207 202
rect 5243 198 5247 202
rect 5371 198 5375 202
rect 5379 198 5383 202
rect 5515 198 5519 202
rect 5663 198 5667 202
rect 1975 186 1979 190
rect 1995 186 1999 190
rect 2131 186 2135 190
rect 2267 186 2271 190
rect 2403 186 2407 190
rect 2539 186 2543 190
rect 2675 186 2679 190
rect 2811 186 2815 190
rect 2947 186 2951 190
rect 3083 186 3087 190
rect 3219 186 3223 190
rect 3355 186 3359 190
rect 3491 186 3495 190
rect 3627 186 3631 190
rect 3799 186 3803 190
rect 111 94 115 98
rect 159 94 163 98
rect 295 94 299 98
rect 431 94 435 98
rect 567 94 571 98
rect 703 94 707 98
rect 839 94 843 98
rect 975 94 979 98
rect 1111 94 1115 98
rect 1935 94 1939 98
rect 3839 86 3843 90
rect 4319 86 4323 90
rect 4455 86 4459 90
rect 4591 86 4595 90
rect 4727 86 4731 90
rect 4863 86 4867 90
rect 4999 86 5003 90
rect 5135 86 5139 90
rect 5271 86 5275 90
rect 5407 86 5411 90
rect 5543 86 5547 90
rect 5663 86 5667 90
rect 1975 74 1979 78
rect 2023 74 2027 78
rect 2159 74 2163 78
rect 2295 74 2299 78
rect 2431 74 2435 78
rect 2567 74 2571 78
rect 2703 74 2707 78
rect 2839 74 2843 78
rect 2975 74 2979 78
rect 3111 74 3115 78
rect 3247 74 3251 78
rect 3383 74 3387 78
rect 3519 74 3523 78
rect 3655 74 3659 78
rect 3799 74 3803 78
<< m4 >>
rect 1946 5753 1947 5759
rect 1953 5758 3811 5759
rect 1953 5754 1975 5758
rect 1979 5754 2375 5758
rect 2379 5754 2511 5758
rect 2515 5754 2655 5758
rect 2659 5754 2807 5758
rect 2811 5754 2959 5758
rect 2963 5754 3119 5758
rect 3123 5754 3799 5758
rect 3803 5754 3811 5758
rect 1953 5753 3811 5754
rect 3817 5753 3818 5759
rect 84 5713 85 5719
rect 91 5718 1947 5719
rect 91 5714 111 5718
rect 115 5714 159 5718
rect 163 5714 295 5718
rect 299 5714 431 5718
rect 435 5714 567 5718
rect 571 5714 703 5718
rect 707 5714 839 5718
rect 843 5714 975 5718
rect 979 5714 1935 5718
rect 1939 5714 1947 5718
rect 91 5713 1947 5714
rect 1953 5713 1954 5719
rect 3810 5677 3811 5683
rect 3817 5682 5695 5683
rect 3817 5678 3839 5682
rect 3843 5678 4335 5682
rect 4339 5678 4471 5682
rect 4475 5678 4607 5682
rect 4611 5678 4743 5682
rect 4747 5678 4879 5682
rect 4883 5678 5015 5682
rect 5019 5678 5663 5682
rect 5667 5678 5695 5682
rect 3817 5677 5695 5678
rect 5701 5677 5702 5683
rect 1958 5641 1959 5647
rect 1965 5646 3823 5647
rect 1965 5642 1975 5646
rect 1979 5642 1995 5646
rect 1999 5642 2203 5646
rect 2207 5642 2347 5646
rect 2351 5642 2427 5646
rect 2431 5642 2483 5646
rect 2487 5642 2627 5646
rect 2631 5642 2651 5646
rect 2655 5642 2779 5646
rect 2783 5642 2867 5646
rect 2871 5642 2931 5646
rect 2935 5642 3075 5646
rect 3079 5642 3091 5646
rect 3095 5642 3275 5646
rect 3279 5642 3475 5646
rect 3479 5642 3651 5646
rect 3655 5642 3799 5646
rect 3803 5642 3823 5646
rect 1965 5641 3823 5642
rect 3829 5641 3830 5647
rect 96 5573 97 5579
rect 103 5578 1959 5579
rect 103 5574 111 5578
rect 115 5574 131 5578
rect 135 5574 267 5578
rect 271 5574 403 5578
rect 407 5574 539 5578
rect 543 5574 619 5578
rect 623 5574 675 5578
rect 679 5574 755 5578
rect 759 5574 811 5578
rect 815 5574 899 5578
rect 903 5574 947 5578
rect 951 5574 1051 5578
rect 1055 5574 1203 5578
rect 1207 5574 1355 5578
rect 1359 5574 1507 5578
rect 1511 5574 1651 5578
rect 1655 5574 1787 5578
rect 1791 5574 1935 5578
rect 1939 5574 1959 5578
rect 103 5573 1959 5574
rect 1965 5573 1966 5579
rect 3822 5565 3823 5571
rect 3829 5570 5707 5571
rect 3829 5566 3839 5570
rect 3843 5566 4211 5570
rect 4215 5566 4307 5570
rect 4311 5566 4403 5570
rect 4407 5566 4443 5570
rect 4447 5566 4579 5570
rect 4583 5566 4595 5570
rect 4599 5566 4715 5570
rect 4719 5566 4795 5570
rect 4799 5566 4851 5570
rect 4855 5566 4987 5570
rect 4991 5566 4995 5570
rect 4999 5566 5195 5570
rect 5199 5566 5663 5570
rect 5667 5566 5707 5570
rect 3829 5565 5707 5566
rect 5713 5565 5714 5571
rect 1946 5529 1947 5535
rect 1953 5534 3811 5535
rect 1953 5530 1975 5534
rect 1979 5530 2023 5534
rect 2027 5530 2231 5534
rect 2235 5530 2455 5534
rect 2459 5530 2679 5534
rect 2683 5530 2895 5534
rect 2899 5530 2951 5534
rect 2955 5530 3103 5534
rect 3107 5530 3255 5534
rect 3259 5530 3303 5534
rect 3307 5530 3415 5534
rect 3419 5530 3503 5534
rect 3507 5530 3679 5534
rect 3683 5530 3799 5534
rect 3803 5530 3811 5534
rect 1953 5529 3811 5530
rect 3817 5529 3818 5535
rect 84 5453 85 5459
rect 91 5458 1947 5459
rect 91 5454 111 5458
rect 115 5454 591 5458
rect 595 5454 647 5458
rect 651 5454 727 5458
rect 731 5454 783 5458
rect 787 5454 863 5458
rect 867 5454 927 5458
rect 931 5454 999 5458
rect 1003 5454 1079 5458
rect 1083 5454 1135 5458
rect 1139 5454 1231 5458
rect 1235 5454 1271 5458
rect 1275 5454 1383 5458
rect 1387 5454 1407 5458
rect 1411 5454 1535 5458
rect 1539 5454 1543 5458
rect 1547 5454 1679 5458
rect 1683 5454 1815 5458
rect 1819 5454 1935 5458
rect 1939 5454 1947 5458
rect 91 5453 1947 5454
rect 1953 5453 1954 5459
rect 3810 5417 3811 5423
rect 3817 5422 5695 5423
rect 3817 5418 3839 5422
rect 3843 5418 4239 5422
rect 4243 5418 4303 5422
rect 4307 5418 4431 5422
rect 4435 5418 4519 5422
rect 4523 5418 4623 5422
rect 4627 5418 4735 5422
rect 4739 5418 4823 5422
rect 4827 5418 4951 5422
rect 4955 5418 5023 5422
rect 5027 5418 5175 5422
rect 5179 5418 5223 5422
rect 5227 5418 5399 5422
rect 5403 5418 5663 5422
rect 5667 5418 5695 5422
rect 3817 5417 5695 5418
rect 5701 5417 5702 5423
rect 1958 5369 1959 5375
rect 1965 5374 3823 5375
rect 1965 5370 1975 5374
rect 1979 5370 2643 5374
rect 2647 5370 2811 5374
rect 2815 5370 2923 5374
rect 2927 5370 2979 5374
rect 2983 5370 3075 5374
rect 3079 5370 3139 5374
rect 3143 5370 3227 5374
rect 3231 5370 3307 5374
rect 3311 5370 3387 5374
rect 3391 5370 3475 5374
rect 3479 5370 3643 5374
rect 3647 5370 3799 5374
rect 3803 5370 3823 5374
rect 1965 5369 3823 5370
rect 3829 5369 3830 5375
rect 96 5317 97 5323
rect 103 5322 1959 5323
rect 103 5318 111 5322
rect 115 5318 411 5322
rect 415 5318 563 5322
rect 567 5318 587 5322
rect 591 5318 699 5322
rect 703 5318 763 5322
rect 767 5318 835 5322
rect 839 5318 939 5322
rect 943 5318 971 5322
rect 975 5318 1107 5322
rect 1111 5318 1243 5322
rect 1247 5318 1275 5322
rect 1279 5318 1379 5322
rect 1383 5318 1443 5322
rect 1447 5318 1515 5322
rect 1519 5318 1611 5322
rect 1615 5318 1651 5322
rect 1655 5318 1787 5322
rect 1791 5318 1935 5322
rect 1939 5318 1959 5322
rect 103 5317 1959 5318
rect 1965 5317 1966 5323
rect 3822 5273 3823 5279
rect 3829 5278 5707 5279
rect 3829 5274 3839 5278
rect 3843 5274 4275 5278
rect 4279 5274 4371 5278
rect 4375 5274 4491 5278
rect 4495 5274 4563 5278
rect 4567 5274 4707 5278
rect 4711 5274 4771 5278
rect 4775 5274 4923 5278
rect 4927 5274 4979 5278
rect 4983 5274 5147 5278
rect 5151 5274 5195 5278
rect 5199 5274 5371 5278
rect 5375 5274 5419 5278
rect 5423 5274 5663 5278
rect 5667 5274 5707 5278
rect 3829 5273 5707 5274
rect 5713 5273 5714 5279
rect 1946 5257 1947 5263
rect 1953 5262 3811 5263
rect 1953 5258 1975 5262
rect 1979 5258 2511 5262
rect 2515 5258 2671 5262
rect 2675 5258 2687 5262
rect 2691 5258 2839 5262
rect 2843 5258 2863 5262
rect 2867 5258 3007 5262
rect 3011 5258 3039 5262
rect 3043 5258 3167 5262
rect 3171 5258 3207 5262
rect 3211 5258 3335 5262
rect 3339 5258 3367 5262
rect 3371 5258 3503 5262
rect 3507 5258 3535 5262
rect 3539 5258 3671 5262
rect 3675 5258 3679 5262
rect 3683 5258 3799 5262
rect 3803 5258 3811 5262
rect 1953 5257 3811 5258
rect 3817 5257 3818 5263
rect 84 5197 85 5203
rect 91 5202 1947 5203
rect 91 5198 111 5202
rect 115 5198 207 5202
rect 211 5198 343 5202
rect 347 5198 439 5202
rect 443 5198 479 5202
rect 483 5198 615 5202
rect 619 5198 751 5202
rect 755 5198 791 5202
rect 795 5198 887 5202
rect 891 5198 967 5202
rect 971 5198 1023 5202
rect 1027 5198 1135 5202
rect 1139 5198 1303 5202
rect 1307 5198 1471 5202
rect 1475 5198 1639 5202
rect 1643 5198 1815 5202
rect 1819 5198 1935 5202
rect 1939 5198 1947 5202
rect 91 5197 1947 5198
rect 1953 5197 1954 5203
rect 3810 5147 3811 5153
rect 3817 5147 3842 5153
rect 3836 5143 3842 5147
rect 1958 5137 1959 5143
rect 1965 5142 3823 5143
rect 1965 5138 1975 5142
rect 1979 5138 2139 5142
rect 2143 5138 2307 5142
rect 2311 5138 2483 5142
rect 2487 5138 2491 5142
rect 2495 5138 2659 5142
rect 2663 5138 2691 5142
rect 2695 5138 2835 5142
rect 2839 5138 2915 5142
rect 2919 5138 3011 5142
rect 3015 5138 3163 5142
rect 3167 5138 3179 5142
rect 3183 5138 3339 5142
rect 3343 5138 3419 5142
rect 3423 5138 3507 5142
rect 3511 5138 3651 5142
rect 3655 5138 3799 5142
rect 3803 5138 3823 5142
rect 1965 5137 3823 5138
rect 3829 5137 3830 5143
rect 3836 5142 5695 5143
rect 3836 5138 3839 5142
rect 3843 5138 3887 5142
rect 3891 5138 4087 5142
rect 4091 5138 4311 5142
rect 4315 5138 4399 5142
rect 4403 5138 4535 5142
rect 4539 5138 4591 5142
rect 4595 5138 4759 5142
rect 4763 5138 4799 5142
rect 4803 5138 4983 5142
rect 4987 5138 5007 5142
rect 5011 5138 5207 5142
rect 5211 5138 5223 5142
rect 5227 5138 5439 5142
rect 5443 5138 5447 5142
rect 5451 5138 5663 5142
rect 5667 5138 5695 5142
rect 3836 5137 5695 5138
rect 5701 5137 5702 5143
rect 96 5065 97 5071
rect 103 5070 1959 5071
rect 103 5066 111 5070
rect 115 5066 147 5070
rect 151 5066 179 5070
rect 183 5066 315 5070
rect 319 5066 339 5070
rect 343 5066 451 5070
rect 455 5066 531 5070
rect 535 5066 587 5070
rect 591 5066 723 5070
rect 727 5066 731 5070
rect 735 5066 859 5070
rect 863 5066 931 5070
rect 935 5066 995 5070
rect 999 5066 1131 5070
rect 1135 5066 1935 5070
rect 1939 5066 1959 5070
rect 103 5065 1959 5066
rect 1965 5065 1966 5071
rect 3822 5009 3823 5015
rect 3829 5014 5707 5015
rect 3829 5010 3839 5014
rect 3843 5010 3859 5014
rect 3863 5010 3995 5014
rect 3999 5010 4059 5014
rect 4063 5010 4131 5014
rect 4135 5010 4283 5014
rect 4287 5010 4443 5014
rect 4447 5010 4507 5014
rect 4511 5010 4611 5014
rect 4615 5010 4731 5014
rect 4735 5010 4787 5014
rect 4791 5010 4955 5014
rect 4959 5010 4971 5014
rect 4975 5010 5155 5014
rect 5159 5010 5179 5014
rect 5183 5010 5339 5014
rect 5343 5010 5411 5014
rect 5415 5010 5515 5014
rect 5519 5010 5663 5014
rect 5667 5010 5707 5014
rect 3829 5009 5707 5010
rect 5713 5009 5714 5015
rect 1946 5001 1947 5007
rect 1953 5006 3811 5007
rect 1953 5002 1975 5006
rect 1979 5002 2023 5006
rect 2027 5002 2167 5006
rect 2171 5002 2335 5006
rect 2339 5002 2351 5006
rect 2355 5002 2519 5006
rect 2523 5002 2543 5006
rect 2547 5002 2719 5006
rect 2723 5002 2751 5006
rect 2755 5002 2943 5006
rect 2947 5002 2967 5006
rect 2971 5002 3183 5006
rect 3187 5002 3191 5006
rect 3195 5002 3447 5006
rect 3451 5002 3679 5006
rect 3683 5002 3799 5006
rect 3803 5002 3811 5006
rect 1953 5001 3811 5002
rect 3817 5001 3818 5007
rect 84 4941 85 4947
rect 91 4946 1947 4947
rect 91 4942 111 4946
rect 115 4942 159 4946
rect 163 4942 175 4946
rect 179 4942 367 4946
rect 371 4942 391 4946
rect 395 4942 559 4946
rect 563 4942 647 4946
rect 651 4942 759 4946
rect 763 4942 895 4946
rect 899 4942 959 4946
rect 963 4942 1135 4946
rect 1139 4942 1159 4946
rect 1163 4942 1367 4946
rect 1371 4942 1599 4946
rect 1603 4942 1815 4946
rect 1819 4942 1935 4946
rect 1939 4942 1947 4946
rect 91 4941 1947 4942
rect 1953 4941 1954 4947
rect 3810 4891 3811 4897
rect 3817 4891 3842 4897
rect 3836 4887 3842 4891
rect 1958 4881 1959 4887
rect 1965 4886 3823 4887
rect 1965 4882 1975 4886
rect 1979 4882 1995 4886
rect 1999 4882 2139 4886
rect 2143 4882 2323 4886
rect 2327 4882 2515 4886
rect 2519 4882 2667 4886
rect 2671 4882 2723 4886
rect 2727 4882 2939 4886
rect 2943 4882 3019 4886
rect 3023 4882 3155 4886
rect 3159 4882 3371 4886
rect 3375 4882 3799 4886
rect 3803 4882 3823 4886
rect 1965 4881 3823 4882
rect 3829 4881 3830 4887
rect 3836 4886 5695 4887
rect 3836 4882 3839 4886
rect 3843 4882 3887 4886
rect 3891 4882 3943 4886
rect 3947 4882 4023 4886
rect 4027 4882 4159 4886
rect 4163 4882 4183 4886
rect 4187 4882 4311 4886
rect 4315 4882 4431 4886
rect 4435 4882 4471 4886
rect 4475 4882 4639 4886
rect 4643 4882 4687 4886
rect 4691 4882 4815 4886
rect 4819 4882 4959 4886
rect 4963 4882 4999 4886
rect 5003 4882 5183 4886
rect 5187 4882 5239 4886
rect 5243 4882 5367 4886
rect 5371 4882 5519 4886
rect 5523 4882 5543 4886
rect 5547 4882 5663 4886
rect 5667 4882 5695 4886
rect 3836 4881 5695 4882
rect 5701 4881 5702 4887
rect 96 4829 97 4835
rect 103 4834 1959 4835
rect 103 4830 111 4834
rect 115 4830 131 4834
rect 135 4830 363 4834
rect 367 4830 475 4834
rect 479 4830 619 4834
rect 623 4830 859 4834
rect 863 4830 867 4834
rect 871 4830 1107 4834
rect 1111 4830 1251 4834
rect 1255 4830 1339 4834
rect 1343 4830 1571 4834
rect 1575 4830 1643 4834
rect 1647 4830 1787 4834
rect 1791 4830 1935 4834
rect 1939 4830 1959 4834
rect 103 4829 1959 4830
rect 1965 4829 1966 4835
rect 3822 4761 3823 4767
rect 3829 4766 5707 4767
rect 3829 4762 3839 4766
rect 3843 4762 3915 4766
rect 3919 4762 3939 4766
rect 3943 4762 4155 4766
rect 4159 4762 4179 4766
rect 4183 4762 4403 4766
rect 4407 4762 4435 4766
rect 4439 4762 4659 4766
rect 4663 4762 4691 4766
rect 4695 4762 4931 4766
rect 4935 4762 4955 4766
rect 4959 4762 5211 4766
rect 5215 4762 5227 4766
rect 5231 4762 5491 4766
rect 5495 4762 5507 4766
rect 5511 4762 5663 4766
rect 5667 4762 5707 4766
rect 3829 4761 5707 4762
rect 5713 4761 5714 4767
rect 1946 4721 1947 4727
rect 1953 4726 3811 4727
rect 1953 4722 1975 4726
rect 1979 4722 2023 4726
rect 2027 4722 2079 4726
rect 2083 4722 2231 4726
rect 2235 4722 2351 4726
rect 2355 4722 2391 4726
rect 2395 4722 2559 4726
rect 2563 4722 2695 4726
rect 2699 4722 2727 4726
rect 2731 4722 2903 4726
rect 2907 4722 3047 4726
rect 3051 4722 3079 4726
rect 3083 4722 3255 4726
rect 3259 4722 3399 4726
rect 3403 4722 3439 4726
rect 3443 4722 3623 4726
rect 3627 4722 3799 4726
rect 3803 4722 3811 4726
rect 1953 4721 3811 4722
rect 3817 4721 3818 4727
rect 84 4697 85 4703
rect 91 4702 1947 4703
rect 91 4698 111 4702
rect 115 4698 159 4702
rect 163 4698 295 4702
rect 299 4698 431 4702
rect 435 4698 503 4702
rect 507 4698 567 4702
rect 571 4698 703 4702
rect 707 4698 887 4702
rect 891 4698 1279 4702
rect 1283 4698 1671 4702
rect 1675 4698 1935 4702
rect 1939 4698 1947 4702
rect 91 4697 1947 4698
rect 1953 4697 1954 4703
rect 3810 4645 3811 4651
rect 3817 4650 5695 4651
rect 3817 4646 3839 4650
rect 3843 4646 3967 4650
rect 3971 4646 4175 4650
rect 4179 4646 4207 4650
rect 4211 4646 4455 4650
rect 4459 4646 4463 4650
rect 4467 4646 4719 4650
rect 4723 4646 4735 4650
rect 4739 4646 4983 4650
rect 4987 4646 5015 4650
rect 5019 4646 5255 4650
rect 5259 4646 5303 4650
rect 5307 4646 5535 4650
rect 5539 4646 5663 4650
rect 5667 4646 5695 4650
rect 3817 4645 5695 4646
rect 5701 4645 5702 4651
rect 1958 4605 1959 4611
rect 1965 4610 3823 4611
rect 1965 4606 1975 4610
rect 1979 4606 2051 4610
rect 2055 4606 2123 4610
rect 2127 4606 2203 4610
rect 2207 4606 2275 4610
rect 2279 4606 2363 4610
rect 2367 4606 2443 4610
rect 2447 4606 2531 4610
rect 2535 4606 2611 4610
rect 2615 4606 2699 4610
rect 2703 4606 2787 4610
rect 2791 4606 2875 4610
rect 2879 4606 2963 4610
rect 2967 4606 3051 4610
rect 3055 4606 3139 4610
rect 3143 4606 3227 4610
rect 3231 4606 3315 4610
rect 3319 4606 3411 4610
rect 3415 4606 3491 4610
rect 3495 4606 3595 4610
rect 3599 4606 3651 4610
rect 3655 4606 3799 4610
rect 3803 4606 3823 4610
rect 1965 4605 3823 4606
rect 3829 4605 3830 4611
rect 96 4569 97 4575
rect 103 4574 1959 4575
rect 103 4570 111 4574
rect 115 4570 131 4574
rect 135 4570 267 4574
rect 271 4570 291 4574
rect 295 4570 403 4574
rect 407 4570 427 4574
rect 431 4570 539 4574
rect 543 4570 563 4574
rect 567 4570 675 4574
rect 679 4570 699 4574
rect 703 4570 835 4574
rect 839 4570 1935 4574
rect 1939 4570 1959 4574
rect 103 4569 1959 4570
rect 1965 4569 1966 4575
rect 3822 4529 3823 4535
rect 3829 4534 5707 4535
rect 3829 4530 3839 4534
rect 3843 4530 3859 4534
rect 3863 4530 4147 4534
rect 4151 4530 4155 4534
rect 4159 4530 4427 4534
rect 4431 4530 4483 4534
rect 4487 4530 4707 4534
rect 4711 4530 4819 4534
rect 4823 4530 4987 4534
rect 4991 4530 5163 4534
rect 5167 4530 5275 4534
rect 5279 4530 5515 4534
rect 5519 4530 5663 4534
rect 5667 4530 5707 4534
rect 3829 4529 5707 4530
rect 5713 4529 5714 4535
rect 1946 4485 1947 4491
rect 1953 4490 3811 4491
rect 1953 4486 1975 4490
rect 1979 4486 2023 4490
rect 2027 4486 2151 4490
rect 2155 4486 2159 4490
rect 2163 4486 2295 4490
rect 2299 4486 2303 4490
rect 2307 4486 2431 4490
rect 2435 4486 2471 4490
rect 2475 4486 2567 4490
rect 2571 4486 2639 4490
rect 2643 4486 2703 4490
rect 2707 4486 2815 4490
rect 2819 4486 2839 4490
rect 2843 4486 2975 4490
rect 2979 4486 2991 4490
rect 2995 4486 3167 4490
rect 3171 4486 3343 4490
rect 3347 4486 3519 4490
rect 3523 4486 3679 4490
rect 3683 4486 3799 4490
rect 3803 4486 3811 4490
rect 1953 4485 3811 4486
rect 3817 4485 3818 4491
rect 84 4441 85 4447
rect 91 4446 1947 4447
rect 91 4442 111 4446
rect 115 4442 319 4446
rect 323 4442 455 4446
rect 459 4442 519 4446
rect 523 4442 591 4446
rect 595 4442 727 4446
rect 731 4442 743 4446
rect 747 4442 863 4446
rect 867 4442 991 4446
rect 995 4442 1263 4446
rect 1267 4442 1551 4446
rect 1555 4442 1815 4446
rect 1819 4442 1935 4446
rect 1939 4442 1947 4446
rect 91 4441 1947 4442
rect 1953 4441 1954 4447
rect 3810 4417 3811 4423
rect 3817 4422 5695 4423
rect 3817 4418 3839 4422
rect 3843 4418 3887 4422
rect 3891 4418 4143 4422
rect 4147 4418 4183 4422
rect 4187 4418 4423 4422
rect 4427 4418 4511 4422
rect 4515 4418 4703 4422
rect 4707 4418 4847 4422
rect 4851 4418 4983 4422
rect 4987 4418 5191 4422
rect 5195 4418 5263 4422
rect 5267 4418 5543 4422
rect 5547 4418 5663 4422
rect 5667 4418 5695 4422
rect 3817 4417 5695 4418
rect 5701 4417 5702 4423
rect 1958 4357 1959 4363
rect 1965 4362 3823 4363
rect 1965 4358 1975 4362
rect 1979 4358 1995 4362
rect 1999 4358 2131 4362
rect 2135 4358 2267 4362
rect 2271 4358 2403 4362
rect 2407 4358 2539 4362
rect 2543 4358 2675 4362
rect 2679 4358 2779 4362
rect 2783 4358 2811 4362
rect 2815 4358 2947 4362
rect 2951 4358 2995 4362
rect 2999 4358 3219 4362
rect 3223 4358 3443 4362
rect 3447 4358 3651 4362
rect 3655 4358 3799 4362
rect 3803 4358 3823 4362
rect 1965 4357 3823 4358
rect 3829 4357 3830 4363
rect 96 4329 97 4335
rect 103 4334 1959 4335
rect 103 4330 111 4334
rect 115 4330 491 4334
rect 495 4330 563 4334
rect 567 4330 699 4334
rect 703 4330 715 4334
rect 719 4330 835 4334
rect 839 4330 963 4334
rect 967 4330 971 4334
rect 975 4330 1107 4334
rect 1111 4330 1235 4334
rect 1239 4330 1243 4334
rect 1247 4330 1379 4334
rect 1383 4330 1515 4334
rect 1519 4330 1523 4334
rect 1527 4330 1651 4334
rect 1655 4330 1787 4334
rect 1791 4330 1935 4334
rect 1939 4330 1959 4334
rect 103 4329 1959 4330
rect 1965 4329 1966 4335
rect 3822 4293 3823 4299
rect 3829 4298 5707 4299
rect 3829 4294 3839 4298
rect 3843 4294 3859 4298
rect 3863 4294 4115 4298
rect 4119 4294 4395 4298
rect 4399 4294 4571 4298
rect 4575 4294 4675 4298
rect 4679 4294 4739 4298
rect 4743 4294 4915 4298
rect 4919 4294 4955 4298
rect 4959 4294 5107 4298
rect 5111 4294 5235 4298
rect 5239 4294 5307 4298
rect 5311 4294 5515 4298
rect 5519 4294 5663 4298
rect 5667 4294 5707 4298
rect 3829 4293 5707 4294
rect 5713 4293 5714 4299
rect 1946 4217 1947 4223
rect 1953 4222 3811 4223
rect 1953 4218 1975 4222
rect 1979 4218 2807 4222
rect 2811 4218 2951 4222
rect 2955 4218 3023 4222
rect 3027 4218 3095 4222
rect 3099 4218 3239 4222
rect 3243 4218 3247 4222
rect 3251 4218 3391 4222
rect 3395 4218 3471 4222
rect 3475 4218 3543 4222
rect 3547 4218 3679 4222
rect 3683 4218 3799 4222
rect 3803 4218 3811 4222
rect 1953 4217 3811 4218
rect 3817 4217 3818 4223
rect 84 4205 85 4211
rect 91 4210 1947 4211
rect 91 4206 111 4210
rect 115 4206 591 4210
rect 595 4206 727 4210
rect 731 4206 863 4210
rect 867 4206 999 4210
rect 1003 4206 1135 4210
rect 1139 4206 1271 4210
rect 1275 4206 1407 4210
rect 1411 4206 1543 4210
rect 1547 4206 1679 4210
rect 1683 4206 1815 4210
rect 1819 4206 1935 4210
rect 1939 4206 1947 4210
rect 91 4205 1947 4206
rect 1953 4205 1954 4211
rect 3810 4181 3811 4187
rect 3817 4186 5695 4187
rect 3817 4182 3839 4186
rect 3843 4182 4599 4186
rect 4603 4182 4655 4186
rect 4659 4182 4767 4186
rect 4771 4182 4815 4186
rect 4819 4182 4943 4186
rect 4947 4182 4983 4186
rect 4987 4182 5135 4186
rect 5139 4182 5167 4186
rect 5171 4182 5335 4186
rect 5339 4182 5359 4186
rect 5363 4182 5543 4186
rect 5547 4182 5663 4186
rect 5667 4182 5695 4186
rect 3817 4181 5695 4182
rect 5701 4181 5702 4187
rect 96 4093 97 4099
rect 103 4098 1959 4099
rect 103 4094 111 4098
rect 115 4094 563 4098
rect 567 4094 699 4098
rect 703 4094 835 4098
rect 839 4094 971 4098
rect 975 4094 1107 4098
rect 1111 4094 1243 4098
rect 1247 4094 1379 4098
rect 1383 4094 1515 4098
rect 1519 4094 1651 4098
rect 1655 4094 1787 4098
rect 1791 4094 1935 4098
rect 1939 4094 1959 4098
rect 103 4093 1959 4094
rect 1965 4093 1966 4099
rect 1958 4069 1959 4075
rect 1965 4074 3823 4075
rect 1965 4070 1975 4074
rect 1979 4070 2899 4074
rect 2903 4070 2923 4074
rect 2927 4070 3043 4074
rect 3047 4070 3067 4074
rect 3071 4070 3187 4074
rect 3191 4070 3211 4074
rect 3215 4070 3339 4074
rect 3343 4070 3363 4074
rect 3367 4070 3491 4074
rect 3495 4070 3515 4074
rect 3519 4070 3643 4074
rect 3647 4070 3651 4074
rect 3655 4070 3799 4074
rect 3803 4070 3823 4074
rect 1965 4069 3823 4070
rect 3829 4069 3830 4075
rect 3822 4033 3823 4039
rect 3829 4038 5707 4039
rect 3829 4034 3839 4038
rect 3843 4034 4627 4038
rect 4631 4034 4787 4038
rect 4791 4034 4939 4038
rect 4943 4034 4955 4038
rect 4959 4034 5075 4038
rect 5079 4034 5139 4038
rect 5143 4034 5211 4038
rect 5215 4034 5331 4038
rect 5335 4034 5347 4038
rect 5351 4034 5515 4038
rect 5519 4034 5663 4038
rect 5667 4034 5707 4038
rect 3829 4033 5707 4034
rect 5713 4033 5714 4039
rect 84 3977 85 3983
rect 91 3982 1947 3983
rect 91 3978 111 3982
rect 115 3978 695 3982
rect 699 3978 727 3982
rect 731 3978 831 3982
rect 835 3978 863 3982
rect 867 3978 967 3982
rect 971 3978 999 3982
rect 1003 3978 1111 3982
rect 1115 3978 1135 3982
rect 1139 3978 1255 3982
rect 1259 3978 1271 3982
rect 1275 3978 1399 3982
rect 1403 3978 1407 3982
rect 1411 3978 1543 3982
rect 1547 3978 1679 3982
rect 1683 3978 1815 3982
rect 1819 3978 1935 3982
rect 1939 3978 1947 3982
rect 91 3977 1947 3978
rect 1953 3977 1954 3983
rect 1946 3929 1947 3935
rect 1953 3934 3811 3935
rect 1953 3930 1975 3934
rect 1979 3930 2759 3934
rect 2763 3930 2911 3934
rect 2915 3930 2927 3934
rect 2931 3930 3071 3934
rect 3075 3930 3215 3934
rect 3219 3930 3239 3934
rect 3243 3930 3367 3934
rect 3371 3930 3415 3934
rect 3419 3930 3519 3934
rect 3523 3930 3591 3934
rect 3595 3930 3671 3934
rect 3675 3930 3799 3934
rect 3803 3930 3811 3934
rect 1953 3929 3811 3930
rect 3817 3929 3818 3935
rect 3810 3927 3818 3929
rect 3810 3921 3811 3927
rect 3817 3926 5695 3927
rect 3817 3922 3839 3926
rect 3843 3922 4687 3926
rect 4691 3922 4847 3926
rect 4851 3922 4967 3926
rect 4971 3922 5015 3926
rect 5019 3922 5103 3926
rect 5107 3922 5191 3926
rect 5195 3922 5239 3926
rect 5243 3922 5375 3926
rect 5379 3922 5543 3926
rect 5547 3922 5663 3926
rect 5667 3922 5695 3926
rect 3817 3921 5695 3922
rect 5701 3921 5702 3927
rect 96 3861 97 3867
rect 103 3866 1959 3867
rect 103 3862 111 3866
rect 115 3862 435 3866
rect 439 3862 619 3866
rect 623 3862 667 3866
rect 671 3862 803 3866
rect 807 3862 819 3866
rect 823 3862 939 3866
rect 943 3862 1027 3866
rect 1031 3862 1083 3866
rect 1087 3862 1227 3866
rect 1231 3862 1251 3866
rect 1255 3862 1371 3866
rect 1375 3862 1483 3866
rect 1487 3862 1515 3866
rect 1519 3862 1651 3866
rect 1655 3862 1723 3866
rect 1727 3862 1787 3866
rect 1791 3862 1935 3866
rect 1939 3862 1959 3866
rect 103 3861 1959 3862
rect 1965 3861 1966 3867
rect 1958 3809 1959 3815
rect 1965 3814 3823 3815
rect 1965 3810 1975 3814
rect 1979 3810 2115 3814
rect 2119 3810 2251 3814
rect 2255 3810 2387 3814
rect 2391 3810 2523 3814
rect 2527 3810 2659 3814
rect 2663 3810 2731 3814
rect 2735 3810 2795 3814
rect 2799 3810 2883 3814
rect 2887 3810 2939 3814
rect 2943 3810 3043 3814
rect 3047 3810 3083 3814
rect 3087 3810 3211 3814
rect 3215 3810 3235 3814
rect 3239 3810 3387 3814
rect 3391 3810 3395 3814
rect 3399 3810 3555 3814
rect 3559 3810 3563 3814
rect 3567 3810 3799 3814
rect 3803 3810 3823 3814
rect 1965 3809 3823 3810
rect 3829 3814 5714 3815
rect 3829 3810 3839 3814
rect 3843 3810 4411 3814
rect 4415 3810 4619 3814
rect 4623 3810 4659 3814
rect 4663 3810 4819 3814
rect 4823 3810 4835 3814
rect 4839 3810 4987 3814
rect 4991 3810 5067 3814
rect 5071 3810 5163 3814
rect 5167 3810 5299 3814
rect 5303 3810 5347 3814
rect 5351 3810 5515 3814
rect 5519 3810 5663 3814
rect 5667 3810 5714 3814
rect 3829 3809 5714 3810
rect 84 3745 85 3751
rect 91 3750 1947 3751
rect 91 3746 111 3750
rect 115 3746 231 3750
rect 235 3746 431 3750
rect 435 3746 463 3750
rect 467 3746 647 3750
rect 651 3746 655 3750
rect 659 3746 847 3750
rect 851 3746 895 3750
rect 899 3746 1055 3750
rect 1059 3746 1151 3750
rect 1155 3746 1279 3750
rect 1283 3746 1415 3750
rect 1419 3746 1511 3750
rect 1515 3746 1679 3750
rect 1683 3746 1751 3750
rect 1755 3746 1935 3750
rect 1939 3746 1947 3750
rect 91 3745 1947 3746
rect 1953 3745 1954 3751
rect 1946 3689 1947 3695
rect 1953 3694 3811 3695
rect 1953 3690 1975 3694
rect 1979 3690 2143 3694
rect 2147 3690 2231 3694
rect 2235 3690 2279 3694
rect 2283 3690 2415 3694
rect 2419 3690 2447 3694
rect 2451 3690 2551 3694
rect 2555 3690 2663 3694
rect 2667 3690 2687 3694
rect 2691 3690 2823 3694
rect 2827 3690 2871 3694
rect 2875 3690 2967 3694
rect 2971 3690 3079 3694
rect 3083 3690 3111 3694
rect 3115 3690 3263 3694
rect 3267 3690 3287 3694
rect 3291 3690 3423 3694
rect 3427 3690 3495 3694
rect 3499 3690 3583 3694
rect 3587 3690 3679 3694
rect 3683 3690 3799 3694
rect 3803 3690 3811 3694
rect 1953 3689 3811 3690
rect 3817 3689 3818 3695
rect 3810 3673 3811 3679
rect 3817 3678 5695 3679
rect 3817 3674 3839 3678
rect 3843 3674 3887 3678
rect 3891 3674 4047 3678
rect 4051 3674 4247 3678
rect 4251 3674 4439 3678
rect 4443 3674 4479 3678
rect 4483 3674 4647 3678
rect 4651 3674 4727 3678
rect 4731 3674 4863 3678
rect 4867 3674 4999 3678
rect 5003 3674 5095 3678
rect 5099 3674 5279 3678
rect 5283 3674 5327 3678
rect 5331 3674 5543 3678
rect 5547 3674 5663 3678
rect 5667 3674 5695 3678
rect 3817 3673 5695 3674
rect 5701 3673 5702 3679
rect 96 3625 97 3631
rect 103 3630 1959 3631
rect 103 3626 111 3630
rect 115 3626 131 3630
rect 135 3626 203 3630
rect 207 3626 315 3630
rect 319 3626 403 3630
rect 407 3626 539 3630
rect 543 3626 627 3630
rect 631 3626 787 3630
rect 791 3626 867 3630
rect 871 3626 1043 3630
rect 1047 3626 1123 3630
rect 1127 3626 1315 3630
rect 1319 3626 1387 3630
rect 1391 3626 1587 3630
rect 1591 3626 1651 3630
rect 1655 3626 1935 3630
rect 1939 3626 1959 3630
rect 103 3625 1959 3626
rect 1965 3625 1966 3631
rect 1958 3561 1959 3567
rect 1965 3566 3823 3567
rect 1965 3562 1975 3566
rect 1979 3562 2163 3566
rect 2167 3562 2203 3566
rect 2207 3562 2299 3566
rect 2303 3562 2419 3566
rect 2423 3562 2435 3566
rect 2439 3562 2571 3566
rect 2575 3562 2635 3566
rect 2639 3562 2843 3566
rect 2847 3562 3051 3566
rect 3055 3562 3259 3566
rect 3263 3562 3467 3566
rect 3471 3562 3651 3566
rect 3655 3562 3799 3566
rect 3803 3562 3823 3566
rect 1965 3561 3823 3562
rect 3829 3561 3830 3567
rect 3822 3549 3823 3555
rect 3829 3554 5707 3555
rect 3829 3550 3839 3554
rect 3843 3550 3859 3554
rect 3863 3550 3995 3554
rect 3999 3550 4019 3554
rect 4023 3550 4131 3554
rect 4135 3550 4219 3554
rect 4223 3550 4267 3554
rect 4271 3550 4403 3554
rect 4407 3550 4451 3554
rect 4455 3550 4539 3554
rect 4543 3550 4699 3554
rect 4703 3550 4891 3554
rect 4895 3550 4971 3554
rect 4975 3550 5099 3554
rect 5103 3550 5251 3554
rect 5255 3550 5315 3554
rect 5319 3550 5515 3554
rect 5519 3550 5663 3554
rect 5667 3550 5707 3554
rect 3829 3549 5707 3550
rect 5713 3549 5714 3555
rect 84 3501 85 3507
rect 91 3506 1947 3507
rect 91 3502 111 3506
rect 115 3502 159 3506
rect 163 3502 335 3506
rect 339 3502 343 3506
rect 347 3502 551 3506
rect 555 3502 567 3506
rect 571 3502 791 3506
rect 795 3502 815 3506
rect 819 3502 1039 3506
rect 1043 3502 1071 3506
rect 1075 3502 1295 3506
rect 1299 3502 1343 3506
rect 1347 3502 1559 3506
rect 1563 3502 1615 3506
rect 1619 3502 1935 3506
rect 1939 3502 1947 3506
rect 91 3501 1947 3502
rect 1953 3501 1954 3507
rect 3810 3429 3811 3435
rect 3817 3434 5695 3435
rect 3817 3430 3839 3434
rect 3843 3430 3887 3434
rect 3891 3430 4023 3434
rect 4027 3430 4159 3434
rect 4163 3430 4295 3434
rect 4299 3430 4431 3434
rect 4435 3430 4567 3434
rect 4571 3430 4583 3434
rect 4587 3430 4727 3434
rect 4731 3430 4759 3434
rect 4763 3430 4919 3434
rect 4923 3430 4951 3434
rect 4955 3430 5127 3434
rect 5131 3430 5151 3434
rect 5155 3430 5343 3434
rect 5347 3430 5359 3434
rect 5363 3430 5543 3434
rect 5547 3430 5663 3434
rect 5667 3430 5695 3434
rect 3817 3429 5695 3430
rect 5701 3429 5702 3435
rect 1946 3413 1947 3419
rect 1953 3418 3811 3419
rect 1953 3414 1975 3418
rect 1979 3414 2191 3418
rect 2195 3414 2231 3418
rect 2235 3414 2327 3418
rect 2331 3414 2463 3418
rect 2467 3414 2583 3418
rect 2587 3414 2599 3418
rect 2603 3414 2951 3418
rect 2955 3414 3327 3418
rect 3331 3414 3679 3418
rect 3683 3414 3799 3418
rect 3803 3414 3811 3418
rect 1953 3413 3811 3414
rect 3817 3413 3818 3419
rect 96 3381 97 3387
rect 103 3386 1959 3387
rect 103 3382 111 3386
rect 115 3382 131 3386
rect 135 3382 299 3386
rect 303 3382 307 3386
rect 311 3382 507 3386
rect 511 3382 523 3386
rect 527 3382 731 3386
rect 735 3382 763 3386
rect 767 3382 971 3386
rect 975 3382 1011 3386
rect 1015 3382 1219 3386
rect 1223 3382 1267 3386
rect 1271 3382 1475 3386
rect 1479 3382 1531 3386
rect 1535 3382 1935 3386
rect 1939 3382 1959 3386
rect 103 3381 1959 3382
rect 1965 3381 1966 3387
rect 1958 3301 1959 3307
rect 1965 3306 3823 3307
rect 1965 3302 1975 3306
rect 1979 3302 2203 3306
rect 2207 3302 2251 3306
rect 2255 3302 2475 3306
rect 2479 3302 2555 3306
rect 2559 3302 2691 3306
rect 2695 3302 2899 3306
rect 2903 3302 2923 3306
rect 2927 3302 3099 3306
rect 3103 3302 3291 3306
rect 3295 3302 3299 3306
rect 3303 3302 3483 3306
rect 3487 3302 3651 3306
rect 3655 3302 3799 3306
rect 3803 3302 3823 3306
rect 1965 3301 3823 3302
rect 3829 3306 5714 3307
rect 3829 3302 3839 3306
rect 3843 3302 3859 3306
rect 3863 3302 3995 3306
rect 3999 3302 4131 3306
rect 4135 3302 4267 3306
rect 4271 3302 4403 3306
rect 4407 3302 4555 3306
rect 4559 3302 4691 3306
rect 4695 3302 4731 3306
rect 4735 3302 4827 3306
rect 4831 3302 4923 3306
rect 4927 3302 4963 3306
rect 4967 3302 5099 3306
rect 5103 3302 5123 3306
rect 5127 3302 5235 3306
rect 5239 3302 5331 3306
rect 5335 3302 5515 3306
rect 5519 3302 5663 3306
rect 5667 3302 5714 3306
rect 3829 3301 5714 3302
rect 84 3265 85 3271
rect 91 3270 1947 3271
rect 91 3266 111 3270
rect 115 3266 159 3270
rect 163 3266 239 3270
rect 243 3266 327 3270
rect 331 3266 463 3270
rect 467 3266 535 3270
rect 539 3266 703 3270
rect 707 3266 759 3270
rect 763 3266 951 3270
rect 955 3266 999 3270
rect 1003 3266 1199 3270
rect 1203 3266 1247 3270
rect 1251 3266 1455 3270
rect 1459 3266 1503 3270
rect 1507 3266 1935 3270
rect 1939 3266 1947 3270
rect 91 3265 1947 3266
rect 1953 3265 1954 3271
rect 1946 3181 1947 3187
rect 1953 3186 3811 3187
rect 1953 3182 1975 3186
rect 1979 3182 2095 3186
rect 2099 3182 2279 3186
rect 2283 3182 2295 3186
rect 2299 3182 2487 3186
rect 2491 3182 2503 3186
rect 2507 3182 2679 3186
rect 2683 3182 2719 3186
rect 2723 3182 2871 3186
rect 2875 3182 2927 3186
rect 2931 3182 3055 3186
rect 3059 3182 3127 3186
rect 3131 3182 3231 3186
rect 3235 3182 3319 3186
rect 3323 3182 3415 3186
rect 3419 3182 3511 3186
rect 3515 3182 3599 3186
rect 3603 3182 3679 3186
rect 3683 3182 3799 3186
rect 3803 3182 3811 3186
rect 1953 3181 3811 3182
rect 3817 3186 5702 3187
rect 3817 3182 3839 3186
rect 3843 3182 4719 3186
rect 4723 3182 4855 3186
rect 4859 3182 4863 3186
rect 4867 3182 4991 3186
rect 4995 3182 4999 3186
rect 5003 3182 5127 3186
rect 5131 3182 5135 3186
rect 5139 3182 5263 3186
rect 5267 3182 5271 3186
rect 5275 3182 5407 3186
rect 5411 3182 5543 3186
rect 5547 3182 5663 3186
rect 5667 3182 5702 3186
rect 3817 3181 5702 3182
rect 96 3149 97 3155
rect 103 3154 1959 3155
rect 103 3150 111 3154
rect 115 3150 211 3154
rect 215 3150 379 3154
rect 383 3150 435 3154
rect 439 3150 563 3154
rect 567 3150 675 3154
rect 679 3150 755 3154
rect 759 3150 923 3154
rect 927 3150 955 3154
rect 959 3150 1163 3154
rect 1167 3150 1171 3154
rect 1175 3150 1371 3154
rect 1375 3150 1427 3154
rect 1431 3150 1935 3154
rect 1939 3150 1959 3154
rect 103 3149 1959 3150
rect 1965 3149 1966 3155
rect 1958 3057 1959 3063
rect 1965 3062 3823 3063
rect 1965 3058 1975 3062
rect 1979 3058 1995 3062
rect 1999 3058 2067 3062
rect 2071 3058 2131 3062
rect 2135 3058 2267 3062
rect 2271 3058 2403 3062
rect 2407 3058 2459 3062
rect 2463 3058 2539 3062
rect 2543 3058 2651 3062
rect 2655 3058 2683 3062
rect 2687 3058 2835 3062
rect 2839 3058 2843 3062
rect 2847 3058 2987 3062
rect 2991 3058 3027 3062
rect 3031 3058 3139 3062
rect 3143 3058 3203 3062
rect 3207 3058 3291 3062
rect 3295 3058 3387 3062
rect 3391 3058 3571 3062
rect 3575 3058 3799 3062
rect 3803 3058 3823 3062
rect 1965 3057 3823 3058
rect 3829 3062 5714 3063
rect 3829 3058 3839 3062
rect 3843 3058 4483 3062
rect 4487 3058 4635 3062
rect 4639 3058 4803 3062
rect 4807 3058 4835 3062
rect 4839 3058 4971 3062
rect 4975 3058 4979 3062
rect 4983 3058 5107 3062
rect 5111 3058 5163 3062
rect 5167 3058 5243 3062
rect 5247 3058 5347 3062
rect 5351 3058 5379 3062
rect 5383 3058 5515 3062
rect 5519 3058 5663 3062
rect 5667 3058 5714 3062
rect 3829 3057 5714 3058
rect 84 3021 85 3027
rect 91 3026 1947 3027
rect 91 3022 111 3026
rect 115 3022 407 3026
rect 411 3022 575 3026
rect 579 3022 591 3026
rect 595 3022 783 3026
rect 787 3022 799 3026
rect 803 3022 983 3026
rect 987 3022 1047 3026
rect 1051 3022 1191 3026
rect 1195 3022 1303 3026
rect 1307 3022 1399 3026
rect 1403 3022 1567 3026
rect 1571 3022 1815 3026
rect 1819 3022 1935 3026
rect 1939 3022 1947 3026
rect 91 3021 1947 3022
rect 1953 3021 1954 3027
rect 1946 2945 1947 2951
rect 1953 2950 3811 2951
rect 1953 2946 1975 2950
rect 1979 2946 2023 2950
rect 2027 2946 2159 2950
rect 2163 2946 2295 2950
rect 2299 2946 2431 2950
rect 2435 2946 2567 2950
rect 2571 2946 2591 2950
rect 2595 2946 2711 2950
rect 2715 2946 2863 2950
rect 2867 2946 2887 2950
rect 2891 2946 3015 2950
rect 3019 2946 3167 2950
rect 3171 2946 3183 2950
rect 3187 2946 3319 2950
rect 3323 2946 3799 2950
rect 3803 2946 3811 2950
rect 1953 2945 3811 2946
rect 3817 2945 3818 2951
rect 3810 2921 3811 2927
rect 3817 2926 5695 2927
rect 3817 2922 3839 2926
rect 3843 2922 4047 2926
rect 4051 2922 4295 2926
rect 4299 2922 4511 2926
rect 4515 2922 4583 2926
rect 4587 2922 4663 2926
rect 4667 2922 4831 2926
rect 4835 2922 4895 2926
rect 4899 2922 5007 2926
rect 5011 2922 5191 2926
rect 5195 2922 5231 2926
rect 5235 2922 5375 2926
rect 5379 2922 5543 2926
rect 5547 2922 5663 2926
rect 5667 2922 5695 2926
rect 3817 2921 5695 2922
rect 5701 2921 5702 2927
rect 96 2901 97 2907
rect 103 2906 1959 2907
rect 103 2902 111 2906
rect 115 2902 427 2906
rect 431 2902 547 2906
rect 551 2902 563 2906
rect 567 2902 699 2906
rect 703 2902 771 2906
rect 775 2902 835 2906
rect 839 2902 971 2906
rect 975 2902 1019 2906
rect 1023 2902 1107 2906
rect 1111 2902 1243 2906
rect 1247 2902 1275 2906
rect 1279 2902 1379 2906
rect 1383 2902 1515 2906
rect 1519 2902 1539 2906
rect 1543 2902 1651 2906
rect 1655 2902 1787 2906
rect 1791 2902 1935 2906
rect 1939 2902 1959 2906
rect 103 2901 1959 2902
rect 1965 2901 1966 2907
rect 3822 2805 3823 2811
rect 3829 2810 5707 2811
rect 3829 2806 3839 2810
rect 3843 2806 3859 2810
rect 3863 2806 3995 2810
rect 3999 2806 4019 2810
rect 4023 2806 4131 2810
rect 4135 2806 4267 2810
rect 4271 2806 4403 2810
rect 4407 2806 4539 2810
rect 4543 2806 4555 2810
rect 4559 2806 4675 2810
rect 4679 2806 4811 2810
rect 4815 2806 4867 2810
rect 4871 2806 5203 2810
rect 5207 2806 5515 2810
rect 5519 2806 5663 2810
rect 5667 2806 5707 2810
rect 3829 2805 5707 2806
rect 5713 2805 5714 2811
rect 84 2781 85 2787
rect 91 2786 1947 2787
rect 91 2782 111 2786
rect 115 2782 455 2786
rect 459 2782 463 2786
rect 467 2782 591 2786
rect 595 2782 623 2786
rect 627 2782 727 2786
rect 731 2782 783 2786
rect 787 2782 863 2786
rect 867 2782 935 2786
rect 939 2782 999 2786
rect 1003 2782 1087 2786
rect 1091 2782 1135 2786
rect 1139 2782 1239 2786
rect 1243 2782 1271 2786
rect 1275 2782 1383 2786
rect 1387 2782 1407 2786
rect 1411 2782 1535 2786
rect 1539 2782 1543 2786
rect 1547 2782 1679 2786
rect 1683 2782 1815 2786
rect 1819 2782 1935 2786
rect 1939 2782 1947 2786
rect 91 2781 1947 2782
rect 1953 2781 1954 2787
rect 1958 2777 1959 2783
rect 1965 2782 3823 2783
rect 1965 2778 1975 2782
rect 1979 2778 1995 2782
rect 1999 2778 2267 2782
rect 2271 2778 2563 2782
rect 2567 2778 2859 2782
rect 2863 2778 3059 2782
rect 3063 2778 3155 2782
rect 3159 2778 3195 2782
rect 3199 2778 3331 2782
rect 3335 2778 3799 2782
rect 3803 2778 3823 2782
rect 1965 2777 3823 2778
rect 3829 2777 3830 2783
rect 3810 2693 3811 2699
rect 3817 2698 5695 2699
rect 3817 2694 3839 2698
rect 3843 2694 3887 2698
rect 3891 2694 4023 2698
rect 4027 2694 4055 2698
rect 4059 2694 4159 2698
rect 4163 2694 4295 2698
rect 4299 2694 4303 2698
rect 4307 2694 4431 2698
rect 4435 2694 4567 2698
rect 4571 2694 4583 2698
rect 4587 2694 4703 2698
rect 4707 2694 4839 2698
rect 4843 2694 4895 2698
rect 4899 2694 5231 2698
rect 5235 2694 5543 2698
rect 5547 2694 5663 2698
rect 5667 2694 5695 2698
rect 3817 2693 5695 2694
rect 5701 2693 5702 2699
rect 96 2665 97 2671
rect 103 2670 1959 2671
rect 103 2666 111 2670
rect 115 2666 355 2670
rect 359 2666 435 2670
rect 439 2666 539 2670
rect 543 2666 595 2670
rect 599 2666 715 2670
rect 719 2666 755 2670
rect 759 2666 883 2670
rect 887 2666 907 2670
rect 911 2666 1043 2670
rect 1047 2666 1059 2670
rect 1063 2666 1203 2670
rect 1207 2666 1211 2670
rect 1215 2666 1355 2670
rect 1359 2666 1507 2670
rect 1511 2666 1651 2670
rect 1655 2666 1787 2670
rect 1791 2666 1935 2670
rect 1939 2666 1959 2670
rect 103 2665 1959 2666
rect 1965 2665 1966 2671
rect 1946 2641 1947 2647
rect 1953 2646 3811 2647
rect 1953 2642 1975 2646
rect 1979 2642 3087 2646
rect 3091 2642 3135 2646
rect 3139 2642 3223 2646
rect 3227 2642 3271 2646
rect 3275 2642 3359 2646
rect 3363 2642 3407 2646
rect 3411 2642 3543 2646
rect 3547 2642 3679 2646
rect 3683 2642 3799 2646
rect 3803 2642 3811 2646
rect 1953 2641 3811 2642
rect 3817 2641 3818 2647
rect 3822 2577 3823 2583
rect 3829 2582 5707 2583
rect 3829 2578 3839 2582
rect 3843 2578 4027 2582
rect 4031 2578 4259 2582
rect 4263 2578 4275 2582
rect 4279 2578 4475 2582
rect 4479 2578 4555 2582
rect 4559 2578 4715 2582
rect 4719 2578 4867 2582
rect 4871 2578 4979 2582
rect 4983 2578 5203 2582
rect 5207 2578 5259 2582
rect 5263 2578 5515 2582
rect 5519 2578 5663 2582
rect 5667 2578 5707 2582
rect 3829 2577 5707 2578
rect 5713 2577 5714 2583
rect 84 2553 85 2559
rect 91 2558 1947 2559
rect 91 2554 111 2558
rect 115 2554 231 2558
rect 235 2554 383 2558
rect 387 2554 423 2558
rect 427 2554 567 2558
rect 571 2554 623 2558
rect 627 2554 743 2558
rect 747 2554 823 2558
rect 827 2554 911 2558
rect 915 2554 1023 2558
rect 1027 2554 1071 2558
rect 1075 2554 1223 2558
rect 1227 2554 1231 2558
rect 1235 2554 1383 2558
rect 1387 2554 1423 2558
rect 1427 2554 1535 2558
rect 1539 2554 1631 2558
rect 1635 2554 1679 2558
rect 1683 2554 1815 2558
rect 1819 2554 1935 2558
rect 1939 2554 1947 2558
rect 91 2553 1947 2554
rect 1953 2553 1954 2559
rect 1958 2521 1959 2527
rect 1965 2526 3823 2527
rect 1965 2522 1975 2526
rect 1979 2522 1995 2526
rect 1999 2522 2235 2526
rect 2239 2522 2483 2526
rect 2487 2522 2715 2526
rect 2719 2522 2939 2526
rect 2943 2522 3107 2526
rect 3111 2522 3155 2526
rect 3159 2522 3243 2526
rect 3247 2522 3363 2526
rect 3367 2522 3379 2526
rect 3383 2522 3515 2526
rect 3519 2522 3579 2526
rect 3583 2522 3651 2526
rect 3655 2522 3799 2526
rect 3803 2522 3823 2526
rect 1965 2521 3823 2522
rect 3829 2521 3830 2527
rect 3810 2461 3811 2467
rect 3817 2466 5695 2467
rect 3817 2462 3839 2466
rect 3843 2462 4287 2466
rect 4291 2462 4503 2466
rect 4507 2462 4663 2466
rect 4667 2462 4743 2466
rect 4747 2462 4847 2466
rect 4851 2462 5007 2466
rect 5011 2462 5023 2466
rect 5027 2462 5199 2466
rect 5203 2462 5287 2466
rect 5291 2462 5383 2466
rect 5387 2462 5543 2466
rect 5547 2462 5663 2466
rect 5667 2462 5695 2466
rect 3817 2461 5695 2462
rect 5701 2461 5702 2467
rect 96 2421 97 2427
rect 103 2426 1959 2427
rect 103 2422 111 2426
rect 115 2422 203 2426
rect 207 2422 219 2426
rect 223 2422 395 2426
rect 399 2422 403 2426
rect 407 2422 595 2426
rect 599 2422 787 2426
rect 791 2422 795 2426
rect 799 2422 979 2426
rect 983 2422 995 2426
rect 999 2422 1195 2426
rect 1199 2422 1395 2426
rect 1399 2422 1603 2426
rect 1607 2422 1787 2426
rect 1791 2422 1935 2426
rect 1939 2422 1959 2426
rect 103 2421 1959 2422
rect 1965 2421 1966 2427
rect 1946 2409 1947 2415
rect 1953 2414 3811 2415
rect 1953 2410 1975 2414
rect 1979 2410 2023 2414
rect 2027 2410 2159 2414
rect 2163 2410 2263 2414
rect 2267 2410 2295 2414
rect 2299 2410 2431 2414
rect 2435 2410 2511 2414
rect 2515 2410 2567 2414
rect 2571 2410 2711 2414
rect 2715 2410 2743 2414
rect 2747 2410 2855 2414
rect 2859 2410 2967 2414
rect 2971 2410 3007 2414
rect 3011 2410 3159 2414
rect 3163 2410 3183 2414
rect 3187 2410 3311 2414
rect 3315 2410 3391 2414
rect 3395 2410 3607 2414
rect 3611 2410 3799 2414
rect 3803 2410 3811 2414
rect 1953 2409 3811 2410
rect 3817 2409 3818 2415
rect 3822 2345 3823 2351
rect 3829 2350 5707 2351
rect 3829 2346 3839 2350
rect 3843 2346 4635 2350
rect 4639 2346 4675 2350
rect 4679 2346 4819 2350
rect 4823 2346 4963 2350
rect 4967 2346 4995 2350
rect 4999 2346 5115 2350
rect 5119 2346 5171 2350
rect 5175 2346 5267 2350
rect 5271 2346 5355 2350
rect 5359 2346 5419 2350
rect 5423 2346 5515 2350
rect 5519 2346 5663 2350
rect 5667 2346 5707 2350
rect 3829 2345 5707 2346
rect 5713 2345 5714 2351
rect 84 2305 85 2311
rect 91 2310 1947 2311
rect 91 2306 111 2310
rect 115 2306 247 2310
rect 251 2306 399 2310
rect 403 2306 431 2310
rect 435 2306 535 2310
rect 539 2306 623 2310
rect 627 2306 671 2310
rect 675 2306 807 2310
rect 811 2306 815 2310
rect 819 2306 943 2310
rect 947 2306 1007 2310
rect 1011 2306 1935 2310
rect 1939 2306 1947 2310
rect 91 2305 1947 2306
rect 1953 2305 1954 2311
rect 1958 2293 1959 2299
rect 1965 2298 3823 2299
rect 1965 2294 1975 2298
rect 1979 2294 1995 2298
rect 1999 2294 2043 2298
rect 2047 2294 2131 2298
rect 2135 2294 2179 2298
rect 2183 2294 2267 2298
rect 2271 2294 2315 2298
rect 2319 2294 2403 2298
rect 2407 2294 2451 2298
rect 2455 2294 2539 2298
rect 2543 2294 2587 2298
rect 2591 2294 2683 2298
rect 2687 2294 2723 2298
rect 2727 2294 2827 2298
rect 2831 2294 2859 2298
rect 2863 2294 2979 2298
rect 2983 2294 2995 2298
rect 2999 2294 3131 2298
rect 3135 2294 3283 2298
rect 3287 2294 3799 2298
rect 3803 2294 3823 2298
rect 1965 2293 3823 2294
rect 3829 2293 3830 2299
rect 3810 2221 3811 2227
rect 3817 2226 5695 2227
rect 3817 2222 3839 2226
rect 3843 2222 3887 2226
rect 3891 2222 4167 2226
rect 4171 2222 4455 2226
rect 4459 2222 4703 2226
rect 4707 2222 4719 2226
rect 4723 2222 4847 2226
rect 4851 2222 4975 2226
rect 4979 2222 4991 2226
rect 4995 2222 5143 2226
rect 5147 2222 5231 2226
rect 5235 2222 5295 2226
rect 5299 2222 5447 2226
rect 5451 2222 5487 2226
rect 5491 2222 5663 2226
rect 5667 2222 5695 2226
rect 3817 2221 5695 2222
rect 5701 2221 5702 2227
rect 1946 2195 1947 2201
rect 1953 2195 1978 2201
rect 96 2185 97 2191
rect 103 2190 1959 2191
rect 103 2186 111 2190
rect 115 2186 323 2190
rect 327 2186 371 2190
rect 375 2186 459 2190
rect 463 2186 507 2190
rect 511 2186 595 2190
rect 599 2186 643 2190
rect 647 2186 731 2190
rect 735 2186 779 2190
rect 783 2186 867 2190
rect 871 2186 915 2190
rect 919 2186 1935 2190
rect 1939 2186 1959 2190
rect 103 2185 1959 2186
rect 1965 2185 1966 2191
rect 1972 2187 1978 2195
rect 1972 2186 3811 2187
rect 1972 2182 1975 2186
rect 1979 2182 2023 2186
rect 2027 2182 2071 2186
rect 2075 2182 2207 2186
rect 2211 2182 2239 2186
rect 2243 2182 2343 2186
rect 2347 2182 2479 2186
rect 2483 2182 2487 2186
rect 2491 2182 2615 2186
rect 2619 2182 2727 2186
rect 2731 2182 2751 2186
rect 2755 2182 2887 2186
rect 2891 2182 2967 2186
rect 2971 2182 3023 2186
rect 3027 2182 3159 2186
rect 3163 2182 3207 2186
rect 3211 2182 3455 2186
rect 3459 2182 3679 2186
rect 3683 2182 3799 2186
rect 3803 2182 3811 2186
rect 1972 2181 3811 2182
rect 3817 2181 3818 2187
rect 3822 2109 3823 2115
rect 3829 2114 5707 2115
rect 3829 2110 3839 2114
rect 3843 2110 3859 2114
rect 3863 2110 4083 2114
rect 4087 2110 4139 2114
rect 4143 2110 4323 2114
rect 4327 2110 4427 2114
rect 4431 2110 4547 2114
rect 4551 2110 4691 2114
rect 4695 2110 4755 2114
rect 4759 2110 4947 2114
rect 4951 2110 5139 2114
rect 5143 2110 5203 2114
rect 5207 2110 5323 2114
rect 5327 2110 5459 2114
rect 5463 2110 5515 2114
rect 5519 2110 5663 2114
rect 5667 2110 5707 2114
rect 3829 2109 5707 2110
rect 5713 2109 5714 2115
rect 1958 2053 1959 2059
rect 1965 2058 3823 2059
rect 1965 2054 1975 2058
rect 1979 2054 1995 2058
rect 1999 2054 2211 2058
rect 2215 2054 2459 2058
rect 2463 2054 2699 2058
rect 2703 2054 2707 2058
rect 2711 2054 2939 2058
rect 2943 2054 2963 2058
rect 2967 2054 3179 2058
rect 3183 2054 3219 2058
rect 3223 2054 3427 2058
rect 3431 2054 3483 2058
rect 3487 2054 3651 2058
rect 3655 2054 3799 2058
rect 3803 2054 3823 2058
rect 1965 2053 3823 2054
rect 3829 2053 3830 2059
rect 84 2041 85 2047
rect 91 2046 1947 2047
rect 91 2042 111 2046
rect 115 2042 319 2046
rect 323 2042 351 2046
rect 355 2042 479 2046
rect 483 2042 487 2046
rect 491 2042 623 2046
rect 627 2042 663 2046
rect 667 2042 759 2046
rect 763 2042 871 2046
rect 875 2042 895 2046
rect 899 2042 1095 2046
rect 1099 2042 1335 2046
rect 1339 2042 1583 2046
rect 1587 2042 1815 2046
rect 1819 2042 1935 2046
rect 1939 2042 1947 2046
rect 91 2041 1947 2042
rect 1953 2041 1954 2047
rect 3810 1997 3811 2003
rect 3817 2002 5695 2003
rect 3817 1998 3839 2002
rect 3843 1998 3887 2002
rect 3891 1998 4111 2002
rect 4115 1998 4167 2002
rect 4171 1998 4351 2002
rect 4355 1998 4463 2002
rect 4467 1998 4575 2002
rect 4579 1998 4743 2002
rect 4747 1998 4783 2002
rect 4787 1998 4975 2002
rect 4979 1998 5007 2002
rect 5011 1998 5167 2002
rect 5171 1998 5271 2002
rect 5275 1998 5351 2002
rect 5355 1998 5543 2002
rect 5547 1998 5663 2002
rect 5667 1998 5695 2002
rect 3817 1997 5695 1998
rect 5701 1997 5702 2003
rect 1946 1933 1947 1939
rect 1953 1938 3811 1939
rect 1953 1934 1975 1938
rect 1979 1934 2023 1938
rect 2027 1934 2159 1938
rect 2163 1934 2239 1938
rect 2243 1934 2439 1938
rect 2443 1934 2487 1938
rect 2491 1934 2703 1938
rect 2707 1934 2735 1938
rect 2739 1934 2959 1938
rect 2963 1934 2991 1938
rect 2995 1934 3207 1938
rect 3211 1934 3247 1938
rect 3251 1934 3455 1938
rect 3459 1934 3511 1938
rect 3515 1934 3679 1938
rect 3683 1934 3799 1938
rect 3803 1934 3811 1938
rect 1953 1933 3811 1934
rect 3817 1933 3818 1939
rect 96 1921 97 1927
rect 103 1926 1959 1927
rect 103 1922 111 1926
rect 115 1922 187 1926
rect 191 1922 291 1926
rect 295 1922 419 1926
rect 423 1922 451 1926
rect 455 1922 635 1926
rect 639 1922 651 1926
rect 655 1922 843 1926
rect 847 1922 883 1926
rect 887 1922 1067 1926
rect 1071 1922 1115 1926
rect 1119 1922 1307 1926
rect 1311 1922 1347 1926
rect 1351 1922 1555 1926
rect 1559 1922 1579 1926
rect 1583 1922 1787 1926
rect 1791 1922 1935 1926
rect 1939 1922 1959 1926
rect 103 1921 1959 1922
rect 1965 1921 1966 1927
rect 3822 1873 3823 1879
rect 3829 1878 5707 1879
rect 3829 1874 3839 1878
rect 3843 1874 3859 1878
rect 3863 1874 4139 1878
rect 4143 1874 4435 1878
rect 4439 1874 4539 1878
rect 4543 1874 4715 1878
rect 4719 1874 4723 1878
rect 4727 1874 4915 1878
rect 4919 1874 4979 1878
rect 4983 1874 5115 1878
rect 5119 1874 5243 1878
rect 5247 1874 5323 1878
rect 5327 1874 5515 1878
rect 5519 1874 5663 1878
rect 5667 1874 5707 1878
rect 3829 1873 5707 1874
rect 5713 1873 5714 1879
rect 1958 1813 1959 1819
rect 1965 1818 3823 1819
rect 1965 1814 1975 1818
rect 1979 1814 2131 1818
rect 2135 1814 2307 1818
rect 2311 1814 2411 1818
rect 2415 1814 2499 1818
rect 2503 1814 2675 1818
rect 2679 1814 2691 1818
rect 2695 1814 2883 1818
rect 2887 1814 2931 1818
rect 2935 1814 3067 1818
rect 3071 1814 3179 1818
rect 3183 1814 3251 1818
rect 3255 1814 3427 1818
rect 3431 1814 3443 1818
rect 3447 1814 3635 1818
rect 3639 1814 3651 1818
rect 3655 1814 3799 1818
rect 3803 1814 3823 1818
rect 1965 1813 3823 1814
rect 3829 1813 3830 1819
rect 84 1797 85 1803
rect 91 1802 1947 1803
rect 91 1798 111 1802
rect 115 1798 159 1802
rect 163 1798 215 1802
rect 219 1798 367 1802
rect 371 1798 447 1802
rect 451 1798 591 1802
rect 595 1798 679 1802
rect 683 1798 799 1802
rect 803 1798 911 1802
rect 915 1798 999 1802
rect 1003 1798 1143 1802
rect 1147 1798 1191 1802
rect 1195 1798 1375 1802
rect 1379 1798 1559 1802
rect 1563 1798 1607 1802
rect 1611 1798 1751 1802
rect 1755 1798 1815 1802
rect 1819 1798 1935 1802
rect 1939 1798 1947 1802
rect 91 1797 1947 1798
rect 1953 1797 1954 1803
rect 3810 1753 3811 1759
rect 3817 1758 5695 1759
rect 3817 1754 3839 1758
rect 3843 1754 4383 1758
rect 4387 1754 4567 1758
rect 4571 1754 4599 1758
rect 4603 1754 4751 1758
rect 4755 1754 4831 1758
rect 4835 1754 4943 1758
rect 4947 1754 5071 1758
rect 5075 1754 5143 1758
rect 5147 1754 5319 1758
rect 5323 1754 5351 1758
rect 5355 1754 5543 1758
rect 5547 1754 5663 1758
rect 5667 1754 5695 1758
rect 3817 1753 5695 1754
rect 5701 1753 5702 1759
rect 1946 1701 1947 1707
rect 1953 1706 3811 1707
rect 1953 1702 1975 1706
rect 1979 1702 2335 1706
rect 2339 1702 2471 1706
rect 2475 1702 2527 1706
rect 2531 1702 2607 1706
rect 2611 1702 2719 1706
rect 2723 1702 2743 1706
rect 2747 1702 2879 1706
rect 2883 1702 2911 1706
rect 2915 1702 3023 1706
rect 3027 1702 3095 1706
rect 3099 1702 3175 1706
rect 3179 1702 3279 1706
rect 3283 1702 3327 1706
rect 3331 1702 3471 1706
rect 3475 1702 3663 1706
rect 3667 1702 3799 1706
rect 3803 1702 3811 1706
rect 1953 1701 3811 1702
rect 3817 1701 3818 1707
rect 96 1677 97 1683
rect 103 1682 1959 1683
rect 103 1678 111 1682
rect 115 1678 131 1682
rect 135 1678 339 1682
rect 343 1678 355 1682
rect 359 1678 563 1682
rect 567 1678 595 1682
rect 599 1678 771 1682
rect 775 1678 835 1682
rect 839 1678 971 1682
rect 975 1678 1067 1682
rect 1071 1678 1163 1682
rect 1167 1678 1307 1682
rect 1311 1678 1347 1682
rect 1351 1678 1531 1682
rect 1535 1678 1547 1682
rect 1551 1678 1723 1682
rect 1727 1678 1935 1682
rect 1939 1678 1959 1682
rect 103 1677 1959 1678
rect 1965 1677 1966 1683
rect 3822 1629 3823 1635
rect 3829 1634 5707 1635
rect 3829 1630 3839 1634
rect 3843 1630 3907 1634
rect 3911 1630 4123 1634
rect 4127 1630 4355 1634
rect 4359 1630 4363 1634
rect 4367 1630 4571 1634
rect 4575 1630 4627 1634
rect 4631 1630 4803 1634
rect 4807 1630 4907 1634
rect 4911 1630 5043 1634
rect 5047 1630 5195 1634
rect 5199 1630 5291 1634
rect 5295 1630 5491 1634
rect 5495 1630 5515 1634
rect 5519 1630 5663 1634
rect 5667 1630 5707 1634
rect 3829 1629 5707 1630
rect 5713 1629 5714 1635
rect 1958 1589 1959 1595
rect 1965 1594 3823 1595
rect 1965 1590 1975 1594
rect 1979 1590 2355 1594
rect 2359 1590 2443 1594
rect 2447 1590 2563 1594
rect 2567 1590 2579 1594
rect 2583 1590 2715 1594
rect 2719 1590 2779 1594
rect 2783 1590 2851 1594
rect 2855 1590 2995 1594
rect 2999 1590 3003 1594
rect 3007 1590 3147 1594
rect 3151 1590 3227 1594
rect 3231 1590 3299 1594
rect 3303 1590 3459 1594
rect 3463 1590 3799 1594
rect 3803 1590 3823 1594
rect 1965 1589 3823 1590
rect 3829 1589 3830 1595
rect 84 1561 85 1567
rect 91 1566 1947 1567
rect 91 1562 111 1566
rect 115 1562 159 1566
rect 163 1562 359 1566
rect 363 1562 383 1566
rect 387 1562 575 1566
rect 579 1562 623 1566
rect 627 1562 783 1566
rect 787 1562 863 1566
rect 867 1562 983 1566
rect 987 1562 1095 1566
rect 1099 1562 1183 1566
rect 1187 1562 1335 1566
rect 1339 1562 1375 1566
rect 1379 1562 1575 1566
rect 1579 1562 1935 1566
rect 1939 1562 1947 1566
rect 91 1561 1947 1562
rect 1953 1561 1954 1567
rect 3810 1517 3811 1523
rect 3817 1522 5695 1523
rect 3817 1518 3839 1522
rect 3843 1518 3887 1522
rect 3891 1518 3935 1522
rect 3939 1518 4023 1522
rect 4027 1518 4151 1522
rect 4155 1518 4159 1522
rect 4163 1518 4295 1522
rect 4299 1518 4391 1522
rect 4395 1518 4479 1522
rect 4483 1518 4655 1522
rect 4659 1518 4695 1522
rect 4699 1518 4935 1522
rect 4939 1518 5191 1522
rect 5195 1518 5223 1522
rect 5227 1518 5447 1522
rect 5451 1518 5519 1522
rect 5523 1518 5663 1522
rect 5667 1518 5695 1522
rect 3817 1517 5695 1518
rect 5701 1517 5702 1523
rect 1946 1477 1947 1483
rect 1953 1482 3811 1483
rect 1953 1478 1975 1482
rect 1979 1478 2023 1482
rect 2027 1478 2159 1482
rect 2163 1478 2327 1482
rect 2331 1478 2383 1482
rect 2387 1478 2543 1482
rect 2547 1478 2591 1482
rect 2595 1478 2799 1482
rect 2803 1478 2807 1482
rect 2811 1478 3031 1482
rect 3035 1478 3087 1482
rect 3091 1478 3255 1482
rect 3259 1478 3391 1482
rect 3395 1478 3487 1482
rect 3491 1478 3679 1482
rect 3683 1478 3799 1482
rect 3803 1478 3811 1482
rect 1953 1477 3811 1478
rect 3817 1477 3818 1483
rect 96 1429 97 1435
rect 103 1434 1959 1435
rect 103 1430 111 1434
rect 115 1430 131 1434
rect 135 1430 235 1434
rect 239 1430 331 1434
rect 335 1430 507 1434
rect 511 1430 547 1434
rect 551 1430 755 1434
rect 759 1430 779 1434
rect 783 1430 955 1434
rect 959 1430 1059 1434
rect 1063 1430 1155 1434
rect 1159 1430 1339 1434
rect 1343 1430 1347 1434
rect 1351 1430 1547 1434
rect 1551 1430 1935 1434
rect 1939 1430 1959 1434
rect 103 1429 1959 1430
rect 1965 1429 1966 1435
rect 3822 1393 3823 1399
rect 3829 1398 5707 1399
rect 3829 1394 3839 1398
rect 3843 1394 3859 1398
rect 3863 1394 3995 1398
rect 3999 1394 4131 1398
rect 4135 1394 4147 1398
rect 4151 1394 4267 1398
rect 4271 1394 4363 1398
rect 4367 1394 4451 1398
rect 4455 1394 4611 1398
rect 4615 1394 4667 1398
rect 4671 1394 4891 1398
rect 4895 1394 4907 1398
rect 4911 1394 5163 1398
rect 5167 1394 5195 1398
rect 5199 1394 5419 1398
rect 5423 1394 5499 1398
rect 5503 1394 5663 1398
rect 5667 1394 5707 1398
rect 3829 1393 5707 1394
rect 5713 1393 5714 1399
rect 1958 1365 1959 1371
rect 1965 1370 3823 1371
rect 1965 1366 1975 1370
rect 1979 1366 1995 1370
rect 1999 1366 2131 1370
rect 2135 1366 2299 1370
rect 2303 1366 2491 1370
rect 2495 1366 2515 1370
rect 2519 1366 2771 1370
rect 2775 1366 3019 1370
rect 3023 1366 3059 1370
rect 3063 1366 3363 1370
rect 3367 1366 3555 1370
rect 3559 1366 3651 1370
rect 3655 1366 3799 1370
rect 3803 1366 3823 1370
rect 1965 1365 3823 1366
rect 3829 1365 3830 1371
rect 84 1313 85 1319
rect 91 1318 1947 1319
rect 91 1314 111 1318
rect 115 1314 159 1318
rect 163 1314 263 1318
rect 267 1314 383 1318
rect 387 1314 535 1318
rect 539 1314 599 1318
rect 603 1314 799 1318
rect 803 1314 807 1318
rect 811 1314 991 1318
rect 995 1314 1087 1318
rect 1091 1314 1167 1318
rect 1171 1314 1335 1318
rect 1339 1314 1367 1318
rect 1371 1314 1503 1318
rect 1507 1314 1671 1318
rect 1675 1314 1815 1318
rect 1819 1314 1935 1318
rect 1939 1314 1947 1318
rect 91 1313 1947 1314
rect 1953 1313 1954 1319
rect 3810 1281 3811 1287
rect 3817 1286 5695 1287
rect 3817 1282 3839 1286
rect 3843 1282 3887 1286
rect 3891 1282 4023 1286
rect 4027 1282 4167 1286
rect 4171 1282 4175 1286
rect 4179 1282 4335 1286
rect 4339 1282 4391 1286
rect 4395 1282 4511 1286
rect 4515 1282 4639 1286
rect 4643 1282 4703 1286
rect 4707 1282 4903 1286
rect 4907 1282 4919 1286
rect 4923 1282 5119 1286
rect 5123 1282 5223 1286
rect 5227 1282 5343 1286
rect 5347 1282 5527 1286
rect 5531 1282 5543 1286
rect 5547 1282 5663 1286
rect 5667 1282 5695 1286
rect 3817 1281 5695 1282
rect 5701 1281 5702 1287
rect 1946 1203 1947 1209
rect 1953 1203 1978 1209
rect 96 1193 97 1199
rect 103 1198 1959 1199
rect 103 1194 111 1198
rect 115 1194 131 1198
rect 135 1194 147 1198
rect 151 1194 323 1198
rect 327 1194 355 1198
rect 359 1194 499 1198
rect 503 1194 571 1198
rect 575 1194 675 1198
rect 679 1194 771 1198
rect 775 1194 851 1198
rect 855 1194 963 1198
rect 967 1194 1019 1198
rect 1023 1194 1139 1198
rect 1143 1194 1179 1198
rect 1183 1194 1307 1198
rect 1311 1194 1331 1198
rect 1335 1194 1475 1198
rect 1479 1194 1483 1198
rect 1487 1194 1643 1198
rect 1647 1194 1787 1198
rect 1791 1194 1935 1198
rect 1939 1194 1959 1198
rect 103 1193 1959 1194
rect 1965 1193 1966 1199
rect 1972 1195 1978 1203
rect 1972 1194 3811 1195
rect 1972 1190 1975 1194
rect 1979 1190 2023 1194
rect 2027 1190 2519 1194
rect 2523 1190 2743 1194
rect 2747 1190 3047 1194
rect 3051 1190 3359 1194
rect 3363 1190 3583 1194
rect 3587 1190 3679 1194
rect 3683 1190 3799 1194
rect 3803 1190 3811 1194
rect 1972 1189 3811 1190
rect 3817 1189 3818 1195
rect 3822 1165 3823 1171
rect 3829 1170 5707 1171
rect 3829 1166 3839 1170
rect 3843 1166 3859 1170
rect 3863 1166 3995 1170
rect 3999 1166 4139 1170
rect 4143 1166 4307 1170
rect 4311 1166 4483 1170
rect 4487 1166 4675 1170
rect 4679 1166 4811 1170
rect 4815 1166 4875 1170
rect 4879 1166 4947 1170
rect 4951 1166 5083 1170
rect 5087 1166 5091 1170
rect 5095 1166 5227 1170
rect 5231 1166 5315 1170
rect 5319 1166 5379 1170
rect 5383 1166 5515 1170
rect 5519 1166 5663 1170
rect 5667 1166 5707 1170
rect 3829 1165 5707 1166
rect 5713 1165 5714 1171
rect 1958 1077 1959 1083
rect 1965 1082 3823 1083
rect 1965 1078 1975 1082
rect 1979 1078 2243 1082
rect 2247 1078 2379 1082
rect 2383 1078 2523 1082
rect 2527 1078 2675 1082
rect 2679 1078 2715 1082
rect 2719 1078 2827 1082
rect 2831 1078 2987 1082
rect 2991 1078 3019 1082
rect 3023 1078 3155 1082
rect 3159 1078 3323 1082
rect 3327 1078 3331 1082
rect 3335 1078 3499 1082
rect 3503 1078 3651 1082
rect 3655 1078 3799 1082
rect 3803 1078 3823 1082
rect 1965 1077 3823 1078
rect 3829 1077 3830 1083
rect 84 1061 85 1067
rect 91 1066 1947 1067
rect 91 1062 111 1066
rect 115 1062 159 1066
rect 163 1062 175 1066
rect 179 1062 351 1066
rect 355 1062 447 1066
rect 451 1062 527 1066
rect 531 1062 703 1066
rect 707 1062 775 1066
rect 779 1062 879 1066
rect 883 1062 1047 1066
rect 1051 1062 1111 1066
rect 1115 1062 1207 1066
rect 1211 1062 1359 1066
rect 1363 1062 1455 1066
rect 1459 1062 1511 1066
rect 1515 1062 1671 1066
rect 1675 1062 1807 1066
rect 1811 1062 1815 1066
rect 1819 1062 1935 1066
rect 1939 1062 1947 1066
rect 91 1061 1947 1062
rect 1953 1061 1954 1067
rect 3810 1049 3811 1055
rect 3817 1054 5695 1055
rect 3817 1050 3839 1054
rect 3843 1050 4807 1054
rect 4811 1050 4839 1054
rect 4843 1050 4943 1054
rect 4947 1050 4975 1054
rect 4979 1050 5079 1054
rect 5083 1050 5111 1054
rect 5115 1050 5215 1054
rect 5219 1050 5255 1054
rect 5259 1050 5351 1054
rect 5355 1050 5407 1054
rect 5411 1050 5487 1054
rect 5491 1050 5543 1054
rect 5547 1050 5663 1054
rect 5667 1050 5695 1054
rect 3817 1049 5695 1050
rect 5701 1049 5702 1055
rect 1946 961 1947 967
rect 1953 966 3811 967
rect 1953 962 1975 966
rect 1979 962 2271 966
rect 2275 962 2279 966
rect 2283 962 2407 966
rect 2411 962 2495 966
rect 2499 962 2551 966
rect 2555 962 2703 966
rect 2707 962 2711 966
rect 2715 962 2855 966
rect 2859 962 2911 966
rect 2915 962 3015 966
rect 3019 962 3103 966
rect 3107 962 3183 966
rect 3187 962 3295 966
rect 3299 962 3351 966
rect 3355 962 3479 966
rect 3483 962 3527 966
rect 3531 962 3671 966
rect 3675 962 3679 966
rect 3683 962 3799 966
rect 3803 962 3811 966
rect 1953 961 3811 962
rect 3817 961 3818 967
rect 96 945 97 951
rect 103 950 1959 951
rect 103 946 111 950
rect 115 946 131 950
rect 135 946 339 950
rect 343 946 419 950
rect 423 946 595 950
rect 599 946 747 950
rect 751 946 875 950
rect 879 946 1083 950
rect 1087 946 1179 950
rect 1183 946 1427 950
rect 1431 946 1491 950
rect 1495 946 1779 950
rect 1783 946 1787 950
rect 1791 946 1935 950
rect 1939 946 1959 950
rect 103 945 1959 946
rect 1965 945 1966 951
rect 3822 933 3823 939
rect 3829 938 5707 939
rect 3829 934 3839 938
rect 3843 934 4355 938
rect 4359 934 4571 938
rect 4575 934 4779 938
rect 4783 934 4803 938
rect 4807 934 4915 938
rect 4919 934 5043 938
rect 5047 934 5051 938
rect 5055 934 5187 938
rect 5191 934 5291 938
rect 5295 934 5323 938
rect 5327 934 5459 938
rect 5463 934 5515 938
rect 5519 934 5663 938
rect 5667 934 5707 938
rect 3829 933 5707 934
rect 5713 933 5714 939
rect 1958 845 1959 851
rect 1965 850 3823 851
rect 1965 846 1975 850
rect 1979 846 1995 850
rect 1999 846 2131 850
rect 2135 846 2251 850
rect 2255 846 2283 850
rect 2287 846 2443 850
rect 2447 846 2467 850
rect 2471 846 2603 850
rect 2607 846 2683 850
rect 2687 846 2763 850
rect 2767 846 2883 850
rect 2887 846 2923 850
rect 2927 846 3075 850
rect 3079 846 3083 850
rect 3087 846 3243 850
rect 3247 846 3267 850
rect 3271 846 3403 850
rect 3407 846 3451 850
rect 3455 846 3643 850
rect 3647 846 3799 850
rect 3803 846 3823 850
rect 1965 845 3823 846
rect 3829 845 3830 851
rect 84 821 85 827
rect 91 826 1947 827
rect 91 822 111 826
rect 115 822 159 826
rect 163 822 367 826
rect 371 822 383 826
rect 387 822 623 826
rect 627 822 631 826
rect 635 822 887 826
rect 891 822 903 826
rect 907 822 1143 826
rect 1147 822 1207 826
rect 1211 822 1519 826
rect 1523 822 1815 826
rect 1819 822 1935 826
rect 1939 822 1947 826
rect 91 821 1947 822
rect 1953 821 1954 827
rect 3810 817 3811 823
rect 3817 822 5695 823
rect 3817 818 3839 822
rect 3843 818 3959 822
rect 3963 818 4207 822
rect 4211 818 4383 822
rect 4387 818 4495 822
rect 4499 818 4599 822
rect 4603 818 4815 822
rect 4819 818 4831 822
rect 4835 818 5071 822
rect 5075 818 5151 822
rect 5155 818 5319 822
rect 5323 818 5487 822
rect 5491 818 5543 822
rect 5547 818 5663 822
rect 5667 818 5695 822
rect 3817 817 5695 818
rect 5701 817 5702 823
rect 1946 733 1947 739
rect 1953 738 3811 739
rect 1953 734 1975 738
rect 1979 734 2023 738
rect 2027 734 2159 738
rect 2163 734 2183 738
rect 2187 734 2311 738
rect 2315 734 2439 738
rect 2443 734 2471 738
rect 2475 734 2631 738
rect 2635 734 2679 738
rect 2683 734 2791 738
rect 2795 734 2903 738
rect 2907 734 2951 738
rect 2955 734 3111 738
rect 3115 734 3271 738
rect 3275 734 3311 738
rect 3315 734 3431 738
rect 3435 734 3503 738
rect 3507 734 3679 738
rect 3683 734 3799 738
rect 3803 734 3811 738
rect 1953 733 3811 734
rect 3817 733 3818 739
rect 96 709 97 715
rect 103 714 1959 715
rect 103 710 111 714
rect 115 710 131 714
rect 135 710 355 714
rect 359 710 603 714
rect 607 710 699 714
rect 703 710 835 714
rect 839 710 859 714
rect 863 710 971 714
rect 975 710 1107 714
rect 1111 710 1115 714
rect 1119 710 1243 714
rect 1247 710 1379 714
rect 1383 710 1515 714
rect 1519 710 1651 714
rect 1655 710 1787 714
rect 1791 710 1935 714
rect 1939 710 1959 714
rect 103 709 1959 710
rect 1965 709 1966 715
rect 3822 693 3823 699
rect 3829 698 5707 699
rect 3829 694 3839 698
rect 3843 694 3859 698
rect 3863 694 3931 698
rect 3935 694 3995 698
rect 3999 694 4147 698
rect 4151 694 4179 698
rect 4183 694 4355 698
rect 4359 694 4467 698
rect 4471 694 4595 698
rect 4599 694 4787 698
rect 4791 694 4867 698
rect 4871 694 5123 698
rect 5127 694 5163 698
rect 5167 694 5459 698
rect 5463 694 5663 698
rect 5667 694 5707 698
rect 3829 693 5707 694
rect 5713 693 5714 699
rect 84 597 85 603
rect 91 602 1947 603
rect 91 598 111 602
rect 115 598 159 602
rect 163 598 375 602
rect 379 598 599 602
rect 603 598 727 602
rect 731 598 807 602
rect 811 598 863 602
rect 867 598 999 602
rect 1003 598 1135 602
rect 1139 598 1175 602
rect 1179 598 1271 602
rect 1275 598 1343 602
rect 1347 598 1407 602
rect 1411 598 1511 602
rect 1515 598 1543 602
rect 1547 598 1671 602
rect 1675 598 1679 602
rect 1683 598 1815 602
rect 1819 598 1935 602
rect 1939 598 1947 602
rect 91 597 1947 598
rect 1953 597 1954 603
rect 3810 581 3811 587
rect 3817 586 5695 587
rect 3817 582 3839 586
rect 3843 582 3887 586
rect 3891 582 4023 586
rect 4027 582 4159 586
rect 4163 582 4175 586
rect 4179 582 4295 586
rect 4299 582 4383 586
rect 4387 582 4431 586
rect 4435 582 4567 586
rect 4571 582 4623 586
rect 4627 582 4711 586
rect 4715 582 4879 586
rect 4883 582 4895 586
rect 4899 582 5063 586
rect 5067 582 5191 586
rect 5195 582 5255 586
rect 5259 582 5447 586
rect 5451 582 5487 586
rect 5491 582 5663 586
rect 5667 582 5695 586
rect 3817 581 5695 582
rect 5701 581 5702 587
rect 96 485 97 491
rect 103 490 1959 491
rect 103 486 111 490
rect 115 486 131 490
rect 135 486 347 490
rect 351 486 355 490
rect 359 486 571 490
rect 575 486 603 490
rect 607 486 779 490
rect 783 486 843 490
rect 847 486 971 490
rect 975 486 1083 490
rect 1087 486 1147 490
rect 1151 486 1315 490
rect 1319 486 1323 490
rect 1327 486 1483 490
rect 1487 486 1563 490
rect 1567 486 1643 490
rect 1647 486 1787 490
rect 1791 486 1935 490
rect 1939 486 1959 490
rect 103 485 1959 486
rect 1965 485 1966 491
rect 3822 469 3823 475
rect 3829 474 5707 475
rect 3829 470 3839 474
rect 3843 470 3859 474
rect 3863 470 3995 474
rect 3999 470 4115 474
rect 4119 470 4131 474
rect 4135 470 4267 474
rect 4271 470 4395 474
rect 4399 470 4403 474
rect 4407 470 4539 474
rect 4543 470 4675 474
rect 4679 470 4683 474
rect 4687 470 4851 474
rect 4855 470 4947 474
rect 4951 470 5035 474
rect 5039 470 5227 474
rect 5231 470 5419 474
rect 5423 470 5507 474
rect 5511 470 5663 474
rect 5667 470 5707 474
rect 3829 469 5707 470
rect 5713 469 5714 475
rect 1958 445 1959 451
rect 1965 450 3823 451
rect 1965 446 1975 450
rect 1979 446 1995 450
rect 1999 446 2155 450
rect 2159 446 2251 450
rect 2255 446 2411 450
rect 2415 446 2523 450
rect 2527 446 2651 450
rect 2655 446 2771 450
rect 2775 446 2875 450
rect 2879 446 3003 450
rect 3007 446 3083 450
rect 3087 446 3227 450
rect 3231 446 3283 450
rect 3287 446 3451 450
rect 3455 446 3475 450
rect 3479 446 3651 450
rect 3655 446 3799 450
rect 3803 446 3823 450
rect 1965 445 3823 446
rect 3829 445 3830 451
rect 84 357 85 363
rect 91 362 1947 363
rect 91 358 111 362
rect 115 358 159 362
rect 163 358 303 362
rect 307 358 383 362
rect 387 358 479 362
rect 483 358 631 362
rect 635 358 655 362
rect 659 358 831 362
rect 835 358 871 362
rect 875 358 1111 362
rect 1115 358 1351 362
rect 1355 358 1591 362
rect 1595 358 1815 362
rect 1819 358 1935 362
rect 1939 358 1947 362
rect 91 357 1947 358
rect 1953 357 1954 363
rect 3810 349 3811 355
rect 3817 354 5695 355
rect 3817 350 3839 354
rect 3843 350 3887 354
rect 3891 350 4143 354
rect 4147 350 4423 354
rect 4427 350 4703 354
rect 4707 350 4727 354
rect 4731 350 4895 354
rect 4899 350 4975 354
rect 4979 350 5063 354
rect 5067 350 5231 354
rect 5235 350 5255 354
rect 5259 350 5399 354
rect 5403 350 5535 354
rect 5539 350 5543 354
rect 5547 350 5663 354
rect 5667 350 5695 354
rect 3817 349 5695 350
rect 5701 349 5702 355
rect 1946 329 1947 335
rect 1953 334 3811 335
rect 1953 330 1975 334
rect 1979 330 2023 334
rect 2027 330 2159 334
rect 2163 330 2279 334
rect 2283 330 2295 334
rect 2299 330 2431 334
rect 2435 330 2551 334
rect 2555 330 2567 334
rect 2571 330 2703 334
rect 2707 330 2799 334
rect 2803 330 2839 334
rect 2843 330 2975 334
rect 2979 330 3031 334
rect 3035 330 3111 334
rect 3115 330 3247 334
rect 3251 330 3255 334
rect 3259 330 3383 334
rect 3387 330 3479 334
rect 3483 330 3519 334
rect 3523 330 3655 334
rect 3659 330 3679 334
rect 3683 330 3799 334
rect 3803 330 3811 334
rect 1953 329 3811 330
rect 3817 329 3818 335
rect 96 205 97 211
rect 103 210 1959 211
rect 103 206 111 210
rect 115 206 131 210
rect 135 206 267 210
rect 271 206 275 210
rect 279 206 403 210
rect 407 206 451 210
rect 455 206 539 210
rect 543 206 627 210
rect 631 206 675 210
rect 679 206 803 210
rect 807 206 811 210
rect 815 206 947 210
rect 951 206 1083 210
rect 1087 206 1935 210
rect 1939 206 1959 210
rect 103 205 1959 206
rect 1965 205 1966 211
rect 3822 197 3823 203
rect 3829 202 5707 203
rect 3829 198 3839 202
rect 3843 198 4291 202
rect 4295 198 4427 202
rect 4431 198 4563 202
rect 4567 198 4699 202
rect 4703 198 4835 202
rect 4839 198 4867 202
rect 4871 198 4971 202
rect 4975 198 5035 202
rect 5039 198 5107 202
rect 5111 198 5203 202
rect 5207 198 5243 202
rect 5247 198 5371 202
rect 5375 198 5379 202
rect 5383 198 5515 202
rect 5519 198 5663 202
rect 5667 198 5707 202
rect 3829 197 5707 198
rect 5713 197 5714 203
rect 1958 185 1959 191
rect 1965 190 3823 191
rect 1965 186 1975 190
rect 1979 186 1995 190
rect 1999 186 2131 190
rect 2135 186 2267 190
rect 2271 186 2403 190
rect 2407 186 2539 190
rect 2543 186 2675 190
rect 2679 186 2811 190
rect 2815 186 2947 190
rect 2951 186 3083 190
rect 3087 186 3219 190
rect 3223 186 3355 190
rect 3359 186 3491 190
rect 3495 186 3627 190
rect 3631 186 3799 190
rect 3803 186 3823 190
rect 1965 185 3823 186
rect 3829 185 3830 191
rect 84 93 85 99
rect 91 98 1947 99
rect 91 94 111 98
rect 115 94 159 98
rect 163 94 295 98
rect 299 94 431 98
rect 435 94 567 98
rect 571 94 703 98
rect 707 94 839 98
rect 843 94 975 98
rect 979 94 1111 98
rect 1115 94 1935 98
rect 1939 94 1947 98
rect 91 93 1947 94
rect 1953 93 1954 99
rect 3810 85 3811 91
rect 3817 90 5695 91
rect 3817 86 3839 90
rect 3843 86 4319 90
rect 4323 86 4455 90
rect 4459 86 4591 90
rect 4595 86 4727 90
rect 4731 86 4863 90
rect 4867 86 4999 90
rect 5003 86 5135 90
rect 5139 86 5271 90
rect 5275 86 5407 90
rect 5411 86 5543 90
rect 5547 86 5663 90
rect 5667 86 5695 90
rect 3817 85 5695 86
rect 5701 85 5702 91
rect 1946 73 1947 79
rect 1953 78 3811 79
rect 1953 74 1975 78
rect 1979 74 2023 78
rect 2027 74 2159 78
rect 2163 74 2295 78
rect 2299 74 2431 78
rect 2435 74 2567 78
rect 2571 74 2703 78
rect 2707 74 2839 78
rect 2843 74 2975 78
rect 2979 74 3111 78
rect 3115 74 3247 78
rect 3251 74 3383 78
rect 3387 74 3519 78
rect 3523 74 3655 78
rect 3659 74 3799 78
rect 3803 74 3811 78
rect 1953 73 3811 74
rect 3817 73 3818 79
<< m5c >>
rect 1947 5753 1953 5759
rect 3811 5753 3817 5759
rect 85 5713 91 5719
rect 1947 5713 1953 5719
rect 3811 5677 3817 5683
rect 5695 5677 5701 5683
rect 1959 5641 1965 5647
rect 3823 5641 3829 5647
rect 97 5573 103 5579
rect 1959 5573 1965 5579
rect 3823 5565 3829 5571
rect 5707 5565 5713 5571
rect 1947 5529 1953 5535
rect 3811 5529 3817 5535
rect 85 5453 91 5459
rect 1947 5453 1953 5459
rect 3811 5417 3817 5423
rect 5695 5417 5701 5423
rect 1959 5369 1965 5375
rect 3823 5369 3829 5375
rect 97 5317 103 5323
rect 1959 5317 1965 5323
rect 3823 5273 3829 5279
rect 5707 5273 5713 5279
rect 1947 5257 1953 5263
rect 3811 5257 3817 5263
rect 85 5197 91 5203
rect 1947 5197 1953 5203
rect 3811 5147 3817 5153
rect 1959 5137 1965 5143
rect 3823 5137 3829 5143
rect 5695 5137 5701 5143
rect 97 5065 103 5071
rect 1959 5065 1965 5071
rect 3823 5009 3829 5015
rect 5707 5009 5713 5015
rect 1947 5001 1953 5007
rect 3811 5001 3817 5007
rect 85 4941 91 4947
rect 1947 4941 1953 4947
rect 3811 4891 3817 4897
rect 1959 4881 1965 4887
rect 3823 4881 3829 4887
rect 5695 4881 5701 4887
rect 97 4829 103 4835
rect 1959 4829 1965 4835
rect 3823 4761 3829 4767
rect 5707 4761 5713 4767
rect 1947 4721 1953 4727
rect 3811 4721 3817 4727
rect 85 4697 91 4703
rect 1947 4697 1953 4703
rect 3811 4645 3817 4651
rect 5695 4645 5701 4651
rect 1959 4605 1965 4611
rect 3823 4605 3829 4611
rect 97 4569 103 4575
rect 1959 4569 1965 4575
rect 3823 4529 3829 4535
rect 5707 4529 5713 4535
rect 1947 4485 1953 4491
rect 3811 4485 3817 4491
rect 85 4441 91 4447
rect 1947 4441 1953 4447
rect 3811 4417 3817 4423
rect 5695 4417 5701 4423
rect 1959 4357 1965 4363
rect 3823 4357 3829 4363
rect 97 4329 103 4335
rect 1959 4329 1965 4335
rect 3823 4293 3829 4299
rect 5707 4293 5713 4299
rect 1947 4217 1953 4223
rect 3811 4217 3817 4223
rect 85 4205 91 4211
rect 1947 4205 1953 4211
rect 3811 4181 3817 4187
rect 5695 4181 5701 4187
rect 97 4093 103 4099
rect 1959 4093 1965 4099
rect 1959 4069 1965 4075
rect 3823 4069 3829 4075
rect 3823 4033 3829 4039
rect 5707 4033 5713 4039
rect 85 3977 91 3983
rect 1947 3977 1953 3983
rect 1947 3929 1953 3935
rect 3811 3929 3817 3935
rect 3811 3921 3817 3927
rect 5695 3921 5701 3927
rect 97 3861 103 3867
rect 1959 3861 1965 3867
rect 1959 3809 1965 3815
rect 3823 3809 3829 3815
rect 85 3745 91 3751
rect 1947 3745 1953 3751
rect 1947 3689 1953 3695
rect 3811 3689 3817 3695
rect 3811 3673 3817 3679
rect 5695 3673 5701 3679
rect 97 3625 103 3631
rect 1959 3625 1965 3631
rect 1959 3561 1965 3567
rect 3823 3561 3829 3567
rect 3823 3549 3829 3555
rect 5707 3549 5713 3555
rect 85 3501 91 3507
rect 1947 3501 1953 3507
rect 3811 3429 3817 3435
rect 5695 3429 5701 3435
rect 1947 3413 1953 3419
rect 3811 3413 3817 3419
rect 97 3381 103 3387
rect 1959 3381 1965 3387
rect 1959 3301 1965 3307
rect 3823 3301 3829 3307
rect 85 3265 91 3271
rect 1947 3265 1953 3271
rect 1947 3181 1953 3187
rect 3811 3181 3817 3187
rect 97 3149 103 3155
rect 1959 3149 1965 3155
rect 1959 3057 1965 3063
rect 3823 3057 3829 3063
rect 85 3021 91 3027
rect 1947 3021 1953 3027
rect 1947 2945 1953 2951
rect 3811 2945 3817 2951
rect 3811 2921 3817 2927
rect 5695 2921 5701 2927
rect 97 2901 103 2907
rect 1959 2901 1965 2907
rect 3823 2805 3829 2811
rect 5707 2805 5713 2811
rect 85 2781 91 2787
rect 1947 2781 1953 2787
rect 1959 2777 1965 2783
rect 3823 2777 3829 2783
rect 3811 2693 3817 2699
rect 5695 2693 5701 2699
rect 97 2665 103 2671
rect 1959 2665 1965 2671
rect 1947 2641 1953 2647
rect 3811 2641 3817 2647
rect 3823 2577 3829 2583
rect 5707 2577 5713 2583
rect 85 2553 91 2559
rect 1947 2553 1953 2559
rect 1959 2521 1965 2527
rect 3823 2521 3829 2527
rect 3811 2461 3817 2467
rect 5695 2461 5701 2467
rect 97 2421 103 2427
rect 1959 2421 1965 2427
rect 1947 2409 1953 2415
rect 3811 2409 3817 2415
rect 3823 2345 3829 2351
rect 5707 2345 5713 2351
rect 85 2305 91 2311
rect 1947 2305 1953 2311
rect 1959 2293 1965 2299
rect 3823 2293 3829 2299
rect 3811 2221 3817 2227
rect 5695 2221 5701 2227
rect 1947 2195 1953 2201
rect 97 2185 103 2191
rect 1959 2185 1965 2191
rect 3811 2181 3817 2187
rect 3823 2109 3829 2115
rect 5707 2109 5713 2115
rect 1959 2053 1965 2059
rect 3823 2053 3829 2059
rect 85 2041 91 2047
rect 1947 2041 1953 2047
rect 3811 1997 3817 2003
rect 5695 1997 5701 2003
rect 1947 1933 1953 1939
rect 3811 1933 3817 1939
rect 97 1921 103 1927
rect 1959 1921 1965 1927
rect 3823 1873 3829 1879
rect 5707 1873 5713 1879
rect 1959 1813 1965 1819
rect 3823 1813 3829 1819
rect 85 1797 91 1803
rect 1947 1797 1953 1803
rect 3811 1753 3817 1759
rect 5695 1753 5701 1759
rect 1947 1701 1953 1707
rect 3811 1701 3817 1707
rect 97 1677 103 1683
rect 1959 1677 1965 1683
rect 3823 1629 3829 1635
rect 5707 1629 5713 1635
rect 1959 1589 1965 1595
rect 3823 1589 3829 1595
rect 85 1561 91 1567
rect 1947 1561 1953 1567
rect 3811 1517 3817 1523
rect 5695 1517 5701 1523
rect 1947 1477 1953 1483
rect 3811 1477 3817 1483
rect 97 1429 103 1435
rect 1959 1429 1965 1435
rect 3823 1393 3829 1399
rect 5707 1393 5713 1399
rect 1959 1365 1965 1371
rect 3823 1365 3829 1371
rect 85 1313 91 1319
rect 1947 1313 1953 1319
rect 3811 1281 3817 1287
rect 5695 1281 5701 1287
rect 1947 1203 1953 1209
rect 97 1193 103 1199
rect 1959 1193 1965 1199
rect 3811 1189 3817 1195
rect 3823 1165 3829 1171
rect 5707 1165 5713 1171
rect 1959 1077 1965 1083
rect 3823 1077 3829 1083
rect 85 1061 91 1067
rect 1947 1061 1953 1067
rect 3811 1049 3817 1055
rect 5695 1049 5701 1055
rect 1947 961 1953 967
rect 3811 961 3817 967
rect 97 945 103 951
rect 1959 945 1965 951
rect 3823 933 3829 939
rect 5707 933 5713 939
rect 1959 845 1965 851
rect 3823 845 3829 851
rect 85 821 91 827
rect 1947 821 1953 827
rect 3811 817 3817 823
rect 5695 817 5701 823
rect 1947 733 1953 739
rect 3811 733 3817 739
rect 97 709 103 715
rect 1959 709 1965 715
rect 3823 693 3829 699
rect 5707 693 5713 699
rect 85 597 91 603
rect 1947 597 1953 603
rect 3811 581 3817 587
rect 5695 581 5701 587
rect 97 485 103 491
rect 1959 485 1965 491
rect 3823 469 3829 475
rect 5707 469 5713 475
rect 1959 445 1965 451
rect 3823 445 3829 451
rect 85 357 91 363
rect 1947 357 1953 363
rect 3811 349 3817 355
rect 5695 349 5701 355
rect 1947 329 1953 335
rect 3811 329 3817 335
rect 97 205 103 211
rect 1959 205 1965 211
rect 3823 197 3829 203
rect 5707 197 5713 203
rect 1959 185 1965 191
rect 3823 185 3829 191
rect 85 93 91 99
rect 1947 93 1953 99
rect 3811 85 3817 91
rect 5695 85 5701 91
rect 1947 73 1953 79
rect 3811 73 3817 79
<< m5 >>
rect 84 5719 92 5760
rect 84 5713 85 5719
rect 91 5713 92 5719
rect 84 5459 92 5713
rect 84 5453 85 5459
rect 91 5453 92 5459
rect 84 5203 92 5453
rect 84 5197 85 5203
rect 91 5197 92 5203
rect 84 4947 92 5197
rect 84 4941 85 4947
rect 91 4941 92 4947
rect 84 4703 92 4941
rect 84 4697 85 4703
rect 91 4697 92 4703
rect 84 4447 92 4697
rect 84 4441 85 4447
rect 91 4441 92 4447
rect 84 4211 92 4441
rect 84 4205 85 4211
rect 91 4205 92 4211
rect 84 3983 92 4205
rect 84 3977 85 3983
rect 91 3977 92 3983
rect 84 3751 92 3977
rect 84 3745 85 3751
rect 91 3745 92 3751
rect 84 3507 92 3745
rect 84 3501 85 3507
rect 91 3501 92 3507
rect 84 3271 92 3501
rect 84 3265 85 3271
rect 91 3265 92 3271
rect 84 3027 92 3265
rect 84 3021 85 3027
rect 91 3021 92 3027
rect 84 2787 92 3021
rect 84 2781 85 2787
rect 91 2781 92 2787
rect 84 2559 92 2781
rect 84 2553 85 2559
rect 91 2553 92 2559
rect 84 2311 92 2553
rect 84 2305 85 2311
rect 91 2305 92 2311
rect 84 2047 92 2305
rect 84 2041 85 2047
rect 91 2041 92 2047
rect 84 1803 92 2041
rect 84 1797 85 1803
rect 91 1797 92 1803
rect 84 1567 92 1797
rect 84 1561 85 1567
rect 91 1561 92 1567
rect 84 1319 92 1561
rect 84 1313 85 1319
rect 91 1313 92 1319
rect 84 1067 92 1313
rect 84 1061 85 1067
rect 91 1061 92 1067
rect 84 827 92 1061
rect 84 821 85 827
rect 91 821 92 827
rect 84 603 92 821
rect 84 597 85 603
rect 91 597 92 603
rect 84 363 92 597
rect 84 357 85 363
rect 91 357 92 363
rect 84 99 92 357
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 5579 104 5760
rect 96 5573 97 5579
rect 103 5573 104 5579
rect 96 5323 104 5573
rect 96 5317 97 5323
rect 103 5317 104 5323
rect 96 5071 104 5317
rect 96 5065 97 5071
rect 103 5065 104 5071
rect 96 4835 104 5065
rect 96 4829 97 4835
rect 103 4829 104 4835
rect 96 4575 104 4829
rect 96 4569 97 4575
rect 103 4569 104 4575
rect 96 4335 104 4569
rect 96 4329 97 4335
rect 103 4329 104 4335
rect 96 4099 104 4329
rect 96 4093 97 4099
rect 103 4093 104 4099
rect 96 3867 104 4093
rect 96 3861 97 3867
rect 103 3861 104 3867
rect 96 3631 104 3861
rect 96 3625 97 3631
rect 103 3625 104 3631
rect 96 3387 104 3625
rect 96 3381 97 3387
rect 103 3381 104 3387
rect 96 3155 104 3381
rect 96 3149 97 3155
rect 103 3149 104 3155
rect 96 2907 104 3149
rect 96 2901 97 2907
rect 103 2901 104 2907
rect 96 2671 104 2901
rect 96 2665 97 2671
rect 103 2665 104 2671
rect 96 2427 104 2665
rect 96 2421 97 2427
rect 103 2421 104 2427
rect 96 2191 104 2421
rect 96 2185 97 2191
rect 103 2185 104 2191
rect 96 1927 104 2185
rect 96 1921 97 1927
rect 103 1921 104 1927
rect 96 1683 104 1921
rect 96 1677 97 1683
rect 103 1677 104 1683
rect 96 1435 104 1677
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1199 104 1429
rect 96 1193 97 1199
rect 103 1193 104 1199
rect 96 951 104 1193
rect 96 945 97 951
rect 103 945 104 951
rect 96 715 104 945
rect 96 709 97 715
rect 103 709 104 715
rect 96 491 104 709
rect 96 485 97 491
rect 103 485 104 491
rect 96 211 104 485
rect 96 205 97 211
rect 103 205 104 211
rect 96 72 104 205
rect 1946 5759 1954 5760
rect 1946 5753 1947 5759
rect 1953 5753 1954 5759
rect 1946 5719 1954 5753
rect 1946 5713 1947 5719
rect 1953 5713 1954 5719
rect 1946 5535 1954 5713
rect 1946 5529 1947 5535
rect 1953 5529 1954 5535
rect 1946 5459 1954 5529
rect 1946 5453 1947 5459
rect 1953 5453 1954 5459
rect 1946 5263 1954 5453
rect 1946 5257 1947 5263
rect 1953 5257 1954 5263
rect 1946 5203 1954 5257
rect 1946 5197 1947 5203
rect 1953 5197 1954 5203
rect 1946 5007 1954 5197
rect 1946 5001 1947 5007
rect 1953 5001 1954 5007
rect 1946 4947 1954 5001
rect 1946 4941 1947 4947
rect 1953 4941 1954 4947
rect 1946 4727 1954 4941
rect 1946 4721 1947 4727
rect 1953 4721 1954 4727
rect 1946 4703 1954 4721
rect 1946 4697 1947 4703
rect 1953 4697 1954 4703
rect 1946 4491 1954 4697
rect 1946 4485 1947 4491
rect 1953 4485 1954 4491
rect 1946 4447 1954 4485
rect 1946 4441 1947 4447
rect 1953 4441 1954 4447
rect 1946 4223 1954 4441
rect 1946 4217 1947 4223
rect 1953 4217 1954 4223
rect 1946 4211 1954 4217
rect 1946 4205 1947 4211
rect 1953 4205 1954 4211
rect 1946 3983 1954 4205
rect 1946 3977 1947 3983
rect 1953 3977 1954 3983
rect 1946 3935 1954 3977
rect 1946 3929 1947 3935
rect 1953 3929 1954 3935
rect 1946 3751 1954 3929
rect 1946 3745 1947 3751
rect 1953 3745 1954 3751
rect 1946 3695 1954 3745
rect 1946 3689 1947 3695
rect 1953 3689 1954 3695
rect 1946 3507 1954 3689
rect 1946 3501 1947 3507
rect 1953 3501 1954 3507
rect 1946 3419 1954 3501
rect 1946 3413 1947 3419
rect 1953 3413 1954 3419
rect 1946 3271 1954 3413
rect 1946 3265 1947 3271
rect 1953 3265 1954 3271
rect 1946 3187 1954 3265
rect 1946 3181 1947 3187
rect 1953 3181 1954 3187
rect 1946 3027 1954 3181
rect 1946 3021 1947 3027
rect 1953 3021 1954 3027
rect 1946 2951 1954 3021
rect 1946 2945 1947 2951
rect 1953 2945 1954 2951
rect 1946 2787 1954 2945
rect 1946 2781 1947 2787
rect 1953 2781 1954 2787
rect 1946 2647 1954 2781
rect 1946 2641 1947 2647
rect 1953 2641 1954 2647
rect 1946 2559 1954 2641
rect 1946 2553 1947 2559
rect 1953 2553 1954 2559
rect 1946 2415 1954 2553
rect 1946 2409 1947 2415
rect 1953 2409 1954 2415
rect 1946 2311 1954 2409
rect 1946 2305 1947 2311
rect 1953 2305 1954 2311
rect 1946 2201 1954 2305
rect 1946 2195 1947 2201
rect 1953 2195 1954 2201
rect 1946 2047 1954 2195
rect 1946 2041 1947 2047
rect 1953 2041 1954 2047
rect 1946 1939 1954 2041
rect 1946 1933 1947 1939
rect 1953 1933 1954 1939
rect 1946 1803 1954 1933
rect 1946 1797 1947 1803
rect 1953 1797 1954 1803
rect 1946 1707 1954 1797
rect 1946 1701 1947 1707
rect 1953 1701 1954 1707
rect 1946 1567 1954 1701
rect 1946 1561 1947 1567
rect 1953 1561 1954 1567
rect 1946 1483 1954 1561
rect 1946 1477 1947 1483
rect 1953 1477 1954 1483
rect 1946 1319 1954 1477
rect 1946 1313 1947 1319
rect 1953 1313 1954 1319
rect 1946 1209 1954 1313
rect 1946 1203 1947 1209
rect 1953 1203 1954 1209
rect 1946 1067 1954 1203
rect 1946 1061 1947 1067
rect 1953 1061 1954 1067
rect 1946 967 1954 1061
rect 1946 961 1947 967
rect 1953 961 1954 967
rect 1946 827 1954 961
rect 1946 821 1947 827
rect 1953 821 1954 827
rect 1946 739 1954 821
rect 1946 733 1947 739
rect 1953 733 1954 739
rect 1946 603 1954 733
rect 1946 597 1947 603
rect 1953 597 1954 603
rect 1946 363 1954 597
rect 1946 357 1947 363
rect 1953 357 1954 363
rect 1946 335 1954 357
rect 1946 329 1947 335
rect 1953 329 1954 335
rect 1946 99 1954 329
rect 1946 93 1947 99
rect 1953 93 1954 99
rect 1946 79 1954 93
rect 1946 73 1947 79
rect 1953 73 1954 79
rect 1946 72 1954 73
rect 1958 5647 1966 5760
rect 1958 5641 1959 5647
rect 1965 5641 1966 5647
rect 1958 5579 1966 5641
rect 1958 5573 1959 5579
rect 1965 5573 1966 5579
rect 1958 5375 1966 5573
rect 1958 5369 1959 5375
rect 1965 5369 1966 5375
rect 1958 5323 1966 5369
rect 1958 5317 1959 5323
rect 1965 5317 1966 5323
rect 1958 5143 1966 5317
rect 1958 5137 1959 5143
rect 1965 5137 1966 5143
rect 1958 5071 1966 5137
rect 1958 5065 1959 5071
rect 1965 5065 1966 5071
rect 1958 4887 1966 5065
rect 1958 4881 1959 4887
rect 1965 4881 1966 4887
rect 1958 4835 1966 4881
rect 1958 4829 1959 4835
rect 1965 4829 1966 4835
rect 1958 4611 1966 4829
rect 1958 4605 1959 4611
rect 1965 4605 1966 4611
rect 1958 4575 1966 4605
rect 1958 4569 1959 4575
rect 1965 4569 1966 4575
rect 1958 4363 1966 4569
rect 1958 4357 1959 4363
rect 1965 4357 1966 4363
rect 1958 4335 1966 4357
rect 1958 4329 1959 4335
rect 1965 4329 1966 4335
rect 1958 4099 1966 4329
rect 1958 4093 1959 4099
rect 1965 4093 1966 4099
rect 1958 4075 1966 4093
rect 1958 4069 1959 4075
rect 1965 4069 1966 4075
rect 1958 3867 1966 4069
rect 1958 3861 1959 3867
rect 1965 3861 1966 3867
rect 1958 3815 1966 3861
rect 1958 3809 1959 3815
rect 1965 3809 1966 3815
rect 1958 3631 1966 3809
rect 1958 3625 1959 3631
rect 1965 3625 1966 3631
rect 1958 3567 1966 3625
rect 1958 3561 1959 3567
rect 1965 3561 1966 3567
rect 1958 3387 1966 3561
rect 1958 3381 1959 3387
rect 1965 3381 1966 3387
rect 1958 3307 1966 3381
rect 1958 3301 1959 3307
rect 1965 3301 1966 3307
rect 1958 3155 1966 3301
rect 1958 3149 1959 3155
rect 1965 3149 1966 3155
rect 1958 3063 1966 3149
rect 1958 3057 1959 3063
rect 1965 3057 1966 3063
rect 1958 2907 1966 3057
rect 1958 2901 1959 2907
rect 1965 2901 1966 2907
rect 1958 2783 1966 2901
rect 1958 2777 1959 2783
rect 1965 2777 1966 2783
rect 1958 2671 1966 2777
rect 1958 2665 1959 2671
rect 1965 2665 1966 2671
rect 1958 2527 1966 2665
rect 1958 2521 1959 2527
rect 1965 2521 1966 2527
rect 1958 2427 1966 2521
rect 1958 2421 1959 2427
rect 1965 2421 1966 2427
rect 1958 2299 1966 2421
rect 1958 2293 1959 2299
rect 1965 2293 1966 2299
rect 1958 2191 1966 2293
rect 1958 2185 1959 2191
rect 1965 2185 1966 2191
rect 1958 2059 1966 2185
rect 1958 2053 1959 2059
rect 1965 2053 1966 2059
rect 1958 1927 1966 2053
rect 1958 1921 1959 1927
rect 1965 1921 1966 1927
rect 1958 1819 1966 1921
rect 1958 1813 1959 1819
rect 1965 1813 1966 1819
rect 1958 1683 1966 1813
rect 1958 1677 1959 1683
rect 1965 1677 1966 1683
rect 1958 1595 1966 1677
rect 1958 1589 1959 1595
rect 1965 1589 1966 1595
rect 1958 1435 1966 1589
rect 1958 1429 1959 1435
rect 1965 1429 1966 1435
rect 1958 1371 1966 1429
rect 1958 1365 1959 1371
rect 1965 1365 1966 1371
rect 1958 1199 1966 1365
rect 1958 1193 1959 1199
rect 1965 1193 1966 1199
rect 1958 1083 1966 1193
rect 1958 1077 1959 1083
rect 1965 1077 1966 1083
rect 1958 951 1966 1077
rect 1958 945 1959 951
rect 1965 945 1966 951
rect 1958 851 1966 945
rect 1958 845 1959 851
rect 1965 845 1966 851
rect 1958 715 1966 845
rect 1958 709 1959 715
rect 1965 709 1966 715
rect 1958 491 1966 709
rect 1958 485 1959 491
rect 1965 485 1966 491
rect 1958 451 1966 485
rect 1958 445 1959 451
rect 1965 445 1966 451
rect 1958 211 1966 445
rect 1958 205 1959 211
rect 1965 205 1966 211
rect 1958 191 1966 205
rect 1958 185 1959 191
rect 1965 185 1966 191
rect 1958 72 1966 185
rect 3810 5759 3818 5760
rect 3810 5753 3811 5759
rect 3817 5753 3818 5759
rect 3810 5683 3818 5753
rect 3810 5677 3811 5683
rect 3817 5677 3818 5683
rect 3810 5535 3818 5677
rect 3810 5529 3811 5535
rect 3817 5529 3818 5535
rect 3810 5423 3818 5529
rect 3810 5417 3811 5423
rect 3817 5417 3818 5423
rect 3810 5263 3818 5417
rect 3810 5257 3811 5263
rect 3817 5257 3818 5263
rect 3810 5153 3818 5257
rect 3810 5147 3811 5153
rect 3817 5147 3818 5153
rect 3810 5007 3818 5147
rect 3810 5001 3811 5007
rect 3817 5001 3818 5007
rect 3810 4897 3818 5001
rect 3810 4891 3811 4897
rect 3817 4891 3818 4897
rect 3810 4727 3818 4891
rect 3810 4721 3811 4727
rect 3817 4721 3818 4727
rect 3810 4651 3818 4721
rect 3810 4645 3811 4651
rect 3817 4645 3818 4651
rect 3810 4491 3818 4645
rect 3810 4485 3811 4491
rect 3817 4485 3818 4491
rect 3810 4423 3818 4485
rect 3810 4417 3811 4423
rect 3817 4417 3818 4423
rect 3810 4223 3818 4417
rect 3810 4217 3811 4223
rect 3817 4217 3818 4223
rect 3810 4187 3818 4217
rect 3810 4181 3811 4187
rect 3817 4181 3818 4187
rect 3810 3935 3818 4181
rect 3810 3929 3811 3935
rect 3817 3929 3818 3935
rect 3810 3927 3818 3929
rect 3810 3921 3811 3927
rect 3817 3921 3818 3927
rect 3810 3695 3818 3921
rect 3810 3689 3811 3695
rect 3817 3689 3818 3695
rect 3810 3679 3818 3689
rect 3810 3673 3811 3679
rect 3817 3673 3818 3679
rect 3810 3435 3818 3673
rect 3810 3429 3811 3435
rect 3817 3429 3818 3435
rect 3810 3419 3818 3429
rect 3810 3413 3811 3419
rect 3817 3413 3818 3419
rect 3810 3187 3818 3413
rect 3810 3181 3811 3187
rect 3817 3181 3818 3187
rect 3810 2951 3818 3181
rect 3810 2945 3811 2951
rect 3817 2945 3818 2951
rect 3810 2927 3818 2945
rect 3810 2921 3811 2927
rect 3817 2921 3818 2927
rect 3810 2699 3818 2921
rect 3810 2693 3811 2699
rect 3817 2693 3818 2699
rect 3810 2647 3818 2693
rect 3810 2641 3811 2647
rect 3817 2641 3818 2647
rect 3810 2467 3818 2641
rect 3810 2461 3811 2467
rect 3817 2461 3818 2467
rect 3810 2415 3818 2461
rect 3810 2409 3811 2415
rect 3817 2409 3818 2415
rect 3810 2227 3818 2409
rect 3810 2221 3811 2227
rect 3817 2221 3818 2227
rect 3810 2187 3818 2221
rect 3810 2181 3811 2187
rect 3817 2181 3818 2187
rect 3810 2003 3818 2181
rect 3810 1997 3811 2003
rect 3817 1997 3818 2003
rect 3810 1939 3818 1997
rect 3810 1933 3811 1939
rect 3817 1933 3818 1939
rect 3810 1759 3818 1933
rect 3810 1753 3811 1759
rect 3817 1753 3818 1759
rect 3810 1707 3818 1753
rect 3810 1701 3811 1707
rect 3817 1701 3818 1707
rect 3810 1523 3818 1701
rect 3810 1517 3811 1523
rect 3817 1517 3818 1523
rect 3810 1483 3818 1517
rect 3810 1477 3811 1483
rect 3817 1477 3818 1483
rect 3810 1287 3818 1477
rect 3810 1281 3811 1287
rect 3817 1281 3818 1287
rect 3810 1195 3818 1281
rect 3810 1189 3811 1195
rect 3817 1189 3818 1195
rect 3810 1055 3818 1189
rect 3810 1049 3811 1055
rect 3817 1049 3818 1055
rect 3810 967 3818 1049
rect 3810 961 3811 967
rect 3817 961 3818 967
rect 3810 823 3818 961
rect 3810 817 3811 823
rect 3817 817 3818 823
rect 3810 739 3818 817
rect 3810 733 3811 739
rect 3817 733 3818 739
rect 3810 587 3818 733
rect 3810 581 3811 587
rect 3817 581 3818 587
rect 3810 355 3818 581
rect 3810 349 3811 355
rect 3817 349 3818 355
rect 3810 335 3818 349
rect 3810 329 3811 335
rect 3817 329 3818 335
rect 3810 91 3818 329
rect 3810 85 3811 91
rect 3817 85 3818 91
rect 3810 79 3818 85
rect 3810 73 3811 79
rect 3817 73 3818 79
rect 3810 72 3818 73
rect 3822 5647 3830 5760
rect 3822 5641 3823 5647
rect 3829 5641 3830 5647
rect 3822 5571 3830 5641
rect 3822 5565 3823 5571
rect 3829 5565 3830 5571
rect 3822 5375 3830 5565
rect 3822 5369 3823 5375
rect 3829 5369 3830 5375
rect 3822 5279 3830 5369
rect 3822 5273 3823 5279
rect 3829 5273 3830 5279
rect 3822 5143 3830 5273
rect 3822 5137 3823 5143
rect 3829 5137 3830 5143
rect 3822 5015 3830 5137
rect 3822 5009 3823 5015
rect 3829 5009 3830 5015
rect 3822 4887 3830 5009
rect 3822 4881 3823 4887
rect 3829 4881 3830 4887
rect 3822 4767 3830 4881
rect 3822 4761 3823 4767
rect 3829 4761 3830 4767
rect 3822 4611 3830 4761
rect 3822 4605 3823 4611
rect 3829 4605 3830 4611
rect 3822 4535 3830 4605
rect 3822 4529 3823 4535
rect 3829 4529 3830 4535
rect 3822 4363 3830 4529
rect 3822 4357 3823 4363
rect 3829 4357 3830 4363
rect 3822 4299 3830 4357
rect 3822 4293 3823 4299
rect 3829 4293 3830 4299
rect 3822 4075 3830 4293
rect 3822 4069 3823 4075
rect 3829 4069 3830 4075
rect 3822 4039 3830 4069
rect 3822 4033 3823 4039
rect 3829 4033 3830 4039
rect 3822 3815 3830 4033
rect 3822 3809 3823 3815
rect 3829 3809 3830 3815
rect 3822 3567 3830 3809
rect 3822 3561 3823 3567
rect 3829 3561 3830 3567
rect 3822 3555 3830 3561
rect 3822 3549 3823 3555
rect 3829 3549 3830 3555
rect 3822 3307 3830 3549
rect 3822 3301 3823 3307
rect 3829 3301 3830 3307
rect 3822 3063 3830 3301
rect 3822 3057 3823 3063
rect 3829 3057 3830 3063
rect 3822 2811 3830 3057
rect 3822 2805 3823 2811
rect 3829 2805 3830 2811
rect 3822 2783 3830 2805
rect 3822 2777 3823 2783
rect 3829 2777 3830 2783
rect 3822 2583 3830 2777
rect 3822 2577 3823 2583
rect 3829 2577 3830 2583
rect 3822 2527 3830 2577
rect 3822 2521 3823 2527
rect 3829 2521 3830 2527
rect 3822 2351 3830 2521
rect 3822 2345 3823 2351
rect 3829 2345 3830 2351
rect 3822 2299 3830 2345
rect 3822 2293 3823 2299
rect 3829 2293 3830 2299
rect 3822 2115 3830 2293
rect 3822 2109 3823 2115
rect 3829 2109 3830 2115
rect 3822 2059 3830 2109
rect 3822 2053 3823 2059
rect 3829 2053 3830 2059
rect 3822 1879 3830 2053
rect 3822 1873 3823 1879
rect 3829 1873 3830 1879
rect 3822 1819 3830 1873
rect 3822 1813 3823 1819
rect 3829 1813 3830 1819
rect 3822 1635 3830 1813
rect 3822 1629 3823 1635
rect 3829 1629 3830 1635
rect 3822 1595 3830 1629
rect 3822 1589 3823 1595
rect 3829 1589 3830 1595
rect 3822 1399 3830 1589
rect 3822 1393 3823 1399
rect 3829 1393 3830 1399
rect 3822 1371 3830 1393
rect 3822 1365 3823 1371
rect 3829 1365 3830 1371
rect 3822 1171 3830 1365
rect 3822 1165 3823 1171
rect 3829 1165 3830 1171
rect 3822 1083 3830 1165
rect 3822 1077 3823 1083
rect 3829 1077 3830 1083
rect 3822 939 3830 1077
rect 3822 933 3823 939
rect 3829 933 3830 939
rect 3822 851 3830 933
rect 3822 845 3823 851
rect 3829 845 3830 851
rect 3822 699 3830 845
rect 3822 693 3823 699
rect 3829 693 3830 699
rect 3822 475 3830 693
rect 3822 469 3823 475
rect 3829 469 3830 475
rect 3822 451 3830 469
rect 3822 445 3823 451
rect 3829 445 3830 451
rect 3822 203 3830 445
rect 3822 197 3823 203
rect 3829 197 3830 203
rect 3822 191 3830 197
rect 3822 185 3823 191
rect 3829 185 3830 191
rect 3822 72 3830 185
rect 5694 5683 5702 5760
rect 5694 5677 5695 5683
rect 5701 5677 5702 5683
rect 5694 5423 5702 5677
rect 5694 5417 5695 5423
rect 5701 5417 5702 5423
rect 5694 5143 5702 5417
rect 5694 5137 5695 5143
rect 5701 5137 5702 5143
rect 5694 4887 5702 5137
rect 5694 4881 5695 4887
rect 5701 4881 5702 4887
rect 5694 4651 5702 4881
rect 5694 4645 5695 4651
rect 5701 4645 5702 4651
rect 5694 4423 5702 4645
rect 5694 4417 5695 4423
rect 5701 4417 5702 4423
rect 5694 4187 5702 4417
rect 5694 4181 5695 4187
rect 5701 4181 5702 4187
rect 5694 3927 5702 4181
rect 5694 3921 5695 3927
rect 5701 3921 5702 3927
rect 5694 3679 5702 3921
rect 5694 3673 5695 3679
rect 5701 3673 5702 3679
rect 5694 3435 5702 3673
rect 5694 3429 5695 3435
rect 5701 3429 5702 3435
rect 5694 2927 5702 3429
rect 5694 2921 5695 2927
rect 5701 2921 5702 2927
rect 5694 2699 5702 2921
rect 5694 2693 5695 2699
rect 5701 2693 5702 2699
rect 5694 2467 5702 2693
rect 5694 2461 5695 2467
rect 5701 2461 5702 2467
rect 5694 2227 5702 2461
rect 5694 2221 5695 2227
rect 5701 2221 5702 2227
rect 5694 2003 5702 2221
rect 5694 1997 5695 2003
rect 5701 1997 5702 2003
rect 5694 1759 5702 1997
rect 5694 1753 5695 1759
rect 5701 1753 5702 1759
rect 5694 1523 5702 1753
rect 5694 1517 5695 1523
rect 5701 1517 5702 1523
rect 5694 1287 5702 1517
rect 5694 1281 5695 1287
rect 5701 1281 5702 1287
rect 5694 1055 5702 1281
rect 5694 1049 5695 1055
rect 5701 1049 5702 1055
rect 5694 823 5702 1049
rect 5694 817 5695 823
rect 5701 817 5702 823
rect 5694 587 5702 817
rect 5694 581 5695 587
rect 5701 581 5702 587
rect 5694 355 5702 581
rect 5694 349 5695 355
rect 5701 349 5702 355
rect 5694 91 5702 349
rect 5694 85 5695 91
rect 5701 85 5702 91
rect 5694 72 5702 85
rect 5706 5571 5714 5760
rect 5706 5565 5707 5571
rect 5713 5565 5714 5571
rect 5706 5279 5714 5565
rect 5706 5273 5707 5279
rect 5713 5273 5714 5279
rect 5706 5015 5714 5273
rect 5706 5009 5707 5015
rect 5713 5009 5714 5015
rect 5706 4767 5714 5009
rect 5706 4761 5707 4767
rect 5713 4761 5714 4767
rect 5706 4535 5714 4761
rect 5706 4529 5707 4535
rect 5713 4529 5714 4535
rect 5706 4299 5714 4529
rect 5706 4293 5707 4299
rect 5713 4293 5714 4299
rect 5706 4039 5714 4293
rect 5706 4033 5707 4039
rect 5713 4033 5714 4039
rect 5706 3555 5714 4033
rect 5706 3549 5707 3555
rect 5713 3549 5714 3555
rect 5706 2811 5714 3549
rect 5706 2805 5707 2811
rect 5713 2805 5714 2811
rect 5706 2583 5714 2805
rect 5706 2577 5707 2583
rect 5713 2577 5714 2583
rect 5706 2351 5714 2577
rect 5706 2345 5707 2351
rect 5713 2345 5714 2351
rect 5706 2115 5714 2345
rect 5706 2109 5707 2115
rect 5713 2109 5714 2115
rect 5706 1879 5714 2109
rect 5706 1873 5707 1879
rect 5713 1873 5714 1879
rect 5706 1635 5714 1873
rect 5706 1629 5707 1635
rect 5713 1629 5714 1635
rect 5706 1399 5714 1629
rect 5706 1393 5707 1399
rect 5713 1393 5714 1399
rect 5706 1171 5714 1393
rect 5706 1165 5707 1171
rect 5713 1165 5714 1171
rect 5706 939 5714 1165
rect 5706 933 5707 939
rect 5713 933 5714 939
rect 5706 699 5714 933
rect 5706 693 5707 699
rect 5713 693 5714 699
rect 5706 475 5714 693
rect 5706 469 5707 475
rect 5713 469 5714 475
rect 5706 203 5714 469
rect 5706 197 5707 203
rect 5713 197 5714 203
rect 5706 72 5714 197
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__271
timestamp 1731220447
transform 1 0 5656 0 -1 5656
box 7 3 12 24
use welltap_svt  __well_tap__270
timestamp 1731220447
transform 1 0 3832 0 -1 5656
box 7 3 12 24
use welltap_svt  __well_tap__269
timestamp 1731220447
transform 1 0 5656 0 1 5480
box 7 3 12 24
use welltap_svt  __well_tap__268
timestamp 1731220447
transform 1 0 3832 0 1 5480
box 7 3 12 24
use welltap_svt  __well_tap__267
timestamp 1731220447
transform 1 0 5656 0 -1 5396
box 7 3 12 24
use welltap_svt  __well_tap__266
timestamp 1731220447
transform 1 0 3832 0 -1 5396
box 7 3 12 24
use welltap_svt  __well_tap__265
timestamp 1731220447
transform 1 0 5656 0 1 5188
box 7 3 12 24
use welltap_svt  __well_tap__264
timestamp 1731220447
transform 1 0 3832 0 1 5188
box 7 3 12 24
use welltap_svt  __well_tap__263
timestamp 1731220447
transform 1 0 5656 0 -1 5116
box 7 3 12 24
use welltap_svt  __well_tap__262
timestamp 1731220447
transform 1 0 3832 0 -1 5116
box 7 3 12 24
use welltap_svt  __well_tap__261
timestamp 1731220447
transform 1 0 5656 0 1 4924
box 7 3 12 24
use welltap_svt  __well_tap__260
timestamp 1731220447
transform 1 0 3832 0 1 4924
box 7 3 12 24
use welltap_svt  __well_tap__259
timestamp 1731220447
transform 1 0 5656 0 -1 4860
box 7 3 12 24
use welltap_svt  __well_tap__258
timestamp 1731220447
transform 1 0 3832 0 -1 4860
box 7 3 12 24
use welltap_svt  __well_tap__257
timestamp 1731220447
transform 1 0 5656 0 1 4676
box 7 3 12 24
use welltap_svt  __well_tap__256
timestamp 1731220447
transform 1 0 3832 0 1 4676
box 7 3 12 24
use welltap_svt  __well_tap__255
timestamp 1731220447
transform 1 0 5656 0 -1 4624
box 7 3 12 24
use welltap_svt  __well_tap__254
timestamp 1731220447
transform 1 0 3832 0 -1 4624
box 7 3 12 24
use welltap_svt  __well_tap__253
timestamp 1731220447
transform 1 0 5656 0 1 4444
box 7 3 12 24
use welltap_svt  __well_tap__252
timestamp 1731220447
transform 1 0 3832 0 1 4444
box 7 3 12 24
use welltap_svt  __well_tap__251
timestamp 1731220447
transform 1 0 5656 0 -1 4396
box 7 3 12 24
use welltap_svt  __well_tap__250
timestamp 1731220447
transform 1 0 3832 0 -1 4396
box 7 3 12 24
use welltap_svt  __well_tap__249
timestamp 1731220447
transform 1 0 5656 0 1 4208
box 7 3 12 24
use welltap_svt  __well_tap__248
timestamp 1731220447
transform 1 0 3832 0 1 4208
box 7 3 12 24
use welltap_svt  __well_tap__247
timestamp 1731220447
transform 1 0 5656 0 -1 4160
box 7 3 12 24
use welltap_svt  __well_tap__246
timestamp 1731220447
transform 1 0 3832 0 -1 4160
box 7 3 12 24
use welltap_svt  __well_tap__245
timestamp 1731220447
transform 1 0 5656 0 1 3948
box 7 3 12 24
use welltap_svt  __well_tap__244
timestamp 1731220447
transform 1 0 3832 0 1 3948
box 7 3 12 24
use welltap_svt  __well_tap__243
timestamp 1731220447
transform 1 0 5656 0 -1 3900
box 7 3 12 24
use welltap_svt  __well_tap__242
timestamp 1731220447
transform 1 0 3832 0 -1 3900
box 7 3 12 24
use welltap_svt  __well_tap__241
timestamp 1731220447
transform 1 0 5656 0 1 3724
box 7 3 12 24
use welltap_svt  __well_tap__240
timestamp 1731220447
transform 1 0 3832 0 1 3724
box 7 3 12 24
use welltap_svt  __well_tap__239
timestamp 1731220447
transform 1 0 5656 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__238
timestamp 1731220447
transform 1 0 3832 0 -1 3652
box 7 3 12 24
use welltap_svt  __well_tap__237
timestamp 1731220447
transform 1 0 5656 0 1 3464
box 7 3 12 24
use welltap_svt  __well_tap__236
timestamp 1731220447
transform 1 0 3832 0 1 3464
box 7 3 12 24
use welltap_svt  __well_tap__235
timestamp 1731220447
transform 1 0 5656 0 -1 3408
box 7 3 12 24
use welltap_svt  __well_tap__234
timestamp 1731220447
transform 1 0 3832 0 -1 3408
box 7 3 12 24
use welltap_svt  __well_tap__233
timestamp 1731220447
transform 1 0 5656 0 1 3216
box 7 3 12 24
use welltap_svt  __well_tap__232
timestamp 1731220447
transform 1 0 3832 0 1 3216
box 7 3 12 24
use welltap_svt  __well_tap__231
timestamp 1731220447
transform 1 0 5656 0 -1 3160
box 7 3 12 24
use welltap_svt  __well_tap__230
timestamp 1731220447
transform 1 0 3832 0 -1 3160
box 7 3 12 24
use welltap_svt  __well_tap__229
timestamp 1731220447
transform 1 0 5656 0 1 2972
box 7 3 12 24
use welltap_svt  __well_tap__228
timestamp 1731220447
transform 1 0 3832 0 1 2972
box 7 3 12 24
use welltap_svt  __well_tap__227
timestamp 1731220447
transform 1 0 5656 0 -1 2900
box 7 3 12 24
use welltap_svt  __well_tap__226
timestamp 1731220447
transform 1 0 3832 0 -1 2900
box 7 3 12 24
use welltap_svt  __well_tap__225
timestamp 1731220447
transform 1 0 5656 0 1 2720
box 7 3 12 24
use welltap_svt  __well_tap__224
timestamp 1731220447
transform 1 0 3832 0 1 2720
box 7 3 12 24
use welltap_svt  __well_tap__223
timestamp 1731220447
transform 1 0 5656 0 -1 2672
box 7 3 12 24
use welltap_svt  __well_tap__222
timestamp 1731220447
transform 1 0 3832 0 -1 2672
box 7 3 12 24
use welltap_svt  __well_tap__221
timestamp 1731220447
transform 1 0 5656 0 1 2492
box 7 3 12 24
use welltap_svt  __well_tap__220
timestamp 1731220447
transform 1 0 3832 0 1 2492
box 7 3 12 24
use welltap_svt  __well_tap__219
timestamp 1731220447
transform 1 0 5656 0 -1 2440
box 7 3 12 24
use welltap_svt  __well_tap__218
timestamp 1731220447
transform 1 0 3832 0 -1 2440
box 7 3 12 24
use welltap_svt  __well_tap__217
timestamp 1731220447
transform 1 0 5656 0 1 2260
box 7 3 12 24
use welltap_svt  __well_tap__216
timestamp 1731220447
transform 1 0 3832 0 1 2260
box 7 3 12 24
use welltap_svt  __well_tap__215
timestamp 1731220447
transform 1 0 5656 0 -1 2200
box 7 3 12 24
use welltap_svt  __well_tap__214
timestamp 1731220447
transform 1 0 3832 0 -1 2200
box 7 3 12 24
use welltap_svt  __well_tap__213
timestamp 1731220447
transform 1 0 5656 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__212
timestamp 1731220447
transform 1 0 3832 0 1 2024
box 7 3 12 24
use welltap_svt  __well_tap__211
timestamp 1731220447
transform 1 0 5656 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__210
timestamp 1731220447
transform 1 0 3832 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__209
timestamp 1731220447
transform 1 0 5656 0 1 1788
box 7 3 12 24
use welltap_svt  __well_tap__208
timestamp 1731220447
transform 1 0 3832 0 1 1788
box 7 3 12 24
use welltap_svt  __well_tap__207
timestamp 1731220447
transform 1 0 5656 0 -1 1732
box 7 3 12 24
use welltap_svt  __well_tap__206
timestamp 1731220447
transform 1 0 3832 0 -1 1732
box 7 3 12 24
use welltap_svt  __well_tap__205
timestamp 1731220447
transform 1 0 5656 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__204
timestamp 1731220447
transform 1 0 3832 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__203
timestamp 1731220447
transform 1 0 5656 0 -1 1496
box 7 3 12 24
use welltap_svt  __well_tap__202
timestamp 1731220447
transform 1 0 3832 0 -1 1496
box 7 3 12 24
use welltap_svt  __well_tap__201
timestamp 1731220447
transform 1 0 5656 0 1 1308
box 7 3 12 24
use welltap_svt  __well_tap__200
timestamp 1731220447
transform 1 0 3832 0 1 1308
box 7 3 12 24
use welltap_svt  __well_tap__199
timestamp 1731220447
transform 1 0 5656 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220447
transform 1 0 3832 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220447
transform 1 0 5656 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220447
transform 1 0 3832 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220447
transform 1 0 5656 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220447
transform 1 0 3832 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220447
transform 1 0 5656 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220447
transform 1 0 3832 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220447
transform 1 0 5656 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220447
transform 1 0 3832 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220447
transform 1 0 5656 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220447
transform 1 0 3832 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220447
transform 1 0 5656 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220447
transform 1 0 3832 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220447
transform 1 0 5656 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220447
transform 1 0 3832 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220447
transform 1 0 5656 0 -1 328
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220447
transform 1 0 3832 0 -1 328
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220447
transform 1 0 5656 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220447
transform 1 0 3832 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220447
transform 1 0 3792 0 -1 5732
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220447
transform 1 0 1968 0 -1 5732
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220447
transform 1 0 3792 0 1 5556
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220447
transform 1 0 1968 0 1 5556
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220447
transform 1 0 3792 0 -1 5508
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220447
transform 1 0 1968 0 -1 5508
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220447
transform 1 0 3792 0 1 5284
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220447
transform 1 0 1968 0 1 5284
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220447
transform 1 0 3792 0 -1 5236
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220447
transform 1 0 1968 0 -1 5236
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220447
transform 1 0 3792 0 1 5052
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220447
transform 1 0 1968 0 1 5052
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220447
transform 1 0 3792 0 -1 4980
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220447
transform 1 0 1968 0 -1 4980
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220447
transform 1 0 3792 0 1 4796
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220447
transform 1 0 1968 0 1 4796
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220447
transform 1 0 3792 0 -1 4700
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220447
transform 1 0 1968 0 -1 4700
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220447
transform 1 0 3792 0 1 4520
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220447
transform 1 0 1968 0 1 4520
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220447
transform 1 0 3792 0 -1 4464
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220447
transform 1 0 1968 0 -1 4464
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220447
transform 1 0 3792 0 1 4272
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220447
transform 1 0 1968 0 1 4272
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220447
transform 1 0 3792 0 -1 4196
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220447
transform 1 0 1968 0 -1 4196
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220447
transform 1 0 3792 0 1 3984
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220447
transform 1 0 1968 0 1 3984
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220447
transform 1 0 3792 0 -1 3908
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220447
transform 1 0 1968 0 -1 3908
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220447
transform 1 0 3792 0 1 3724
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220447
transform 1 0 1968 0 1 3724
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220447
transform 1 0 3792 0 -1 3668
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220447
transform 1 0 1968 0 -1 3668
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220447
transform 1 0 3792 0 1 3476
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220447
transform 1 0 1968 0 1 3476
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220447
transform 1 0 3792 0 -1 3392
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220447
transform 1 0 1968 0 -1 3392
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220447
transform 1 0 3792 0 1 3216
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220447
transform 1 0 1968 0 1 3216
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220447
transform 1 0 3792 0 -1 3160
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220447
transform 1 0 1968 0 -1 3160
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220447
transform 1 0 3792 0 1 2972
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220447
transform 1 0 1968 0 1 2972
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220447
transform 1 0 3792 0 -1 2924
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220447
transform 1 0 1968 0 -1 2924
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220447
transform 1 0 3792 0 1 2692
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220447
transform 1 0 1968 0 1 2692
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220447
transform 1 0 3792 0 -1 2620
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220447
transform 1 0 1968 0 -1 2620
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220447
transform 1 0 3792 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220447
transform 1 0 1968 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220447
transform 1 0 3792 0 -1 2388
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220447
transform 1 0 1968 0 -1 2388
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220447
transform 1 0 3792 0 1 2208
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220447
transform 1 0 1968 0 1 2208
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220447
transform 1 0 3792 0 -1 2160
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220447
transform 1 0 1968 0 -1 2160
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220447
transform 1 0 3792 0 1 1968
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220447
transform 1 0 1968 0 1 1968
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220447
transform 1 0 3792 0 -1 1912
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220447
transform 1 0 1968 0 -1 1912
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220447
transform 1 0 3792 0 1 1728
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220447
transform 1 0 1968 0 1 1728
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220447
transform 1 0 3792 0 -1 1680
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220447
transform 1 0 1968 0 -1 1680
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220447
transform 1 0 3792 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220447
transform 1 0 1968 0 1 1504
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220447
transform 1 0 3792 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220447
transform 1 0 1968 0 -1 1456
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220447
transform 1 0 3792 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220447
transform 1 0 1968 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220447
transform 1 0 3792 0 -1 1168
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220447
transform 1 0 1968 0 -1 1168
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220447
transform 1 0 3792 0 1 992
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220447
transform 1 0 1968 0 1 992
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220447
transform 1 0 3792 0 -1 940
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220447
transform 1 0 1968 0 -1 940
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220447
transform 1 0 3792 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220447
transform 1 0 1968 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220447
transform 1 0 3792 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220447
transform 1 0 1968 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220447
transform 1 0 3792 0 1 360
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220447
transform 1 0 1968 0 1 360
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220447
transform 1 0 3792 0 -1 308
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220447
transform 1 0 1968 0 -1 308
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220447
transform 1 0 3792 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220447
transform 1 0 1968 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220447
transform 1 0 1928 0 -1 5692
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220447
transform 1 0 104 0 -1 5692
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220447
transform 1 0 1928 0 1 5488
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220447
transform 1 0 104 0 1 5488
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220447
transform 1 0 1928 0 -1 5432
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220447
transform 1 0 104 0 -1 5432
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220447
transform 1 0 1928 0 1 5232
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220447
transform 1 0 104 0 1 5232
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220447
transform 1 0 1928 0 -1 5176
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220447
transform 1 0 104 0 -1 5176
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220447
transform 1 0 1928 0 1 4980
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220447
transform 1 0 104 0 1 4980
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220447
transform 1 0 1928 0 -1 4920
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220447
transform 1 0 104 0 -1 4920
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220447
transform 1 0 1928 0 1 4744
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220447
transform 1 0 104 0 1 4744
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220447
transform 1 0 1928 0 -1 4676
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220447
transform 1 0 104 0 -1 4676
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220447
transform 1 0 1928 0 1 4484
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220447
transform 1 0 104 0 1 4484
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220447
transform 1 0 1928 0 -1 4420
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220447
transform 1 0 104 0 -1 4420
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220447
transform 1 0 1928 0 1 4244
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220447
transform 1 0 104 0 1 4244
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220447
transform 1 0 1928 0 -1 4184
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220447
transform 1 0 104 0 -1 4184
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220447
transform 1 0 1928 0 1 4008
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220447
transform 1 0 104 0 1 4008
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220447
transform 1 0 1928 0 -1 3956
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220447
transform 1 0 104 0 -1 3956
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220447
transform 1 0 1928 0 1 3776
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220447
transform 1 0 104 0 1 3776
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220447
transform 1 0 1928 0 -1 3724
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220447
transform 1 0 104 0 -1 3724
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220447
transform 1 0 1928 0 1 3540
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220447
transform 1 0 104 0 1 3540
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220447
transform 1 0 1928 0 -1 3480
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220447
transform 1 0 104 0 -1 3480
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220447
transform 1 0 1928 0 1 3296
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220447
transform 1 0 104 0 1 3296
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220447
transform 1 0 1928 0 -1 3244
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220447
transform 1 0 104 0 -1 3244
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220447
transform 1 0 1928 0 1 3064
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220447
transform 1 0 104 0 1 3064
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220447
transform 1 0 1928 0 -1 3000
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220447
transform 1 0 104 0 -1 3000
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220447
transform 1 0 1928 0 1 2816
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220447
transform 1 0 104 0 1 2816
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220447
transform 1 0 1928 0 -1 2760
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220447
transform 1 0 104 0 -1 2760
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220447
transform 1 0 1928 0 1 2580
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220447
transform 1 0 104 0 1 2580
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220447
transform 1 0 1928 0 -1 2532
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220447
transform 1 0 104 0 -1 2532
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220447
transform 1 0 1928 0 1 2336
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220447
transform 1 0 104 0 1 2336
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220447
transform 1 0 1928 0 -1 2284
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220447
transform 1 0 104 0 -1 2284
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220447
transform 1 0 1928 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220447
transform 1 0 104 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220447
transform 1 0 1928 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220447
transform 1 0 104 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220447
transform 1 0 1928 0 1 1836
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220447
transform 1 0 104 0 1 1836
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220447
transform 1 0 1928 0 -1 1776
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220447
transform 1 0 104 0 -1 1776
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220447
transform 1 0 1928 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220447
transform 1 0 104 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220447
transform 1 0 1928 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220447
transform 1 0 104 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220447
transform 1 0 1928 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220447
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220447
transform 1 0 1928 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220447
transform 1 0 104 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220447
transform 1 0 1928 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220447
transform 1 0 104 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220447
transform 1 0 1928 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220447
transform 1 0 104 0 -1 1040
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220447
transform 1 0 1928 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220447
transform 1 0 104 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220447
transform 1 0 1928 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220447
transform 1 0 104 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220447
transform 1 0 1928 0 1 624
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220447
transform 1 0 104 0 1 624
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220447
transform 1 0 1928 0 -1 576
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220447
transform 1 0 104 0 -1 576
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220447
transform 1 0 1928 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220447
transform 1 0 104 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220447
transform 1 0 1928 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220447
transform 1 0 104 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220447
transform 1 0 1928 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220447
transform 1 0 104 0 1 120
box 7 3 12 24
use _0_0std_0_0cells_0_0FAX1  tst_5999_6
timestamp 1731220447
transform 1 0 5376 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5998_6
timestamp 1731220447
transform 1 0 5512 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5997_6
timestamp 1731220447
transform 1 0 5512 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5996_6
timestamp 1731220447
transform 1 0 5504 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5995_6
timestamp 1731220447
transform 1 0 5456 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5994_6
timestamp 1731220447
transform 1 0 5416 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5993_6
timestamp 1731220447
transform 1 0 5224 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5992_6
timestamp 1731220447
transform 1 0 5200 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5991_6
timestamp 1731220447
transform 1 0 5368 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5990_6
timestamp 1731220447
transform 1 0 5240 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5989_6
timestamp 1731220447
transform 1 0 5104 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5988_6
timestamp 1731220447
transform 1 0 4968 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5987_6
timestamp 1731220447
transform 1 0 4832 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5986_6
timestamp 1731220447
transform 1 0 4696 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5985_6
timestamp 1731220447
transform 1 0 4560 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5984_6
timestamp 1731220447
transform 1 0 4424 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5983_6
timestamp 1731220447
transform 1 0 4288 0 1 88
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5982_6
timestamp 1731220447
transform 1 0 4696 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5981_6
timestamp 1731220447
transform 1 0 4864 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5980_6
timestamp 1731220447
transform 1 0 5032 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5979_6
timestamp 1731220447
transform 1 0 4944 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5978_6
timestamp 1731220447
transform 1 0 4672 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5977_6
timestamp 1731220447
transform 1 0 4392 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5976_6
timestamp 1731220447
transform 1 0 4112 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5975_6
timestamp 1731220447
transform 1 0 5032 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5974_6
timestamp 1731220447
transform 1 0 5224 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5973_6
timestamp 1731220447
transform 1 0 5160 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5972_6
timestamp 1731220447
transform 1 0 4864 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5971_6
timestamp 1731220447
transform 1 0 4176 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5970_6
timestamp 1731220447
transform 1 0 3928 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5969_6
timestamp 1731220447
transform 1 0 3992 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5968_6
timestamp 1731220447
transform 1 0 4144 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5967_6
timestamp 1731220447
transform 1 0 4536 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5966_6
timestamp 1731220447
transform 1 0 4848 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5965_6
timestamp 1731220447
transform 1 0 4680 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5964_6
timestamp 1731220447
transform 1 0 4592 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5963_6
timestamp 1731220447
transform 1 0 4352 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5962_6
timestamp 1731220447
transform 1 0 4464 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5961_6
timestamp 1731220447
transform 1 0 4784 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5960_6
timestamp 1731220447
transform 1 0 5120 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5959_6
timestamp 1731220447
transform 1 0 5040 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5958_6
timestamp 1731220447
transform 1 0 4800 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5957_6
timestamp 1731220447
transform 1 0 4568 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5956_6
timestamp 1731220447
transform 1 0 4352 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5955_6
timestamp 1731220447
transform 1 0 4776 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5954_6
timestamp 1731220447
transform 1 0 4912 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5953_6
timestamp 1731220447
transform 1 0 5048 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5952_6
timestamp 1731220447
transform 1 0 5184 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5951_6
timestamp 1731220447
transform 1 0 5376 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5950_6
timestamp 1731220447
transform 1 0 5224 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5949_6
timestamp 1731220447
transform 1 0 5080 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5948_6
timestamp 1731220447
transform 1 0 4944 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5947_6
timestamp 1731220447
transform 1 0 4808 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5946_6
timestamp 1731220447
transform 1 0 5088 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5945_6
timestamp 1731220447
transform 1 0 4872 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5944_6
timestamp 1731220447
transform 1 0 4672 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5943_6
timestamp 1731220447
transform 1 0 4480 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5942_6
timestamp 1731220447
transform 1 0 5192 0 1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5941_6
timestamp 1731220447
transform 1 0 4888 0 1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5940_6
timestamp 1731220447
transform 1 0 4608 0 1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5939_6
timestamp 1731220447
transform 1 0 4360 0 1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5938_6
timestamp 1731220447
transform 1 0 4448 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5937_6
timestamp 1731220447
transform 1 0 4664 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5936_6
timestamp 1731220447
transform 1 0 5160 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5935_6
timestamp 1731220447
transform 1 0 4904 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5934_6
timestamp 1731220447
transform 1 0 4904 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5933_6
timestamp 1731220447
transform 1 0 4264 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5932_6
timestamp 1731220447
transform 1 0 4144 0 1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5931_6
timestamp 1731220447
transform 1 0 3992 0 1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5930_6
timestamp 1731220447
transform 1 0 4304 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5929_6
timestamp 1731220447
transform 1 0 4136 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5928_6
timestamp 1731220447
transform 1 0 3992 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5927_6
timestamp 1731220447
transform 1 0 3856 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5926_6
timestamp 1731220447
transform 1 0 3856 0 1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5925_6
timestamp 1731220447
transform 1 0 3648 0 -1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5924_6
timestamp 1731220447
transform 1 0 3856 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5923_6
timestamp 1731220447
transform 1 0 4128 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5922_6
timestamp 1731220447
transform 1 0 3992 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5921_6
timestamp 1731220447
transform 1 0 3904 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5920_6
timestamp 1731220447
transform 1 0 4120 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5919_6
timestamp 1731220447
transform 1 0 4360 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5918_6
timestamp 1731220447
transform 1 0 4624 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5917_6
timestamp 1731220447
transform 1 0 4568 0 -1 1756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5916_6
timestamp 1731220447
transform 1 0 4352 0 -1 1756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5915_6
timestamp 1731220447
transform 1 0 5040 0 -1 1756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5914_6
timestamp 1731220447
transform 1 0 4800 0 -1 1756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5913_6
timestamp 1731220447
transform 1 0 4720 0 1 1764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5912_6
timestamp 1731220447
transform 1 0 4536 0 1 1764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5911_6
timestamp 1731220447
transform 1 0 5112 0 1 1764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5910_6
timestamp 1731220447
transform 1 0 4912 0 1 1764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5909_6
timestamp 1731220447
transform 1 0 4712 0 -1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5908_6
timestamp 1731220447
transform 1 0 4432 0 -1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5907_6
timestamp 1731220447
transform 1 0 4136 0 -1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5906_6
timestamp 1731220447
transform 1 0 4976 0 -1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5905_6
timestamp 1731220447
transform 1 0 4944 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5904_6
timestamp 1731220447
transform 1 0 4752 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5903_6
timestamp 1731220447
transform 1 0 4544 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5902_6
timestamp 1731220447
transform 1 0 5200 0 -1 2224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5901_6
timestamp 1731220447
transform 1 0 5136 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5900_6
timestamp 1731220447
transform 1 0 5320 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5899_6
timestamp 1731220447
transform 1 0 5240 0 -1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5898_6
timestamp 1731220447
transform 1 0 5320 0 1 1764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5897_6
timestamp 1731220447
transform 1 0 5288 0 -1 1756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5896_6
timestamp 1731220447
transform 1 0 5192 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5895_6
timestamp 1731220447
transform 1 0 5312 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5894_6
timestamp 1731220447
transform 1 0 5320 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5893_6
timestamp 1731220447
transform 1 0 5288 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5892_6
timestamp 1731220447
transform 1 0 5456 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5891_6
timestamp 1731220447
transform 1 0 5456 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5890_6
timestamp 1731220447
transform 1 0 5512 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5889_6
timestamp 1731220447
transform 1 0 5512 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5888_6
timestamp 1731220447
transform 1 0 5512 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5887_6
timestamp 1731220447
transform 1 0 5496 0 1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5886_6
timestamp 1731220447
transform 1 0 5416 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5885_6
timestamp 1731220447
transform 1 0 5488 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5884_6
timestamp 1731220447
transform 1 0 5512 0 -1 1756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5883_6
timestamp 1731220447
transform 1 0 5512 0 1 1764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5882_6
timestamp 1731220447
transform 1 0 5512 0 -1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5881_6
timestamp 1731220447
transform 1 0 5512 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5880_6
timestamp 1731220447
transform 1 0 5456 0 -1 2224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5879_6
timestamp 1731220447
transform 1 0 5416 0 1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5878_6
timestamp 1731220447
transform 1 0 5352 0 -1 2464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5877_6
timestamp 1731220447
transform 1 0 5168 0 -1 2464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5876_6
timestamp 1731220447
transform 1 0 4992 0 -1 2464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5875_6
timestamp 1731220447
transform 1 0 5264 0 1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5874_6
timestamp 1731220447
transform 1 0 5112 0 1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5873_6
timestamp 1731220447
transform 1 0 4944 0 -1 2224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5872_6
timestamp 1731220447
transform 1 0 4688 0 -1 2224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5871_6
timestamp 1731220447
transform 1 0 4424 0 -1 2224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5870_6
timestamp 1731220447
transform 1 0 4136 0 -1 2224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5869_6
timestamp 1731220447
transform 1 0 4960 0 1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5868_6
timestamp 1731220447
transform 1 0 4816 0 1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5867_6
timestamp 1731220447
transform 1 0 4672 0 1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5866_6
timestamp 1731220447
transform 1 0 4632 0 -1 2464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5865_6
timestamp 1731220447
transform 1 0 4816 0 -1 2464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5864_6
timestamp 1731220447
transform 1 0 5256 0 1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5863_6
timestamp 1731220447
transform 1 0 4976 0 1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5862_6
timestamp 1731220447
transform 1 0 4712 0 1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5861_6
timestamp 1731220447
transform 1 0 4472 0 1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5860_6
timestamp 1731220447
transform 1 0 4256 0 1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5859_6
timestamp 1731220447
transform 1 0 5200 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5858_6
timestamp 1731220447
transform 1 0 4864 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5857_6
timestamp 1731220447
transform 1 0 4552 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5856_6
timestamp 1731220447
transform 1 0 4272 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5855_6
timestamp 1731220447
transform 1 0 4024 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5854_6
timestamp 1731220447
transform 1 0 4808 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5853_6
timestamp 1731220447
transform 1 0 4672 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5852_6
timestamp 1731220447
transform 1 0 4536 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5851_6
timestamp 1731220447
transform 1 0 4400 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5850_6
timestamp 1731220447
transform 1 0 4264 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5849_6
timestamp 1731220447
transform 1 0 4128 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5848_6
timestamp 1731220447
transform 1 0 3992 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5847_6
timestamp 1731220447
transform 1 0 3856 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5846_6
timestamp 1731220447
transform 1 0 4016 0 -1 2924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5845_6
timestamp 1731220447
transform 1 0 4264 0 -1 2924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5844_6
timestamp 1731220447
transform 1 0 4552 0 -1 2924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5843_6
timestamp 1731220447
transform 1 0 4864 0 -1 2924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5842_6
timestamp 1731220447
transform 1 0 5200 0 -1 2924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5841_6
timestamp 1731220447
transform 1 0 5160 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5840_6
timestamp 1731220447
transform 1 0 4976 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5839_6
timestamp 1731220447
transform 1 0 4800 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5838_6
timestamp 1731220447
transform 1 0 4632 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5837_6
timestamp 1731220447
transform 1 0 4480 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5836_6
timestamp 1731220447
transform 1 0 4832 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5835_6
timestamp 1731220447
transform 1 0 4968 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5834_6
timestamp 1731220447
transform 1 0 5104 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5833_6
timestamp 1731220447
transform 1 0 5376 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5832_6
timestamp 1731220447
transform 1 0 5240 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5831_6
timestamp 1731220447
transform 1 0 5232 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5830_6
timestamp 1731220447
transform 1 0 5096 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5829_6
timestamp 1731220447
transform 1 0 4960 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5828_6
timestamp 1731220447
transform 1 0 4824 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5827_6
timestamp 1731220447
transform 1 0 4688 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5826_6
timestamp 1731220447
transform 1 0 5120 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5825_6
timestamp 1731220447
transform 1 0 4920 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5824_6
timestamp 1731220447
transform 1 0 4728 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5823_6
timestamp 1731220447
transform 1 0 4552 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5822_6
timestamp 1731220447
transform 1 0 4400 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5821_6
timestamp 1731220447
transform 1 0 5312 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5820_6
timestamp 1731220447
transform 1 0 5096 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5819_6
timestamp 1731220447
transform 1 0 4888 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5818_6
timestamp 1731220447
transform 1 0 4696 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5817_6
timestamp 1731220447
transform 1 0 4536 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5816_6
timestamp 1731220447
transform 1 0 4448 0 -1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5815_6
timestamp 1731220447
transform 1 0 4216 0 -1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5814_6
timestamp 1731220447
transform 1 0 4016 0 -1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5813_6
timestamp 1731220447
transform 1 0 4968 0 -1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5812_6
timestamp 1731220447
transform 1 0 4696 0 -1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5811_6
timestamp 1731220447
transform 1 0 4616 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5810_6
timestamp 1731220447
transform 1 0 4408 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5809_6
timestamp 1731220447
transform 1 0 5064 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5808_6
timestamp 1731220447
transform 1 0 4832 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5807_6
timestamp 1731220447
transform 1 0 4816 0 -1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5806_6
timestamp 1731220447
transform 1 0 4656 0 -1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5805_6
timestamp 1731220447
transform 1 0 4984 0 -1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5804_6
timestamp 1731220447
transform 1 0 5160 0 -1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5803_6
timestamp 1731220447
transform 1 0 5072 0 1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5802_6
timestamp 1731220447
transform 1 0 4936 0 1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5801_6
timestamp 1731220447
transform 1 0 5208 0 1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5800_6
timestamp 1731220447
transform 1 0 5344 0 1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5799_6
timestamp 1731220447
transform 1 0 5344 0 -1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5798_6
timestamp 1731220447
transform 1 0 5296 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5797_6
timestamp 1731220447
transform 1 0 5248 0 -1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5796_6
timestamp 1731220447
transform 1 0 5328 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5795_6
timestamp 1731220447
transform 1 0 5344 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5794_6
timestamp 1731220447
transform 1 0 5512 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5793_6
timestamp 1731220447
transform 1 0 5512 0 -1 2464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5792_6
timestamp 1731220447
transform 1 0 5512 0 1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5791_6
timestamp 1731220447
transform 1 0 5512 0 -1 2924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5790_6
timestamp 1731220447
transform 1 0 5512 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5789_6
timestamp 1731220447
transform 1 0 5512 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5788_6
timestamp 1731220447
transform 1 0 5512 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5787_6
timestamp 1731220447
transform 1 0 5512 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5786_6
timestamp 1731220447
transform 1 0 5512 0 -1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5785_6
timestamp 1731220447
transform 1 0 5512 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5784_6
timestamp 1731220447
transform 1 0 5512 0 -1 3924
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5783_6
timestamp 1731220447
transform 1 0 5512 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5782_6
timestamp 1731220447
transform 1 0 5512 0 1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5781_6
timestamp 1731220447
transform 1 0 5512 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5780_6
timestamp 1731220447
transform 1 0 5512 0 1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5779_6
timestamp 1731220447
transform 1 0 5504 0 1 4652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5778_6
timestamp 1731220447
transform 1 0 5488 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5777_6
timestamp 1731220447
transform 1 0 5512 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5776_6
timestamp 1731220447
transform 1 0 5336 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5775_6
timestamp 1731220447
transform 1 0 5408 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5774_6
timestamp 1731220447
transform 1 0 5192 0 1 5164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5773_6
timestamp 1731220447
transform 1 0 5416 0 1 5164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5772_6
timestamp 1731220447
transform 1 0 5368 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5771_6
timestamp 1731220447
transform 1 0 5144 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5770_6
timestamp 1731220447
transform 1 0 4920 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5769_6
timestamp 1731220447
transform 1 0 4792 0 1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5768_6
timestamp 1731220447
transform 1 0 5192 0 1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5767_6
timestamp 1731220447
transform 1 0 4992 0 1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5766_6
timestamp 1731220447
transform 1 0 4984 0 -1 5680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5765_6
timestamp 1731220447
transform 1 0 4848 0 -1 5680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5764_6
timestamp 1731220447
transform 1 0 4712 0 -1 5680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5763_6
timestamp 1731220447
transform 1 0 4576 0 -1 5680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5762_6
timestamp 1731220447
transform 1 0 4440 0 -1 5680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5761_6
timestamp 1731220447
transform 1 0 4304 0 -1 5680
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5760_6
timestamp 1731220447
transform 1 0 4208 0 1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5759_6
timestamp 1731220447
transform 1 0 4592 0 1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5758_6
timestamp 1731220447
transform 1 0 4400 0 1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5757_6
timestamp 1731220447
transform 1 0 4272 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5756_6
timestamp 1731220447
transform 1 0 4704 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5755_6
timestamp 1731220447
transform 1 0 4488 0 -1 5420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5754_6
timestamp 1731220447
transform 1 0 4368 0 1 5164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5753_6
timestamp 1731220447
transform 1 0 4976 0 1 5164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5752_6
timestamp 1731220447
transform 1 0 4768 0 1 5164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5751_6
timestamp 1731220447
transform 1 0 4560 0 1 5164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5750_6
timestamp 1731220447
transform 1 0 4504 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5749_6
timestamp 1731220447
transform 1 0 4280 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5748_6
timestamp 1731220447
transform 1 0 4728 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5747_6
timestamp 1731220447
transform 1 0 4952 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5746_6
timestamp 1731220447
transform 1 0 5176 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5745_6
timestamp 1731220447
transform 1 0 5152 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5744_6
timestamp 1731220447
transform 1 0 4968 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5743_6
timestamp 1731220447
transform 1 0 4784 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5742_6
timestamp 1731220447
transform 1 0 4928 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5741_6
timestamp 1731220447
transform 1 0 5208 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5740_6
timestamp 1731220447
transform 1 0 5224 0 1 4652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5739_6
timestamp 1731220447
transform 1 0 4952 0 1 4652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5738_6
timestamp 1731220447
transform 1 0 4984 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5737_6
timestamp 1731220447
transform 1 0 5272 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5736_6
timestamp 1731220447
transform 1 0 5160 0 1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5735_6
timestamp 1731220447
transform 1 0 4952 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5734_6
timestamp 1731220447
transform 1 0 5232 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5733_6
timestamp 1731220447
transform 1 0 5104 0 1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5732_6
timestamp 1731220447
transform 1 0 5304 0 1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5731_6
timestamp 1731220447
transform 1 0 5328 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5730_6
timestamp 1731220447
transform 1 0 5136 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5729_6
timestamp 1731220447
transform 1 0 4952 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5728_6
timestamp 1731220447
transform 1 0 4784 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5727_6
timestamp 1731220447
transform 1 0 4624 0 -1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5726_6
timestamp 1731220447
transform 1 0 4568 0 1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5725_6
timestamp 1731220447
transform 1 0 4912 0 1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5724_6
timestamp 1731220447
transform 1 0 4736 0 1 4184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5723_6
timestamp 1731220447
transform 1 0 4672 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5722_6
timestamp 1731220447
transform 1 0 4392 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5721_6
timestamp 1731220447
transform 1 0 4112 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5720_6
timestamp 1731220447
transform 1 0 4152 0 1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5719_6
timestamp 1731220447
transform 1 0 4480 0 1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5718_6
timestamp 1731220447
transform 1 0 4816 0 1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5717_6
timestamp 1731220447
transform 1 0 4704 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5716_6
timestamp 1731220447
transform 1 0 4424 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5715_6
timestamp 1731220447
transform 1 0 4144 0 -1 4648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5714_6
timestamp 1731220447
transform 1 0 4688 0 1 4652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5713_6
timestamp 1731220447
transform 1 0 4432 0 1 4652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5712_6
timestamp 1731220447
transform 1 0 4176 0 1 4652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5711_6
timestamp 1731220447
transform 1 0 3936 0 1 4652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5710_6
timestamp 1731220447
transform 1 0 3912 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5709_6
timestamp 1731220447
transform 1 0 4152 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5708_6
timestamp 1731220447
transform 1 0 4400 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5707_6
timestamp 1731220447
transform 1 0 4656 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5706_6
timestamp 1731220447
transform 1 0 4608 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5705_6
timestamp 1731220447
transform 1 0 4440 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5704_6
timestamp 1731220447
transform 1 0 4280 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5703_6
timestamp 1731220447
transform 1 0 4128 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5702_6
timestamp 1731220447
transform 1 0 3992 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5701_6
timestamp 1731220447
transform 1 0 3856 0 1 4900
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5700_6
timestamp 1731220447
transform 1 0 4056 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5699_6
timestamp 1731220447
transform 1 0 3856 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5698_6
timestamp 1731220447
transform 1 0 3648 0 1 5028
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5697_6
timestamp 1731220447
transform 1 0 3648 0 -1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5696_6
timestamp 1731220447
transform 1 0 3504 0 -1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5695_6
timestamp 1731220447
transform 1 0 3336 0 -1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5694_6
timestamp 1731220447
transform 1 0 3640 0 1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5693_6
timestamp 1731220447
transform 1 0 3472 0 1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5692_6
timestamp 1731220447
transform 1 0 3304 0 1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5691_6
timestamp 1731220447
transform 1 0 3136 0 1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5690_6
timestamp 1731220447
transform 1 0 3008 0 -1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5689_6
timestamp 1731220447
transform 1 0 3176 0 -1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5688_6
timestamp 1731220447
transform 1 0 3416 0 1 5028
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5687_6
timestamp 1731220447
transform 1 0 3160 0 1 5028
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5686_6
timestamp 1731220447
transform 1 0 3152 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5685_6
timestamp 1731220447
transform 1 0 2936 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5684_6
timestamp 1731220447
transform 1 0 2664 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5683_6
timestamp 1731220447
transform 1 0 2320 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5682_6
timestamp 1731220447
transform 1 0 3016 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5681_6
timestamp 1731220447
transform 1 0 3368 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5680_6
timestamp 1731220447
transform 1 0 3224 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5679_6
timestamp 1731220447
transform 1 0 3048 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5678_6
timestamp 1731220447
transform 1 0 3408 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5677_6
timestamp 1731220447
transform 1 0 3592 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5676_6
timestamp 1731220447
transform 1 0 3488 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5675_6
timestamp 1731220447
transform 1 0 3312 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5674_6
timestamp 1731220447
transform 1 0 3136 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5673_6
timestamp 1731220447
transform 1 0 3648 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5672_6
timestamp 1731220447
transform 1 0 3856 0 1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5671_6
timestamp 1731220447
transform 1 0 3856 0 -1 4420
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5670_6
timestamp 1731220447
transform 1 0 3648 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5669_6
timestamp 1731220447
transform 1 0 3648 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5668_6
timestamp 1731220447
transform 1 0 3512 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5667_6
timestamp 1731220447
transform 1 0 3488 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5666_6
timestamp 1731220447
transform 1 0 3640 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5665_6
timestamp 1731220447
transform 1 0 3560 0 -1 3932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5664_6
timestamp 1731220447
transform 1 0 3384 0 -1 3932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5663_6
timestamp 1731220447
transform 1 0 3392 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5662_6
timestamp 1731220447
transform 1 0 3552 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5661_6
timestamp 1731220447
transform 1 0 3464 0 -1 3692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5660_6
timestamp 1731220447
transform 1 0 3256 0 -1 3692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5659_6
timestamp 1731220447
transform 1 0 3048 0 -1 3692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5658_6
timestamp 1731220447
transform 1 0 3648 0 -1 3692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5657_6
timestamp 1731220447
transform 1 0 3856 0 -1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5656_6
timestamp 1731220447
transform 1 0 3856 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5655_6
timestamp 1731220447
transform 1 0 3992 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5654_6
timestamp 1731220447
transform 1 0 4128 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5653_6
timestamp 1731220447
transform 1 0 4400 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5652_6
timestamp 1731220447
transform 1 0 4264 0 1 3440
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5651_6
timestamp 1731220447
transform 1 0 4264 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5650_6
timestamp 1731220447
transform 1 0 4128 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5649_6
timestamp 1731220447
transform 1 0 3992 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5648_6
timestamp 1731220447
transform 1 0 3856 0 -1 3432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5647_6
timestamp 1731220447
transform 1 0 3648 0 -1 3416
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5646_6
timestamp 1731220447
transform 1 0 3648 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5645_6
timestamp 1731220447
transform 1 0 3480 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5644_6
timestamp 1731220447
transform 1 0 3288 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5643_6
timestamp 1731220447
transform 1 0 3096 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5642_6
timestamp 1731220447
transform 1 0 2896 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5641_6
timestamp 1731220447
transform 1 0 3568 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5640_6
timestamp 1731220447
transform 1 0 3384 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5639_6
timestamp 1731220447
transform 1 0 3200 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5638_6
timestamp 1731220447
transform 1 0 3024 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5637_6
timestamp 1731220447
transform 1 0 2840 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5636_6
timestamp 1731220447
transform 1 0 3288 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5635_6
timestamp 1731220447
transform 1 0 3136 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5634_6
timestamp 1731220447
transform 1 0 2984 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5633_6
timestamp 1731220447
transform 1 0 2832 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5632_6
timestamp 1731220447
transform 1 0 2680 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5631_6
timestamp 1731220447
transform 1 0 2560 0 -1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5630_6
timestamp 1731220447
transform 1 0 2264 0 -1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5629_6
timestamp 1731220447
transform 1 0 2856 0 -1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5628_6
timestamp 1731220447
transform 1 0 3152 0 -1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5627_6
timestamp 1731220447
transform 1 0 3056 0 1 2668
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5626_6
timestamp 1731220447
transform 1 0 3192 0 1 2668
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5625_6
timestamp 1731220447
transform 1 0 3328 0 1 2668
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5624_6
timestamp 1731220447
transform 1 0 3240 0 -1 2644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5623_6
timestamp 1731220447
transform 1 0 3104 0 -1 2644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5622_6
timestamp 1731220447
transform 1 0 3376 0 -1 2644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5621_6
timestamp 1731220447
transform 1 0 3512 0 -1 2644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5620_6
timestamp 1731220447
transform 1 0 3648 0 -1 2644
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5619_6
timestamp 1731220447
transform 1 0 3576 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5618_6
timestamp 1731220447
transform 1 0 3360 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5617_6
timestamp 1731220447
transform 1 0 3152 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5616_6
timestamp 1731220447
transform 1 0 2936 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5615_6
timestamp 1731220447
transform 1 0 2712 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5614_6
timestamp 1731220447
transform 1 0 3280 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5613_6
timestamp 1731220447
transform 1 0 3128 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5612_6
timestamp 1731220447
transform 1 0 2976 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5611_6
timestamp 1731220447
transform 1 0 2824 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5610_6
timestamp 1731220447
transform 1 0 2680 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5609_6
timestamp 1731220447
transform 1 0 3128 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5608_6
timestamp 1731220447
transform 1 0 2992 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5607_6
timestamp 1731220447
transform 1 0 2856 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5606_6
timestamp 1731220447
transform 1 0 2720 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5605_6
timestamp 1731220447
transform 1 0 2584 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5604_6
timestamp 1731220447
transform 1 0 2936 0 -1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5603_6
timestamp 1731220447
transform 1 0 2696 0 -1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5602_6
timestamp 1731220447
transform 1 0 2456 0 -1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5601_6
timestamp 1731220447
transform 1 0 2208 0 -1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5600_6
timestamp 1731220447
transform 1 0 2448 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5599_6
timestamp 1731220447
transform 1 0 2312 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5598_6
timestamp 1731220447
transform 1 0 2176 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5597_6
timestamp 1731220447
transform 1 0 2040 0 1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5596_6
timestamp 1731220447
transform 1 0 2536 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5595_6
timestamp 1731220447
transform 1 0 2400 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5594_6
timestamp 1731220447
transform 1 0 2264 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5593_6
timestamp 1731220447
transform 1 0 2128 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5592_6
timestamp 1731220447
transform 1 0 1992 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5591_6
timestamp 1731220447
transform 1 0 2480 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5590_6
timestamp 1731220447
transform 1 0 2232 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5589_6
timestamp 1731220447
transform 1 0 1992 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5588_6
timestamp 1731220447
transform 1 0 1784 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5587_6
timestamp 1731220447
transform 1 0 1600 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5586_6
timestamp 1731220447
transform 1 0 1392 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5585_6
timestamp 1731220447
transform 1 0 1784 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5584_6
timestamp 1731220447
transform 1 0 1648 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5583_6
timestamp 1731220447
transform 1 0 1504 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5582_6
timestamp 1731220447
transform 1 0 1352 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5581_6
timestamp 1731220447
transform 1 0 1200 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5580_6
timestamp 1731220447
transform 1 0 1208 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5579_6
timestamp 1731220447
transform 1 0 1352 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5578_6
timestamp 1731220447
transform 1 0 1784 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5577_6
timestamp 1731220447
transform 1 0 1648 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5576_6
timestamp 1731220447
transform 1 0 1504 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5575_6
timestamp 1731220447
transform 1 0 1376 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5574_6
timestamp 1731220447
transform 1 0 1240 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5573_6
timestamp 1731220447
transform 1 0 1512 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5572_6
timestamp 1731220447
transform 1 0 1648 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5571_6
timestamp 1731220447
transform 1 0 1784 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5570_6
timestamp 1731220447
transform 1 0 1784 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5569_6
timestamp 1731220447
transform 1 0 1992 0 -1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5568_6
timestamp 1731220447
transform 1 0 1992 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5567_6
timestamp 1731220447
transform 1 0 2128 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5566_6
timestamp 1731220447
transform 1 0 2536 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5565_6
timestamp 1731220447
transform 1 0 2400 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5564_6
timestamp 1731220447
transform 1 0 2264 0 1 2948
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5563_6
timestamp 1731220447
transform 1 0 2064 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5562_6
timestamp 1731220447
transform 1 0 2648 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5561_6
timestamp 1731220447
transform 1 0 2456 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5560_6
timestamp 1731220447
transform 1 0 2264 0 -1 3184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5559_6
timestamp 1731220447
transform 1 0 2248 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5558_6
timestamp 1731220447
transform 1 0 2472 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5557_6
timestamp 1731220447
transform 1 0 2688 0 1 3192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5556_6
timestamp 1731220447
transform 1 0 3296 0 -1 3416
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5555_6
timestamp 1731220447
transform 1 0 2920 0 -1 3416
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5554_6
timestamp 1731220447
transform 1 0 2552 0 -1 3416
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5553_6
timestamp 1731220447
transform 1 0 2200 0 -1 3416
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5552_6
timestamp 1731220447
transform 1 0 2568 0 1 3452
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5551_6
timestamp 1731220447
transform 1 0 2432 0 1 3452
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5550_6
timestamp 1731220447
transform 1 0 2296 0 1 3452
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5549_6
timestamp 1731220447
transform 1 0 2160 0 1 3452
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5548_6
timestamp 1731220447
transform 1 0 2200 0 -1 3692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5547_6
timestamp 1731220447
transform 1 0 2840 0 -1 3692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5546_6
timestamp 1731220447
transform 1 0 2632 0 -1 3692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5545_6
timestamp 1731220447
transform 1 0 2416 0 -1 3692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5544_6
timestamp 1731220447
transform 1 0 2384 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5543_6
timestamp 1731220447
transform 1 0 2248 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5542_6
timestamp 1731220447
transform 1 0 2112 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5541_6
timestamp 1731220447
transform 1 0 2520 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5540_6
timestamp 1731220447
transform 1 0 2656 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5539_6
timestamp 1731220447
transform 1 0 2792 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5538_6
timestamp 1731220447
transform 1 0 3232 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5537_6
timestamp 1731220447
transform 1 0 3080 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5536_6
timestamp 1731220447
transform 1 0 2936 0 1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5535_6
timestamp 1731220447
transform 1 0 2880 0 -1 3932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5534_6
timestamp 1731220447
transform 1 0 2728 0 -1 3932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5533_6
timestamp 1731220447
transform 1 0 3208 0 -1 3932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5532_6
timestamp 1731220447
transform 1 0 3040 0 -1 3932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5531_6
timestamp 1731220447
transform 1 0 2896 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5530_6
timestamp 1731220447
transform 1 0 3040 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5529_6
timestamp 1731220447
transform 1 0 3184 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5528_6
timestamp 1731220447
transform 1 0 3336 0 1 3960
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5527_6
timestamp 1731220447
transform 1 0 3360 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5526_6
timestamp 1731220447
transform 1 0 3208 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5525_6
timestamp 1731220447
transform 1 0 3064 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5524_6
timestamp 1731220447
transform 1 0 2920 0 -1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5523_6
timestamp 1731220447
transform 1 0 3440 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5522_6
timestamp 1731220447
transform 1 0 3216 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5521_6
timestamp 1731220447
transform 1 0 2992 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5520_6
timestamp 1731220447
transform 1 0 2776 0 1 4248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5519_6
timestamp 1731220447
transform 1 0 2672 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5518_6
timestamp 1731220447
transform 1 0 2808 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5517_6
timestamp 1731220447
transform 1 0 2944 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5516_6
timestamp 1731220447
transform 1 0 2960 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5515_6
timestamp 1731220447
transform 1 0 2784 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5514_6
timestamp 1731220447
transform 1 0 2608 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5513_6
timestamp 1731220447
transform 1 0 2440 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5512_6
timestamp 1731220447
transform 1 0 2872 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5511_6
timestamp 1731220447
transform 1 0 2696 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5510_6
timestamp 1731220447
transform 1 0 2528 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5509_6
timestamp 1731220447
transform 1 0 2360 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5508_6
timestamp 1731220447
transform 1 0 2200 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5507_6
timestamp 1731220447
transform 1 0 2048 0 -1 4724
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5506_6
timestamp 1731220447
transform 1 0 2120 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5505_6
timestamp 1731220447
transform 1 0 2272 0 1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5504_6
timestamp 1731220447
transform 1 0 2536 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5503_6
timestamp 1731220447
transform 1 0 2400 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5502_6
timestamp 1731220447
transform 1 0 2264 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5501_6
timestamp 1731220447
transform 1 0 2128 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5500_6
timestamp 1731220447
transform 1 0 1992 0 -1 4488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5499_6
timestamp 1731220447
transform 1 0 1784 0 -1 4444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5498_6
timestamp 1731220447
transform 1 0 1784 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5497_6
timestamp 1731220447
transform 1 0 1648 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5496_6
timestamp 1731220447
transform 1 0 1512 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5495_6
timestamp 1731220447
transform 1 0 1376 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5494_6
timestamp 1731220447
transform 1 0 1240 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5493_6
timestamp 1731220447
transform 1 0 1240 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5492_6
timestamp 1731220447
transform 1 0 1376 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5491_6
timestamp 1731220447
transform 1 0 1512 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5490_6
timestamp 1731220447
transform 1 0 1784 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5489_6
timestamp 1731220447
transform 1 0 1648 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5488_6
timestamp 1731220447
transform 1 0 1512 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5487_6
timestamp 1731220447
transform 1 0 1376 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5486_6
timestamp 1731220447
transform 1 0 1648 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5485_6
timestamp 1731220447
transform 1 0 1784 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5484_6
timestamp 1731220447
transform 1 0 1784 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5483_6
timestamp 1731220447
transform 1 0 1648 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5482_6
timestamp 1731220447
transform 1 0 1512 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5481_6
timestamp 1731220447
transform 1 0 1368 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5480_6
timestamp 1731220447
transform 1 0 1480 0 1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5479_6
timestamp 1731220447
transform 1 0 1720 0 1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5478_6
timestamp 1731220447
transform 1 0 1648 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5477_6
timestamp 1731220447
transform 1 0 1384 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5476_6
timestamp 1731220447
transform 1 0 1312 0 1 3516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5475_6
timestamp 1731220447
transform 1 0 1584 0 1 3516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5474_6
timestamp 1731220447
transform 1 0 1528 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5473_6
timestamp 1731220447
transform 1 0 1264 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5472_6
timestamp 1731220447
transform 1 0 1216 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5471_6
timestamp 1731220447
transform 1 0 1472 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5470_6
timestamp 1731220447
transform 1 0 1424 0 -1 3268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5469_6
timestamp 1731220447
transform 1 0 1168 0 -1 3268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5468_6
timestamp 1731220447
transform 1 0 1160 0 1 3040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5467_6
timestamp 1731220447
transform 1 0 1368 0 1 3040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5466_6
timestamp 1731220447
transform 1 0 1536 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5465_6
timestamp 1731220447
transform 1 0 1272 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5464_6
timestamp 1731220447
transform 1 0 1104 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5463_6
timestamp 1731220447
transform 1 0 968 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5462_6
timestamp 1731220447
transform 1 0 832 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5461_6
timestamp 1731220447
transform 1 0 904 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5460_6
timestamp 1731220447
transform 1 0 1056 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5459_6
timestamp 1731220447
transform 1 0 1040 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5458_6
timestamp 1731220447
transform 1 0 880 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5457_6
timestamp 1731220447
transform 1 0 712 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5456_6
timestamp 1731220447
transform 1 0 792 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5455_6
timestamp 1731220447
transform 1 0 1192 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5454_6
timestamp 1731220447
transform 1 0 992 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5453_6
timestamp 1731220447
transform 1 0 976 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5452_6
timestamp 1731220447
transform 1 0 784 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5451_6
timestamp 1731220447
transform 1 0 776 0 -1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5450_6
timestamp 1731220447
transform 1 0 640 0 -1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5449_6
timestamp 1731220447
transform 1 0 912 0 -1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5448_6
timestamp 1731220447
transform 1 0 864 0 1 2076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5447_6
timestamp 1731220447
transform 1 0 728 0 1 2076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5446_6
timestamp 1731220447
transform 1 0 632 0 -1 2044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5445_6
timestamp 1731220447
transform 1 0 448 0 -1 2044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5444_6
timestamp 1731220447
transform 1 0 288 0 -1 2044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5443_6
timestamp 1731220447
transform 1 0 648 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5442_6
timestamp 1731220447
transform 1 0 416 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5441_6
timestamp 1731220447
transform 1 0 184 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5440_6
timestamp 1731220447
transform 1 0 128 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5439_6
timestamp 1731220447
transform 1 0 336 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5438_6
timestamp 1731220447
transform 1 0 560 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5437_6
timestamp 1731220447
transform 1 0 352 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5436_6
timestamp 1731220447
transform 1 0 128 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5435_6
timestamp 1731220447
transform 1 0 128 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5434_6
timestamp 1731220447
transform 1 0 232 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5433_6
timestamp 1731220447
transform 1 0 352 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5432_6
timestamp 1731220447
transform 1 0 128 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5431_6
timestamp 1731220447
transform 1 0 144 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5430_6
timestamp 1731220447
transform 1 0 128 0 -1 1064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5429_6
timestamp 1731220447
transform 1 0 128 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5428_6
timestamp 1731220447
transform 1 0 128 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5427_6
timestamp 1731220447
transform 1 0 128 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5426_6
timestamp 1731220447
transform 1 0 128 0 1 376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5425_6
timestamp 1731220447
transform 1 0 352 0 1 376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5424_6
timestamp 1731220447
transform 1 0 272 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5423_6
timestamp 1731220447
transform 1 0 128 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5422_6
timestamp 1731220447
transform 1 0 128 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5421_6
timestamp 1731220447
transform 1 0 264 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5420_6
timestamp 1731220447
transform 1 0 400 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5419_6
timestamp 1731220447
transform 1 0 536 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5418_6
timestamp 1731220447
transform 1 0 672 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5417_6
timestamp 1731220447
transform 1 0 808 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5416_6
timestamp 1731220447
transform 1 0 1080 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5415_6
timestamp 1731220447
transform 1 0 944 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5414_6
timestamp 1731220447
transform 1 0 800 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5413_6
timestamp 1731220447
transform 1 0 624 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5412_6
timestamp 1731220447
transform 1 0 448 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5411_6
timestamp 1731220447
transform 1 0 1080 0 1 376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5410_6
timestamp 1731220447
transform 1 0 840 0 1 376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5409_6
timestamp 1731220447
transform 1 0 600 0 1 376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5408_6
timestamp 1731220447
transform 1 0 344 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5407_6
timestamp 1731220447
transform 1 0 968 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5406_6
timestamp 1731220447
transform 1 0 1104 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5405_6
timestamp 1731220447
transform 1 0 1112 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5404_6
timestamp 1731220447
transform 1 0 1176 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5403_6
timestamp 1731220447
transform 1 0 1488 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5402_6
timestamp 1731220447
transform 1 0 1424 0 -1 1064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5401_6
timestamp 1731220447
transform 1 0 1080 0 -1 1064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5400_6
timestamp 1731220447
transform 1 0 1016 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5399_6
timestamp 1731220447
transform 1 0 848 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5398_6
timestamp 1731220447
transform 1 0 768 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5397_6
timestamp 1731220447
transform 1 0 960 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5396_6
timestamp 1731220447
transform 1 0 1056 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5395_6
timestamp 1731220447
transform 1 0 1336 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5394_6
timestamp 1731220447
transform 1 0 1152 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5393_6
timestamp 1731220447
transform 1 0 952 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5392_6
timestamp 1731220447
transform 1 0 1344 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5391_6
timestamp 1731220447
transform 1 0 1544 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5390_6
timestamp 1731220447
transform 1 0 1544 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5389_6
timestamp 1731220447
transform 1 0 1304 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5388_6
timestamp 1731220447
transform 1 0 1720 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5387_6
timestamp 1731220447
transform 1 0 1528 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5386_6
timestamp 1731220447
transform 1 0 1344 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5385_6
timestamp 1731220447
transform 1 0 1344 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5384_6
timestamp 1731220447
transform 1 0 1784 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5383_6
timestamp 1731220447
transform 1 0 1576 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5382_6
timestamp 1731220447
transform 1 0 1552 0 -1 2044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5381_6
timestamp 1731220447
transform 1 0 1784 0 -1 2044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5380_6
timestamp 1731220447
transform 1 0 1992 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5379_6
timestamp 1731220447
transform 1 0 1992 0 -1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5378_6
timestamp 1731220447
transform 1 0 2208 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5377_6
timestamp 1731220447
transform 1 0 2704 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5376_6
timestamp 1731220447
transform 1 0 2456 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5375_6
timestamp 1731220447
transform 1 0 2408 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5374_6
timestamp 1731220447
transform 1 0 2128 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5373_6
timestamp 1731220447
transform 1 0 2304 0 1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5372_6
timestamp 1731220447
transform 1 0 2496 0 1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5371_6
timestamp 1731220447
transform 1 0 2688 0 1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5370_6
timestamp 1731220447
transform 1 0 2576 0 -1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5369_6
timestamp 1731220447
transform 1 0 2440 0 -1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5368_6
timestamp 1731220447
transform 1 0 2352 0 1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5367_6
timestamp 1731220447
transform 1 0 2560 0 1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5366_6
timestamp 1731220447
transform 1 0 2776 0 1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5365_6
timestamp 1731220447
transform 1 0 2768 0 -1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5364_6
timestamp 1731220447
transform 1 0 2512 0 -1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5363_6
timestamp 1731220447
transform 1 0 2296 0 -1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5362_6
timestamp 1731220447
transform 1 0 2128 0 -1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5361_6
timestamp 1731220447
transform 1 0 1992 0 -1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5360_6
timestamp 1731220447
transform 1 0 2488 0 1 1256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5359_6
timestamp 1731220447
transform 1 0 1992 0 1 1256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5358_6
timestamp 1731220447
transform 1 0 1784 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5357_6
timestamp 1731220447
transform 1 0 1640 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5356_6
timestamp 1731220447
transform 1 0 1472 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5355_6
timestamp 1731220447
transform 1 0 1304 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5354_6
timestamp 1731220447
transform 1 0 1136 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5353_6
timestamp 1731220447
transform 1 0 1176 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5352_6
timestamp 1731220447
transform 1 0 1328 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5351_6
timestamp 1731220447
transform 1 0 1480 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5350_6
timestamp 1731220447
transform 1 0 1640 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5349_6
timestamp 1731220447
transform 1 0 1784 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5348_6
timestamp 1731220447
transform 1 0 1776 0 -1 1064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5347_6
timestamp 1731220447
transform 1 0 1784 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5346_6
timestamp 1731220447
transform 1 0 1992 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5345_6
timestamp 1731220447
transform 1 0 2128 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5344_6
timestamp 1731220447
transform 1 0 2152 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5343_6
timestamp 1731220447
transform 1 0 2408 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5342_6
timestamp 1731220447
transform 1 0 2280 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5341_6
timestamp 1731220447
transform 1 0 2440 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5340_6
timestamp 1731220447
transform 1 0 2600 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5339_6
timestamp 1731220447
transform 1 0 2680 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5338_6
timestamp 1731220447
transform 1 0 2464 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5337_6
timestamp 1731220447
transform 1 0 2248 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5336_6
timestamp 1731220447
transform 1 0 2240 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5335_6
timestamp 1731220447
transform 1 0 2376 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5334_6
timestamp 1731220447
transform 1 0 2520 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5333_6
timestamp 1731220447
transform 1 0 2672 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5332_6
timestamp 1731220447
transform 1 0 2824 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5331_6
timestamp 1731220447
transform 1 0 2712 0 -1 1192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5330_6
timestamp 1731220447
transform 1 0 2984 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5329_6
timestamp 1731220447
transform 1 0 3152 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5328_6
timestamp 1731220447
transform 1 0 3328 0 -1 1192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5327_6
timestamp 1731220447
transform 1 0 3016 0 -1 1192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5326_6
timestamp 1731220447
transform 1 0 3016 0 1 1256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5325_6
timestamp 1731220447
transform 1 0 3360 0 -1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5324_6
timestamp 1731220447
transform 1 0 3056 0 -1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5323_6
timestamp 1731220447
transform 1 0 3000 0 1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5322_6
timestamp 1731220447
transform 1 0 2848 0 -1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5321_6
timestamp 1731220447
transform 1 0 2712 0 -1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5320_6
timestamp 1731220447
transform 1 0 3144 0 -1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5319_6
timestamp 1731220447
transform 1 0 2992 0 -1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5318_6
timestamp 1731220447
transform 1 0 2880 0 1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5317_6
timestamp 1731220447
transform 1 0 3064 0 1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5316_6
timestamp 1731220447
transform 1 0 3176 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5315_6
timestamp 1731220447
transform 1 0 2928 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5314_6
timestamp 1731220447
transform 1 0 2672 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5313_6
timestamp 1731220447
transform 1 0 2960 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5312_6
timestamp 1731220447
transform 1 0 3216 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5311_6
timestamp 1731220447
transform 1 0 3480 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5310_6
timestamp 1731220447
transform 1 0 3424 0 -1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5309_6
timestamp 1731220447
transform 1 0 3176 0 -1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5308_6
timestamp 1731220447
transform 1 0 3648 0 -1 2184
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5307_6
timestamp 1731220447
transform 1 0 3856 0 -1 2224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5306_6
timestamp 1731220447
transform 1 0 4320 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5305_6
timestamp 1731220447
transform 1 0 4080 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5304_6
timestamp 1731220447
transform 1 0 3856 0 1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5303_6
timestamp 1731220447
transform 1 0 3856 0 -1 2000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5302_6
timestamp 1731220447
transform 1 0 3648 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5301_6
timestamp 1731220447
transform 1 0 3424 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5300_6
timestamp 1731220447
transform 1 0 3632 0 1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5299_6
timestamp 1731220447
transform 1 0 3440 0 1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5298_6
timestamp 1731220447
transform 1 0 3248 0 1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5297_6
timestamp 1731220447
transform 1 0 3296 0 -1 1704
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5296_6
timestamp 1731220447
transform 1 0 3224 0 1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5295_6
timestamp 1731220447
transform 1 0 3456 0 1 1480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5294_6
timestamp 1731220447
transform 1 0 3552 0 1 1256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5293_6
timestamp 1731220447
transform 1 0 3648 0 -1 1192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5292_6
timestamp 1731220447
transform 1 0 3496 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5291_6
timestamp 1731220447
transform 1 0 3320 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5290_6
timestamp 1731220447
transform 1 0 3648 0 1 968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5289_6
timestamp 1731220447
transform 1 0 3640 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5288_6
timestamp 1731220447
transform 1 0 3448 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5287_6
timestamp 1731220447
transform 1 0 3264 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5286_6
timestamp 1731220447
transform 1 0 3072 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5285_6
timestamp 1731220447
transform 1 0 2880 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5284_6
timestamp 1731220447
transform 1 0 3400 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5283_6
timestamp 1731220447
transform 1 0 3240 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5282_6
timestamp 1731220447
transform 1 0 3080 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5281_6
timestamp 1731220447
transform 1 0 2920 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5280_6
timestamp 1731220447
transform 1 0 2760 0 1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5279_6
timestamp 1731220447
transform 1 0 2648 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5278_6
timestamp 1731220447
transform 1 0 2872 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5277_6
timestamp 1731220447
transform 1 0 3080 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5276_6
timestamp 1731220447
transform 1 0 3280 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5275_6
timestamp 1731220447
transform 1 0 3472 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5274_6
timestamp 1731220447
transform 1 0 3648 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5273_6
timestamp 1731220447
transform 1 0 3856 0 1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5272_6
timestamp 1731220447
transform 1 0 3856 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5271_6
timestamp 1731220447
transform 1 0 4400 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5270_6
timestamp 1731220447
transform 1 0 4264 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5269_6
timestamp 1731220447
transform 1 0 4128 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5268_6
timestamp 1731220447
transform 1 0 3992 0 -1 584
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5267_6
timestamp 1731220447
transform 1 0 3856 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5266_6
timestamp 1731220447
transform 1 0 3648 0 1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5265_6
timestamp 1731220447
transform 1 0 3448 0 1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5264_6
timestamp 1731220447
transform 1 0 3224 0 1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5263_6
timestamp 1731220447
transform 1 0 3000 0 1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5262_6
timestamp 1731220447
transform 1 0 2768 0 1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5261_6
timestamp 1731220447
transform 1 0 3624 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5260_6
timestamp 1731220447
transform 1 0 3488 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5259_6
timestamp 1731220447
transform 1 0 3352 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5258_6
timestamp 1731220447
transform 1 0 3216 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5257_6
timestamp 1731220447
transform 1 0 3080 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5256_6
timestamp 1731220447
transform 1 0 2944 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5255_6
timestamp 1731220447
transform 1 0 3624 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5254_6
timestamp 1731220447
transform 1 0 3488 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5253_6
timestamp 1731220447
transform 1 0 3352 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5252_6
timestamp 1731220447
transform 1 0 3216 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5251_6
timestamp 1731220447
transform 1 0 3080 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5250_6
timestamp 1731220447
transform 1 0 2944 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5249_6
timestamp 1731220447
transform 1 0 2808 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5248_6
timestamp 1731220447
transform 1 0 2672 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5247_6
timestamp 1731220447
transform 1 0 2536 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5246_6
timestamp 1731220447
transform 1 0 2400 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5245_6
timestamp 1731220447
transform 1 0 2264 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5244_6
timestamp 1731220447
transform 1 0 2128 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5243_6
timestamp 1731220447
transform 1 0 1992 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5242_6
timestamp 1731220447
transform 1 0 2808 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5241_6
timestamp 1731220447
transform 1 0 2672 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5240_6
timestamp 1731220447
transform 1 0 2536 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5239_6
timestamp 1731220447
transform 1 0 2400 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5238_6
timestamp 1731220447
transform 1 0 2264 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5237_6
timestamp 1731220447
transform 1 0 2128 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5236_6
timestamp 1731220447
transform 1 0 1992 0 -1 332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5235_6
timestamp 1731220447
transform 1 0 2520 0 1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5234_6
timestamp 1731220447
transform 1 0 2248 0 1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5233_6
timestamp 1731220447
transform 1 0 1992 0 1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5232_6
timestamp 1731220447
transform 1 0 1784 0 1 376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5231_6
timestamp 1731220447
transform 1 0 1560 0 1 376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5230_6
timestamp 1731220447
transform 1 0 1320 0 1 376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5229_6
timestamp 1731220447
transform 1 0 1784 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5228_6
timestamp 1731220447
transform 1 0 1640 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5227_6
timestamp 1731220447
transform 1 0 1480 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5226_6
timestamp 1731220447
transform 1 0 1312 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5225_6
timestamp 1731220447
transform 1 0 1144 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5224_6
timestamp 1731220447
transform 1 0 1784 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5223_6
timestamp 1731220447
transform 1 0 1648 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5222_6
timestamp 1731220447
transform 1 0 1512 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5221_6
timestamp 1731220447
transform 1 0 1376 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5220_6
timestamp 1731220447
transform 1 0 1240 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5219_6
timestamp 1731220447
transform 1 0 968 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5218_6
timestamp 1731220447
transform 1 0 776 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5217_6
timestamp 1731220447
transform 1 0 568 0 -1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5216_6
timestamp 1731220447
transform 1 0 696 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5215_6
timestamp 1731220447
transform 1 0 832 0 1 600
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5214_6
timestamp 1731220447
transform 1 0 856 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5213_6
timestamp 1731220447
transform 1 0 600 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5212_6
timestamp 1731220447
transform 1 0 352 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5211_6
timestamp 1731220447
transform 1 0 336 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5210_6
timestamp 1731220447
transform 1 0 592 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5209_6
timestamp 1731220447
transform 1 0 872 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5208_6
timestamp 1731220447
transform 1 0 744 0 -1 1064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5207_6
timestamp 1731220447
transform 1 0 416 0 -1 1064
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5206_6
timestamp 1731220447
transform 1 0 320 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5205_6
timestamp 1731220447
transform 1 0 496 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5204_6
timestamp 1731220447
transform 1 0 672 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5203_6
timestamp 1731220447
transform 1 0 568 0 -1 1316
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5202_6
timestamp 1731220447
transform 1 0 776 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5201_6
timestamp 1731220447
transform 1 0 504 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5200_6
timestamp 1731220447
transform 1 0 328 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5199_6
timestamp 1731220447
transform 1 0 544 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5198_6
timestamp 1731220447
transform 1 0 752 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5197_6
timestamp 1731220447
transform 1 0 592 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5196_6
timestamp 1731220447
transform 1 0 832 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5195_6
timestamp 1731220447
transform 1 0 1064 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5194_6
timestamp 1731220447
transform 1 0 1160 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5193_6
timestamp 1731220447
transform 1 0 968 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5192_6
timestamp 1731220447
transform 1 0 768 0 -1 1800
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5191_6
timestamp 1731220447
transform 1 0 880 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5190_6
timestamp 1731220447
transform 1 0 1112 0 1 1812
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5189_6
timestamp 1731220447
transform 1 0 1304 0 -1 2044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5188_6
timestamp 1731220447
transform 1 0 1064 0 -1 2044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5187_6
timestamp 1731220447
transform 1 0 840 0 -1 2044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5186_6
timestamp 1731220447
transform 1 0 592 0 1 2076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5185_6
timestamp 1731220447
transform 1 0 456 0 1 2076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5184_6
timestamp 1731220447
transform 1 0 320 0 1 2076
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5183_6
timestamp 1731220447
transform 1 0 368 0 -1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5182_6
timestamp 1731220447
transform 1 0 504 0 -1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5181_6
timestamp 1731220447
transform 1 0 592 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5180_6
timestamp 1731220447
transform 1 0 400 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5179_6
timestamp 1731220447
transform 1 0 216 0 1 2312
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5178_6
timestamp 1731220447
transform 1 0 200 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5177_6
timestamp 1731220447
transform 1 0 392 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5176_6
timestamp 1731220447
transform 1 0 592 0 -1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5175_6
timestamp 1731220447
transform 1 0 536 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5174_6
timestamp 1731220447
transform 1 0 352 0 1 2556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5173_6
timestamp 1731220447
transform 1 0 432 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5172_6
timestamp 1731220447
transform 1 0 592 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5171_6
timestamp 1731220447
transform 1 0 752 0 -1 2784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5170_6
timestamp 1731220447
transform 1 0 696 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5169_6
timestamp 1731220447
transform 1 0 560 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5168_6
timestamp 1731220447
transform 1 0 424 0 1 2792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5167_6
timestamp 1731220447
transform 1 0 544 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5166_6
timestamp 1731220447
transform 1 0 768 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5165_6
timestamp 1731220447
transform 1 0 1016 0 -1 3024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5164_6
timestamp 1731220447
transform 1 0 952 0 1 3040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5163_6
timestamp 1731220447
transform 1 0 752 0 1 3040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5162_6
timestamp 1731220447
transform 1 0 560 0 1 3040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5161_6
timestamp 1731220447
transform 1 0 376 0 1 3040
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5160_6
timestamp 1731220447
transform 1 0 920 0 -1 3268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5159_6
timestamp 1731220447
transform 1 0 672 0 -1 3268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5158_6
timestamp 1731220447
transform 1 0 432 0 -1 3268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5157_6
timestamp 1731220447
transform 1 0 208 0 -1 3268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5156_6
timestamp 1731220447
transform 1 0 968 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5155_6
timestamp 1731220447
transform 1 0 728 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5154_6
timestamp 1731220447
transform 1 0 504 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5153_6
timestamp 1731220447
transform 1 0 296 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5152_6
timestamp 1731220447
transform 1 0 128 0 1 3272
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5151_6
timestamp 1731220447
transform 1 0 1008 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5150_6
timestamp 1731220447
transform 1 0 760 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5149_6
timestamp 1731220447
transform 1 0 520 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5148_6
timestamp 1731220447
transform 1 0 304 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5147_6
timestamp 1731220447
transform 1 0 128 0 -1 3504
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5146_6
timestamp 1731220447
transform 1 0 128 0 1 3516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5145_6
timestamp 1731220447
transform 1 0 312 0 1 3516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5144_6
timestamp 1731220447
transform 1 0 1040 0 1 3516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5143_6
timestamp 1731220447
transform 1 0 784 0 1 3516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5142_6
timestamp 1731220447
transform 1 0 536 0 1 3516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5141_6
timestamp 1731220447
transform 1 0 400 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5140_6
timestamp 1731220447
transform 1 0 200 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5139_6
timestamp 1731220447
transform 1 0 1120 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5138_6
timestamp 1731220447
transform 1 0 864 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5137_6
timestamp 1731220447
transform 1 0 624 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5136_6
timestamp 1731220447
transform 1 0 616 0 1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5135_6
timestamp 1731220447
transform 1 0 432 0 1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5134_6
timestamp 1731220447
transform 1 0 1248 0 1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5133_6
timestamp 1731220447
transform 1 0 1024 0 1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5132_6
timestamp 1731220447
transform 1 0 816 0 1 3752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5131_6
timestamp 1731220447
transform 1 0 800 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5130_6
timestamp 1731220447
transform 1 0 664 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5129_6
timestamp 1731220447
transform 1 0 1224 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5128_6
timestamp 1731220447
transform 1 0 1080 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5127_6
timestamp 1731220447
transform 1 0 936 0 -1 3980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5126_6
timestamp 1731220447
transform 1 0 832 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5125_6
timestamp 1731220447
transform 1 0 696 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5124_6
timestamp 1731220447
transform 1 0 968 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5123_6
timestamp 1731220447
transform 1 0 1104 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5122_6
timestamp 1731220447
transform 1 0 1240 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5121_6
timestamp 1731220447
transform 1 0 1104 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5120_6
timestamp 1731220447
transform 1 0 968 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5119_6
timestamp 1731220447
transform 1 0 832 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5118_6
timestamp 1731220447
transform 1 0 696 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5117_6
timestamp 1731220447
transform 1 0 560 0 -1 4208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5116_6
timestamp 1731220447
transform 1 0 1104 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5115_6
timestamp 1731220447
transform 1 0 968 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5114_6
timestamp 1731220447
transform 1 0 832 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5113_6
timestamp 1731220447
transform 1 0 696 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5112_6
timestamp 1731220447
transform 1 0 560 0 1 4220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5111_6
timestamp 1731220447
transform 1 0 1520 0 -1 4444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5110_6
timestamp 1731220447
transform 1 0 1232 0 -1 4444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5109_6
timestamp 1731220447
transform 1 0 960 0 -1 4444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5108_6
timestamp 1731220447
transform 1 0 712 0 -1 4444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5107_6
timestamp 1731220447
transform 1 0 488 0 -1 4444
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5106_6
timestamp 1731220447
transform 1 0 832 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5105_6
timestamp 1731220447
transform 1 0 696 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5104_6
timestamp 1731220447
transform 1 0 560 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5103_6
timestamp 1731220447
transform 1 0 424 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5102_6
timestamp 1731220447
transform 1 0 288 0 1 4460
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5101_6
timestamp 1731220447
transform 1 0 672 0 -1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5100_6
timestamp 1731220447
transform 1 0 536 0 -1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_599_6
timestamp 1731220447
transform 1 0 400 0 -1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_598_6
timestamp 1731220447
transform 1 0 264 0 -1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_597_6
timestamp 1731220447
transform 1 0 128 0 -1 4700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_596_6
timestamp 1731220447
transform 1 0 1248 0 1 4720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_595_6
timestamp 1731220447
transform 1 0 856 0 1 4720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_594_6
timestamp 1731220447
transform 1 0 472 0 1 4720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_593_6
timestamp 1731220447
transform 1 0 128 0 1 4720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_592_6
timestamp 1731220447
transform 1 0 128 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_591_6
timestamp 1731220447
transform 1 0 360 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_590_6
timestamp 1731220447
transform 1 0 616 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_589_6
timestamp 1731220447
transform 1 0 528 0 1 4956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_588_6
timestamp 1731220447
transform 1 0 336 0 1 4956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_587_6
timestamp 1731220447
transform 1 0 144 0 1 4956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_586_6
timestamp 1731220447
transform 1 0 176 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_585_6
timestamp 1731220447
transform 1 0 312 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_584_6
timestamp 1731220447
transform 1 0 584 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_583_6
timestamp 1731220447
transform 1 0 448 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_582_6
timestamp 1731220447
transform 1 0 408 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_581_6
timestamp 1731220447
transform 1 0 584 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_580_6
timestamp 1731220447
transform 1 0 760 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_579_6
timestamp 1731220447
transform 1 0 936 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_578_6
timestamp 1731220447
transform 1 0 856 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_577_6
timestamp 1731220447
transform 1 0 720 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_576_6
timestamp 1731220447
transform 1 0 992 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_575_6
timestamp 1731220447
transform 1 0 1128 0 1 4956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_574_6
timestamp 1731220447
transform 1 0 928 0 1 4956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_573_6
timestamp 1731220447
transform 1 0 728 0 1 4956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_572_6
timestamp 1731220447
transform 1 0 864 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_571_6
timestamp 1731220447
transform 1 0 1104 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_570_6
timestamp 1731220447
transform 1 0 1336 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_569_6
timestamp 1731220447
transform 1 0 1568 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_568_6
timestamp 1731220447
transform 1 0 1640 0 1 4720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_567_6
timestamp 1731220447
transform 1 0 1784 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_566_6
timestamp 1731220447
transform 1 0 1992 0 1 4772
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_565_6
timestamp 1731220447
transform 1 0 1992 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_564_6
timestamp 1731220447
transform 1 0 2136 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_563_6
timestamp 1731220447
transform 1 0 2720 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_562_6
timestamp 1731220447
transform 1 0 2512 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_561_6
timestamp 1731220447
transform 1 0 2320 0 -1 5004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_560_6
timestamp 1731220447
transform 1 0 2304 0 1 5028
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_559_6
timestamp 1731220447
transform 1 0 2136 0 1 5028
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_558_6
timestamp 1731220447
transform 1 0 2488 0 1 5028
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_557_6
timestamp 1731220447
transform 1 0 2912 0 1 5028
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_556_6
timestamp 1731220447
transform 1 0 2688 0 1 5028
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_555_6
timestamp 1731220447
transform 1 0 2656 0 -1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_554_6
timestamp 1731220447
transform 1 0 2480 0 -1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_553_6
timestamp 1731220447
transform 1 0 2832 0 -1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_552_6
timestamp 1731220447
transform 1 0 2808 0 1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_551_6
timestamp 1731220447
transform 1 0 2640 0 1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_550_6
timestamp 1731220447
transform 1 0 2976 0 1 5260
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_549_6
timestamp 1731220447
transform 1 0 2920 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_548_6
timestamp 1731220447
transform 1 0 3072 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_547_6
timestamp 1731220447
transform 1 0 3224 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_546_6
timestamp 1731220447
transform 1 0 3384 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_545_6
timestamp 1731220447
transform 1 0 3648 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_544_6
timestamp 1731220447
transform 1 0 3472 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_543_6
timestamp 1731220447
transform 1 0 3272 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_542_6
timestamp 1731220447
transform 1 0 3072 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_541_6
timestamp 1731220447
transform 1 0 2864 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_540_6
timestamp 1731220447
transform 1 0 3088 0 -1 5756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_539_6
timestamp 1731220447
transform 1 0 2928 0 -1 5756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_538_6
timestamp 1731220447
transform 1 0 2776 0 -1 5756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_537_6
timestamp 1731220447
transform 1 0 2624 0 -1 5756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_536_6
timestamp 1731220447
transform 1 0 2480 0 -1 5756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_535_6
timestamp 1731220447
transform 1 0 2344 0 -1 5756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_534_6
timestamp 1731220447
transform 1 0 2648 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_533_6
timestamp 1731220447
transform 1 0 2424 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_532_6
timestamp 1731220447
transform 1 0 2200 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_531_6
timestamp 1731220447
transform 1 0 1992 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_530_6
timestamp 1731220447
transform 1 0 1784 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_529_6
timestamp 1731220447
transform 1 0 1648 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_528_6
timestamp 1731220447
transform 1 0 1504 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_527_6
timestamp 1731220447
transform 1 0 1352 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_526_6
timestamp 1731220447
transform 1 0 1240 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_525_6
timestamp 1731220447
transform 1 0 1784 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_524_6
timestamp 1731220447
transform 1 0 1648 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_523_6
timestamp 1731220447
transform 1 0 1512 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_522_6
timestamp 1731220447
transform 1 0 1376 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_521_6
timestamp 1731220447
transform 1 0 1784 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_520_6
timestamp 1731220447
transform 1 0 1608 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_519_6
timestamp 1731220447
transform 1 0 1440 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_518_6
timestamp 1731220447
transform 1 0 1272 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_517_6
timestamp 1731220447
transform 1 0 1104 0 1 5208
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_516_6
timestamp 1731220447
transform 1 0 1104 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_515_6
timestamp 1731220447
transform 1 0 968 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_514_6
timestamp 1731220447
transform 1 0 832 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_513_6
timestamp 1731220447
transform 1 0 696 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_512_6
timestamp 1731220447
transform 1 0 560 0 -1 5456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_511_6
timestamp 1731220447
transform 1 0 1200 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_510_6
timestamp 1731220447
transform 1 0 1048 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_59_6
timestamp 1731220447
transform 1 0 896 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_58_6
timestamp 1731220447
transform 1 0 752 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_57_6
timestamp 1731220447
transform 1 0 616 0 1 5464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_56_6
timestamp 1731220447
transform 1 0 944 0 -1 5716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_55_6
timestamp 1731220447
transform 1 0 808 0 -1 5716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_54_6
timestamp 1731220447
transform 1 0 672 0 -1 5716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_53_6
timestamp 1731220447
transform 1 0 536 0 -1 5716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_52_6
timestamp 1731220447
transform 1 0 400 0 -1 5716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_51_6
timestamp 1731220447
transform 1 0 264 0 -1 5716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_50_6
timestamp 1731220447
transform 1 0 128 0 -1 5716
box 3 5 132 108
<< end >>
