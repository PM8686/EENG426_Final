magic
tech sky130l
timestamp 1730592110
<< m1 >>
rect 704 563 708 607
rect 528 467 532 531
rect 592 443 596 547
rect 704 467 708 511
rect 128 359 132 411
rect 704 359 708 411
rect 704 263 708 307
<< m2c >>
rect 111 801 115 805
rect 775 801 779 805
rect 111 783 115 787
rect 775 783 779 787
rect 203 771 207 775
rect 259 771 263 775
rect 315 771 319 775
rect 371 771 375 775
rect 427 771 431 775
rect 483 771 487 775
rect 547 771 551 775
rect 610 771 614 775
rect 730 771 734 775
rect 402 755 406 759
rect 730 755 734 759
rect 186 751 190 755
rect 250 751 254 755
rect 322 751 326 755
rect 490 751 494 755
rect 578 751 582 755
rect 666 751 670 755
rect 111 741 115 745
rect 775 741 779 745
rect 111 723 115 727
rect 775 723 779 727
rect 111 689 115 693
rect 775 689 779 693
rect 111 671 115 675
rect 775 671 779 675
rect 234 659 238 663
rect 338 659 342 663
rect 442 659 446 663
rect 547 659 551 663
rect 651 659 655 663
rect 730 659 734 663
rect 482 647 486 651
rect 730 647 734 651
rect 290 643 294 647
rect 346 643 350 647
rect 410 643 414 647
rect 562 643 566 647
rect 650 643 654 647
rect 111 633 115 637
rect 775 633 779 637
rect 111 615 115 619
rect 775 615 779 619
rect 704 607 708 611
rect 111 589 115 593
rect 111 571 115 575
rect 775 589 779 593
rect 775 571 779 575
rect 354 559 358 563
rect 418 559 422 563
rect 490 559 494 563
rect 570 559 574 563
rect 658 559 662 563
rect 704 559 708 563
rect 730 559 734 563
rect 562 551 566 555
rect 730 551 734 555
rect 330 547 334 551
rect 402 547 406 551
rect 482 547 486 551
rect 592 547 596 551
rect 650 547 654 551
rect 111 537 115 541
rect 528 531 532 535
rect 111 519 115 523
rect 111 493 115 497
rect 111 475 115 479
rect 203 463 207 467
rect 291 463 295 467
rect 387 463 391 467
rect 499 463 503 467
rect 528 463 532 467
rect 458 451 462 455
rect 154 447 158 451
rect 210 447 214 451
rect 282 447 286 451
rect 370 447 374 451
rect 554 447 558 451
rect 775 537 779 541
rect 775 519 779 523
rect 704 511 708 515
rect 775 493 779 497
rect 775 475 779 479
rect 618 463 622 467
rect 704 463 708 467
rect 730 463 734 467
rect 650 451 654 455
rect 730 447 734 451
rect 111 437 115 441
rect 592 439 596 443
rect 775 437 779 441
rect 111 419 115 423
rect 775 419 779 423
rect 128 411 132 415
rect 111 385 115 389
rect 111 367 115 371
rect 704 411 708 415
rect 775 385 779 389
rect 775 367 779 371
rect 128 355 132 359
rect 154 355 158 359
rect 234 355 238 359
rect 322 355 326 359
rect 418 355 422 359
rect 522 355 526 359
rect 634 355 638 359
rect 704 355 708 359
rect 730 355 734 359
rect 546 347 550 351
rect 674 347 678 351
rect 298 343 302 347
rect 354 343 358 347
rect 418 343 422 347
rect 482 343 486 347
rect 610 343 614 347
rect 730 343 734 347
rect 111 333 115 337
rect 775 333 779 337
rect 111 315 115 319
rect 775 315 779 319
rect 704 307 708 311
rect 111 289 115 293
rect 111 271 115 275
rect 775 289 779 293
rect 775 271 779 275
rect 227 259 231 263
rect 283 259 287 263
rect 339 259 343 263
rect 395 259 399 263
rect 450 259 454 263
rect 507 259 511 263
rect 563 259 567 263
rect 619 259 623 263
rect 675 259 679 263
rect 704 259 708 263
rect 730 259 734 263
rect 514 239 518 243
rect 290 235 294 239
rect 346 235 350 239
rect 402 235 406 239
rect 458 235 462 239
rect 111 225 115 229
rect 775 225 779 229
rect 111 207 115 211
rect 775 207 779 211
rect 111 177 115 181
rect 775 177 779 181
rect 111 159 115 163
rect 775 159 779 163
rect 171 147 175 151
rect 227 147 231 151
rect 283 147 287 151
rect 339 147 343 151
rect 394 147 398 151
rect 546 127 550 131
rect 154 123 158 127
rect 210 123 214 127
rect 266 123 270 127
rect 322 123 326 127
rect 378 123 382 127
rect 434 123 438 127
rect 490 123 494 127
rect 111 113 115 117
rect 775 113 779 117
rect 111 95 115 99
rect 775 95 779 99
<< m2 >>
rect 194 813 200 814
rect 194 809 195 813
rect 199 809 200 813
rect 194 808 200 809
rect 250 813 256 814
rect 250 809 251 813
rect 255 809 256 813
rect 250 808 256 809
rect 306 813 312 814
rect 306 809 307 813
rect 311 809 312 813
rect 306 808 312 809
rect 362 813 368 814
rect 362 809 363 813
rect 367 809 368 813
rect 362 808 368 809
rect 418 813 424 814
rect 418 809 419 813
rect 423 809 424 813
rect 418 808 424 809
rect 474 813 480 814
rect 474 809 475 813
rect 479 809 480 813
rect 474 808 480 809
rect 538 813 544 814
rect 538 809 539 813
rect 543 809 544 813
rect 538 808 544 809
rect 602 813 608 814
rect 602 809 603 813
rect 607 809 608 813
rect 602 808 608 809
rect 666 813 672 814
rect 666 809 667 813
rect 671 809 672 813
rect 666 808 672 809
rect 722 813 728 814
rect 722 809 723 813
rect 727 809 728 813
rect 722 808 728 809
rect 110 805 116 806
rect 110 801 111 805
rect 115 801 116 805
rect 110 800 116 801
rect 774 805 780 806
rect 774 801 775 805
rect 779 801 780 805
rect 774 800 780 801
rect 110 787 116 788
rect 110 783 111 787
rect 115 783 116 787
rect 110 782 116 783
rect 194 787 200 788
rect 194 783 195 787
rect 199 783 200 787
rect 734 787 740 788
rect 734 786 735 787
rect 194 782 200 783
rect 208 784 249 786
rect 264 784 305 786
rect 319 784 361 786
rect 376 784 417 786
rect 432 784 473 786
rect 488 784 537 786
rect 552 784 601 786
rect 673 784 718 786
rect 729 784 735 786
rect 208 776 210 784
rect 264 776 266 784
rect 319 776 321 784
rect 376 776 378 784
rect 432 776 434 784
rect 488 776 490 784
rect 552 776 554 784
rect 202 775 210 776
rect 202 771 203 775
rect 207 772 210 775
rect 218 775 224 776
rect 207 771 208 772
rect 202 770 208 771
rect 218 771 219 775
rect 223 771 224 775
rect 218 770 224 771
rect 258 775 266 776
rect 258 771 259 775
rect 263 772 266 775
rect 274 775 280 776
rect 263 771 264 772
rect 258 770 264 771
rect 274 771 275 775
rect 279 771 280 775
rect 274 770 280 771
rect 314 775 321 776
rect 314 771 315 775
rect 319 772 321 775
rect 330 775 336 776
rect 319 771 320 772
rect 314 770 320 771
rect 330 771 331 775
rect 335 771 336 775
rect 330 770 336 771
rect 370 775 378 776
rect 370 771 371 775
rect 375 772 378 775
rect 386 775 392 776
rect 375 771 376 772
rect 370 770 376 771
rect 386 771 387 775
rect 391 771 392 775
rect 386 770 392 771
rect 426 775 434 776
rect 426 771 427 775
rect 431 772 434 775
rect 442 775 448 776
rect 431 771 432 772
rect 426 770 432 771
rect 442 771 443 775
rect 447 771 448 775
rect 442 770 448 771
rect 482 775 490 776
rect 482 771 483 775
rect 487 772 490 775
rect 498 775 504 776
rect 487 771 488 772
rect 482 770 488 771
rect 498 771 499 775
rect 503 771 504 775
rect 498 770 504 771
rect 546 775 554 776
rect 546 771 547 775
rect 551 772 554 775
rect 562 775 568 776
rect 551 771 552 772
rect 546 770 552 771
rect 562 771 563 775
rect 567 771 568 775
rect 562 770 568 771
rect 574 775 580 776
rect 574 771 575 775
rect 579 774 580 775
rect 609 775 615 776
rect 609 774 610 775
rect 579 772 610 774
rect 579 771 580 772
rect 574 770 580 771
rect 609 771 610 772
rect 614 771 615 775
rect 609 770 615 771
rect 626 775 632 776
rect 626 771 627 775
rect 631 771 632 775
rect 626 770 632 771
rect 690 775 696 776
rect 690 771 691 775
rect 695 771 696 775
rect 716 774 718 784
rect 734 783 735 784
rect 739 783 740 787
rect 734 782 740 783
rect 774 787 780 788
rect 774 783 775 787
rect 779 783 780 787
rect 774 782 780 783
rect 729 775 735 776
rect 729 774 730 775
rect 716 772 730 774
rect 690 770 696 771
rect 729 771 730 772
rect 734 771 735 775
rect 729 770 735 771
rect 746 775 752 776
rect 746 771 747 775
rect 751 771 752 775
rect 746 770 752 771
rect 194 763 200 764
rect 194 759 195 763
rect 199 762 200 763
rect 199 760 366 762
rect 199 759 200 760
rect 194 758 200 759
rect 364 758 366 760
rect 401 759 407 760
rect 401 758 402 759
rect 202 757 208 758
rect 185 755 191 756
rect 185 751 186 755
rect 190 754 191 755
rect 190 752 198 754
rect 202 753 203 757
rect 207 753 208 757
rect 266 757 272 758
rect 202 752 208 753
rect 249 755 255 756
rect 190 751 191 752
rect 185 750 191 751
rect 196 750 198 752
rect 249 751 250 755
rect 254 754 255 755
rect 254 752 262 754
rect 266 753 267 757
rect 271 753 272 757
rect 338 757 344 758
rect 266 752 272 753
rect 321 755 327 756
rect 254 751 255 752
rect 249 750 255 751
rect 260 750 262 752
rect 321 751 322 755
rect 326 754 327 755
rect 326 752 334 754
rect 338 753 339 757
rect 343 753 344 757
rect 364 756 402 758
rect 401 755 402 756
rect 406 755 407 759
rect 729 759 740 760
rect 401 754 407 755
rect 418 757 424 758
rect 338 752 344 753
rect 418 753 419 757
rect 423 753 424 757
rect 506 757 512 758
rect 418 752 424 753
rect 489 755 496 756
rect 326 751 327 752
rect 321 750 327 751
rect 332 750 334 752
rect 489 751 490 755
rect 495 751 496 755
rect 506 753 507 757
rect 511 753 512 757
rect 594 757 600 758
rect 577 755 583 756
rect 577 754 578 755
rect 506 752 512 753
rect 524 752 578 754
rect 489 750 496 751
rect 196 748 242 750
rect 260 748 314 750
rect 332 748 394 750
rect 110 745 116 746
rect 240 745 242 748
rect 312 745 314 748
rect 392 745 394 748
rect 524 746 526 752
rect 577 751 578 752
rect 582 751 583 755
rect 594 753 595 757
rect 599 753 600 757
rect 682 757 688 758
rect 594 752 600 753
rect 665 755 671 756
rect 577 750 583 751
rect 665 751 666 755
rect 670 754 671 755
rect 670 752 678 754
rect 682 753 683 757
rect 687 753 688 757
rect 729 755 730 759
rect 734 755 735 759
rect 739 755 740 759
rect 729 754 740 755
rect 746 757 752 758
rect 682 752 688 753
rect 746 753 747 757
rect 751 753 752 757
rect 746 752 752 753
rect 670 751 671 752
rect 665 750 671 751
rect 676 750 678 752
rect 676 748 722 750
rect 110 741 111 745
rect 115 741 116 745
rect 489 744 526 746
rect 574 747 580 748
rect 198 743 204 744
rect 198 742 199 743
rect 110 740 116 741
rect 185 740 199 742
rect 198 739 199 740
rect 203 739 204 743
rect 574 743 575 747
rect 579 743 580 747
rect 720 745 722 748
rect 774 745 780 746
rect 574 742 580 743
rect 774 741 775 745
rect 779 741 780 745
rect 774 740 780 741
rect 198 738 204 739
rect 110 727 116 728
rect 110 723 111 727
rect 115 723 116 727
rect 110 722 116 723
rect 774 727 780 728
rect 774 723 775 727
rect 779 723 780 727
rect 774 722 780 723
rect 178 719 184 720
rect 178 715 179 719
rect 183 715 184 719
rect 178 714 184 715
rect 242 719 248 720
rect 242 715 243 719
rect 247 715 248 719
rect 242 714 248 715
rect 314 719 320 720
rect 314 715 315 719
rect 319 715 320 719
rect 314 714 320 715
rect 394 719 400 720
rect 394 715 395 719
rect 399 715 400 719
rect 394 714 400 715
rect 482 719 488 720
rect 482 715 483 719
rect 487 715 488 719
rect 482 714 488 715
rect 570 719 576 720
rect 570 715 571 719
rect 575 715 576 719
rect 658 719 664 720
rect 570 714 576 715
rect 648 712 650 717
rect 658 715 659 719
rect 663 715 664 719
rect 658 714 664 715
rect 722 719 728 720
rect 722 715 723 719
rect 727 715 728 719
rect 722 714 728 715
rect 648 711 656 712
rect 648 708 651 711
rect 650 707 651 708
rect 655 707 656 711
rect 650 706 656 707
rect 490 703 496 704
rect 226 701 232 702
rect 226 697 227 701
rect 231 697 232 701
rect 226 696 232 697
rect 330 701 336 702
rect 330 697 331 701
rect 335 697 336 701
rect 330 696 336 697
rect 434 701 440 702
rect 434 697 435 701
rect 439 697 440 701
rect 490 699 491 703
rect 495 702 496 703
rect 495 700 529 702
rect 538 701 544 702
rect 495 699 496 700
rect 490 698 496 699
rect 434 696 440 697
rect 538 697 539 701
rect 543 697 544 701
rect 538 696 544 697
rect 642 701 648 702
rect 642 697 643 701
rect 647 697 648 701
rect 642 696 648 697
rect 722 701 728 702
rect 722 697 723 701
rect 727 697 728 701
rect 722 696 728 697
rect 110 693 116 694
rect 110 689 111 693
rect 115 689 116 693
rect 110 688 116 689
rect 774 693 780 694
rect 774 689 775 693
rect 779 689 780 693
rect 774 688 780 689
rect 110 675 116 676
rect 110 671 111 675
rect 115 671 116 675
rect 478 675 484 676
rect 478 674 479 675
rect 233 672 321 674
rect 337 672 430 674
rect 441 672 479 674
rect 110 670 116 671
rect 198 663 204 664
rect 198 659 199 663
rect 203 662 204 663
rect 233 663 239 664
rect 233 662 234 663
rect 203 660 234 662
rect 203 659 204 660
rect 198 658 204 659
rect 233 659 234 660
rect 238 659 239 663
rect 233 658 239 659
rect 250 663 256 664
rect 250 659 251 663
rect 255 659 256 663
rect 319 662 321 672
rect 337 663 343 664
rect 337 662 338 663
rect 319 660 338 662
rect 250 658 256 659
rect 337 659 338 660
rect 342 659 343 663
rect 337 658 343 659
rect 354 663 360 664
rect 354 659 355 663
rect 359 659 360 663
rect 428 662 430 672
rect 478 671 479 672
rect 483 671 484 675
rect 734 675 740 676
rect 734 674 735 675
rect 649 672 718 674
rect 729 672 735 674
rect 478 670 484 671
rect 441 663 447 664
rect 441 662 442 663
rect 428 660 442 662
rect 354 658 360 659
rect 441 659 442 660
rect 446 659 447 663
rect 441 658 447 659
rect 458 663 464 664
rect 458 659 459 663
rect 463 659 464 663
rect 458 658 464 659
rect 546 663 556 664
rect 546 659 547 663
rect 555 659 556 663
rect 546 658 556 659
rect 562 663 568 664
rect 562 659 563 663
rect 567 659 568 663
rect 562 658 568 659
rect 650 663 656 664
rect 650 659 651 663
rect 655 659 656 663
rect 650 658 656 659
rect 666 663 672 664
rect 666 659 667 663
rect 671 659 672 663
rect 716 662 718 672
rect 734 671 735 672
rect 739 671 740 675
rect 734 670 740 671
rect 774 675 780 676
rect 774 671 775 675
rect 779 671 780 675
rect 774 670 780 671
rect 729 663 735 664
rect 729 662 730 663
rect 716 660 730 662
rect 666 658 672 659
rect 729 659 730 660
rect 734 659 735 663
rect 729 658 735 659
rect 746 663 752 664
rect 746 659 747 663
rect 751 659 752 663
rect 746 658 752 659
rect 478 651 487 652
rect 306 649 312 650
rect 289 647 295 648
rect 289 643 290 647
rect 294 646 295 647
rect 294 644 302 646
rect 306 645 307 649
rect 311 645 312 649
rect 362 649 368 650
rect 306 644 312 645
rect 345 647 351 648
rect 294 643 295 644
rect 289 642 295 643
rect 300 642 302 644
rect 345 643 346 647
rect 350 646 351 647
rect 350 644 358 646
rect 362 645 363 649
rect 367 645 368 649
rect 426 649 432 650
rect 362 644 368 645
rect 409 647 415 648
rect 350 643 351 644
rect 345 642 351 643
rect 356 642 358 644
rect 409 643 410 647
rect 414 646 415 647
rect 414 644 422 646
rect 426 645 427 649
rect 431 645 432 649
rect 478 647 479 651
rect 486 647 487 651
rect 729 651 740 652
rect 478 646 487 647
rect 498 649 504 650
rect 426 644 432 645
rect 498 645 499 649
rect 503 645 504 649
rect 578 649 584 650
rect 498 644 504 645
rect 561 647 567 648
rect 414 643 415 644
rect 409 642 415 643
rect 420 642 422 644
rect 561 643 562 647
rect 566 646 567 647
rect 566 644 574 646
rect 578 645 579 649
rect 583 645 584 649
rect 666 649 672 650
rect 578 644 584 645
rect 630 647 636 648
rect 566 643 567 644
rect 561 642 567 643
rect 300 640 338 642
rect 356 640 402 642
rect 420 640 474 642
rect 110 637 116 638
rect 336 637 338 640
rect 400 637 402 640
rect 472 637 474 640
rect 550 639 556 640
rect 110 633 111 637
rect 115 633 116 637
rect 294 635 300 636
rect 294 634 295 635
rect 110 632 116 633
rect 289 632 295 634
rect 294 631 295 632
rect 299 631 300 635
rect 550 635 551 639
rect 555 635 556 639
rect 550 634 556 635
rect 572 634 574 644
rect 630 643 631 647
rect 635 646 636 647
rect 649 647 655 648
rect 649 646 650 647
rect 635 644 650 646
rect 635 643 636 644
rect 630 642 636 643
rect 649 643 650 644
rect 654 643 655 647
rect 666 645 667 649
rect 671 645 672 649
rect 729 647 730 651
rect 734 647 735 651
rect 739 647 740 651
rect 729 646 740 647
rect 746 649 752 650
rect 666 644 672 645
rect 746 645 747 649
rect 751 645 752 649
rect 746 644 752 645
rect 649 642 655 643
rect 774 637 780 638
rect 572 632 641 634
rect 774 633 775 637
rect 779 633 780 637
rect 774 632 780 633
rect 294 630 300 631
rect 110 619 116 620
rect 110 615 111 619
rect 115 615 116 619
rect 110 614 116 615
rect 774 619 780 620
rect 774 615 775 619
rect 779 615 780 619
rect 774 614 780 615
rect 282 611 288 612
rect 282 607 283 611
rect 287 607 288 611
rect 282 606 288 607
rect 338 611 344 612
rect 338 607 339 611
rect 343 607 344 611
rect 338 606 344 607
rect 402 611 408 612
rect 402 607 403 611
rect 407 607 408 611
rect 402 606 408 607
rect 474 611 480 612
rect 474 607 475 611
rect 479 607 480 611
rect 474 606 480 607
rect 554 611 560 612
rect 554 607 555 611
rect 559 607 560 611
rect 554 606 560 607
rect 642 611 648 612
rect 642 607 643 611
rect 647 607 648 611
rect 642 606 648 607
rect 703 611 709 612
rect 703 607 704 611
rect 708 610 709 611
rect 722 611 728 612
rect 708 608 713 610
rect 708 607 709 608
rect 703 606 709 607
rect 722 607 723 611
rect 727 607 728 611
rect 722 606 728 607
rect 630 603 636 604
rect 346 601 352 602
rect 346 597 347 601
rect 351 597 352 601
rect 346 596 352 597
rect 410 601 416 602
rect 410 597 411 601
rect 415 597 416 601
rect 410 596 416 597
rect 482 601 488 602
rect 482 597 483 601
rect 487 597 488 601
rect 482 596 488 597
rect 562 601 568 602
rect 562 597 563 601
rect 567 597 568 601
rect 630 599 631 603
rect 635 602 636 603
rect 635 600 641 602
rect 650 601 656 602
rect 635 599 636 600
rect 630 598 636 599
rect 562 596 568 597
rect 650 597 651 601
rect 655 597 656 601
rect 650 596 656 597
rect 722 601 728 602
rect 722 597 723 601
rect 727 597 728 601
rect 722 596 728 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 110 588 116 589
rect 774 593 780 594
rect 774 589 775 593
rect 779 589 780 593
rect 774 588 780 589
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 562 575 568 576
rect 353 572 406 574
rect 417 572 478 574
rect 489 572 558 574
rect 110 570 116 571
rect 294 563 300 564
rect 294 559 295 563
rect 299 562 300 563
rect 353 563 359 564
rect 353 562 354 563
rect 299 560 354 562
rect 299 559 300 560
rect 294 558 300 559
rect 353 559 354 560
rect 358 559 359 563
rect 353 558 359 559
rect 370 563 376 564
rect 370 559 371 563
rect 375 559 376 563
rect 404 562 406 572
rect 417 563 423 564
rect 417 562 418 563
rect 404 560 418 562
rect 370 558 376 559
rect 417 559 418 560
rect 422 559 423 563
rect 417 558 423 559
rect 434 563 440 564
rect 434 559 435 563
rect 439 559 440 563
rect 476 562 478 572
rect 489 563 495 564
rect 489 562 490 563
rect 476 560 490 562
rect 434 558 440 559
rect 489 559 490 560
rect 494 559 495 563
rect 489 558 495 559
rect 506 563 512 564
rect 506 559 507 563
rect 511 559 512 563
rect 556 562 558 572
rect 562 571 563 575
rect 567 571 568 575
rect 734 575 740 576
rect 734 574 735 575
rect 729 572 735 574
rect 562 570 568 571
rect 734 571 735 572
rect 739 571 740 575
rect 734 570 740 571
rect 774 575 780 576
rect 774 571 775 575
rect 779 571 780 575
rect 774 570 780 571
rect 569 563 575 564
rect 569 562 570 563
rect 556 560 570 562
rect 506 558 512 559
rect 569 559 570 560
rect 574 559 575 563
rect 569 558 575 559
rect 586 563 592 564
rect 586 559 587 563
rect 591 559 592 563
rect 586 558 592 559
rect 646 563 652 564
rect 646 559 647 563
rect 651 562 652 563
rect 657 563 663 564
rect 657 562 658 563
rect 651 560 658 562
rect 651 559 652 560
rect 646 558 652 559
rect 657 559 658 560
rect 662 559 663 563
rect 657 558 663 559
rect 674 563 680 564
rect 674 559 675 563
rect 679 559 680 563
rect 674 558 680 559
rect 703 563 709 564
rect 703 559 704 563
rect 708 562 709 563
rect 729 563 735 564
rect 729 562 730 563
rect 708 560 730 562
rect 708 559 709 560
rect 703 558 709 559
rect 729 559 730 560
rect 734 559 735 563
rect 729 558 735 559
rect 746 563 752 564
rect 746 559 747 563
rect 751 559 752 563
rect 746 558 752 559
rect 561 555 568 556
rect 346 553 352 554
rect 329 551 335 552
rect 329 547 330 551
rect 334 550 335 551
rect 334 548 342 550
rect 346 549 347 553
rect 351 549 352 553
rect 418 553 424 554
rect 346 548 352 549
rect 401 551 407 552
rect 334 547 335 548
rect 329 546 335 547
rect 340 546 342 548
rect 401 547 402 551
rect 406 550 407 551
rect 406 548 414 550
rect 418 549 419 553
rect 423 549 424 553
rect 498 553 504 554
rect 418 548 424 549
rect 481 551 487 552
rect 406 547 407 548
rect 401 546 407 547
rect 412 546 414 548
rect 481 547 482 551
rect 486 550 487 551
rect 486 548 494 550
rect 498 549 499 553
rect 503 549 504 553
rect 561 551 562 555
rect 567 551 568 555
rect 729 555 740 556
rect 561 550 568 551
rect 578 553 584 554
rect 498 548 504 549
rect 578 549 579 553
rect 583 549 584 553
rect 666 553 672 554
rect 578 548 584 549
rect 591 551 597 552
rect 486 547 487 548
rect 481 546 487 547
rect 492 546 494 548
rect 591 547 592 551
rect 596 550 597 551
rect 649 551 655 552
rect 649 550 650 551
rect 596 548 650 550
rect 596 547 597 548
rect 591 546 597 547
rect 649 547 650 548
rect 654 547 655 551
rect 666 549 667 553
rect 671 549 672 553
rect 729 551 730 555
rect 734 551 735 555
rect 739 551 740 555
rect 729 550 740 551
rect 746 553 752 554
rect 666 548 672 549
rect 746 549 747 553
rect 751 549 752 553
rect 746 548 752 549
rect 649 546 655 547
rect 340 544 394 546
rect 412 544 474 546
rect 492 544 554 546
rect 110 541 116 542
rect 392 541 394 544
rect 472 541 474 544
rect 552 541 554 544
rect 646 543 652 544
rect 110 537 111 541
rect 115 537 116 541
rect 646 539 647 543
rect 651 539 652 543
rect 646 538 652 539
rect 774 541 780 542
rect 774 537 775 541
rect 779 537 780 541
rect 110 536 116 537
rect 328 534 330 537
rect 774 536 780 537
rect 527 535 533 536
rect 527 534 528 535
rect 328 532 528 534
rect 527 531 528 532
rect 532 531 533 535
rect 527 530 533 531
rect 110 523 116 524
rect 110 519 111 523
rect 115 519 116 523
rect 110 518 116 519
rect 774 523 780 524
rect 774 519 775 523
rect 779 519 780 523
rect 774 518 780 519
rect 322 515 328 516
rect 322 511 323 515
rect 327 511 328 515
rect 322 510 328 511
rect 394 515 400 516
rect 394 511 395 515
rect 399 511 400 515
rect 394 510 400 511
rect 474 515 480 516
rect 474 511 475 515
rect 479 511 480 515
rect 474 510 480 511
rect 554 515 560 516
rect 554 511 555 515
rect 559 511 560 515
rect 554 510 560 511
rect 642 515 648 516
rect 642 511 643 515
rect 647 511 648 515
rect 642 510 648 511
rect 703 515 709 516
rect 703 511 704 515
rect 708 514 709 515
rect 722 515 728 516
rect 708 512 713 514
rect 708 511 709 512
rect 703 510 709 511
rect 722 511 723 515
rect 727 511 728 515
rect 722 510 728 511
rect 194 505 200 506
rect 194 501 195 505
rect 199 501 200 505
rect 194 500 200 501
rect 282 505 288 506
rect 282 501 283 505
rect 287 501 288 505
rect 282 500 288 501
rect 378 505 384 506
rect 378 501 379 505
rect 383 501 384 505
rect 378 500 384 501
rect 490 505 496 506
rect 490 501 491 505
rect 495 501 496 505
rect 490 500 496 501
rect 610 505 616 506
rect 610 501 611 505
rect 615 501 616 505
rect 610 500 616 501
rect 722 505 728 506
rect 722 501 723 505
rect 727 501 728 505
rect 722 500 728 501
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 110 492 116 493
rect 774 497 780 498
rect 774 493 775 497
rect 779 493 780 497
rect 774 492 780 493
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 194 479 200 480
rect 194 475 195 479
rect 199 475 200 479
rect 650 479 656 480
rect 194 474 200 475
rect 208 476 281 478
rect 300 476 377 478
rect 392 476 489 478
rect 504 476 609 478
rect 208 468 210 476
rect 202 467 210 468
rect 202 463 203 467
rect 207 464 210 467
rect 218 467 224 468
rect 207 463 208 464
rect 202 462 208 463
rect 218 463 219 467
rect 223 463 224 467
rect 218 462 224 463
rect 290 467 296 468
rect 290 463 291 467
rect 295 466 296 467
rect 300 466 302 476
rect 392 468 394 476
rect 504 468 506 476
rect 650 475 651 479
rect 655 478 656 479
rect 774 479 780 480
rect 655 476 721 478
rect 655 475 656 476
rect 650 474 656 475
rect 774 475 775 479
rect 779 475 780 479
rect 774 474 780 475
rect 295 464 302 466
rect 306 467 312 468
rect 295 463 296 464
rect 290 462 296 463
rect 306 463 307 467
rect 311 463 312 467
rect 306 462 312 463
rect 386 467 394 468
rect 386 463 387 467
rect 391 464 394 467
rect 402 467 408 468
rect 391 463 392 464
rect 386 462 392 463
rect 402 463 403 467
rect 407 463 408 467
rect 402 462 408 463
rect 498 467 506 468
rect 498 463 499 467
rect 503 464 506 467
rect 514 467 520 468
rect 503 463 504 464
rect 498 462 504 463
rect 514 463 515 467
rect 519 463 520 467
rect 514 462 520 463
rect 527 467 533 468
rect 527 463 528 467
rect 532 466 533 467
rect 617 467 623 468
rect 617 466 618 467
rect 532 464 618 466
rect 532 463 533 464
rect 527 462 533 463
rect 617 463 618 464
rect 622 463 623 467
rect 617 462 623 463
rect 634 467 640 468
rect 634 463 635 467
rect 639 463 640 467
rect 634 462 640 463
rect 703 467 709 468
rect 703 463 704 467
rect 708 466 709 467
rect 729 467 735 468
rect 729 466 730 467
rect 708 464 730 466
rect 708 463 709 464
rect 703 462 709 463
rect 729 463 730 464
rect 734 463 735 467
rect 729 462 735 463
rect 746 467 752 468
rect 746 463 747 467
rect 751 463 752 467
rect 746 462 752 463
rect 194 459 200 460
rect 194 455 195 459
rect 199 458 200 459
rect 199 456 398 458
rect 199 455 200 456
rect 194 454 200 455
rect 396 454 398 456
rect 457 455 463 456
rect 457 454 458 455
rect 170 453 176 454
rect 153 451 159 452
rect 153 447 154 451
rect 158 450 159 451
rect 158 448 166 450
rect 170 449 171 453
rect 175 449 176 453
rect 226 453 232 454
rect 170 448 176 449
rect 209 451 215 452
rect 158 447 159 448
rect 153 446 159 447
rect 164 446 166 448
rect 209 447 210 451
rect 214 450 215 451
rect 214 448 222 450
rect 226 449 227 453
rect 231 449 232 453
rect 298 453 304 454
rect 226 448 232 449
rect 281 451 287 452
rect 214 447 215 448
rect 209 446 215 447
rect 220 446 222 448
rect 281 447 282 451
rect 286 450 287 451
rect 286 448 294 450
rect 298 449 299 453
rect 303 449 304 453
rect 386 453 392 454
rect 298 448 304 449
rect 369 451 375 452
rect 286 447 287 448
rect 281 446 287 447
rect 292 446 294 448
rect 369 447 370 451
rect 374 450 375 451
rect 374 448 382 450
rect 386 449 387 453
rect 391 449 392 453
rect 396 452 458 454
rect 457 451 458 452
rect 462 451 463 455
rect 649 455 656 456
rect 457 450 463 451
rect 474 453 480 454
rect 386 448 392 449
rect 474 449 475 453
rect 479 449 480 453
rect 570 453 576 454
rect 474 448 480 449
rect 553 451 559 452
rect 374 447 375 448
rect 369 446 375 447
rect 380 446 382 448
rect 553 447 554 451
rect 558 450 559 451
rect 562 451 568 452
rect 562 450 563 451
rect 558 448 563 450
rect 558 447 559 448
rect 553 446 559 447
rect 562 447 563 448
rect 567 447 568 451
rect 570 449 571 453
rect 575 449 576 453
rect 649 451 650 455
rect 655 451 656 455
rect 649 450 656 451
rect 666 453 672 454
rect 570 448 576 449
rect 666 449 667 453
rect 671 449 672 453
rect 746 453 752 454
rect 729 451 735 452
rect 729 450 730 451
rect 666 448 672 449
rect 680 448 730 450
rect 562 446 568 447
rect 164 444 202 446
rect 220 444 274 446
rect 292 444 362 446
rect 380 444 450 446
rect 110 441 116 442
rect 200 441 202 444
rect 272 441 274 444
rect 360 441 362 444
rect 448 441 450 444
rect 591 443 597 444
rect 591 442 592 443
rect 110 437 111 441
rect 115 437 116 441
rect 553 440 592 442
rect 591 439 592 440
rect 596 439 597 443
rect 680 442 682 448
rect 729 447 730 448
rect 734 447 735 451
rect 746 449 747 453
rect 751 449 752 453
rect 746 448 752 449
rect 729 446 735 447
rect 649 440 682 442
rect 774 441 780 442
rect 591 438 597 439
rect 110 436 116 437
rect 774 437 775 441
rect 779 437 780 441
rect 774 436 780 437
rect 110 423 116 424
rect 110 419 111 423
rect 115 419 116 423
rect 110 418 116 419
rect 774 423 780 424
rect 774 419 775 423
rect 779 419 780 423
rect 774 418 780 419
rect 127 415 133 416
rect 127 411 128 415
rect 132 414 133 415
rect 146 415 152 416
rect 132 412 137 414
rect 132 411 133 412
rect 127 410 133 411
rect 146 411 147 415
rect 151 411 152 415
rect 146 410 152 411
rect 202 415 208 416
rect 202 411 203 415
rect 207 411 208 415
rect 202 410 208 411
rect 274 415 280 416
rect 274 411 275 415
rect 279 411 280 415
rect 274 410 280 411
rect 362 415 368 416
rect 362 411 363 415
rect 367 411 368 415
rect 362 410 368 411
rect 450 415 456 416
rect 450 411 451 415
rect 455 411 456 415
rect 450 410 456 411
rect 546 415 552 416
rect 546 411 547 415
rect 551 411 552 415
rect 546 410 552 411
rect 642 415 648 416
rect 642 411 643 415
rect 647 411 648 415
rect 642 410 648 411
rect 703 415 709 416
rect 703 411 704 415
rect 708 414 709 415
rect 722 415 728 416
rect 708 412 713 414
rect 708 411 709 412
rect 703 410 709 411
rect 722 411 723 415
rect 727 411 728 415
rect 722 410 728 411
rect 562 399 568 400
rect 146 397 152 398
rect 146 393 147 397
rect 151 393 152 397
rect 146 392 152 393
rect 226 397 232 398
rect 226 393 227 397
rect 231 393 232 397
rect 226 392 232 393
rect 314 397 320 398
rect 314 393 315 397
rect 319 393 320 397
rect 314 392 320 393
rect 410 397 416 398
rect 410 393 411 397
rect 415 393 416 397
rect 410 392 416 393
rect 514 397 520 398
rect 514 393 515 397
rect 519 393 520 397
rect 562 395 563 399
rect 567 398 568 399
rect 567 396 617 398
rect 626 397 632 398
rect 567 395 568 396
rect 562 394 568 395
rect 514 392 520 393
rect 626 393 627 397
rect 631 393 632 397
rect 626 392 632 393
rect 722 397 728 398
rect 722 393 723 397
rect 727 393 728 397
rect 722 392 728 393
rect 110 389 116 390
rect 110 385 111 389
rect 115 385 116 389
rect 110 384 116 385
rect 774 389 780 390
rect 774 385 775 389
rect 779 385 780 389
rect 774 384 780 385
rect 110 371 116 372
rect 110 367 111 371
rect 115 367 116 371
rect 530 371 536 372
rect 530 370 531 371
rect 153 368 222 370
rect 233 368 310 370
rect 321 368 370 370
rect 417 368 510 370
rect 521 368 531 370
rect 110 366 116 367
rect 127 359 133 360
rect 127 355 128 359
rect 132 358 133 359
rect 153 359 159 360
rect 153 358 154 359
rect 132 356 154 358
rect 132 355 133 356
rect 127 354 133 355
rect 153 355 154 356
rect 158 355 159 359
rect 153 354 159 355
rect 170 359 176 360
rect 170 355 171 359
rect 175 355 176 359
rect 220 358 222 368
rect 233 359 239 360
rect 233 358 234 359
rect 220 356 234 358
rect 170 354 176 355
rect 233 355 234 356
rect 238 355 239 359
rect 233 354 239 355
rect 250 359 256 360
rect 250 355 251 359
rect 255 355 256 359
rect 308 358 310 368
rect 321 359 327 360
rect 321 358 322 359
rect 308 356 322 358
rect 250 354 256 355
rect 321 355 322 356
rect 326 355 327 359
rect 321 354 327 355
rect 338 359 344 360
rect 338 355 339 359
rect 343 355 344 359
rect 368 358 370 368
rect 417 359 423 360
rect 417 358 418 359
rect 368 356 418 358
rect 338 354 344 355
rect 417 355 418 356
rect 422 355 423 359
rect 417 354 423 355
rect 434 359 440 360
rect 434 355 435 359
rect 439 355 440 359
rect 508 358 510 368
rect 530 367 531 368
rect 535 367 536 371
rect 530 366 536 367
rect 674 371 680 372
rect 674 367 675 371
rect 679 370 680 371
rect 774 371 780 372
rect 679 368 721 370
rect 679 367 680 368
rect 674 366 680 367
rect 774 367 775 371
rect 779 367 780 371
rect 774 366 780 367
rect 521 359 527 360
rect 521 358 522 359
rect 508 356 522 358
rect 434 354 440 355
rect 521 355 522 356
rect 526 355 527 359
rect 521 354 527 355
rect 538 359 544 360
rect 538 355 539 359
rect 543 355 544 359
rect 538 354 544 355
rect 606 359 612 360
rect 606 355 607 359
rect 611 358 612 359
rect 633 359 639 360
rect 633 358 634 359
rect 611 356 634 358
rect 611 355 612 356
rect 606 354 612 355
rect 633 355 634 356
rect 638 355 639 359
rect 633 354 639 355
rect 650 359 656 360
rect 650 355 651 359
rect 655 355 656 359
rect 650 354 656 355
rect 703 359 709 360
rect 703 355 704 359
rect 708 358 709 359
rect 729 359 735 360
rect 729 358 730 359
rect 708 356 730 358
rect 708 355 709 356
rect 703 354 709 355
rect 729 355 730 356
rect 734 355 735 359
rect 729 354 735 355
rect 746 359 752 360
rect 746 355 747 359
rect 751 355 752 359
rect 746 354 752 355
rect 530 351 536 352
rect 314 349 320 350
rect 297 347 303 348
rect 297 343 298 347
rect 302 346 303 347
rect 302 344 310 346
rect 314 345 315 349
rect 319 345 320 349
rect 370 349 376 350
rect 314 344 320 345
rect 353 347 359 348
rect 302 343 303 344
rect 297 342 303 343
rect 308 342 310 344
rect 353 343 354 347
rect 358 346 359 347
rect 358 344 366 346
rect 370 345 371 349
rect 375 345 376 349
rect 434 349 440 350
rect 370 344 376 345
rect 417 347 423 348
rect 358 343 359 344
rect 353 342 359 343
rect 364 342 366 344
rect 417 343 418 347
rect 422 346 423 347
rect 422 344 430 346
rect 434 345 435 349
rect 439 345 440 349
rect 498 349 504 350
rect 434 344 440 345
rect 481 347 487 348
rect 422 343 423 344
rect 417 342 423 343
rect 428 342 430 344
rect 481 343 482 347
rect 486 346 487 347
rect 486 344 494 346
rect 498 345 499 349
rect 503 345 504 349
rect 530 347 531 351
rect 535 350 536 351
rect 545 351 551 352
rect 545 350 546 351
rect 535 348 546 350
rect 535 347 536 348
rect 530 346 536 347
rect 545 347 546 348
rect 550 347 551 351
rect 673 351 680 352
rect 545 346 551 347
rect 562 349 568 350
rect 498 344 504 345
rect 562 345 563 349
rect 567 345 568 349
rect 626 349 632 350
rect 562 344 568 345
rect 570 347 576 348
rect 486 343 487 344
rect 481 342 487 343
rect 492 342 494 344
rect 570 343 571 347
rect 575 346 576 347
rect 609 347 615 348
rect 609 346 610 347
rect 575 344 610 346
rect 575 343 576 344
rect 570 342 576 343
rect 609 343 610 344
rect 614 343 615 347
rect 626 345 627 349
rect 631 345 632 349
rect 673 347 674 351
rect 679 347 680 351
rect 673 346 680 347
rect 690 349 696 350
rect 626 344 632 345
rect 690 345 691 349
rect 695 345 696 349
rect 746 349 752 350
rect 729 347 735 348
rect 729 346 730 347
rect 690 344 696 345
rect 700 344 730 346
rect 609 342 615 343
rect 308 340 346 342
rect 364 340 410 342
rect 428 340 474 342
rect 492 340 538 342
rect 110 337 116 338
rect 344 337 346 340
rect 408 337 410 340
rect 472 337 474 340
rect 536 337 538 340
rect 606 339 612 340
rect 110 333 111 337
rect 115 333 116 337
rect 606 335 607 339
rect 611 335 612 339
rect 700 338 702 344
rect 729 343 730 344
rect 734 343 735 347
rect 746 345 747 349
rect 751 345 752 349
rect 746 344 752 345
rect 729 342 735 343
rect 673 336 702 338
rect 774 337 780 338
rect 606 334 612 335
rect 110 332 116 333
rect 297 332 321 334
rect 774 333 775 337
rect 779 333 780 337
rect 774 332 780 333
rect 319 330 321 332
rect 434 331 440 332
rect 434 330 435 331
rect 319 328 435 330
rect 434 327 435 328
rect 439 327 440 331
rect 434 326 440 327
rect 110 319 116 320
rect 110 315 111 319
rect 115 315 116 319
rect 110 314 116 315
rect 774 319 780 320
rect 774 315 775 319
rect 779 315 780 319
rect 774 314 780 315
rect 290 311 296 312
rect 290 307 291 311
rect 295 307 296 311
rect 290 306 296 307
rect 346 311 352 312
rect 346 307 347 311
rect 351 307 352 311
rect 346 306 352 307
rect 410 311 416 312
rect 410 307 411 311
rect 415 307 416 311
rect 410 306 416 307
rect 474 311 480 312
rect 474 307 475 311
rect 479 307 480 311
rect 474 306 480 307
rect 538 311 544 312
rect 538 307 539 311
rect 543 307 544 311
rect 538 306 544 307
rect 602 311 608 312
rect 602 307 603 311
rect 607 307 608 311
rect 602 306 608 307
rect 666 311 672 312
rect 666 307 667 311
rect 671 307 672 311
rect 666 306 672 307
rect 703 311 709 312
rect 703 307 704 311
rect 708 310 709 311
rect 722 311 728 312
rect 708 308 713 310
rect 708 307 709 308
rect 703 306 709 307
rect 722 307 723 311
rect 727 307 728 311
rect 722 306 728 307
rect 218 301 224 302
rect 218 297 219 301
rect 223 297 224 301
rect 218 296 224 297
rect 274 301 280 302
rect 274 297 275 301
rect 279 297 280 301
rect 274 296 280 297
rect 330 301 336 302
rect 330 297 331 301
rect 335 297 336 301
rect 330 296 336 297
rect 386 301 392 302
rect 386 297 387 301
rect 391 297 392 301
rect 386 296 392 297
rect 442 301 448 302
rect 442 297 443 301
rect 447 297 448 301
rect 442 296 448 297
rect 498 301 504 302
rect 498 297 499 301
rect 503 297 504 301
rect 498 296 504 297
rect 554 301 560 302
rect 554 297 555 301
rect 559 297 560 301
rect 554 296 560 297
rect 610 301 616 302
rect 610 297 611 301
rect 615 297 616 301
rect 610 296 616 297
rect 666 301 672 302
rect 666 297 667 301
rect 671 297 672 301
rect 666 296 672 297
rect 722 301 728 302
rect 722 297 723 301
rect 727 297 728 301
rect 722 296 728 297
rect 110 293 116 294
rect 110 289 111 293
rect 115 289 116 293
rect 110 288 116 289
rect 774 293 780 294
rect 774 289 775 293
rect 779 289 780 293
rect 774 288 780 289
rect 570 283 576 284
rect 570 282 571 283
rect 532 280 571 282
rect 532 278 534 280
rect 570 279 571 280
rect 575 279 576 283
rect 570 278 576 279
rect 504 276 534 278
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 110 270 116 271
rect 218 275 224 276
rect 218 271 219 275
rect 223 271 224 275
rect 218 270 224 271
rect 232 272 273 274
rect 292 272 329 274
rect 344 272 385 274
rect 400 272 441 274
rect 504 273 506 276
rect 774 275 780 276
rect 512 272 553 274
rect 568 272 609 274
rect 624 272 665 274
rect 680 272 721 274
rect 232 264 234 272
rect 226 263 234 264
rect 226 259 227 263
rect 231 260 234 263
rect 242 263 248 264
rect 231 259 232 260
rect 226 258 232 259
rect 242 259 243 263
rect 247 259 248 263
rect 242 258 248 259
rect 282 263 288 264
rect 282 259 283 263
rect 287 262 288 263
rect 292 262 294 272
rect 344 264 346 272
rect 400 264 402 272
rect 512 264 514 272
rect 568 264 570 272
rect 624 264 626 272
rect 680 264 682 272
rect 774 271 775 275
rect 779 271 780 275
rect 774 270 780 271
rect 287 260 294 262
rect 298 263 304 264
rect 287 259 288 260
rect 282 258 288 259
rect 298 259 299 263
rect 303 259 304 263
rect 298 258 304 259
rect 338 263 346 264
rect 338 259 339 263
rect 343 260 346 263
rect 354 263 360 264
rect 343 259 344 260
rect 338 258 344 259
rect 354 259 355 263
rect 359 259 360 263
rect 354 258 360 259
rect 394 263 402 264
rect 394 259 395 263
rect 399 260 402 263
rect 410 263 416 264
rect 399 259 400 260
rect 394 258 400 259
rect 410 259 411 263
rect 415 259 416 263
rect 410 258 416 259
rect 434 263 440 264
rect 434 259 435 263
rect 439 262 440 263
rect 449 263 455 264
rect 449 262 450 263
rect 439 260 450 262
rect 439 259 440 260
rect 434 258 440 259
rect 449 259 450 260
rect 454 259 455 263
rect 449 258 455 259
rect 466 263 472 264
rect 466 259 467 263
rect 471 259 472 263
rect 466 258 472 259
rect 506 263 514 264
rect 506 259 507 263
rect 511 260 514 263
rect 522 263 528 264
rect 511 259 512 260
rect 506 258 512 259
rect 522 259 523 263
rect 527 259 528 263
rect 522 258 528 259
rect 562 263 570 264
rect 562 259 563 263
rect 567 260 570 263
rect 578 263 584 264
rect 567 259 568 260
rect 562 258 568 259
rect 578 259 579 263
rect 583 259 584 263
rect 578 258 584 259
rect 618 263 626 264
rect 618 259 619 263
rect 623 260 626 263
rect 634 263 640 264
rect 623 259 624 260
rect 618 258 624 259
rect 634 259 635 263
rect 639 259 640 263
rect 634 258 640 259
rect 674 263 682 264
rect 674 259 675 263
rect 679 260 682 263
rect 690 263 696 264
rect 679 259 680 260
rect 674 258 680 259
rect 690 259 691 263
rect 695 259 696 263
rect 690 258 696 259
rect 703 263 709 264
rect 703 259 704 263
rect 708 262 709 263
rect 729 263 735 264
rect 729 262 730 263
rect 708 260 730 262
rect 708 259 709 260
rect 703 258 709 259
rect 729 259 730 260
rect 734 259 735 263
rect 729 258 735 259
rect 746 263 752 264
rect 746 259 747 263
rect 751 259 752 263
rect 746 258 752 259
rect 218 247 224 248
rect 218 243 219 247
rect 223 246 224 247
rect 223 244 486 246
rect 223 243 224 244
rect 218 242 224 243
rect 484 242 486 244
rect 513 243 519 244
rect 513 242 514 243
rect 306 241 312 242
rect 289 239 295 240
rect 289 235 290 239
rect 294 238 295 239
rect 294 236 302 238
rect 306 237 307 241
rect 311 237 312 241
rect 362 241 368 242
rect 306 236 312 237
rect 345 239 351 240
rect 294 235 295 236
rect 289 234 295 235
rect 300 234 302 236
rect 345 235 346 239
rect 350 238 351 239
rect 350 236 358 238
rect 362 237 363 241
rect 367 237 368 241
rect 418 241 424 242
rect 362 236 368 237
rect 401 239 407 240
rect 350 235 351 236
rect 345 234 351 235
rect 356 234 358 236
rect 401 235 402 239
rect 406 238 407 239
rect 406 236 414 238
rect 418 237 419 241
rect 423 237 424 241
rect 474 241 480 242
rect 418 236 424 237
rect 457 239 463 240
rect 406 235 407 236
rect 401 234 407 235
rect 412 234 414 236
rect 457 235 458 239
rect 462 238 463 239
rect 462 236 470 238
rect 474 237 475 241
rect 479 237 480 241
rect 484 240 514 242
rect 513 239 514 240
rect 518 239 519 243
rect 513 238 519 239
rect 530 241 536 242
rect 474 236 480 237
rect 530 237 531 241
rect 535 237 536 241
rect 530 236 536 237
rect 462 235 463 236
rect 457 234 463 235
rect 468 234 470 236
rect 300 232 338 234
rect 356 232 394 234
rect 412 232 450 234
rect 468 232 506 234
rect 110 229 116 230
rect 336 229 338 232
rect 392 229 394 232
rect 448 229 450 232
rect 504 229 506 232
rect 774 229 780 230
rect 110 225 111 229
rect 115 225 116 229
rect 774 225 775 229
rect 779 225 780 229
rect 110 224 116 225
rect 288 222 290 225
rect 774 224 780 225
rect 362 223 368 224
rect 362 222 363 223
rect 288 220 363 222
rect 362 219 363 220
rect 367 219 368 223
rect 362 218 368 219
rect 110 211 116 212
rect 110 207 111 211
rect 115 207 116 211
rect 110 206 116 207
rect 774 211 780 212
rect 774 207 775 211
rect 779 207 780 211
rect 774 206 780 207
rect 282 203 288 204
rect 282 199 283 203
rect 287 199 288 203
rect 282 198 288 199
rect 338 203 344 204
rect 338 199 339 203
rect 343 199 344 203
rect 338 198 344 199
rect 394 203 400 204
rect 394 199 395 203
rect 399 199 400 203
rect 394 198 400 199
rect 450 203 456 204
rect 450 199 451 203
rect 455 199 456 203
rect 450 198 456 199
rect 506 203 512 204
rect 506 199 507 203
rect 511 199 512 203
rect 506 198 512 199
rect 162 189 168 190
rect 162 185 163 189
rect 167 185 168 189
rect 162 184 168 185
rect 218 189 224 190
rect 218 185 219 189
rect 223 185 224 189
rect 218 184 224 185
rect 274 189 280 190
rect 274 185 275 189
rect 279 185 280 189
rect 274 184 280 185
rect 330 189 336 190
rect 330 185 331 189
rect 335 185 336 189
rect 330 184 336 185
rect 386 189 392 190
rect 386 185 387 189
rect 391 185 392 189
rect 386 184 392 185
rect 110 181 116 182
rect 110 177 111 181
rect 115 177 116 181
rect 110 176 116 177
rect 774 181 780 182
rect 774 177 775 181
rect 779 177 780 181
rect 774 176 780 177
rect 110 163 116 164
rect 110 159 111 163
rect 115 159 116 163
rect 110 158 116 159
rect 162 163 168 164
rect 162 159 163 163
rect 167 159 168 163
rect 774 163 780 164
rect 162 158 168 159
rect 176 160 217 162
rect 232 160 273 162
rect 292 160 329 162
rect 344 160 385 162
rect 176 152 178 160
rect 232 152 234 160
rect 170 151 178 152
rect 170 147 171 151
rect 175 148 178 151
rect 186 151 192 152
rect 175 147 176 148
rect 170 146 176 147
rect 186 147 187 151
rect 191 147 192 151
rect 186 146 192 147
rect 226 151 234 152
rect 226 147 227 151
rect 231 148 234 151
rect 242 151 248 152
rect 231 147 232 148
rect 226 146 232 147
rect 242 147 243 151
rect 247 147 248 151
rect 242 146 248 147
rect 282 151 288 152
rect 282 147 283 151
rect 287 150 288 151
rect 292 150 294 160
rect 344 152 346 160
rect 774 159 775 163
rect 779 159 780 163
rect 774 158 780 159
rect 287 148 294 150
rect 298 151 304 152
rect 287 147 288 148
rect 282 146 288 147
rect 298 147 299 151
rect 303 147 304 151
rect 298 146 304 147
rect 338 151 346 152
rect 338 147 339 151
rect 343 148 346 151
rect 354 151 360 152
rect 343 147 344 148
rect 338 146 344 147
rect 354 147 355 151
rect 359 147 360 151
rect 354 146 360 147
rect 362 151 368 152
rect 362 147 363 151
rect 367 150 368 151
rect 393 151 399 152
rect 393 150 394 151
rect 367 148 394 150
rect 367 147 368 148
rect 362 146 368 147
rect 393 147 394 148
rect 398 147 399 151
rect 393 146 399 147
rect 410 151 416 152
rect 410 147 411 151
rect 415 147 416 151
rect 410 146 416 147
rect 542 131 551 132
rect 170 129 176 130
rect 153 127 159 128
rect 153 123 154 127
rect 158 126 159 127
rect 158 124 166 126
rect 170 125 171 129
rect 175 125 176 129
rect 226 129 232 130
rect 170 124 176 125
rect 209 127 215 128
rect 158 123 159 124
rect 153 122 159 123
rect 164 122 166 124
rect 209 123 210 127
rect 214 126 215 127
rect 214 124 222 126
rect 226 125 227 129
rect 231 125 232 129
rect 282 129 288 130
rect 226 124 232 125
rect 265 127 271 128
rect 214 123 215 124
rect 209 122 215 123
rect 220 122 222 124
rect 265 123 266 127
rect 270 126 271 127
rect 270 124 278 126
rect 282 125 283 129
rect 287 125 288 129
rect 338 129 344 130
rect 282 124 288 125
rect 321 127 327 128
rect 270 123 271 124
rect 265 122 271 123
rect 276 122 278 124
rect 321 123 322 127
rect 326 126 327 127
rect 326 124 334 126
rect 338 125 339 129
rect 343 125 344 129
rect 394 129 400 130
rect 338 124 344 125
rect 377 127 383 128
rect 326 123 327 124
rect 321 122 327 123
rect 332 122 334 124
rect 377 123 378 127
rect 382 126 383 127
rect 382 124 390 126
rect 394 125 395 129
rect 399 125 400 129
rect 450 129 456 130
rect 394 124 400 125
rect 433 127 439 128
rect 382 123 383 124
rect 377 122 383 123
rect 388 122 390 124
rect 433 123 434 127
rect 438 126 439 127
rect 438 124 446 126
rect 450 125 451 129
rect 455 125 456 129
rect 506 129 512 130
rect 450 124 456 125
rect 489 127 495 128
rect 438 123 439 124
rect 433 122 439 123
rect 444 122 446 124
rect 489 123 490 127
rect 494 126 495 127
rect 494 124 502 126
rect 506 125 507 129
rect 511 125 512 129
rect 542 127 543 131
rect 550 127 551 131
rect 542 126 551 127
rect 562 129 568 130
rect 506 124 512 125
rect 562 125 563 129
rect 567 125 568 129
rect 562 124 568 125
rect 494 123 495 124
rect 489 122 495 123
rect 500 122 502 124
rect 164 120 202 122
rect 220 120 258 122
rect 276 120 314 122
rect 332 120 370 122
rect 388 120 426 122
rect 444 120 482 122
rect 500 120 538 122
rect 110 117 116 118
rect 200 117 202 120
rect 256 117 258 120
rect 312 117 314 120
rect 368 117 370 120
rect 424 117 426 120
rect 480 117 482 120
rect 536 117 538 120
rect 774 117 780 118
rect 110 113 111 117
rect 115 113 116 117
rect 110 112 116 113
rect 774 113 775 117
rect 779 113 780 117
rect 774 112 780 113
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 774 99 780 100
rect 774 95 775 99
rect 779 95 780 99
rect 774 94 780 95
rect 146 91 152 92
rect 146 87 147 91
rect 151 87 152 91
rect 146 86 152 87
rect 202 91 208 92
rect 202 87 203 91
rect 207 87 208 91
rect 202 86 208 87
rect 258 91 264 92
rect 258 87 259 91
rect 263 87 264 91
rect 258 86 264 87
rect 314 91 320 92
rect 314 87 315 91
rect 319 87 320 91
rect 314 86 320 87
rect 370 91 376 92
rect 370 87 371 91
rect 375 87 376 91
rect 370 86 376 87
rect 426 91 432 92
rect 426 87 427 91
rect 431 87 432 91
rect 426 86 432 87
rect 482 91 488 92
rect 482 87 483 91
rect 487 87 488 91
rect 482 86 488 87
rect 538 91 544 92
rect 538 87 539 91
rect 543 87 544 91
rect 538 86 544 87
<< m3c >>
rect 195 809 199 813
rect 251 809 255 813
rect 307 809 311 813
rect 363 809 367 813
rect 419 809 423 813
rect 475 809 479 813
rect 539 809 543 813
rect 603 809 607 813
rect 667 809 671 813
rect 723 809 727 813
rect 111 801 115 805
rect 775 801 779 805
rect 111 783 115 787
rect 195 783 199 787
rect 219 771 223 775
rect 275 771 279 775
rect 331 771 335 775
rect 387 771 391 775
rect 443 771 447 775
rect 499 771 503 775
rect 563 771 567 775
rect 575 771 579 775
rect 627 771 631 775
rect 691 771 695 775
rect 735 783 739 787
rect 775 783 779 787
rect 747 771 751 775
rect 195 759 199 763
rect 203 753 207 757
rect 267 753 271 757
rect 339 753 343 757
rect 419 753 423 757
rect 491 751 494 755
rect 494 751 495 755
rect 507 753 511 757
rect 595 753 599 757
rect 683 753 687 757
rect 735 755 739 759
rect 747 753 751 757
rect 111 741 115 745
rect 199 739 203 743
rect 575 743 579 747
rect 775 741 779 745
rect 111 723 115 727
rect 775 723 779 727
rect 179 715 183 719
rect 243 715 247 719
rect 315 715 319 719
rect 395 715 399 719
rect 483 715 487 719
rect 571 715 575 719
rect 659 715 663 719
rect 723 715 727 719
rect 651 707 655 711
rect 227 697 231 701
rect 331 697 335 701
rect 435 697 439 701
rect 491 699 495 703
rect 539 697 543 701
rect 643 697 647 701
rect 723 697 727 701
rect 111 689 115 693
rect 775 689 779 693
rect 111 671 115 675
rect 199 659 203 663
rect 251 659 255 663
rect 355 659 359 663
rect 479 671 483 675
rect 459 659 463 663
rect 551 659 555 663
rect 563 659 567 663
rect 651 659 655 663
rect 667 659 671 663
rect 735 671 739 675
rect 775 671 779 675
rect 747 659 751 663
rect 307 645 311 649
rect 363 645 367 649
rect 427 645 431 649
rect 479 647 482 651
rect 482 647 483 651
rect 499 645 503 649
rect 579 645 583 649
rect 111 633 115 637
rect 295 631 299 635
rect 551 635 555 639
rect 631 643 635 647
rect 667 645 671 649
rect 735 647 739 651
rect 747 645 751 649
rect 775 633 779 637
rect 111 615 115 619
rect 775 615 779 619
rect 283 607 287 611
rect 339 607 343 611
rect 403 607 407 611
rect 475 607 479 611
rect 555 607 559 611
rect 643 607 647 611
rect 723 607 727 611
rect 347 597 351 601
rect 411 597 415 601
rect 483 597 487 601
rect 563 597 567 601
rect 631 599 635 603
rect 651 597 655 601
rect 723 597 727 601
rect 111 589 115 593
rect 775 589 779 593
rect 111 571 115 575
rect 295 559 299 563
rect 371 559 375 563
rect 435 559 439 563
rect 507 559 511 563
rect 563 571 567 575
rect 735 571 739 575
rect 775 571 779 575
rect 587 559 591 563
rect 647 559 651 563
rect 675 559 679 563
rect 747 559 751 563
rect 347 549 351 553
rect 419 549 423 553
rect 499 549 503 553
rect 563 551 566 555
rect 566 551 567 555
rect 579 549 583 553
rect 667 549 671 553
rect 735 551 739 555
rect 747 549 751 553
rect 111 537 115 541
rect 647 539 651 543
rect 775 537 779 541
rect 111 519 115 523
rect 775 519 779 523
rect 323 511 327 515
rect 395 511 399 515
rect 475 511 479 515
rect 555 511 559 515
rect 643 511 647 515
rect 723 511 727 515
rect 195 501 199 505
rect 283 501 287 505
rect 379 501 383 505
rect 491 501 495 505
rect 611 501 615 505
rect 723 501 727 505
rect 111 493 115 497
rect 775 493 779 497
rect 111 475 115 479
rect 195 475 199 479
rect 219 463 223 467
rect 651 475 655 479
rect 775 475 779 479
rect 307 463 311 467
rect 403 463 407 467
rect 515 463 519 467
rect 635 463 639 467
rect 747 463 751 467
rect 195 455 199 459
rect 171 449 175 453
rect 227 449 231 453
rect 299 449 303 453
rect 387 449 391 453
rect 475 449 479 453
rect 563 447 567 451
rect 571 449 575 453
rect 651 451 654 455
rect 654 451 655 455
rect 667 449 671 453
rect 111 437 115 441
rect 747 449 751 453
rect 775 437 779 441
rect 111 419 115 423
rect 775 419 779 423
rect 147 411 151 415
rect 203 411 207 415
rect 275 411 279 415
rect 363 411 367 415
rect 451 411 455 415
rect 547 411 551 415
rect 643 411 647 415
rect 723 411 727 415
rect 147 393 151 397
rect 227 393 231 397
rect 315 393 319 397
rect 411 393 415 397
rect 515 393 519 397
rect 563 395 567 399
rect 627 393 631 397
rect 723 393 727 397
rect 111 385 115 389
rect 775 385 779 389
rect 111 367 115 371
rect 171 355 175 359
rect 251 355 255 359
rect 339 355 343 359
rect 435 355 439 359
rect 531 367 535 371
rect 675 367 679 371
rect 775 367 779 371
rect 539 355 543 359
rect 607 355 611 359
rect 651 355 655 359
rect 747 355 751 359
rect 315 345 319 349
rect 371 345 375 349
rect 435 345 439 349
rect 499 345 503 349
rect 531 347 535 351
rect 563 345 567 349
rect 571 343 575 347
rect 627 345 631 349
rect 675 347 678 351
rect 678 347 679 351
rect 691 345 695 349
rect 111 333 115 337
rect 607 335 611 339
rect 747 345 751 349
rect 775 333 779 337
rect 435 327 439 331
rect 111 315 115 319
rect 775 315 779 319
rect 291 307 295 311
rect 347 307 351 311
rect 411 307 415 311
rect 475 307 479 311
rect 539 307 543 311
rect 603 307 607 311
rect 667 307 671 311
rect 723 307 727 311
rect 219 297 223 301
rect 275 297 279 301
rect 331 297 335 301
rect 387 297 391 301
rect 443 297 447 301
rect 499 297 503 301
rect 555 297 559 301
rect 611 297 615 301
rect 667 297 671 301
rect 723 297 727 301
rect 111 289 115 293
rect 775 289 779 293
rect 571 279 575 283
rect 111 271 115 275
rect 219 271 223 275
rect 243 259 247 263
rect 775 271 779 275
rect 299 259 303 263
rect 355 259 359 263
rect 411 259 415 263
rect 435 259 439 263
rect 467 259 471 263
rect 523 259 527 263
rect 579 259 583 263
rect 635 259 639 263
rect 691 259 695 263
rect 747 259 751 263
rect 219 243 223 247
rect 307 237 311 241
rect 363 237 367 241
rect 419 237 423 241
rect 475 237 479 241
rect 531 237 535 241
rect 111 225 115 229
rect 775 225 779 229
rect 363 219 367 223
rect 111 207 115 211
rect 775 207 779 211
rect 283 199 287 203
rect 339 199 343 203
rect 395 199 399 203
rect 451 199 455 203
rect 507 199 511 203
rect 163 185 167 189
rect 219 185 223 189
rect 275 185 279 189
rect 331 185 335 189
rect 387 185 391 189
rect 111 177 115 181
rect 775 177 779 181
rect 111 159 115 163
rect 163 159 167 163
rect 187 147 191 151
rect 243 147 247 151
rect 775 159 779 163
rect 299 147 303 151
rect 355 147 359 151
rect 363 147 367 151
rect 411 147 415 151
rect 171 125 175 129
rect 227 125 231 129
rect 283 125 287 129
rect 339 125 343 129
rect 395 125 399 129
rect 451 125 455 129
rect 507 125 511 129
rect 543 127 546 131
rect 546 127 547 131
rect 563 125 567 129
rect 111 113 115 117
rect 775 113 779 117
rect 111 95 115 99
rect 775 95 779 99
rect 147 87 151 91
rect 203 87 207 91
rect 259 87 263 91
rect 315 87 319 91
rect 371 87 375 91
rect 427 87 431 91
rect 483 87 487 91
rect 539 87 543 91
<< m3 >>
rect 111 818 115 819
rect 195 818 199 819
rect 251 818 255 819
rect 307 818 311 819
rect 363 818 367 819
rect 419 818 423 819
rect 475 818 479 819
rect 539 818 543 819
rect 603 818 607 819
rect 667 818 671 819
rect 723 818 727 819
rect 775 818 779 819
rect 111 813 115 814
rect 194 813 200 814
rect 112 806 114 813
rect 194 809 195 813
rect 199 809 200 813
rect 194 808 200 809
rect 250 813 256 814
rect 250 809 251 813
rect 255 809 256 813
rect 250 808 256 809
rect 306 813 312 814
rect 306 809 307 813
rect 311 809 312 813
rect 306 808 312 809
rect 362 813 368 814
rect 362 809 363 813
rect 367 809 368 813
rect 362 808 368 809
rect 418 813 424 814
rect 418 809 419 813
rect 423 809 424 813
rect 418 808 424 809
rect 474 813 480 814
rect 474 809 475 813
rect 479 809 480 813
rect 474 808 480 809
rect 538 813 544 814
rect 538 809 539 813
rect 543 809 544 813
rect 538 808 544 809
rect 602 813 608 814
rect 602 809 603 813
rect 607 809 608 813
rect 602 808 608 809
rect 666 813 672 814
rect 666 809 667 813
rect 671 809 672 813
rect 666 808 672 809
rect 722 813 728 814
rect 775 813 779 814
rect 722 809 723 813
rect 727 809 728 813
rect 722 808 728 809
rect 776 806 778 813
rect 110 805 116 806
rect 110 801 111 805
rect 115 801 116 805
rect 110 800 116 801
rect 774 805 780 806
rect 774 801 775 805
rect 779 801 780 805
rect 774 800 780 801
rect 110 787 116 788
rect 110 783 111 787
rect 115 783 116 787
rect 110 782 116 783
rect 194 787 200 788
rect 194 783 195 787
rect 199 783 200 787
rect 194 782 200 783
rect 734 787 740 788
rect 734 783 735 787
rect 739 783 740 787
rect 734 782 740 783
rect 774 787 780 788
rect 774 783 775 787
rect 779 783 780 787
rect 774 782 780 783
rect 112 763 114 782
rect 196 764 198 782
rect 218 775 224 776
rect 218 771 219 775
rect 223 771 224 775
rect 218 770 224 771
rect 274 775 280 776
rect 274 771 275 775
rect 279 771 280 775
rect 274 770 280 771
rect 330 775 336 776
rect 330 771 331 775
rect 335 771 336 775
rect 330 770 336 771
rect 386 775 392 776
rect 386 771 387 775
rect 391 771 392 775
rect 386 770 392 771
rect 442 775 448 776
rect 442 771 443 775
rect 447 771 448 775
rect 442 770 448 771
rect 498 775 504 776
rect 498 771 499 775
rect 503 771 504 775
rect 498 770 504 771
rect 562 775 568 776
rect 562 771 563 775
rect 567 771 568 775
rect 562 770 568 771
rect 574 775 580 776
rect 574 771 575 775
rect 579 771 580 775
rect 574 770 580 771
rect 626 775 632 776
rect 626 771 627 775
rect 631 771 632 775
rect 626 770 632 771
rect 690 775 696 776
rect 690 771 691 775
rect 695 771 696 775
rect 690 770 696 771
rect 194 763 200 764
rect 220 763 222 770
rect 276 763 278 770
rect 332 763 334 770
rect 388 763 390 770
rect 444 763 446 770
rect 500 763 502 770
rect 564 763 566 770
rect 111 762 115 763
rect 194 759 195 763
rect 199 759 200 763
rect 194 758 200 759
rect 203 762 207 763
rect 219 762 223 763
rect 267 762 271 763
rect 275 762 279 763
rect 111 757 115 758
rect 202 757 208 758
rect 219 757 223 758
rect 266 757 272 758
rect 275 757 279 758
rect 331 762 335 763
rect 339 762 343 763
rect 387 762 391 763
rect 419 762 423 763
rect 443 762 447 763
rect 331 757 335 758
rect 338 757 344 758
rect 387 757 391 758
rect 418 757 424 758
rect 443 757 447 758
rect 499 762 503 763
rect 507 762 511 763
rect 563 762 567 763
rect 499 757 503 758
rect 506 757 512 758
rect 563 757 567 758
rect 112 746 114 757
rect 202 753 203 757
rect 207 753 208 757
rect 202 752 208 753
rect 266 753 267 757
rect 271 753 272 757
rect 266 752 272 753
rect 338 753 339 757
rect 343 753 344 757
rect 338 752 344 753
rect 418 753 419 757
rect 423 753 424 757
rect 418 752 424 753
rect 490 755 496 756
rect 490 751 491 755
rect 495 751 496 755
rect 506 753 507 757
rect 511 753 512 757
rect 506 752 512 753
rect 490 750 496 751
rect 110 745 116 746
rect 110 741 111 745
rect 115 741 116 745
rect 110 740 116 741
rect 198 743 204 744
rect 198 739 199 743
rect 203 739 204 743
rect 198 738 204 739
rect 110 727 116 728
rect 110 723 111 727
rect 115 723 116 727
rect 110 722 116 723
rect 112 707 114 722
rect 178 719 184 720
rect 178 715 179 719
rect 183 715 184 719
rect 178 714 184 715
rect 180 707 182 714
rect 111 706 115 707
rect 111 701 115 702
rect 179 706 183 707
rect 179 701 183 702
rect 112 694 114 701
rect 110 693 116 694
rect 110 689 111 693
rect 115 689 116 693
rect 110 688 116 689
rect 110 675 116 676
rect 110 671 111 675
rect 115 671 116 675
rect 110 670 116 671
rect 112 655 114 670
rect 200 664 202 738
rect 242 719 248 720
rect 242 715 243 719
rect 247 715 248 719
rect 242 714 248 715
rect 314 719 320 720
rect 314 715 315 719
rect 319 715 320 719
rect 314 714 320 715
rect 394 719 400 720
rect 394 715 395 719
rect 399 715 400 719
rect 394 714 400 715
rect 482 719 488 720
rect 482 715 483 719
rect 487 715 488 719
rect 482 714 488 715
rect 244 707 246 714
rect 316 707 318 714
rect 396 707 398 714
rect 484 707 486 714
rect 227 706 231 707
rect 243 706 247 707
rect 226 701 232 702
rect 243 701 247 702
rect 315 706 319 707
rect 331 706 335 707
rect 395 706 399 707
rect 435 706 439 707
rect 483 706 487 707
rect 492 704 494 750
rect 576 748 578 770
rect 628 763 630 770
rect 692 763 694 770
rect 595 762 599 763
rect 627 762 631 763
rect 683 762 687 763
rect 691 762 695 763
rect 736 760 738 782
rect 746 775 752 776
rect 746 771 747 775
rect 751 771 752 775
rect 746 770 752 771
rect 748 763 750 770
rect 776 763 778 782
rect 747 762 751 763
rect 594 757 600 758
rect 627 757 631 758
rect 682 757 688 758
rect 691 757 695 758
rect 734 759 740 760
rect 594 753 595 757
rect 599 753 600 757
rect 594 752 600 753
rect 682 753 683 757
rect 687 753 688 757
rect 734 755 735 759
rect 739 755 740 759
rect 775 762 779 763
rect 734 754 740 755
rect 746 757 752 758
rect 775 757 779 758
rect 682 752 688 753
rect 746 753 747 757
rect 751 753 752 757
rect 746 752 752 753
rect 574 747 580 748
rect 574 743 575 747
rect 579 743 580 747
rect 776 746 778 757
rect 574 742 580 743
rect 774 745 780 746
rect 774 741 775 745
rect 779 741 780 745
rect 774 740 780 741
rect 774 727 780 728
rect 774 723 775 727
rect 779 723 780 727
rect 774 722 780 723
rect 570 719 576 720
rect 570 715 571 719
rect 575 715 576 719
rect 570 714 576 715
rect 658 719 664 720
rect 658 715 659 719
rect 663 715 664 719
rect 658 714 664 715
rect 722 719 728 720
rect 722 715 723 719
rect 727 715 728 719
rect 722 714 728 715
rect 572 707 574 714
rect 650 711 656 712
rect 650 707 651 711
rect 655 707 656 711
rect 660 707 662 714
rect 724 707 726 714
rect 776 707 778 722
rect 539 706 543 707
rect 315 701 319 702
rect 330 701 336 702
rect 395 701 399 702
rect 434 701 440 702
rect 483 701 487 702
rect 490 703 496 704
rect 226 697 227 701
rect 231 697 232 701
rect 226 696 232 697
rect 330 697 331 701
rect 335 697 336 701
rect 330 696 336 697
rect 434 697 435 701
rect 439 697 440 701
rect 490 699 491 703
rect 495 699 496 703
rect 571 706 575 707
rect 643 706 647 707
rect 650 706 656 707
rect 659 706 663 707
rect 490 698 496 699
rect 538 701 544 702
rect 571 701 575 702
rect 642 701 648 702
rect 434 696 440 697
rect 538 697 539 701
rect 543 697 544 701
rect 538 696 544 697
rect 642 697 643 701
rect 647 697 648 701
rect 642 696 648 697
rect 478 675 484 676
rect 478 671 479 675
rect 483 671 484 675
rect 478 670 484 671
rect 198 663 204 664
rect 198 659 199 663
rect 203 659 204 663
rect 198 658 204 659
rect 250 663 256 664
rect 250 659 251 663
rect 255 659 256 663
rect 250 658 256 659
rect 354 663 360 664
rect 354 659 355 663
rect 359 659 360 663
rect 354 658 360 659
rect 458 663 464 664
rect 458 659 459 663
rect 463 659 464 663
rect 458 658 464 659
rect 252 655 254 658
rect 356 655 358 658
rect 460 655 462 658
rect 111 654 115 655
rect 111 649 115 650
rect 251 654 255 655
rect 307 654 311 655
rect 355 654 359 655
rect 363 654 367 655
rect 427 654 431 655
rect 459 654 463 655
rect 480 652 482 670
rect 652 664 654 706
rect 723 706 727 707
rect 775 706 779 707
rect 659 701 663 702
rect 722 701 728 702
rect 775 701 779 702
rect 722 697 723 701
rect 727 697 728 701
rect 722 696 728 697
rect 776 694 778 701
rect 774 693 780 694
rect 774 689 775 693
rect 779 689 780 693
rect 774 688 780 689
rect 734 675 740 676
rect 734 671 735 675
rect 739 671 740 675
rect 734 670 740 671
rect 774 675 780 676
rect 774 671 775 675
rect 779 671 780 675
rect 774 670 780 671
rect 550 663 556 664
rect 550 659 551 663
rect 555 659 556 663
rect 550 658 556 659
rect 562 663 568 664
rect 562 659 563 663
rect 567 659 568 663
rect 562 658 568 659
rect 650 663 656 664
rect 650 659 651 663
rect 655 659 656 663
rect 650 658 656 659
rect 666 663 672 664
rect 666 659 667 663
rect 671 659 672 663
rect 666 658 672 659
rect 499 654 503 655
rect 251 649 255 650
rect 306 649 312 650
rect 355 649 359 650
rect 362 649 368 650
rect 112 638 114 649
rect 306 645 307 649
rect 311 645 312 649
rect 306 644 312 645
rect 362 645 363 649
rect 367 645 368 649
rect 362 644 368 645
rect 426 649 432 650
rect 459 649 463 650
rect 478 651 484 652
rect 426 645 427 649
rect 431 645 432 649
rect 478 647 479 651
rect 483 647 484 651
rect 478 646 484 647
rect 498 649 504 650
rect 426 644 432 645
rect 498 645 499 649
rect 503 645 504 649
rect 498 644 504 645
rect 552 640 554 658
rect 564 655 566 658
rect 668 655 670 658
rect 563 654 567 655
rect 579 654 583 655
rect 667 654 671 655
rect 736 652 738 670
rect 746 663 752 664
rect 746 659 747 663
rect 751 659 752 663
rect 746 658 752 659
rect 748 655 750 658
rect 776 655 778 670
rect 747 654 751 655
rect 734 651 740 652
rect 563 649 567 650
rect 578 649 584 650
rect 578 645 579 649
rect 583 645 584 649
rect 666 649 672 650
rect 578 644 584 645
rect 630 647 636 648
rect 630 643 631 647
rect 635 643 636 647
rect 666 645 667 649
rect 671 645 672 649
rect 734 647 735 651
rect 739 647 740 651
rect 775 654 779 655
rect 734 646 740 647
rect 746 649 752 650
rect 775 649 779 650
rect 666 644 672 645
rect 746 645 747 649
rect 751 645 752 649
rect 746 644 752 645
rect 630 642 636 643
rect 550 639 556 640
rect 110 637 116 638
rect 110 633 111 637
rect 115 633 116 637
rect 110 632 116 633
rect 294 635 300 636
rect 294 631 295 635
rect 299 631 300 635
rect 550 635 551 639
rect 555 635 556 639
rect 550 634 556 635
rect 294 630 300 631
rect 110 619 116 620
rect 110 615 111 619
rect 115 615 116 619
rect 110 614 116 615
rect 112 607 114 614
rect 282 611 288 612
rect 282 607 283 611
rect 287 607 288 611
rect 111 606 115 607
rect 282 606 288 607
rect 111 601 115 602
rect 283 601 287 602
rect 112 594 114 601
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 110 588 116 589
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 110 570 116 571
rect 112 559 114 570
rect 296 564 298 630
rect 338 611 344 612
rect 338 607 339 611
rect 343 607 344 611
rect 402 611 408 612
rect 402 607 403 611
rect 407 607 408 611
rect 474 611 480 612
rect 474 607 475 611
rect 479 607 480 611
rect 554 611 560 612
rect 554 607 555 611
rect 559 607 560 611
rect 338 606 344 607
rect 347 606 351 607
rect 402 606 408 607
rect 411 606 415 607
rect 474 606 480 607
rect 483 606 487 607
rect 554 606 560 607
rect 563 606 567 607
rect 632 604 634 642
rect 776 638 778 649
rect 774 637 780 638
rect 774 633 775 637
rect 779 633 780 637
rect 774 632 780 633
rect 774 619 780 620
rect 774 615 775 619
rect 779 615 780 619
rect 774 614 780 615
rect 642 611 648 612
rect 642 607 643 611
rect 647 607 648 611
rect 722 611 728 612
rect 722 607 723 611
rect 727 607 728 611
rect 776 607 778 614
rect 642 606 648 607
rect 651 606 655 607
rect 722 606 728 607
rect 775 606 779 607
rect 630 603 636 604
rect 339 601 343 602
rect 346 601 352 602
rect 403 601 407 602
rect 410 601 416 602
rect 475 601 479 602
rect 482 601 488 602
rect 555 601 559 602
rect 562 601 568 602
rect 346 597 347 601
rect 351 597 352 601
rect 346 596 352 597
rect 410 597 411 601
rect 415 597 416 601
rect 410 596 416 597
rect 482 597 483 601
rect 487 597 488 601
rect 482 596 488 597
rect 562 597 563 601
rect 567 597 568 601
rect 630 599 631 603
rect 635 599 636 603
rect 643 601 647 602
rect 650 601 656 602
rect 630 598 636 599
rect 562 596 568 597
rect 650 597 651 601
rect 655 597 656 601
rect 650 596 656 597
rect 722 601 728 602
rect 775 601 779 602
rect 722 597 723 601
rect 727 597 728 601
rect 722 596 728 597
rect 776 594 778 601
rect 774 593 780 594
rect 774 589 775 593
rect 779 589 780 593
rect 774 588 780 589
rect 562 575 568 576
rect 562 571 563 575
rect 567 571 568 575
rect 562 570 568 571
rect 734 575 740 576
rect 734 571 735 575
rect 739 571 740 575
rect 734 570 740 571
rect 774 575 780 576
rect 774 571 775 575
rect 779 571 780 575
rect 774 570 780 571
rect 294 563 300 564
rect 294 559 295 563
rect 299 559 300 563
rect 370 563 376 564
rect 370 559 371 563
rect 375 559 376 563
rect 434 563 440 564
rect 434 559 435 563
rect 439 559 440 563
rect 506 563 512 564
rect 506 559 507 563
rect 511 559 512 563
rect 111 558 115 559
rect 294 558 300 559
rect 347 558 351 559
rect 370 558 376 559
rect 419 558 423 559
rect 434 558 440 559
rect 499 558 503 559
rect 506 558 512 559
rect 564 556 566 570
rect 586 563 592 564
rect 586 559 587 563
rect 591 559 592 563
rect 579 558 583 559
rect 586 558 592 559
rect 646 563 652 564
rect 646 559 647 563
rect 651 559 652 563
rect 674 563 680 564
rect 674 559 675 563
rect 679 559 680 563
rect 646 558 652 559
rect 667 558 671 559
rect 674 558 680 559
rect 111 553 115 554
rect 346 553 352 554
rect 371 553 375 554
rect 418 553 424 554
rect 435 553 439 554
rect 498 553 504 554
rect 507 553 511 554
rect 562 555 568 556
rect 112 542 114 553
rect 346 549 347 553
rect 351 549 352 553
rect 346 548 352 549
rect 418 549 419 553
rect 423 549 424 553
rect 418 548 424 549
rect 498 549 499 553
rect 503 549 504 553
rect 562 551 563 555
rect 567 551 568 555
rect 562 550 568 551
rect 578 553 584 554
rect 587 553 591 554
rect 498 548 504 549
rect 578 549 579 553
rect 583 549 584 553
rect 578 548 584 549
rect 648 544 650 558
rect 736 556 738 570
rect 746 563 752 564
rect 746 559 747 563
rect 751 559 752 563
rect 776 559 778 570
rect 746 558 752 559
rect 775 558 779 559
rect 666 553 672 554
rect 675 553 679 554
rect 734 555 740 556
rect 666 549 667 553
rect 671 549 672 553
rect 734 551 735 555
rect 739 551 740 555
rect 734 550 740 551
rect 746 553 752 554
rect 775 553 779 554
rect 666 548 672 549
rect 746 549 747 553
rect 751 549 752 553
rect 746 548 752 549
rect 646 543 652 544
rect 110 541 116 542
rect 110 537 111 541
rect 115 537 116 541
rect 646 539 647 543
rect 651 539 652 543
rect 776 542 778 553
rect 646 538 652 539
rect 774 541 780 542
rect 110 536 116 537
rect 774 537 775 541
rect 779 537 780 541
rect 774 536 780 537
rect 110 523 116 524
rect 110 519 111 523
rect 115 519 116 523
rect 110 518 116 519
rect 774 523 780 524
rect 774 519 775 523
rect 779 519 780 523
rect 774 518 780 519
rect 112 511 114 518
rect 322 515 328 516
rect 322 511 323 515
rect 327 511 328 515
rect 394 515 400 516
rect 394 511 395 515
rect 399 511 400 515
rect 111 510 115 511
rect 195 510 199 511
rect 283 510 287 511
rect 322 510 328 511
rect 379 510 383 511
rect 394 510 400 511
rect 474 515 480 516
rect 474 511 475 515
rect 479 511 480 515
rect 554 515 560 516
rect 554 511 555 515
rect 559 511 560 515
rect 642 515 648 516
rect 642 511 643 515
rect 647 511 648 515
rect 474 510 480 511
rect 491 510 495 511
rect 554 510 560 511
rect 611 510 615 511
rect 642 510 648 511
rect 722 515 728 516
rect 722 511 723 515
rect 727 511 728 515
rect 776 511 778 518
rect 722 510 728 511
rect 775 510 779 511
rect 111 505 115 506
rect 194 505 200 506
rect 112 498 114 505
rect 194 501 195 505
rect 199 501 200 505
rect 194 500 200 501
rect 282 505 288 506
rect 323 505 327 506
rect 378 505 384 506
rect 395 505 399 506
rect 475 505 479 506
rect 490 505 496 506
rect 555 505 559 506
rect 610 505 616 506
rect 643 505 647 506
rect 722 505 728 506
rect 775 505 779 506
rect 282 501 283 505
rect 287 501 288 505
rect 282 500 288 501
rect 378 501 379 505
rect 383 501 384 505
rect 378 500 384 501
rect 490 501 491 505
rect 495 501 496 505
rect 490 500 496 501
rect 610 501 611 505
rect 615 501 616 505
rect 610 500 616 501
rect 722 501 723 505
rect 727 501 728 505
rect 722 500 728 501
rect 776 498 778 505
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 110 492 116 493
rect 774 497 780 498
rect 774 493 775 497
rect 779 493 780 497
rect 774 492 780 493
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 194 479 200 480
rect 194 475 195 479
rect 199 475 200 479
rect 194 474 200 475
rect 650 479 656 480
rect 650 475 651 479
rect 655 475 656 479
rect 650 474 656 475
rect 774 479 780 480
rect 774 475 775 479
rect 779 475 780 479
rect 774 474 780 475
rect 112 459 114 474
rect 196 460 198 474
rect 218 467 224 468
rect 218 463 219 467
rect 223 463 224 467
rect 218 462 224 463
rect 306 467 312 468
rect 306 463 307 467
rect 311 463 312 467
rect 306 462 312 463
rect 402 467 408 468
rect 402 463 403 467
rect 407 463 408 467
rect 402 462 408 463
rect 514 467 520 468
rect 514 463 515 467
rect 519 463 520 467
rect 514 462 520 463
rect 634 467 640 468
rect 634 463 635 467
rect 639 463 640 467
rect 634 462 640 463
rect 194 459 200 460
rect 220 459 222 462
rect 308 459 310 462
rect 404 459 406 462
rect 516 459 518 462
rect 636 459 638 462
rect 111 458 115 459
rect 171 458 175 459
rect 194 455 195 459
rect 199 455 200 459
rect 194 454 200 455
rect 219 458 223 459
rect 227 458 231 459
rect 299 458 303 459
rect 307 458 311 459
rect 387 458 391 459
rect 403 458 407 459
rect 475 458 479 459
rect 515 458 519 459
rect 571 458 575 459
rect 635 458 639 459
rect 652 456 654 474
rect 746 467 752 468
rect 746 463 747 467
rect 751 463 752 467
rect 746 462 752 463
rect 748 459 750 462
rect 776 459 778 474
rect 667 458 671 459
rect 111 453 115 454
rect 170 453 176 454
rect 219 453 223 454
rect 226 453 232 454
rect 112 442 114 453
rect 170 449 171 453
rect 175 449 176 453
rect 170 448 176 449
rect 226 449 227 453
rect 231 449 232 453
rect 226 448 232 449
rect 298 453 304 454
rect 307 453 311 454
rect 386 453 392 454
rect 403 453 407 454
rect 474 453 480 454
rect 515 453 519 454
rect 570 453 576 454
rect 635 453 639 454
rect 650 455 656 456
rect 298 449 299 453
rect 303 449 304 453
rect 298 448 304 449
rect 386 449 387 453
rect 391 449 392 453
rect 386 448 392 449
rect 474 449 475 453
rect 479 449 480 453
rect 474 448 480 449
rect 562 451 568 452
rect 562 447 563 451
rect 567 447 568 451
rect 570 449 571 453
rect 575 449 576 453
rect 650 451 651 455
rect 655 451 656 455
rect 747 458 751 459
rect 775 458 779 459
rect 650 450 656 451
rect 666 453 672 454
rect 570 448 576 449
rect 666 449 667 453
rect 671 449 672 453
rect 666 448 672 449
rect 746 453 752 454
rect 775 453 779 454
rect 746 449 747 453
rect 751 449 752 453
rect 746 448 752 449
rect 562 446 568 447
rect 110 441 116 442
rect 110 437 111 441
rect 115 437 116 441
rect 110 436 116 437
rect 110 423 116 424
rect 110 419 111 423
rect 115 419 116 423
rect 110 418 116 419
rect 112 403 114 418
rect 146 415 152 416
rect 146 411 147 415
rect 151 411 152 415
rect 146 410 152 411
rect 202 415 208 416
rect 202 411 203 415
rect 207 411 208 415
rect 202 410 208 411
rect 274 415 280 416
rect 274 411 275 415
rect 279 411 280 415
rect 274 410 280 411
rect 362 415 368 416
rect 362 411 363 415
rect 367 411 368 415
rect 362 410 368 411
rect 450 415 456 416
rect 450 411 451 415
rect 455 411 456 415
rect 450 410 456 411
rect 546 415 552 416
rect 546 411 547 415
rect 551 411 552 415
rect 546 410 552 411
rect 148 403 150 410
rect 204 403 206 410
rect 276 403 278 410
rect 364 403 366 410
rect 452 403 454 410
rect 548 403 550 410
rect 111 402 115 403
rect 147 402 151 403
rect 203 402 207 403
rect 227 402 231 403
rect 275 402 279 403
rect 315 402 319 403
rect 363 402 367 403
rect 411 402 415 403
rect 451 402 455 403
rect 515 402 519 403
rect 547 402 551 403
rect 564 400 566 446
rect 776 442 778 453
rect 774 441 780 442
rect 774 437 775 441
rect 779 437 780 441
rect 774 436 780 437
rect 774 423 780 424
rect 774 419 775 423
rect 779 419 780 423
rect 774 418 780 419
rect 642 415 648 416
rect 642 411 643 415
rect 647 411 648 415
rect 642 410 648 411
rect 722 415 728 416
rect 722 411 723 415
rect 727 411 728 415
rect 722 410 728 411
rect 644 403 646 410
rect 724 403 726 410
rect 776 403 778 418
rect 627 402 631 403
rect 111 397 115 398
rect 146 397 152 398
rect 203 397 207 398
rect 226 397 232 398
rect 275 397 279 398
rect 314 397 320 398
rect 363 397 367 398
rect 410 397 416 398
rect 451 397 455 398
rect 514 397 520 398
rect 547 397 551 398
rect 562 399 568 400
rect 112 390 114 397
rect 146 393 147 397
rect 151 393 152 397
rect 146 392 152 393
rect 226 393 227 397
rect 231 393 232 397
rect 226 392 232 393
rect 314 393 315 397
rect 319 393 320 397
rect 314 392 320 393
rect 410 393 411 397
rect 415 393 416 397
rect 410 392 416 393
rect 514 393 515 397
rect 519 393 520 397
rect 562 395 563 399
rect 567 395 568 399
rect 643 402 647 403
rect 723 402 727 403
rect 775 402 779 403
rect 562 394 568 395
rect 626 397 632 398
rect 643 397 647 398
rect 722 397 728 398
rect 775 397 779 398
rect 514 392 520 393
rect 626 393 627 397
rect 631 393 632 397
rect 626 392 632 393
rect 722 393 723 397
rect 727 393 728 397
rect 722 392 728 393
rect 776 390 778 397
rect 110 389 116 390
rect 110 385 111 389
rect 115 385 116 389
rect 110 384 116 385
rect 774 389 780 390
rect 774 385 775 389
rect 779 385 780 389
rect 774 384 780 385
rect 110 371 116 372
rect 110 367 111 371
rect 115 367 116 371
rect 110 366 116 367
rect 530 371 536 372
rect 530 367 531 371
rect 535 367 536 371
rect 530 366 536 367
rect 674 371 680 372
rect 674 367 675 371
rect 679 367 680 371
rect 674 366 680 367
rect 774 371 780 372
rect 774 367 775 371
rect 779 367 780 371
rect 774 366 780 367
rect 112 355 114 366
rect 170 359 176 360
rect 170 355 171 359
rect 175 355 176 359
rect 111 354 115 355
rect 170 354 176 355
rect 250 359 256 360
rect 250 355 251 359
rect 255 355 256 359
rect 338 359 344 360
rect 338 355 339 359
rect 343 355 344 359
rect 434 359 440 360
rect 434 355 435 359
rect 439 355 440 359
rect 250 354 256 355
rect 315 354 319 355
rect 338 354 344 355
rect 371 354 375 355
rect 434 354 440 355
rect 499 354 503 355
rect 111 349 115 350
rect 171 349 175 350
rect 532 352 534 366
rect 538 359 544 360
rect 538 355 539 359
rect 543 355 544 359
rect 606 359 612 360
rect 606 355 607 359
rect 611 355 612 359
rect 650 359 656 360
rect 650 355 651 359
rect 655 355 656 359
rect 538 354 544 355
rect 563 354 567 355
rect 606 354 612 355
rect 627 354 631 355
rect 650 354 656 355
rect 530 351 536 352
rect 251 349 255 350
rect 314 349 320 350
rect 339 349 343 350
rect 370 349 376 350
rect 112 338 114 349
rect 314 345 315 349
rect 319 345 320 349
rect 314 344 320 345
rect 370 345 371 349
rect 375 345 376 349
rect 370 344 376 345
rect 434 349 440 350
rect 434 345 435 349
rect 439 345 440 349
rect 434 344 440 345
rect 498 349 504 350
rect 498 345 499 349
rect 503 345 504 349
rect 530 347 531 351
rect 535 347 536 351
rect 539 349 543 350
rect 562 349 568 350
rect 530 346 536 347
rect 498 344 504 345
rect 562 345 563 349
rect 567 345 568 349
rect 562 344 568 345
rect 570 347 576 348
rect 570 343 571 347
rect 575 343 576 347
rect 570 342 576 343
rect 110 337 116 338
rect 110 333 111 337
rect 115 333 116 337
rect 110 332 116 333
rect 434 331 440 332
rect 434 327 435 331
rect 439 327 440 331
rect 434 326 440 327
rect 110 319 116 320
rect 110 315 111 319
rect 115 315 116 319
rect 110 314 116 315
rect 112 307 114 314
rect 290 311 296 312
rect 290 307 291 311
rect 295 307 296 311
rect 346 311 352 312
rect 346 307 347 311
rect 351 307 352 311
rect 410 311 416 312
rect 410 307 411 311
rect 415 307 416 311
rect 111 306 115 307
rect 219 306 223 307
rect 275 306 279 307
rect 290 306 296 307
rect 331 306 335 307
rect 346 306 352 307
rect 387 306 391 307
rect 410 306 416 307
rect 111 301 115 302
rect 218 301 224 302
rect 112 294 114 301
rect 218 297 219 301
rect 223 297 224 301
rect 218 296 224 297
rect 274 301 280 302
rect 291 301 295 302
rect 330 301 336 302
rect 347 301 351 302
rect 386 301 392 302
rect 411 301 415 302
rect 274 297 275 301
rect 279 297 280 301
rect 274 296 280 297
rect 330 297 331 301
rect 335 297 336 301
rect 330 296 336 297
rect 386 297 387 301
rect 391 297 392 301
rect 386 296 392 297
rect 110 293 116 294
rect 110 289 111 293
rect 115 289 116 293
rect 110 288 116 289
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 110 270 116 271
rect 218 275 224 276
rect 218 271 219 275
rect 223 271 224 275
rect 218 270 224 271
rect 112 247 114 270
rect 220 248 222 270
rect 436 264 438 326
rect 474 311 480 312
rect 474 307 475 311
rect 479 307 480 311
rect 538 311 544 312
rect 538 307 539 311
rect 543 307 544 311
rect 443 306 447 307
rect 474 306 480 307
rect 499 306 503 307
rect 538 306 544 307
rect 555 306 559 307
rect 442 301 448 302
rect 475 301 479 302
rect 498 301 504 302
rect 539 301 543 302
rect 554 301 560 302
rect 442 297 443 301
rect 447 297 448 301
rect 442 296 448 297
rect 498 297 499 301
rect 503 297 504 301
rect 498 296 504 297
rect 554 297 555 301
rect 559 297 560 301
rect 554 296 560 297
rect 572 284 574 342
rect 608 340 610 354
rect 676 352 678 366
rect 746 359 752 360
rect 746 355 747 359
rect 751 355 752 359
rect 776 355 778 366
rect 691 354 695 355
rect 746 354 752 355
rect 775 354 779 355
rect 626 349 632 350
rect 651 349 655 350
rect 674 351 680 352
rect 626 345 627 349
rect 631 345 632 349
rect 674 347 675 351
rect 679 347 680 351
rect 674 346 680 347
rect 690 349 696 350
rect 626 344 632 345
rect 690 345 691 349
rect 695 345 696 349
rect 690 344 696 345
rect 746 349 752 350
rect 775 349 779 350
rect 746 345 747 349
rect 751 345 752 349
rect 746 344 752 345
rect 606 339 612 340
rect 606 335 607 339
rect 611 335 612 339
rect 776 338 778 349
rect 606 334 612 335
rect 774 337 780 338
rect 774 333 775 337
rect 779 333 780 337
rect 774 332 780 333
rect 774 319 780 320
rect 774 315 775 319
rect 779 315 780 319
rect 774 314 780 315
rect 602 311 608 312
rect 602 307 603 311
rect 607 307 608 311
rect 666 311 672 312
rect 666 307 667 311
rect 671 307 672 311
rect 602 306 608 307
rect 611 306 615 307
rect 666 306 672 307
rect 722 311 728 312
rect 722 307 723 311
rect 727 307 728 311
rect 776 307 778 314
rect 722 306 728 307
rect 775 306 779 307
rect 603 301 607 302
rect 610 301 616 302
rect 610 297 611 301
rect 615 297 616 301
rect 610 296 616 297
rect 666 301 672 302
rect 666 297 667 301
rect 671 297 672 301
rect 666 296 672 297
rect 722 301 728 302
rect 775 301 779 302
rect 722 297 723 301
rect 727 297 728 301
rect 722 296 728 297
rect 776 294 778 301
rect 774 293 780 294
rect 774 289 775 293
rect 779 289 780 293
rect 774 288 780 289
rect 570 283 576 284
rect 570 279 571 283
rect 575 279 576 283
rect 570 278 576 279
rect 774 275 780 276
rect 774 271 775 275
rect 779 271 780 275
rect 774 270 780 271
rect 242 263 248 264
rect 242 259 243 263
rect 247 259 248 263
rect 242 258 248 259
rect 298 263 304 264
rect 298 259 299 263
rect 303 259 304 263
rect 298 258 304 259
rect 354 263 360 264
rect 354 259 355 263
rect 359 259 360 263
rect 354 258 360 259
rect 410 263 416 264
rect 410 259 411 263
rect 415 259 416 263
rect 410 258 416 259
rect 434 263 440 264
rect 434 259 435 263
rect 439 259 440 263
rect 434 258 440 259
rect 466 263 472 264
rect 466 259 467 263
rect 471 259 472 263
rect 466 258 472 259
rect 522 263 528 264
rect 522 259 523 263
rect 527 259 528 263
rect 522 258 528 259
rect 578 263 584 264
rect 578 259 579 263
rect 583 259 584 263
rect 578 258 584 259
rect 634 263 640 264
rect 634 259 635 263
rect 639 259 640 263
rect 634 258 640 259
rect 690 263 696 264
rect 690 259 691 263
rect 695 259 696 263
rect 690 258 696 259
rect 746 263 752 264
rect 746 259 747 263
rect 751 259 752 263
rect 746 258 752 259
rect 218 247 224 248
rect 244 247 246 258
rect 300 247 302 258
rect 356 247 358 258
rect 412 247 414 258
rect 468 247 470 258
rect 524 247 526 258
rect 580 247 582 258
rect 636 247 638 258
rect 692 247 694 258
rect 748 247 750 258
rect 776 247 778 270
rect 111 246 115 247
rect 218 243 219 247
rect 223 243 224 247
rect 218 242 224 243
rect 243 246 247 247
rect 111 241 115 242
rect 243 241 247 242
rect 299 246 303 247
rect 307 246 311 247
rect 355 246 359 247
rect 363 246 367 247
rect 411 246 415 247
rect 419 246 423 247
rect 467 246 471 247
rect 475 246 479 247
rect 523 246 527 247
rect 531 246 535 247
rect 579 246 583 247
rect 299 241 303 242
rect 306 241 312 242
rect 355 241 359 242
rect 362 241 368 242
rect 411 241 415 242
rect 418 241 424 242
rect 467 241 471 242
rect 474 241 480 242
rect 523 241 527 242
rect 530 241 536 242
rect 579 241 583 242
rect 635 246 639 247
rect 635 241 639 242
rect 691 246 695 247
rect 691 241 695 242
rect 747 246 751 247
rect 747 241 751 242
rect 775 246 779 247
rect 775 241 779 242
rect 112 230 114 241
rect 306 237 307 241
rect 311 237 312 241
rect 306 236 312 237
rect 362 237 363 241
rect 367 237 368 241
rect 362 236 368 237
rect 418 237 419 241
rect 423 237 424 241
rect 418 236 424 237
rect 474 237 475 241
rect 479 237 480 241
rect 474 236 480 237
rect 530 237 531 241
rect 535 237 536 241
rect 530 236 536 237
rect 776 230 778 241
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 774 229 780 230
rect 774 225 775 229
rect 779 225 780 229
rect 774 224 780 225
rect 362 223 368 224
rect 362 219 363 223
rect 367 219 368 223
rect 362 218 368 219
rect 110 211 116 212
rect 110 207 111 211
rect 115 207 116 211
rect 110 206 116 207
rect 112 195 114 206
rect 282 203 288 204
rect 282 199 283 203
rect 287 199 288 203
rect 282 198 288 199
rect 338 203 344 204
rect 338 199 339 203
rect 343 199 344 203
rect 338 198 344 199
rect 284 195 286 198
rect 340 195 342 198
rect 111 194 115 195
rect 163 194 167 195
rect 219 194 223 195
rect 275 194 279 195
rect 283 194 287 195
rect 331 194 335 195
rect 339 194 343 195
rect 111 189 115 190
rect 162 189 168 190
rect 112 182 114 189
rect 162 185 163 189
rect 167 185 168 189
rect 162 184 168 185
rect 218 189 224 190
rect 218 185 219 189
rect 223 185 224 189
rect 218 184 224 185
rect 274 189 280 190
rect 283 189 287 190
rect 330 189 336 190
rect 339 189 343 190
rect 274 185 275 189
rect 279 185 280 189
rect 274 184 280 185
rect 330 185 331 189
rect 335 185 336 189
rect 330 184 336 185
rect 110 181 116 182
rect 110 177 111 181
rect 115 177 116 181
rect 110 176 116 177
rect 110 163 116 164
rect 110 159 111 163
rect 115 159 116 163
rect 110 158 116 159
rect 162 163 168 164
rect 162 159 163 163
rect 167 159 168 163
rect 162 158 168 159
rect 112 135 114 158
rect 164 149 166 158
rect 364 152 366 218
rect 774 211 780 212
rect 774 207 775 211
rect 779 207 780 211
rect 774 206 780 207
rect 394 203 400 204
rect 394 199 395 203
rect 399 199 400 203
rect 394 198 400 199
rect 450 203 456 204
rect 450 199 451 203
rect 455 199 456 203
rect 450 198 456 199
rect 506 203 512 204
rect 506 199 507 203
rect 511 199 512 203
rect 506 198 512 199
rect 396 195 398 198
rect 452 195 454 198
rect 508 195 510 198
rect 776 195 778 206
rect 387 194 391 195
rect 395 194 399 195
rect 386 189 392 190
rect 395 189 399 190
rect 451 194 455 195
rect 451 189 455 190
rect 507 194 511 195
rect 507 189 511 190
rect 775 194 779 195
rect 775 189 779 190
rect 386 185 387 189
rect 391 185 392 189
rect 386 184 392 185
rect 776 182 778 189
rect 774 181 780 182
rect 774 177 775 181
rect 779 177 780 181
rect 774 176 780 177
rect 774 163 780 164
rect 774 159 775 163
rect 779 159 780 163
rect 774 158 780 159
rect 186 151 192 152
rect 163 148 167 149
rect 186 147 187 151
rect 191 147 192 151
rect 186 146 192 147
rect 242 151 248 152
rect 242 147 243 151
rect 247 147 248 151
rect 242 146 248 147
rect 298 151 304 152
rect 298 147 299 151
rect 303 147 304 151
rect 298 146 304 147
rect 354 151 360 152
rect 354 147 355 151
rect 359 147 360 151
rect 354 146 360 147
rect 362 151 368 152
rect 362 147 363 151
rect 367 147 368 151
rect 362 146 368 147
rect 410 151 416 152
rect 410 147 411 151
rect 415 147 416 151
rect 410 146 416 147
rect 543 148 547 149
rect 163 143 167 144
rect 188 135 190 146
rect 244 135 246 146
rect 300 135 302 146
rect 356 135 358 146
rect 412 135 414 146
rect 543 143 547 144
rect 111 134 115 135
rect 171 134 175 135
rect 187 134 191 135
rect 227 134 231 135
rect 243 134 247 135
rect 283 134 287 135
rect 299 134 303 135
rect 339 134 343 135
rect 355 134 359 135
rect 395 134 399 135
rect 411 134 415 135
rect 451 134 455 135
rect 507 134 511 135
rect 544 132 546 143
rect 776 135 778 158
rect 563 134 567 135
rect 542 131 548 132
rect 111 129 115 130
rect 170 129 176 130
rect 187 129 191 130
rect 226 129 232 130
rect 243 129 247 130
rect 282 129 288 130
rect 299 129 303 130
rect 338 129 344 130
rect 355 129 359 130
rect 394 129 400 130
rect 411 129 415 130
rect 450 129 456 130
rect 112 118 114 129
rect 170 125 171 129
rect 175 125 176 129
rect 170 124 176 125
rect 226 125 227 129
rect 231 125 232 129
rect 226 124 232 125
rect 282 125 283 129
rect 287 125 288 129
rect 282 124 288 125
rect 338 125 339 129
rect 343 125 344 129
rect 338 124 344 125
rect 394 125 395 129
rect 399 125 400 129
rect 394 124 400 125
rect 450 125 451 129
rect 455 125 456 129
rect 450 124 456 125
rect 506 129 512 130
rect 506 125 507 129
rect 511 125 512 129
rect 542 127 543 131
rect 547 127 548 131
rect 775 134 779 135
rect 542 126 548 127
rect 562 129 568 130
rect 775 129 779 130
rect 506 124 512 125
rect 562 125 563 129
rect 567 125 568 129
rect 562 124 568 125
rect 776 118 778 129
rect 110 117 116 118
rect 110 113 111 117
rect 115 113 116 117
rect 110 112 116 113
rect 774 117 780 118
rect 774 113 775 117
rect 779 113 780 117
rect 774 112 780 113
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 774 99 780 100
rect 774 95 775 99
rect 779 95 780 99
rect 774 94 780 95
rect 112 87 114 94
rect 146 91 152 92
rect 146 87 147 91
rect 151 87 152 91
rect 111 86 115 87
rect 146 86 152 87
rect 202 91 208 92
rect 202 87 203 91
rect 207 87 208 91
rect 202 86 208 87
rect 258 91 264 92
rect 258 87 259 91
rect 263 87 264 91
rect 258 86 264 87
rect 314 91 320 92
rect 314 87 315 91
rect 319 87 320 91
rect 314 86 320 87
rect 370 91 376 92
rect 370 87 371 91
rect 375 87 376 91
rect 370 86 376 87
rect 426 91 432 92
rect 426 87 427 91
rect 431 87 432 91
rect 426 86 432 87
rect 482 91 488 92
rect 482 87 483 91
rect 487 87 488 91
rect 482 86 488 87
rect 538 91 544 92
rect 538 87 539 91
rect 543 87 544 91
rect 776 87 778 94
rect 538 86 544 87
rect 775 86 779 87
rect 111 81 115 82
rect 147 81 151 82
rect 203 81 207 82
rect 259 81 263 82
rect 315 81 319 82
rect 371 81 375 82
rect 427 81 431 82
rect 483 81 487 82
rect 539 81 543 82
rect 775 81 779 82
<< m4c >>
rect 111 814 115 818
rect 195 814 199 818
rect 251 814 255 818
rect 307 814 311 818
rect 363 814 367 818
rect 419 814 423 818
rect 475 814 479 818
rect 539 814 543 818
rect 603 814 607 818
rect 667 814 671 818
rect 723 814 727 818
rect 775 814 779 818
rect 111 758 115 762
rect 203 758 207 762
rect 219 758 223 762
rect 267 758 271 762
rect 275 758 279 762
rect 331 758 335 762
rect 339 758 343 762
rect 387 758 391 762
rect 419 758 423 762
rect 443 758 447 762
rect 499 758 503 762
rect 507 758 511 762
rect 563 758 567 762
rect 111 702 115 706
rect 179 702 183 706
rect 227 702 231 706
rect 243 702 247 706
rect 315 702 319 706
rect 331 702 335 706
rect 395 702 399 706
rect 435 702 439 706
rect 483 702 487 706
rect 595 758 599 762
rect 627 758 631 762
rect 683 758 687 762
rect 691 758 695 762
rect 747 758 751 762
rect 775 758 779 762
rect 539 702 543 706
rect 571 702 575 706
rect 643 702 647 706
rect 111 650 115 654
rect 251 650 255 654
rect 307 650 311 654
rect 355 650 359 654
rect 363 650 367 654
rect 427 650 431 654
rect 459 650 463 654
rect 659 702 663 706
rect 723 702 727 706
rect 775 702 779 706
rect 499 650 503 654
rect 563 650 567 654
rect 579 650 583 654
rect 667 650 671 654
rect 747 650 751 654
rect 775 650 779 654
rect 111 602 115 606
rect 283 602 287 606
rect 339 602 343 606
rect 347 602 351 606
rect 403 602 407 606
rect 411 602 415 606
rect 475 602 479 606
rect 483 602 487 606
rect 555 602 559 606
rect 563 602 567 606
rect 643 602 647 606
rect 651 602 655 606
rect 723 602 727 606
rect 775 602 779 606
rect 111 554 115 558
rect 347 554 351 558
rect 371 554 375 558
rect 419 554 423 558
rect 435 554 439 558
rect 499 554 503 558
rect 507 554 511 558
rect 579 554 583 558
rect 587 554 591 558
rect 667 554 671 558
rect 675 554 679 558
rect 747 554 751 558
rect 775 554 779 558
rect 111 506 115 510
rect 195 506 199 510
rect 283 506 287 510
rect 323 506 327 510
rect 379 506 383 510
rect 395 506 399 510
rect 475 506 479 510
rect 491 506 495 510
rect 555 506 559 510
rect 611 506 615 510
rect 643 506 647 510
rect 723 506 727 510
rect 775 506 779 510
rect 111 454 115 458
rect 171 454 175 458
rect 219 454 223 458
rect 227 454 231 458
rect 299 454 303 458
rect 307 454 311 458
rect 387 454 391 458
rect 403 454 407 458
rect 475 454 479 458
rect 515 454 519 458
rect 571 454 575 458
rect 635 454 639 458
rect 667 454 671 458
rect 747 454 751 458
rect 775 454 779 458
rect 111 398 115 402
rect 147 398 151 402
rect 203 398 207 402
rect 227 398 231 402
rect 275 398 279 402
rect 315 398 319 402
rect 363 398 367 402
rect 411 398 415 402
rect 451 398 455 402
rect 515 398 519 402
rect 547 398 551 402
rect 627 398 631 402
rect 643 398 647 402
rect 723 398 727 402
rect 775 398 779 402
rect 111 350 115 354
rect 171 350 175 354
rect 251 350 255 354
rect 315 350 319 354
rect 339 350 343 354
rect 371 350 375 354
rect 435 350 439 354
rect 499 350 503 354
rect 539 350 543 354
rect 563 350 567 354
rect 111 302 115 306
rect 219 302 223 306
rect 275 302 279 306
rect 291 302 295 306
rect 331 302 335 306
rect 347 302 351 306
rect 387 302 391 306
rect 411 302 415 306
rect 443 302 447 306
rect 475 302 479 306
rect 499 302 503 306
rect 539 302 543 306
rect 555 302 559 306
rect 627 350 631 354
rect 651 350 655 354
rect 691 350 695 354
rect 747 350 751 354
rect 775 350 779 354
rect 603 302 607 306
rect 611 302 615 306
rect 667 302 671 306
rect 723 302 727 306
rect 775 302 779 306
rect 111 242 115 246
rect 243 242 247 246
rect 299 242 303 246
rect 307 242 311 246
rect 355 242 359 246
rect 363 242 367 246
rect 411 242 415 246
rect 419 242 423 246
rect 467 242 471 246
rect 475 242 479 246
rect 523 242 527 246
rect 531 242 535 246
rect 579 242 583 246
rect 635 242 639 246
rect 691 242 695 246
rect 747 242 751 246
rect 775 242 779 246
rect 111 190 115 194
rect 163 190 167 194
rect 219 190 223 194
rect 275 190 279 194
rect 283 190 287 194
rect 331 190 335 194
rect 339 190 343 194
rect 387 190 391 194
rect 395 190 399 194
rect 451 190 455 194
rect 507 190 511 194
rect 775 190 779 194
rect 163 144 167 148
rect 543 144 547 148
rect 111 130 115 134
rect 171 130 175 134
rect 187 130 191 134
rect 227 130 231 134
rect 243 130 247 134
rect 283 130 287 134
rect 299 130 303 134
rect 339 130 343 134
rect 355 130 359 134
rect 395 130 399 134
rect 411 130 415 134
rect 451 130 455 134
rect 507 130 511 134
rect 563 130 567 134
rect 775 130 779 134
rect 111 82 115 86
rect 147 82 151 86
rect 203 82 207 86
rect 259 82 263 86
rect 315 82 319 86
rect 371 82 375 86
rect 427 82 431 86
rect 483 82 487 86
rect 539 82 543 86
rect 775 82 779 86
<< m4 >>
rect 84 813 85 819
rect 91 818 799 819
rect 91 814 111 818
rect 115 814 195 818
rect 199 814 251 818
rect 255 814 307 818
rect 311 814 363 818
rect 367 814 419 818
rect 423 814 475 818
rect 479 814 539 818
rect 543 814 603 818
rect 607 814 667 818
rect 671 814 723 818
rect 727 814 775 818
rect 779 814 799 818
rect 91 813 799 814
rect 805 813 806 819
rect 96 757 97 763
rect 103 762 811 763
rect 103 758 111 762
rect 115 758 203 762
rect 207 758 219 762
rect 223 758 267 762
rect 271 758 275 762
rect 279 758 331 762
rect 335 758 339 762
rect 343 758 387 762
rect 391 758 419 762
rect 423 758 443 762
rect 447 758 499 762
rect 503 758 507 762
rect 511 758 563 762
rect 567 758 595 762
rect 599 758 627 762
rect 631 758 683 762
rect 687 758 691 762
rect 695 758 747 762
rect 751 758 775 762
rect 779 758 811 762
rect 103 757 811 758
rect 817 757 818 763
rect 84 701 85 707
rect 91 706 799 707
rect 91 702 111 706
rect 115 702 179 706
rect 183 702 227 706
rect 231 702 243 706
rect 247 702 315 706
rect 319 702 331 706
rect 335 702 395 706
rect 399 702 435 706
rect 439 702 483 706
rect 487 702 539 706
rect 543 702 571 706
rect 575 702 643 706
rect 647 702 659 706
rect 663 702 723 706
rect 727 702 775 706
rect 779 702 799 706
rect 91 701 799 702
rect 805 701 806 707
rect 96 649 97 655
rect 103 654 811 655
rect 103 650 111 654
rect 115 650 251 654
rect 255 650 307 654
rect 311 650 355 654
rect 359 650 363 654
rect 367 650 427 654
rect 431 650 459 654
rect 463 650 499 654
rect 503 650 563 654
rect 567 650 579 654
rect 583 650 667 654
rect 671 650 747 654
rect 751 650 775 654
rect 779 650 811 654
rect 103 649 811 650
rect 817 649 818 655
rect 84 601 85 607
rect 91 606 799 607
rect 91 602 111 606
rect 115 602 283 606
rect 287 602 339 606
rect 343 602 347 606
rect 351 602 403 606
rect 407 602 411 606
rect 415 602 475 606
rect 479 602 483 606
rect 487 602 555 606
rect 559 602 563 606
rect 567 602 643 606
rect 647 602 651 606
rect 655 602 723 606
rect 727 602 775 606
rect 779 602 799 606
rect 91 601 799 602
rect 805 601 806 607
rect 96 553 97 559
rect 103 558 811 559
rect 103 554 111 558
rect 115 554 347 558
rect 351 554 371 558
rect 375 554 419 558
rect 423 554 435 558
rect 439 554 499 558
rect 503 554 507 558
rect 511 554 579 558
rect 583 554 587 558
rect 591 554 667 558
rect 671 554 675 558
rect 679 554 747 558
rect 751 554 775 558
rect 779 554 811 558
rect 103 553 811 554
rect 817 553 818 559
rect 84 505 85 511
rect 91 510 799 511
rect 91 506 111 510
rect 115 506 195 510
rect 199 506 283 510
rect 287 506 323 510
rect 327 506 379 510
rect 383 506 395 510
rect 399 506 475 510
rect 479 506 491 510
rect 495 506 555 510
rect 559 506 611 510
rect 615 506 643 510
rect 647 506 723 510
rect 727 506 775 510
rect 779 506 799 510
rect 91 505 799 506
rect 805 505 806 511
rect 96 453 97 459
rect 103 458 811 459
rect 103 454 111 458
rect 115 454 171 458
rect 175 454 219 458
rect 223 454 227 458
rect 231 454 299 458
rect 303 454 307 458
rect 311 454 387 458
rect 391 454 403 458
rect 407 454 475 458
rect 479 454 515 458
rect 519 454 571 458
rect 575 454 635 458
rect 639 454 667 458
rect 671 454 747 458
rect 751 454 775 458
rect 779 454 811 458
rect 103 453 811 454
rect 817 453 818 459
rect 84 397 85 403
rect 91 402 799 403
rect 91 398 111 402
rect 115 398 147 402
rect 151 398 203 402
rect 207 398 227 402
rect 231 398 275 402
rect 279 398 315 402
rect 319 398 363 402
rect 367 398 411 402
rect 415 398 451 402
rect 455 398 515 402
rect 519 398 547 402
rect 551 398 627 402
rect 631 398 643 402
rect 647 398 723 402
rect 727 398 775 402
rect 779 398 799 402
rect 91 397 799 398
rect 805 397 806 403
rect 96 349 97 355
rect 103 354 811 355
rect 103 350 111 354
rect 115 350 171 354
rect 175 350 251 354
rect 255 350 315 354
rect 319 350 339 354
rect 343 350 371 354
rect 375 350 435 354
rect 439 350 499 354
rect 503 350 539 354
rect 543 350 563 354
rect 567 350 627 354
rect 631 350 651 354
rect 655 350 691 354
rect 695 350 747 354
rect 751 350 775 354
rect 779 350 811 354
rect 103 349 811 350
rect 817 349 818 355
rect 84 301 85 307
rect 91 306 799 307
rect 91 302 111 306
rect 115 302 219 306
rect 223 302 275 306
rect 279 302 291 306
rect 295 302 331 306
rect 335 302 347 306
rect 351 302 387 306
rect 391 302 411 306
rect 415 302 443 306
rect 447 302 475 306
rect 479 302 499 306
rect 503 302 539 306
rect 543 302 555 306
rect 559 302 603 306
rect 607 302 611 306
rect 615 302 667 306
rect 671 302 723 306
rect 727 302 775 306
rect 779 302 799 306
rect 91 301 799 302
rect 805 301 806 307
rect 96 241 97 247
rect 103 246 811 247
rect 103 242 111 246
rect 115 242 243 246
rect 247 242 299 246
rect 303 242 307 246
rect 311 242 355 246
rect 359 242 363 246
rect 367 242 411 246
rect 415 242 419 246
rect 423 242 467 246
rect 471 242 475 246
rect 479 242 523 246
rect 527 242 531 246
rect 535 242 579 246
rect 583 242 635 246
rect 639 242 691 246
rect 695 242 747 246
rect 751 242 775 246
rect 779 242 811 246
rect 103 241 811 242
rect 817 241 818 247
rect 84 189 85 195
rect 91 194 799 195
rect 91 190 111 194
rect 115 190 163 194
rect 167 190 219 194
rect 223 190 275 194
rect 279 190 283 194
rect 287 190 331 194
rect 335 190 339 194
rect 343 190 387 194
rect 391 190 395 194
rect 399 190 451 194
rect 455 190 507 194
rect 511 190 775 194
rect 779 190 799 194
rect 91 189 799 190
rect 805 189 806 195
rect 162 148 168 149
rect 542 148 548 149
rect 162 144 163 148
rect 167 144 543 148
rect 547 144 548 148
rect 162 143 168 144
rect 542 143 548 144
rect 96 129 97 135
rect 103 134 811 135
rect 103 130 111 134
rect 115 130 171 134
rect 175 130 187 134
rect 191 130 227 134
rect 231 130 243 134
rect 247 130 283 134
rect 287 130 299 134
rect 303 130 339 134
rect 343 130 355 134
rect 359 130 395 134
rect 399 130 411 134
rect 415 130 451 134
rect 455 130 507 134
rect 511 130 563 134
rect 567 130 775 134
rect 779 130 811 134
rect 103 129 811 130
rect 817 129 818 135
rect 84 81 85 87
rect 91 86 799 87
rect 91 82 111 86
rect 115 82 147 86
rect 151 82 203 86
rect 207 82 259 86
rect 263 82 315 86
rect 319 82 371 86
rect 375 82 427 86
rect 431 82 483 86
rect 487 82 539 86
rect 543 82 775 86
rect 779 82 799 86
rect 91 81 799 82
rect 805 81 806 87
<< m5c >>
rect 85 813 91 819
rect 799 813 805 819
rect 97 757 103 763
rect 811 757 817 763
rect 85 701 91 707
rect 799 701 805 707
rect 97 649 103 655
rect 811 649 817 655
rect 85 601 91 607
rect 799 601 805 607
rect 97 553 103 559
rect 811 553 817 559
rect 85 505 91 511
rect 799 505 805 511
rect 97 453 103 459
rect 811 453 817 459
rect 85 397 91 403
rect 799 397 805 403
rect 97 349 103 355
rect 811 349 817 355
rect 85 301 91 307
rect 799 301 805 307
rect 97 241 103 247
rect 811 241 817 247
rect 85 189 91 195
rect 799 189 805 195
rect 97 129 103 135
rect 811 129 817 135
rect 85 81 91 87
rect 799 81 805 87
<< m5 >>
rect 84 819 92 864
rect 84 813 85 819
rect 91 813 92 819
rect 84 707 92 813
rect 84 701 85 707
rect 91 701 92 707
rect 84 607 92 701
rect 84 601 85 607
rect 91 601 92 607
rect 84 511 92 601
rect 84 505 85 511
rect 91 505 92 511
rect 84 403 92 505
rect 84 397 85 403
rect 91 397 92 403
rect 84 307 92 397
rect 84 301 85 307
rect 91 301 92 307
rect 84 195 92 301
rect 84 189 85 195
rect 91 189 92 195
rect 84 87 92 189
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 763 104 864
rect 96 757 97 763
rect 103 757 104 763
rect 96 655 104 757
rect 96 649 97 655
rect 103 649 104 655
rect 96 559 104 649
rect 96 553 97 559
rect 103 553 104 559
rect 96 459 104 553
rect 96 453 97 459
rect 103 453 104 459
rect 96 355 104 453
rect 96 349 97 355
rect 103 349 104 355
rect 96 247 104 349
rect 96 241 97 247
rect 103 241 104 247
rect 96 135 104 241
rect 96 129 97 135
rect 103 129 104 135
rect 96 72 104 129
rect 798 819 806 864
rect 798 813 799 819
rect 805 813 806 819
rect 798 707 806 813
rect 798 701 799 707
rect 805 701 806 707
rect 798 607 806 701
rect 798 601 799 607
rect 805 601 806 607
rect 798 511 806 601
rect 798 505 799 511
rect 805 505 806 511
rect 798 403 806 505
rect 798 397 799 403
rect 805 397 806 403
rect 798 307 806 397
rect 798 301 799 307
rect 805 301 806 307
rect 798 195 806 301
rect 798 189 799 195
rect 805 189 806 195
rect 798 87 806 189
rect 798 81 799 87
rect 805 81 806 87
rect 798 72 806 81
rect 810 763 818 864
rect 810 757 811 763
rect 817 757 818 763
rect 810 655 818 757
rect 810 649 811 655
rect 817 649 818 655
rect 810 559 818 649
rect 810 553 811 559
rect 817 553 818 559
rect 810 459 818 553
rect 810 453 811 459
rect 817 453 818 459
rect 810 355 818 453
rect 810 349 811 355
rect 817 349 818 355
rect 810 247 818 349
rect 810 241 811 247
rect 817 241 818 247
rect 810 135 818 241
rect 810 129 811 135
rect 817 129 818 135
rect 810 72 818 129
use welltap_svt  __well_tap__0
timestamp 1730592110
transform 1 0 104 0 1 92
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730592110
transform 1 0 104 0 1 92
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0NOR2X1  nor_599_6
timestamp 1730592110
transform 1 0 128 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_599_6
timestamp 1730592110
transform 1 0 128 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_598_6
timestamp 1730592110
transform 1 0 184 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_598_6
timestamp 1730592110
transform 1 0 184 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_597_6
timestamp 1730592110
transform 1 0 240 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_597_6
timestamp 1730592110
transform 1 0 240 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_596_6
timestamp 1730592110
transform 1 0 296 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_596_6
timestamp 1730592110
transform 1 0 296 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_595_6
timestamp 1730592110
transform 1 0 352 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_595_6
timestamp 1730592110
transform 1 0 352 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_594_6
timestamp 1730592110
transform 1 0 408 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_594_6
timestamp 1730592110
transform 1 0 408 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_593_6
timestamp 1730592110
transform 1 0 464 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_593_6
timestamp 1730592110
transform 1 0 464 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_592_6
timestamp 1730592110
transform 1 0 520 0 1 84
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_592_6
timestamp 1730592110
transform 1 0 520 0 1 84
box 9 2 47 46
use welltap_svt  __well_tap__1
timestamp 1730592110
transform 1 0 768 0 1 92
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730592110
transform 1 0 768 0 1 92
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730592110
transform 1 0 104 0 -1 184
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730592110
transform 1 0 104 0 -1 184
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_591_6
timestamp 1730592110
transform 1 0 144 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_591_6
timestamp 1730592110
transform 1 0 144 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_590_6
timestamp 1730592110
transform 1 0 200 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_590_6
timestamp 1730592110
transform 1 0 200 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_589_6
timestamp 1730592110
transform 1 0 256 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_589_6
timestamp 1730592110
transform 1 0 256 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_588_6
timestamp 1730592110
transform 1 0 312 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_588_6
timestamp 1730592110
transform 1 0 312 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_587_6
timestamp 1730592110
transform 1 0 368 0 -1 192
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_587_6
timestamp 1730592110
transform 1 0 368 0 -1 192
box 9 2 47 46
use welltap_svt  __well_tap__3
timestamp 1730592110
transform 1 0 768 0 -1 184
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730592110
transform 1 0 768 0 -1 184
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_586_6
timestamp 1730592110
transform 1 0 264 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_586_6
timestamp 1730592110
transform 1 0 264 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_585_6
timestamp 1730592110
transform 1 0 320 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_585_6
timestamp 1730592110
transform 1 0 320 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_584_6
timestamp 1730592110
transform 1 0 376 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_584_6
timestamp 1730592110
transform 1 0 376 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_583_6
timestamp 1730592110
transform 1 0 432 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_583_6
timestamp 1730592110
transform 1 0 432 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_582_6
timestamp 1730592110
transform 1 0 488 0 1 196
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_582_6
timestamp 1730592110
transform 1 0 488 0 1 196
box 9 2 47 46
use welltap_svt  __well_tap__4
timestamp 1730592110
transform 1 0 104 0 1 204
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730592110
transform 1 0 104 0 1 204
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730592110
transform 1 0 768 0 1 204
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730592110
transform 1 0 768 0 1 204
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730592110
transform 1 0 104 0 -1 296
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730592110
transform 1 0 104 0 -1 296
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_581_6
timestamp 1730592110
transform 1 0 200 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_581_6
timestamp 1730592110
transform 1 0 200 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_580_6
timestamp 1730592110
transform 1 0 256 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_580_6
timestamp 1730592110
transform 1 0 256 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_579_6
timestamp 1730592110
transform 1 0 312 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_579_6
timestamp 1730592110
transform 1 0 312 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_578_6
timestamp 1730592110
transform 1 0 368 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_578_6
timestamp 1730592110
transform 1 0 368 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_577_6
timestamp 1730592110
transform 1 0 424 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_577_6
timestamp 1730592110
transform 1 0 424 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_519_6
timestamp 1730592110
transform 1 0 480 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_519_6
timestamp 1730592110
transform 1 0 480 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_518_6
timestamp 1730592110
transform 1 0 536 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_518_6
timestamp 1730592110
transform 1 0 536 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_517_6
timestamp 1730592110
transform 1 0 592 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_517_6
timestamp 1730592110
transform 1 0 592 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_516_6
timestamp 1730592110
transform 1 0 648 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_516_6
timestamp 1730592110
transform 1 0 648 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_515_6
timestamp 1730592110
transform 1 0 704 0 -1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_515_6
timestamp 1730592110
transform 1 0 704 0 -1 304
box 9 2 47 46
use welltap_svt  __well_tap__7
timestamp 1730592110
transform 1 0 768 0 -1 296
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730592110
transform 1 0 768 0 -1 296
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730592110
transform 1 0 104 0 1 312
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730592110
transform 1 0 104 0 1 312
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_576_6
timestamp 1730592110
transform 1 0 272 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_576_6
timestamp 1730592110
transform 1 0 272 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_575_6
timestamp 1730592110
transform 1 0 328 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_575_6
timestamp 1730592110
transform 1 0 328 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_574_6
timestamp 1730592110
transform 1 0 392 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_574_6
timestamp 1730592110
transform 1 0 392 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_573_6
timestamp 1730592110
transform 1 0 456 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_573_6
timestamp 1730592110
transform 1 0 456 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_572_6
timestamp 1730592110
transform 1 0 520 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_572_6
timestamp 1730592110
transform 1 0 520 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_520_6
timestamp 1730592110
transform 1 0 584 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_520_6
timestamp 1730592110
transform 1 0 584 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_513_6
timestamp 1730592110
transform 1 0 648 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_513_6
timestamp 1730592110
transform 1 0 648 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_514_6
timestamp 1730592110
transform 1 0 704 0 1 304
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_514_6
timestamp 1730592110
transform 1 0 704 0 1 304
box 9 2 47 46
use welltap_svt  __well_tap__9
timestamp 1730592110
transform 1 0 768 0 1 312
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730592110
transform 1 0 768 0 1 312
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730592110
transform 1 0 104 0 -1 392
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730592110
transform 1 0 104 0 -1 392
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_567_6
timestamp 1730592110
transform 1 0 128 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_567_6
timestamp 1730592110
transform 1 0 128 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_568_6
timestamp 1730592110
transform 1 0 208 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_568_6
timestamp 1730592110
transform 1 0 208 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_569_6
timestamp 1730592110
transform 1 0 296 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_569_6
timestamp 1730592110
transform 1 0 296 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_570_6
timestamp 1730592110
transform 1 0 392 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_570_6
timestamp 1730592110
transform 1 0 392 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_571_6
timestamp 1730592110
transform 1 0 496 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_571_6
timestamp 1730592110
transform 1 0 496 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_521_6
timestamp 1730592110
transform 1 0 608 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_521_6
timestamp 1730592110
transform 1 0 608 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_512_6
timestamp 1730592110
transform 1 0 704 0 -1 400
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_512_6
timestamp 1730592110
transform 1 0 704 0 -1 400
box 9 2 47 46
use welltap_svt  __well_tap__11
timestamp 1730592110
transform 1 0 768 0 -1 392
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730592110
transform 1 0 768 0 -1 392
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730592110
transform 1 0 104 0 1 416
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730592110
transform 1 0 104 0 1 416
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_566_6
timestamp 1730592110
transform 1 0 128 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_566_6
timestamp 1730592110
transform 1 0 128 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_565_6
timestamp 1730592110
transform 1 0 184 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_565_6
timestamp 1730592110
transform 1 0 184 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_564_6
timestamp 1730592110
transform 1 0 256 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_564_6
timestamp 1730592110
transform 1 0 256 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_563_6
timestamp 1730592110
transform 1 0 344 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_563_6
timestamp 1730592110
transform 1 0 344 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_562_6
timestamp 1730592110
transform 1 0 432 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_562_6
timestamp 1730592110
transform 1 0 432 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_522_6
timestamp 1730592110
transform 1 0 528 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_522_6
timestamp 1730592110
transform 1 0 528 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_510_6
timestamp 1730592110
transform 1 0 624 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_510_6
timestamp 1730592110
transform 1 0 624 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_511_6
timestamp 1730592110
transform 1 0 704 0 1 408
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_511_6
timestamp 1730592110
transform 1 0 704 0 1 408
box 9 2 47 46
use welltap_svt  __well_tap__13
timestamp 1730592110
transform 1 0 768 0 1 416
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730592110
transform 1 0 768 0 1 416
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730592110
transform 1 0 104 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730592110
transform 1 0 104 0 -1 500
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_561_6
timestamp 1730592110
transform 1 0 176 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_561_6
timestamp 1730592110
transform 1 0 176 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_560_6
timestamp 1730592110
transform 1 0 264 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_560_6
timestamp 1730592110
transform 1 0 264 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_559_6
timestamp 1730592110
transform 1 0 360 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_559_6
timestamp 1730592110
transform 1 0 360 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_558_6
timestamp 1730592110
transform 1 0 472 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_558_6
timestamp 1730592110
transform 1 0 472 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_557_6
timestamp 1730592110
transform 1 0 592 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_557_6
timestamp 1730592110
transform 1 0 592 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_59_6
timestamp 1730592110
transform 1 0 704 0 -1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_59_6
timestamp 1730592110
transform 1 0 704 0 -1 508
box 9 2 47 46
use welltap_svt  __well_tap__15
timestamp 1730592110
transform 1 0 768 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730592110
transform 1 0 768 0 -1 500
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730592110
transform 1 0 104 0 1 516
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730592110
transform 1 0 104 0 1 516
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_556_6
timestamp 1730592110
transform 1 0 304 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_556_6
timestamp 1730592110
transform 1 0 304 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_555_6
timestamp 1730592110
transform 1 0 376 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_555_6
timestamp 1730592110
transform 1 0 376 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_554_6
timestamp 1730592110
transform 1 0 456 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_554_6
timestamp 1730592110
transform 1 0 456 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_553_6
timestamp 1730592110
transform 1 0 536 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_553_6
timestamp 1730592110
transform 1 0 536 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_523_6
timestamp 1730592110
transform 1 0 624 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_523_6
timestamp 1730592110
transform 1 0 624 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_58_6
timestamp 1730592110
transform 1 0 704 0 1 508
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_58_6
timestamp 1730592110
transform 1 0 704 0 1 508
box 9 2 47 46
use welltap_svt  __well_tap__17
timestamp 1730592110
transform 1 0 768 0 1 516
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730592110
transform 1 0 768 0 1 516
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_549_6
timestamp 1730592110
transform 1 0 328 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_549_6
timestamp 1730592110
transform 1 0 328 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_550_6
timestamp 1730592110
transform 1 0 392 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_550_6
timestamp 1730592110
transform 1 0 392 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_551_6
timestamp 1730592110
transform 1 0 464 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_551_6
timestamp 1730592110
transform 1 0 464 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_552_6
timestamp 1730592110
transform 1 0 544 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_552_6
timestamp 1730592110
transform 1 0 544 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_524_6
timestamp 1730592110
transform 1 0 632 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_524_6
timestamp 1730592110
transform 1 0 632 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_57_6
timestamp 1730592110
transform 1 0 704 0 -1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_57_6
timestamp 1730592110
transform 1 0 704 0 -1 604
box 9 2 47 46
use welltap_svt  __well_tap__18
timestamp 1730592110
transform 1 0 104 0 -1 596
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730592110
transform 1 0 104 0 -1 596
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_548_6
timestamp 1730592110
transform 1 0 264 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_548_6
timestamp 1730592110
transform 1 0 264 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_547_6
timestamp 1730592110
transform 1 0 320 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_547_6
timestamp 1730592110
transform 1 0 320 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_546_6
timestamp 1730592110
transform 1 0 384 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_546_6
timestamp 1730592110
transform 1 0 384 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_545_6
timestamp 1730592110
transform 1 0 456 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_545_6
timestamp 1730592110
transform 1 0 456 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_526_6
timestamp 1730592110
transform 1 0 536 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_526_6
timestamp 1730592110
transform 1 0 536 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_525_6
timestamp 1730592110
transform 1 0 624 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_525_6
timestamp 1730592110
transform 1 0 624 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_56_6
timestamp 1730592110
transform 1 0 704 0 1 604
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_56_6
timestamp 1730592110
transform 1 0 704 0 1 604
box 9 2 47 46
use welltap_svt  __well_tap__19
timestamp 1730592110
transform 1 0 768 0 -1 596
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730592110
transform 1 0 768 0 -1 596
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730592110
transform 1 0 104 0 1 612
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730592110
transform 1 0 104 0 1 612
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730592110
transform 1 0 768 0 1 612
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730592110
transform 1 0 768 0 1 612
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730592110
transform 1 0 104 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730592110
transform 1 0 104 0 -1 696
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_542_6
timestamp 1730592110
transform 1 0 208 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_542_6
timestamp 1730592110
transform 1 0 208 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_543_6
timestamp 1730592110
transform 1 0 312 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_543_6
timestamp 1730592110
transform 1 0 312 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_544_6
timestamp 1730592110
transform 1 0 416 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_544_6
timestamp 1730592110
transform 1 0 416 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_527_6
timestamp 1730592110
transform 1 0 520 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_527_6
timestamp 1730592110
transform 1 0 520 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_54_6
timestamp 1730592110
transform 1 0 624 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_54_6
timestamp 1730592110
transform 1 0 624 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_55_6
timestamp 1730592110
transform 1 0 704 0 -1 704
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_55_6
timestamp 1730592110
transform 1 0 704 0 -1 704
box 9 2 47 46
use welltap_svt  __well_tap__23
timestamp 1730592110
transform 1 0 768 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730592110
transform 1 0 768 0 -1 696
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730592110
transform 1 0 104 0 1 720
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730592110
transform 1 0 104 0 1 720
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_541_6
timestamp 1730592110
transform 1 0 160 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_541_6
timestamp 1730592110
transform 1 0 160 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_540_6
timestamp 1730592110
transform 1 0 224 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_540_6
timestamp 1730592110
transform 1 0 224 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_539_6
timestamp 1730592110
transform 1 0 296 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_539_6
timestamp 1730592110
transform 1 0 296 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_538_6
timestamp 1730592110
transform 1 0 376 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_538_6
timestamp 1730592110
transform 1 0 376 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_528_6
timestamp 1730592110
transform 1 0 464 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_528_6
timestamp 1730592110
transform 1 0 464 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_529_6
timestamp 1730592110
transform 1 0 552 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_529_6
timestamp 1730592110
transform 1 0 552 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_53_6
timestamp 1730592110
transform 1 0 640 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_53_6
timestamp 1730592110
transform 1 0 640 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_52_6
timestamp 1730592110
transform 1 0 704 0 1 712
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_52_6
timestamp 1730592110
transform 1 0 704 0 1 712
box 9 2 47 46
use welltap_svt  __well_tap__25
timestamp 1730592110
transform 1 0 768 0 1 720
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730592110
transform 1 0 768 0 1 720
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730592110
transform 1 0 104 0 -1 808
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730592110
transform 1 0 104 0 -1 808
box 8 4 12 24
use _0_0std_0_0cells_0_0NOR2X1  nor_537_6
timestamp 1730592110
transform 1 0 176 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_537_6
timestamp 1730592110
transform 1 0 176 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_536_6
timestamp 1730592110
transform 1 0 232 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_536_6
timestamp 1730592110
transform 1 0 232 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_535_6
timestamp 1730592110
transform 1 0 288 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_535_6
timestamp 1730592110
transform 1 0 288 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_534_6
timestamp 1730592110
transform 1 0 344 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_534_6
timestamp 1730592110
transform 1 0 344 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_533_6
timestamp 1730592110
transform 1 0 400 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_533_6
timestamp 1730592110
transform 1 0 400 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_532_6
timestamp 1730592110
transform 1 0 456 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_532_6
timestamp 1730592110
transform 1 0 456 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_531_6
timestamp 1730592110
transform 1 0 520 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_531_6
timestamp 1730592110
transform 1 0 520 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_530_6
timestamp 1730592110
transform 1 0 584 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_530_6
timestamp 1730592110
transform 1 0 584 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_50_6
timestamp 1730592110
transform 1 0 648 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_50_6
timestamp 1730592110
transform 1 0 648 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_51_6
timestamp 1730592110
transform 1 0 704 0 -1 816
box 9 2 47 46
use _0_0std_0_0cells_0_0NOR2X1  nor_51_6
timestamp 1730592110
transform 1 0 704 0 -1 816
box 9 2 47 46
use welltap_svt  __well_tap__27
timestamp 1730592110
transform 1 0 768 0 -1 808
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730592110
transform 1 0 768 0 -1 808
box 8 4 12 24
<< end >>
